* NGSPICE file created from opamp_corec.ext - technology: sky130A

.subckt opamp_corec gp dp out dn gn xn vdda vssa
X0 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X1 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X2 n2 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X3 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X4 n7 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X5 p7 gp vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X6 vdda gp p8 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X7 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X8 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X9 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X10 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X11 xn gn n7 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X12 p1 gp vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X13 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X14 xn gn n5 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X15 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X16 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X17 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X18 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X19 n6 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X20 xp gp p3 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X21 p2 gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X22 p8 gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X23 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X24 n1 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X25 n4 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X26 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X27 p5 gp vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X28 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X29 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X30 xp gp p1 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X31 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X32 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X33 vssa gn n2 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X34 vssa gn n6 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X35 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X36 vssa gn n4 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X37 p3 gp vdda vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.95e+12p ps=5.05e+06u w=3e+06u l=2e+06u
X38 vdda gp p6 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X39 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X40 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X41 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X42 n5 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X43 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X44 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X45 n3 gn vssa vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.5e+11p ps=2.55e+06u w=1e+06u l=2e+06u
X46 vdda gp p2 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X47 p6 gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X48 vdda gp p4 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.95e+12p pd=5.05e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X49 dn gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.25e+11p pd=2.375e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X50 n8 gn xn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X51 xn gn n3 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X52 p4 gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X53 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X54 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X55 vssa gn n8 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6.5e+11p pd=2.55e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
X56 xp gp p7 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X57 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X58 xn gn dn vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6.25e+11p ps=2.375e+06u w=1e+06u l=2e+06u
X59 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X60 xp gp p5 vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X61 xp gp dp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.85e+12p pd=4.48333e+06u as=1.8e+12p ps=4.2e+06u w=3e+06u l=2e+06u
X62 dp gp xp vdda sky130_fd_pr__pfet_g5v0d10v5 ad=1.8e+12p pd=4.2e+06u as=1.85e+12p ps=4.48333e+06u w=3e+06u l=2e+06u
X63 xn gn n1 vssa sky130_fd_pr__nfet_g5v0d10v5 ad=6e+11p pd=2.2e+06u as=6e+11p ps=2.2e+06u w=1e+06u l=2e+06u
.ends

