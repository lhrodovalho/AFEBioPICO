magic
tech sky130A
timestamp 1634672824
<< nwell >>
rect -2870 -3290 -2820 -460
rect 23500 -3290 23550 -460
<< pwell >>
rect -2910 -440 -2820 -410
rect 23500 -440 23590 -410
rect -2920 -5150 -2810 -5120
rect 23500 -5150 23600 -5120
rect -2920 -6280 -2890 -5150
rect 23570 -6280 23600 -5150
<< psubdiff >>
rect -2920 -440 -2820 -410
rect 23500 -440 23600 -410
rect -2920 -3310 -2890 -440
rect 23570 -3310 23600 -440
rect -2920 -3340 -1810 -3310
rect 10270 -3340 10410 -3310
rect 22490 -3340 23600 -3310
rect -2920 -5120 -2890 -3340
rect 23570 -5120 23600 -3340
rect -2920 -5150 -2810 -5120
rect 23500 -5150 23600 -5120
rect -2920 -6280 -2890 -5150
rect 23570 -6280 23600 -5150
rect -2920 -6310 23600 -6280
<< psubdiffcont >>
rect -1810 -3340 10270 -3310
rect 10410 -3340 22490 -3310
<< locali >>
rect -6280 -4120 -6110 -220
rect -6080 -4120 -5910 -220
rect -5880 -4120 -5710 -220
rect -5680 -4120 -5510 -220
rect -5480 -4120 -5310 -220
rect -5280 -4120 -5110 -220
rect -5080 -4120 -4710 -220
rect -4680 -4120 -4510 -220
rect -4480 -4120 -4310 -220
rect -4280 -4120 -4110 -220
rect -4080 -4120 -3910 -220
rect -3880 -4120 -3710 -220
rect -3680 -3400 -3510 -220
rect -2920 -440 -2820 -410
rect 23500 -440 23600 -410
rect -2920 -3310 -2890 -440
rect -1010 -480 -960 -470
rect -2850 -3270 -2820 -480
rect -1010 -510 -1000 -480
rect -970 -510 -960 -480
rect -1010 -520 -960 -510
rect 21640 -480 21690 -470
rect 21640 -510 21650 -480
rect 21680 -510 21690 -480
rect 21640 -520 21690 -510
rect 23500 -3270 23530 -480
rect 23570 -3310 23600 -440
rect -2920 -3340 -1850 -3310
rect -1820 -3340 -1810 -3310
rect 10270 -3340 10410 -3310
rect 22490 -3340 22500 -3310
rect 22530 -3340 23600 -3310
rect -3680 -3490 23560 -3400
rect -3680 -3520 -3510 -3490
rect -3680 -3610 23560 -3520
rect -3680 -3640 -3510 -3610
rect -3680 -3730 23560 -3640
rect -3680 -3760 -3510 -3730
rect -3680 -3850 23560 -3760
rect -3680 -3880 -3510 -3850
rect -3680 -3970 23560 -3880
rect -3680 -4000 -3510 -3970
rect -3680 -4090 23560 -4000
rect -3680 -4120 -3510 -4090
rect -6280 -4160 24420 -4120
rect -6280 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect -6280 -4340 24420 -4300
rect -6280 -6500 -6110 -4340
rect -6080 -6500 -5910 -4340
rect -5880 -6500 -5710 -4340
rect -5680 -6500 -5510 -4340
rect -5480 -6500 -5310 -4340
rect -5280 -6500 -5110 -4340
rect -5080 -6500 -4710 -4340
rect -4680 -6500 -4510 -4340
rect -4480 -6500 -4310 -4340
rect -4280 -6500 -4110 -4340
rect -4080 -6500 -3910 -4340
rect -3880 -6500 -3710 -4340
rect -3680 -4370 -3510 -4340
rect -3680 -4460 23560 -4370
rect -3680 -4490 -3510 -4460
rect -3680 -4580 23560 -4490
rect -3680 -4610 -3510 -4580
rect -3680 -4700 23560 -4610
rect -3680 -4730 -3510 -4700
rect -3680 -4820 23560 -4730
rect -3680 -4850 -3510 -4820
rect -3680 -4940 23560 -4850
rect -3680 -4970 -3510 -4940
rect -3680 -5060 23560 -4970
rect -3680 -6500 -3510 -5060
rect -2920 -5150 -2810 -5120
rect 23500 -5150 23600 -5120
rect -2920 -6280 -2890 -5150
rect -1860 -6280 -1810 -6270
rect 22490 -6280 22540 -6270
rect 23570 -6280 23600 -5150
rect -2920 -6310 -1850 -6280
rect -1820 -6310 22500 -6280
rect 22530 -6310 23600 -6280
rect -1860 -6320 -1810 -6310
rect 22490 -6320 22540 -6310
<< viali >>
rect -1000 -510 -970 -480
rect 21650 -510 21680 -480
rect -1850 -3340 -1820 -3310
rect 22500 -3340 22530 -3310
rect 24270 -4300 24410 -4160
rect -1850 -6310 -1820 -6280
rect 22500 -6310 22530 -6280
<< metal1 >>
rect -6310 -3360 -6280 -220
rect -6110 -3360 -6080 -220
rect -5910 -3360 -5880 -220
rect -5710 -3360 -5680 -220
rect -5510 -3360 -5480 -220
rect -5310 -3360 -5280 -220
rect -5110 -3360 -5080 -220
rect -4710 -3360 -4680 -220
rect -4510 -3360 -4480 -220
rect -4310 -3360 -4280 -220
rect -4110 -3360 -4080 -220
rect -3910 -3360 -3880 -220
rect -3710 -3360 -3680 -220
rect -3510 -3360 -3480 -220
rect -2790 -230 -2760 -220
rect -2790 -3360 -2760 -370
rect -1940 -230 -1910 -220
rect -1940 -390 -1910 -370
rect -1000 -230 -970 -220
rect -1000 -390 -970 -370
rect 880 -230 910 -220
rect 880 -450 910 -370
rect 1820 -230 1850 -220
rect 1820 -450 1850 -370
rect 3700 -230 3730 -220
rect 3700 -390 3730 -370
rect 5580 -230 5610 -220
rect 5580 -390 5610 -370
rect 7460 -230 7490 -220
rect 7460 -390 7490 -370
rect 10280 -230 10310 -220
rect 10280 -390 10310 -370
rect 10370 -230 10400 -220
rect 10370 -390 10400 -370
rect 13190 -230 13220 -220
rect 13190 -390 13220 -370
rect 15070 -230 15100 -220
rect 15070 -390 15100 -370
rect 16950 -230 16980 -220
rect 16950 -390 16980 -370
rect 18830 -230 18860 -220
rect 18830 -450 18860 -370
rect 19770 -230 19800 -220
rect 19770 -450 19800 -370
rect 21650 -230 21680 -220
rect 21650 -390 21680 -370
rect 22590 -230 22620 -220
rect 22590 -390 22620 -370
rect 23440 -230 23470 -220
rect -1010 -480 -960 -470
rect -1010 -510 -1000 -480
rect -970 -510 -960 -480
rect -1010 -520 -960 -510
rect 21640 -480 21690 -470
rect 21640 -510 21650 -480
rect 21680 -510 21690 -480
rect 21640 -520 21690 -510
rect 23440 -540 23470 -370
rect -1860 -3310 -1810 -3300
rect -1860 -3340 -1850 -3310
rect -1820 -3340 -1810 -3310
rect -1860 -3350 -1810 -3340
rect -6320 -3370 -6270 -3360
rect -6320 -3400 -6310 -3370
rect -6280 -3400 -6270 -3370
rect -6320 -3410 -6270 -3400
rect -6120 -3370 -6070 -3360
rect -6120 -3400 -6110 -3370
rect -6080 -3400 -6070 -3370
rect -6120 -3410 -6070 -3400
rect -5920 -3370 -5870 -3360
rect -5920 -3400 -5910 -3370
rect -5880 -3400 -5870 -3370
rect -5920 -3410 -5870 -3400
rect -5720 -3370 -5670 -3360
rect -5720 -3400 -5710 -3370
rect -5680 -3400 -5670 -3370
rect -5720 -3410 -5670 -3400
rect -5520 -3370 -5470 -3360
rect -5520 -3400 -5510 -3370
rect -5480 -3400 -5470 -3370
rect -5520 -3410 -5470 -3400
rect -5320 -3370 -5270 -3360
rect -5320 -3400 -5310 -3370
rect -5280 -3400 -5270 -3370
rect -5320 -3410 -5270 -3400
rect -5120 -3370 -5070 -3360
rect -5120 -3400 -5110 -3370
rect -5080 -3400 -5070 -3370
rect -5120 -3410 -5070 -3400
rect -4720 -3370 -4670 -3360
rect -4720 -3400 -4710 -3370
rect -4680 -3400 -4670 -3370
rect -4720 -3410 -4670 -3400
rect -4520 -3370 -4470 -3360
rect -4520 -3400 -4510 -3370
rect -4480 -3400 -4470 -3370
rect -4520 -3410 -4470 -3400
rect -4320 -3370 -4270 -3360
rect -4320 -3400 -4310 -3370
rect -4280 -3400 -4270 -3370
rect -4320 -3410 -4270 -3400
rect -4120 -3370 -4070 -3360
rect -4120 -3400 -4110 -3370
rect -4080 -3400 -4070 -3370
rect -4120 -3410 -4070 -3400
rect -3920 -3370 -3870 -3360
rect -3920 -3400 -3910 -3370
rect -3880 -3400 -3870 -3370
rect -3920 -3410 -3870 -3400
rect -3720 -3370 -3670 -3360
rect -3720 -3400 -3710 -3370
rect -3680 -3400 -3670 -3370
rect -3720 -3410 -3670 -3400
rect -3520 -3370 -3470 -3360
rect -3520 -3400 -3510 -3370
rect -3480 -3400 -3470 -3370
rect -3520 -3410 -3470 -3400
rect -6310 -3480 -6280 -3410
rect -6320 -3490 -6270 -3480
rect -6320 -3520 -6310 -3490
rect -6280 -3520 -6270 -3490
rect -6320 -3530 -6270 -3520
rect -6310 -3600 -6280 -3530
rect -6320 -3610 -6270 -3600
rect -6320 -3640 -6310 -3610
rect -6280 -3640 -6270 -3610
rect -6320 -3650 -6270 -3640
rect -6310 -3720 -6280 -3650
rect -6320 -3730 -6270 -3720
rect -6320 -3760 -6310 -3730
rect -6280 -3760 -6270 -3730
rect -6320 -3770 -6270 -3760
rect -6310 -3840 -6280 -3770
rect -6320 -3850 -6270 -3840
rect -6320 -3880 -6310 -3850
rect -6280 -3880 -6270 -3850
rect -6320 -3890 -6270 -3880
rect -6310 -3960 -6280 -3890
rect -6320 -3970 -6270 -3960
rect -6320 -4000 -6310 -3970
rect -6280 -4000 -6270 -3970
rect -6320 -4010 -6270 -4000
rect -6310 -4080 -6280 -4010
rect -6320 -4090 -6270 -4080
rect -6320 -4120 -6310 -4090
rect -6280 -4120 -6270 -4090
rect -6320 -4130 -6270 -4120
rect -6310 -4330 -6280 -4130
rect -6320 -4340 -6270 -4330
rect -6320 -4370 -6310 -4340
rect -6280 -4370 -6270 -4340
rect -6320 -4380 -6270 -4370
rect -6310 -4450 -6280 -4380
rect -6320 -4460 -6270 -4450
rect -6320 -4490 -6310 -4460
rect -6280 -4490 -6270 -4460
rect -6320 -4500 -6270 -4490
rect -6310 -4570 -6280 -4500
rect -6320 -4580 -6270 -4570
rect -6320 -4610 -6310 -4580
rect -6280 -4610 -6270 -4580
rect -6320 -4620 -6270 -4610
rect -6310 -4690 -6280 -4620
rect -6320 -4700 -6270 -4690
rect -6320 -4730 -6310 -4700
rect -6280 -4730 -6270 -4700
rect -6320 -4740 -6270 -4730
rect -6310 -4810 -6280 -4740
rect -6320 -4820 -6270 -4810
rect -6320 -4850 -6310 -4820
rect -6280 -4850 -6270 -4820
rect -6320 -4860 -6270 -4850
rect -6310 -4930 -6280 -4860
rect -6320 -4940 -6270 -4930
rect -6320 -4970 -6310 -4940
rect -6280 -4970 -6270 -4940
rect -6320 -4980 -6270 -4970
rect -6310 -5050 -6280 -4980
rect -6110 -5050 -6080 -3410
rect -5910 -5050 -5880 -3410
rect -5710 -5050 -5680 -3410
rect -5510 -5050 -5480 -3410
rect -5310 -5050 -5280 -3410
rect -5110 -5050 -5080 -3410
rect -4710 -5050 -4680 -3410
rect -4510 -5050 -4480 -3410
rect -4310 -5050 -4280 -3410
rect -4110 -5050 -4080 -3410
rect -3910 -5050 -3880 -3410
rect -3710 -5050 -3680 -3410
rect -3510 -5050 -3480 -3410
rect -2670 -3430 -2640 -3360
rect -2670 -3470 -2640 -3460
rect -2060 -5000 -2030 -4990
rect -6400 -5060 -6350 -5050
rect -6400 -5090 -6390 -5060
rect -6360 -5090 -6350 -5060
rect -6400 -5100 -6350 -5090
rect -6320 -5060 -6270 -5050
rect -6320 -5090 -6310 -5060
rect -6280 -5090 -6270 -5060
rect -6320 -5100 -6270 -5090
rect -6120 -5060 -6070 -5050
rect -6120 -5090 -6110 -5060
rect -6080 -5090 -6070 -5060
rect -6120 -5100 -6070 -5090
rect -5920 -5060 -5870 -5050
rect -5920 -5090 -5910 -5060
rect -5880 -5090 -5870 -5060
rect -5920 -5100 -5870 -5090
rect -5720 -5060 -5670 -5050
rect -5720 -5090 -5710 -5060
rect -5680 -5090 -5670 -5060
rect -5720 -5100 -5670 -5090
rect -5520 -5060 -5470 -5050
rect -5520 -5090 -5510 -5060
rect -5480 -5090 -5470 -5060
rect -5520 -5100 -5470 -5090
rect -5320 -5060 -5270 -5050
rect -5320 -5090 -5310 -5060
rect -5280 -5090 -5270 -5060
rect -5320 -5100 -5270 -5090
rect -5120 -5060 -5070 -5050
rect -5120 -5090 -5110 -5060
rect -5080 -5090 -5070 -5060
rect -5120 -5100 -5070 -5090
rect -4720 -5060 -4670 -5050
rect -4720 -5090 -4710 -5060
rect -4680 -5090 -4670 -5060
rect -4720 -5100 -4670 -5090
rect -4520 -5060 -4470 -5050
rect -4520 -5090 -4510 -5060
rect -4480 -5090 -4470 -5060
rect -4520 -5100 -4470 -5090
rect -4320 -5060 -4270 -5050
rect -4320 -5090 -4310 -5060
rect -4280 -5090 -4270 -5060
rect -4320 -5100 -4270 -5090
rect -4120 -5060 -4070 -5050
rect -4120 -5090 -4110 -5060
rect -4080 -5090 -4070 -5060
rect -4120 -5100 -4070 -5090
rect -3920 -5060 -3870 -5050
rect -3920 -5090 -3910 -5060
rect -3880 -5090 -3870 -5060
rect -3920 -5100 -3870 -5090
rect -3720 -5060 -3670 -5050
rect -3720 -5090 -3710 -5060
rect -3680 -5090 -3670 -5060
rect -3720 -5100 -3670 -5090
rect -3520 -5060 -3470 -5050
rect -3520 -5090 -3510 -5060
rect -3480 -5090 -3470 -5060
rect -3520 -5100 -3470 -5090
rect -6310 -6500 -6280 -5100
rect -6110 -6500 -6080 -5100
rect -5910 -6500 -5880 -5100
rect -5710 -6500 -5680 -5100
rect -5510 -6500 -5480 -5100
rect -5310 -6500 -5280 -5100
rect -5110 -6500 -5080 -5100
rect -4710 -6500 -4680 -5100
rect -4510 -6500 -4480 -5100
rect -4310 -6500 -4280 -5100
rect -4110 -6500 -4080 -5100
rect -3910 -6500 -3880 -5100
rect -3710 -6500 -3680 -5100
rect -3510 -6500 -3480 -5100
rect -2790 -6350 -2760 -5100
rect -2060 -5110 -2030 -5030
rect -2790 -6500 -2760 -6490
rect -1940 -6350 -1910 -5100
rect -1850 -6270 -1820 -3350
rect -1730 -3430 -1700 -3360
rect -1730 -3470 -1700 -3460
rect -1000 -3430 -970 -3360
rect -1000 -3470 -970 -3460
rect -910 -3550 -880 -3360
rect -910 -3590 -880 -3580
rect -790 -3550 -760 -3360
rect -60 -3430 -30 -3150
rect 1820 -3160 1850 -3150
rect -60 -3470 -30 -3460
rect 150 -3430 180 -3360
rect 150 -3470 180 -3460
rect -790 -3590 -760 -3580
rect 760 -4880 790 -4870
rect -1120 -5000 -1090 -4990
rect -1120 -5100 -1090 -5030
rect -910 -5000 -880 -4990
rect -910 -5100 -880 -5030
rect -180 -5000 -150 -4990
rect -180 -5100 -150 -5030
rect 30 -5000 60 -4990
rect 30 -5240 60 -5030
rect 760 -5100 790 -4910
rect 880 -4880 910 -3360
rect 1090 -3430 1120 -3360
rect 1090 -3470 1120 -3460
rect 1820 -3670 1850 -3360
rect 1820 -3710 1850 -3700
rect 1910 -3670 1940 -3360
rect 1910 -3710 1940 -3700
rect 2030 -3790 2060 -3360
rect 2030 -3830 2060 -3820
rect 880 -5100 910 -4910
rect 970 -4030 1000 -4020
rect 970 -5100 1000 -4060
rect 1910 -4030 1940 -4020
rect 1700 -4520 1730 -4510
rect 1700 -5100 1730 -4550
rect 1910 -5240 1940 -4060
rect 2760 -4030 2790 -3150
rect 2970 -3430 3000 -3360
rect 2970 -3470 3000 -3460
rect 3700 -3670 3730 -3360
rect 3700 -3710 3730 -3700
rect 3790 -3670 3820 -3360
rect 3790 -3710 3820 -3700
rect 3910 -3910 3940 -3350
rect 3910 -3950 3940 -3940
rect 2760 -4070 2790 -4060
rect 2850 -4400 2880 -4390
rect 2640 -4520 2670 -4510
rect 2640 -5100 2670 -4550
rect 2760 -4520 2790 -4510
rect 2760 -5100 2790 -4550
rect 2850 -5100 2880 -4430
rect 3790 -4400 3820 -4390
rect 3580 -4520 3610 -4510
rect 3580 -5100 3610 -4550
rect 3790 -5240 3820 -4430
rect 4640 -4400 4670 -3150
rect 4850 -3430 4880 -3360
rect 4850 -3470 4880 -3460
rect 4640 -4440 4670 -4430
rect 4730 -4400 4760 -4390
rect 4520 -4520 4550 -4510
rect 4520 -5100 4550 -4550
rect 4640 -4760 4670 -4750
rect 4640 -5100 4670 -4790
rect 4730 -5100 4760 -4430
rect 5460 -4520 5490 -4510
rect 5460 -5100 5490 -4550
rect 5580 -4520 5610 -3360
rect 5670 -3670 5700 -3360
rect 5670 -3710 5700 -3700
rect 5790 -3910 5820 -3360
rect 5790 -3950 5820 -3940
rect 5580 -4560 5610 -4550
rect 5670 -4400 5700 -4390
rect 5670 -5240 5700 -4430
rect 6520 -4400 6550 -3150
rect 6730 -3430 6760 -3360
rect 6730 -3470 6760 -3460
rect 6520 -4440 6550 -4430
rect 6610 -4030 6640 -4020
rect 6400 -4520 6430 -4510
rect 6400 -5100 6430 -4550
rect 6520 -4760 6550 -4750
rect 6520 -5100 6550 -4790
rect 6610 -5100 6640 -4060
rect 7340 -4520 7370 -4510
rect 7340 -5100 7370 -4550
rect 7460 -4640 7490 -3360
rect 7550 -3670 7580 -3360
rect 7550 -3710 7580 -3700
rect 7670 -3790 7700 -3360
rect 7670 -3830 7700 -3820
rect 7460 -4680 7490 -4670
rect 7550 -4030 7580 -4020
rect 7550 -5240 7580 -4060
rect 8400 -4030 8430 -3150
rect 8400 -4070 8430 -4060
rect 8280 -4520 8310 -4510
rect 8280 -5100 8310 -4550
rect 8400 -4520 8430 -4510
rect 8400 -5100 8430 -4550
rect 8490 -4640 8520 -3360
rect 8610 -3550 8640 -3360
rect 8610 -3590 8640 -3580
rect 8490 -5240 8520 -4670
rect 9340 -4760 9370 -3150
rect 9220 -4880 9250 -4870
rect 9220 -5100 9250 -4910
rect 9340 -5100 9370 -4790
rect 9430 -4160 9460 -4150
rect 9430 -5100 9460 -4300
rect 9550 -4640 9580 -3350
rect 10280 -4160 10310 -2570
rect 10280 -4310 10310 -4300
rect 10370 -4160 10400 -3360
rect 10370 -4310 10400 -4300
rect 9550 -4680 9580 -4670
rect 11100 -4640 11130 -3360
rect 11100 -4680 11130 -4670
rect 11220 -4160 11250 -4150
rect 10160 -4760 10190 -4750
rect 10160 -5100 10190 -4790
rect 10490 -4760 10520 -4750
rect 10490 -5100 10520 -4790
rect 11220 -5100 11250 -4300
rect 11310 -4760 11340 -3150
rect 12040 -3550 12070 -3360
rect 12040 -3590 12070 -3580
rect 11310 -5100 11340 -4790
rect 12160 -4640 12190 -3360
rect 12250 -4030 12280 -3150
rect 12980 -3790 13010 -3360
rect 13100 -3670 13130 -3360
rect 13100 -3710 13130 -3700
rect 12980 -3830 13010 -3820
rect 12250 -4070 12280 -4060
rect 13100 -4030 13130 -4020
rect 11430 -4880 11460 -4870
rect 11430 -5100 11460 -4910
rect 12160 -5240 12190 -4670
rect 12250 -4520 12280 -4510
rect 12250 -5100 12280 -4550
rect 12370 -4520 12400 -4510
rect 12370 -5100 12400 -4550
rect 13100 -5240 13130 -4060
rect 13190 -4640 13220 -3360
rect 13920 -3430 13950 -3360
rect 13920 -3470 13950 -3460
rect 14040 -4030 14070 -4020
rect 13190 -4680 13220 -4670
rect 13310 -4520 13340 -4510
rect 13310 -5100 13340 -4550
rect 14040 -5100 14070 -4060
rect 14130 -4400 14160 -3150
rect 14860 -3910 14890 -3360
rect 14980 -3670 15010 -3360
rect 14980 -3710 15010 -3700
rect 14860 -3950 14890 -3940
rect 14130 -4440 14160 -4430
rect 14980 -4400 15010 -4390
rect 14250 -4520 14280 -4510
rect 14130 -4760 14160 -4750
rect 14130 -5100 14160 -4790
rect 14250 -5100 14280 -4550
rect 14980 -5240 15010 -4430
rect 15070 -4520 15100 -3360
rect 15800 -3430 15830 -3360
rect 15800 -3470 15830 -3460
rect 15920 -4400 15950 -4390
rect 15070 -4560 15100 -4550
rect 15190 -4520 15220 -4510
rect 15190 -5100 15220 -4550
rect 15920 -5100 15950 -4430
rect 16010 -4400 16040 -3150
rect 16740 -3910 16770 -3350
rect 16860 -3670 16890 -3360
rect 16860 -3710 16890 -3700
rect 16950 -3670 16980 -3360
rect 17680 -3430 17710 -3360
rect 17680 -3470 17710 -3460
rect 16950 -3710 16980 -3700
rect 16740 -3950 16770 -3940
rect 17890 -4030 17920 -3150
rect 18830 -3160 18860 -3150
rect 18620 -3790 18650 -3360
rect 18740 -3670 18770 -3360
rect 18740 -3710 18770 -3700
rect 18830 -3670 18860 -3360
rect 19560 -3430 19590 -3360
rect 19560 -3470 19590 -3460
rect 18830 -3710 18860 -3700
rect 18620 -3830 18650 -3820
rect 17890 -4070 17920 -4060
rect 18740 -4030 18770 -4020
rect 16010 -4440 16040 -4430
rect 16860 -4400 16890 -4390
rect 16130 -4520 16160 -4510
rect 16010 -4760 16040 -4750
rect 16010 -5100 16040 -4790
rect 16130 -5100 16160 -4550
rect 16860 -5240 16890 -4430
rect 17800 -4400 17830 -4390
rect 17070 -4520 17100 -4510
rect 17070 -5100 17100 -4550
rect 17800 -5100 17830 -4430
rect 17890 -4520 17920 -4510
rect 17890 -5100 17920 -4550
rect 18010 -4520 18040 -4510
rect 18010 -5100 18040 -4550
rect 18740 -5240 18770 -4060
rect 19680 -4030 19710 -4020
rect 18950 -4520 18980 -4510
rect 18950 -5100 18980 -4550
rect 19680 -5100 19710 -4060
rect 19770 -4880 19800 -3360
rect 20500 -3430 20530 -3360
rect 20500 -3470 20530 -3460
rect 20710 -3430 20740 -3150
rect 22490 -3310 22540 -3300
rect 22490 -3340 22500 -3310
rect 22530 -3340 22540 -3310
rect 22490 -3350 22540 -3340
rect 20710 -3470 20740 -3460
rect 21440 -3550 21470 -3360
rect 21440 -3590 21470 -3580
rect 21560 -3550 21590 -3360
rect 21650 -3430 21680 -3360
rect 21650 -3470 21680 -3460
rect 22380 -3430 22410 -3360
rect 22380 -3470 22410 -3460
rect 21560 -3590 21590 -3580
rect 19770 -5100 19800 -4910
rect 19890 -4880 19920 -4870
rect 19890 -5100 19920 -4910
rect 20620 -5000 20650 -4990
rect 20620 -5240 20650 -5030
rect 20830 -5000 20860 -4990
rect 20830 -5100 20860 -5030
rect 21560 -5000 21590 -4990
rect 21560 -5100 21590 -5030
rect 21770 -5000 21800 -4990
rect 21770 -5100 21800 -5030
rect 22500 -6270 22530 -3350
rect 23320 -3430 23350 -3330
rect 23320 -3470 23350 -3460
rect 24260 -4160 24420 -4150
rect 24260 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect 24260 -4310 24420 -4300
rect 22710 -5000 22740 -4990
rect 22710 -5100 22740 -5030
rect -1860 -6280 -1810 -6270
rect -1860 -6310 -1850 -6280
rect -1820 -6310 -1810 -6280
rect -1860 -6320 -1810 -6310
rect 22490 -6280 22540 -6270
rect 22490 -6310 22500 -6280
rect 22530 -6310 22540 -6280
rect 22490 -6320 22540 -6310
rect -1940 -6500 -1910 -6490
rect -1850 -6350 -1820 -6320
rect -1850 -6500 -1820 -6490
rect -910 -6350 -880 -6330
rect -910 -6500 -880 -6490
rect 970 -6350 1000 -6330
rect 970 -6500 1000 -6490
rect 2850 -6350 2880 -6330
rect 2850 -6500 2880 -6490
rect 4730 -6350 4760 -6330
rect 4730 -6500 4760 -6490
rect 6610 -6350 6640 -6330
rect 6610 -6500 6640 -6490
rect 9430 -6350 9460 -6330
rect 9430 -6500 9460 -6490
rect 11220 -6350 11250 -6330
rect 11220 -6500 11250 -6490
rect 14040 -6350 14070 -6330
rect 14040 -6500 14070 -6490
rect 15920 -6350 15950 -6330
rect 15920 -6500 15950 -6490
rect 17800 -6350 17830 -6330
rect 17800 -6500 17830 -6490
rect 19680 -6350 19710 -6330
rect 19680 -6500 19710 -6490
rect 21560 -6350 21590 -6330
rect 21560 -6500 21590 -6490
rect 22500 -6350 22530 -6320
rect 22500 -6500 22530 -6490
rect 22590 -6350 22620 -6250
rect 22590 -6500 22620 -6490
rect 23440 -6350 23470 -6330
rect 23440 -6500 23470 -6490
<< via1 >>
rect -2790 -370 -2760 -230
rect -1940 -370 -1910 -230
rect -1000 -370 -970 -230
rect 880 -370 910 -230
rect 1820 -370 1850 -230
rect 3700 -370 3730 -230
rect 5580 -370 5610 -230
rect 7460 -370 7490 -230
rect 10280 -370 10310 -230
rect 10370 -370 10400 -230
rect 13190 -370 13220 -230
rect 15070 -370 15100 -230
rect 16950 -370 16980 -230
rect 18830 -370 18860 -230
rect 19770 -370 19800 -230
rect 21650 -370 21680 -230
rect 22590 -370 22620 -230
rect 23440 -370 23470 -230
rect -6310 -3400 -6280 -3370
rect -6110 -3400 -6080 -3370
rect -5910 -3400 -5880 -3370
rect -5710 -3400 -5680 -3370
rect -5510 -3400 -5480 -3370
rect -5310 -3400 -5280 -3370
rect -5110 -3400 -5080 -3370
rect -4710 -3400 -4680 -3370
rect -4510 -3400 -4480 -3370
rect -4310 -3400 -4280 -3370
rect -4110 -3400 -4080 -3370
rect -3910 -3400 -3880 -3370
rect -3710 -3400 -3680 -3370
rect -3510 -3400 -3480 -3370
rect -6310 -3520 -6280 -3490
rect -6310 -3640 -6280 -3610
rect -6310 -3760 -6280 -3730
rect -6310 -3880 -6280 -3850
rect -6310 -4000 -6280 -3970
rect -6310 -4120 -6280 -4090
rect -6310 -4370 -6280 -4340
rect -6310 -4490 -6280 -4460
rect -6310 -4610 -6280 -4580
rect -6310 -4730 -6280 -4700
rect -6310 -4850 -6280 -4820
rect -6310 -4970 -6280 -4940
rect -2670 -3460 -2640 -3430
rect -2060 -5030 -2030 -5000
rect -6390 -5090 -6360 -5060
rect -6310 -5090 -6280 -5060
rect -6110 -5090 -6080 -5060
rect -5910 -5090 -5880 -5060
rect -5710 -5090 -5680 -5060
rect -5510 -5090 -5480 -5060
rect -5310 -5090 -5280 -5060
rect -5110 -5090 -5080 -5060
rect -4710 -5090 -4680 -5060
rect -4510 -5090 -4480 -5060
rect -4310 -5090 -4280 -5060
rect -4110 -5090 -4080 -5060
rect -3910 -5090 -3880 -5060
rect -3710 -5090 -3680 -5060
rect -3510 -5090 -3480 -5060
rect -2790 -6490 -2760 -6350
rect -1730 -3460 -1700 -3430
rect -1000 -3460 -970 -3430
rect -910 -3580 -880 -3550
rect -60 -3460 -30 -3430
rect 150 -3460 180 -3430
rect -790 -3580 -760 -3550
rect 760 -4910 790 -4880
rect -1120 -5030 -1090 -5000
rect -910 -5030 -880 -5000
rect -180 -5030 -150 -5000
rect 30 -5030 60 -5000
rect 1090 -3460 1120 -3430
rect 1820 -3700 1850 -3670
rect 1910 -3700 1940 -3670
rect 2030 -3820 2060 -3790
rect 880 -4910 910 -4880
rect 970 -4060 1000 -4030
rect 1910 -4060 1940 -4030
rect 1700 -4550 1730 -4520
rect 2970 -3460 3000 -3430
rect 3700 -3700 3730 -3670
rect 3790 -3700 3820 -3670
rect 3910 -3940 3940 -3910
rect 2760 -4060 2790 -4030
rect 2850 -4430 2880 -4400
rect 2640 -4550 2670 -4520
rect 2760 -4550 2790 -4520
rect 3790 -4430 3820 -4400
rect 3580 -4550 3610 -4520
rect 4850 -3460 4880 -3430
rect 4640 -4430 4670 -4400
rect 4730 -4430 4760 -4400
rect 4520 -4550 4550 -4520
rect 4640 -4790 4670 -4760
rect 5460 -4550 5490 -4520
rect 5670 -3700 5700 -3670
rect 5790 -3940 5820 -3910
rect 5580 -4550 5610 -4520
rect 5670 -4430 5700 -4400
rect 6730 -3460 6760 -3430
rect 6520 -4430 6550 -4400
rect 6610 -4060 6640 -4030
rect 6400 -4550 6430 -4520
rect 6520 -4790 6550 -4760
rect 7340 -4550 7370 -4520
rect 7550 -3700 7580 -3670
rect 7670 -3820 7700 -3790
rect 7460 -4670 7490 -4640
rect 7550 -4060 7580 -4030
rect 8400 -4060 8430 -4030
rect 8280 -4550 8310 -4520
rect 8400 -4550 8430 -4520
rect 8610 -3580 8640 -3550
rect 8490 -4670 8520 -4640
rect 9340 -4790 9370 -4760
rect 9220 -4910 9250 -4880
rect 9430 -4300 9460 -4160
rect 10280 -4300 10310 -4160
rect 10370 -4300 10400 -4160
rect 9550 -4670 9580 -4640
rect 11100 -4670 11130 -4640
rect 11220 -4300 11250 -4160
rect 10160 -4790 10190 -4760
rect 10490 -4790 10520 -4760
rect 12040 -3580 12070 -3550
rect 11310 -4790 11340 -4760
rect 13100 -3700 13130 -3670
rect 12980 -3820 13010 -3790
rect 12250 -4060 12280 -4030
rect 13100 -4060 13130 -4030
rect 12160 -4670 12190 -4640
rect 11430 -4910 11460 -4880
rect 12250 -4550 12280 -4520
rect 12370 -4550 12400 -4520
rect 13920 -3460 13950 -3430
rect 14040 -4060 14070 -4030
rect 13190 -4670 13220 -4640
rect 13310 -4550 13340 -4520
rect 14980 -3700 15010 -3670
rect 14860 -3940 14890 -3910
rect 14130 -4430 14160 -4400
rect 14980 -4430 15010 -4400
rect 14250 -4550 14280 -4520
rect 14130 -4790 14160 -4760
rect 15800 -3460 15830 -3430
rect 15920 -4430 15950 -4400
rect 15070 -4550 15100 -4520
rect 15190 -4550 15220 -4520
rect 16860 -3700 16890 -3670
rect 17680 -3460 17710 -3430
rect 16950 -3700 16980 -3670
rect 16740 -3940 16770 -3910
rect 18740 -3700 18770 -3670
rect 19560 -3460 19590 -3430
rect 18830 -3700 18860 -3670
rect 18620 -3820 18650 -3790
rect 17890 -4060 17920 -4030
rect 18740 -4060 18770 -4030
rect 16010 -4430 16040 -4400
rect 16860 -4430 16890 -4400
rect 16130 -4550 16160 -4520
rect 16010 -4790 16040 -4760
rect 17800 -4430 17830 -4400
rect 17070 -4550 17100 -4520
rect 17890 -4550 17920 -4520
rect 18010 -4550 18040 -4520
rect 19680 -4060 19710 -4030
rect 18950 -4550 18980 -4520
rect 20500 -3460 20530 -3430
rect 20710 -3460 20740 -3430
rect 21440 -3580 21470 -3550
rect 21650 -3460 21680 -3430
rect 22380 -3460 22410 -3430
rect 21560 -3580 21590 -3550
rect 19770 -4910 19800 -4880
rect 19890 -4910 19920 -4880
rect 20620 -5030 20650 -5000
rect 20830 -5030 20860 -5000
rect 21560 -5030 21590 -5000
rect 21770 -5030 21800 -5000
rect 23320 -3460 23350 -3430
rect 24270 -4300 24410 -4160
rect 22710 -5030 22740 -5000
rect -1940 -6490 -1910 -6350
rect -1850 -6490 -1820 -6350
rect -910 -6490 -880 -6350
rect 970 -6490 1000 -6350
rect 2850 -6490 2880 -6350
rect 4730 -6490 4760 -6350
rect 6610 -6490 6640 -6350
rect 9430 -6490 9460 -6350
rect 11220 -6490 11250 -6350
rect 14040 -6490 14070 -6350
rect 15920 -6490 15950 -6350
rect 17800 -6490 17830 -6350
rect 19680 -6490 19710 -6350
rect 21560 -6490 21590 -6350
rect 22500 -6490 22530 -6350
rect 22590 -6490 22620 -6350
rect 23440 -6490 23470 -6350
<< metal2 >>
rect -3420 -230 24420 -220
rect -3420 -370 -3410 -230
rect -3270 -370 -2790 -230
rect -2760 -370 -1940 -230
rect -1910 -370 -1000 -230
rect -970 -370 880 -230
rect 910 -370 1820 -230
rect 1850 -370 3700 -230
rect 3730 -370 5580 -230
rect 5610 -370 7460 -230
rect 7490 -370 10280 -230
rect 10310 -370 10370 -230
rect 10400 -370 13190 -230
rect 13220 -370 15070 -230
rect 15100 -370 16950 -230
rect 16980 -370 18830 -230
rect 18860 -370 19770 -230
rect 19800 -370 21650 -230
rect 21680 -370 22590 -230
rect 22620 -370 23440 -230
rect 23470 -370 23950 -230
rect 24090 -370 24420 -230
rect -3420 -380 24420 -370
rect -6320 -3370 -6270 -3360
rect -6120 -3370 -6070 -3360
rect -5920 -3370 -5870 -3360
rect -5720 -3370 -5670 -3360
rect -5520 -3370 -5470 -3360
rect -5320 -3370 -5270 -3360
rect -5120 -3370 -5070 -3360
rect -4720 -3370 -4670 -3360
rect -4520 -3370 -4470 -3360
rect -4320 -3370 -4270 -3360
rect -4120 -3370 -4070 -3360
rect -3920 -3370 -3870 -3360
rect -3720 -3370 -3670 -3360
rect -3520 -3370 -3470 -3360
rect -6320 -3400 -6310 -3370
rect -6280 -3400 -6110 -3370
rect -6080 -3400 -5910 -3370
rect -5880 -3400 -5710 -3370
rect -5680 -3400 -5510 -3370
rect -5480 -3400 -5310 -3370
rect -5280 -3400 -5110 -3370
rect -5080 -3400 -4710 -3370
rect -4680 -3400 -4510 -3370
rect -4480 -3400 -4310 -3370
rect -4280 -3400 -4110 -3370
rect -4080 -3400 -3910 -3370
rect -3880 -3400 -3710 -3370
rect -3680 -3400 -3510 -3370
rect -3480 -3400 23620 -3370
rect -6320 -3410 -6270 -3400
rect -6120 -3410 -6070 -3400
rect -5920 -3410 -5870 -3400
rect -5720 -3410 -5670 -3400
rect -5520 -3410 -5470 -3400
rect -5320 -3410 -5270 -3400
rect -5120 -3410 -5070 -3400
rect -4720 -3410 -4670 -3400
rect -4520 -3410 -4470 -3400
rect -4320 -3410 -4270 -3400
rect -4120 -3410 -4070 -3400
rect -3920 -3410 -3870 -3400
rect -3720 -3410 -3670 -3400
rect -3520 -3410 -3470 -3400
rect -6220 -3430 -6170 -3420
rect -6310 -3460 -6210 -3430
rect -6180 -3460 -2670 -3430
rect -2640 -3460 -1730 -3430
rect -1700 -3460 -1000 -3430
rect -970 -3460 -60 -3430
rect -30 -3460 150 -3430
rect 180 -3460 1090 -3430
rect 1120 -3460 2970 -3430
rect 3000 -3460 4850 -3430
rect 4880 -3460 6730 -3430
rect 6760 -3460 13920 -3430
rect 13950 -3460 15800 -3430
rect 15830 -3460 17680 -3430
rect 17710 -3460 19560 -3430
rect 19590 -3460 20500 -3430
rect 20530 -3460 20710 -3430
rect 20740 -3460 21650 -3430
rect 21680 -3460 22380 -3430
rect 22410 -3460 23320 -3430
rect 23350 -3460 23620 -3430
rect -6220 -3470 -6170 -3460
rect -6320 -3490 -6270 -3480
rect -6320 -3520 -6310 -3490
rect -6280 -3520 23620 -3490
rect -6320 -3530 -6270 -3520
rect -6020 -3550 -5970 -3540
rect -6310 -3580 -6010 -3550
rect -5980 -3580 -910 -3550
rect -880 -3580 -790 -3550
rect -760 -3580 8610 -3550
rect 8640 -3580 12040 -3550
rect 12070 -3580 21440 -3550
rect 21470 -3580 21560 -3550
rect 21590 -3580 23620 -3550
rect -6020 -3590 -5970 -3580
rect -6320 -3610 -6270 -3600
rect -6320 -3640 -6310 -3610
rect -6280 -3640 23620 -3610
rect -6320 -3650 -6270 -3640
rect -5820 -3670 -5770 -3660
rect -6310 -3700 -5810 -3670
rect -5780 -3700 1820 -3670
rect 1850 -3700 1910 -3670
rect 1940 -3700 3700 -3670
rect 3730 -3700 3790 -3670
rect 3820 -3700 5670 -3670
rect 5700 -3700 7550 -3670
rect 7580 -3700 13100 -3670
rect 13130 -3700 14980 -3670
rect 15010 -3700 16860 -3670
rect 16890 -3700 16950 -3670
rect 16980 -3700 18740 -3670
rect 18770 -3700 18830 -3670
rect 18860 -3700 23620 -3670
rect -5820 -3710 -5770 -3700
rect -6320 -3730 -6270 -3720
rect -6320 -3760 -6310 -3730
rect -6280 -3760 23620 -3730
rect -6320 -3770 -6270 -3760
rect -5620 -3790 -5570 -3780
rect -6310 -3820 -5610 -3790
rect -5580 -3820 2030 -3790
rect 2060 -3820 7670 -3790
rect 7700 -3820 12980 -3790
rect 13010 -3820 18620 -3790
rect 18650 -3820 23620 -3790
rect -5620 -3830 -5570 -3820
rect -6320 -3850 -6270 -3840
rect -6320 -3880 -6310 -3850
rect -6280 -3880 23620 -3850
rect -6320 -3890 -6270 -3880
rect -5420 -3910 -5370 -3900
rect -6310 -3940 -5410 -3910
rect -5380 -3940 3910 -3910
rect 3940 -3940 5790 -3910
rect 5820 -3940 14860 -3910
rect 14890 -3940 16740 -3910
rect 16770 -3940 23620 -3910
rect -5420 -3950 -5370 -3940
rect -6320 -3970 -6270 -3960
rect -6320 -4000 -6310 -3970
rect -6280 -4000 23620 -3970
rect -6320 -4010 -6270 -4000
rect -5220 -4030 -5170 -4020
rect -6310 -4060 -5210 -4030
rect -5180 -4060 970 -4030
rect 1000 -4060 1910 -4030
rect 1940 -4060 2760 -4030
rect 2790 -4060 6610 -4030
rect 6640 -4060 7550 -4030
rect 7580 -4060 8400 -4030
rect 8430 -4060 12250 -4030
rect 12280 -4060 13100 -4030
rect 13130 -4060 14040 -4030
rect 14070 -4060 17890 -4030
rect 17920 -4060 18740 -4030
rect 18770 -4060 19680 -4030
rect 19710 -4060 23620 -4030
rect -5220 -4070 -5170 -4060
rect -6320 -4090 -6270 -4080
rect -6320 -4120 -6310 -4090
rect -6280 -4120 23620 -4090
rect -6320 -4130 -6270 -4120
rect -6310 -4160 23620 -4150
rect -6310 -4300 -5000 -4160
rect -4790 -4300 9430 -4160
rect 9460 -4300 10280 -4160
rect 10310 -4300 10370 -4160
rect 10400 -4300 11220 -4160
rect 11250 -4300 23620 -4160
rect -6310 -4310 23620 -4300
rect 24260 -4160 24420 -4150
rect 24260 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect 24260 -4310 24420 -4300
rect -6320 -4340 -6270 -4330
rect -6320 -4370 -6310 -4340
rect -6280 -4370 23620 -4340
rect -6320 -4380 -6270 -4370
rect -4620 -4400 -4570 -4390
rect -6310 -4430 -4610 -4400
rect -4580 -4430 2850 -4400
rect 2880 -4430 3790 -4400
rect 3820 -4430 4640 -4400
rect 4670 -4430 4730 -4400
rect 4760 -4430 5670 -4400
rect 5700 -4430 6520 -4400
rect 6550 -4430 14130 -4400
rect 14160 -4430 14980 -4400
rect 15010 -4430 15920 -4400
rect 15950 -4430 16010 -4400
rect 16040 -4430 16860 -4400
rect 16890 -4430 17800 -4400
rect 17830 -4430 23620 -4400
rect -4620 -4440 -4570 -4430
rect -6320 -4460 -6270 -4450
rect -6320 -4490 -6310 -4460
rect -6280 -4490 23620 -4460
rect -6320 -4500 -6270 -4490
rect -4420 -4520 -4370 -4510
rect -6310 -4550 -4410 -4520
rect -4380 -4550 1700 -4520
rect 1730 -4550 2640 -4520
rect 2670 -4550 2760 -4520
rect 2790 -4550 3580 -4520
rect 3610 -4550 4520 -4520
rect 4550 -4550 5460 -4520
rect 5490 -4550 5580 -4520
rect 5610 -4550 6400 -4520
rect 6430 -4550 7340 -4520
rect 7370 -4550 8280 -4520
rect 8310 -4550 8400 -4520
rect 8430 -4550 12250 -4520
rect 12280 -4550 12370 -4520
rect 12400 -4550 13310 -4520
rect 13340 -4550 14250 -4520
rect 14280 -4550 15070 -4520
rect 15100 -4550 15190 -4520
rect 15220 -4550 16130 -4520
rect 16160 -4550 17070 -4520
rect 17100 -4550 17890 -4520
rect 17920 -4550 18010 -4520
rect 18040 -4550 18950 -4520
rect 18980 -4550 23620 -4520
rect -4420 -4560 -4370 -4550
rect -6320 -4580 -6270 -4570
rect -6320 -4610 -6310 -4580
rect -6280 -4610 23620 -4580
rect -6320 -4620 -6270 -4610
rect -4220 -4640 -4170 -4630
rect -6310 -4670 -4210 -4640
rect -4180 -4670 7460 -4640
rect 7490 -4670 8490 -4640
rect 8520 -4670 9550 -4640
rect 9580 -4670 11100 -4640
rect 11130 -4670 12160 -4640
rect 12190 -4670 13190 -4640
rect 13220 -4670 23620 -4640
rect -4220 -4680 -4170 -4670
rect -6320 -4700 -6270 -4690
rect -6320 -4730 -6310 -4700
rect -6280 -4730 23620 -4700
rect -6320 -4740 -6270 -4730
rect -4020 -4760 -3970 -4750
rect -6310 -4790 -4010 -4760
rect -3980 -4790 4640 -4760
rect 4670 -4790 6520 -4760
rect 6550 -4790 9340 -4760
rect 9370 -4790 10160 -4760
rect 10190 -4790 10490 -4760
rect 10520 -4790 11310 -4760
rect 11340 -4790 14130 -4760
rect 14160 -4790 16010 -4760
rect 16040 -4790 23620 -4760
rect -4020 -4800 -3970 -4790
rect -6320 -4820 -6270 -4810
rect -6320 -4850 -6310 -4820
rect -6280 -4850 23620 -4820
rect -6320 -4860 -6270 -4850
rect -3820 -4880 -3770 -4870
rect -6310 -4910 -3810 -4880
rect -3780 -4910 760 -4880
rect 790 -4910 880 -4880
rect 910 -4910 9220 -4880
rect 9250 -4910 11430 -4880
rect 11460 -4910 19770 -4880
rect 19800 -4910 19890 -4880
rect 19920 -4910 23620 -4880
rect -3820 -4920 -3770 -4910
rect -6320 -4940 -6270 -4930
rect -6320 -4970 -6310 -4940
rect -6280 -4970 23620 -4940
rect -6320 -4980 -6270 -4970
rect -3620 -5000 -3570 -4990
rect -6310 -5030 -3610 -5000
rect -3580 -5030 -2060 -5000
rect -2030 -5030 -1120 -5000
rect -1090 -5030 -910 -5000
rect -880 -5030 -180 -5000
rect -150 -5030 30 -5000
rect 60 -5030 20620 -5000
rect 20650 -5030 20830 -5000
rect 20860 -5030 21560 -5000
rect 21590 -5030 21770 -5000
rect 21800 -5030 22710 -5000
rect 22740 -5030 23620 -5000
rect -3620 -5040 -3570 -5030
rect -6400 -5060 -6350 -5050
rect -6400 -5090 -6390 -5060
rect -6360 -5090 -6350 -5060
rect -6400 -5100 -6350 -5090
rect -6320 -5060 -6270 -5050
rect -6120 -5060 -6070 -5050
rect -5920 -5060 -5870 -5050
rect -5720 -5060 -5670 -5050
rect -5520 -5060 -5470 -5050
rect -5320 -5060 -5270 -5050
rect -5120 -5060 -5070 -5050
rect -4720 -5060 -4670 -5050
rect -4520 -5060 -4470 -5050
rect -4320 -5060 -4270 -5050
rect -4120 -5060 -4070 -5050
rect -3920 -5060 -3870 -5050
rect -3720 -5060 -3670 -5050
rect -3520 -5060 -3470 -5050
rect -6320 -5090 -6310 -5060
rect -6280 -5090 -6110 -5060
rect -6080 -5090 -5910 -5060
rect -5880 -5090 -5710 -5060
rect -5680 -5090 -5510 -5060
rect -5480 -5090 -5310 -5060
rect -5280 -5090 -5110 -5060
rect -5080 -5090 -4710 -5060
rect -4680 -5090 -4510 -5060
rect -4480 -5090 -4310 -5060
rect -4280 -5090 -4110 -5060
rect -4080 -5090 -3910 -5060
rect -3880 -5090 -3710 -5060
rect -3680 -5090 -3510 -5060
rect -3480 -5090 23620 -5060
rect -6320 -5100 -6270 -5090
rect -6120 -5100 -6070 -5090
rect -5920 -5100 -5870 -5090
rect -5720 -5100 -5670 -5090
rect -5520 -5100 -5470 -5090
rect -5320 -5100 -5270 -5090
rect -5120 -5100 -5070 -5090
rect -4720 -5100 -4670 -5090
rect -4520 -5100 -4470 -5090
rect -4320 -5100 -4270 -5090
rect -4120 -5100 -4070 -5090
rect -3920 -5100 -3870 -5090
rect -3720 -5100 -3670 -5090
rect -3520 -5100 -3470 -5090
rect -3100 -6350 24420 -6340
rect -3100 -6490 -3090 -6350
rect -2950 -6490 -2790 -6350
rect -2760 -6490 -1940 -6350
rect -1910 -6490 -1850 -6350
rect -1820 -6490 -910 -6350
rect -880 -6490 970 -6350
rect 1000 -6490 2850 -6350
rect 2880 -6490 4730 -6350
rect 4760 -6490 6610 -6350
rect 6640 -6490 9430 -6350
rect 9460 -6490 11220 -6350
rect 11250 -6490 14040 -6350
rect 14070 -6490 15920 -6350
rect 15950 -6490 17800 -6350
rect 17830 -6490 19680 -6350
rect 19710 -6490 21560 -6350
rect 21590 -6490 22500 -6350
rect 22530 -6490 22590 -6350
rect 22620 -6490 23440 -6350
rect 23470 -6490 23630 -6350
rect 23770 -6490 24420 -6350
rect -3100 -6500 24420 -6490
<< via2 >>
rect -3410 -370 -3270 -230
rect 23950 -370 24090 -230
rect -6310 -3400 -6280 -3370
rect -6110 -3400 -6080 -3370
rect -5910 -3400 -5880 -3370
rect -5710 -3400 -5680 -3370
rect -5510 -3400 -5480 -3370
rect -5310 -3400 -5280 -3370
rect -5110 -3400 -5080 -3370
rect -4710 -3400 -4680 -3370
rect -4510 -3400 -4480 -3370
rect -4310 -3400 -4280 -3370
rect -4110 -3400 -4080 -3370
rect -3910 -3400 -3880 -3370
rect -3710 -3400 -3680 -3370
rect -3510 -3400 -3480 -3370
rect -6210 -3460 -6180 -3430
rect -6310 -3520 -6280 -3490
rect -6010 -3580 -5980 -3550
rect -6310 -3640 -6280 -3610
rect -5810 -3700 -5780 -3670
rect -6310 -3760 -6280 -3730
rect -5610 -3820 -5580 -3790
rect -6310 -3880 -6280 -3850
rect -5410 -3940 -5380 -3910
rect -6310 -4000 -6280 -3970
rect -5210 -4060 -5180 -4030
rect -6310 -4120 -6280 -4090
rect -5000 -4300 -4790 -4160
rect 24270 -4300 24410 -4160
rect -6310 -4370 -6280 -4340
rect -4610 -4430 -4580 -4400
rect -6310 -4490 -6280 -4460
rect -4410 -4550 -4380 -4520
rect -6310 -4610 -6280 -4580
rect -4210 -4670 -4180 -4640
rect -6310 -4730 -6280 -4700
rect -4010 -4790 -3980 -4760
rect -6310 -4850 -6280 -4820
rect -3810 -4910 -3780 -4880
rect -6310 -4970 -6280 -4940
rect -3610 -5030 -3580 -5000
rect -6390 -5090 -6360 -5060
rect -6310 -5090 -6280 -5060
rect -6110 -5090 -6080 -5060
rect -5910 -5090 -5880 -5060
rect -5710 -5090 -5680 -5060
rect -5510 -5090 -5480 -5060
rect -5310 -5090 -5280 -5060
rect -5110 -5090 -5080 -5060
rect -4710 -5090 -4680 -5060
rect -4510 -5090 -4480 -5060
rect -4310 -5090 -4280 -5060
rect -4110 -5090 -4080 -5060
rect -3910 -5090 -3880 -5060
rect -3710 -5090 -3680 -5060
rect -3510 -5090 -3480 -5060
rect -3090 -6490 -2950 -6350
rect 23630 -6490 23770 -6350
<< metal3 >>
rect -6310 -3360 -6280 -220
rect -6320 -3370 -6270 -3360
rect -6320 -3400 -6310 -3370
rect -6280 -3400 -6270 -3370
rect -6320 -3410 -6270 -3400
rect -6310 -3480 -6280 -3410
rect -6210 -3420 -6180 -190
rect -6110 -3360 -6080 -220
rect -6120 -3370 -6070 -3360
rect -6120 -3400 -6110 -3370
rect -6080 -3400 -6070 -3370
rect -6120 -3410 -6070 -3400
rect -6220 -3430 -6170 -3420
rect -6220 -3460 -6210 -3430
rect -6180 -3460 -6170 -3430
rect -6220 -3470 -6170 -3460
rect -6320 -3490 -6270 -3480
rect -6320 -3520 -6310 -3490
rect -6280 -3520 -6270 -3490
rect -6320 -3530 -6270 -3520
rect -6310 -3600 -6280 -3530
rect -6320 -3610 -6270 -3600
rect -6320 -3640 -6310 -3610
rect -6280 -3640 -6270 -3610
rect -6320 -3650 -6270 -3640
rect -6310 -3720 -6280 -3650
rect -6320 -3730 -6270 -3720
rect -6320 -3760 -6310 -3730
rect -6280 -3760 -6270 -3730
rect -6320 -3770 -6270 -3760
rect -6310 -3840 -6280 -3770
rect -6320 -3850 -6270 -3840
rect -6320 -3880 -6310 -3850
rect -6280 -3880 -6270 -3850
rect -6320 -3890 -6270 -3880
rect -6310 -3960 -6280 -3890
rect -6320 -3970 -6270 -3960
rect -6320 -4000 -6310 -3970
rect -6280 -4000 -6270 -3970
rect -6320 -4010 -6270 -4000
rect -6310 -4080 -6280 -4010
rect -6320 -4090 -6270 -4080
rect -6320 -4120 -6310 -4090
rect -6280 -4120 -6270 -4090
rect -6320 -4130 -6270 -4120
rect -6310 -4330 -6280 -4130
rect -6320 -4340 -6270 -4330
rect -6320 -4370 -6310 -4340
rect -6280 -4370 -6270 -4340
rect -6320 -4380 -6270 -4370
rect -6310 -4450 -6280 -4380
rect -6320 -4460 -6270 -4450
rect -6320 -4490 -6310 -4460
rect -6280 -4490 -6270 -4460
rect -6320 -4500 -6270 -4490
rect -6310 -4570 -6280 -4500
rect -6320 -4580 -6270 -4570
rect -6320 -4610 -6310 -4580
rect -6280 -4610 -6270 -4580
rect -6320 -4620 -6270 -4610
rect -6310 -4690 -6280 -4620
rect -6320 -4700 -6270 -4690
rect -6320 -4730 -6310 -4700
rect -6280 -4730 -6270 -4700
rect -6320 -4740 -6270 -4730
rect -6310 -4810 -6280 -4740
rect -6320 -4820 -6270 -4810
rect -6320 -4850 -6310 -4820
rect -6280 -4850 -6270 -4820
rect -6320 -4860 -6270 -4850
rect -6310 -4930 -6280 -4860
rect -6320 -4940 -6270 -4930
rect -6320 -4970 -6310 -4940
rect -6280 -4970 -6270 -4940
rect -6320 -4980 -6270 -4970
rect -6310 -5050 -6280 -4980
rect -6400 -5060 -6350 -5050
rect -6400 -5090 -6390 -5060
rect -6360 -5090 -6350 -5060
rect -6400 -5100 -6350 -5090
rect -6320 -5060 -6270 -5050
rect -6320 -5090 -6310 -5060
rect -6280 -5090 -6270 -5060
rect -6320 -5100 -6270 -5090
rect -6310 -6500 -6280 -5100
rect -6210 -6500 -6180 -3470
rect -6110 -5050 -6080 -3410
rect -6010 -3540 -5980 -190
rect -5910 -3360 -5880 -220
rect -5920 -3370 -5870 -3360
rect -5920 -3400 -5910 -3370
rect -5880 -3400 -5870 -3370
rect -5920 -3410 -5870 -3400
rect -6020 -3550 -5970 -3540
rect -6020 -3580 -6010 -3550
rect -5980 -3580 -5970 -3550
rect -6020 -3590 -5970 -3580
rect -6120 -5060 -6070 -5050
rect -6120 -5090 -6110 -5060
rect -6080 -5090 -6070 -5060
rect -6120 -5100 -6070 -5090
rect -6110 -6500 -6080 -5100
rect -6010 -6500 -5980 -3590
rect -5910 -5050 -5880 -3410
rect -5810 -3660 -5780 -190
rect -5710 -3360 -5680 -220
rect -5720 -3370 -5670 -3360
rect -5720 -3400 -5710 -3370
rect -5680 -3400 -5670 -3370
rect -5720 -3410 -5670 -3400
rect -5820 -3670 -5770 -3660
rect -5820 -3700 -5810 -3670
rect -5780 -3700 -5770 -3670
rect -5820 -3710 -5770 -3700
rect -5920 -5060 -5870 -5050
rect -5920 -5090 -5910 -5060
rect -5880 -5090 -5870 -5060
rect -5920 -5100 -5870 -5090
rect -5910 -6500 -5880 -5100
rect -5810 -6500 -5780 -3710
rect -5710 -5050 -5680 -3410
rect -5610 -3780 -5580 -190
rect -5510 -3360 -5480 -220
rect -5520 -3370 -5470 -3360
rect -5520 -3400 -5510 -3370
rect -5480 -3400 -5470 -3370
rect -5520 -3410 -5470 -3400
rect -5620 -3790 -5570 -3780
rect -5620 -3820 -5610 -3790
rect -5580 -3820 -5570 -3790
rect -5620 -3830 -5570 -3820
rect -5720 -5060 -5670 -5050
rect -5720 -5090 -5710 -5060
rect -5680 -5090 -5670 -5060
rect -5720 -5100 -5670 -5090
rect -5710 -6500 -5680 -5100
rect -5610 -6500 -5580 -3830
rect -5510 -5050 -5480 -3410
rect -5410 -3900 -5380 -190
rect -5310 -3360 -5280 -220
rect -5320 -3370 -5270 -3360
rect -5320 -3400 -5310 -3370
rect -5280 -3400 -5270 -3370
rect -5320 -3410 -5270 -3400
rect -5420 -3910 -5370 -3900
rect -5420 -3940 -5410 -3910
rect -5380 -3940 -5370 -3910
rect -5420 -3950 -5370 -3940
rect -5520 -5060 -5470 -5050
rect -5520 -5090 -5510 -5060
rect -5480 -5090 -5470 -5060
rect -5520 -5100 -5470 -5090
rect -5510 -6500 -5480 -5100
rect -5410 -6500 -5380 -3950
rect -5310 -5050 -5280 -3410
rect -5210 -4020 -5180 -190
rect -5110 -3360 -5080 -220
rect -5120 -3370 -5070 -3360
rect -5120 -3400 -5110 -3370
rect -5080 -3400 -5070 -3370
rect -5120 -3410 -5070 -3400
rect -5220 -4030 -5170 -4020
rect -5220 -4060 -5210 -4030
rect -5180 -4060 -5170 -4030
rect -5220 -4070 -5170 -4060
rect -5320 -5060 -5270 -5050
rect -5320 -5090 -5310 -5060
rect -5280 -5090 -5270 -5060
rect -5320 -5100 -5270 -5090
rect -5310 -6500 -5280 -5100
rect -5210 -6500 -5180 -4070
rect -5110 -5050 -5080 -3410
rect -5010 -4160 -4780 -190
rect -4710 -3360 -4680 -220
rect -4720 -3370 -4670 -3360
rect -4720 -3400 -4710 -3370
rect -4680 -3400 -4670 -3370
rect -4720 -3410 -4670 -3400
rect -5010 -4300 -5000 -4160
rect -4790 -4300 -4780 -4160
rect -5120 -5060 -5070 -5050
rect -5120 -5090 -5110 -5060
rect -5080 -5090 -5070 -5060
rect -5120 -5100 -5070 -5090
rect -5110 -6500 -5080 -5100
rect -5010 -6500 -4780 -4300
rect -4710 -5050 -4680 -3410
rect -4610 -4390 -4580 -190
rect -4510 -3360 -4480 -220
rect -4520 -3370 -4470 -3360
rect -4520 -3400 -4510 -3370
rect -4480 -3400 -4470 -3370
rect -4520 -3410 -4470 -3400
rect -4620 -4400 -4570 -4390
rect -4620 -4430 -4610 -4400
rect -4580 -4430 -4570 -4400
rect -4620 -4440 -4570 -4430
rect -4720 -5060 -4670 -5050
rect -4720 -5090 -4710 -5060
rect -4680 -5090 -4670 -5060
rect -4720 -5100 -4670 -5090
rect -4710 -6500 -4680 -5100
rect -4610 -6500 -4580 -4440
rect -4510 -5050 -4480 -3410
rect -4410 -4510 -4380 -190
rect -4310 -3360 -4280 -220
rect -4320 -3370 -4270 -3360
rect -4320 -3400 -4310 -3370
rect -4280 -3400 -4270 -3370
rect -4320 -3410 -4270 -3400
rect -4420 -4520 -4370 -4510
rect -4420 -4550 -4410 -4520
rect -4380 -4550 -4370 -4520
rect -4420 -4560 -4370 -4550
rect -4520 -5060 -4470 -5050
rect -4520 -5090 -4510 -5060
rect -4480 -5090 -4470 -5060
rect -4520 -5100 -4470 -5090
rect -4510 -6500 -4480 -5100
rect -4410 -6500 -4380 -4560
rect -4310 -5050 -4280 -3410
rect -4210 -4630 -4180 -190
rect -4110 -3360 -4080 -220
rect -4120 -3370 -4070 -3360
rect -4120 -3400 -4110 -3370
rect -4080 -3400 -4070 -3370
rect -4120 -3410 -4070 -3400
rect -4220 -4640 -4170 -4630
rect -4220 -4670 -4210 -4640
rect -4180 -4670 -4170 -4640
rect -4220 -4680 -4170 -4670
rect -4320 -5060 -4270 -5050
rect -4320 -5090 -4310 -5060
rect -4280 -5090 -4270 -5060
rect -4320 -5100 -4270 -5090
rect -4310 -6500 -4280 -5100
rect -4210 -6500 -4180 -4680
rect -4110 -5050 -4080 -3410
rect -4010 -4750 -3980 -190
rect -3910 -3360 -3880 -220
rect -3920 -3370 -3870 -3360
rect -3920 -3400 -3910 -3370
rect -3880 -3400 -3870 -3370
rect -3920 -3410 -3870 -3400
rect -4020 -4760 -3970 -4750
rect -4020 -4790 -4010 -4760
rect -3980 -4790 -3970 -4760
rect -4020 -4800 -3970 -4790
rect -4120 -5060 -4070 -5050
rect -4120 -5090 -4110 -5060
rect -4080 -5090 -4070 -5060
rect -4120 -5100 -4070 -5090
rect -4110 -6500 -4080 -5100
rect -4010 -6500 -3980 -4800
rect -3910 -5050 -3880 -3410
rect -3810 -4870 -3780 -190
rect -3710 -3360 -3680 -220
rect -3720 -3370 -3670 -3360
rect -3720 -3400 -3710 -3370
rect -3680 -3400 -3670 -3370
rect -3720 -3410 -3670 -3400
rect -3820 -4880 -3770 -4870
rect -3820 -4910 -3810 -4880
rect -3780 -4910 -3770 -4880
rect -3820 -4920 -3770 -4910
rect -3920 -5060 -3870 -5050
rect -3920 -5090 -3910 -5060
rect -3880 -5090 -3870 -5060
rect -3920 -5100 -3870 -5090
rect -3910 -6500 -3880 -5100
rect -3810 -6500 -3780 -4920
rect -3710 -5050 -3680 -3410
rect -3610 -4990 -3580 -190
rect -3510 -3360 -3480 -220
rect -3420 -230 -3260 -220
rect -3420 -370 -3410 -230
rect -3270 -370 -3260 -230
rect -3520 -3370 -3470 -3360
rect -3520 -3400 -3510 -3370
rect -3480 -3400 -3470 -3370
rect -3520 -3410 -3470 -3400
rect -3620 -5000 -3570 -4990
rect -3620 -5030 -3610 -5000
rect -3580 -5030 -3570 -5000
rect -3620 -5040 -3570 -5030
rect -3720 -5060 -3670 -5050
rect -3720 -5090 -3710 -5060
rect -3680 -5090 -3670 -5060
rect -3720 -5100 -3670 -5090
rect -3710 -6500 -3680 -5100
rect -3610 -6500 -3580 -5040
rect -3510 -5050 -3480 -3410
rect -3520 -5060 -3470 -5050
rect -3520 -5090 -3510 -5060
rect -3480 -5090 -3470 -5060
rect -3520 -5100 -3470 -5090
rect -3510 -6500 -3480 -5100
rect -3420 -6500 -3260 -370
rect -3100 -6350 -2940 -220
rect -3100 -6490 -3090 -6350
rect -2950 -6490 -2940 -6350
rect -3100 -6500 -2940 -6490
rect 23620 -6350 23780 -190
rect 23620 -6490 23630 -6350
rect 23770 -6490 23780 -6350
rect 23620 -6500 23780 -6490
rect 23940 -230 24100 -190
rect 23940 -370 23950 -230
rect 24090 -370 24100 -230
rect 23940 -6500 24100 -370
rect 24260 -3440 24420 -190
rect 24260 -3570 24270 -3440
rect 24410 -3570 24420 -3440
rect 24260 -3680 24420 -3570
rect 24260 -3810 24270 -3680
rect 24410 -3810 24420 -3680
rect 24260 -3920 24420 -3810
rect 24260 -4050 24270 -3920
rect 24410 -4050 24420 -3920
rect 24260 -4160 24420 -4050
rect 24260 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect 24260 -4410 24420 -4300
rect 24260 -4540 24270 -4410
rect 24410 -4540 24420 -4410
rect 24260 -4650 24420 -4540
rect 24260 -4780 24270 -4650
rect 24410 -4780 24420 -4650
rect 24260 -4890 24420 -4780
rect 24260 -5020 24270 -4890
rect 24410 -5020 24420 -4890
rect 24260 -6500 24420 -5020
<< via3 >>
rect 24270 -3570 24410 -3440
rect 24270 -3810 24410 -3680
rect 24270 -4050 24410 -3920
rect 24270 -4300 24410 -4160
rect 24270 -4540 24410 -4410
rect 24270 -4780 24410 -4650
rect 24270 -5020 24410 -4890
<< metal4 >>
rect -3510 -3440 24420 -3430
rect -3510 -3570 24270 -3440
rect 24410 -3570 24420 -3440
rect -3510 -3580 24420 -3570
rect -3510 -3680 24420 -3670
rect -3510 -3810 24270 -3680
rect 24410 -3810 24420 -3680
rect -3510 -3820 24420 -3810
rect -3510 -3920 24420 -3910
rect -3510 -4050 24270 -3920
rect 24410 -4050 24420 -3920
rect -3510 -4060 24420 -4050
rect -3510 -4160 24420 -4150
rect -3510 -4300 24270 -4160
rect 24410 -4300 24420 -4160
rect -3510 -4310 24420 -4300
rect -3510 -4410 24420 -4400
rect -3510 -4540 24270 -4410
rect 24410 -4540 24420 -4410
rect -3510 -4550 24420 -4540
rect -3510 -4650 24420 -4640
rect -3510 -4780 24270 -4650
rect 24410 -4780 24420 -4650
rect -3510 -4790 24420 -4780
rect -3510 -4890 24420 -4880
rect -3510 -5020 24270 -4890
rect 24410 -5020 24420 -4890
rect -3510 -5030 24420 -5020
<< metal5 >>
rect -6180 -6500 -5950 -220
rect -5780 -6500 -5550 -220
rect -5380 -6500 -5150 -220
rect -4980 -6500 -4750 -220
rect -4580 -6500 -4350 -220
rect -4180 -6500 -3950 -220
rect -3780 -6500 -3550 -220
use n8_1  n8_1_8
timestamp 1634429522
transform 1 0 -2820 0 1 -6330
box 0 0 940 1230
use n1_8  na4_1
timestamp 1634337365
transform 1 0 -1880 0 1 -6330
box 0 0 940 1230
use p1_8  pa1_1
timestamp 1634440922
transform 1 0 -1880 0 1 -3360
box 0 0 940 2970
use p8_1  p8_1_7
timestamp 1634440961
transform 1 0 -2820 0 1 -3360
box 0 0 940 2970
use n1_8  nb4_1
timestamp 1634337365
transform 1 0 -940 0 1 -6330
box 0 0 940 1230
use p8_1  pa2_1
timestamp 1634440961
transform 1 0 -940 0 1 -3360
box 0 0 940 2970
use n8_1  nb3_1
timestamp 1634429522
transform 1 0 0 0 1 -6330
box 0 0 940 1230
use p1_8  pb1_1
timestamp 1634440922
transform 1 0 0 0 1 -3360
box 0 0 940 2970
use n1_8  ne4_1
timestamp 1634337365
transform 1 0 940 0 1 -6330
box 0 0 940 1230
use p1_8  pc1_1
timestamp 1634440922
transform 1 0 940 0 1 -3360
box 0 0 940 2970
use n8_1  ne3_1
timestamp 1634429522
transform 1 0 1880 0 1 -6330
box 0 0 940 1230
use p8_1  pc2_1
timestamp 1634440961
transform 1 0 1880 0 1 -3360
box 0 0 940 2970
use n1_8  nf4_1
timestamp 1634337365
transform 1 0 2820 0 1 -6330
box 0 0 940 1230
use p1_8  pd1_1
timestamp 1634440922
transform 1 0 2820 0 1 -3360
box 0 0 940 2970
use n8_1  nf3_1
timestamp 1634429522
transform 1 0 3760 0 1 -6330
box 0 0 940 1230
use p8_1  pd2_1
timestamp 1634440961
transform 1 0 3760 0 1 -3360
box 0 0 940 2970
use n1_8  nf4_2
timestamp 1634337365
transform 1 0 4700 0 1 -6330
box 0 0 940 1230
use p1_8  pe1_1
timestamp 1634440922
transform 1 0 4700 0 1 -3360
box 0 0 940 2970
use n8_1  nf3_2
timestamp 1634429522
transform 1 0 5640 0 1 -6330
box 0 0 940 1230
use p8_1  pd2_2
timestamp 1634440961
transform 1 0 5640 0 1 -3360
box 0 0 940 2970
use n1_8  ne4_2
timestamp 1634337365
transform 1 0 6580 0 1 -6330
box 0 0 940 1230
use p1_8  pf1_1
timestamp 1634440922
transform 1 0 6580 0 1 -3360
box 0 0 940 2970
use n8_1  ne3_2
timestamp 1634429522
transform 1 0 7520 0 1 -6330
box 0 0 940 1230
use p8_1  pc2_2
timestamp 1634440961
transform 1 0 7520 0 1 -3360
box 0 0 940 2970
use n8_1  nf2_1
timestamp 1634429522
transform 1 0 8460 0 1 -6330
box 0 0 940 1230
use p8_1  pf2_1
timestamp 1634440961
transform 1 0 8460 0 1 -3360
box 0 0 940 2970
use p4_2  p4_2_0
timestamp 1634665005
transform 1 0 9400 0 1 -3360
box 0 0 940 2970
use n4_2  n4_2_0
timestamp 1634664854
transform 1 0 9400 0 1 -6330
box 0 0 940 1230
use p4_2  p4_2_1
timestamp 1634665005
transform -1 0 11280 0 1 -3360
box 0 0 940 2970
use n4_2  n4_2_1
timestamp 1634664854
transform -1 0 11280 0 1 -6330
box 0 0 940 1230
use n8_1  n8_1_5
timestamp 1634429522
transform -1 0 12220 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_5
timestamp 1634440961
transform -1 0 12220 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_4
timestamp 1634429522
transform -1 0 13160 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_4
timestamp 1634440961
transform -1 0 13160 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_5
timestamp 1634337365
transform -1 0 14100 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_5
timestamp 1634440922
transform -1 0 14100 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_3
timestamp 1634429522
transform -1 0 15040 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_3
timestamp 1634440961
transform -1 0 15040 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_4
timestamp 1634337365
transform -1 0 15980 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_4
timestamp 1634440922
transform -1 0 15980 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_2
timestamp 1634429522
transform -1 0 16920 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_2
timestamp 1634440961
transform -1 0 16920 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_3
timestamp 1634337365
transform -1 0 17860 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_3
timestamp 1634440922
transform -1 0 17860 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_1
timestamp 1634429522
transform -1 0 18800 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_1
timestamp 1634440961
transform -1 0 18800 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_2
timestamp 1634337365
transform -1 0 19740 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_2
timestamp 1634440922
transform -1 0 19740 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_0
timestamp 1634429522
transform -1 0 20680 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_1
timestamp 1634440922
transform -1 0 20680 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_0
timestamp 1634337365
transform -1 0 21620 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_0
timestamp 1634440961
transform -1 0 21620 0 1 -3360
box 0 0 940 2970
use n1_8  n1_8_1
timestamp 1634337365
transform -1 0 22560 0 1 -6330
box 0 0 940 1230
use p1_8  p1_8_0
timestamp 1634440922
transform -1 0 22560 0 1 -3360
box 0 0 940 2970
use n8_1  n8_1_7
timestamp 1634429522
transform -1 0 23500 0 1 -6330
box 0 0 940 1230
use p8_1  p8_1_8
timestamp 1634440961
transform -1 0 23500 0 1 -3360
box 0 0 940 2970
<< labels >>
rlabel metal3 23940 -220 24100 -190 1 vdda
port 5 n
rlabel metal3 24260 -220 24420 -190 1 gnda
port 6 n
rlabel metal3 23620 -220 23780 -190 1 vssa
port 7 n
rlabel metal3 -3610 -220 -3580 -190 1 n1
rlabel metal3 -3810 -220 -3780 -190 1 n2
rlabel metal3 -4010 -220 -3980 -190 1 c
rlabel metal3 -4210 -220 -4180 -190 1 b
rlabel metal3 -4410 -220 -4380 -190 1 a
rlabel metal3 -4610 -220 -4580 -190 1 xp
rlabel metal3 -5010 -220 -4780 -190 1 out
port 3 n
rlabel metal3 -5610 -220 -5580 -190 1 inm
port 1 n
rlabel metal3 -5410 -220 -5380 -190 1 inp
port 2 n
rlabel metal3 -5210 -220 -5180 -190 1 xm
rlabel metal3 -5810 -220 -5780 -190 1 x
rlabel metal3 -6210 -220 -6180 -190 1 p1
rlabel metal3 -6010 -220 -5980 -190 1 ib
port 4 n
rlabel metal2 -6310 -3820 -6300 -3790 3 inm
<< end >>
