magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_p >>
rect 8 10000 8392 10072
rect 8 9920 80 10000
rect 94 9960 8306 9986
rect 94 8840 120 9960
rect 160 9894 8240 9920
rect 160 8952 232 9894
rect 8214 8952 8240 9894
rect 160 8880 8240 8952
rect 8280 8840 8306 9960
rect 8320 8880 8392 10000
rect 94 8814 8306 8840
rect 8 5360 8392 5432
rect 8 5280 80 5360
rect 94 5320 8306 5346
rect 94 4200 120 5320
rect 160 5254 8240 5280
rect 160 4312 232 5254
rect 8214 4312 8240 5254
rect 160 4240 8240 4312
rect 8280 4200 8306 5320
rect 8320 4240 8392 5360
rect 94 4174 8306 4200
rect 8 3920 8392 3992
rect 8 3840 80 3920
rect 94 3880 8306 3906
rect 94 2760 120 3880
rect 160 3814 8240 3840
rect 160 2872 232 3814
rect 8214 2872 8240 3814
rect 160 2800 8240 2872
rect 8280 2760 8306 3880
rect 8320 2800 8392 3920
rect 94 2734 8306 2760
rect 8 2480 8392 2552
rect 8 2400 80 2480
rect 94 2440 8306 2466
rect 94 1320 120 2440
rect 160 2374 8240 2400
rect 160 1432 232 2374
rect 8214 1432 8240 2374
rect 160 1360 8240 1432
rect 8280 1320 8306 2440
rect 8320 1360 8392 2480
rect 94 1294 8306 1320
<< nwell >>
rect 120 8840 8280 9960
rect 120 4200 8280 5320
rect 120 2760 8280 3880
rect 120 1320 8280 2440
<< pwell >>
rect -26 9974 8426 10106
rect -26 8826 106 9974
rect 8294 8826 8426 9974
rect -26 8694 8426 8826
rect -26 8026 106 8694
rect 8294 8026 8426 8694
rect -26 7894 8426 8026
rect -26 7466 106 7894
rect 294 7466 8106 7894
rect 8294 7466 8426 7894
rect -26 7174 8426 7466
rect -26 6746 106 7174
rect 294 6746 8106 7174
rect 8294 6746 8426 7174
rect -26 6614 8426 6746
rect -26 5466 106 6614
rect 8294 5466 8426 6614
rect -26 5334 8426 5466
rect -26 4186 106 5334
rect 8294 4186 8426 5334
rect -26 3894 8426 4186
rect -26 2746 106 3894
rect 8294 2746 8426 3894
rect -26 2454 8426 2746
rect -26 1306 106 2454
rect 8294 1306 8426 2454
rect -26 1174 8426 1306
rect 8294 666 8426 1174
rect -26 534 8426 666
rect -26 106 106 534
rect 294 106 8106 534
rect 8294 106 8426 534
rect -26 -26 8426 106
rect -26 -506 8426 -374
rect -26 -934 106 -506
rect 294 -934 8106 -506
rect 8294 -934 8426 -506
rect -26 -1066 8426 -934
<< mvnmos >>
rect 520 7520 2120 7720
rect 2440 7520 4040 7720
rect 4360 7520 5960 7720
rect 6280 7520 7880 7720
rect 520 6920 2120 7120
rect 2440 6920 4040 7120
rect 4360 6920 5960 7120
rect 6280 6920 7880 7120
rect 520 160 2120 360
rect 2440 160 4040 360
rect 4360 160 5960 360
rect 6280 160 7880 360
rect 520 -880 2120 -680
rect 2440 -880 4040 -680
rect 4360 -880 5960 -680
rect 6280 -880 7880 -680
<< mvpmos >>
rect 520 9160 2120 9760
rect 2440 9160 4040 9760
rect 4360 9160 5960 9760
rect 6280 9160 7880 9760
rect 520 4400 2120 5000
rect 2440 4400 4040 5000
rect 4360 4400 5960 5000
rect 6280 4400 7880 5000
rect 520 3080 2120 3680
rect 2440 3080 4040 3680
rect 4360 3080 5960 3680
rect 6280 3080 7880 3680
rect 520 1640 2120 2240
rect 2440 1640 4040 2240
rect 4360 1640 5960 2240
rect 6280 1640 7880 2240
<< mvndiff >>
rect 320 7671 520 7720
rect 320 7637 343 7671
rect 377 7637 520 7671
rect 320 7603 520 7637
rect 320 7569 343 7603
rect 377 7569 520 7603
rect 320 7520 520 7569
rect 2120 7671 2440 7720
rect 2120 7637 2263 7671
rect 2297 7637 2440 7671
rect 2120 7603 2440 7637
rect 2120 7569 2263 7603
rect 2297 7569 2440 7603
rect 2120 7520 2440 7569
rect 4040 7671 4360 7720
rect 4040 7637 4183 7671
rect 4217 7637 4360 7671
rect 4040 7603 4360 7637
rect 4040 7569 4183 7603
rect 4217 7569 4360 7603
rect 4040 7520 4360 7569
rect 5960 7671 6280 7720
rect 5960 7637 6103 7671
rect 6137 7637 6280 7671
rect 5960 7603 6280 7637
rect 5960 7569 6103 7603
rect 6137 7569 6280 7603
rect 5960 7520 6280 7569
rect 7880 7671 8080 7720
rect 7880 7637 8023 7671
rect 8057 7637 8080 7671
rect 7880 7603 8080 7637
rect 7880 7569 8023 7603
rect 8057 7569 8080 7603
rect 7880 7520 8080 7569
rect 320 7071 520 7120
rect 320 7037 343 7071
rect 377 7037 520 7071
rect 320 7003 520 7037
rect 320 6969 343 7003
rect 377 6969 520 7003
rect 320 6920 520 6969
rect 2120 7071 2440 7120
rect 2120 7037 2263 7071
rect 2297 7037 2440 7071
rect 2120 7003 2440 7037
rect 2120 6969 2263 7003
rect 2297 6969 2440 7003
rect 2120 6920 2440 6969
rect 4040 7071 4360 7120
rect 4040 7037 4183 7071
rect 4217 7037 4360 7071
rect 4040 7003 4360 7037
rect 4040 6969 4183 7003
rect 4217 6969 4360 7003
rect 4040 6920 4360 6969
rect 5960 7071 6280 7120
rect 5960 7037 6103 7071
rect 6137 7037 6280 7071
rect 5960 7003 6280 7037
rect 5960 6969 6103 7003
rect 6137 6969 6280 7003
rect 5960 6920 6280 6969
rect 7880 7071 8080 7120
rect 7880 7037 8023 7071
rect 8057 7037 8080 7071
rect 7880 7003 8080 7037
rect 7880 6969 8023 7003
rect 8057 6969 8080 7003
rect 7880 6920 8080 6969
rect 320 311 520 360
rect 320 277 343 311
rect 377 277 520 311
rect 320 243 520 277
rect 320 209 343 243
rect 377 209 520 243
rect 320 160 520 209
rect 2120 311 2440 360
rect 2120 277 2263 311
rect 2297 277 2440 311
rect 2120 243 2440 277
rect 2120 209 2263 243
rect 2297 209 2440 243
rect 2120 160 2440 209
rect 4040 311 4360 360
rect 4040 277 4183 311
rect 4217 277 4360 311
rect 4040 243 4360 277
rect 4040 209 4183 243
rect 4217 209 4360 243
rect 4040 160 4360 209
rect 5960 311 6280 360
rect 5960 277 6103 311
rect 6137 277 6280 311
rect 5960 243 6280 277
rect 5960 209 6103 243
rect 6137 209 6280 243
rect 5960 160 6280 209
rect 7880 311 8080 360
rect 7880 277 8023 311
rect 8057 277 8080 311
rect 7880 243 8080 277
rect 7880 209 8023 243
rect 8057 209 8080 243
rect 7880 160 8080 209
rect 320 -729 520 -680
rect 320 -763 343 -729
rect 377 -763 520 -729
rect 320 -797 520 -763
rect 320 -831 343 -797
rect 377 -831 520 -797
rect 320 -880 520 -831
rect 2120 -729 2440 -680
rect 2120 -763 2263 -729
rect 2297 -763 2440 -729
rect 2120 -797 2440 -763
rect 2120 -831 2263 -797
rect 2297 -831 2440 -797
rect 2120 -880 2440 -831
rect 4040 -729 4360 -680
rect 4040 -763 4183 -729
rect 4217 -763 4360 -729
rect 4040 -797 4360 -763
rect 4040 -831 4183 -797
rect 4217 -831 4360 -797
rect 4040 -880 4360 -831
rect 5960 -729 6280 -680
rect 5960 -763 6103 -729
rect 6137 -763 6280 -729
rect 5960 -797 6280 -763
rect 5960 -831 6103 -797
rect 6137 -831 6280 -797
rect 5960 -880 6280 -831
rect 7880 -729 8080 -680
rect 7880 -763 8023 -729
rect 8057 -763 8080 -729
rect 7880 -797 8080 -763
rect 7880 -831 8023 -797
rect 8057 -831 8080 -797
rect 7880 -880 8080 -831
<< mvpdiff >>
rect 320 9715 520 9760
rect 320 9681 343 9715
rect 377 9681 520 9715
rect 320 9647 520 9681
rect 320 9613 343 9647
rect 377 9613 520 9647
rect 320 9579 520 9613
rect 320 9545 343 9579
rect 377 9545 520 9579
rect 320 9511 520 9545
rect 320 9477 343 9511
rect 377 9477 520 9511
rect 320 9443 520 9477
rect 320 9409 343 9443
rect 377 9409 520 9443
rect 320 9375 520 9409
rect 320 9341 343 9375
rect 377 9341 520 9375
rect 320 9307 520 9341
rect 320 9273 343 9307
rect 377 9273 520 9307
rect 320 9239 520 9273
rect 320 9205 343 9239
rect 377 9205 520 9239
rect 320 9160 520 9205
rect 2120 9715 2440 9760
rect 2120 9681 2263 9715
rect 2297 9681 2440 9715
rect 2120 9647 2440 9681
rect 2120 9613 2263 9647
rect 2297 9613 2440 9647
rect 2120 9579 2440 9613
rect 2120 9545 2263 9579
rect 2297 9545 2440 9579
rect 2120 9511 2440 9545
rect 2120 9477 2263 9511
rect 2297 9477 2440 9511
rect 2120 9443 2440 9477
rect 2120 9409 2263 9443
rect 2297 9409 2440 9443
rect 2120 9375 2440 9409
rect 2120 9341 2263 9375
rect 2297 9341 2440 9375
rect 2120 9307 2440 9341
rect 2120 9273 2263 9307
rect 2297 9273 2440 9307
rect 2120 9239 2440 9273
rect 2120 9205 2263 9239
rect 2297 9205 2440 9239
rect 2120 9160 2440 9205
rect 4040 9715 4360 9760
rect 4040 9681 4183 9715
rect 4217 9681 4360 9715
rect 4040 9647 4360 9681
rect 4040 9613 4183 9647
rect 4217 9613 4360 9647
rect 4040 9579 4360 9613
rect 4040 9545 4183 9579
rect 4217 9545 4360 9579
rect 4040 9511 4360 9545
rect 4040 9477 4183 9511
rect 4217 9477 4360 9511
rect 4040 9443 4360 9477
rect 4040 9409 4183 9443
rect 4217 9409 4360 9443
rect 4040 9375 4360 9409
rect 4040 9341 4183 9375
rect 4217 9341 4360 9375
rect 4040 9307 4360 9341
rect 4040 9273 4183 9307
rect 4217 9273 4360 9307
rect 4040 9239 4360 9273
rect 4040 9205 4183 9239
rect 4217 9205 4360 9239
rect 4040 9160 4360 9205
rect 5960 9715 6280 9760
rect 5960 9681 6103 9715
rect 6137 9681 6280 9715
rect 5960 9647 6280 9681
rect 5960 9613 6103 9647
rect 6137 9613 6280 9647
rect 5960 9579 6280 9613
rect 5960 9545 6103 9579
rect 6137 9545 6280 9579
rect 5960 9511 6280 9545
rect 5960 9477 6103 9511
rect 6137 9477 6280 9511
rect 5960 9443 6280 9477
rect 5960 9409 6103 9443
rect 6137 9409 6280 9443
rect 5960 9375 6280 9409
rect 5960 9341 6103 9375
rect 6137 9341 6280 9375
rect 5960 9307 6280 9341
rect 5960 9273 6103 9307
rect 6137 9273 6280 9307
rect 5960 9239 6280 9273
rect 5960 9205 6103 9239
rect 6137 9205 6280 9239
rect 5960 9160 6280 9205
rect 7880 9715 8080 9760
rect 7880 9681 8023 9715
rect 8057 9681 8080 9715
rect 7880 9647 8080 9681
rect 7880 9613 8023 9647
rect 8057 9613 8080 9647
rect 7880 9579 8080 9613
rect 7880 9545 8023 9579
rect 8057 9545 8080 9579
rect 7880 9511 8080 9545
rect 7880 9477 8023 9511
rect 8057 9477 8080 9511
rect 7880 9443 8080 9477
rect 7880 9409 8023 9443
rect 8057 9409 8080 9443
rect 7880 9375 8080 9409
rect 7880 9341 8023 9375
rect 8057 9341 8080 9375
rect 7880 9307 8080 9341
rect 7880 9273 8023 9307
rect 8057 9273 8080 9307
rect 7880 9239 8080 9273
rect 7880 9205 8023 9239
rect 8057 9205 8080 9239
rect 7880 9160 8080 9205
rect 320 4955 520 5000
rect 320 4921 343 4955
rect 377 4921 520 4955
rect 320 4887 520 4921
rect 320 4853 343 4887
rect 377 4853 520 4887
rect 320 4819 520 4853
rect 320 4785 343 4819
rect 377 4785 520 4819
rect 320 4751 520 4785
rect 320 4717 343 4751
rect 377 4717 520 4751
rect 320 4683 520 4717
rect 320 4649 343 4683
rect 377 4649 520 4683
rect 320 4615 520 4649
rect 320 4581 343 4615
rect 377 4581 520 4615
rect 320 4547 520 4581
rect 320 4513 343 4547
rect 377 4513 520 4547
rect 320 4479 520 4513
rect 320 4445 343 4479
rect 377 4445 520 4479
rect 320 4400 520 4445
rect 2120 4955 2440 5000
rect 2120 4921 2263 4955
rect 2297 4921 2440 4955
rect 2120 4887 2440 4921
rect 2120 4853 2263 4887
rect 2297 4853 2440 4887
rect 2120 4819 2440 4853
rect 2120 4785 2263 4819
rect 2297 4785 2440 4819
rect 2120 4751 2440 4785
rect 2120 4717 2263 4751
rect 2297 4717 2440 4751
rect 2120 4683 2440 4717
rect 2120 4649 2263 4683
rect 2297 4649 2440 4683
rect 2120 4615 2440 4649
rect 2120 4581 2263 4615
rect 2297 4581 2440 4615
rect 2120 4547 2440 4581
rect 2120 4513 2263 4547
rect 2297 4513 2440 4547
rect 2120 4479 2440 4513
rect 2120 4445 2263 4479
rect 2297 4445 2440 4479
rect 2120 4400 2440 4445
rect 4040 4955 4360 5000
rect 4040 4921 4183 4955
rect 4217 4921 4360 4955
rect 4040 4887 4360 4921
rect 4040 4853 4183 4887
rect 4217 4853 4360 4887
rect 4040 4819 4360 4853
rect 4040 4785 4183 4819
rect 4217 4785 4360 4819
rect 4040 4751 4360 4785
rect 4040 4717 4183 4751
rect 4217 4717 4360 4751
rect 4040 4683 4360 4717
rect 4040 4649 4183 4683
rect 4217 4649 4360 4683
rect 4040 4615 4360 4649
rect 4040 4581 4183 4615
rect 4217 4581 4360 4615
rect 4040 4547 4360 4581
rect 4040 4513 4183 4547
rect 4217 4513 4360 4547
rect 4040 4479 4360 4513
rect 4040 4445 4183 4479
rect 4217 4445 4360 4479
rect 4040 4400 4360 4445
rect 5960 4955 6280 5000
rect 5960 4921 6103 4955
rect 6137 4921 6280 4955
rect 5960 4887 6280 4921
rect 5960 4853 6103 4887
rect 6137 4853 6280 4887
rect 5960 4819 6280 4853
rect 5960 4785 6103 4819
rect 6137 4785 6280 4819
rect 5960 4751 6280 4785
rect 5960 4717 6103 4751
rect 6137 4717 6280 4751
rect 5960 4683 6280 4717
rect 5960 4649 6103 4683
rect 6137 4649 6280 4683
rect 5960 4615 6280 4649
rect 5960 4581 6103 4615
rect 6137 4581 6280 4615
rect 5960 4547 6280 4581
rect 5960 4513 6103 4547
rect 6137 4513 6280 4547
rect 5960 4479 6280 4513
rect 5960 4445 6103 4479
rect 6137 4445 6280 4479
rect 5960 4400 6280 4445
rect 7880 4955 8080 5000
rect 7880 4921 8023 4955
rect 8057 4921 8080 4955
rect 7880 4887 8080 4921
rect 7880 4853 8023 4887
rect 8057 4853 8080 4887
rect 7880 4819 8080 4853
rect 7880 4785 8023 4819
rect 8057 4785 8080 4819
rect 7880 4751 8080 4785
rect 7880 4717 8023 4751
rect 8057 4717 8080 4751
rect 7880 4683 8080 4717
rect 7880 4649 8023 4683
rect 8057 4649 8080 4683
rect 7880 4615 8080 4649
rect 7880 4581 8023 4615
rect 8057 4581 8080 4615
rect 7880 4547 8080 4581
rect 7880 4513 8023 4547
rect 8057 4513 8080 4547
rect 7880 4479 8080 4513
rect 7880 4445 8023 4479
rect 8057 4445 8080 4479
rect 7880 4400 8080 4445
rect 320 3635 520 3680
rect 320 3601 343 3635
rect 377 3601 520 3635
rect 320 3567 520 3601
rect 320 3533 343 3567
rect 377 3533 520 3567
rect 320 3499 520 3533
rect 320 3465 343 3499
rect 377 3465 520 3499
rect 320 3431 520 3465
rect 320 3397 343 3431
rect 377 3397 520 3431
rect 320 3363 520 3397
rect 320 3329 343 3363
rect 377 3329 520 3363
rect 320 3295 520 3329
rect 320 3261 343 3295
rect 377 3261 520 3295
rect 320 3227 520 3261
rect 320 3193 343 3227
rect 377 3193 520 3227
rect 320 3159 520 3193
rect 320 3125 343 3159
rect 377 3125 520 3159
rect 320 3080 520 3125
rect 2120 3635 2440 3680
rect 2120 3601 2263 3635
rect 2297 3601 2440 3635
rect 2120 3567 2440 3601
rect 2120 3533 2263 3567
rect 2297 3533 2440 3567
rect 2120 3499 2440 3533
rect 2120 3465 2263 3499
rect 2297 3465 2440 3499
rect 2120 3431 2440 3465
rect 2120 3397 2263 3431
rect 2297 3397 2440 3431
rect 2120 3363 2440 3397
rect 2120 3329 2263 3363
rect 2297 3329 2440 3363
rect 2120 3295 2440 3329
rect 2120 3261 2263 3295
rect 2297 3261 2440 3295
rect 2120 3227 2440 3261
rect 2120 3193 2263 3227
rect 2297 3193 2440 3227
rect 2120 3159 2440 3193
rect 2120 3125 2263 3159
rect 2297 3125 2440 3159
rect 2120 3080 2440 3125
rect 4040 3635 4360 3680
rect 4040 3601 4183 3635
rect 4217 3601 4360 3635
rect 4040 3567 4360 3601
rect 4040 3533 4183 3567
rect 4217 3533 4360 3567
rect 4040 3499 4360 3533
rect 4040 3465 4183 3499
rect 4217 3465 4360 3499
rect 4040 3431 4360 3465
rect 4040 3397 4183 3431
rect 4217 3397 4360 3431
rect 4040 3363 4360 3397
rect 4040 3329 4183 3363
rect 4217 3329 4360 3363
rect 4040 3295 4360 3329
rect 4040 3261 4183 3295
rect 4217 3261 4360 3295
rect 4040 3227 4360 3261
rect 4040 3193 4183 3227
rect 4217 3193 4360 3227
rect 4040 3159 4360 3193
rect 4040 3125 4183 3159
rect 4217 3125 4360 3159
rect 4040 3080 4360 3125
rect 5960 3635 6280 3680
rect 5960 3601 6103 3635
rect 6137 3601 6280 3635
rect 5960 3567 6280 3601
rect 5960 3533 6103 3567
rect 6137 3533 6280 3567
rect 5960 3499 6280 3533
rect 5960 3465 6103 3499
rect 6137 3465 6280 3499
rect 5960 3431 6280 3465
rect 5960 3397 6103 3431
rect 6137 3397 6280 3431
rect 5960 3363 6280 3397
rect 5960 3329 6103 3363
rect 6137 3329 6280 3363
rect 5960 3295 6280 3329
rect 5960 3261 6103 3295
rect 6137 3261 6280 3295
rect 5960 3227 6280 3261
rect 5960 3193 6103 3227
rect 6137 3193 6280 3227
rect 5960 3159 6280 3193
rect 5960 3125 6103 3159
rect 6137 3125 6280 3159
rect 5960 3080 6280 3125
rect 7880 3635 8080 3680
rect 7880 3601 8023 3635
rect 8057 3601 8080 3635
rect 7880 3567 8080 3601
rect 7880 3533 8023 3567
rect 8057 3533 8080 3567
rect 7880 3499 8080 3533
rect 7880 3465 8023 3499
rect 8057 3465 8080 3499
rect 7880 3431 8080 3465
rect 7880 3397 8023 3431
rect 8057 3397 8080 3431
rect 7880 3363 8080 3397
rect 7880 3329 8023 3363
rect 8057 3329 8080 3363
rect 7880 3295 8080 3329
rect 7880 3261 8023 3295
rect 8057 3261 8080 3295
rect 7880 3227 8080 3261
rect 7880 3193 8023 3227
rect 8057 3193 8080 3227
rect 7880 3159 8080 3193
rect 7880 3125 8023 3159
rect 8057 3125 8080 3159
rect 7880 3080 8080 3125
rect 320 2195 520 2240
rect 320 2161 343 2195
rect 377 2161 520 2195
rect 320 2127 520 2161
rect 320 2093 343 2127
rect 377 2093 520 2127
rect 320 2059 520 2093
rect 320 2025 343 2059
rect 377 2025 520 2059
rect 320 1991 520 2025
rect 320 1957 343 1991
rect 377 1957 520 1991
rect 320 1923 520 1957
rect 320 1889 343 1923
rect 377 1889 520 1923
rect 320 1855 520 1889
rect 320 1821 343 1855
rect 377 1821 520 1855
rect 320 1787 520 1821
rect 320 1753 343 1787
rect 377 1753 520 1787
rect 320 1719 520 1753
rect 320 1685 343 1719
rect 377 1685 520 1719
rect 320 1640 520 1685
rect 2120 2195 2440 2240
rect 2120 2161 2263 2195
rect 2297 2161 2440 2195
rect 2120 2127 2440 2161
rect 2120 2093 2263 2127
rect 2297 2093 2440 2127
rect 2120 2059 2440 2093
rect 2120 2025 2263 2059
rect 2297 2025 2440 2059
rect 2120 1991 2440 2025
rect 2120 1957 2263 1991
rect 2297 1957 2440 1991
rect 2120 1923 2440 1957
rect 2120 1889 2263 1923
rect 2297 1889 2440 1923
rect 2120 1855 2440 1889
rect 2120 1821 2263 1855
rect 2297 1821 2440 1855
rect 2120 1787 2440 1821
rect 2120 1753 2263 1787
rect 2297 1753 2440 1787
rect 2120 1719 2440 1753
rect 2120 1685 2263 1719
rect 2297 1685 2440 1719
rect 2120 1640 2440 1685
rect 4040 2195 4360 2240
rect 4040 2161 4183 2195
rect 4217 2161 4360 2195
rect 4040 2127 4360 2161
rect 4040 2093 4183 2127
rect 4217 2093 4360 2127
rect 4040 2059 4360 2093
rect 4040 2025 4183 2059
rect 4217 2025 4360 2059
rect 4040 1991 4360 2025
rect 4040 1957 4183 1991
rect 4217 1957 4360 1991
rect 4040 1923 4360 1957
rect 4040 1889 4183 1923
rect 4217 1889 4360 1923
rect 4040 1855 4360 1889
rect 4040 1821 4183 1855
rect 4217 1821 4360 1855
rect 4040 1787 4360 1821
rect 4040 1753 4183 1787
rect 4217 1753 4360 1787
rect 4040 1719 4360 1753
rect 4040 1685 4183 1719
rect 4217 1685 4360 1719
rect 4040 1640 4360 1685
rect 5960 2195 6280 2240
rect 5960 2161 6103 2195
rect 6137 2161 6280 2195
rect 5960 2127 6280 2161
rect 5960 2093 6103 2127
rect 6137 2093 6280 2127
rect 5960 2059 6280 2093
rect 5960 2025 6103 2059
rect 6137 2025 6280 2059
rect 5960 1991 6280 2025
rect 5960 1957 6103 1991
rect 6137 1957 6280 1991
rect 5960 1923 6280 1957
rect 5960 1889 6103 1923
rect 6137 1889 6280 1923
rect 5960 1855 6280 1889
rect 5960 1821 6103 1855
rect 6137 1821 6280 1855
rect 5960 1787 6280 1821
rect 5960 1753 6103 1787
rect 6137 1753 6280 1787
rect 5960 1719 6280 1753
rect 5960 1685 6103 1719
rect 6137 1685 6280 1719
rect 5960 1640 6280 1685
rect 7880 2195 8080 2240
rect 7880 2161 8023 2195
rect 8057 2161 8080 2195
rect 7880 2127 8080 2161
rect 7880 2093 8023 2127
rect 8057 2093 8080 2127
rect 7880 2059 8080 2093
rect 7880 2025 8023 2059
rect 8057 2025 8080 2059
rect 7880 1991 8080 2025
rect 7880 1957 8023 1991
rect 8057 1957 8080 1991
rect 7880 1923 8080 1957
rect 7880 1889 8023 1923
rect 8057 1889 8080 1923
rect 7880 1855 8080 1889
rect 7880 1821 8023 1855
rect 8057 1821 8080 1855
rect 7880 1787 8080 1821
rect 7880 1753 8023 1787
rect 8057 1753 8080 1787
rect 7880 1719 8080 1753
rect 7880 1685 8023 1719
rect 8057 1685 8080 1719
rect 7880 1640 8080 1685
<< mvndiffc >>
rect 343 7637 377 7671
rect 343 7569 377 7603
rect 2263 7637 2297 7671
rect 2263 7569 2297 7603
rect 4183 7637 4217 7671
rect 4183 7569 4217 7603
rect 6103 7637 6137 7671
rect 6103 7569 6137 7603
rect 8023 7637 8057 7671
rect 8023 7569 8057 7603
rect 343 7037 377 7071
rect 343 6969 377 7003
rect 2263 7037 2297 7071
rect 2263 6969 2297 7003
rect 4183 7037 4217 7071
rect 4183 6969 4217 7003
rect 6103 7037 6137 7071
rect 6103 6969 6137 7003
rect 8023 7037 8057 7071
rect 8023 6969 8057 7003
rect 343 277 377 311
rect 343 209 377 243
rect 2263 277 2297 311
rect 2263 209 2297 243
rect 4183 277 4217 311
rect 4183 209 4217 243
rect 6103 277 6137 311
rect 6103 209 6137 243
rect 8023 277 8057 311
rect 8023 209 8057 243
rect 343 -763 377 -729
rect 343 -831 377 -797
rect 2263 -763 2297 -729
rect 2263 -831 2297 -797
rect 4183 -763 4217 -729
rect 4183 -831 4217 -797
rect 6103 -763 6137 -729
rect 6103 -831 6137 -797
rect 8023 -763 8057 -729
rect 8023 -831 8057 -797
<< mvpdiffc >>
rect 343 9681 377 9715
rect 343 9613 377 9647
rect 343 9545 377 9579
rect 343 9477 377 9511
rect 343 9409 377 9443
rect 343 9341 377 9375
rect 343 9273 377 9307
rect 343 9205 377 9239
rect 2263 9681 2297 9715
rect 2263 9613 2297 9647
rect 2263 9545 2297 9579
rect 2263 9477 2297 9511
rect 2263 9409 2297 9443
rect 2263 9341 2297 9375
rect 2263 9273 2297 9307
rect 2263 9205 2297 9239
rect 4183 9681 4217 9715
rect 4183 9613 4217 9647
rect 4183 9545 4217 9579
rect 4183 9477 4217 9511
rect 4183 9409 4217 9443
rect 4183 9341 4217 9375
rect 4183 9273 4217 9307
rect 4183 9205 4217 9239
rect 6103 9681 6137 9715
rect 6103 9613 6137 9647
rect 6103 9545 6137 9579
rect 6103 9477 6137 9511
rect 6103 9409 6137 9443
rect 6103 9341 6137 9375
rect 6103 9273 6137 9307
rect 6103 9205 6137 9239
rect 8023 9681 8057 9715
rect 8023 9613 8057 9647
rect 8023 9545 8057 9579
rect 8023 9477 8057 9511
rect 8023 9409 8057 9443
rect 8023 9341 8057 9375
rect 8023 9273 8057 9307
rect 8023 9205 8057 9239
rect 343 4921 377 4955
rect 343 4853 377 4887
rect 343 4785 377 4819
rect 343 4717 377 4751
rect 343 4649 377 4683
rect 343 4581 377 4615
rect 343 4513 377 4547
rect 343 4445 377 4479
rect 2263 4921 2297 4955
rect 2263 4853 2297 4887
rect 2263 4785 2297 4819
rect 2263 4717 2297 4751
rect 2263 4649 2297 4683
rect 2263 4581 2297 4615
rect 2263 4513 2297 4547
rect 2263 4445 2297 4479
rect 4183 4921 4217 4955
rect 4183 4853 4217 4887
rect 4183 4785 4217 4819
rect 4183 4717 4217 4751
rect 4183 4649 4217 4683
rect 4183 4581 4217 4615
rect 4183 4513 4217 4547
rect 4183 4445 4217 4479
rect 6103 4921 6137 4955
rect 6103 4853 6137 4887
rect 6103 4785 6137 4819
rect 6103 4717 6137 4751
rect 6103 4649 6137 4683
rect 6103 4581 6137 4615
rect 6103 4513 6137 4547
rect 6103 4445 6137 4479
rect 8023 4921 8057 4955
rect 8023 4853 8057 4887
rect 8023 4785 8057 4819
rect 8023 4717 8057 4751
rect 8023 4649 8057 4683
rect 8023 4581 8057 4615
rect 8023 4513 8057 4547
rect 8023 4445 8057 4479
rect 343 3601 377 3635
rect 343 3533 377 3567
rect 343 3465 377 3499
rect 343 3397 377 3431
rect 343 3329 377 3363
rect 343 3261 377 3295
rect 343 3193 377 3227
rect 343 3125 377 3159
rect 2263 3601 2297 3635
rect 2263 3533 2297 3567
rect 2263 3465 2297 3499
rect 2263 3397 2297 3431
rect 2263 3329 2297 3363
rect 2263 3261 2297 3295
rect 2263 3193 2297 3227
rect 2263 3125 2297 3159
rect 4183 3601 4217 3635
rect 4183 3533 4217 3567
rect 4183 3465 4217 3499
rect 4183 3397 4217 3431
rect 4183 3329 4217 3363
rect 4183 3261 4217 3295
rect 4183 3193 4217 3227
rect 4183 3125 4217 3159
rect 6103 3601 6137 3635
rect 6103 3533 6137 3567
rect 6103 3465 6137 3499
rect 6103 3397 6137 3431
rect 6103 3329 6137 3363
rect 6103 3261 6137 3295
rect 6103 3193 6137 3227
rect 6103 3125 6137 3159
rect 8023 3601 8057 3635
rect 8023 3533 8057 3567
rect 8023 3465 8057 3499
rect 8023 3397 8057 3431
rect 8023 3329 8057 3363
rect 8023 3261 8057 3295
rect 8023 3193 8057 3227
rect 8023 3125 8057 3159
rect 343 2161 377 2195
rect 343 2093 377 2127
rect 343 2025 377 2059
rect 343 1957 377 1991
rect 343 1889 377 1923
rect 343 1821 377 1855
rect 343 1753 377 1787
rect 343 1685 377 1719
rect 2263 2161 2297 2195
rect 2263 2093 2297 2127
rect 2263 2025 2297 2059
rect 2263 1957 2297 1991
rect 2263 1889 2297 1923
rect 2263 1821 2297 1855
rect 2263 1753 2297 1787
rect 2263 1685 2297 1719
rect 4183 2161 4217 2195
rect 4183 2093 4217 2127
rect 4183 2025 4217 2059
rect 4183 1957 4217 1991
rect 4183 1889 4217 1923
rect 4183 1821 4217 1855
rect 4183 1753 4217 1787
rect 4183 1685 4217 1719
rect 6103 2161 6137 2195
rect 6103 2093 6137 2127
rect 6103 2025 6137 2059
rect 6103 1957 6137 1991
rect 6103 1889 6137 1923
rect 6103 1821 6137 1855
rect 6103 1753 6137 1787
rect 6103 1685 6137 1719
rect 8023 2161 8057 2195
rect 8023 2093 8057 2127
rect 8023 2025 8057 2059
rect 8023 1957 8057 1991
rect 8023 1889 8057 1923
rect 8023 1821 8057 1855
rect 8023 1753 8057 1787
rect 8023 1685 8057 1719
<< psubdiff >>
rect 0 10057 8400 10080
rect 0 10023 137 10057
rect 171 10023 205 10057
rect 239 10023 273 10057
rect 307 10023 341 10057
rect 375 10023 409 10057
rect 443 10023 477 10057
rect 511 10023 545 10057
rect 579 10023 613 10057
rect 647 10023 681 10057
rect 715 10023 749 10057
rect 783 10023 817 10057
rect 851 10023 885 10057
rect 919 10023 953 10057
rect 987 10023 1021 10057
rect 1055 10023 1089 10057
rect 1123 10023 1157 10057
rect 1191 10023 1225 10057
rect 1259 10023 1293 10057
rect 1327 10023 1361 10057
rect 1395 10023 1429 10057
rect 1463 10023 1497 10057
rect 1531 10023 1565 10057
rect 1599 10023 1633 10057
rect 1667 10023 1701 10057
rect 1735 10023 1769 10057
rect 1803 10023 1837 10057
rect 1871 10023 1905 10057
rect 1939 10023 1973 10057
rect 2007 10023 2041 10057
rect 2075 10023 2109 10057
rect 2143 10023 2177 10057
rect 2211 10023 2245 10057
rect 2279 10023 2313 10057
rect 2347 10023 2381 10057
rect 2415 10023 2449 10057
rect 2483 10023 2517 10057
rect 2551 10023 2585 10057
rect 2619 10023 2653 10057
rect 2687 10023 2721 10057
rect 2755 10023 2789 10057
rect 2823 10023 2857 10057
rect 2891 10023 2925 10057
rect 2959 10023 2993 10057
rect 3027 10023 3061 10057
rect 3095 10023 3129 10057
rect 3163 10023 3197 10057
rect 3231 10023 3265 10057
rect 3299 10023 3333 10057
rect 3367 10023 3401 10057
rect 3435 10023 3469 10057
rect 3503 10023 3537 10057
rect 3571 10023 3605 10057
rect 3639 10023 3673 10057
rect 3707 10023 3741 10057
rect 3775 10023 3809 10057
rect 3843 10023 3877 10057
rect 3911 10023 3945 10057
rect 3979 10023 4013 10057
rect 4047 10023 4081 10057
rect 4115 10023 4149 10057
rect 4183 10023 4217 10057
rect 4251 10023 4285 10057
rect 4319 10023 4353 10057
rect 4387 10023 4421 10057
rect 4455 10023 4489 10057
rect 4523 10023 4557 10057
rect 4591 10023 4625 10057
rect 4659 10023 4693 10057
rect 4727 10023 4761 10057
rect 4795 10023 4829 10057
rect 4863 10023 4897 10057
rect 4931 10023 4965 10057
rect 4999 10023 5033 10057
rect 5067 10023 5101 10057
rect 5135 10023 5169 10057
rect 5203 10023 5237 10057
rect 5271 10023 5305 10057
rect 5339 10023 5373 10057
rect 5407 10023 5441 10057
rect 5475 10023 5509 10057
rect 5543 10023 5577 10057
rect 5611 10023 5645 10057
rect 5679 10023 5713 10057
rect 5747 10023 5781 10057
rect 5815 10023 5849 10057
rect 5883 10023 5917 10057
rect 5951 10023 5985 10057
rect 6019 10023 6053 10057
rect 6087 10023 6121 10057
rect 6155 10023 6189 10057
rect 6223 10023 6257 10057
rect 6291 10023 6325 10057
rect 6359 10023 6393 10057
rect 6427 10023 6461 10057
rect 6495 10023 6529 10057
rect 6563 10023 6597 10057
rect 6631 10023 6665 10057
rect 6699 10023 6733 10057
rect 6767 10023 6801 10057
rect 6835 10023 6869 10057
rect 6903 10023 6937 10057
rect 6971 10023 7005 10057
rect 7039 10023 7073 10057
rect 7107 10023 7141 10057
rect 7175 10023 7209 10057
rect 7243 10023 7277 10057
rect 7311 10023 7345 10057
rect 7379 10023 7413 10057
rect 7447 10023 7481 10057
rect 7515 10023 7549 10057
rect 7583 10023 7617 10057
rect 7651 10023 7685 10057
rect 7719 10023 7753 10057
rect 7787 10023 7821 10057
rect 7855 10023 7889 10057
rect 7923 10023 7957 10057
rect 7991 10023 8025 10057
rect 8059 10023 8093 10057
rect 8127 10023 8161 10057
rect 8195 10023 8229 10057
rect 8263 10023 8400 10057
rect 0 10000 8400 10023
rect 0 9927 80 10000
rect 0 9893 23 9927
rect 57 9893 80 9927
rect 8320 9927 8400 10000
rect 0 9859 80 9893
rect 0 9825 23 9859
rect 57 9825 80 9859
rect 0 9791 80 9825
rect 0 9757 23 9791
rect 57 9757 80 9791
rect 0 9723 80 9757
rect 0 9689 23 9723
rect 57 9689 80 9723
rect 0 9655 80 9689
rect 0 9621 23 9655
rect 57 9621 80 9655
rect 0 9587 80 9621
rect 0 9553 23 9587
rect 57 9553 80 9587
rect 0 9519 80 9553
rect 0 9485 23 9519
rect 57 9485 80 9519
rect 0 9451 80 9485
rect 0 9417 23 9451
rect 57 9417 80 9451
rect 0 9383 80 9417
rect 0 9349 23 9383
rect 57 9349 80 9383
rect 0 9315 80 9349
rect 0 9281 23 9315
rect 57 9281 80 9315
rect 0 9247 80 9281
rect 0 9213 23 9247
rect 57 9213 80 9247
rect 0 9179 80 9213
rect 0 9145 23 9179
rect 57 9145 80 9179
rect 0 9111 80 9145
rect 0 9077 23 9111
rect 57 9077 80 9111
rect 0 9043 80 9077
rect 0 9009 23 9043
rect 57 9009 80 9043
rect 0 8975 80 9009
rect 0 8941 23 8975
rect 57 8941 80 8975
rect 0 8907 80 8941
rect 0 8873 23 8907
rect 57 8873 80 8907
rect 8320 9893 8343 9927
rect 8377 9893 8400 9927
rect 8320 9859 8400 9893
rect 8320 9825 8343 9859
rect 8377 9825 8400 9859
rect 8320 9791 8400 9825
rect 8320 9757 8343 9791
rect 8377 9757 8400 9791
rect 8320 9723 8400 9757
rect 8320 9689 8343 9723
rect 8377 9689 8400 9723
rect 8320 9655 8400 9689
rect 8320 9621 8343 9655
rect 8377 9621 8400 9655
rect 8320 9587 8400 9621
rect 8320 9553 8343 9587
rect 8377 9553 8400 9587
rect 8320 9519 8400 9553
rect 8320 9485 8343 9519
rect 8377 9485 8400 9519
rect 8320 9451 8400 9485
rect 8320 9417 8343 9451
rect 8377 9417 8400 9451
rect 8320 9383 8400 9417
rect 8320 9349 8343 9383
rect 8377 9349 8400 9383
rect 8320 9315 8400 9349
rect 8320 9281 8343 9315
rect 8377 9281 8400 9315
rect 8320 9247 8400 9281
rect 8320 9213 8343 9247
rect 8377 9213 8400 9247
rect 8320 9179 8400 9213
rect 8320 9145 8343 9179
rect 8377 9145 8400 9179
rect 8320 9111 8400 9145
rect 8320 9077 8343 9111
rect 8377 9077 8400 9111
rect 8320 9043 8400 9077
rect 8320 9009 8343 9043
rect 8377 9009 8400 9043
rect 8320 8975 8400 9009
rect 8320 8941 8343 8975
rect 8377 8941 8400 8975
rect 8320 8907 8400 8941
rect 0 8800 80 8873
rect 8320 8873 8343 8907
rect 8377 8873 8400 8907
rect 8320 8800 8400 8873
rect 0 8777 8400 8800
rect 0 8743 137 8777
rect 171 8743 205 8777
rect 239 8743 273 8777
rect 307 8743 341 8777
rect 375 8743 409 8777
rect 443 8743 477 8777
rect 511 8743 545 8777
rect 579 8743 613 8777
rect 647 8743 681 8777
rect 715 8743 749 8777
rect 783 8743 817 8777
rect 851 8743 885 8777
rect 919 8743 953 8777
rect 987 8743 1021 8777
rect 1055 8743 1089 8777
rect 1123 8743 1157 8777
rect 1191 8743 1225 8777
rect 1259 8743 1293 8777
rect 1327 8743 1361 8777
rect 1395 8743 1429 8777
rect 1463 8743 1497 8777
rect 1531 8743 1565 8777
rect 1599 8743 1633 8777
rect 1667 8743 1701 8777
rect 1735 8743 1769 8777
rect 1803 8743 1837 8777
rect 1871 8743 1905 8777
rect 1939 8743 1973 8777
rect 2007 8743 2041 8777
rect 2075 8743 2109 8777
rect 2143 8743 2177 8777
rect 2211 8743 2245 8777
rect 2279 8743 2313 8777
rect 2347 8743 2381 8777
rect 2415 8743 2449 8777
rect 2483 8743 2517 8777
rect 2551 8743 2585 8777
rect 2619 8743 2653 8777
rect 2687 8743 2721 8777
rect 2755 8743 2789 8777
rect 2823 8743 2857 8777
rect 2891 8743 2925 8777
rect 2959 8743 2993 8777
rect 3027 8743 3061 8777
rect 3095 8743 3129 8777
rect 3163 8743 3197 8777
rect 3231 8743 3265 8777
rect 3299 8743 3333 8777
rect 3367 8743 3401 8777
rect 3435 8743 3469 8777
rect 3503 8743 3537 8777
rect 3571 8743 3605 8777
rect 3639 8743 3673 8777
rect 3707 8743 3741 8777
rect 3775 8743 3809 8777
rect 3843 8743 3877 8777
rect 3911 8743 3945 8777
rect 3979 8743 4013 8777
rect 4047 8743 4081 8777
rect 4115 8743 4149 8777
rect 4183 8743 4217 8777
rect 4251 8743 4285 8777
rect 4319 8743 4353 8777
rect 4387 8743 4421 8777
rect 4455 8743 4489 8777
rect 4523 8743 4557 8777
rect 4591 8743 4625 8777
rect 4659 8743 4693 8777
rect 4727 8743 4761 8777
rect 4795 8743 4829 8777
rect 4863 8743 4897 8777
rect 4931 8743 4965 8777
rect 4999 8743 5033 8777
rect 5067 8743 5101 8777
rect 5135 8743 5169 8777
rect 5203 8743 5237 8777
rect 5271 8743 5305 8777
rect 5339 8743 5373 8777
rect 5407 8743 5441 8777
rect 5475 8743 5509 8777
rect 5543 8743 5577 8777
rect 5611 8743 5645 8777
rect 5679 8743 5713 8777
rect 5747 8743 5781 8777
rect 5815 8743 5849 8777
rect 5883 8743 5917 8777
rect 5951 8743 5985 8777
rect 6019 8743 6053 8777
rect 6087 8743 6121 8777
rect 6155 8743 6189 8777
rect 6223 8743 6257 8777
rect 6291 8743 6325 8777
rect 6359 8743 6393 8777
rect 6427 8743 6461 8777
rect 6495 8743 6529 8777
rect 6563 8743 6597 8777
rect 6631 8743 6665 8777
rect 6699 8743 6733 8777
rect 6767 8743 6801 8777
rect 6835 8743 6869 8777
rect 6903 8743 6937 8777
rect 6971 8743 7005 8777
rect 7039 8743 7073 8777
rect 7107 8743 7141 8777
rect 7175 8743 7209 8777
rect 7243 8743 7277 8777
rect 7311 8743 7345 8777
rect 7379 8743 7413 8777
rect 7447 8743 7481 8777
rect 7515 8743 7549 8777
rect 7583 8743 7617 8777
rect 7651 8743 7685 8777
rect 7719 8743 7753 8777
rect 7787 8743 7821 8777
rect 7855 8743 7889 8777
rect 7923 8743 7957 8777
rect 7991 8743 8025 8777
rect 8059 8743 8093 8777
rect 8127 8743 8161 8777
rect 8195 8743 8229 8777
rect 8263 8743 8400 8777
rect 0 8720 8400 8743
rect 0 8000 80 8720
rect 8320 8000 8400 8720
rect 0 7977 8400 8000
rect 0 7943 137 7977
rect 171 7943 205 7977
rect 239 7943 273 7977
rect 307 7943 341 7977
rect 375 7943 409 7977
rect 443 7943 477 7977
rect 511 7943 545 7977
rect 579 7943 613 7977
rect 647 7943 681 7977
rect 715 7943 749 7977
rect 783 7943 817 7977
rect 851 7943 885 7977
rect 919 7943 953 7977
rect 987 7943 1021 7977
rect 1055 7943 1089 7977
rect 1123 7943 1157 7977
rect 1191 7943 1225 7977
rect 1259 7943 1293 7977
rect 1327 7943 1361 7977
rect 1395 7943 1429 7977
rect 1463 7943 1497 7977
rect 1531 7943 1565 7977
rect 1599 7943 1633 7977
rect 1667 7943 1701 7977
rect 1735 7943 1769 7977
rect 1803 7943 1837 7977
rect 1871 7943 1905 7977
rect 1939 7943 1973 7977
rect 2007 7943 2041 7977
rect 2075 7943 2109 7977
rect 2143 7943 2177 7977
rect 2211 7943 2245 7977
rect 2279 7943 2313 7977
rect 2347 7943 2381 7977
rect 2415 7943 2449 7977
rect 2483 7943 2517 7977
rect 2551 7943 2585 7977
rect 2619 7943 2653 7977
rect 2687 7943 2721 7977
rect 2755 7943 2789 7977
rect 2823 7943 2857 7977
rect 2891 7943 2925 7977
rect 2959 7943 2993 7977
rect 3027 7943 3061 7977
rect 3095 7943 3129 7977
rect 3163 7943 3197 7977
rect 3231 7943 3265 7977
rect 3299 7943 3333 7977
rect 3367 7943 3401 7977
rect 3435 7943 3469 7977
rect 3503 7943 3537 7977
rect 3571 7943 3605 7977
rect 3639 7943 3673 7977
rect 3707 7943 3741 7977
rect 3775 7943 3809 7977
rect 3843 7943 3877 7977
rect 3911 7943 3945 7977
rect 3979 7943 4013 7977
rect 4047 7943 4081 7977
rect 4115 7943 4149 7977
rect 4183 7943 4217 7977
rect 4251 7943 4285 7977
rect 4319 7943 4353 7977
rect 4387 7943 4421 7977
rect 4455 7943 4489 7977
rect 4523 7943 4557 7977
rect 4591 7943 4625 7977
rect 4659 7943 4693 7977
rect 4727 7943 4761 7977
rect 4795 7943 4829 7977
rect 4863 7943 4897 7977
rect 4931 7943 4965 7977
rect 4999 7943 5033 7977
rect 5067 7943 5101 7977
rect 5135 7943 5169 7977
rect 5203 7943 5237 7977
rect 5271 7943 5305 7977
rect 5339 7943 5373 7977
rect 5407 7943 5441 7977
rect 5475 7943 5509 7977
rect 5543 7943 5577 7977
rect 5611 7943 5645 7977
rect 5679 7943 5713 7977
rect 5747 7943 5781 7977
rect 5815 7943 5849 7977
rect 5883 7943 5917 7977
rect 5951 7943 5985 7977
rect 6019 7943 6053 7977
rect 6087 7943 6121 7977
rect 6155 7943 6189 7977
rect 6223 7943 6257 7977
rect 6291 7943 6325 7977
rect 6359 7943 6393 7977
rect 6427 7943 6461 7977
rect 6495 7943 6529 7977
rect 6563 7943 6597 7977
rect 6631 7943 6665 7977
rect 6699 7943 6733 7977
rect 6767 7943 6801 7977
rect 6835 7943 6869 7977
rect 6903 7943 6937 7977
rect 6971 7943 7005 7977
rect 7039 7943 7073 7977
rect 7107 7943 7141 7977
rect 7175 7943 7209 7977
rect 7243 7943 7277 7977
rect 7311 7943 7345 7977
rect 7379 7943 7413 7977
rect 7447 7943 7481 7977
rect 7515 7943 7549 7977
rect 7583 7943 7617 7977
rect 7651 7943 7685 7977
rect 7719 7943 7753 7977
rect 7787 7943 7821 7977
rect 7855 7943 7889 7977
rect 7923 7943 7957 7977
rect 7991 7943 8025 7977
rect 8059 7943 8093 7977
rect 8127 7943 8161 7977
rect 8195 7943 8229 7977
rect 8263 7943 8400 7977
rect 0 7920 8400 7943
rect 0 7867 80 7920
rect 0 7833 23 7867
rect 57 7833 80 7867
rect 0 7799 80 7833
rect 0 7765 23 7799
rect 57 7765 80 7799
rect 0 7731 80 7765
rect 0 7697 23 7731
rect 57 7697 80 7731
rect 0 7663 80 7697
rect 0 7629 23 7663
rect 57 7629 80 7663
rect 0 7595 80 7629
rect 0 7561 23 7595
rect 57 7561 80 7595
rect 0 7527 80 7561
rect 0 7493 23 7527
rect 57 7493 80 7527
rect 0 7440 80 7493
rect 8320 7440 8400 7920
rect 0 7417 8400 7440
rect 0 7383 137 7417
rect 171 7383 205 7417
rect 239 7383 273 7417
rect 307 7383 341 7417
rect 375 7383 409 7417
rect 443 7383 477 7417
rect 511 7383 545 7417
rect 579 7383 613 7417
rect 647 7383 681 7417
rect 715 7383 749 7417
rect 783 7383 817 7417
rect 851 7383 885 7417
rect 919 7383 953 7417
rect 987 7383 1021 7417
rect 1055 7383 1089 7417
rect 1123 7383 1157 7417
rect 1191 7383 1225 7417
rect 1259 7383 1293 7417
rect 1327 7383 1361 7417
rect 1395 7383 1429 7417
rect 1463 7383 1497 7417
rect 1531 7383 1565 7417
rect 1599 7383 1633 7417
rect 1667 7383 1701 7417
rect 1735 7383 1769 7417
rect 1803 7383 1837 7417
rect 1871 7383 1905 7417
rect 1939 7383 1973 7417
rect 2007 7383 2041 7417
rect 2075 7383 2109 7417
rect 2143 7383 2177 7417
rect 2211 7383 2245 7417
rect 2279 7383 2313 7417
rect 2347 7383 2381 7417
rect 2415 7383 2449 7417
rect 2483 7383 2517 7417
rect 2551 7383 2585 7417
rect 2619 7383 2653 7417
rect 2687 7383 2721 7417
rect 2755 7383 2789 7417
rect 2823 7383 2857 7417
rect 2891 7383 2925 7417
rect 2959 7383 2993 7417
rect 3027 7383 3061 7417
rect 3095 7383 3129 7417
rect 3163 7383 3197 7417
rect 3231 7383 3265 7417
rect 3299 7383 3333 7417
rect 3367 7383 3401 7417
rect 3435 7383 3469 7417
rect 3503 7383 3537 7417
rect 3571 7383 3605 7417
rect 3639 7383 3673 7417
rect 3707 7383 3741 7417
rect 3775 7383 3809 7417
rect 3843 7383 3877 7417
rect 3911 7383 3945 7417
rect 3979 7383 4013 7417
rect 4047 7383 4081 7417
rect 4115 7383 4149 7417
rect 4183 7383 4217 7417
rect 4251 7383 4285 7417
rect 4319 7383 4353 7417
rect 4387 7383 4421 7417
rect 4455 7383 4489 7417
rect 4523 7383 4557 7417
rect 4591 7383 4625 7417
rect 4659 7383 4693 7417
rect 4727 7383 4761 7417
rect 4795 7383 4829 7417
rect 4863 7383 4897 7417
rect 4931 7383 4965 7417
rect 4999 7383 5033 7417
rect 5067 7383 5101 7417
rect 5135 7383 5169 7417
rect 5203 7383 5237 7417
rect 5271 7383 5305 7417
rect 5339 7383 5373 7417
rect 5407 7383 5441 7417
rect 5475 7383 5509 7417
rect 5543 7383 5577 7417
rect 5611 7383 5645 7417
rect 5679 7383 5713 7417
rect 5747 7383 5781 7417
rect 5815 7383 5849 7417
rect 5883 7383 5917 7417
rect 5951 7383 5985 7417
rect 6019 7383 6053 7417
rect 6087 7383 6121 7417
rect 6155 7383 6189 7417
rect 6223 7383 6257 7417
rect 6291 7383 6325 7417
rect 6359 7383 6393 7417
rect 6427 7383 6461 7417
rect 6495 7383 6529 7417
rect 6563 7383 6597 7417
rect 6631 7383 6665 7417
rect 6699 7383 6733 7417
rect 6767 7383 6801 7417
rect 6835 7383 6869 7417
rect 6903 7383 6937 7417
rect 6971 7383 7005 7417
rect 7039 7383 7073 7417
rect 7107 7383 7141 7417
rect 7175 7383 7209 7417
rect 7243 7383 7277 7417
rect 7311 7383 7345 7417
rect 7379 7383 7413 7417
rect 7447 7383 7481 7417
rect 7515 7383 7549 7417
rect 7583 7383 7617 7417
rect 7651 7383 7685 7417
rect 7719 7383 7753 7417
rect 7787 7383 7821 7417
rect 7855 7383 7889 7417
rect 7923 7383 7957 7417
rect 7991 7383 8025 7417
rect 8059 7383 8093 7417
rect 8127 7383 8161 7417
rect 8195 7383 8229 7417
rect 8263 7383 8400 7417
rect 0 7360 8400 7383
rect 0 7257 8400 7280
rect 0 7223 137 7257
rect 171 7223 205 7257
rect 239 7223 273 7257
rect 307 7223 341 7257
rect 375 7223 409 7257
rect 443 7223 477 7257
rect 511 7223 545 7257
rect 579 7223 613 7257
rect 647 7223 681 7257
rect 715 7223 749 7257
rect 783 7223 817 7257
rect 851 7223 885 7257
rect 919 7223 953 7257
rect 987 7223 1021 7257
rect 1055 7223 1089 7257
rect 1123 7223 1157 7257
rect 1191 7223 1225 7257
rect 1259 7223 1293 7257
rect 1327 7223 1361 7257
rect 1395 7223 1429 7257
rect 1463 7223 1497 7257
rect 1531 7223 1565 7257
rect 1599 7223 1633 7257
rect 1667 7223 1701 7257
rect 1735 7223 1769 7257
rect 1803 7223 1837 7257
rect 1871 7223 1905 7257
rect 1939 7223 1973 7257
rect 2007 7223 2041 7257
rect 2075 7223 2109 7257
rect 2143 7223 2177 7257
rect 2211 7223 2245 7257
rect 2279 7223 2313 7257
rect 2347 7223 2381 7257
rect 2415 7223 2449 7257
rect 2483 7223 2517 7257
rect 2551 7223 2585 7257
rect 2619 7223 2653 7257
rect 2687 7223 2721 7257
rect 2755 7223 2789 7257
rect 2823 7223 2857 7257
rect 2891 7223 2925 7257
rect 2959 7223 2993 7257
rect 3027 7223 3061 7257
rect 3095 7223 3129 7257
rect 3163 7223 3197 7257
rect 3231 7223 3265 7257
rect 3299 7223 3333 7257
rect 3367 7223 3401 7257
rect 3435 7223 3469 7257
rect 3503 7223 3537 7257
rect 3571 7223 3605 7257
rect 3639 7223 3673 7257
rect 3707 7223 3741 7257
rect 3775 7223 3809 7257
rect 3843 7223 3877 7257
rect 3911 7223 3945 7257
rect 3979 7223 4013 7257
rect 4047 7223 4081 7257
rect 4115 7223 4149 7257
rect 4183 7223 4217 7257
rect 4251 7223 4285 7257
rect 4319 7223 4353 7257
rect 4387 7223 4421 7257
rect 4455 7223 4489 7257
rect 4523 7223 4557 7257
rect 4591 7223 4625 7257
rect 4659 7223 4693 7257
rect 4727 7223 4761 7257
rect 4795 7223 4829 7257
rect 4863 7223 4897 7257
rect 4931 7223 4965 7257
rect 4999 7223 5033 7257
rect 5067 7223 5101 7257
rect 5135 7223 5169 7257
rect 5203 7223 5237 7257
rect 5271 7223 5305 7257
rect 5339 7223 5373 7257
rect 5407 7223 5441 7257
rect 5475 7223 5509 7257
rect 5543 7223 5577 7257
rect 5611 7223 5645 7257
rect 5679 7223 5713 7257
rect 5747 7223 5781 7257
rect 5815 7223 5849 7257
rect 5883 7223 5917 7257
rect 5951 7223 5985 7257
rect 6019 7223 6053 7257
rect 6087 7223 6121 7257
rect 6155 7223 6189 7257
rect 6223 7223 6257 7257
rect 6291 7223 6325 7257
rect 6359 7223 6393 7257
rect 6427 7223 6461 7257
rect 6495 7223 6529 7257
rect 6563 7223 6597 7257
rect 6631 7223 6665 7257
rect 6699 7223 6733 7257
rect 6767 7223 6801 7257
rect 6835 7223 6869 7257
rect 6903 7223 6937 7257
rect 6971 7223 7005 7257
rect 7039 7223 7073 7257
rect 7107 7223 7141 7257
rect 7175 7223 7209 7257
rect 7243 7223 7277 7257
rect 7311 7223 7345 7257
rect 7379 7223 7413 7257
rect 7447 7223 7481 7257
rect 7515 7223 7549 7257
rect 7583 7223 7617 7257
rect 7651 7223 7685 7257
rect 7719 7223 7753 7257
rect 7787 7223 7821 7257
rect 7855 7223 7889 7257
rect 7923 7223 7957 7257
rect 7991 7223 8025 7257
rect 8059 7223 8093 7257
rect 8127 7223 8161 7257
rect 8195 7223 8229 7257
rect 8263 7223 8400 7257
rect 0 7200 8400 7223
rect 0 7147 80 7200
rect 0 7113 23 7147
rect 57 7113 80 7147
rect 0 7079 80 7113
rect 0 7045 23 7079
rect 57 7045 80 7079
rect 0 7011 80 7045
rect 0 6977 23 7011
rect 57 6977 80 7011
rect 0 6943 80 6977
rect 0 6909 23 6943
rect 57 6909 80 6943
rect 0 6875 80 6909
rect 0 6841 23 6875
rect 57 6841 80 6875
rect 0 6807 80 6841
rect 0 6773 23 6807
rect 57 6773 80 6807
rect 0 6720 80 6773
rect 8320 6720 8400 7200
rect 0 6697 8400 6720
rect 0 6663 137 6697
rect 171 6663 205 6697
rect 239 6663 273 6697
rect 307 6663 341 6697
rect 375 6663 409 6697
rect 443 6663 477 6697
rect 511 6663 545 6697
rect 579 6663 613 6697
rect 647 6663 681 6697
rect 715 6663 749 6697
rect 783 6663 817 6697
rect 851 6663 885 6697
rect 919 6663 953 6697
rect 987 6663 1021 6697
rect 1055 6663 1089 6697
rect 1123 6663 1157 6697
rect 1191 6663 1225 6697
rect 1259 6663 1293 6697
rect 1327 6663 1361 6697
rect 1395 6663 1429 6697
rect 1463 6663 1497 6697
rect 1531 6663 1565 6697
rect 1599 6663 1633 6697
rect 1667 6663 1701 6697
rect 1735 6663 1769 6697
rect 1803 6663 1837 6697
rect 1871 6663 1905 6697
rect 1939 6663 1973 6697
rect 2007 6663 2041 6697
rect 2075 6663 2109 6697
rect 2143 6663 2177 6697
rect 2211 6663 2245 6697
rect 2279 6663 2313 6697
rect 2347 6663 2381 6697
rect 2415 6663 2449 6697
rect 2483 6663 2517 6697
rect 2551 6663 2585 6697
rect 2619 6663 2653 6697
rect 2687 6663 2721 6697
rect 2755 6663 2789 6697
rect 2823 6663 2857 6697
rect 2891 6663 2925 6697
rect 2959 6663 2993 6697
rect 3027 6663 3061 6697
rect 3095 6663 3129 6697
rect 3163 6663 3197 6697
rect 3231 6663 3265 6697
rect 3299 6663 3333 6697
rect 3367 6663 3401 6697
rect 3435 6663 3469 6697
rect 3503 6663 3537 6697
rect 3571 6663 3605 6697
rect 3639 6663 3673 6697
rect 3707 6663 3741 6697
rect 3775 6663 3809 6697
rect 3843 6663 3877 6697
rect 3911 6663 3945 6697
rect 3979 6663 4013 6697
rect 4047 6663 4081 6697
rect 4115 6663 4149 6697
rect 4183 6663 4217 6697
rect 4251 6663 4285 6697
rect 4319 6663 4353 6697
rect 4387 6663 4421 6697
rect 4455 6663 4489 6697
rect 4523 6663 4557 6697
rect 4591 6663 4625 6697
rect 4659 6663 4693 6697
rect 4727 6663 4761 6697
rect 4795 6663 4829 6697
rect 4863 6663 4897 6697
rect 4931 6663 4965 6697
rect 4999 6663 5033 6697
rect 5067 6663 5101 6697
rect 5135 6663 5169 6697
rect 5203 6663 5237 6697
rect 5271 6663 5305 6697
rect 5339 6663 5373 6697
rect 5407 6663 5441 6697
rect 5475 6663 5509 6697
rect 5543 6663 5577 6697
rect 5611 6663 5645 6697
rect 5679 6663 5713 6697
rect 5747 6663 5781 6697
rect 5815 6663 5849 6697
rect 5883 6663 5917 6697
rect 5951 6663 5985 6697
rect 6019 6663 6053 6697
rect 6087 6663 6121 6697
rect 6155 6663 6189 6697
rect 6223 6663 6257 6697
rect 6291 6663 6325 6697
rect 6359 6663 6393 6697
rect 6427 6663 6461 6697
rect 6495 6663 6529 6697
rect 6563 6663 6597 6697
rect 6631 6663 6665 6697
rect 6699 6663 6733 6697
rect 6767 6663 6801 6697
rect 6835 6663 6869 6697
rect 6903 6663 6937 6697
rect 6971 6663 7005 6697
rect 7039 6663 7073 6697
rect 7107 6663 7141 6697
rect 7175 6663 7209 6697
rect 7243 6663 7277 6697
rect 7311 6663 7345 6697
rect 7379 6663 7413 6697
rect 7447 6663 7481 6697
rect 7515 6663 7549 6697
rect 7583 6663 7617 6697
rect 7651 6663 7685 6697
rect 7719 6663 7753 6697
rect 7787 6663 7821 6697
rect 7855 6663 7889 6697
rect 7923 6663 7957 6697
rect 7991 6663 8025 6697
rect 8059 6663 8093 6697
rect 8127 6663 8161 6697
rect 8195 6663 8229 6697
rect 8263 6663 8400 6697
rect 0 6640 8400 6663
rect 0 5440 80 6640
rect 8320 5440 8400 6640
rect 0 5417 8400 5440
rect 0 5383 137 5417
rect 171 5383 205 5417
rect 239 5383 273 5417
rect 307 5383 341 5417
rect 375 5383 409 5417
rect 443 5383 477 5417
rect 511 5383 545 5417
rect 579 5383 613 5417
rect 647 5383 681 5417
rect 715 5383 749 5417
rect 783 5383 817 5417
rect 851 5383 885 5417
rect 919 5383 953 5417
rect 987 5383 1021 5417
rect 1055 5383 1089 5417
rect 1123 5383 1157 5417
rect 1191 5383 1225 5417
rect 1259 5383 1293 5417
rect 1327 5383 1361 5417
rect 1395 5383 1429 5417
rect 1463 5383 1497 5417
rect 1531 5383 1565 5417
rect 1599 5383 1633 5417
rect 1667 5383 1701 5417
rect 1735 5383 1769 5417
rect 1803 5383 1837 5417
rect 1871 5383 1905 5417
rect 1939 5383 1973 5417
rect 2007 5383 2041 5417
rect 2075 5383 2109 5417
rect 2143 5383 2177 5417
rect 2211 5383 2245 5417
rect 2279 5383 2313 5417
rect 2347 5383 2381 5417
rect 2415 5383 2449 5417
rect 2483 5383 2517 5417
rect 2551 5383 2585 5417
rect 2619 5383 2653 5417
rect 2687 5383 2721 5417
rect 2755 5383 2789 5417
rect 2823 5383 2857 5417
rect 2891 5383 2925 5417
rect 2959 5383 2993 5417
rect 3027 5383 3061 5417
rect 3095 5383 3129 5417
rect 3163 5383 3197 5417
rect 3231 5383 3265 5417
rect 3299 5383 3333 5417
rect 3367 5383 3401 5417
rect 3435 5383 3469 5417
rect 3503 5383 3537 5417
rect 3571 5383 3605 5417
rect 3639 5383 3673 5417
rect 3707 5383 3741 5417
rect 3775 5383 3809 5417
rect 3843 5383 3877 5417
rect 3911 5383 3945 5417
rect 3979 5383 4013 5417
rect 4047 5383 4081 5417
rect 4115 5383 4149 5417
rect 4183 5383 4217 5417
rect 4251 5383 4285 5417
rect 4319 5383 4353 5417
rect 4387 5383 4421 5417
rect 4455 5383 4489 5417
rect 4523 5383 4557 5417
rect 4591 5383 4625 5417
rect 4659 5383 4693 5417
rect 4727 5383 4761 5417
rect 4795 5383 4829 5417
rect 4863 5383 4897 5417
rect 4931 5383 4965 5417
rect 4999 5383 5033 5417
rect 5067 5383 5101 5417
rect 5135 5383 5169 5417
rect 5203 5383 5237 5417
rect 5271 5383 5305 5417
rect 5339 5383 5373 5417
rect 5407 5383 5441 5417
rect 5475 5383 5509 5417
rect 5543 5383 5577 5417
rect 5611 5383 5645 5417
rect 5679 5383 5713 5417
rect 5747 5383 5781 5417
rect 5815 5383 5849 5417
rect 5883 5383 5917 5417
rect 5951 5383 5985 5417
rect 6019 5383 6053 5417
rect 6087 5383 6121 5417
rect 6155 5383 6189 5417
rect 6223 5383 6257 5417
rect 6291 5383 6325 5417
rect 6359 5383 6393 5417
rect 6427 5383 6461 5417
rect 6495 5383 6529 5417
rect 6563 5383 6597 5417
rect 6631 5383 6665 5417
rect 6699 5383 6733 5417
rect 6767 5383 6801 5417
rect 6835 5383 6869 5417
rect 6903 5383 6937 5417
rect 6971 5383 7005 5417
rect 7039 5383 7073 5417
rect 7107 5383 7141 5417
rect 7175 5383 7209 5417
rect 7243 5383 7277 5417
rect 7311 5383 7345 5417
rect 7379 5383 7413 5417
rect 7447 5383 7481 5417
rect 7515 5383 7549 5417
rect 7583 5383 7617 5417
rect 7651 5383 7685 5417
rect 7719 5383 7753 5417
rect 7787 5383 7821 5417
rect 7855 5383 7889 5417
rect 7923 5383 7957 5417
rect 7991 5383 8025 5417
rect 8059 5383 8093 5417
rect 8127 5383 8161 5417
rect 8195 5383 8229 5417
rect 8263 5383 8400 5417
rect 0 5360 8400 5383
rect 0 5287 80 5360
rect 0 5253 23 5287
rect 57 5253 80 5287
rect 8320 5287 8400 5360
rect 0 5219 80 5253
rect 0 5185 23 5219
rect 57 5185 80 5219
rect 0 5151 80 5185
rect 0 5117 23 5151
rect 57 5117 80 5151
rect 0 5083 80 5117
rect 0 5049 23 5083
rect 57 5049 80 5083
rect 0 5015 80 5049
rect 0 4981 23 5015
rect 57 4981 80 5015
rect 0 4947 80 4981
rect 0 4913 23 4947
rect 57 4913 80 4947
rect 0 4879 80 4913
rect 0 4845 23 4879
rect 57 4845 80 4879
rect 0 4811 80 4845
rect 0 4777 23 4811
rect 57 4777 80 4811
rect 0 4743 80 4777
rect 0 4709 23 4743
rect 57 4709 80 4743
rect 0 4675 80 4709
rect 0 4641 23 4675
rect 57 4641 80 4675
rect 0 4607 80 4641
rect 0 4573 23 4607
rect 57 4573 80 4607
rect 0 4539 80 4573
rect 0 4505 23 4539
rect 57 4505 80 4539
rect 0 4471 80 4505
rect 0 4437 23 4471
rect 57 4437 80 4471
rect 0 4403 80 4437
rect 0 4369 23 4403
rect 57 4369 80 4403
rect 0 4335 80 4369
rect 0 4301 23 4335
rect 57 4301 80 4335
rect 0 4267 80 4301
rect 0 4233 23 4267
rect 57 4233 80 4267
rect 8320 5253 8343 5287
rect 8377 5253 8400 5287
rect 8320 5219 8400 5253
rect 8320 5185 8343 5219
rect 8377 5185 8400 5219
rect 8320 5151 8400 5185
rect 8320 5117 8343 5151
rect 8377 5117 8400 5151
rect 8320 5083 8400 5117
rect 8320 5049 8343 5083
rect 8377 5049 8400 5083
rect 8320 5015 8400 5049
rect 8320 4981 8343 5015
rect 8377 4981 8400 5015
rect 8320 4947 8400 4981
rect 8320 4913 8343 4947
rect 8377 4913 8400 4947
rect 8320 4879 8400 4913
rect 8320 4845 8343 4879
rect 8377 4845 8400 4879
rect 8320 4811 8400 4845
rect 8320 4777 8343 4811
rect 8377 4777 8400 4811
rect 8320 4743 8400 4777
rect 8320 4709 8343 4743
rect 8377 4709 8400 4743
rect 8320 4675 8400 4709
rect 8320 4641 8343 4675
rect 8377 4641 8400 4675
rect 8320 4607 8400 4641
rect 8320 4573 8343 4607
rect 8377 4573 8400 4607
rect 8320 4539 8400 4573
rect 8320 4505 8343 4539
rect 8377 4505 8400 4539
rect 8320 4471 8400 4505
rect 8320 4437 8343 4471
rect 8377 4437 8400 4471
rect 8320 4403 8400 4437
rect 8320 4369 8343 4403
rect 8377 4369 8400 4403
rect 8320 4335 8400 4369
rect 8320 4301 8343 4335
rect 8377 4301 8400 4335
rect 8320 4267 8400 4301
rect 0 4160 80 4233
rect 8320 4233 8343 4267
rect 8377 4233 8400 4267
rect 8320 4160 8400 4233
rect 0 4137 8400 4160
rect 0 4103 137 4137
rect 171 4103 205 4137
rect 239 4103 273 4137
rect 307 4103 341 4137
rect 375 4103 409 4137
rect 443 4103 477 4137
rect 511 4103 545 4137
rect 579 4103 613 4137
rect 647 4103 681 4137
rect 715 4103 749 4137
rect 783 4103 817 4137
rect 851 4103 885 4137
rect 919 4103 953 4137
rect 987 4103 1021 4137
rect 1055 4103 1089 4137
rect 1123 4103 1157 4137
rect 1191 4103 1225 4137
rect 1259 4103 1293 4137
rect 1327 4103 1361 4137
rect 1395 4103 1429 4137
rect 1463 4103 1497 4137
rect 1531 4103 1565 4137
rect 1599 4103 1633 4137
rect 1667 4103 1701 4137
rect 1735 4103 1769 4137
rect 1803 4103 1837 4137
rect 1871 4103 1905 4137
rect 1939 4103 1973 4137
rect 2007 4103 2041 4137
rect 2075 4103 2109 4137
rect 2143 4103 2177 4137
rect 2211 4103 2245 4137
rect 2279 4103 2313 4137
rect 2347 4103 2381 4137
rect 2415 4103 2449 4137
rect 2483 4103 2517 4137
rect 2551 4103 2585 4137
rect 2619 4103 2653 4137
rect 2687 4103 2721 4137
rect 2755 4103 2789 4137
rect 2823 4103 2857 4137
rect 2891 4103 2925 4137
rect 2959 4103 2993 4137
rect 3027 4103 3061 4137
rect 3095 4103 3129 4137
rect 3163 4103 3197 4137
rect 3231 4103 3265 4137
rect 3299 4103 3333 4137
rect 3367 4103 3401 4137
rect 3435 4103 3469 4137
rect 3503 4103 3537 4137
rect 3571 4103 3605 4137
rect 3639 4103 3673 4137
rect 3707 4103 3741 4137
rect 3775 4103 3809 4137
rect 3843 4103 3877 4137
rect 3911 4103 3945 4137
rect 3979 4103 4013 4137
rect 4047 4103 4081 4137
rect 4115 4103 4149 4137
rect 4183 4103 4217 4137
rect 4251 4103 4285 4137
rect 4319 4103 4353 4137
rect 4387 4103 4421 4137
rect 4455 4103 4489 4137
rect 4523 4103 4557 4137
rect 4591 4103 4625 4137
rect 4659 4103 4693 4137
rect 4727 4103 4761 4137
rect 4795 4103 4829 4137
rect 4863 4103 4897 4137
rect 4931 4103 4965 4137
rect 4999 4103 5033 4137
rect 5067 4103 5101 4137
rect 5135 4103 5169 4137
rect 5203 4103 5237 4137
rect 5271 4103 5305 4137
rect 5339 4103 5373 4137
rect 5407 4103 5441 4137
rect 5475 4103 5509 4137
rect 5543 4103 5577 4137
rect 5611 4103 5645 4137
rect 5679 4103 5713 4137
rect 5747 4103 5781 4137
rect 5815 4103 5849 4137
rect 5883 4103 5917 4137
rect 5951 4103 5985 4137
rect 6019 4103 6053 4137
rect 6087 4103 6121 4137
rect 6155 4103 6189 4137
rect 6223 4103 6257 4137
rect 6291 4103 6325 4137
rect 6359 4103 6393 4137
rect 6427 4103 6461 4137
rect 6495 4103 6529 4137
rect 6563 4103 6597 4137
rect 6631 4103 6665 4137
rect 6699 4103 6733 4137
rect 6767 4103 6801 4137
rect 6835 4103 6869 4137
rect 6903 4103 6937 4137
rect 6971 4103 7005 4137
rect 7039 4103 7073 4137
rect 7107 4103 7141 4137
rect 7175 4103 7209 4137
rect 7243 4103 7277 4137
rect 7311 4103 7345 4137
rect 7379 4103 7413 4137
rect 7447 4103 7481 4137
rect 7515 4103 7549 4137
rect 7583 4103 7617 4137
rect 7651 4103 7685 4137
rect 7719 4103 7753 4137
rect 7787 4103 7821 4137
rect 7855 4103 7889 4137
rect 7923 4103 7957 4137
rect 7991 4103 8025 4137
rect 8059 4103 8093 4137
rect 8127 4103 8161 4137
rect 8195 4103 8229 4137
rect 8263 4103 8400 4137
rect 0 4080 8400 4103
rect 0 3977 8400 4000
rect 0 3943 137 3977
rect 171 3943 205 3977
rect 239 3943 273 3977
rect 307 3943 341 3977
rect 375 3943 409 3977
rect 443 3943 477 3977
rect 511 3943 545 3977
rect 579 3943 613 3977
rect 647 3943 681 3977
rect 715 3943 749 3977
rect 783 3943 817 3977
rect 851 3943 885 3977
rect 919 3943 953 3977
rect 987 3943 1021 3977
rect 1055 3943 1089 3977
rect 1123 3943 1157 3977
rect 1191 3943 1225 3977
rect 1259 3943 1293 3977
rect 1327 3943 1361 3977
rect 1395 3943 1429 3977
rect 1463 3943 1497 3977
rect 1531 3943 1565 3977
rect 1599 3943 1633 3977
rect 1667 3943 1701 3977
rect 1735 3943 1769 3977
rect 1803 3943 1837 3977
rect 1871 3943 1905 3977
rect 1939 3943 1973 3977
rect 2007 3943 2041 3977
rect 2075 3943 2109 3977
rect 2143 3943 2177 3977
rect 2211 3943 2245 3977
rect 2279 3943 2313 3977
rect 2347 3943 2381 3977
rect 2415 3943 2449 3977
rect 2483 3943 2517 3977
rect 2551 3943 2585 3977
rect 2619 3943 2653 3977
rect 2687 3943 2721 3977
rect 2755 3943 2789 3977
rect 2823 3943 2857 3977
rect 2891 3943 2925 3977
rect 2959 3943 2993 3977
rect 3027 3943 3061 3977
rect 3095 3943 3129 3977
rect 3163 3943 3197 3977
rect 3231 3943 3265 3977
rect 3299 3943 3333 3977
rect 3367 3943 3401 3977
rect 3435 3943 3469 3977
rect 3503 3943 3537 3977
rect 3571 3943 3605 3977
rect 3639 3943 3673 3977
rect 3707 3943 3741 3977
rect 3775 3943 3809 3977
rect 3843 3943 3877 3977
rect 3911 3943 3945 3977
rect 3979 3943 4013 3977
rect 4047 3943 4081 3977
rect 4115 3943 4149 3977
rect 4183 3943 4217 3977
rect 4251 3943 4285 3977
rect 4319 3943 4353 3977
rect 4387 3943 4421 3977
rect 4455 3943 4489 3977
rect 4523 3943 4557 3977
rect 4591 3943 4625 3977
rect 4659 3943 4693 3977
rect 4727 3943 4761 3977
rect 4795 3943 4829 3977
rect 4863 3943 4897 3977
rect 4931 3943 4965 3977
rect 4999 3943 5033 3977
rect 5067 3943 5101 3977
rect 5135 3943 5169 3977
rect 5203 3943 5237 3977
rect 5271 3943 5305 3977
rect 5339 3943 5373 3977
rect 5407 3943 5441 3977
rect 5475 3943 5509 3977
rect 5543 3943 5577 3977
rect 5611 3943 5645 3977
rect 5679 3943 5713 3977
rect 5747 3943 5781 3977
rect 5815 3943 5849 3977
rect 5883 3943 5917 3977
rect 5951 3943 5985 3977
rect 6019 3943 6053 3977
rect 6087 3943 6121 3977
rect 6155 3943 6189 3977
rect 6223 3943 6257 3977
rect 6291 3943 6325 3977
rect 6359 3943 6393 3977
rect 6427 3943 6461 3977
rect 6495 3943 6529 3977
rect 6563 3943 6597 3977
rect 6631 3943 6665 3977
rect 6699 3943 6733 3977
rect 6767 3943 6801 3977
rect 6835 3943 6869 3977
rect 6903 3943 6937 3977
rect 6971 3943 7005 3977
rect 7039 3943 7073 3977
rect 7107 3943 7141 3977
rect 7175 3943 7209 3977
rect 7243 3943 7277 3977
rect 7311 3943 7345 3977
rect 7379 3943 7413 3977
rect 7447 3943 7481 3977
rect 7515 3943 7549 3977
rect 7583 3943 7617 3977
rect 7651 3943 7685 3977
rect 7719 3943 7753 3977
rect 7787 3943 7821 3977
rect 7855 3943 7889 3977
rect 7923 3943 7957 3977
rect 7991 3943 8025 3977
rect 8059 3943 8093 3977
rect 8127 3943 8161 3977
rect 8195 3943 8229 3977
rect 8263 3943 8400 3977
rect 0 3920 8400 3943
rect 0 3847 80 3920
rect 0 3813 23 3847
rect 57 3813 80 3847
rect 8320 3847 8400 3920
rect 0 3779 80 3813
rect 0 3745 23 3779
rect 57 3745 80 3779
rect 0 3711 80 3745
rect 0 3677 23 3711
rect 57 3677 80 3711
rect 0 3643 80 3677
rect 0 3609 23 3643
rect 57 3609 80 3643
rect 0 3575 80 3609
rect 0 3541 23 3575
rect 57 3541 80 3575
rect 0 3507 80 3541
rect 0 3473 23 3507
rect 57 3473 80 3507
rect 0 3439 80 3473
rect 0 3405 23 3439
rect 57 3405 80 3439
rect 0 3371 80 3405
rect 0 3337 23 3371
rect 57 3337 80 3371
rect 0 3303 80 3337
rect 0 3269 23 3303
rect 57 3269 80 3303
rect 0 3235 80 3269
rect 0 3201 23 3235
rect 57 3201 80 3235
rect 0 3167 80 3201
rect 0 3133 23 3167
rect 57 3133 80 3167
rect 0 3099 80 3133
rect 0 3065 23 3099
rect 57 3065 80 3099
rect 0 3031 80 3065
rect 0 2997 23 3031
rect 57 2997 80 3031
rect 0 2963 80 2997
rect 0 2929 23 2963
rect 57 2929 80 2963
rect 0 2895 80 2929
rect 0 2861 23 2895
rect 57 2861 80 2895
rect 0 2827 80 2861
rect 0 2793 23 2827
rect 57 2793 80 2827
rect 8320 3813 8343 3847
rect 8377 3813 8400 3847
rect 8320 3779 8400 3813
rect 8320 3745 8343 3779
rect 8377 3745 8400 3779
rect 8320 3711 8400 3745
rect 8320 3677 8343 3711
rect 8377 3677 8400 3711
rect 8320 3643 8400 3677
rect 8320 3609 8343 3643
rect 8377 3609 8400 3643
rect 8320 3575 8400 3609
rect 8320 3541 8343 3575
rect 8377 3541 8400 3575
rect 8320 3507 8400 3541
rect 8320 3473 8343 3507
rect 8377 3473 8400 3507
rect 8320 3439 8400 3473
rect 8320 3405 8343 3439
rect 8377 3405 8400 3439
rect 8320 3371 8400 3405
rect 8320 3337 8343 3371
rect 8377 3337 8400 3371
rect 8320 3303 8400 3337
rect 8320 3269 8343 3303
rect 8377 3269 8400 3303
rect 8320 3235 8400 3269
rect 8320 3201 8343 3235
rect 8377 3201 8400 3235
rect 8320 3167 8400 3201
rect 8320 3133 8343 3167
rect 8377 3133 8400 3167
rect 8320 3099 8400 3133
rect 8320 3065 8343 3099
rect 8377 3065 8400 3099
rect 8320 3031 8400 3065
rect 8320 2997 8343 3031
rect 8377 2997 8400 3031
rect 8320 2963 8400 2997
rect 8320 2929 8343 2963
rect 8377 2929 8400 2963
rect 8320 2895 8400 2929
rect 8320 2861 8343 2895
rect 8377 2861 8400 2895
rect 8320 2827 8400 2861
rect 0 2720 80 2793
rect 8320 2793 8343 2827
rect 8377 2793 8400 2827
rect 8320 2720 8400 2793
rect 0 2697 8400 2720
rect 0 2663 151 2697
rect 185 2663 219 2697
rect 253 2663 287 2697
rect 321 2663 355 2697
rect 389 2663 423 2697
rect 457 2663 491 2697
rect 525 2663 559 2697
rect 593 2663 627 2697
rect 661 2663 695 2697
rect 729 2663 763 2697
rect 797 2663 831 2697
rect 865 2663 899 2697
rect 933 2663 967 2697
rect 1001 2663 1035 2697
rect 1069 2663 1103 2697
rect 1137 2663 1171 2697
rect 1205 2663 1239 2697
rect 1273 2663 1307 2697
rect 1341 2663 1375 2697
rect 1409 2663 1443 2697
rect 1477 2663 1511 2697
rect 1545 2663 1579 2697
rect 1613 2663 1647 2697
rect 1681 2663 1715 2697
rect 1749 2663 1783 2697
rect 1817 2663 1851 2697
rect 1885 2663 1919 2697
rect 1953 2663 1987 2697
rect 2021 2663 2055 2697
rect 2089 2663 2123 2697
rect 2157 2663 2191 2697
rect 2225 2663 2259 2697
rect 2293 2663 2327 2697
rect 2361 2663 2395 2697
rect 2429 2663 2463 2697
rect 2497 2663 2531 2697
rect 2565 2663 2599 2697
rect 2633 2663 2667 2697
rect 2701 2663 2735 2697
rect 2769 2663 2803 2697
rect 2837 2663 2871 2697
rect 2905 2663 2939 2697
rect 2973 2663 3007 2697
rect 3041 2663 3075 2697
rect 3109 2663 3143 2697
rect 3177 2663 3211 2697
rect 3245 2663 3279 2697
rect 3313 2663 3347 2697
rect 3381 2663 3415 2697
rect 3449 2663 3483 2697
rect 3517 2663 3551 2697
rect 3585 2663 3619 2697
rect 3653 2663 3687 2697
rect 3721 2663 3755 2697
rect 3789 2663 3823 2697
rect 3857 2663 3891 2697
rect 3925 2663 3959 2697
rect 3993 2663 4027 2697
rect 4061 2663 4095 2697
rect 4129 2663 4163 2697
rect 4197 2663 4231 2697
rect 4265 2663 4299 2697
rect 4333 2663 4367 2697
rect 4401 2663 4435 2697
rect 4469 2663 4503 2697
rect 4537 2663 4571 2697
rect 4605 2663 4639 2697
rect 4673 2663 4707 2697
rect 4741 2663 4775 2697
rect 4809 2663 4843 2697
rect 4877 2663 4911 2697
rect 4945 2663 4979 2697
rect 5013 2663 5047 2697
rect 5081 2663 5115 2697
rect 5149 2663 5183 2697
rect 5217 2663 5251 2697
rect 5285 2663 5319 2697
rect 5353 2663 5387 2697
rect 5421 2663 5455 2697
rect 5489 2663 5523 2697
rect 5557 2663 5591 2697
rect 5625 2663 5659 2697
rect 5693 2663 5727 2697
rect 5761 2663 5795 2697
rect 5829 2663 5863 2697
rect 5897 2663 5931 2697
rect 5965 2663 5999 2697
rect 6033 2663 6067 2697
rect 6101 2663 6135 2697
rect 6169 2663 6203 2697
rect 6237 2663 6271 2697
rect 6305 2663 6339 2697
rect 6373 2663 6407 2697
rect 6441 2663 6475 2697
rect 6509 2663 6543 2697
rect 6577 2663 6611 2697
rect 6645 2663 6679 2697
rect 6713 2663 6747 2697
rect 6781 2663 6815 2697
rect 6849 2663 6883 2697
rect 6917 2663 6951 2697
rect 6985 2663 7019 2697
rect 7053 2663 7087 2697
rect 7121 2663 7155 2697
rect 7189 2663 7223 2697
rect 7257 2663 7291 2697
rect 7325 2663 7359 2697
rect 7393 2663 7427 2697
rect 7461 2663 7495 2697
rect 7529 2663 7563 2697
rect 7597 2663 7631 2697
rect 7665 2663 7699 2697
rect 7733 2663 7767 2697
rect 7801 2663 7835 2697
rect 7869 2663 7903 2697
rect 7937 2663 7971 2697
rect 8005 2663 8039 2697
rect 8073 2663 8107 2697
rect 8141 2663 8175 2697
rect 8209 2663 8400 2697
rect 0 2640 8400 2663
rect 0 2537 8400 2560
rect 0 2503 151 2537
rect 185 2503 219 2537
rect 253 2503 287 2537
rect 321 2503 355 2537
rect 389 2503 423 2537
rect 457 2503 491 2537
rect 525 2503 559 2537
rect 593 2503 627 2537
rect 661 2503 695 2537
rect 729 2503 763 2537
rect 797 2503 831 2537
rect 865 2503 899 2537
rect 933 2503 967 2537
rect 1001 2503 1035 2537
rect 1069 2503 1103 2537
rect 1137 2503 1171 2537
rect 1205 2503 1239 2537
rect 1273 2503 1307 2537
rect 1341 2503 1375 2537
rect 1409 2503 1443 2537
rect 1477 2503 1511 2537
rect 1545 2503 1579 2537
rect 1613 2503 1647 2537
rect 1681 2503 1715 2537
rect 1749 2503 1783 2537
rect 1817 2503 1851 2537
rect 1885 2503 1919 2537
rect 1953 2503 1987 2537
rect 2021 2503 2055 2537
rect 2089 2503 2123 2537
rect 2157 2503 2191 2537
rect 2225 2503 2259 2537
rect 2293 2503 2327 2537
rect 2361 2503 2395 2537
rect 2429 2503 2463 2537
rect 2497 2503 2531 2537
rect 2565 2503 2599 2537
rect 2633 2503 2667 2537
rect 2701 2503 2735 2537
rect 2769 2503 2803 2537
rect 2837 2503 2871 2537
rect 2905 2503 2939 2537
rect 2973 2503 3007 2537
rect 3041 2503 3075 2537
rect 3109 2503 3143 2537
rect 3177 2503 3211 2537
rect 3245 2503 3279 2537
rect 3313 2503 3347 2537
rect 3381 2503 3415 2537
rect 3449 2503 3483 2537
rect 3517 2503 3551 2537
rect 3585 2503 3619 2537
rect 3653 2503 3687 2537
rect 3721 2503 3755 2537
rect 3789 2503 3823 2537
rect 3857 2503 3891 2537
rect 3925 2503 3959 2537
rect 3993 2503 4027 2537
rect 4061 2503 4095 2537
rect 4129 2503 4163 2537
rect 4197 2503 4231 2537
rect 4265 2503 4299 2537
rect 4333 2503 4367 2537
rect 4401 2503 4435 2537
rect 4469 2503 4503 2537
rect 4537 2503 4571 2537
rect 4605 2503 4639 2537
rect 4673 2503 4707 2537
rect 4741 2503 4775 2537
rect 4809 2503 4843 2537
rect 4877 2503 4911 2537
rect 4945 2503 4979 2537
rect 5013 2503 5047 2537
rect 5081 2503 5115 2537
rect 5149 2503 5183 2537
rect 5217 2503 5251 2537
rect 5285 2503 5319 2537
rect 5353 2503 5387 2537
rect 5421 2503 5455 2537
rect 5489 2503 5523 2537
rect 5557 2503 5591 2537
rect 5625 2503 5659 2537
rect 5693 2503 5727 2537
rect 5761 2503 5795 2537
rect 5829 2503 5863 2537
rect 5897 2503 5931 2537
rect 5965 2503 5999 2537
rect 6033 2503 6067 2537
rect 6101 2503 6135 2537
rect 6169 2503 6203 2537
rect 6237 2503 6271 2537
rect 6305 2503 6339 2537
rect 6373 2503 6407 2537
rect 6441 2503 6475 2537
rect 6509 2503 6543 2537
rect 6577 2503 6611 2537
rect 6645 2503 6679 2537
rect 6713 2503 6747 2537
rect 6781 2503 6815 2537
rect 6849 2503 6883 2537
rect 6917 2503 6951 2537
rect 6985 2503 7019 2537
rect 7053 2503 7087 2537
rect 7121 2503 7155 2537
rect 7189 2503 7223 2537
rect 7257 2503 7291 2537
rect 7325 2503 7359 2537
rect 7393 2503 7427 2537
rect 7461 2503 7495 2537
rect 7529 2503 7563 2537
rect 7597 2503 7631 2537
rect 7665 2503 7699 2537
rect 7733 2503 7767 2537
rect 7801 2503 7835 2537
rect 7869 2503 7903 2537
rect 7937 2503 7971 2537
rect 8005 2503 8039 2537
rect 8073 2503 8107 2537
rect 8141 2503 8175 2537
rect 8209 2503 8400 2537
rect 0 2480 8400 2503
rect 0 2407 80 2480
rect 0 2373 23 2407
rect 57 2373 80 2407
rect 8320 2419 8400 2480
rect 0 2339 80 2373
rect 0 2305 23 2339
rect 57 2305 80 2339
rect 0 2271 80 2305
rect 0 2237 23 2271
rect 57 2237 80 2271
rect 0 2203 80 2237
rect 0 2169 23 2203
rect 57 2169 80 2203
rect 0 2135 80 2169
rect 0 2101 23 2135
rect 57 2101 80 2135
rect 0 2067 80 2101
rect 0 2033 23 2067
rect 57 2033 80 2067
rect 0 1999 80 2033
rect 0 1965 23 1999
rect 57 1965 80 1999
rect 0 1931 80 1965
rect 0 1897 23 1931
rect 57 1897 80 1931
rect 0 1863 80 1897
rect 0 1829 23 1863
rect 57 1829 80 1863
rect 0 1795 80 1829
rect 0 1761 23 1795
rect 57 1761 80 1795
rect 0 1727 80 1761
rect 0 1693 23 1727
rect 57 1693 80 1727
rect 0 1659 80 1693
rect 0 1625 23 1659
rect 57 1625 80 1659
rect 0 1591 80 1625
rect 0 1557 23 1591
rect 57 1557 80 1591
rect 0 1523 80 1557
rect 0 1489 23 1523
rect 57 1489 80 1523
rect 0 1455 80 1489
rect 0 1421 23 1455
rect 57 1421 80 1455
rect 0 1387 80 1421
rect 0 1353 23 1387
rect 57 1353 80 1387
rect 8320 2385 8343 2419
rect 8377 2385 8400 2419
rect 8320 2351 8400 2385
rect 8320 2317 8343 2351
rect 8377 2317 8400 2351
rect 8320 2283 8400 2317
rect 8320 2249 8343 2283
rect 8377 2249 8400 2283
rect 8320 2215 8400 2249
rect 8320 2181 8343 2215
rect 8377 2181 8400 2215
rect 8320 2147 8400 2181
rect 8320 2113 8343 2147
rect 8377 2113 8400 2147
rect 8320 2079 8400 2113
rect 8320 2045 8343 2079
rect 8377 2045 8400 2079
rect 8320 2011 8400 2045
rect 8320 1977 8343 2011
rect 8377 1977 8400 2011
rect 8320 1943 8400 1977
rect 8320 1909 8343 1943
rect 8377 1909 8400 1943
rect 8320 1875 8400 1909
rect 8320 1841 8343 1875
rect 8377 1841 8400 1875
rect 8320 1807 8400 1841
rect 8320 1773 8343 1807
rect 8377 1773 8400 1807
rect 8320 1739 8400 1773
rect 8320 1705 8343 1739
rect 8377 1705 8400 1739
rect 8320 1671 8400 1705
rect 8320 1637 8343 1671
rect 8377 1637 8400 1671
rect 8320 1603 8400 1637
rect 8320 1569 8343 1603
rect 8377 1569 8400 1603
rect 8320 1535 8400 1569
rect 8320 1501 8343 1535
rect 8377 1501 8400 1535
rect 8320 1467 8400 1501
rect 8320 1433 8343 1467
rect 8377 1433 8400 1467
rect 8320 1399 8400 1433
rect 8320 1365 8343 1399
rect 8377 1365 8400 1399
rect 0 1280 80 1353
rect 8320 1331 8400 1365
rect 8320 1297 8343 1331
rect 8377 1297 8400 1331
rect 8320 1280 8400 1297
rect 0 1263 8400 1280
rect 0 1257 8343 1263
rect 0 1223 137 1257
rect 171 1223 205 1257
rect 239 1223 273 1257
rect 307 1223 341 1257
rect 375 1223 409 1257
rect 443 1223 477 1257
rect 511 1223 545 1257
rect 579 1223 613 1257
rect 647 1223 681 1257
rect 715 1223 749 1257
rect 783 1223 817 1257
rect 851 1223 885 1257
rect 919 1223 953 1257
rect 987 1223 1021 1257
rect 1055 1223 1089 1257
rect 1123 1223 1157 1257
rect 1191 1223 1225 1257
rect 1259 1223 1293 1257
rect 1327 1223 1361 1257
rect 1395 1223 1429 1257
rect 1463 1223 1497 1257
rect 1531 1223 1565 1257
rect 1599 1223 1633 1257
rect 1667 1223 1701 1257
rect 1735 1223 1769 1257
rect 1803 1223 1837 1257
rect 1871 1223 1905 1257
rect 1939 1223 1973 1257
rect 2007 1223 2041 1257
rect 2075 1223 2109 1257
rect 2143 1223 2177 1257
rect 2211 1223 2245 1257
rect 2279 1223 2313 1257
rect 2347 1223 2381 1257
rect 2415 1223 2449 1257
rect 2483 1223 2517 1257
rect 2551 1223 2585 1257
rect 2619 1223 2653 1257
rect 2687 1223 2721 1257
rect 2755 1223 2789 1257
rect 2823 1223 2857 1257
rect 2891 1223 2925 1257
rect 2959 1223 2993 1257
rect 3027 1223 3061 1257
rect 3095 1223 3129 1257
rect 3163 1223 3197 1257
rect 3231 1223 3265 1257
rect 3299 1223 3333 1257
rect 3367 1223 3401 1257
rect 3435 1223 3469 1257
rect 3503 1223 3537 1257
rect 3571 1223 3605 1257
rect 3639 1223 3673 1257
rect 3707 1223 3741 1257
rect 3775 1223 3809 1257
rect 3843 1223 3877 1257
rect 3911 1223 3945 1257
rect 3979 1223 4013 1257
rect 4047 1223 4081 1257
rect 4115 1223 4149 1257
rect 4183 1223 4217 1257
rect 4251 1223 4285 1257
rect 4319 1223 4353 1257
rect 4387 1223 4421 1257
rect 4455 1223 4489 1257
rect 4523 1223 4557 1257
rect 4591 1223 4625 1257
rect 4659 1223 4693 1257
rect 4727 1223 4761 1257
rect 4795 1223 4829 1257
rect 4863 1223 4897 1257
rect 4931 1223 4965 1257
rect 4999 1223 5033 1257
rect 5067 1223 5101 1257
rect 5135 1223 5169 1257
rect 5203 1223 5237 1257
rect 5271 1223 5305 1257
rect 5339 1223 5373 1257
rect 5407 1223 5441 1257
rect 5475 1223 5509 1257
rect 5543 1223 5577 1257
rect 5611 1223 5645 1257
rect 5679 1223 5713 1257
rect 5747 1223 5781 1257
rect 5815 1223 5849 1257
rect 5883 1223 5917 1257
rect 5951 1223 5985 1257
rect 6019 1223 6053 1257
rect 6087 1223 6121 1257
rect 6155 1223 6189 1257
rect 6223 1223 6257 1257
rect 6291 1223 6325 1257
rect 6359 1223 6393 1257
rect 6427 1223 6461 1257
rect 6495 1223 6529 1257
rect 6563 1223 6597 1257
rect 6631 1223 6665 1257
rect 6699 1223 6733 1257
rect 6767 1223 6801 1257
rect 6835 1223 6869 1257
rect 6903 1223 6937 1257
rect 6971 1223 7005 1257
rect 7039 1223 7073 1257
rect 7107 1223 7141 1257
rect 7175 1223 7209 1257
rect 7243 1223 7277 1257
rect 7311 1223 7345 1257
rect 7379 1223 7413 1257
rect 7447 1223 7481 1257
rect 7515 1223 7549 1257
rect 7583 1223 7617 1257
rect 7651 1223 7685 1257
rect 7719 1223 7753 1257
rect 7787 1223 7821 1257
rect 7855 1223 7889 1257
rect 7923 1223 7957 1257
rect 7991 1223 8025 1257
rect 8059 1223 8093 1257
rect 8127 1223 8161 1257
rect 8195 1223 8229 1257
rect 8263 1229 8343 1257
rect 8377 1229 8400 1263
rect 8263 1223 8400 1229
rect 0 1200 8400 1223
rect 8320 1195 8400 1200
rect 8320 1161 8343 1195
rect 8377 1161 8400 1195
rect 8320 1127 8400 1161
rect 8320 1093 8343 1127
rect 8377 1093 8400 1127
rect 8320 1059 8400 1093
rect 8320 1025 8343 1059
rect 8377 1025 8400 1059
rect 8320 991 8400 1025
rect 8320 957 8343 991
rect 8377 957 8400 991
rect 8320 923 8400 957
rect 8320 889 8343 923
rect 8377 889 8400 923
rect 8320 855 8400 889
rect 8320 821 8343 855
rect 8377 821 8400 855
rect 8320 787 8400 821
rect 8320 753 8343 787
rect 8377 753 8400 787
rect 8320 719 8400 753
rect 8320 685 8343 719
rect 8377 685 8400 719
rect 8320 651 8400 685
rect 8320 640 8343 651
rect 0 617 8343 640
rect 8377 617 8400 651
rect 0 583 137 617
rect 171 583 205 617
rect 239 583 273 617
rect 307 583 341 617
rect 375 583 409 617
rect 443 583 477 617
rect 511 583 545 617
rect 579 583 613 617
rect 647 583 681 617
rect 715 583 749 617
rect 783 583 817 617
rect 851 583 885 617
rect 919 583 953 617
rect 987 583 1021 617
rect 1055 583 1089 617
rect 1123 583 1157 617
rect 1191 583 1225 617
rect 1259 583 1293 617
rect 1327 583 1361 617
rect 1395 583 1429 617
rect 1463 583 1497 617
rect 1531 583 1565 617
rect 1599 583 1633 617
rect 1667 583 1701 617
rect 1735 583 1769 617
rect 1803 583 1837 617
rect 1871 583 1905 617
rect 1939 583 1973 617
rect 2007 583 2041 617
rect 2075 583 2109 617
rect 2143 583 2177 617
rect 2211 583 2245 617
rect 2279 583 2313 617
rect 2347 583 2381 617
rect 2415 583 2449 617
rect 2483 583 2517 617
rect 2551 583 2585 617
rect 2619 583 2653 617
rect 2687 583 2721 617
rect 2755 583 2789 617
rect 2823 583 2857 617
rect 2891 583 2925 617
rect 2959 583 2993 617
rect 3027 583 3061 617
rect 3095 583 3129 617
rect 3163 583 3197 617
rect 3231 583 3265 617
rect 3299 583 3333 617
rect 3367 583 3401 617
rect 3435 583 3469 617
rect 3503 583 3537 617
rect 3571 583 3605 617
rect 3639 583 3673 617
rect 3707 583 3741 617
rect 3775 583 3809 617
rect 3843 583 3877 617
rect 3911 583 3945 617
rect 3979 583 4013 617
rect 4047 583 4081 617
rect 4115 583 4149 617
rect 4183 583 4217 617
rect 4251 583 4285 617
rect 4319 583 4353 617
rect 4387 583 4421 617
rect 4455 583 4489 617
rect 4523 583 4557 617
rect 4591 583 4625 617
rect 4659 583 4693 617
rect 4727 583 4761 617
rect 4795 583 4829 617
rect 4863 583 4897 617
rect 4931 583 4965 617
rect 4999 583 5033 617
rect 5067 583 5101 617
rect 5135 583 5169 617
rect 5203 583 5237 617
rect 5271 583 5305 617
rect 5339 583 5373 617
rect 5407 583 5441 617
rect 5475 583 5509 617
rect 5543 583 5577 617
rect 5611 583 5645 617
rect 5679 583 5713 617
rect 5747 583 5781 617
rect 5815 583 5849 617
rect 5883 583 5917 617
rect 5951 583 5985 617
rect 6019 583 6053 617
rect 6087 583 6121 617
rect 6155 583 6189 617
rect 6223 583 6257 617
rect 6291 583 6325 617
rect 6359 583 6393 617
rect 6427 583 6461 617
rect 6495 583 6529 617
rect 6563 583 6597 617
rect 6631 583 6665 617
rect 6699 583 6733 617
rect 6767 583 6801 617
rect 6835 583 6869 617
rect 6903 583 6937 617
rect 6971 583 7005 617
rect 7039 583 7073 617
rect 7107 583 7141 617
rect 7175 583 7209 617
rect 7243 583 7277 617
rect 7311 583 7345 617
rect 7379 583 7413 617
rect 7447 583 7481 617
rect 7515 583 7549 617
rect 7583 583 7617 617
rect 7651 583 7685 617
rect 7719 583 7753 617
rect 7787 583 7821 617
rect 7855 583 7889 617
rect 7923 583 7957 617
rect 7991 583 8025 617
rect 8059 583 8093 617
rect 8127 583 8161 617
rect 8195 583 8229 617
rect 8263 583 8400 617
rect 0 560 8343 583
rect 0 507 80 560
rect 0 473 23 507
rect 57 473 80 507
rect 8320 549 8343 560
rect 8377 549 8400 583
rect 8320 515 8400 549
rect 8320 481 8343 515
rect 8377 481 8400 515
rect 0 439 80 473
rect 0 405 23 439
rect 57 405 80 439
rect 0 371 80 405
rect 0 337 23 371
rect 57 337 80 371
rect 8320 447 8400 481
rect 8320 413 8343 447
rect 8377 413 8400 447
rect 8320 379 8400 413
rect 0 303 80 337
rect 0 269 23 303
rect 57 269 80 303
rect 0 235 80 269
rect 0 201 23 235
rect 57 201 80 235
rect 0 167 80 201
rect 0 133 23 167
rect 57 133 80 167
rect 8320 345 8343 379
rect 8377 345 8400 379
rect 8320 311 8400 345
rect 8320 277 8343 311
rect 8377 277 8400 311
rect 8320 243 8400 277
rect 8320 209 8343 243
rect 8377 209 8400 243
rect 8320 175 8400 209
rect 0 80 80 133
rect 8320 141 8343 175
rect 8377 141 8400 175
rect 8320 80 8400 141
rect 0 57 8400 80
rect 0 23 137 57
rect 171 23 205 57
rect 239 23 273 57
rect 307 23 341 57
rect 375 23 409 57
rect 443 23 477 57
rect 511 23 545 57
rect 579 23 613 57
rect 647 23 681 57
rect 715 23 749 57
rect 783 23 817 57
rect 851 23 885 57
rect 919 23 953 57
rect 987 23 1021 57
rect 1055 23 1089 57
rect 1123 23 1157 57
rect 1191 23 1225 57
rect 1259 23 1293 57
rect 1327 23 1361 57
rect 1395 23 1429 57
rect 1463 23 1497 57
rect 1531 23 1565 57
rect 1599 23 1633 57
rect 1667 23 1701 57
rect 1735 23 1769 57
rect 1803 23 1837 57
rect 1871 23 1905 57
rect 1939 23 1973 57
rect 2007 23 2041 57
rect 2075 23 2109 57
rect 2143 23 2177 57
rect 2211 23 2245 57
rect 2279 23 2313 57
rect 2347 23 2381 57
rect 2415 23 2449 57
rect 2483 23 2517 57
rect 2551 23 2585 57
rect 2619 23 2653 57
rect 2687 23 2721 57
rect 2755 23 2789 57
rect 2823 23 2857 57
rect 2891 23 2925 57
rect 2959 23 2993 57
rect 3027 23 3061 57
rect 3095 23 3129 57
rect 3163 23 3197 57
rect 3231 23 3265 57
rect 3299 23 3333 57
rect 3367 23 3401 57
rect 3435 23 3469 57
rect 3503 23 3537 57
rect 3571 23 3605 57
rect 3639 23 3673 57
rect 3707 23 3741 57
rect 3775 23 3809 57
rect 3843 23 3877 57
rect 3911 23 3945 57
rect 3979 23 4013 57
rect 4047 23 4081 57
rect 4115 23 4149 57
rect 4183 23 4217 57
rect 4251 23 4285 57
rect 4319 23 4353 57
rect 4387 23 4421 57
rect 4455 23 4489 57
rect 4523 23 4557 57
rect 4591 23 4625 57
rect 4659 23 4693 57
rect 4727 23 4761 57
rect 4795 23 4829 57
rect 4863 23 4897 57
rect 4931 23 4965 57
rect 4999 23 5033 57
rect 5067 23 5101 57
rect 5135 23 5169 57
rect 5203 23 5237 57
rect 5271 23 5305 57
rect 5339 23 5373 57
rect 5407 23 5441 57
rect 5475 23 5509 57
rect 5543 23 5577 57
rect 5611 23 5645 57
rect 5679 23 5713 57
rect 5747 23 5781 57
rect 5815 23 5849 57
rect 5883 23 5917 57
rect 5951 23 5985 57
rect 6019 23 6053 57
rect 6087 23 6121 57
rect 6155 23 6189 57
rect 6223 23 6257 57
rect 6291 23 6325 57
rect 6359 23 6393 57
rect 6427 23 6461 57
rect 6495 23 6529 57
rect 6563 23 6597 57
rect 6631 23 6665 57
rect 6699 23 6733 57
rect 6767 23 6801 57
rect 6835 23 6869 57
rect 6903 23 6937 57
rect 6971 23 7005 57
rect 7039 23 7073 57
rect 7107 23 7141 57
rect 7175 23 7209 57
rect 7243 23 7277 57
rect 7311 23 7345 57
rect 7379 23 7413 57
rect 7447 23 7481 57
rect 7515 23 7549 57
rect 7583 23 7617 57
rect 7651 23 7685 57
rect 7719 23 7753 57
rect 7787 23 7821 57
rect 7855 23 7889 57
rect 7923 23 7957 57
rect 7991 23 8025 57
rect 8059 23 8093 57
rect 8127 23 8161 57
rect 8195 23 8229 57
rect 8263 23 8400 57
rect 0 0 8400 23
rect 0 -423 8400 -400
rect 0 -457 137 -423
rect 171 -457 205 -423
rect 239 -457 273 -423
rect 307 -457 341 -423
rect 375 -457 409 -423
rect 443 -457 477 -423
rect 511 -457 545 -423
rect 579 -457 613 -423
rect 647 -457 681 -423
rect 715 -457 749 -423
rect 783 -457 817 -423
rect 851 -457 885 -423
rect 919 -457 953 -423
rect 987 -457 1021 -423
rect 1055 -457 1089 -423
rect 1123 -457 1157 -423
rect 1191 -457 1225 -423
rect 1259 -457 1293 -423
rect 1327 -457 1361 -423
rect 1395 -457 1429 -423
rect 1463 -457 1497 -423
rect 1531 -457 1565 -423
rect 1599 -457 1633 -423
rect 1667 -457 1701 -423
rect 1735 -457 1769 -423
rect 1803 -457 1837 -423
rect 1871 -457 1905 -423
rect 1939 -457 1973 -423
rect 2007 -457 2041 -423
rect 2075 -457 2109 -423
rect 2143 -457 2177 -423
rect 2211 -457 2245 -423
rect 2279 -457 2313 -423
rect 2347 -457 2381 -423
rect 2415 -457 2449 -423
rect 2483 -457 2517 -423
rect 2551 -457 2585 -423
rect 2619 -457 2653 -423
rect 2687 -457 2721 -423
rect 2755 -457 2789 -423
rect 2823 -457 2857 -423
rect 2891 -457 2925 -423
rect 2959 -457 2993 -423
rect 3027 -457 3061 -423
rect 3095 -457 3129 -423
rect 3163 -457 3197 -423
rect 3231 -457 3265 -423
rect 3299 -457 3333 -423
rect 3367 -457 3401 -423
rect 3435 -457 3469 -423
rect 3503 -457 3537 -423
rect 3571 -457 3605 -423
rect 3639 -457 3673 -423
rect 3707 -457 3741 -423
rect 3775 -457 3809 -423
rect 3843 -457 3877 -423
rect 3911 -457 3945 -423
rect 3979 -457 4013 -423
rect 4047 -457 4081 -423
rect 4115 -457 4149 -423
rect 4183 -457 4217 -423
rect 4251 -457 4285 -423
rect 4319 -457 4353 -423
rect 4387 -457 4421 -423
rect 4455 -457 4489 -423
rect 4523 -457 4557 -423
rect 4591 -457 4625 -423
rect 4659 -457 4693 -423
rect 4727 -457 4761 -423
rect 4795 -457 4829 -423
rect 4863 -457 4897 -423
rect 4931 -457 4965 -423
rect 4999 -457 5033 -423
rect 5067 -457 5101 -423
rect 5135 -457 5169 -423
rect 5203 -457 5237 -423
rect 5271 -457 5305 -423
rect 5339 -457 5373 -423
rect 5407 -457 5441 -423
rect 5475 -457 5509 -423
rect 5543 -457 5577 -423
rect 5611 -457 5645 -423
rect 5679 -457 5713 -423
rect 5747 -457 5781 -423
rect 5815 -457 5849 -423
rect 5883 -457 5917 -423
rect 5951 -457 5985 -423
rect 6019 -457 6053 -423
rect 6087 -457 6121 -423
rect 6155 -457 6189 -423
rect 6223 -457 6257 -423
rect 6291 -457 6325 -423
rect 6359 -457 6393 -423
rect 6427 -457 6461 -423
rect 6495 -457 6529 -423
rect 6563 -457 6597 -423
rect 6631 -457 6665 -423
rect 6699 -457 6733 -423
rect 6767 -457 6801 -423
rect 6835 -457 6869 -423
rect 6903 -457 6937 -423
rect 6971 -457 7005 -423
rect 7039 -457 7073 -423
rect 7107 -457 7141 -423
rect 7175 -457 7209 -423
rect 7243 -457 7277 -423
rect 7311 -457 7345 -423
rect 7379 -457 7413 -423
rect 7447 -457 7481 -423
rect 7515 -457 7549 -423
rect 7583 -457 7617 -423
rect 7651 -457 7685 -423
rect 7719 -457 7753 -423
rect 7787 -457 7821 -423
rect 7855 -457 7889 -423
rect 7923 -457 7957 -423
rect 7991 -457 8025 -423
rect 8059 -457 8093 -423
rect 8127 -457 8161 -423
rect 8195 -457 8229 -423
rect 8263 -457 8400 -423
rect 0 -480 8400 -457
rect 0 -533 80 -480
rect 0 -567 23 -533
rect 57 -567 80 -533
rect 8320 -533 8400 -480
rect 0 -601 80 -567
rect 0 -635 23 -601
rect 57 -635 80 -601
rect 0 -669 80 -635
rect 0 -703 23 -669
rect 57 -703 80 -669
rect 8320 -567 8343 -533
rect 8377 -567 8400 -533
rect 8320 -601 8400 -567
rect 8320 -635 8343 -601
rect 8377 -635 8400 -601
rect 8320 -669 8400 -635
rect 0 -737 80 -703
rect 0 -771 23 -737
rect 57 -771 80 -737
rect 0 -805 80 -771
rect 0 -839 23 -805
rect 57 -839 80 -805
rect 0 -873 80 -839
rect 0 -907 23 -873
rect 57 -907 80 -873
rect 8320 -703 8343 -669
rect 8377 -703 8400 -669
rect 8320 -737 8400 -703
rect 8320 -771 8343 -737
rect 8377 -771 8400 -737
rect 8320 -805 8400 -771
rect 8320 -839 8343 -805
rect 8377 -839 8400 -805
rect 8320 -873 8400 -839
rect 0 -960 80 -907
rect 8320 -907 8343 -873
rect 8377 -907 8400 -873
rect 8320 -960 8400 -907
rect 0 -983 8400 -960
rect 0 -1017 137 -983
rect 171 -1017 205 -983
rect 239 -1017 273 -983
rect 307 -1017 341 -983
rect 375 -1017 409 -983
rect 443 -1017 477 -983
rect 511 -1017 545 -983
rect 579 -1017 613 -983
rect 647 -1017 681 -983
rect 715 -1017 749 -983
rect 783 -1017 817 -983
rect 851 -1017 885 -983
rect 919 -1017 953 -983
rect 987 -1017 1021 -983
rect 1055 -1017 1089 -983
rect 1123 -1017 1157 -983
rect 1191 -1017 1225 -983
rect 1259 -1017 1293 -983
rect 1327 -1017 1361 -983
rect 1395 -1017 1429 -983
rect 1463 -1017 1497 -983
rect 1531 -1017 1565 -983
rect 1599 -1017 1633 -983
rect 1667 -1017 1701 -983
rect 1735 -1017 1769 -983
rect 1803 -1017 1837 -983
rect 1871 -1017 1905 -983
rect 1939 -1017 1973 -983
rect 2007 -1017 2041 -983
rect 2075 -1017 2109 -983
rect 2143 -1017 2177 -983
rect 2211 -1017 2245 -983
rect 2279 -1017 2313 -983
rect 2347 -1017 2381 -983
rect 2415 -1017 2449 -983
rect 2483 -1017 2517 -983
rect 2551 -1017 2585 -983
rect 2619 -1017 2653 -983
rect 2687 -1017 2721 -983
rect 2755 -1017 2789 -983
rect 2823 -1017 2857 -983
rect 2891 -1017 2925 -983
rect 2959 -1017 2993 -983
rect 3027 -1017 3061 -983
rect 3095 -1017 3129 -983
rect 3163 -1017 3197 -983
rect 3231 -1017 3265 -983
rect 3299 -1017 3333 -983
rect 3367 -1017 3401 -983
rect 3435 -1017 3469 -983
rect 3503 -1017 3537 -983
rect 3571 -1017 3605 -983
rect 3639 -1017 3673 -983
rect 3707 -1017 3741 -983
rect 3775 -1017 3809 -983
rect 3843 -1017 3877 -983
rect 3911 -1017 3945 -983
rect 3979 -1017 4013 -983
rect 4047 -1017 4081 -983
rect 4115 -1017 4149 -983
rect 4183 -1017 4217 -983
rect 4251 -1017 4285 -983
rect 4319 -1017 4353 -983
rect 4387 -1017 4421 -983
rect 4455 -1017 4489 -983
rect 4523 -1017 4557 -983
rect 4591 -1017 4625 -983
rect 4659 -1017 4693 -983
rect 4727 -1017 4761 -983
rect 4795 -1017 4829 -983
rect 4863 -1017 4897 -983
rect 4931 -1017 4965 -983
rect 4999 -1017 5033 -983
rect 5067 -1017 5101 -983
rect 5135 -1017 5169 -983
rect 5203 -1017 5237 -983
rect 5271 -1017 5305 -983
rect 5339 -1017 5373 -983
rect 5407 -1017 5441 -983
rect 5475 -1017 5509 -983
rect 5543 -1017 5577 -983
rect 5611 -1017 5645 -983
rect 5679 -1017 5713 -983
rect 5747 -1017 5781 -983
rect 5815 -1017 5849 -983
rect 5883 -1017 5917 -983
rect 5951 -1017 5985 -983
rect 6019 -1017 6053 -983
rect 6087 -1017 6121 -983
rect 6155 -1017 6189 -983
rect 6223 -1017 6257 -983
rect 6291 -1017 6325 -983
rect 6359 -1017 6393 -983
rect 6427 -1017 6461 -983
rect 6495 -1017 6529 -983
rect 6563 -1017 6597 -983
rect 6631 -1017 6665 -983
rect 6699 -1017 6733 -983
rect 6767 -1017 6801 -983
rect 6835 -1017 6869 -983
rect 6903 -1017 6937 -983
rect 6971 -1017 7005 -983
rect 7039 -1017 7073 -983
rect 7107 -1017 7141 -983
rect 7175 -1017 7209 -983
rect 7243 -1017 7277 -983
rect 7311 -1017 7345 -983
rect 7379 -1017 7413 -983
rect 7447 -1017 7481 -983
rect 7515 -1017 7549 -983
rect 7583 -1017 7617 -983
rect 7651 -1017 7685 -983
rect 7719 -1017 7753 -983
rect 7787 -1017 7821 -983
rect 7855 -1017 7889 -983
rect 7923 -1017 7957 -983
rect 7991 -1017 8025 -983
rect 8059 -1017 8093 -983
rect 8127 -1017 8161 -983
rect 8195 -1017 8229 -983
rect 8263 -1017 8400 -983
rect 0 -1040 8400 -1017
<< mvnsubdiff >>
rect 160 9897 8240 9920
rect 160 9863 307 9897
rect 341 9863 375 9897
rect 409 9863 443 9897
rect 477 9863 511 9897
rect 545 9863 579 9897
rect 613 9863 647 9897
rect 681 9863 715 9897
rect 749 9863 783 9897
rect 817 9863 851 9897
rect 885 9863 919 9897
rect 953 9863 987 9897
rect 1021 9863 1055 9897
rect 1089 9863 1123 9897
rect 1157 9863 1191 9897
rect 1225 9863 1259 9897
rect 1293 9863 1327 9897
rect 1361 9863 1395 9897
rect 1429 9863 1463 9897
rect 1497 9863 1531 9897
rect 1565 9863 1599 9897
rect 1633 9863 1667 9897
rect 1701 9863 1735 9897
rect 1769 9863 1803 9897
rect 1837 9863 1871 9897
rect 1905 9863 1939 9897
rect 1973 9863 2007 9897
rect 2041 9863 2075 9897
rect 2109 9863 2143 9897
rect 2177 9863 2211 9897
rect 2245 9863 2279 9897
rect 2313 9863 2347 9897
rect 2381 9863 2415 9897
rect 2449 9863 2483 9897
rect 2517 9863 2551 9897
rect 2585 9863 2619 9897
rect 2653 9863 2687 9897
rect 2721 9863 2755 9897
rect 2789 9863 2823 9897
rect 2857 9863 2891 9897
rect 2925 9863 2959 9897
rect 2993 9863 3027 9897
rect 3061 9863 3095 9897
rect 3129 9863 3163 9897
rect 3197 9863 3231 9897
rect 3265 9863 3299 9897
rect 3333 9863 3367 9897
rect 3401 9863 3435 9897
rect 3469 9863 3503 9897
rect 3537 9863 3571 9897
rect 3605 9863 3639 9897
rect 3673 9863 3707 9897
rect 3741 9863 3775 9897
rect 3809 9863 3843 9897
rect 3877 9863 3911 9897
rect 3945 9863 3979 9897
rect 4013 9863 4047 9897
rect 4081 9863 4115 9897
rect 4149 9863 4183 9897
rect 4217 9863 4251 9897
rect 4285 9863 4319 9897
rect 4353 9863 4387 9897
rect 4421 9863 4455 9897
rect 4489 9863 4523 9897
rect 4557 9863 4591 9897
rect 4625 9863 4659 9897
rect 4693 9863 4727 9897
rect 4761 9863 4795 9897
rect 4829 9863 4863 9897
rect 4897 9863 4931 9897
rect 4965 9863 4999 9897
rect 5033 9863 5067 9897
rect 5101 9863 5135 9897
rect 5169 9863 5203 9897
rect 5237 9863 5271 9897
rect 5305 9863 5339 9897
rect 5373 9863 5407 9897
rect 5441 9863 5475 9897
rect 5509 9863 5543 9897
rect 5577 9863 5611 9897
rect 5645 9863 5679 9897
rect 5713 9863 5747 9897
rect 5781 9863 5815 9897
rect 5849 9863 5883 9897
rect 5917 9863 5951 9897
rect 5985 9863 6019 9897
rect 6053 9863 6087 9897
rect 6121 9863 6155 9897
rect 6189 9863 6223 9897
rect 6257 9863 6291 9897
rect 6325 9863 6359 9897
rect 6393 9863 6427 9897
rect 6461 9863 6495 9897
rect 6529 9863 6563 9897
rect 6597 9863 6631 9897
rect 6665 9863 6699 9897
rect 6733 9863 6767 9897
rect 6801 9863 6835 9897
rect 6869 9863 6903 9897
rect 6937 9863 6971 9897
rect 7005 9863 7039 9897
rect 7073 9863 7107 9897
rect 7141 9863 7175 9897
rect 7209 9863 7243 9897
rect 7277 9863 7311 9897
rect 7345 9863 7379 9897
rect 7413 9863 7447 9897
rect 7481 9863 7515 9897
rect 7549 9863 7583 9897
rect 7617 9863 7651 9897
rect 7685 9863 7719 9897
rect 7753 9863 7787 9897
rect 7821 9863 7855 9897
rect 7889 9863 7923 9897
rect 7957 9863 7991 9897
rect 8025 9863 8059 9897
rect 8093 9863 8240 9897
rect 160 9840 8240 9863
rect 160 9791 240 9840
rect 160 9757 183 9791
rect 217 9757 240 9791
rect 8160 9791 8240 9840
rect 160 9723 240 9757
rect 160 9689 183 9723
rect 217 9689 240 9723
rect 160 9655 240 9689
rect 160 9621 183 9655
rect 217 9621 240 9655
rect 160 9587 240 9621
rect 160 9553 183 9587
rect 217 9553 240 9587
rect 160 9519 240 9553
rect 160 9485 183 9519
rect 217 9485 240 9519
rect 160 9451 240 9485
rect 160 9417 183 9451
rect 217 9417 240 9451
rect 160 9383 240 9417
rect 160 9349 183 9383
rect 217 9349 240 9383
rect 160 9315 240 9349
rect 160 9281 183 9315
rect 217 9281 240 9315
rect 160 9247 240 9281
rect 160 9213 183 9247
rect 217 9213 240 9247
rect 160 9179 240 9213
rect 160 9145 183 9179
rect 217 9145 240 9179
rect 8160 9757 8183 9791
rect 8217 9757 8240 9791
rect 8160 9723 8240 9757
rect 8160 9689 8183 9723
rect 8217 9689 8240 9723
rect 8160 9655 8240 9689
rect 8160 9621 8183 9655
rect 8217 9621 8240 9655
rect 8160 9587 8240 9621
rect 8160 9553 8183 9587
rect 8217 9553 8240 9587
rect 8160 9519 8240 9553
rect 8160 9485 8183 9519
rect 8217 9485 8240 9519
rect 8160 9451 8240 9485
rect 8160 9417 8183 9451
rect 8217 9417 8240 9451
rect 8160 9383 8240 9417
rect 8160 9349 8183 9383
rect 8217 9349 8240 9383
rect 8160 9315 8240 9349
rect 8160 9281 8183 9315
rect 8217 9281 8240 9315
rect 8160 9247 8240 9281
rect 8160 9213 8183 9247
rect 8217 9213 8240 9247
rect 8160 9179 8240 9213
rect 160 9111 240 9145
rect 160 9077 183 9111
rect 217 9077 240 9111
rect 160 9043 240 9077
rect 160 9009 183 9043
rect 217 9009 240 9043
rect 8160 9145 8183 9179
rect 8217 9145 8240 9179
rect 8160 9111 8240 9145
rect 8160 9077 8183 9111
rect 8217 9077 8240 9111
rect 8160 9043 8240 9077
rect 160 8960 240 9009
rect 8160 9009 8183 9043
rect 8217 9009 8240 9043
rect 8160 8960 8240 9009
rect 160 8937 8240 8960
rect 160 8903 307 8937
rect 341 8903 375 8937
rect 409 8903 443 8937
rect 477 8903 511 8937
rect 545 8903 579 8937
rect 613 8903 647 8937
rect 681 8903 715 8937
rect 749 8903 783 8937
rect 817 8903 851 8937
rect 885 8903 919 8937
rect 953 8903 987 8937
rect 1021 8903 1055 8937
rect 1089 8903 1123 8937
rect 1157 8903 1191 8937
rect 1225 8903 1259 8937
rect 1293 8903 1327 8937
rect 1361 8903 1395 8937
rect 1429 8903 1463 8937
rect 1497 8903 1531 8937
rect 1565 8903 1599 8937
rect 1633 8903 1667 8937
rect 1701 8903 1735 8937
rect 1769 8903 1803 8937
rect 1837 8903 1871 8937
rect 1905 8903 1939 8937
rect 1973 8903 2007 8937
rect 2041 8903 2075 8937
rect 2109 8903 2143 8937
rect 2177 8903 2211 8937
rect 2245 8903 2279 8937
rect 2313 8903 2347 8937
rect 2381 8903 2415 8937
rect 2449 8903 2483 8937
rect 2517 8903 2551 8937
rect 2585 8903 2619 8937
rect 2653 8903 2687 8937
rect 2721 8903 2755 8937
rect 2789 8903 2823 8937
rect 2857 8903 2891 8937
rect 2925 8903 2959 8937
rect 2993 8903 3027 8937
rect 3061 8903 3095 8937
rect 3129 8903 3163 8937
rect 3197 8903 3231 8937
rect 3265 8903 3299 8937
rect 3333 8903 3367 8937
rect 3401 8903 3435 8937
rect 3469 8903 3503 8937
rect 3537 8903 3571 8937
rect 3605 8903 3639 8937
rect 3673 8903 3707 8937
rect 3741 8903 3775 8937
rect 3809 8903 3843 8937
rect 3877 8903 3911 8937
rect 3945 8903 3979 8937
rect 4013 8903 4047 8937
rect 4081 8903 4115 8937
rect 4149 8903 4183 8937
rect 4217 8903 4251 8937
rect 4285 8903 4319 8937
rect 4353 8903 4387 8937
rect 4421 8903 4455 8937
rect 4489 8903 4523 8937
rect 4557 8903 4591 8937
rect 4625 8903 4659 8937
rect 4693 8903 4727 8937
rect 4761 8903 4795 8937
rect 4829 8903 4863 8937
rect 4897 8903 4931 8937
rect 4965 8903 4999 8937
rect 5033 8903 5067 8937
rect 5101 8903 5135 8937
rect 5169 8903 5203 8937
rect 5237 8903 5271 8937
rect 5305 8903 5339 8937
rect 5373 8903 5407 8937
rect 5441 8903 5475 8937
rect 5509 8903 5543 8937
rect 5577 8903 5611 8937
rect 5645 8903 5679 8937
rect 5713 8903 5747 8937
rect 5781 8903 5815 8937
rect 5849 8903 5883 8937
rect 5917 8903 5951 8937
rect 5985 8903 6019 8937
rect 6053 8903 6087 8937
rect 6121 8903 6155 8937
rect 6189 8903 6223 8937
rect 6257 8903 6291 8937
rect 6325 8903 6359 8937
rect 6393 8903 6427 8937
rect 6461 8903 6495 8937
rect 6529 8903 6563 8937
rect 6597 8903 6631 8937
rect 6665 8903 6699 8937
rect 6733 8903 6767 8937
rect 6801 8903 6835 8937
rect 6869 8903 6903 8937
rect 6937 8903 6971 8937
rect 7005 8903 7039 8937
rect 7073 8903 7107 8937
rect 7141 8903 7175 8937
rect 7209 8903 7243 8937
rect 7277 8903 7311 8937
rect 7345 8903 7379 8937
rect 7413 8903 7447 8937
rect 7481 8903 7515 8937
rect 7549 8903 7583 8937
rect 7617 8903 7651 8937
rect 7685 8903 7719 8937
rect 7753 8903 7787 8937
rect 7821 8903 7855 8937
rect 7889 8903 7923 8937
rect 7957 8903 7991 8937
rect 8025 8903 8059 8937
rect 8093 8903 8240 8937
rect 160 8880 8240 8903
rect 160 5257 8240 5280
rect 160 5223 307 5257
rect 341 5223 375 5257
rect 409 5223 443 5257
rect 477 5223 511 5257
rect 545 5223 579 5257
rect 613 5223 647 5257
rect 681 5223 715 5257
rect 749 5223 783 5257
rect 817 5223 851 5257
rect 885 5223 919 5257
rect 953 5223 987 5257
rect 1021 5223 1055 5257
rect 1089 5223 1123 5257
rect 1157 5223 1191 5257
rect 1225 5223 1259 5257
rect 1293 5223 1327 5257
rect 1361 5223 1395 5257
rect 1429 5223 1463 5257
rect 1497 5223 1531 5257
rect 1565 5223 1599 5257
rect 1633 5223 1667 5257
rect 1701 5223 1735 5257
rect 1769 5223 1803 5257
rect 1837 5223 1871 5257
rect 1905 5223 1939 5257
rect 1973 5223 2007 5257
rect 2041 5223 2075 5257
rect 2109 5223 2143 5257
rect 2177 5223 2211 5257
rect 2245 5223 2279 5257
rect 2313 5223 2347 5257
rect 2381 5223 2415 5257
rect 2449 5223 2483 5257
rect 2517 5223 2551 5257
rect 2585 5223 2619 5257
rect 2653 5223 2687 5257
rect 2721 5223 2755 5257
rect 2789 5223 2823 5257
rect 2857 5223 2891 5257
rect 2925 5223 2959 5257
rect 2993 5223 3027 5257
rect 3061 5223 3095 5257
rect 3129 5223 3163 5257
rect 3197 5223 3231 5257
rect 3265 5223 3299 5257
rect 3333 5223 3367 5257
rect 3401 5223 3435 5257
rect 3469 5223 3503 5257
rect 3537 5223 3571 5257
rect 3605 5223 3639 5257
rect 3673 5223 3707 5257
rect 3741 5223 3775 5257
rect 3809 5223 3843 5257
rect 3877 5223 3911 5257
rect 3945 5223 3979 5257
rect 4013 5223 4047 5257
rect 4081 5223 4115 5257
rect 4149 5223 4183 5257
rect 4217 5223 4251 5257
rect 4285 5223 4319 5257
rect 4353 5223 4387 5257
rect 4421 5223 4455 5257
rect 4489 5223 4523 5257
rect 4557 5223 4591 5257
rect 4625 5223 4659 5257
rect 4693 5223 4727 5257
rect 4761 5223 4795 5257
rect 4829 5223 4863 5257
rect 4897 5223 4931 5257
rect 4965 5223 4999 5257
rect 5033 5223 5067 5257
rect 5101 5223 5135 5257
rect 5169 5223 5203 5257
rect 5237 5223 5271 5257
rect 5305 5223 5339 5257
rect 5373 5223 5407 5257
rect 5441 5223 5475 5257
rect 5509 5223 5543 5257
rect 5577 5223 5611 5257
rect 5645 5223 5679 5257
rect 5713 5223 5747 5257
rect 5781 5223 5815 5257
rect 5849 5223 5883 5257
rect 5917 5223 5951 5257
rect 5985 5223 6019 5257
rect 6053 5223 6087 5257
rect 6121 5223 6155 5257
rect 6189 5223 6223 5257
rect 6257 5223 6291 5257
rect 6325 5223 6359 5257
rect 6393 5223 6427 5257
rect 6461 5223 6495 5257
rect 6529 5223 6563 5257
rect 6597 5223 6631 5257
rect 6665 5223 6699 5257
rect 6733 5223 6767 5257
rect 6801 5223 6835 5257
rect 6869 5223 6903 5257
rect 6937 5223 6971 5257
rect 7005 5223 7039 5257
rect 7073 5223 7107 5257
rect 7141 5223 7175 5257
rect 7209 5223 7243 5257
rect 7277 5223 7311 5257
rect 7345 5223 7379 5257
rect 7413 5223 7447 5257
rect 7481 5223 7515 5257
rect 7549 5223 7583 5257
rect 7617 5223 7651 5257
rect 7685 5223 7719 5257
rect 7753 5223 7787 5257
rect 7821 5223 7855 5257
rect 7889 5223 7923 5257
rect 7957 5223 7991 5257
rect 8025 5223 8059 5257
rect 8093 5223 8240 5257
rect 160 5200 8240 5223
rect 160 5151 240 5200
rect 160 5117 183 5151
rect 217 5117 240 5151
rect 8160 5151 8240 5200
rect 160 5083 240 5117
rect 160 5049 183 5083
rect 217 5049 240 5083
rect 160 5015 240 5049
rect 160 4981 183 5015
rect 217 4981 240 5015
rect 8160 5117 8183 5151
rect 8217 5117 8240 5151
rect 8160 5083 8240 5117
rect 8160 5049 8183 5083
rect 8217 5049 8240 5083
rect 8160 5015 8240 5049
rect 160 4947 240 4981
rect 160 4913 183 4947
rect 217 4913 240 4947
rect 160 4879 240 4913
rect 160 4845 183 4879
rect 217 4845 240 4879
rect 160 4811 240 4845
rect 160 4777 183 4811
rect 217 4777 240 4811
rect 160 4743 240 4777
rect 160 4709 183 4743
rect 217 4709 240 4743
rect 160 4675 240 4709
rect 160 4641 183 4675
rect 217 4641 240 4675
rect 160 4607 240 4641
rect 160 4573 183 4607
rect 217 4573 240 4607
rect 160 4539 240 4573
rect 160 4505 183 4539
rect 217 4505 240 4539
rect 160 4471 240 4505
rect 160 4437 183 4471
rect 217 4437 240 4471
rect 160 4403 240 4437
rect 160 4369 183 4403
rect 217 4369 240 4403
rect 8160 4981 8183 5015
rect 8217 4981 8240 5015
rect 8160 4947 8240 4981
rect 8160 4913 8183 4947
rect 8217 4913 8240 4947
rect 8160 4879 8240 4913
rect 8160 4845 8183 4879
rect 8217 4845 8240 4879
rect 8160 4811 8240 4845
rect 8160 4777 8183 4811
rect 8217 4777 8240 4811
rect 8160 4743 8240 4777
rect 8160 4709 8183 4743
rect 8217 4709 8240 4743
rect 8160 4675 8240 4709
rect 8160 4641 8183 4675
rect 8217 4641 8240 4675
rect 8160 4607 8240 4641
rect 8160 4573 8183 4607
rect 8217 4573 8240 4607
rect 8160 4539 8240 4573
rect 8160 4505 8183 4539
rect 8217 4505 8240 4539
rect 8160 4471 8240 4505
rect 8160 4437 8183 4471
rect 8217 4437 8240 4471
rect 8160 4403 8240 4437
rect 160 4320 240 4369
rect 8160 4369 8183 4403
rect 8217 4369 8240 4403
rect 8160 4320 8240 4369
rect 160 4297 8240 4320
rect 160 4263 307 4297
rect 341 4263 375 4297
rect 409 4263 443 4297
rect 477 4263 511 4297
rect 545 4263 579 4297
rect 613 4263 647 4297
rect 681 4263 715 4297
rect 749 4263 783 4297
rect 817 4263 851 4297
rect 885 4263 919 4297
rect 953 4263 987 4297
rect 1021 4263 1055 4297
rect 1089 4263 1123 4297
rect 1157 4263 1191 4297
rect 1225 4263 1259 4297
rect 1293 4263 1327 4297
rect 1361 4263 1395 4297
rect 1429 4263 1463 4297
rect 1497 4263 1531 4297
rect 1565 4263 1599 4297
rect 1633 4263 1667 4297
rect 1701 4263 1735 4297
rect 1769 4263 1803 4297
rect 1837 4263 1871 4297
rect 1905 4263 1939 4297
rect 1973 4263 2007 4297
rect 2041 4263 2075 4297
rect 2109 4263 2143 4297
rect 2177 4263 2211 4297
rect 2245 4263 2279 4297
rect 2313 4263 2347 4297
rect 2381 4263 2415 4297
rect 2449 4263 2483 4297
rect 2517 4263 2551 4297
rect 2585 4263 2619 4297
rect 2653 4263 2687 4297
rect 2721 4263 2755 4297
rect 2789 4263 2823 4297
rect 2857 4263 2891 4297
rect 2925 4263 2959 4297
rect 2993 4263 3027 4297
rect 3061 4263 3095 4297
rect 3129 4263 3163 4297
rect 3197 4263 3231 4297
rect 3265 4263 3299 4297
rect 3333 4263 3367 4297
rect 3401 4263 3435 4297
rect 3469 4263 3503 4297
rect 3537 4263 3571 4297
rect 3605 4263 3639 4297
rect 3673 4263 3707 4297
rect 3741 4263 3775 4297
rect 3809 4263 3843 4297
rect 3877 4263 3911 4297
rect 3945 4263 3979 4297
rect 4013 4263 4047 4297
rect 4081 4263 4115 4297
rect 4149 4263 4183 4297
rect 4217 4263 4251 4297
rect 4285 4263 4319 4297
rect 4353 4263 4387 4297
rect 4421 4263 4455 4297
rect 4489 4263 4523 4297
rect 4557 4263 4591 4297
rect 4625 4263 4659 4297
rect 4693 4263 4727 4297
rect 4761 4263 4795 4297
rect 4829 4263 4863 4297
rect 4897 4263 4931 4297
rect 4965 4263 4999 4297
rect 5033 4263 5067 4297
rect 5101 4263 5135 4297
rect 5169 4263 5203 4297
rect 5237 4263 5271 4297
rect 5305 4263 5339 4297
rect 5373 4263 5407 4297
rect 5441 4263 5475 4297
rect 5509 4263 5543 4297
rect 5577 4263 5611 4297
rect 5645 4263 5679 4297
rect 5713 4263 5747 4297
rect 5781 4263 5815 4297
rect 5849 4263 5883 4297
rect 5917 4263 5951 4297
rect 5985 4263 6019 4297
rect 6053 4263 6087 4297
rect 6121 4263 6155 4297
rect 6189 4263 6223 4297
rect 6257 4263 6291 4297
rect 6325 4263 6359 4297
rect 6393 4263 6427 4297
rect 6461 4263 6495 4297
rect 6529 4263 6563 4297
rect 6597 4263 6631 4297
rect 6665 4263 6699 4297
rect 6733 4263 6767 4297
rect 6801 4263 6835 4297
rect 6869 4263 6903 4297
rect 6937 4263 6971 4297
rect 7005 4263 7039 4297
rect 7073 4263 7107 4297
rect 7141 4263 7175 4297
rect 7209 4263 7243 4297
rect 7277 4263 7311 4297
rect 7345 4263 7379 4297
rect 7413 4263 7447 4297
rect 7481 4263 7515 4297
rect 7549 4263 7583 4297
rect 7617 4263 7651 4297
rect 7685 4263 7719 4297
rect 7753 4263 7787 4297
rect 7821 4263 7855 4297
rect 7889 4263 7923 4297
rect 7957 4263 7991 4297
rect 8025 4263 8059 4297
rect 8093 4263 8240 4297
rect 160 4240 8240 4263
rect 160 3817 8240 3840
rect 160 3783 307 3817
rect 341 3783 375 3817
rect 409 3783 443 3817
rect 477 3783 511 3817
rect 545 3783 579 3817
rect 613 3783 647 3817
rect 681 3783 715 3817
rect 749 3783 783 3817
rect 817 3783 851 3817
rect 885 3783 919 3817
rect 953 3783 987 3817
rect 1021 3783 1055 3817
rect 1089 3783 1123 3817
rect 1157 3783 1191 3817
rect 1225 3783 1259 3817
rect 1293 3783 1327 3817
rect 1361 3783 1395 3817
rect 1429 3783 1463 3817
rect 1497 3783 1531 3817
rect 1565 3783 1599 3817
rect 1633 3783 1667 3817
rect 1701 3783 1735 3817
rect 1769 3783 1803 3817
rect 1837 3783 1871 3817
rect 1905 3783 1939 3817
rect 1973 3783 2007 3817
rect 2041 3783 2075 3817
rect 2109 3783 2143 3817
rect 2177 3783 2211 3817
rect 2245 3783 2279 3817
rect 2313 3783 2347 3817
rect 2381 3783 2415 3817
rect 2449 3783 2483 3817
rect 2517 3783 2551 3817
rect 2585 3783 2619 3817
rect 2653 3783 2687 3817
rect 2721 3783 2755 3817
rect 2789 3783 2823 3817
rect 2857 3783 2891 3817
rect 2925 3783 2959 3817
rect 2993 3783 3027 3817
rect 3061 3783 3095 3817
rect 3129 3783 3163 3817
rect 3197 3783 3231 3817
rect 3265 3783 3299 3817
rect 3333 3783 3367 3817
rect 3401 3783 3435 3817
rect 3469 3783 3503 3817
rect 3537 3783 3571 3817
rect 3605 3783 3639 3817
rect 3673 3783 3707 3817
rect 3741 3783 3775 3817
rect 3809 3783 3843 3817
rect 3877 3783 3911 3817
rect 3945 3783 3979 3817
rect 4013 3783 4047 3817
rect 4081 3783 4115 3817
rect 4149 3783 4183 3817
rect 4217 3783 4251 3817
rect 4285 3783 4319 3817
rect 4353 3783 4387 3817
rect 4421 3783 4455 3817
rect 4489 3783 4523 3817
rect 4557 3783 4591 3817
rect 4625 3783 4659 3817
rect 4693 3783 4727 3817
rect 4761 3783 4795 3817
rect 4829 3783 4863 3817
rect 4897 3783 4931 3817
rect 4965 3783 4999 3817
rect 5033 3783 5067 3817
rect 5101 3783 5135 3817
rect 5169 3783 5203 3817
rect 5237 3783 5271 3817
rect 5305 3783 5339 3817
rect 5373 3783 5407 3817
rect 5441 3783 5475 3817
rect 5509 3783 5543 3817
rect 5577 3783 5611 3817
rect 5645 3783 5679 3817
rect 5713 3783 5747 3817
rect 5781 3783 5815 3817
rect 5849 3783 5883 3817
rect 5917 3783 5951 3817
rect 5985 3783 6019 3817
rect 6053 3783 6087 3817
rect 6121 3783 6155 3817
rect 6189 3783 6223 3817
rect 6257 3783 6291 3817
rect 6325 3783 6359 3817
rect 6393 3783 6427 3817
rect 6461 3783 6495 3817
rect 6529 3783 6563 3817
rect 6597 3783 6631 3817
rect 6665 3783 6699 3817
rect 6733 3783 6767 3817
rect 6801 3783 6835 3817
rect 6869 3783 6903 3817
rect 6937 3783 6971 3817
rect 7005 3783 7039 3817
rect 7073 3783 7107 3817
rect 7141 3783 7175 3817
rect 7209 3783 7243 3817
rect 7277 3783 7311 3817
rect 7345 3783 7379 3817
rect 7413 3783 7447 3817
rect 7481 3783 7515 3817
rect 7549 3783 7583 3817
rect 7617 3783 7651 3817
rect 7685 3783 7719 3817
rect 7753 3783 7787 3817
rect 7821 3783 7855 3817
rect 7889 3783 7923 3817
rect 7957 3783 7991 3817
rect 8025 3783 8059 3817
rect 8093 3783 8240 3817
rect 160 3760 8240 3783
rect 160 3711 240 3760
rect 160 3677 183 3711
rect 217 3677 240 3711
rect 8160 3711 8240 3760
rect 160 3643 240 3677
rect 160 3609 183 3643
rect 217 3609 240 3643
rect 160 3575 240 3609
rect 160 3541 183 3575
rect 217 3541 240 3575
rect 160 3507 240 3541
rect 160 3473 183 3507
rect 217 3473 240 3507
rect 160 3439 240 3473
rect 160 3405 183 3439
rect 217 3405 240 3439
rect 160 3371 240 3405
rect 160 3337 183 3371
rect 217 3337 240 3371
rect 160 3303 240 3337
rect 160 3269 183 3303
rect 217 3269 240 3303
rect 160 3235 240 3269
rect 160 3201 183 3235
rect 217 3201 240 3235
rect 160 3167 240 3201
rect 160 3133 183 3167
rect 217 3133 240 3167
rect 160 3099 240 3133
rect 160 3065 183 3099
rect 217 3065 240 3099
rect 8160 3677 8183 3711
rect 8217 3677 8240 3711
rect 8160 3643 8240 3677
rect 8160 3609 8183 3643
rect 8217 3609 8240 3643
rect 8160 3575 8240 3609
rect 8160 3541 8183 3575
rect 8217 3541 8240 3575
rect 8160 3507 8240 3541
rect 8160 3473 8183 3507
rect 8217 3473 8240 3507
rect 8160 3439 8240 3473
rect 8160 3405 8183 3439
rect 8217 3405 8240 3439
rect 8160 3371 8240 3405
rect 8160 3337 8183 3371
rect 8217 3337 8240 3371
rect 8160 3303 8240 3337
rect 8160 3269 8183 3303
rect 8217 3269 8240 3303
rect 8160 3235 8240 3269
rect 8160 3201 8183 3235
rect 8217 3201 8240 3235
rect 8160 3167 8240 3201
rect 8160 3133 8183 3167
rect 8217 3133 8240 3167
rect 8160 3099 8240 3133
rect 160 3031 240 3065
rect 160 2997 183 3031
rect 217 2997 240 3031
rect 160 2963 240 2997
rect 160 2929 183 2963
rect 217 2929 240 2963
rect 8160 3065 8183 3099
rect 8217 3065 8240 3099
rect 8160 3031 8240 3065
rect 8160 2997 8183 3031
rect 8217 2997 8240 3031
rect 8160 2963 8240 2997
rect 160 2880 240 2929
rect 8160 2929 8183 2963
rect 8217 2929 8240 2963
rect 8160 2880 8240 2929
rect 160 2857 8240 2880
rect 160 2823 307 2857
rect 341 2823 375 2857
rect 409 2823 443 2857
rect 477 2823 511 2857
rect 545 2823 579 2857
rect 613 2823 647 2857
rect 681 2823 715 2857
rect 749 2823 783 2857
rect 817 2823 851 2857
rect 885 2823 919 2857
rect 953 2823 987 2857
rect 1021 2823 1055 2857
rect 1089 2823 1123 2857
rect 1157 2823 1191 2857
rect 1225 2823 1259 2857
rect 1293 2823 1327 2857
rect 1361 2823 1395 2857
rect 1429 2823 1463 2857
rect 1497 2823 1531 2857
rect 1565 2823 1599 2857
rect 1633 2823 1667 2857
rect 1701 2823 1735 2857
rect 1769 2823 1803 2857
rect 1837 2823 1871 2857
rect 1905 2823 1939 2857
rect 1973 2823 2007 2857
rect 2041 2823 2075 2857
rect 2109 2823 2143 2857
rect 2177 2823 2211 2857
rect 2245 2823 2279 2857
rect 2313 2823 2347 2857
rect 2381 2823 2415 2857
rect 2449 2823 2483 2857
rect 2517 2823 2551 2857
rect 2585 2823 2619 2857
rect 2653 2823 2687 2857
rect 2721 2823 2755 2857
rect 2789 2823 2823 2857
rect 2857 2823 2891 2857
rect 2925 2823 2959 2857
rect 2993 2823 3027 2857
rect 3061 2823 3095 2857
rect 3129 2823 3163 2857
rect 3197 2823 3231 2857
rect 3265 2823 3299 2857
rect 3333 2823 3367 2857
rect 3401 2823 3435 2857
rect 3469 2823 3503 2857
rect 3537 2823 3571 2857
rect 3605 2823 3639 2857
rect 3673 2823 3707 2857
rect 3741 2823 3775 2857
rect 3809 2823 3843 2857
rect 3877 2823 3911 2857
rect 3945 2823 3979 2857
rect 4013 2823 4047 2857
rect 4081 2823 4115 2857
rect 4149 2823 4183 2857
rect 4217 2823 4251 2857
rect 4285 2823 4319 2857
rect 4353 2823 4387 2857
rect 4421 2823 4455 2857
rect 4489 2823 4523 2857
rect 4557 2823 4591 2857
rect 4625 2823 4659 2857
rect 4693 2823 4727 2857
rect 4761 2823 4795 2857
rect 4829 2823 4863 2857
rect 4897 2823 4931 2857
rect 4965 2823 4999 2857
rect 5033 2823 5067 2857
rect 5101 2823 5135 2857
rect 5169 2823 5203 2857
rect 5237 2823 5271 2857
rect 5305 2823 5339 2857
rect 5373 2823 5407 2857
rect 5441 2823 5475 2857
rect 5509 2823 5543 2857
rect 5577 2823 5611 2857
rect 5645 2823 5679 2857
rect 5713 2823 5747 2857
rect 5781 2823 5815 2857
rect 5849 2823 5883 2857
rect 5917 2823 5951 2857
rect 5985 2823 6019 2857
rect 6053 2823 6087 2857
rect 6121 2823 6155 2857
rect 6189 2823 6223 2857
rect 6257 2823 6291 2857
rect 6325 2823 6359 2857
rect 6393 2823 6427 2857
rect 6461 2823 6495 2857
rect 6529 2823 6563 2857
rect 6597 2823 6631 2857
rect 6665 2823 6699 2857
rect 6733 2823 6767 2857
rect 6801 2823 6835 2857
rect 6869 2823 6903 2857
rect 6937 2823 6971 2857
rect 7005 2823 7039 2857
rect 7073 2823 7107 2857
rect 7141 2823 7175 2857
rect 7209 2823 7243 2857
rect 7277 2823 7311 2857
rect 7345 2823 7379 2857
rect 7413 2823 7447 2857
rect 7481 2823 7515 2857
rect 7549 2823 7583 2857
rect 7617 2823 7651 2857
rect 7685 2823 7719 2857
rect 7753 2823 7787 2857
rect 7821 2823 7855 2857
rect 7889 2823 7923 2857
rect 7957 2823 7991 2857
rect 8025 2823 8059 2857
rect 8093 2823 8240 2857
rect 160 2800 8240 2823
rect 160 2377 8240 2400
rect 160 2343 307 2377
rect 341 2343 375 2377
rect 409 2343 443 2377
rect 477 2343 511 2377
rect 545 2343 579 2377
rect 613 2343 647 2377
rect 681 2343 715 2377
rect 749 2343 783 2377
rect 817 2343 851 2377
rect 885 2343 919 2377
rect 953 2343 987 2377
rect 1021 2343 1055 2377
rect 1089 2343 1123 2377
rect 1157 2343 1191 2377
rect 1225 2343 1259 2377
rect 1293 2343 1327 2377
rect 1361 2343 1395 2377
rect 1429 2343 1463 2377
rect 1497 2343 1531 2377
rect 1565 2343 1599 2377
rect 1633 2343 1667 2377
rect 1701 2343 1735 2377
rect 1769 2343 1803 2377
rect 1837 2343 1871 2377
rect 1905 2343 1939 2377
rect 1973 2343 2007 2377
rect 2041 2343 2075 2377
rect 2109 2343 2143 2377
rect 2177 2343 2211 2377
rect 2245 2343 2279 2377
rect 2313 2343 2347 2377
rect 2381 2343 2415 2377
rect 2449 2343 2483 2377
rect 2517 2343 2551 2377
rect 2585 2343 2619 2377
rect 2653 2343 2687 2377
rect 2721 2343 2755 2377
rect 2789 2343 2823 2377
rect 2857 2343 2891 2377
rect 2925 2343 2959 2377
rect 2993 2343 3027 2377
rect 3061 2343 3095 2377
rect 3129 2343 3163 2377
rect 3197 2343 3231 2377
rect 3265 2343 3299 2377
rect 3333 2343 3367 2377
rect 3401 2343 3435 2377
rect 3469 2343 3503 2377
rect 3537 2343 3571 2377
rect 3605 2343 3639 2377
rect 3673 2343 3707 2377
rect 3741 2343 3775 2377
rect 3809 2343 3843 2377
rect 3877 2343 3911 2377
rect 3945 2343 3979 2377
rect 4013 2343 4047 2377
rect 4081 2343 4115 2377
rect 4149 2343 4183 2377
rect 4217 2343 4251 2377
rect 4285 2343 4319 2377
rect 4353 2343 4387 2377
rect 4421 2343 4455 2377
rect 4489 2343 4523 2377
rect 4557 2343 4591 2377
rect 4625 2343 4659 2377
rect 4693 2343 4727 2377
rect 4761 2343 4795 2377
rect 4829 2343 4863 2377
rect 4897 2343 4931 2377
rect 4965 2343 4999 2377
rect 5033 2343 5067 2377
rect 5101 2343 5135 2377
rect 5169 2343 5203 2377
rect 5237 2343 5271 2377
rect 5305 2343 5339 2377
rect 5373 2343 5407 2377
rect 5441 2343 5475 2377
rect 5509 2343 5543 2377
rect 5577 2343 5611 2377
rect 5645 2343 5679 2377
rect 5713 2343 5747 2377
rect 5781 2343 5815 2377
rect 5849 2343 5883 2377
rect 5917 2343 5951 2377
rect 5985 2343 6019 2377
rect 6053 2343 6087 2377
rect 6121 2343 6155 2377
rect 6189 2343 6223 2377
rect 6257 2343 6291 2377
rect 6325 2343 6359 2377
rect 6393 2343 6427 2377
rect 6461 2343 6495 2377
rect 6529 2343 6563 2377
rect 6597 2343 6631 2377
rect 6665 2343 6699 2377
rect 6733 2343 6767 2377
rect 6801 2343 6835 2377
rect 6869 2343 6903 2377
rect 6937 2343 6971 2377
rect 7005 2343 7039 2377
rect 7073 2343 7107 2377
rect 7141 2343 7175 2377
rect 7209 2343 7243 2377
rect 7277 2343 7311 2377
rect 7345 2343 7379 2377
rect 7413 2343 7447 2377
rect 7481 2343 7515 2377
rect 7549 2343 7583 2377
rect 7617 2343 7651 2377
rect 7685 2343 7719 2377
rect 7753 2343 7787 2377
rect 7821 2343 7855 2377
rect 7889 2343 7923 2377
rect 7957 2343 7991 2377
rect 8025 2343 8059 2377
rect 8093 2343 8240 2377
rect 160 2320 8240 2343
rect 160 2271 240 2320
rect 160 2237 183 2271
rect 217 2237 240 2271
rect 8160 2271 8240 2320
rect 160 2203 240 2237
rect 160 2169 183 2203
rect 217 2169 240 2203
rect 160 2135 240 2169
rect 160 2101 183 2135
rect 217 2101 240 2135
rect 160 2067 240 2101
rect 160 2033 183 2067
rect 217 2033 240 2067
rect 160 1999 240 2033
rect 160 1965 183 1999
rect 217 1965 240 1999
rect 160 1931 240 1965
rect 160 1897 183 1931
rect 217 1897 240 1931
rect 160 1863 240 1897
rect 160 1829 183 1863
rect 217 1829 240 1863
rect 160 1795 240 1829
rect 160 1761 183 1795
rect 217 1761 240 1795
rect 160 1727 240 1761
rect 160 1693 183 1727
rect 217 1693 240 1727
rect 160 1659 240 1693
rect 160 1625 183 1659
rect 217 1625 240 1659
rect 8160 2237 8183 2271
rect 8217 2237 8240 2271
rect 8160 2203 8240 2237
rect 8160 2169 8183 2203
rect 8217 2169 8240 2203
rect 8160 2135 8240 2169
rect 8160 2101 8183 2135
rect 8217 2101 8240 2135
rect 8160 2067 8240 2101
rect 8160 2033 8183 2067
rect 8217 2033 8240 2067
rect 8160 1999 8240 2033
rect 8160 1965 8183 1999
rect 8217 1965 8240 1999
rect 8160 1931 8240 1965
rect 8160 1897 8183 1931
rect 8217 1897 8240 1931
rect 8160 1863 8240 1897
rect 8160 1829 8183 1863
rect 8217 1829 8240 1863
rect 8160 1795 8240 1829
rect 8160 1761 8183 1795
rect 8217 1761 8240 1795
rect 8160 1727 8240 1761
rect 8160 1693 8183 1727
rect 8217 1693 8240 1727
rect 8160 1659 8240 1693
rect 160 1591 240 1625
rect 160 1557 183 1591
rect 217 1557 240 1591
rect 160 1523 240 1557
rect 160 1489 183 1523
rect 217 1489 240 1523
rect 8160 1625 8183 1659
rect 8217 1625 8240 1659
rect 8160 1591 8240 1625
rect 8160 1557 8183 1591
rect 8217 1557 8240 1591
rect 8160 1523 8240 1557
rect 160 1440 240 1489
rect 8160 1489 8183 1523
rect 8217 1489 8240 1523
rect 8160 1440 8240 1489
rect 160 1417 8240 1440
rect 160 1383 307 1417
rect 341 1383 375 1417
rect 409 1383 443 1417
rect 477 1383 511 1417
rect 545 1383 579 1417
rect 613 1383 647 1417
rect 681 1383 715 1417
rect 749 1383 783 1417
rect 817 1383 851 1417
rect 885 1383 919 1417
rect 953 1383 987 1417
rect 1021 1383 1055 1417
rect 1089 1383 1123 1417
rect 1157 1383 1191 1417
rect 1225 1383 1259 1417
rect 1293 1383 1327 1417
rect 1361 1383 1395 1417
rect 1429 1383 1463 1417
rect 1497 1383 1531 1417
rect 1565 1383 1599 1417
rect 1633 1383 1667 1417
rect 1701 1383 1735 1417
rect 1769 1383 1803 1417
rect 1837 1383 1871 1417
rect 1905 1383 1939 1417
rect 1973 1383 2007 1417
rect 2041 1383 2075 1417
rect 2109 1383 2143 1417
rect 2177 1383 2211 1417
rect 2245 1383 2279 1417
rect 2313 1383 2347 1417
rect 2381 1383 2415 1417
rect 2449 1383 2483 1417
rect 2517 1383 2551 1417
rect 2585 1383 2619 1417
rect 2653 1383 2687 1417
rect 2721 1383 2755 1417
rect 2789 1383 2823 1417
rect 2857 1383 2891 1417
rect 2925 1383 2959 1417
rect 2993 1383 3027 1417
rect 3061 1383 3095 1417
rect 3129 1383 3163 1417
rect 3197 1383 3231 1417
rect 3265 1383 3299 1417
rect 3333 1383 3367 1417
rect 3401 1383 3435 1417
rect 3469 1383 3503 1417
rect 3537 1383 3571 1417
rect 3605 1383 3639 1417
rect 3673 1383 3707 1417
rect 3741 1383 3775 1417
rect 3809 1383 3843 1417
rect 3877 1383 3911 1417
rect 3945 1383 3979 1417
rect 4013 1383 4047 1417
rect 4081 1383 4115 1417
rect 4149 1383 4183 1417
rect 4217 1383 4251 1417
rect 4285 1383 4319 1417
rect 4353 1383 4387 1417
rect 4421 1383 4455 1417
rect 4489 1383 4523 1417
rect 4557 1383 4591 1417
rect 4625 1383 4659 1417
rect 4693 1383 4727 1417
rect 4761 1383 4795 1417
rect 4829 1383 4863 1417
rect 4897 1383 4931 1417
rect 4965 1383 4999 1417
rect 5033 1383 5067 1417
rect 5101 1383 5135 1417
rect 5169 1383 5203 1417
rect 5237 1383 5271 1417
rect 5305 1383 5339 1417
rect 5373 1383 5407 1417
rect 5441 1383 5475 1417
rect 5509 1383 5543 1417
rect 5577 1383 5611 1417
rect 5645 1383 5679 1417
rect 5713 1383 5747 1417
rect 5781 1383 5815 1417
rect 5849 1383 5883 1417
rect 5917 1383 5951 1417
rect 5985 1383 6019 1417
rect 6053 1383 6087 1417
rect 6121 1383 6155 1417
rect 6189 1383 6223 1417
rect 6257 1383 6291 1417
rect 6325 1383 6359 1417
rect 6393 1383 6427 1417
rect 6461 1383 6495 1417
rect 6529 1383 6563 1417
rect 6597 1383 6631 1417
rect 6665 1383 6699 1417
rect 6733 1383 6767 1417
rect 6801 1383 6835 1417
rect 6869 1383 6903 1417
rect 6937 1383 6971 1417
rect 7005 1383 7039 1417
rect 7073 1383 7107 1417
rect 7141 1383 7175 1417
rect 7209 1383 7243 1417
rect 7277 1383 7311 1417
rect 7345 1383 7379 1417
rect 7413 1383 7447 1417
rect 7481 1383 7515 1417
rect 7549 1383 7583 1417
rect 7617 1383 7651 1417
rect 7685 1383 7719 1417
rect 7753 1383 7787 1417
rect 7821 1383 7855 1417
rect 7889 1383 7923 1417
rect 7957 1383 7991 1417
rect 8025 1383 8059 1417
rect 8093 1383 8240 1417
rect 160 1360 8240 1383
<< psubdiffcont >>
rect 137 10023 171 10057
rect 205 10023 239 10057
rect 273 10023 307 10057
rect 341 10023 375 10057
rect 409 10023 443 10057
rect 477 10023 511 10057
rect 545 10023 579 10057
rect 613 10023 647 10057
rect 681 10023 715 10057
rect 749 10023 783 10057
rect 817 10023 851 10057
rect 885 10023 919 10057
rect 953 10023 987 10057
rect 1021 10023 1055 10057
rect 1089 10023 1123 10057
rect 1157 10023 1191 10057
rect 1225 10023 1259 10057
rect 1293 10023 1327 10057
rect 1361 10023 1395 10057
rect 1429 10023 1463 10057
rect 1497 10023 1531 10057
rect 1565 10023 1599 10057
rect 1633 10023 1667 10057
rect 1701 10023 1735 10057
rect 1769 10023 1803 10057
rect 1837 10023 1871 10057
rect 1905 10023 1939 10057
rect 1973 10023 2007 10057
rect 2041 10023 2075 10057
rect 2109 10023 2143 10057
rect 2177 10023 2211 10057
rect 2245 10023 2279 10057
rect 2313 10023 2347 10057
rect 2381 10023 2415 10057
rect 2449 10023 2483 10057
rect 2517 10023 2551 10057
rect 2585 10023 2619 10057
rect 2653 10023 2687 10057
rect 2721 10023 2755 10057
rect 2789 10023 2823 10057
rect 2857 10023 2891 10057
rect 2925 10023 2959 10057
rect 2993 10023 3027 10057
rect 3061 10023 3095 10057
rect 3129 10023 3163 10057
rect 3197 10023 3231 10057
rect 3265 10023 3299 10057
rect 3333 10023 3367 10057
rect 3401 10023 3435 10057
rect 3469 10023 3503 10057
rect 3537 10023 3571 10057
rect 3605 10023 3639 10057
rect 3673 10023 3707 10057
rect 3741 10023 3775 10057
rect 3809 10023 3843 10057
rect 3877 10023 3911 10057
rect 3945 10023 3979 10057
rect 4013 10023 4047 10057
rect 4081 10023 4115 10057
rect 4149 10023 4183 10057
rect 4217 10023 4251 10057
rect 4285 10023 4319 10057
rect 4353 10023 4387 10057
rect 4421 10023 4455 10057
rect 4489 10023 4523 10057
rect 4557 10023 4591 10057
rect 4625 10023 4659 10057
rect 4693 10023 4727 10057
rect 4761 10023 4795 10057
rect 4829 10023 4863 10057
rect 4897 10023 4931 10057
rect 4965 10023 4999 10057
rect 5033 10023 5067 10057
rect 5101 10023 5135 10057
rect 5169 10023 5203 10057
rect 5237 10023 5271 10057
rect 5305 10023 5339 10057
rect 5373 10023 5407 10057
rect 5441 10023 5475 10057
rect 5509 10023 5543 10057
rect 5577 10023 5611 10057
rect 5645 10023 5679 10057
rect 5713 10023 5747 10057
rect 5781 10023 5815 10057
rect 5849 10023 5883 10057
rect 5917 10023 5951 10057
rect 5985 10023 6019 10057
rect 6053 10023 6087 10057
rect 6121 10023 6155 10057
rect 6189 10023 6223 10057
rect 6257 10023 6291 10057
rect 6325 10023 6359 10057
rect 6393 10023 6427 10057
rect 6461 10023 6495 10057
rect 6529 10023 6563 10057
rect 6597 10023 6631 10057
rect 6665 10023 6699 10057
rect 6733 10023 6767 10057
rect 6801 10023 6835 10057
rect 6869 10023 6903 10057
rect 6937 10023 6971 10057
rect 7005 10023 7039 10057
rect 7073 10023 7107 10057
rect 7141 10023 7175 10057
rect 7209 10023 7243 10057
rect 7277 10023 7311 10057
rect 7345 10023 7379 10057
rect 7413 10023 7447 10057
rect 7481 10023 7515 10057
rect 7549 10023 7583 10057
rect 7617 10023 7651 10057
rect 7685 10023 7719 10057
rect 7753 10023 7787 10057
rect 7821 10023 7855 10057
rect 7889 10023 7923 10057
rect 7957 10023 7991 10057
rect 8025 10023 8059 10057
rect 8093 10023 8127 10057
rect 8161 10023 8195 10057
rect 8229 10023 8263 10057
rect 23 9893 57 9927
rect 23 9825 57 9859
rect 23 9757 57 9791
rect 23 9689 57 9723
rect 23 9621 57 9655
rect 23 9553 57 9587
rect 23 9485 57 9519
rect 23 9417 57 9451
rect 23 9349 57 9383
rect 23 9281 57 9315
rect 23 9213 57 9247
rect 23 9145 57 9179
rect 23 9077 57 9111
rect 23 9009 57 9043
rect 23 8941 57 8975
rect 23 8873 57 8907
rect 8343 9893 8377 9927
rect 8343 9825 8377 9859
rect 8343 9757 8377 9791
rect 8343 9689 8377 9723
rect 8343 9621 8377 9655
rect 8343 9553 8377 9587
rect 8343 9485 8377 9519
rect 8343 9417 8377 9451
rect 8343 9349 8377 9383
rect 8343 9281 8377 9315
rect 8343 9213 8377 9247
rect 8343 9145 8377 9179
rect 8343 9077 8377 9111
rect 8343 9009 8377 9043
rect 8343 8941 8377 8975
rect 8343 8873 8377 8907
rect 137 8743 171 8777
rect 205 8743 239 8777
rect 273 8743 307 8777
rect 341 8743 375 8777
rect 409 8743 443 8777
rect 477 8743 511 8777
rect 545 8743 579 8777
rect 613 8743 647 8777
rect 681 8743 715 8777
rect 749 8743 783 8777
rect 817 8743 851 8777
rect 885 8743 919 8777
rect 953 8743 987 8777
rect 1021 8743 1055 8777
rect 1089 8743 1123 8777
rect 1157 8743 1191 8777
rect 1225 8743 1259 8777
rect 1293 8743 1327 8777
rect 1361 8743 1395 8777
rect 1429 8743 1463 8777
rect 1497 8743 1531 8777
rect 1565 8743 1599 8777
rect 1633 8743 1667 8777
rect 1701 8743 1735 8777
rect 1769 8743 1803 8777
rect 1837 8743 1871 8777
rect 1905 8743 1939 8777
rect 1973 8743 2007 8777
rect 2041 8743 2075 8777
rect 2109 8743 2143 8777
rect 2177 8743 2211 8777
rect 2245 8743 2279 8777
rect 2313 8743 2347 8777
rect 2381 8743 2415 8777
rect 2449 8743 2483 8777
rect 2517 8743 2551 8777
rect 2585 8743 2619 8777
rect 2653 8743 2687 8777
rect 2721 8743 2755 8777
rect 2789 8743 2823 8777
rect 2857 8743 2891 8777
rect 2925 8743 2959 8777
rect 2993 8743 3027 8777
rect 3061 8743 3095 8777
rect 3129 8743 3163 8777
rect 3197 8743 3231 8777
rect 3265 8743 3299 8777
rect 3333 8743 3367 8777
rect 3401 8743 3435 8777
rect 3469 8743 3503 8777
rect 3537 8743 3571 8777
rect 3605 8743 3639 8777
rect 3673 8743 3707 8777
rect 3741 8743 3775 8777
rect 3809 8743 3843 8777
rect 3877 8743 3911 8777
rect 3945 8743 3979 8777
rect 4013 8743 4047 8777
rect 4081 8743 4115 8777
rect 4149 8743 4183 8777
rect 4217 8743 4251 8777
rect 4285 8743 4319 8777
rect 4353 8743 4387 8777
rect 4421 8743 4455 8777
rect 4489 8743 4523 8777
rect 4557 8743 4591 8777
rect 4625 8743 4659 8777
rect 4693 8743 4727 8777
rect 4761 8743 4795 8777
rect 4829 8743 4863 8777
rect 4897 8743 4931 8777
rect 4965 8743 4999 8777
rect 5033 8743 5067 8777
rect 5101 8743 5135 8777
rect 5169 8743 5203 8777
rect 5237 8743 5271 8777
rect 5305 8743 5339 8777
rect 5373 8743 5407 8777
rect 5441 8743 5475 8777
rect 5509 8743 5543 8777
rect 5577 8743 5611 8777
rect 5645 8743 5679 8777
rect 5713 8743 5747 8777
rect 5781 8743 5815 8777
rect 5849 8743 5883 8777
rect 5917 8743 5951 8777
rect 5985 8743 6019 8777
rect 6053 8743 6087 8777
rect 6121 8743 6155 8777
rect 6189 8743 6223 8777
rect 6257 8743 6291 8777
rect 6325 8743 6359 8777
rect 6393 8743 6427 8777
rect 6461 8743 6495 8777
rect 6529 8743 6563 8777
rect 6597 8743 6631 8777
rect 6665 8743 6699 8777
rect 6733 8743 6767 8777
rect 6801 8743 6835 8777
rect 6869 8743 6903 8777
rect 6937 8743 6971 8777
rect 7005 8743 7039 8777
rect 7073 8743 7107 8777
rect 7141 8743 7175 8777
rect 7209 8743 7243 8777
rect 7277 8743 7311 8777
rect 7345 8743 7379 8777
rect 7413 8743 7447 8777
rect 7481 8743 7515 8777
rect 7549 8743 7583 8777
rect 7617 8743 7651 8777
rect 7685 8743 7719 8777
rect 7753 8743 7787 8777
rect 7821 8743 7855 8777
rect 7889 8743 7923 8777
rect 7957 8743 7991 8777
rect 8025 8743 8059 8777
rect 8093 8743 8127 8777
rect 8161 8743 8195 8777
rect 8229 8743 8263 8777
rect 137 7943 171 7977
rect 205 7943 239 7977
rect 273 7943 307 7977
rect 341 7943 375 7977
rect 409 7943 443 7977
rect 477 7943 511 7977
rect 545 7943 579 7977
rect 613 7943 647 7977
rect 681 7943 715 7977
rect 749 7943 783 7977
rect 817 7943 851 7977
rect 885 7943 919 7977
rect 953 7943 987 7977
rect 1021 7943 1055 7977
rect 1089 7943 1123 7977
rect 1157 7943 1191 7977
rect 1225 7943 1259 7977
rect 1293 7943 1327 7977
rect 1361 7943 1395 7977
rect 1429 7943 1463 7977
rect 1497 7943 1531 7977
rect 1565 7943 1599 7977
rect 1633 7943 1667 7977
rect 1701 7943 1735 7977
rect 1769 7943 1803 7977
rect 1837 7943 1871 7977
rect 1905 7943 1939 7977
rect 1973 7943 2007 7977
rect 2041 7943 2075 7977
rect 2109 7943 2143 7977
rect 2177 7943 2211 7977
rect 2245 7943 2279 7977
rect 2313 7943 2347 7977
rect 2381 7943 2415 7977
rect 2449 7943 2483 7977
rect 2517 7943 2551 7977
rect 2585 7943 2619 7977
rect 2653 7943 2687 7977
rect 2721 7943 2755 7977
rect 2789 7943 2823 7977
rect 2857 7943 2891 7977
rect 2925 7943 2959 7977
rect 2993 7943 3027 7977
rect 3061 7943 3095 7977
rect 3129 7943 3163 7977
rect 3197 7943 3231 7977
rect 3265 7943 3299 7977
rect 3333 7943 3367 7977
rect 3401 7943 3435 7977
rect 3469 7943 3503 7977
rect 3537 7943 3571 7977
rect 3605 7943 3639 7977
rect 3673 7943 3707 7977
rect 3741 7943 3775 7977
rect 3809 7943 3843 7977
rect 3877 7943 3911 7977
rect 3945 7943 3979 7977
rect 4013 7943 4047 7977
rect 4081 7943 4115 7977
rect 4149 7943 4183 7977
rect 4217 7943 4251 7977
rect 4285 7943 4319 7977
rect 4353 7943 4387 7977
rect 4421 7943 4455 7977
rect 4489 7943 4523 7977
rect 4557 7943 4591 7977
rect 4625 7943 4659 7977
rect 4693 7943 4727 7977
rect 4761 7943 4795 7977
rect 4829 7943 4863 7977
rect 4897 7943 4931 7977
rect 4965 7943 4999 7977
rect 5033 7943 5067 7977
rect 5101 7943 5135 7977
rect 5169 7943 5203 7977
rect 5237 7943 5271 7977
rect 5305 7943 5339 7977
rect 5373 7943 5407 7977
rect 5441 7943 5475 7977
rect 5509 7943 5543 7977
rect 5577 7943 5611 7977
rect 5645 7943 5679 7977
rect 5713 7943 5747 7977
rect 5781 7943 5815 7977
rect 5849 7943 5883 7977
rect 5917 7943 5951 7977
rect 5985 7943 6019 7977
rect 6053 7943 6087 7977
rect 6121 7943 6155 7977
rect 6189 7943 6223 7977
rect 6257 7943 6291 7977
rect 6325 7943 6359 7977
rect 6393 7943 6427 7977
rect 6461 7943 6495 7977
rect 6529 7943 6563 7977
rect 6597 7943 6631 7977
rect 6665 7943 6699 7977
rect 6733 7943 6767 7977
rect 6801 7943 6835 7977
rect 6869 7943 6903 7977
rect 6937 7943 6971 7977
rect 7005 7943 7039 7977
rect 7073 7943 7107 7977
rect 7141 7943 7175 7977
rect 7209 7943 7243 7977
rect 7277 7943 7311 7977
rect 7345 7943 7379 7977
rect 7413 7943 7447 7977
rect 7481 7943 7515 7977
rect 7549 7943 7583 7977
rect 7617 7943 7651 7977
rect 7685 7943 7719 7977
rect 7753 7943 7787 7977
rect 7821 7943 7855 7977
rect 7889 7943 7923 7977
rect 7957 7943 7991 7977
rect 8025 7943 8059 7977
rect 8093 7943 8127 7977
rect 8161 7943 8195 7977
rect 8229 7943 8263 7977
rect 23 7833 57 7867
rect 23 7765 57 7799
rect 23 7697 57 7731
rect 23 7629 57 7663
rect 23 7561 57 7595
rect 23 7493 57 7527
rect 137 7383 171 7417
rect 205 7383 239 7417
rect 273 7383 307 7417
rect 341 7383 375 7417
rect 409 7383 443 7417
rect 477 7383 511 7417
rect 545 7383 579 7417
rect 613 7383 647 7417
rect 681 7383 715 7417
rect 749 7383 783 7417
rect 817 7383 851 7417
rect 885 7383 919 7417
rect 953 7383 987 7417
rect 1021 7383 1055 7417
rect 1089 7383 1123 7417
rect 1157 7383 1191 7417
rect 1225 7383 1259 7417
rect 1293 7383 1327 7417
rect 1361 7383 1395 7417
rect 1429 7383 1463 7417
rect 1497 7383 1531 7417
rect 1565 7383 1599 7417
rect 1633 7383 1667 7417
rect 1701 7383 1735 7417
rect 1769 7383 1803 7417
rect 1837 7383 1871 7417
rect 1905 7383 1939 7417
rect 1973 7383 2007 7417
rect 2041 7383 2075 7417
rect 2109 7383 2143 7417
rect 2177 7383 2211 7417
rect 2245 7383 2279 7417
rect 2313 7383 2347 7417
rect 2381 7383 2415 7417
rect 2449 7383 2483 7417
rect 2517 7383 2551 7417
rect 2585 7383 2619 7417
rect 2653 7383 2687 7417
rect 2721 7383 2755 7417
rect 2789 7383 2823 7417
rect 2857 7383 2891 7417
rect 2925 7383 2959 7417
rect 2993 7383 3027 7417
rect 3061 7383 3095 7417
rect 3129 7383 3163 7417
rect 3197 7383 3231 7417
rect 3265 7383 3299 7417
rect 3333 7383 3367 7417
rect 3401 7383 3435 7417
rect 3469 7383 3503 7417
rect 3537 7383 3571 7417
rect 3605 7383 3639 7417
rect 3673 7383 3707 7417
rect 3741 7383 3775 7417
rect 3809 7383 3843 7417
rect 3877 7383 3911 7417
rect 3945 7383 3979 7417
rect 4013 7383 4047 7417
rect 4081 7383 4115 7417
rect 4149 7383 4183 7417
rect 4217 7383 4251 7417
rect 4285 7383 4319 7417
rect 4353 7383 4387 7417
rect 4421 7383 4455 7417
rect 4489 7383 4523 7417
rect 4557 7383 4591 7417
rect 4625 7383 4659 7417
rect 4693 7383 4727 7417
rect 4761 7383 4795 7417
rect 4829 7383 4863 7417
rect 4897 7383 4931 7417
rect 4965 7383 4999 7417
rect 5033 7383 5067 7417
rect 5101 7383 5135 7417
rect 5169 7383 5203 7417
rect 5237 7383 5271 7417
rect 5305 7383 5339 7417
rect 5373 7383 5407 7417
rect 5441 7383 5475 7417
rect 5509 7383 5543 7417
rect 5577 7383 5611 7417
rect 5645 7383 5679 7417
rect 5713 7383 5747 7417
rect 5781 7383 5815 7417
rect 5849 7383 5883 7417
rect 5917 7383 5951 7417
rect 5985 7383 6019 7417
rect 6053 7383 6087 7417
rect 6121 7383 6155 7417
rect 6189 7383 6223 7417
rect 6257 7383 6291 7417
rect 6325 7383 6359 7417
rect 6393 7383 6427 7417
rect 6461 7383 6495 7417
rect 6529 7383 6563 7417
rect 6597 7383 6631 7417
rect 6665 7383 6699 7417
rect 6733 7383 6767 7417
rect 6801 7383 6835 7417
rect 6869 7383 6903 7417
rect 6937 7383 6971 7417
rect 7005 7383 7039 7417
rect 7073 7383 7107 7417
rect 7141 7383 7175 7417
rect 7209 7383 7243 7417
rect 7277 7383 7311 7417
rect 7345 7383 7379 7417
rect 7413 7383 7447 7417
rect 7481 7383 7515 7417
rect 7549 7383 7583 7417
rect 7617 7383 7651 7417
rect 7685 7383 7719 7417
rect 7753 7383 7787 7417
rect 7821 7383 7855 7417
rect 7889 7383 7923 7417
rect 7957 7383 7991 7417
rect 8025 7383 8059 7417
rect 8093 7383 8127 7417
rect 8161 7383 8195 7417
rect 8229 7383 8263 7417
rect 137 7223 171 7257
rect 205 7223 239 7257
rect 273 7223 307 7257
rect 341 7223 375 7257
rect 409 7223 443 7257
rect 477 7223 511 7257
rect 545 7223 579 7257
rect 613 7223 647 7257
rect 681 7223 715 7257
rect 749 7223 783 7257
rect 817 7223 851 7257
rect 885 7223 919 7257
rect 953 7223 987 7257
rect 1021 7223 1055 7257
rect 1089 7223 1123 7257
rect 1157 7223 1191 7257
rect 1225 7223 1259 7257
rect 1293 7223 1327 7257
rect 1361 7223 1395 7257
rect 1429 7223 1463 7257
rect 1497 7223 1531 7257
rect 1565 7223 1599 7257
rect 1633 7223 1667 7257
rect 1701 7223 1735 7257
rect 1769 7223 1803 7257
rect 1837 7223 1871 7257
rect 1905 7223 1939 7257
rect 1973 7223 2007 7257
rect 2041 7223 2075 7257
rect 2109 7223 2143 7257
rect 2177 7223 2211 7257
rect 2245 7223 2279 7257
rect 2313 7223 2347 7257
rect 2381 7223 2415 7257
rect 2449 7223 2483 7257
rect 2517 7223 2551 7257
rect 2585 7223 2619 7257
rect 2653 7223 2687 7257
rect 2721 7223 2755 7257
rect 2789 7223 2823 7257
rect 2857 7223 2891 7257
rect 2925 7223 2959 7257
rect 2993 7223 3027 7257
rect 3061 7223 3095 7257
rect 3129 7223 3163 7257
rect 3197 7223 3231 7257
rect 3265 7223 3299 7257
rect 3333 7223 3367 7257
rect 3401 7223 3435 7257
rect 3469 7223 3503 7257
rect 3537 7223 3571 7257
rect 3605 7223 3639 7257
rect 3673 7223 3707 7257
rect 3741 7223 3775 7257
rect 3809 7223 3843 7257
rect 3877 7223 3911 7257
rect 3945 7223 3979 7257
rect 4013 7223 4047 7257
rect 4081 7223 4115 7257
rect 4149 7223 4183 7257
rect 4217 7223 4251 7257
rect 4285 7223 4319 7257
rect 4353 7223 4387 7257
rect 4421 7223 4455 7257
rect 4489 7223 4523 7257
rect 4557 7223 4591 7257
rect 4625 7223 4659 7257
rect 4693 7223 4727 7257
rect 4761 7223 4795 7257
rect 4829 7223 4863 7257
rect 4897 7223 4931 7257
rect 4965 7223 4999 7257
rect 5033 7223 5067 7257
rect 5101 7223 5135 7257
rect 5169 7223 5203 7257
rect 5237 7223 5271 7257
rect 5305 7223 5339 7257
rect 5373 7223 5407 7257
rect 5441 7223 5475 7257
rect 5509 7223 5543 7257
rect 5577 7223 5611 7257
rect 5645 7223 5679 7257
rect 5713 7223 5747 7257
rect 5781 7223 5815 7257
rect 5849 7223 5883 7257
rect 5917 7223 5951 7257
rect 5985 7223 6019 7257
rect 6053 7223 6087 7257
rect 6121 7223 6155 7257
rect 6189 7223 6223 7257
rect 6257 7223 6291 7257
rect 6325 7223 6359 7257
rect 6393 7223 6427 7257
rect 6461 7223 6495 7257
rect 6529 7223 6563 7257
rect 6597 7223 6631 7257
rect 6665 7223 6699 7257
rect 6733 7223 6767 7257
rect 6801 7223 6835 7257
rect 6869 7223 6903 7257
rect 6937 7223 6971 7257
rect 7005 7223 7039 7257
rect 7073 7223 7107 7257
rect 7141 7223 7175 7257
rect 7209 7223 7243 7257
rect 7277 7223 7311 7257
rect 7345 7223 7379 7257
rect 7413 7223 7447 7257
rect 7481 7223 7515 7257
rect 7549 7223 7583 7257
rect 7617 7223 7651 7257
rect 7685 7223 7719 7257
rect 7753 7223 7787 7257
rect 7821 7223 7855 7257
rect 7889 7223 7923 7257
rect 7957 7223 7991 7257
rect 8025 7223 8059 7257
rect 8093 7223 8127 7257
rect 8161 7223 8195 7257
rect 8229 7223 8263 7257
rect 23 7113 57 7147
rect 23 7045 57 7079
rect 23 6977 57 7011
rect 23 6909 57 6943
rect 23 6841 57 6875
rect 23 6773 57 6807
rect 137 6663 171 6697
rect 205 6663 239 6697
rect 273 6663 307 6697
rect 341 6663 375 6697
rect 409 6663 443 6697
rect 477 6663 511 6697
rect 545 6663 579 6697
rect 613 6663 647 6697
rect 681 6663 715 6697
rect 749 6663 783 6697
rect 817 6663 851 6697
rect 885 6663 919 6697
rect 953 6663 987 6697
rect 1021 6663 1055 6697
rect 1089 6663 1123 6697
rect 1157 6663 1191 6697
rect 1225 6663 1259 6697
rect 1293 6663 1327 6697
rect 1361 6663 1395 6697
rect 1429 6663 1463 6697
rect 1497 6663 1531 6697
rect 1565 6663 1599 6697
rect 1633 6663 1667 6697
rect 1701 6663 1735 6697
rect 1769 6663 1803 6697
rect 1837 6663 1871 6697
rect 1905 6663 1939 6697
rect 1973 6663 2007 6697
rect 2041 6663 2075 6697
rect 2109 6663 2143 6697
rect 2177 6663 2211 6697
rect 2245 6663 2279 6697
rect 2313 6663 2347 6697
rect 2381 6663 2415 6697
rect 2449 6663 2483 6697
rect 2517 6663 2551 6697
rect 2585 6663 2619 6697
rect 2653 6663 2687 6697
rect 2721 6663 2755 6697
rect 2789 6663 2823 6697
rect 2857 6663 2891 6697
rect 2925 6663 2959 6697
rect 2993 6663 3027 6697
rect 3061 6663 3095 6697
rect 3129 6663 3163 6697
rect 3197 6663 3231 6697
rect 3265 6663 3299 6697
rect 3333 6663 3367 6697
rect 3401 6663 3435 6697
rect 3469 6663 3503 6697
rect 3537 6663 3571 6697
rect 3605 6663 3639 6697
rect 3673 6663 3707 6697
rect 3741 6663 3775 6697
rect 3809 6663 3843 6697
rect 3877 6663 3911 6697
rect 3945 6663 3979 6697
rect 4013 6663 4047 6697
rect 4081 6663 4115 6697
rect 4149 6663 4183 6697
rect 4217 6663 4251 6697
rect 4285 6663 4319 6697
rect 4353 6663 4387 6697
rect 4421 6663 4455 6697
rect 4489 6663 4523 6697
rect 4557 6663 4591 6697
rect 4625 6663 4659 6697
rect 4693 6663 4727 6697
rect 4761 6663 4795 6697
rect 4829 6663 4863 6697
rect 4897 6663 4931 6697
rect 4965 6663 4999 6697
rect 5033 6663 5067 6697
rect 5101 6663 5135 6697
rect 5169 6663 5203 6697
rect 5237 6663 5271 6697
rect 5305 6663 5339 6697
rect 5373 6663 5407 6697
rect 5441 6663 5475 6697
rect 5509 6663 5543 6697
rect 5577 6663 5611 6697
rect 5645 6663 5679 6697
rect 5713 6663 5747 6697
rect 5781 6663 5815 6697
rect 5849 6663 5883 6697
rect 5917 6663 5951 6697
rect 5985 6663 6019 6697
rect 6053 6663 6087 6697
rect 6121 6663 6155 6697
rect 6189 6663 6223 6697
rect 6257 6663 6291 6697
rect 6325 6663 6359 6697
rect 6393 6663 6427 6697
rect 6461 6663 6495 6697
rect 6529 6663 6563 6697
rect 6597 6663 6631 6697
rect 6665 6663 6699 6697
rect 6733 6663 6767 6697
rect 6801 6663 6835 6697
rect 6869 6663 6903 6697
rect 6937 6663 6971 6697
rect 7005 6663 7039 6697
rect 7073 6663 7107 6697
rect 7141 6663 7175 6697
rect 7209 6663 7243 6697
rect 7277 6663 7311 6697
rect 7345 6663 7379 6697
rect 7413 6663 7447 6697
rect 7481 6663 7515 6697
rect 7549 6663 7583 6697
rect 7617 6663 7651 6697
rect 7685 6663 7719 6697
rect 7753 6663 7787 6697
rect 7821 6663 7855 6697
rect 7889 6663 7923 6697
rect 7957 6663 7991 6697
rect 8025 6663 8059 6697
rect 8093 6663 8127 6697
rect 8161 6663 8195 6697
rect 8229 6663 8263 6697
rect 137 5383 171 5417
rect 205 5383 239 5417
rect 273 5383 307 5417
rect 341 5383 375 5417
rect 409 5383 443 5417
rect 477 5383 511 5417
rect 545 5383 579 5417
rect 613 5383 647 5417
rect 681 5383 715 5417
rect 749 5383 783 5417
rect 817 5383 851 5417
rect 885 5383 919 5417
rect 953 5383 987 5417
rect 1021 5383 1055 5417
rect 1089 5383 1123 5417
rect 1157 5383 1191 5417
rect 1225 5383 1259 5417
rect 1293 5383 1327 5417
rect 1361 5383 1395 5417
rect 1429 5383 1463 5417
rect 1497 5383 1531 5417
rect 1565 5383 1599 5417
rect 1633 5383 1667 5417
rect 1701 5383 1735 5417
rect 1769 5383 1803 5417
rect 1837 5383 1871 5417
rect 1905 5383 1939 5417
rect 1973 5383 2007 5417
rect 2041 5383 2075 5417
rect 2109 5383 2143 5417
rect 2177 5383 2211 5417
rect 2245 5383 2279 5417
rect 2313 5383 2347 5417
rect 2381 5383 2415 5417
rect 2449 5383 2483 5417
rect 2517 5383 2551 5417
rect 2585 5383 2619 5417
rect 2653 5383 2687 5417
rect 2721 5383 2755 5417
rect 2789 5383 2823 5417
rect 2857 5383 2891 5417
rect 2925 5383 2959 5417
rect 2993 5383 3027 5417
rect 3061 5383 3095 5417
rect 3129 5383 3163 5417
rect 3197 5383 3231 5417
rect 3265 5383 3299 5417
rect 3333 5383 3367 5417
rect 3401 5383 3435 5417
rect 3469 5383 3503 5417
rect 3537 5383 3571 5417
rect 3605 5383 3639 5417
rect 3673 5383 3707 5417
rect 3741 5383 3775 5417
rect 3809 5383 3843 5417
rect 3877 5383 3911 5417
rect 3945 5383 3979 5417
rect 4013 5383 4047 5417
rect 4081 5383 4115 5417
rect 4149 5383 4183 5417
rect 4217 5383 4251 5417
rect 4285 5383 4319 5417
rect 4353 5383 4387 5417
rect 4421 5383 4455 5417
rect 4489 5383 4523 5417
rect 4557 5383 4591 5417
rect 4625 5383 4659 5417
rect 4693 5383 4727 5417
rect 4761 5383 4795 5417
rect 4829 5383 4863 5417
rect 4897 5383 4931 5417
rect 4965 5383 4999 5417
rect 5033 5383 5067 5417
rect 5101 5383 5135 5417
rect 5169 5383 5203 5417
rect 5237 5383 5271 5417
rect 5305 5383 5339 5417
rect 5373 5383 5407 5417
rect 5441 5383 5475 5417
rect 5509 5383 5543 5417
rect 5577 5383 5611 5417
rect 5645 5383 5679 5417
rect 5713 5383 5747 5417
rect 5781 5383 5815 5417
rect 5849 5383 5883 5417
rect 5917 5383 5951 5417
rect 5985 5383 6019 5417
rect 6053 5383 6087 5417
rect 6121 5383 6155 5417
rect 6189 5383 6223 5417
rect 6257 5383 6291 5417
rect 6325 5383 6359 5417
rect 6393 5383 6427 5417
rect 6461 5383 6495 5417
rect 6529 5383 6563 5417
rect 6597 5383 6631 5417
rect 6665 5383 6699 5417
rect 6733 5383 6767 5417
rect 6801 5383 6835 5417
rect 6869 5383 6903 5417
rect 6937 5383 6971 5417
rect 7005 5383 7039 5417
rect 7073 5383 7107 5417
rect 7141 5383 7175 5417
rect 7209 5383 7243 5417
rect 7277 5383 7311 5417
rect 7345 5383 7379 5417
rect 7413 5383 7447 5417
rect 7481 5383 7515 5417
rect 7549 5383 7583 5417
rect 7617 5383 7651 5417
rect 7685 5383 7719 5417
rect 7753 5383 7787 5417
rect 7821 5383 7855 5417
rect 7889 5383 7923 5417
rect 7957 5383 7991 5417
rect 8025 5383 8059 5417
rect 8093 5383 8127 5417
rect 8161 5383 8195 5417
rect 8229 5383 8263 5417
rect 23 5253 57 5287
rect 23 5185 57 5219
rect 23 5117 57 5151
rect 23 5049 57 5083
rect 23 4981 57 5015
rect 23 4913 57 4947
rect 23 4845 57 4879
rect 23 4777 57 4811
rect 23 4709 57 4743
rect 23 4641 57 4675
rect 23 4573 57 4607
rect 23 4505 57 4539
rect 23 4437 57 4471
rect 23 4369 57 4403
rect 23 4301 57 4335
rect 23 4233 57 4267
rect 8343 5253 8377 5287
rect 8343 5185 8377 5219
rect 8343 5117 8377 5151
rect 8343 5049 8377 5083
rect 8343 4981 8377 5015
rect 8343 4913 8377 4947
rect 8343 4845 8377 4879
rect 8343 4777 8377 4811
rect 8343 4709 8377 4743
rect 8343 4641 8377 4675
rect 8343 4573 8377 4607
rect 8343 4505 8377 4539
rect 8343 4437 8377 4471
rect 8343 4369 8377 4403
rect 8343 4301 8377 4335
rect 8343 4233 8377 4267
rect 137 4103 171 4137
rect 205 4103 239 4137
rect 273 4103 307 4137
rect 341 4103 375 4137
rect 409 4103 443 4137
rect 477 4103 511 4137
rect 545 4103 579 4137
rect 613 4103 647 4137
rect 681 4103 715 4137
rect 749 4103 783 4137
rect 817 4103 851 4137
rect 885 4103 919 4137
rect 953 4103 987 4137
rect 1021 4103 1055 4137
rect 1089 4103 1123 4137
rect 1157 4103 1191 4137
rect 1225 4103 1259 4137
rect 1293 4103 1327 4137
rect 1361 4103 1395 4137
rect 1429 4103 1463 4137
rect 1497 4103 1531 4137
rect 1565 4103 1599 4137
rect 1633 4103 1667 4137
rect 1701 4103 1735 4137
rect 1769 4103 1803 4137
rect 1837 4103 1871 4137
rect 1905 4103 1939 4137
rect 1973 4103 2007 4137
rect 2041 4103 2075 4137
rect 2109 4103 2143 4137
rect 2177 4103 2211 4137
rect 2245 4103 2279 4137
rect 2313 4103 2347 4137
rect 2381 4103 2415 4137
rect 2449 4103 2483 4137
rect 2517 4103 2551 4137
rect 2585 4103 2619 4137
rect 2653 4103 2687 4137
rect 2721 4103 2755 4137
rect 2789 4103 2823 4137
rect 2857 4103 2891 4137
rect 2925 4103 2959 4137
rect 2993 4103 3027 4137
rect 3061 4103 3095 4137
rect 3129 4103 3163 4137
rect 3197 4103 3231 4137
rect 3265 4103 3299 4137
rect 3333 4103 3367 4137
rect 3401 4103 3435 4137
rect 3469 4103 3503 4137
rect 3537 4103 3571 4137
rect 3605 4103 3639 4137
rect 3673 4103 3707 4137
rect 3741 4103 3775 4137
rect 3809 4103 3843 4137
rect 3877 4103 3911 4137
rect 3945 4103 3979 4137
rect 4013 4103 4047 4137
rect 4081 4103 4115 4137
rect 4149 4103 4183 4137
rect 4217 4103 4251 4137
rect 4285 4103 4319 4137
rect 4353 4103 4387 4137
rect 4421 4103 4455 4137
rect 4489 4103 4523 4137
rect 4557 4103 4591 4137
rect 4625 4103 4659 4137
rect 4693 4103 4727 4137
rect 4761 4103 4795 4137
rect 4829 4103 4863 4137
rect 4897 4103 4931 4137
rect 4965 4103 4999 4137
rect 5033 4103 5067 4137
rect 5101 4103 5135 4137
rect 5169 4103 5203 4137
rect 5237 4103 5271 4137
rect 5305 4103 5339 4137
rect 5373 4103 5407 4137
rect 5441 4103 5475 4137
rect 5509 4103 5543 4137
rect 5577 4103 5611 4137
rect 5645 4103 5679 4137
rect 5713 4103 5747 4137
rect 5781 4103 5815 4137
rect 5849 4103 5883 4137
rect 5917 4103 5951 4137
rect 5985 4103 6019 4137
rect 6053 4103 6087 4137
rect 6121 4103 6155 4137
rect 6189 4103 6223 4137
rect 6257 4103 6291 4137
rect 6325 4103 6359 4137
rect 6393 4103 6427 4137
rect 6461 4103 6495 4137
rect 6529 4103 6563 4137
rect 6597 4103 6631 4137
rect 6665 4103 6699 4137
rect 6733 4103 6767 4137
rect 6801 4103 6835 4137
rect 6869 4103 6903 4137
rect 6937 4103 6971 4137
rect 7005 4103 7039 4137
rect 7073 4103 7107 4137
rect 7141 4103 7175 4137
rect 7209 4103 7243 4137
rect 7277 4103 7311 4137
rect 7345 4103 7379 4137
rect 7413 4103 7447 4137
rect 7481 4103 7515 4137
rect 7549 4103 7583 4137
rect 7617 4103 7651 4137
rect 7685 4103 7719 4137
rect 7753 4103 7787 4137
rect 7821 4103 7855 4137
rect 7889 4103 7923 4137
rect 7957 4103 7991 4137
rect 8025 4103 8059 4137
rect 8093 4103 8127 4137
rect 8161 4103 8195 4137
rect 8229 4103 8263 4137
rect 137 3943 171 3977
rect 205 3943 239 3977
rect 273 3943 307 3977
rect 341 3943 375 3977
rect 409 3943 443 3977
rect 477 3943 511 3977
rect 545 3943 579 3977
rect 613 3943 647 3977
rect 681 3943 715 3977
rect 749 3943 783 3977
rect 817 3943 851 3977
rect 885 3943 919 3977
rect 953 3943 987 3977
rect 1021 3943 1055 3977
rect 1089 3943 1123 3977
rect 1157 3943 1191 3977
rect 1225 3943 1259 3977
rect 1293 3943 1327 3977
rect 1361 3943 1395 3977
rect 1429 3943 1463 3977
rect 1497 3943 1531 3977
rect 1565 3943 1599 3977
rect 1633 3943 1667 3977
rect 1701 3943 1735 3977
rect 1769 3943 1803 3977
rect 1837 3943 1871 3977
rect 1905 3943 1939 3977
rect 1973 3943 2007 3977
rect 2041 3943 2075 3977
rect 2109 3943 2143 3977
rect 2177 3943 2211 3977
rect 2245 3943 2279 3977
rect 2313 3943 2347 3977
rect 2381 3943 2415 3977
rect 2449 3943 2483 3977
rect 2517 3943 2551 3977
rect 2585 3943 2619 3977
rect 2653 3943 2687 3977
rect 2721 3943 2755 3977
rect 2789 3943 2823 3977
rect 2857 3943 2891 3977
rect 2925 3943 2959 3977
rect 2993 3943 3027 3977
rect 3061 3943 3095 3977
rect 3129 3943 3163 3977
rect 3197 3943 3231 3977
rect 3265 3943 3299 3977
rect 3333 3943 3367 3977
rect 3401 3943 3435 3977
rect 3469 3943 3503 3977
rect 3537 3943 3571 3977
rect 3605 3943 3639 3977
rect 3673 3943 3707 3977
rect 3741 3943 3775 3977
rect 3809 3943 3843 3977
rect 3877 3943 3911 3977
rect 3945 3943 3979 3977
rect 4013 3943 4047 3977
rect 4081 3943 4115 3977
rect 4149 3943 4183 3977
rect 4217 3943 4251 3977
rect 4285 3943 4319 3977
rect 4353 3943 4387 3977
rect 4421 3943 4455 3977
rect 4489 3943 4523 3977
rect 4557 3943 4591 3977
rect 4625 3943 4659 3977
rect 4693 3943 4727 3977
rect 4761 3943 4795 3977
rect 4829 3943 4863 3977
rect 4897 3943 4931 3977
rect 4965 3943 4999 3977
rect 5033 3943 5067 3977
rect 5101 3943 5135 3977
rect 5169 3943 5203 3977
rect 5237 3943 5271 3977
rect 5305 3943 5339 3977
rect 5373 3943 5407 3977
rect 5441 3943 5475 3977
rect 5509 3943 5543 3977
rect 5577 3943 5611 3977
rect 5645 3943 5679 3977
rect 5713 3943 5747 3977
rect 5781 3943 5815 3977
rect 5849 3943 5883 3977
rect 5917 3943 5951 3977
rect 5985 3943 6019 3977
rect 6053 3943 6087 3977
rect 6121 3943 6155 3977
rect 6189 3943 6223 3977
rect 6257 3943 6291 3977
rect 6325 3943 6359 3977
rect 6393 3943 6427 3977
rect 6461 3943 6495 3977
rect 6529 3943 6563 3977
rect 6597 3943 6631 3977
rect 6665 3943 6699 3977
rect 6733 3943 6767 3977
rect 6801 3943 6835 3977
rect 6869 3943 6903 3977
rect 6937 3943 6971 3977
rect 7005 3943 7039 3977
rect 7073 3943 7107 3977
rect 7141 3943 7175 3977
rect 7209 3943 7243 3977
rect 7277 3943 7311 3977
rect 7345 3943 7379 3977
rect 7413 3943 7447 3977
rect 7481 3943 7515 3977
rect 7549 3943 7583 3977
rect 7617 3943 7651 3977
rect 7685 3943 7719 3977
rect 7753 3943 7787 3977
rect 7821 3943 7855 3977
rect 7889 3943 7923 3977
rect 7957 3943 7991 3977
rect 8025 3943 8059 3977
rect 8093 3943 8127 3977
rect 8161 3943 8195 3977
rect 8229 3943 8263 3977
rect 23 3813 57 3847
rect 23 3745 57 3779
rect 23 3677 57 3711
rect 23 3609 57 3643
rect 23 3541 57 3575
rect 23 3473 57 3507
rect 23 3405 57 3439
rect 23 3337 57 3371
rect 23 3269 57 3303
rect 23 3201 57 3235
rect 23 3133 57 3167
rect 23 3065 57 3099
rect 23 2997 57 3031
rect 23 2929 57 2963
rect 23 2861 57 2895
rect 23 2793 57 2827
rect 8343 3813 8377 3847
rect 8343 3745 8377 3779
rect 8343 3677 8377 3711
rect 8343 3609 8377 3643
rect 8343 3541 8377 3575
rect 8343 3473 8377 3507
rect 8343 3405 8377 3439
rect 8343 3337 8377 3371
rect 8343 3269 8377 3303
rect 8343 3201 8377 3235
rect 8343 3133 8377 3167
rect 8343 3065 8377 3099
rect 8343 2997 8377 3031
rect 8343 2929 8377 2963
rect 8343 2861 8377 2895
rect 8343 2793 8377 2827
rect 151 2663 185 2697
rect 219 2663 253 2697
rect 287 2663 321 2697
rect 355 2663 389 2697
rect 423 2663 457 2697
rect 491 2663 525 2697
rect 559 2663 593 2697
rect 627 2663 661 2697
rect 695 2663 729 2697
rect 763 2663 797 2697
rect 831 2663 865 2697
rect 899 2663 933 2697
rect 967 2663 1001 2697
rect 1035 2663 1069 2697
rect 1103 2663 1137 2697
rect 1171 2663 1205 2697
rect 1239 2663 1273 2697
rect 1307 2663 1341 2697
rect 1375 2663 1409 2697
rect 1443 2663 1477 2697
rect 1511 2663 1545 2697
rect 1579 2663 1613 2697
rect 1647 2663 1681 2697
rect 1715 2663 1749 2697
rect 1783 2663 1817 2697
rect 1851 2663 1885 2697
rect 1919 2663 1953 2697
rect 1987 2663 2021 2697
rect 2055 2663 2089 2697
rect 2123 2663 2157 2697
rect 2191 2663 2225 2697
rect 2259 2663 2293 2697
rect 2327 2663 2361 2697
rect 2395 2663 2429 2697
rect 2463 2663 2497 2697
rect 2531 2663 2565 2697
rect 2599 2663 2633 2697
rect 2667 2663 2701 2697
rect 2735 2663 2769 2697
rect 2803 2663 2837 2697
rect 2871 2663 2905 2697
rect 2939 2663 2973 2697
rect 3007 2663 3041 2697
rect 3075 2663 3109 2697
rect 3143 2663 3177 2697
rect 3211 2663 3245 2697
rect 3279 2663 3313 2697
rect 3347 2663 3381 2697
rect 3415 2663 3449 2697
rect 3483 2663 3517 2697
rect 3551 2663 3585 2697
rect 3619 2663 3653 2697
rect 3687 2663 3721 2697
rect 3755 2663 3789 2697
rect 3823 2663 3857 2697
rect 3891 2663 3925 2697
rect 3959 2663 3993 2697
rect 4027 2663 4061 2697
rect 4095 2663 4129 2697
rect 4163 2663 4197 2697
rect 4231 2663 4265 2697
rect 4299 2663 4333 2697
rect 4367 2663 4401 2697
rect 4435 2663 4469 2697
rect 4503 2663 4537 2697
rect 4571 2663 4605 2697
rect 4639 2663 4673 2697
rect 4707 2663 4741 2697
rect 4775 2663 4809 2697
rect 4843 2663 4877 2697
rect 4911 2663 4945 2697
rect 4979 2663 5013 2697
rect 5047 2663 5081 2697
rect 5115 2663 5149 2697
rect 5183 2663 5217 2697
rect 5251 2663 5285 2697
rect 5319 2663 5353 2697
rect 5387 2663 5421 2697
rect 5455 2663 5489 2697
rect 5523 2663 5557 2697
rect 5591 2663 5625 2697
rect 5659 2663 5693 2697
rect 5727 2663 5761 2697
rect 5795 2663 5829 2697
rect 5863 2663 5897 2697
rect 5931 2663 5965 2697
rect 5999 2663 6033 2697
rect 6067 2663 6101 2697
rect 6135 2663 6169 2697
rect 6203 2663 6237 2697
rect 6271 2663 6305 2697
rect 6339 2663 6373 2697
rect 6407 2663 6441 2697
rect 6475 2663 6509 2697
rect 6543 2663 6577 2697
rect 6611 2663 6645 2697
rect 6679 2663 6713 2697
rect 6747 2663 6781 2697
rect 6815 2663 6849 2697
rect 6883 2663 6917 2697
rect 6951 2663 6985 2697
rect 7019 2663 7053 2697
rect 7087 2663 7121 2697
rect 7155 2663 7189 2697
rect 7223 2663 7257 2697
rect 7291 2663 7325 2697
rect 7359 2663 7393 2697
rect 7427 2663 7461 2697
rect 7495 2663 7529 2697
rect 7563 2663 7597 2697
rect 7631 2663 7665 2697
rect 7699 2663 7733 2697
rect 7767 2663 7801 2697
rect 7835 2663 7869 2697
rect 7903 2663 7937 2697
rect 7971 2663 8005 2697
rect 8039 2663 8073 2697
rect 8107 2663 8141 2697
rect 8175 2663 8209 2697
rect 151 2503 185 2537
rect 219 2503 253 2537
rect 287 2503 321 2537
rect 355 2503 389 2537
rect 423 2503 457 2537
rect 491 2503 525 2537
rect 559 2503 593 2537
rect 627 2503 661 2537
rect 695 2503 729 2537
rect 763 2503 797 2537
rect 831 2503 865 2537
rect 899 2503 933 2537
rect 967 2503 1001 2537
rect 1035 2503 1069 2537
rect 1103 2503 1137 2537
rect 1171 2503 1205 2537
rect 1239 2503 1273 2537
rect 1307 2503 1341 2537
rect 1375 2503 1409 2537
rect 1443 2503 1477 2537
rect 1511 2503 1545 2537
rect 1579 2503 1613 2537
rect 1647 2503 1681 2537
rect 1715 2503 1749 2537
rect 1783 2503 1817 2537
rect 1851 2503 1885 2537
rect 1919 2503 1953 2537
rect 1987 2503 2021 2537
rect 2055 2503 2089 2537
rect 2123 2503 2157 2537
rect 2191 2503 2225 2537
rect 2259 2503 2293 2537
rect 2327 2503 2361 2537
rect 2395 2503 2429 2537
rect 2463 2503 2497 2537
rect 2531 2503 2565 2537
rect 2599 2503 2633 2537
rect 2667 2503 2701 2537
rect 2735 2503 2769 2537
rect 2803 2503 2837 2537
rect 2871 2503 2905 2537
rect 2939 2503 2973 2537
rect 3007 2503 3041 2537
rect 3075 2503 3109 2537
rect 3143 2503 3177 2537
rect 3211 2503 3245 2537
rect 3279 2503 3313 2537
rect 3347 2503 3381 2537
rect 3415 2503 3449 2537
rect 3483 2503 3517 2537
rect 3551 2503 3585 2537
rect 3619 2503 3653 2537
rect 3687 2503 3721 2537
rect 3755 2503 3789 2537
rect 3823 2503 3857 2537
rect 3891 2503 3925 2537
rect 3959 2503 3993 2537
rect 4027 2503 4061 2537
rect 4095 2503 4129 2537
rect 4163 2503 4197 2537
rect 4231 2503 4265 2537
rect 4299 2503 4333 2537
rect 4367 2503 4401 2537
rect 4435 2503 4469 2537
rect 4503 2503 4537 2537
rect 4571 2503 4605 2537
rect 4639 2503 4673 2537
rect 4707 2503 4741 2537
rect 4775 2503 4809 2537
rect 4843 2503 4877 2537
rect 4911 2503 4945 2537
rect 4979 2503 5013 2537
rect 5047 2503 5081 2537
rect 5115 2503 5149 2537
rect 5183 2503 5217 2537
rect 5251 2503 5285 2537
rect 5319 2503 5353 2537
rect 5387 2503 5421 2537
rect 5455 2503 5489 2537
rect 5523 2503 5557 2537
rect 5591 2503 5625 2537
rect 5659 2503 5693 2537
rect 5727 2503 5761 2537
rect 5795 2503 5829 2537
rect 5863 2503 5897 2537
rect 5931 2503 5965 2537
rect 5999 2503 6033 2537
rect 6067 2503 6101 2537
rect 6135 2503 6169 2537
rect 6203 2503 6237 2537
rect 6271 2503 6305 2537
rect 6339 2503 6373 2537
rect 6407 2503 6441 2537
rect 6475 2503 6509 2537
rect 6543 2503 6577 2537
rect 6611 2503 6645 2537
rect 6679 2503 6713 2537
rect 6747 2503 6781 2537
rect 6815 2503 6849 2537
rect 6883 2503 6917 2537
rect 6951 2503 6985 2537
rect 7019 2503 7053 2537
rect 7087 2503 7121 2537
rect 7155 2503 7189 2537
rect 7223 2503 7257 2537
rect 7291 2503 7325 2537
rect 7359 2503 7393 2537
rect 7427 2503 7461 2537
rect 7495 2503 7529 2537
rect 7563 2503 7597 2537
rect 7631 2503 7665 2537
rect 7699 2503 7733 2537
rect 7767 2503 7801 2537
rect 7835 2503 7869 2537
rect 7903 2503 7937 2537
rect 7971 2503 8005 2537
rect 8039 2503 8073 2537
rect 8107 2503 8141 2537
rect 8175 2503 8209 2537
rect 23 2373 57 2407
rect 23 2305 57 2339
rect 23 2237 57 2271
rect 23 2169 57 2203
rect 23 2101 57 2135
rect 23 2033 57 2067
rect 23 1965 57 1999
rect 23 1897 57 1931
rect 23 1829 57 1863
rect 23 1761 57 1795
rect 23 1693 57 1727
rect 23 1625 57 1659
rect 23 1557 57 1591
rect 23 1489 57 1523
rect 23 1421 57 1455
rect 23 1353 57 1387
rect 8343 2385 8377 2419
rect 8343 2317 8377 2351
rect 8343 2249 8377 2283
rect 8343 2181 8377 2215
rect 8343 2113 8377 2147
rect 8343 2045 8377 2079
rect 8343 1977 8377 2011
rect 8343 1909 8377 1943
rect 8343 1841 8377 1875
rect 8343 1773 8377 1807
rect 8343 1705 8377 1739
rect 8343 1637 8377 1671
rect 8343 1569 8377 1603
rect 8343 1501 8377 1535
rect 8343 1433 8377 1467
rect 8343 1365 8377 1399
rect 8343 1297 8377 1331
rect 137 1223 171 1257
rect 205 1223 239 1257
rect 273 1223 307 1257
rect 341 1223 375 1257
rect 409 1223 443 1257
rect 477 1223 511 1257
rect 545 1223 579 1257
rect 613 1223 647 1257
rect 681 1223 715 1257
rect 749 1223 783 1257
rect 817 1223 851 1257
rect 885 1223 919 1257
rect 953 1223 987 1257
rect 1021 1223 1055 1257
rect 1089 1223 1123 1257
rect 1157 1223 1191 1257
rect 1225 1223 1259 1257
rect 1293 1223 1327 1257
rect 1361 1223 1395 1257
rect 1429 1223 1463 1257
rect 1497 1223 1531 1257
rect 1565 1223 1599 1257
rect 1633 1223 1667 1257
rect 1701 1223 1735 1257
rect 1769 1223 1803 1257
rect 1837 1223 1871 1257
rect 1905 1223 1939 1257
rect 1973 1223 2007 1257
rect 2041 1223 2075 1257
rect 2109 1223 2143 1257
rect 2177 1223 2211 1257
rect 2245 1223 2279 1257
rect 2313 1223 2347 1257
rect 2381 1223 2415 1257
rect 2449 1223 2483 1257
rect 2517 1223 2551 1257
rect 2585 1223 2619 1257
rect 2653 1223 2687 1257
rect 2721 1223 2755 1257
rect 2789 1223 2823 1257
rect 2857 1223 2891 1257
rect 2925 1223 2959 1257
rect 2993 1223 3027 1257
rect 3061 1223 3095 1257
rect 3129 1223 3163 1257
rect 3197 1223 3231 1257
rect 3265 1223 3299 1257
rect 3333 1223 3367 1257
rect 3401 1223 3435 1257
rect 3469 1223 3503 1257
rect 3537 1223 3571 1257
rect 3605 1223 3639 1257
rect 3673 1223 3707 1257
rect 3741 1223 3775 1257
rect 3809 1223 3843 1257
rect 3877 1223 3911 1257
rect 3945 1223 3979 1257
rect 4013 1223 4047 1257
rect 4081 1223 4115 1257
rect 4149 1223 4183 1257
rect 4217 1223 4251 1257
rect 4285 1223 4319 1257
rect 4353 1223 4387 1257
rect 4421 1223 4455 1257
rect 4489 1223 4523 1257
rect 4557 1223 4591 1257
rect 4625 1223 4659 1257
rect 4693 1223 4727 1257
rect 4761 1223 4795 1257
rect 4829 1223 4863 1257
rect 4897 1223 4931 1257
rect 4965 1223 4999 1257
rect 5033 1223 5067 1257
rect 5101 1223 5135 1257
rect 5169 1223 5203 1257
rect 5237 1223 5271 1257
rect 5305 1223 5339 1257
rect 5373 1223 5407 1257
rect 5441 1223 5475 1257
rect 5509 1223 5543 1257
rect 5577 1223 5611 1257
rect 5645 1223 5679 1257
rect 5713 1223 5747 1257
rect 5781 1223 5815 1257
rect 5849 1223 5883 1257
rect 5917 1223 5951 1257
rect 5985 1223 6019 1257
rect 6053 1223 6087 1257
rect 6121 1223 6155 1257
rect 6189 1223 6223 1257
rect 6257 1223 6291 1257
rect 6325 1223 6359 1257
rect 6393 1223 6427 1257
rect 6461 1223 6495 1257
rect 6529 1223 6563 1257
rect 6597 1223 6631 1257
rect 6665 1223 6699 1257
rect 6733 1223 6767 1257
rect 6801 1223 6835 1257
rect 6869 1223 6903 1257
rect 6937 1223 6971 1257
rect 7005 1223 7039 1257
rect 7073 1223 7107 1257
rect 7141 1223 7175 1257
rect 7209 1223 7243 1257
rect 7277 1223 7311 1257
rect 7345 1223 7379 1257
rect 7413 1223 7447 1257
rect 7481 1223 7515 1257
rect 7549 1223 7583 1257
rect 7617 1223 7651 1257
rect 7685 1223 7719 1257
rect 7753 1223 7787 1257
rect 7821 1223 7855 1257
rect 7889 1223 7923 1257
rect 7957 1223 7991 1257
rect 8025 1223 8059 1257
rect 8093 1223 8127 1257
rect 8161 1223 8195 1257
rect 8229 1223 8263 1257
rect 8343 1229 8377 1263
rect 8343 1161 8377 1195
rect 8343 1093 8377 1127
rect 8343 1025 8377 1059
rect 8343 957 8377 991
rect 8343 889 8377 923
rect 8343 821 8377 855
rect 8343 753 8377 787
rect 8343 685 8377 719
rect 8343 617 8377 651
rect 137 583 171 617
rect 205 583 239 617
rect 273 583 307 617
rect 341 583 375 617
rect 409 583 443 617
rect 477 583 511 617
rect 545 583 579 617
rect 613 583 647 617
rect 681 583 715 617
rect 749 583 783 617
rect 817 583 851 617
rect 885 583 919 617
rect 953 583 987 617
rect 1021 583 1055 617
rect 1089 583 1123 617
rect 1157 583 1191 617
rect 1225 583 1259 617
rect 1293 583 1327 617
rect 1361 583 1395 617
rect 1429 583 1463 617
rect 1497 583 1531 617
rect 1565 583 1599 617
rect 1633 583 1667 617
rect 1701 583 1735 617
rect 1769 583 1803 617
rect 1837 583 1871 617
rect 1905 583 1939 617
rect 1973 583 2007 617
rect 2041 583 2075 617
rect 2109 583 2143 617
rect 2177 583 2211 617
rect 2245 583 2279 617
rect 2313 583 2347 617
rect 2381 583 2415 617
rect 2449 583 2483 617
rect 2517 583 2551 617
rect 2585 583 2619 617
rect 2653 583 2687 617
rect 2721 583 2755 617
rect 2789 583 2823 617
rect 2857 583 2891 617
rect 2925 583 2959 617
rect 2993 583 3027 617
rect 3061 583 3095 617
rect 3129 583 3163 617
rect 3197 583 3231 617
rect 3265 583 3299 617
rect 3333 583 3367 617
rect 3401 583 3435 617
rect 3469 583 3503 617
rect 3537 583 3571 617
rect 3605 583 3639 617
rect 3673 583 3707 617
rect 3741 583 3775 617
rect 3809 583 3843 617
rect 3877 583 3911 617
rect 3945 583 3979 617
rect 4013 583 4047 617
rect 4081 583 4115 617
rect 4149 583 4183 617
rect 4217 583 4251 617
rect 4285 583 4319 617
rect 4353 583 4387 617
rect 4421 583 4455 617
rect 4489 583 4523 617
rect 4557 583 4591 617
rect 4625 583 4659 617
rect 4693 583 4727 617
rect 4761 583 4795 617
rect 4829 583 4863 617
rect 4897 583 4931 617
rect 4965 583 4999 617
rect 5033 583 5067 617
rect 5101 583 5135 617
rect 5169 583 5203 617
rect 5237 583 5271 617
rect 5305 583 5339 617
rect 5373 583 5407 617
rect 5441 583 5475 617
rect 5509 583 5543 617
rect 5577 583 5611 617
rect 5645 583 5679 617
rect 5713 583 5747 617
rect 5781 583 5815 617
rect 5849 583 5883 617
rect 5917 583 5951 617
rect 5985 583 6019 617
rect 6053 583 6087 617
rect 6121 583 6155 617
rect 6189 583 6223 617
rect 6257 583 6291 617
rect 6325 583 6359 617
rect 6393 583 6427 617
rect 6461 583 6495 617
rect 6529 583 6563 617
rect 6597 583 6631 617
rect 6665 583 6699 617
rect 6733 583 6767 617
rect 6801 583 6835 617
rect 6869 583 6903 617
rect 6937 583 6971 617
rect 7005 583 7039 617
rect 7073 583 7107 617
rect 7141 583 7175 617
rect 7209 583 7243 617
rect 7277 583 7311 617
rect 7345 583 7379 617
rect 7413 583 7447 617
rect 7481 583 7515 617
rect 7549 583 7583 617
rect 7617 583 7651 617
rect 7685 583 7719 617
rect 7753 583 7787 617
rect 7821 583 7855 617
rect 7889 583 7923 617
rect 7957 583 7991 617
rect 8025 583 8059 617
rect 8093 583 8127 617
rect 8161 583 8195 617
rect 8229 583 8263 617
rect 23 473 57 507
rect 8343 549 8377 583
rect 8343 481 8377 515
rect 23 405 57 439
rect 23 337 57 371
rect 8343 413 8377 447
rect 23 269 57 303
rect 23 201 57 235
rect 23 133 57 167
rect 8343 345 8377 379
rect 8343 277 8377 311
rect 8343 209 8377 243
rect 8343 141 8377 175
rect 137 23 171 57
rect 205 23 239 57
rect 273 23 307 57
rect 341 23 375 57
rect 409 23 443 57
rect 477 23 511 57
rect 545 23 579 57
rect 613 23 647 57
rect 681 23 715 57
rect 749 23 783 57
rect 817 23 851 57
rect 885 23 919 57
rect 953 23 987 57
rect 1021 23 1055 57
rect 1089 23 1123 57
rect 1157 23 1191 57
rect 1225 23 1259 57
rect 1293 23 1327 57
rect 1361 23 1395 57
rect 1429 23 1463 57
rect 1497 23 1531 57
rect 1565 23 1599 57
rect 1633 23 1667 57
rect 1701 23 1735 57
rect 1769 23 1803 57
rect 1837 23 1871 57
rect 1905 23 1939 57
rect 1973 23 2007 57
rect 2041 23 2075 57
rect 2109 23 2143 57
rect 2177 23 2211 57
rect 2245 23 2279 57
rect 2313 23 2347 57
rect 2381 23 2415 57
rect 2449 23 2483 57
rect 2517 23 2551 57
rect 2585 23 2619 57
rect 2653 23 2687 57
rect 2721 23 2755 57
rect 2789 23 2823 57
rect 2857 23 2891 57
rect 2925 23 2959 57
rect 2993 23 3027 57
rect 3061 23 3095 57
rect 3129 23 3163 57
rect 3197 23 3231 57
rect 3265 23 3299 57
rect 3333 23 3367 57
rect 3401 23 3435 57
rect 3469 23 3503 57
rect 3537 23 3571 57
rect 3605 23 3639 57
rect 3673 23 3707 57
rect 3741 23 3775 57
rect 3809 23 3843 57
rect 3877 23 3911 57
rect 3945 23 3979 57
rect 4013 23 4047 57
rect 4081 23 4115 57
rect 4149 23 4183 57
rect 4217 23 4251 57
rect 4285 23 4319 57
rect 4353 23 4387 57
rect 4421 23 4455 57
rect 4489 23 4523 57
rect 4557 23 4591 57
rect 4625 23 4659 57
rect 4693 23 4727 57
rect 4761 23 4795 57
rect 4829 23 4863 57
rect 4897 23 4931 57
rect 4965 23 4999 57
rect 5033 23 5067 57
rect 5101 23 5135 57
rect 5169 23 5203 57
rect 5237 23 5271 57
rect 5305 23 5339 57
rect 5373 23 5407 57
rect 5441 23 5475 57
rect 5509 23 5543 57
rect 5577 23 5611 57
rect 5645 23 5679 57
rect 5713 23 5747 57
rect 5781 23 5815 57
rect 5849 23 5883 57
rect 5917 23 5951 57
rect 5985 23 6019 57
rect 6053 23 6087 57
rect 6121 23 6155 57
rect 6189 23 6223 57
rect 6257 23 6291 57
rect 6325 23 6359 57
rect 6393 23 6427 57
rect 6461 23 6495 57
rect 6529 23 6563 57
rect 6597 23 6631 57
rect 6665 23 6699 57
rect 6733 23 6767 57
rect 6801 23 6835 57
rect 6869 23 6903 57
rect 6937 23 6971 57
rect 7005 23 7039 57
rect 7073 23 7107 57
rect 7141 23 7175 57
rect 7209 23 7243 57
rect 7277 23 7311 57
rect 7345 23 7379 57
rect 7413 23 7447 57
rect 7481 23 7515 57
rect 7549 23 7583 57
rect 7617 23 7651 57
rect 7685 23 7719 57
rect 7753 23 7787 57
rect 7821 23 7855 57
rect 7889 23 7923 57
rect 7957 23 7991 57
rect 8025 23 8059 57
rect 8093 23 8127 57
rect 8161 23 8195 57
rect 8229 23 8263 57
rect 137 -457 171 -423
rect 205 -457 239 -423
rect 273 -457 307 -423
rect 341 -457 375 -423
rect 409 -457 443 -423
rect 477 -457 511 -423
rect 545 -457 579 -423
rect 613 -457 647 -423
rect 681 -457 715 -423
rect 749 -457 783 -423
rect 817 -457 851 -423
rect 885 -457 919 -423
rect 953 -457 987 -423
rect 1021 -457 1055 -423
rect 1089 -457 1123 -423
rect 1157 -457 1191 -423
rect 1225 -457 1259 -423
rect 1293 -457 1327 -423
rect 1361 -457 1395 -423
rect 1429 -457 1463 -423
rect 1497 -457 1531 -423
rect 1565 -457 1599 -423
rect 1633 -457 1667 -423
rect 1701 -457 1735 -423
rect 1769 -457 1803 -423
rect 1837 -457 1871 -423
rect 1905 -457 1939 -423
rect 1973 -457 2007 -423
rect 2041 -457 2075 -423
rect 2109 -457 2143 -423
rect 2177 -457 2211 -423
rect 2245 -457 2279 -423
rect 2313 -457 2347 -423
rect 2381 -457 2415 -423
rect 2449 -457 2483 -423
rect 2517 -457 2551 -423
rect 2585 -457 2619 -423
rect 2653 -457 2687 -423
rect 2721 -457 2755 -423
rect 2789 -457 2823 -423
rect 2857 -457 2891 -423
rect 2925 -457 2959 -423
rect 2993 -457 3027 -423
rect 3061 -457 3095 -423
rect 3129 -457 3163 -423
rect 3197 -457 3231 -423
rect 3265 -457 3299 -423
rect 3333 -457 3367 -423
rect 3401 -457 3435 -423
rect 3469 -457 3503 -423
rect 3537 -457 3571 -423
rect 3605 -457 3639 -423
rect 3673 -457 3707 -423
rect 3741 -457 3775 -423
rect 3809 -457 3843 -423
rect 3877 -457 3911 -423
rect 3945 -457 3979 -423
rect 4013 -457 4047 -423
rect 4081 -457 4115 -423
rect 4149 -457 4183 -423
rect 4217 -457 4251 -423
rect 4285 -457 4319 -423
rect 4353 -457 4387 -423
rect 4421 -457 4455 -423
rect 4489 -457 4523 -423
rect 4557 -457 4591 -423
rect 4625 -457 4659 -423
rect 4693 -457 4727 -423
rect 4761 -457 4795 -423
rect 4829 -457 4863 -423
rect 4897 -457 4931 -423
rect 4965 -457 4999 -423
rect 5033 -457 5067 -423
rect 5101 -457 5135 -423
rect 5169 -457 5203 -423
rect 5237 -457 5271 -423
rect 5305 -457 5339 -423
rect 5373 -457 5407 -423
rect 5441 -457 5475 -423
rect 5509 -457 5543 -423
rect 5577 -457 5611 -423
rect 5645 -457 5679 -423
rect 5713 -457 5747 -423
rect 5781 -457 5815 -423
rect 5849 -457 5883 -423
rect 5917 -457 5951 -423
rect 5985 -457 6019 -423
rect 6053 -457 6087 -423
rect 6121 -457 6155 -423
rect 6189 -457 6223 -423
rect 6257 -457 6291 -423
rect 6325 -457 6359 -423
rect 6393 -457 6427 -423
rect 6461 -457 6495 -423
rect 6529 -457 6563 -423
rect 6597 -457 6631 -423
rect 6665 -457 6699 -423
rect 6733 -457 6767 -423
rect 6801 -457 6835 -423
rect 6869 -457 6903 -423
rect 6937 -457 6971 -423
rect 7005 -457 7039 -423
rect 7073 -457 7107 -423
rect 7141 -457 7175 -423
rect 7209 -457 7243 -423
rect 7277 -457 7311 -423
rect 7345 -457 7379 -423
rect 7413 -457 7447 -423
rect 7481 -457 7515 -423
rect 7549 -457 7583 -423
rect 7617 -457 7651 -423
rect 7685 -457 7719 -423
rect 7753 -457 7787 -423
rect 7821 -457 7855 -423
rect 7889 -457 7923 -423
rect 7957 -457 7991 -423
rect 8025 -457 8059 -423
rect 8093 -457 8127 -423
rect 8161 -457 8195 -423
rect 8229 -457 8263 -423
rect 23 -567 57 -533
rect 23 -635 57 -601
rect 23 -703 57 -669
rect 8343 -567 8377 -533
rect 8343 -635 8377 -601
rect 23 -771 57 -737
rect 23 -839 57 -805
rect 23 -907 57 -873
rect 8343 -703 8377 -669
rect 8343 -771 8377 -737
rect 8343 -839 8377 -805
rect 8343 -907 8377 -873
rect 137 -1017 171 -983
rect 205 -1017 239 -983
rect 273 -1017 307 -983
rect 341 -1017 375 -983
rect 409 -1017 443 -983
rect 477 -1017 511 -983
rect 545 -1017 579 -983
rect 613 -1017 647 -983
rect 681 -1017 715 -983
rect 749 -1017 783 -983
rect 817 -1017 851 -983
rect 885 -1017 919 -983
rect 953 -1017 987 -983
rect 1021 -1017 1055 -983
rect 1089 -1017 1123 -983
rect 1157 -1017 1191 -983
rect 1225 -1017 1259 -983
rect 1293 -1017 1327 -983
rect 1361 -1017 1395 -983
rect 1429 -1017 1463 -983
rect 1497 -1017 1531 -983
rect 1565 -1017 1599 -983
rect 1633 -1017 1667 -983
rect 1701 -1017 1735 -983
rect 1769 -1017 1803 -983
rect 1837 -1017 1871 -983
rect 1905 -1017 1939 -983
rect 1973 -1017 2007 -983
rect 2041 -1017 2075 -983
rect 2109 -1017 2143 -983
rect 2177 -1017 2211 -983
rect 2245 -1017 2279 -983
rect 2313 -1017 2347 -983
rect 2381 -1017 2415 -983
rect 2449 -1017 2483 -983
rect 2517 -1017 2551 -983
rect 2585 -1017 2619 -983
rect 2653 -1017 2687 -983
rect 2721 -1017 2755 -983
rect 2789 -1017 2823 -983
rect 2857 -1017 2891 -983
rect 2925 -1017 2959 -983
rect 2993 -1017 3027 -983
rect 3061 -1017 3095 -983
rect 3129 -1017 3163 -983
rect 3197 -1017 3231 -983
rect 3265 -1017 3299 -983
rect 3333 -1017 3367 -983
rect 3401 -1017 3435 -983
rect 3469 -1017 3503 -983
rect 3537 -1017 3571 -983
rect 3605 -1017 3639 -983
rect 3673 -1017 3707 -983
rect 3741 -1017 3775 -983
rect 3809 -1017 3843 -983
rect 3877 -1017 3911 -983
rect 3945 -1017 3979 -983
rect 4013 -1017 4047 -983
rect 4081 -1017 4115 -983
rect 4149 -1017 4183 -983
rect 4217 -1017 4251 -983
rect 4285 -1017 4319 -983
rect 4353 -1017 4387 -983
rect 4421 -1017 4455 -983
rect 4489 -1017 4523 -983
rect 4557 -1017 4591 -983
rect 4625 -1017 4659 -983
rect 4693 -1017 4727 -983
rect 4761 -1017 4795 -983
rect 4829 -1017 4863 -983
rect 4897 -1017 4931 -983
rect 4965 -1017 4999 -983
rect 5033 -1017 5067 -983
rect 5101 -1017 5135 -983
rect 5169 -1017 5203 -983
rect 5237 -1017 5271 -983
rect 5305 -1017 5339 -983
rect 5373 -1017 5407 -983
rect 5441 -1017 5475 -983
rect 5509 -1017 5543 -983
rect 5577 -1017 5611 -983
rect 5645 -1017 5679 -983
rect 5713 -1017 5747 -983
rect 5781 -1017 5815 -983
rect 5849 -1017 5883 -983
rect 5917 -1017 5951 -983
rect 5985 -1017 6019 -983
rect 6053 -1017 6087 -983
rect 6121 -1017 6155 -983
rect 6189 -1017 6223 -983
rect 6257 -1017 6291 -983
rect 6325 -1017 6359 -983
rect 6393 -1017 6427 -983
rect 6461 -1017 6495 -983
rect 6529 -1017 6563 -983
rect 6597 -1017 6631 -983
rect 6665 -1017 6699 -983
rect 6733 -1017 6767 -983
rect 6801 -1017 6835 -983
rect 6869 -1017 6903 -983
rect 6937 -1017 6971 -983
rect 7005 -1017 7039 -983
rect 7073 -1017 7107 -983
rect 7141 -1017 7175 -983
rect 7209 -1017 7243 -983
rect 7277 -1017 7311 -983
rect 7345 -1017 7379 -983
rect 7413 -1017 7447 -983
rect 7481 -1017 7515 -983
rect 7549 -1017 7583 -983
rect 7617 -1017 7651 -983
rect 7685 -1017 7719 -983
rect 7753 -1017 7787 -983
rect 7821 -1017 7855 -983
rect 7889 -1017 7923 -983
rect 7957 -1017 7991 -983
rect 8025 -1017 8059 -983
rect 8093 -1017 8127 -983
rect 8161 -1017 8195 -983
rect 8229 -1017 8263 -983
<< mvnsubdiffcont >>
rect 307 9863 341 9897
rect 375 9863 409 9897
rect 443 9863 477 9897
rect 511 9863 545 9897
rect 579 9863 613 9897
rect 647 9863 681 9897
rect 715 9863 749 9897
rect 783 9863 817 9897
rect 851 9863 885 9897
rect 919 9863 953 9897
rect 987 9863 1021 9897
rect 1055 9863 1089 9897
rect 1123 9863 1157 9897
rect 1191 9863 1225 9897
rect 1259 9863 1293 9897
rect 1327 9863 1361 9897
rect 1395 9863 1429 9897
rect 1463 9863 1497 9897
rect 1531 9863 1565 9897
rect 1599 9863 1633 9897
rect 1667 9863 1701 9897
rect 1735 9863 1769 9897
rect 1803 9863 1837 9897
rect 1871 9863 1905 9897
rect 1939 9863 1973 9897
rect 2007 9863 2041 9897
rect 2075 9863 2109 9897
rect 2143 9863 2177 9897
rect 2211 9863 2245 9897
rect 2279 9863 2313 9897
rect 2347 9863 2381 9897
rect 2415 9863 2449 9897
rect 2483 9863 2517 9897
rect 2551 9863 2585 9897
rect 2619 9863 2653 9897
rect 2687 9863 2721 9897
rect 2755 9863 2789 9897
rect 2823 9863 2857 9897
rect 2891 9863 2925 9897
rect 2959 9863 2993 9897
rect 3027 9863 3061 9897
rect 3095 9863 3129 9897
rect 3163 9863 3197 9897
rect 3231 9863 3265 9897
rect 3299 9863 3333 9897
rect 3367 9863 3401 9897
rect 3435 9863 3469 9897
rect 3503 9863 3537 9897
rect 3571 9863 3605 9897
rect 3639 9863 3673 9897
rect 3707 9863 3741 9897
rect 3775 9863 3809 9897
rect 3843 9863 3877 9897
rect 3911 9863 3945 9897
rect 3979 9863 4013 9897
rect 4047 9863 4081 9897
rect 4115 9863 4149 9897
rect 4183 9863 4217 9897
rect 4251 9863 4285 9897
rect 4319 9863 4353 9897
rect 4387 9863 4421 9897
rect 4455 9863 4489 9897
rect 4523 9863 4557 9897
rect 4591 9863 4625 9897
rect 4659 9863 4693 9897
rect 4727 9863 4761 9897
rect 4795 9863 4829 9897
rect 4863 9863 4897 9897
rect 4931 9863 4965 9897
rect 4999 9863 5033 9897
rect 5067 9863 5101 9897
rect 5135 9863 5169 9897
rect 5203 9863 5237 9897
rect 5271 9863 5305 9897
rect 5339 9863 5373 9897
rect 5407 9863 5441 9897
rect 5475 9863 5509 9897
rect 5543 9863 5577 9897
rect 5611 9863 5645 9897
rect 5679 9863 5713 9897
rect 5747 9863 5781 9897
rect 5815 9863 5849 9897
rect 5883 9863 5917 9897
rect 5951 9863 5985 9897
rect 6019 9863 6053 9897
rect 6087 9863 6121 9897
rect 6155 9863 6189 9897
rect 6223 9863 6257 9897
rect 6291 9863 6325 9897
rect 6359 9863 6393 9897
rect 6427 9863 6461 9897
rect 6495 9863 6529 9897
rect 6563 9863 6597 9897
rect 6631 9863 6665 9897
rect 6699 9863 6733 9897
rect 6767 9863 6801 9897
rect 6835 9863 6869 9897
rect 6903 9863 6937 9897
rect 6971 9863 7005 9897
rect 7039 9863 7073 9897
rect 7107 9863 7141 9897
rect 7175 9863 7209 9897
rect 7243 9863 7277 9897
rect 7311 9863 7345 9897
rect 7379 9863 7413 9897
rect 7447 9863 7481 9897
rect 7515 9863 7549 9897
rect 7583 9863 7617 9897
rect 7651 9863 7685 9897
rect 7719 9863 7753 9897
rect 7787 9863 7821 9897
rect 7855 9863 7889 9897
rect 7923 9863 7957 9897
rect 7991 9863 8025 9897
rect 8059 9863 8093 9897
rect 183 9757 217 9791
rect 183 9689 217 9723
rect 183 9621 217 9655
rect 183 9553 217 9587
rect 183 9485 217 9519
rect 183 9417 217 9451
rect 183 9349 217 9383
rect 183 9281 217 9315
rect 183 9213 217 9247
rect 183 9145 217 9179
rect 8183 9757 8217 9791
rect 8183 9689 8217 9723
rect 8183 9621 8217 9655
rect 8183 9553 8217 9587
rect 8183 9485 8217 9519
rect 8183 9417 8217 9451
rect 8183 9349 8217 9383
rect 8183 9281 8217 9315
rect 8183 9213 8217 9247
rect 183 9077 217 9111
rect 183 9009 217 9043
rect 8183 9145 8217 9179
rect 8183 9077 8217 9111
rect 8183 9009 8217 9043
rect 307 8903 341 8937
rect 375 8903 409 8937
rect 443 8903 477 8937
rect 511 8903 545 8937
rect 579 8903 613 8937
rect 647 8903 681 8937
rect 715 8903 749 8937
rect 783 8903 817 8937
rect 851 8903 885 8937
rect 919 8903 953 8937
rect 987 8903 1021 8937
rect 1055 8903 1089 8937
rect 1123 8903 1157 8937
rect 1191 8903 1225 8937
rect 1259 8903 1293 8937
rect 1327 8903 1361 8937
rect 1395 8903 1429 8937
rect 1463 8903 1497 8937
rect 1531 8903 1565 8937
rect 1599 8903 1633 8937
rect 1667 8903 1701 8937
rect 1735 8903 1769 8937
rect 1803 8903 1837 8937
rect 1871 8903 1905 8937
rect 1939 8903 1973 8937
rect 2007 8903 2041 8937
rect 2075 8903 2109 8937
rect 2143 8903 2177 8937
rect 2211 8903 2245 8937
rect 2279 8903 2313 8937
rect 2347 8903 2381 8937
rect 2415 8903 2449 8937
rect 2483 8903 2517 8937
rect 2551 8903 2585 8937
rect 2619 8903 2653 8937
rect 2687 8903 2721 8937
rect 2755 8903 2789 8937
rect 2823 8903 2857 8937
rect 2891 8903 2925 8937
rect 2959 8903 2993 8937
rect 3027 8903 3061 8937
rect 3095 8903 3129 8937
rect 3163 8903 3197 8937
rect 3231 8903 3265 8937
rect 3299 8903 3333 8937
rect 3367 8903 3401 8937
rect 3435 8903 3469 8937
rect 3503 8903 3537 8937
rect 3571 8903 3605 8937
rect 3639 8903 3673 8937
rect 3707 8903 3741 8937
rect 3775 8903 3809 8937
rect 3843 8903 3877 8937
rect 3911 8903 3945 8937
rect 3979 8903 4013 8937
rect 4047 8903 4081 8937
rect 4115 8903 4149 8937
rect 4183 8903 4217 8937
rect 4251 8903 4285 8937
rect 4319 8903 4353 8937
rect 4387 8903 4421 8937
rect 4455 8903 4489 8937
rect 4523 8903 4557 8937
rect 4591 8903 4625 8937
rect 4659 8903 4693 8937
rect 4727 8903 4761 8937
rect 4795 8903 4829 8937
rect 4863 8903 4897 8937
rect 4931 8903 4965 8937
rect 4999 8903 5033 8937
rect 5067 8903 5101 8937
rect 5135 8903 5169 8937
rect 5203 8903 5237 8937
rect 5271 8903 5305 8937
rect 5339 8903 5373 8937
rect 5407 8903 5441 8937
rect 5475 8903 5509 8937
rect 5543 8903 5577 8937
rect 5611 8903 5645 8937
rect 5679 8903 5713 8937
rect 5747 8903 5781 8937
rect 5815 8903 5849 8937
rect 5883 8903 5917 8937
rect 5951 8903 5985 8937
rect 6019 8903 6053 8937
rect 6087 8903 6121 8937
rect 6155 8903 6189 8937
rect 6223 8903 6257 8937
rect 6291 8903 6325 8937
rect 6359 8903 6393 8937
rect 6427 8903 6461 8937
rect 6495 8903 6529 8937
rect 6563 8903 6597 8937
rect 6631 8903 6665 8937
rect 6699 8903 6733 8937
rect 6767 8903 6801 8937
rect 6835 8903 6869 8937
rect 6903 8903 6937 8937
rect 6971 8903 7005 8937
rect 7039 8903 7073 8937
rect 7107 8903 7141 8937
rect 7175 8903 7209 8937
rect 7243 8903 7277 8937
rect 7311 8903 7345 8937
rect 7379 8903 7413 8937
rect 7447 8903 7481 8937
rect 7515 8903 7549 8937
rect 7583 8903 7617 8937
rect 7651 8903 7685 8937
rect 7719 8903 7753 8937
rect 7787 8903 7821 8937
rect 7855 8903 7889 8937
rect 7923 8903 7957 8937
rect 7991 8903 8025 8937
rect 8059 8903 8093 8937
rect 307 5223 341 5257
rect 375 5223 409 5257
rect 443 5223 477 5257
rect 511 5223 545 5257
rect 579 5223 613 5257
rect 647 5223 681 5257
rect 715 5223 749 5257
rect 783 5223 817 5257
rect 851 5223 885 5257
rect 919 5223 953 5257
rect 987 5223 1021 5257
rect 1055 5223 1089 5257
rect 1123 5223 1157 5257
rect 1191 5223 1225 5257
rect 1259 5223 1293 5257
rect 1327 5223 1361 5257
rect 1395 5223 1429 5257
rect 1463 5223 1497 5257
rect 1531 5223 1565 5257
rect 1599 5223 1633 5257
rect 1667 5223 1701 5257
rect 1735 5223 1769 5257
rect 1803 5223 1837 5257
rect 1871 5223 1905 5257
rect 1939 5223 1973 5257
rect 2007 5223 2041 5257
rect 2075 5223 2109 5257
rect 2143 5223 2177 5257
rect 2211 5223 2245 5257
rect 2279 5223 2313 5257
rect 2347 5223 2381 5257
rect 2415 5223 2449 5257
rect 2483 5223 2517 5257
rect 2551 5223 2585 5257
rect 2619 5223 2653 5257
rect 2687 5223 2721 5257
rect 2755 5223 2789 5257
rect 2823 5223 2857 5257
rect 2891 5223 2925 5257
rect 2959 5223 2993 5257
rect 3027 5223 3061 5257
rect 3095 5223 3129 5257
rect 3163 5223 3197 5257
rect 3231 5223 3265 5257
rect 3299 5223 3333 5257
rect 3367 5223 3401 5257
rect 3435 5223 3469 5257
rect 3503 5223 3537 5257
rect 3571 5223 3605 5257
rect 3639 5223 3673 5257
rect 3707 5223 3741 5257
rect 3775 5223 3809 5257
rect 3843 5223 3877 5257
rect 3911 5223 3945 5257
rect 3979 5223 4013 5257
rect 4047 5223 4081 5257
rect 4115 5223 4149 5257
rect 4183 5223 4217 5257
rect 4251 5223 4285 5257
rect 4319 5223 4353 5257
rect 4387 5223 4421 5257
rect 4455 5223 4489 5257
rect 4523 5223 4557 5257
rect 4591 5223 4625 5257
rect 4659 5223 4693 5257
rect 4727 5223 4761 5257
rect 4795 5223 4829 5257
rect 4863 5223 4897 5257
rect 4931 5223 4965 5257
rect 4999 5223 5033 5257
rect 5067 5223 5101 5257
rect 5135 5223 5169 5257
rect 5203 5223 5237 5257
rect 5271 5223 5305 5257
rect 5339 5223 5373 5257
rect 5407 5223 5441 5257
rect 5475 5223 5509 5257
rect 5543 5223 5577 5257
rect 5611 5223 5645 5257
rect 5679 5223 5713 5257
rect 5747 5223 5781 5257
rect 5815 5223 5849 5257
rect 5883 5223 5917 5257
rect 5951 5223 5985 5257
rect 6019 5223 6053 5257
rect 6087 5223 6121 5257
rect 6155 5223 6189 5257
rect 6223 5223 6257 5257
rect 6291 5223 6325 5257
rect 6359 5223 6393 5257
rect 6427 5223 6461 5257
rect 6495 5223 6529 5257
rect 6563 5223 6597 5257
rect 6631 5223 6665 5257
rect 6699 5223 6733 5257
rect 6767 5223 6801 5257
rect 6835 5223 6869 5257
rect 6903 5223 6937 5257
rect 6971 5223 7005 5257
rect 7039 5223 7073 5257
rect 7107 5223 7141 5257
rect 7175 5223 7209 5257
rect 7243 5223 7277 5257
rect 7311 5223 7345 5257
rect 7379 5223 7413 5257
rect 7447 5223 7481 5257
rect 7515 5223 7549 5257
rect 7583 5223 7617 5257
rect 7651 5223 7685 5257
rect 7719 5223 7753 5257
rect 7787 5223 7821 5257
rect 7855 5223 7889 5257
rect 7923 5223 7957 5257
rect 7991 5223 8025 5257
rect 8059 5223 8093 5257
rect 183 5117 217 5151
rect 183 5049 217 5083
rect 183 4981 217 5015
rect 8183 5117 8217 5151
rect 8183 5049 8217 5083
rect 183 4913 217 4947
rect 183 4845 217 4879
rect 183 4777 217 4811
rect 183 4709 217 4743
rect 183 4641 217 4675
rect 183 4573 217 4607
rect 183 4505 217 4539
rect 183 4437 217 4471
rect 183 4369 217 4403
rect 8183 4981 8217 5015
rect 8183 4913 8217 4947
rect 8183 4845 8217 4879
rect 8183 4777 8217 4811
rect 8183 4709 8217 4743
rect 8183 4641 8217 4675
rect 8183 4573 8217 4607
rect 8183 4505 8217 4539
rect 8183 4437 8217 4471
rect 8183 4369 8217 4403
rect 307 4263 341 4297
rect 375 4263 409 4297
rect 443 4263 477 4297
rect 511 4263 545 4297
rect 579 4263 613 4297
rect 647 4263 681 4297
rect 715 4263 749 4297
rect 783 4263 817 4297
rect 851 4263 885 4297
rect 919 4263 953 4297
rect 987 4263 1021 4297
rect 1055 4263 1089 4297
rect 1123 4263 1157 4297
rect 1191 4263 1225 4297
rect 1259 4263 1293 4297
rect 1327 4263 1361 4297
rect 1395 4263 1429 4297
rect 1463 4263 1497 4297
rect 1531 4263 1565 4297
rect 1599 4263 1633 4297
rect 1667 4263 1701 4297
rect 1735 4263 1769 4297
rect 1803 4263 1837 4297
rect 1871 4263 1905 4297
rect 1939 4263 1973 4297
rect 2007 4263 2041 4297
rect 2075 4263 2109 4297
rect 2143 4263 2177 4297
rect 2211 4263 2245 4297
rect 2279 4263 2313 4297
rect 2347 4263 2381 4297
rect 2415 4263 2449 4297
rect 2483 4263 2517 4297
rect 2551 4263 2585 4297
rect 2619 4263 2653 4297
rect 2687 4263 2721 4297
rect 2755 4263 2789 4297
rect 2823 4263 2857 4297
rect 2891 4263 2925 4297
rect 2959 4263 2993 4297
rect 3027 4263 3061 4297
rect 3095 4263 3129 4297
rect 3163 4263 3197 4297
rect 3231 4263 3265 4297
rect 3299 4263 3333 4297
rect 3367 4263 3401 4297
rect 3435 4263 3469 4297
rect 3503 4263 3537 4297
rect 3571 4263 3605 4297
rect 3639 4263 3673 4297
rect 3707 4263 3741 4297
rect 3775 4263 3809 4297
rect 3843 4263 3877 4297
rect 3911 4263 3945 4297
rect 3979 4263 4013 4297
rect 4047 4263 4081 4297
rect 4115 4263 4149 4297
rect 4183 4263 4217 4297
rect 4251 4263 4285 4297
rect 4319 4263 4353 4297
rect 4387 4263 4421 4297
rect 4455 4263 4489 4297
rect 4523 4263 4557 4297
rect 4591 4263 4625 4297
rect 4659 4263 4693 4297
rect 4727 4263 4761 4297
rect 4795 4263 4829 4297
rect 4863 4263 4897 4297
rect 4931 4263 4965 4297
rect 4999 4263 5033 4297
rect 5067 4263 5101 4297
rect 5135 4263 5169 4297
rect 5203 4263 5237 4297
rect 5271 4263 5305 4297
rect 5339 4263 5373 4297
rect 5407 4263 5441 4297
rect 5475 4263 5509 4297
rect 5543 4263 5577 4297
rect 5611 4263 5645 4297
rect 5679 4263 5713 4297
rect 5747 4263 5781 4297
rect 5815 4263 5849 4297
rect 5883 4263 5917 4297
rect 5951 4263 5985 4297
rect 6019 4263 6053 4297
rect 6087 4263 6121 4297
rect 6155 4263 6189 4297
rect 6223 4263 6257 4297
rect 6291 4263 6325 4297
rect 6359 4263 6393 4297
rect 6427 4263 6461 4297
rect 6495 4263 6529 4297
rect 6563 4263 6597 4297
rect 6631 4263 6665 4297
rect 6699 4263 6733 4297
rect 6767 4263 6801 4297
rect 6835 4263 6869 4297
rect 6903 4263 6937 4297
rect 6971 4263 7005 4297
rect 7039 4263 7073 4297
rect 7107 4263 7141 4297
rect 7175 4263 7209 4297
rect 7243 4263 7277 4297
rect 7311 4263 7345 4297
rect 7379 4263 7413 4297
rect 7447 4263 7481 4297
rect 7515 4263 7549 4297
rect 7583 4263 7617 4297
rect 7651 4263 7685 4297
rect 7719 4263 7753 4297
rect 7787 4263 7821 4297
rect 7855 4263 7889 4297
rect 7923 4263 7957 4297
rect 7991 4263 8025 4297
rect 8059 4263 8093 4297
rect 307 3783 341 3817
rect 375 3783 409 3817
rect 443 3783 477 3817
rect 511 3783 545 3817
rect 579 3783 613 3817
rect 647 3783 681 3817
rect 715 3783 749 3817
rect 783 3783 817 3817
rect 851 3783 885 3817
rect 919 3783 953 3817
rect 987 3783 1021 3817
rect 1055 3783 1089 3817
rect 1123 3783 1157 3817
rect 1191 3783 1225 3817
rect 1259 3783 1293 3817
rect 1327 3783 1361 3817
rect 1395 3783 1429 3817
rect 1463 3783 1497 3817
rect 1531 3783 1565 3817
rect 1599 3783 1633 3817
rect 1667 3783 1701 3817
rect 1735 3783 1769 3817
rect 1803 3783 1837 3817
rect 1871 3783 1905 3817
rect 1939 3783 1973 3817
rect 2007 3783 2041 3817
rect 2075 3783 2109 3817
rect 2143 3783 2177 3817
rect 2211 3783 2245 3817
rect 2279 3783 2313 3817
rect 2347 3783 2381 3817
rect 2415 3783 2449 3817
rect 2483 3783 2517 3817
rect 2551 3783 2585 3817
rect 2619 3783 2653 3817
rect 2687 3783 2721 3817
rect 2755 3783 2789 3817
rect 2823 3783 2857 3817
rect 2891 3783 2925 3817
rect 2959 3783 2993 3817
rect 3027 3783 3061 3817
rect 3095 3783 3129 3817
rect 3163 3783 3197 3817
rect 3231 3783 3265 3817
rect 3299 3783 3333 3817
rect 3367 3783 3401 3817
rect 3435 3783 3469 3817
rect 3503 3783 3537 3817
rect 3571 3783 3605 3817
rect 3639 3783 3673 3817
rect 3707 3783 3741 3817
rect 3775 3783 3809 3817
rect 3843 3783 3877 3817
rect 3911 3783 3945 3817
rect 3979 3783 4013 3817
rect 4047 3783 4081 3817
rect 4115 3783 4149 3817
rect 4183 3783 4217 3817
rect 4251 3783 4285 3817
rect 4319 3783 4353 3817
rect 4387 3783 4421 3817
rect 4455 3783 4489 3817
rect 4523 3783 4557 3817
rect 4591 3783 4625 3817
rect 4659 3783 4693 3817
rect 4727 3783 4761 3817
rect 4795 3783 4829 3817
rect 4863 3783 4897 3817
rect 4931 3783 4965 3817
rect 4999 3783 5033 3817
rect 5067 3783 5101 3817
rect 5135 3783 5169 3817
rect 5203 3783 5237 3817
rect 5271 3783 5305 3817
rect 5339 3783 5373 3817
rect 5407 3783 5441 3817
rect 5475 3783 5509 3817
rect 5543 3783 5577 3817
rect 5611 3783 5645 3817
rect 5679 3783 5713 3817
rect 5747 3783 5781 3817
rect 5815 3783 5849 3817
rect 5883 3783 5917 3817
rect 5951 3783 5985 3817
rect 6019 3783 6053 3817
rect 6087 3783 6121 3817
rect 6155 3783 6189 3817
rect 6223 3783 6257 3817
rect 6291 3783 6325 3817
rect 6359 3783 6393 3817
rect 6427 3783 6461 3817
rect 6495 3783 6529 3817
rect 6563 3783 6597 3817
rect 6631 3783 6665 3817
rect 6699 3783 6733 3817
rect 6767 3783 6801 3817
rect 6835 3783 6869 3817
rect 6903 3783 6937 3817
rect 6971 3783 7005 3817
rect 7039 3783 7073 3817
rect 7107 3783 7141 3817
rect 7175 3783 7209 3817
rect 7243 3783 7277 3817
rect 7311 3783 7345 3817
rect 7379 3783 7413 3817
rect 7447 3783 7481 3817
rect 7515 3783 7549 3817
rect 7583 3783 7617 3817
rect 7651 3783 7685 3817
rect 7719 3783 7753 3817
rect 7787 3783 7821 3817
rect 7855 3783 7889 3817
rect 7923 3783 7957 3817
rect 7991 3783 8025 3817
rect 8059 3783 8093 3817
rect 183 3677 217 3711
rect 183 3609 217 3643
rect 183 3541 217 3575
rect 183 3473 217 3507
rect 183 3405 217 3439
rect 183 3337 217 3371
rect 183 3269 217 3303
rect 183 3201 217 3235
rect 183 3133 217 3167
rect 183 3065 217 3099
rect 8183 3677 8217 3711
rect 8183 3609 8217 3643
rect 8183 3541 8217 3575
rect 8183 3473 8217 3507
rect 8183 3405 8217 3439
rect 8183 3337 8217 3371
rect 8183 3269 8217 3303
rect 8183 3201 8217 3235
rect 8183 3133 8217 3167
rect 183 2997 217 3031
rect 183 2929 217 2963
rect 8183 3065 8217 3099
rect 8183 2997 8217 3031
rect 8183 2929 8217 2963
rect 307 2823 341 2857
rect 375 2823 409 2857
rect 443 2823 477 2857
rect 511 2823 545 2857
rect 579 2823 613 2857
rect 647 2823 681 2857
rect 715 2823 749 2857
rect 783 2823 817 2857
rect 851 2823 885 2857
rect 919 2823 953 2857
rect 987 2823 1021 2857
rect 1055 2823 1089 2857
rect 1123 2823 1157 2857
rect 1191 2823 1225 2857
rect 1259 2823 1293 2857
rect 1327 2823 1361 2857
rect 1395 2823 1429 2857
rect 1463 2823 1497 2857
rect 1531 2823 1565 2857
rect 1599 2823 1633 2857
rect 1667 2823 1701 2857
rect 1735 2823 1769 2857
rect 1803 2823 1837 2857
rect 1871 2823 1905 2857
rect 1939 2823 1973 2857
rect 2007 2823 2041 2857
rect 2075 2823 2109 2857
rect 2143 2823 2177 2857
rect 2211 2823 2245 2857
rect 2279 2823 2313 2857
rect 2347 2823 2381 2857
rect 2415 2823 2449 2857
rect 2483 2823 2517 2857
rect 2551 2823 2585 2857
rect 2619 2823 2653 2857
rect 2687 2823 2721 2857
rect 2755 2823 2789 2857
rect 2823 2823 2857 2857
rect 2891 2823 2925 2857
rect 2959 2823 2993 2857
rect 3027 2823 3061 2857
rect 3095 2823 3129 2857
rect 3163 2823 3197 2857
rect 3231 2823 3265 2857
rect 3299 2823 3333 2857
rect 3367 2823 3401 2857
rect 3435 2823 3469 2857
rect 3503 2823 3537 2857
rect 3571 2823 3605 2857
rect 3639 2823 3673 2857
rect 3707 2823 3741 2857
rect 3775 2823 3809 2857
rect 3843 2823 3877 2857
rect 3911 2823 3945 2857
rect 3979 2823 4013 2857
rect 4047 2823 4081 2857
rect 4115 2823 4149 2857
rect 4183 2823 4217 2857
rect 4251 2823 4285 2857
rect 4319 2823 4353 2857
rect 4387 2823 4421 2857
rect 4455 2823 4489 2857
rect 4523 2823 4557 2857
rect 4591 2823 4625 2857
rect 4659 2823 4693 2857
rect 4727 2823 4761 2857
rect 4795 2823 4829 2857
rect 4863 2823 4897 2857
rect 4931 2823 4965 2857
rect 4999 2823 5033 2857
rect 5067 2823 5101 2857
rect 5135 2823 5169 2857
rect 5203 2823 5237 2857
rect 5271 2823 5305 2857
rect 5339 2823 5373 2857
rect 5407 2823 5441 2857
rect 5475 2823 5509 2857
rect 5543 2823 5577 2857
rect 5611 2823 5645 2857
rect 5679 2823 5713 2857
rect 5747 2823 5781 2857
rect 5815 2823 5849 2857
rect 5883 2823 5917 2857
rect 5951 2823 5985 2857
rect 6019 2823 6053 2857
rect 6087 2823 6121 2857
rect 6155 2823 6189 2857
rect 6223 2823 6257 2857
rect 6291 2823 6325 2857
rect 6359 2823 6393 2857
rect 6427 2823 6461 2857
rect 6495 2823 6529 2857
rect 6563 2823 6597 2857
rect 6631 2823 6665 2857
rect 6699 2823 6733 2857
rect 6767 2823 6801 2857
rect 6835 2823 6869 2857
rect 6903 2823 6937 2857
rect 6971 2823 7005 2857
rect 7039 2823 7073 2857
rect 7107 2823 7141 2857
rect 7175 2823 7209 2857
rect 7243 2823 7277 2857
rect 7311 2823 7345 2857
rect 7379 2823 7413 2857
rect 7447 2823 7481 2857
rect 7515 2823 7549 2857
rect 7583 2823 7617 2857
rect 7651 2823 7685 2857
rect 7719 2823 7753 2857
rect 7787 2823 7821 2857
rect 7855 2823 7889 2857
rect 7923 2823 7957 2857
rect 7991 2823 8025 2857
rect 8059 2823 8093 2857
rect 307 2343 341 2377
rect 375 2343 409 2377
rect 443 2343 477 2377
rect 511 2343 545 2377
rect 579 2343 613 2377
rect 647 2343 681 2377
rect 715 2343 749 2377
rect 783 2343 817 2377
rect 851 2343 885 2377
rect 919 2343 953 2377
rect 987 2343 1021 2377
rect 1055 2343 1089 2377
rect 1123 2343 1157 2377
rect 1191 2343 1225 2377
rect 1259 2343 1293 2377
rect 1327 2343 1361 2377
rect 1395 2343 1429 2377
rect 1463 2343 1497 2377
rect 1531 2343 1565 2377
rect 1599 2343 1633 2377
rect 1667 2343 1701 2377
rect 1735 2343 1769 2377
rect 1803 2343 1837 2377
rect 1871 2343 1905 2377
rect 1939 2343 1973 2377
rect 2007 2343 2041 2377
rect 2075 2343 2109 2377
rect 2143 2343 2177 2377
rect 2211 2343 2245 2377
rect 2279 2343 2313 2377
rect 2347 2343 2381 2377
rect 2415 2343 2449 2377
rect 2483 2343 2517 2377
rect 2551 2343 2585 2377
rect 2619 2343 2653 2377
rect 2687 2343 2721 2377
rect 2755 2343 2789 2377
rect 2823 2343 2857 2377
rect 2891 2343 2925 2377
rect 2959 2343 2993 2377
rect 3027 2343 3061 2377
rect 3095 2343 3129 2377
rect 3163 2343 3197 2377
rect 3231 2343 3265 2377
rect 3299 2343 3333 2377
rect 3367 2343 3401 2377
rect 3435 2343 3469 2377
rect 3503 2343 3537 2377
rect 3571 2343 3605 2377
rect 3639 2343 3673 2377
rect 3707 2343 3741 2377
rect 3775 2343 3809 2377
rect 3843 2343 3877 2377
rect 3911 2343 3945 2377
rect 3979 2343 4013 2377
rect 4047 2343 4081 2377
rect 4115 2343 4149 2377
rect 4183 2343 4217 2377
rect 4251 2343 4285 2377
rect 4319 2343 4353 2377
rect 4387 2343 4421 2377
rect 4455 2343 4489 2377
rect 4523 2343 4557 2377
rect 4591 2343 4625 2377
rect 4659 2343 4693 2377
rect 4727 2343 4761 2377
rect 4795 2343 4829 2377
rect 4863 2343 4897 2377
rect 4931 2343 4965 2377
rect 4999 2343 5033 2377
rect 5067 2343 5101 2377
rect 5135 2343 5169 2377
rect 5203 2343 5237 2377
rect 5271 2343 5305 2377
rect 5339 2343 5373 2377
rect 5407 2343 5441 2377
rect 5475 2343 5509 2377
rect 5543 2343 5577 2377
rect 5611 2343 5645 2377
rect 5679 2343 5713 2377
rect 5747 2343 5781 2377
rect 5815 2343 5849 2377
rect 5883 2343 5917 2377
rect 5951 2343 5985 2377
rect 6019 2343 6053 2377
rect 6087 2343 6121 2377
rect 6155 2343 6189 2377
rect 6223 2343 6257 2377
rect 6291 2343 6325 2377
rect 6359 2343 6393 2377
rect 6427 2343 6461 2377
rect 6495 2343 6529 2377
rect 6563 2343 6597 2377
rect 6631 2343 6665 2377
rect 6699 2343 6733 2377
rect 6767 2343 6801 2377
rect 6835 2343 6869 2377
rect 6903 2343 6937 2377
rect 6971 2343 7005 2377
rect 7039 2343 7073 2377
rect 7107 2343 7141 2377
rect 7175 2343 7209 2377
rect 7243 2343 7277 2377
rect 7311 2343 7345 2377
rect 7379 2343 7413 2377
rect 7447 2343 7481 2377
rect 7515 2343 7549 2377
rect 7583 2343 7617 2377
rect 7651 2343 7685 2377
rect 7719 2343 7753 2377
rect 7787 2343 7821 2377
rect 7855 2343 7889 2377
rect 7923 2343 7957 2377
rect 7991 2343 8025 2377
rect 8059 2343 8093 2377
rect 183 2237 217 2271
rect 183 2169 217 2203
rect 183 2101 217 2135
rect 183 2033 217 2067
rect 183 1965 217 1999
rect 183 1897 217 1931
rect 183 1829 217 1863
rect 183 1761 217 1795
rect 183 1693 217 1727
rect 183 1625 217 1659
rect 8183 2237 8217 2271
rect 8183 2169 8217 2203
rect 8183 2101 8217 2135
rect 8183 2033 8217 2067
rect 8183 1965 8217 1999
rect 8183 1897 8217 1931
rect 8183 1829 8217 1863
rect 8183 1761 8217 1795
rect 8183 1693 8217 1727
rect 183 1557 217 1591
rect 183 1489 217 1523
rect 8183 1625 8217 1659
rect 8183 1557 8217 1591
rect 8183 1489 8217 1523
rect 307 1383 341 1417
rect 375 1383 409 1417
rect 443 1383 477 1417
rect 511 1383 545 1417
rect 579 1383 613 1417
rect 647 1383 681 1417
rect 715 1383 749 1417
rect 783 1383 817 1417
rect 851 1383 885 1417
rect 919 1383 953 1417
rect 987 1383 1021 1417
rect 1055 1383 1089 1417
rect 1123 1383 1157 1417
rect 1191 1383 1225 1417
rect 1259 1383 1293 1417
rect 1327 1383 1361 1417
rect 1395 1383 1429 1417
rect 1463 1383 1497 1417
rect 1531 1383 1565 1417
rect 1599 1383 1633 1417
rect 1667 1383 1701 1417
rect 1735 1383 1769 1417
rect 1803 1383 1837 1417
rect 1871 1383 1905 1417
rect 1939 1383 1973 1417
rect 2007 1383 2041 1417
rect 2075 1383 2109 1417
rect 2143 1383 2177 1417
rect 2211 1383 2245 1417
rect 2279 1383 2313 1417
rect 2347 1383 2381 1417
rect 2415 1383 2449 1417
rect 2483 1383 2517 1417
rect 2551 1383 2585 1417
rect 2619 1383 2653 1417
rect 2687 1383 2721 1417
rect 2755 1383 2789 1417
rect 2823 1383 2857 1417
rect 2891 1383 2925 1417
rect 2959 1383 2993 1417
rect 3027 1383 3061 1417
rect 3095 1383 3129 1417
rect 3163 1383 3197 1417
rect 3231 1383 3265 1417
rect 3299 1383 3333 1417
rect 3367 1383 3401 1417
rect 3435 1383 3469 1417
rect 3503 1383 3537 1417
rect 3571 1383 3605 1417
rect 3639 1383 3673 1417
rect 3707 1383 3741 1417
rect 3775 1383 3809 1417
rect 3843 1383 3877 1417
rect 3911 1383 3945 1417
rect 3979 1383 4013 1417
rect 4047 1383 4081 1417
rect 4115 1383 4149 1417
rect 4183 1383 4217 1417
rect 4251 1383 4285 1417
rect 4319 1383 4353 1417
rect 4387 1383 4421 1417
rect 4455 1383 4489 1417
rect 4523 1383 4557 1417
rect 4591 1383 4625 1417
rect 4659 1383 4693 1417
rect 4727 1383 4761 1417
rect 4795 1383 4829 1417
rect 4863 1383 4897 1417
rect 4931 1383 4965 1417
rect 4999 1383 5033 1417
rect 5067 1383 5101 1417
rect 5135 1383 5169 1417
rect 5203 1383 5237 1417
rect 5271 1383 5305 1417
rect 5339 1383 5373 1417
rect 5407 1383 5441 1417
rect 5475 1383 5509 1417
rect 5543 1383 5577 1417
rect 5611 1383 5645 1417
rect 5679 1383 5713 1417
rect 5747 1383 5781 1417
rect 5815 1383 5849 1417
rect 5883 1383 5917 1417
rect 5951 1383 5985 1417
rect 6019 1383 6053 1417
rect 6087 1383 6121 1417
rect 6155 1383 6189 1417
rect 6223 1383 6257 1417
rect 6291 1383 6325 1417
rect 6359 1383 6393 1417
rect 6427 1383 6461 1417
rect 6495 1383 6529 1417
rect 6563 1383 6597 1417
rect 6631 1383 6665 1417
rect 6699 1383 6733 1417
rect 6767 1383 6801 1417
rect 6835 1383 6869 1417
rect 6903 1383 6937 1417
rect 6971 1383 7005 1417
rect 7039 1383 7073 1417
rect 7107 1383 7141 1417
rect 7175 1383 7209 1417
rect 7243 1383 7277 1417
rect 7311 1383 7345 1417
rect 7379 1383 7413 1417
rect 7447 1383 7481 1417
rect 7515 1383 7549 1417
rect 7583 1383 7617 1417
rect 7651 1383 7685 1417
rect 7719 1383 7753 1417
rect 7787 1383 7821 1417
rect 7855 1383 7889 1417
rect 7923 1383 7957 1417
rect 7991 1383 8025 1417
rect 8059 1383 8093 1417
<< poly >>
rect 520 9760 2120 9800
rect 2440 9760 4040 9800
rect 4360 9760 5960 9800
rect 6280 9760 7880 9800
rect 520 9097 2120 9160
rect 520 9063 555 9097
rect 589 9063 623 9097
rect 657 9063 691 9097
rect 725 9063 759 9097
rect 793 9063 827 9097
rect 861 9063 895 9097
rect 929 9063 963 9097
rect 997 9063 1031 9097
rect 1065 9063 1099 9097
rect 1133 9063 1167 9097
rect 1201 9063 1235 9097
rect 1269 9063 1303 9097
rect 1337 9063 1371 9097
rect 1405 9063 1439 9097
rect 1473 9063 1507 9097
rect 1541 9063 1575 9097
rect 1609 9063 1643 9097
rect 1677 9063 1711 9097
rect 1745 9063 1779 9097
rect 1813 9063 1847 9097
rect 1881 9063 1915 9097
rect 1949 9063 1983 9097
rect 2017 9063 2051 9097
rect 2085 9063 2120 9097
rect 520 9040 2120 9063
rect 2440 9097 4040 9160
rect 2440 9063 2475 9097
rect 2509 9063 2543 9097
rect 2577 9063 2611 9097
rect 2645 9063 2679 9097
rect 2713 9063 2747 9097
rect 2781 9063 2815 9097
rect 2849 9063 2883 9097
rect 2917 9063 2951 9097
rect 2985 9063 3019 9097
rect 3053 9063 3087 9097
rect 3121 9063 3155 9097
rect 3189 9063 3223 9097
rect 3257 9063 3291 9097
rect 3325 9063 3359 9097
rect 3393 9063 3427 9097
rect 3461 9063 3495 9097
rect 3529 9063 3563 9097
rect 3597 9063 3631 9097
rect 3665 9063 3699 9097
rect 3733 9063 3767 9097
rect 3801 9063 3835 9097
rect 3869 9063 3903 9097
rect 3937 9063 3971 9097
rect 4005 9063 4040 9097
rect 2440 9040 4040 9063
rect 4360 9097 5960 9160
rect 4360 9063 4395 9097
rect 4429 9063 4463 9097
rect 4497 9063 4531 9097
rect 4565 9063 4599 9097
rect 4633 9063 4667 9097
rect 4701 9063 4735 9097
rect 4769 9063 4803 9097
rect 4837 9063 4871 9097
rect 4905 9063 4939 9097
rect 4973 9063 5007 9097
rect 5041 9063 5075 9097
rect 5109 9063 5143 9097
rect 5177 9063 5211 9097
rect 5245 9063 5279 9097
rect 5313 9063 5347 9097
rect 5381 9063 5415 9097
rect 5449 9063 5483 9097
rect 5517 9063 5551 9097
rect 5585 9063 5619 9097
rect 5653 9063 5687 9097
rect 5721 9063 5755 9097
rect 5789 9063 5823 9097
rect 5857 9063 5891 9097
rect 5925 9063 5960 9097
rect 4360 9040 5960 9063
rect 6280 9097 7880 9160
rect 6280 9063 6315 9097
rect 6349 9063 6383 9097
rect 6417 9063 6451 9097
rect 6485 9063 6519 9097
rect 6553 9063 6587 9097
rect 6621 9063 6655 9097
rect 6689 9063 6723 9097
rect 6757 9063 6791 9097
rect 6825 9063 6859 9097
rect 6893 9063 6927 9097
rect 6961 9063 6995 9097
rect 7029 9063 7063 9097
rect 7097 9063 7131 9097
rect 7165 9063 7199 9097
rect 7233 9063 7267 9097
rect 7301 9063 7335 9097
rect 7369 9063 7403 9097
rect 7437 9063 7471 9097
rect 7505 9063 7539 9097
rect 7573 9063 7607 9097
rect 7641 9063 7675 9097
rect 7709 9063 7743 9097
rect 7777 9063 7811 9097
rect 7845 9063 7880 9097
rect 6280 9040 7880 9063
rect 520 7817 2120 7840
rect 520 7783 555 7817
rect 589 7783 623 7817
rect 657 7783 691 7817
rect 725 7783 759 7817
rect 793 7783 827 7817
rect 861 7783 895 7817
rect 929 7783 963 7817
rect 997 7783 1031 7817
rect 1065 7783 1099 7817
rect 1133 7783 1167 7817
rect 1201 7783 1235 7817
rect 1269 7783 1303 7817
rect 1337 7783 1371 7817
rect 1405 7783 1439 7817
rect 1473 7783 1507 7817
rect 1541 7783 1575 7817
rect 1609 7783 1643 7817
rect 1677 7783 1711 7817
rect 1745 7783 1779 7817
rect 1813 7783 1847 7817
rect 1881 7783 1915 7817
rect 1949 7783 1983 7817
rect 2017 7783 2051 7817
rect 2085 7783 2120 7817
rect 520 7720 2120 7783
rect 2440 7817 4040 7840
rect 2440 7783 2475 7817
rect 2509 7783 2543 7817
rect 2577 7783 2611 7817
rect 2645 7783 2679 7817
rect 2713 7783 2747 7817
rect 2781 7783 2815 7817
rect 2849 7783 2883 7817
rect 2917 7783 2951 7817
rect 2985 7783 3019 7817
rect 3053 7783 3087 7817
rect 3121 7783 3155 7817
rect 3189 7783 3223 7817
rect 3257 7783 3291 7817
rect 3325 7783 3359 7817
rect 3393 7783 3427 7817
rect 3461 7783 3495 7817
rect 3529 7783 3563 7817
rect 3597 7783 3631 7817
rect 3665 7783 3699 7817
rect 3733 7783 3767 7817
rect 3801 7783 3835 7817
rect 3869 7783 3903 7817
rect 3937 7783 3971 7817
rect 4005 7783 4040 7817
rect 2440 7720 4040 7783
rect 4360 7817 5960 7840
rect 4360 7783 4395 7817
rect 4429 7783 4463 7817
rect 4497 7783 4531 7817
rect 4565 7783 4599 7817
rect 4633 7783 4667 7817
rect 4701 7783 4735 7817
rect 4769 7783 4803 7817
rect 4837 7783 4871 7817
rect 4905 7783 4939 7817
rect 4973 7783 5007 7817
rect 5041 7783 5075 7817
rect 5109 7783 5143 7817
rect 5177 7783 5211 7817
rect 5245 7783 5279 7817
rect 5313 7783 5347 7817
rect 5381 7783 5415 7817
rect 5449 7783 5483 7817
rect 5517 7783 5551 7817
rect 5585 7783 5619 7817
rect 5653 7783 5687 7817
rect 5721 7783 5755 7817
rect 5789 7783 5823 7817
rect 5857 7783 5891 7817
rect 5925 7783 5960 7817
rect 4360 7720 5960 7783
rect 6280 7817 7880 7840
rect 6280 7783 6315 7817
rect 6349 7783 6383 7817
rect 6417 7783 6451 7817
rect 6485 7783 6519 7817
rect 6553 7783 6587 7817
rect 6621 7783 6655 7817
rect 6689 7783 6723 7817
rect 6757 7783 6791 7817
rect 6825 7783 6859 7817
rect 6893 7783 6927 7817
rect 6961 7783 6995 7817
rect 7029 7783 7063 7817
rect 7097 7783 7131 7817
rect 7165 7783 7199 7817
rect 7233 7783 7267 7817
rect 7301 7783 7335 7817
rect 7369 7783 7403 7817
rect 7437 7783 7471 7817
rect 7505 7783 7539 7817
rect 7573 7783 7607 7817
rect 7641 7783 7675 7817
rect 7709 7783 7743 7817
rect 7777 7783 7811 7817
rect 7845 7783 7880 7817
rect 6280 7720 7880 7783
rect 520 7480 2120 7520
rect 2440 7480 4040 7520
rect 4360 7480 5960 7520
rect 6280 7480 7880 7520
rect 520 7120 2120 7160
rect 2440 7120 4040 7160
rect 4360 7120 5960 7160
rect 6280 7120 7880 7160
rect 520 6857 2120 6920
rect 520 6823 555 6857
rect 589 6823 623 6857
rect 657 6823 691 6857
rect 725 6823 759 6857
rect 793 6823 827 6857
rect 861 6823 895 6857
rect 929 6823 963 6857
rect 997 6823 1031 6857
rect 1065 6823 1099 6857
rect 1133 6823 1167 6857
rect 1201 6823 1235 6857
rect 1269 6823 1303 6857
rect 1337 6823 1371 6857
rect 1405 6823 1439 6857
rect 1473 6823 1507 6857
rect 1541 6823 1575 6857
rect 1609 6823 1643 6857
rect 1677 6823 1711 6857
rect 1745 6823 1779 6857
rect 1813 6823 1847 6857
rect 1881 6823 1915 6857
rect 1949 6823 1983 6857
rect 2017 6823 2051 6857
rect 2085 6823 2120 6857
rect 520 6800 2120 6823
rect 2440 6857 4040 6920
rect 2440 6823 2475 6857
rect 2509 6823 2543 6857
rect 2577 6823 2611 6857
rect 2645 6823 2679 6857
rect 2713 6823 2747 6857
rect 2781 6823 2815 6857
rect 2849 6823 2883 6857
rect 2917 6823 2951 6857
rect 2985 6823 3019 6857
rect 3053 6823 3087 6857
rect 3121 6823 3155 6857
rect 3189 6823 3223 6857
rect 3257 6823 3291 6857
rect 3325 6823 3359 6857
rect 3393 6823 3427 6857
rect 3461 6823 3495 6857
rect 3529 6823 3563 6857
rect 3597 6823 3631 6857
rect 3665 6823 3699 6857
rect 3733 6823 3767 6857
rect 3801 6823 3835 6857
rect 3869 6823 3903 6857
rect 3937 6823 3971 6857
rect 4005 6823 4040 6857
rect 2440 6800 4040 6823
rect 4360 6857 5960 6920
rect 4360 6823 4395 6857
rect 4429 6823 4463 6857
rect 4497 6823 4531 6857
rect 4565 6823 4599 6857
rect 4633 6823 4667 6857
rect 4701 6823 4735 6857
rect 4769 6823 4803 6857
rect 4837 6823 4871 6857
rect 4905 6823 4939 6857
rect 4973 6823 5007 6857
rect 5041 6823 5075 6857
rect 5109 6823 5143 6857
rect 5177 6823 5211 6857
rect 5245 6823 5279 6857
rect 5313 6823 5347 6857
rect 5381 6823 5415 6857
rect 5449 6823 5483 6857
rect 5517 6823 5551 6857
rect 5585 6823 5619 6857
rect 5653 6823 5687 6857
rect 5721 6823 5755 6857
rect 5789 6823 5823 6857
rect 5857 6823 5891 6857
rect 5925 6823 5960 6857
rect 4360 6800 5960 6823
rect 6280 6857 7880 6920
rect 6280 6823 6315 6857
rect 6349 6823 6383 6857
rect 6417 6823 6451 6857
rect 6485 6823 6519 6857
rect 6553 6823 6587 6857
rect 6621 6823 6655 6857
rect 6689 6823 6723 6857
rect 6757 6823 6791 6857
rect 6825 6823 6859 6857
rect 6893 6823 6927 6857
rect 6961 6823 6995 6857
rect 7029 6823 7063 6857
rect 7097 6823 7131 6857
rect 7165 6823 7199 6857
rect 7233 6823 7267 6857
rect 7301 6823 7335 6857
rect 7369 6823 7403 6857
rect 7437 6823 7471 6857
rect 7505 6823 7539 6857
rect 7573 6823 7607 6857
rect 7641 6823 7675 6857
rect 7709 6823 7743 6857
rect 7777 6823 7811 6857
rect 7845 6823 7880 6857
rect 6280 6800 7880 6823
rect 520 5097 2120 5120
rect 520 5063 555 5097
rect 589 5063 623 5097
rect 657 5063 691 5097
rect 725 5063 759 5097
rect 793 5063 827 5097
rect 861 5063 895 5097
rect 929 5063 963 5097
rect 997 5063 1031 5097
rect 1065 5063 1099 5097
rect 1133 5063 1167 5097
rect 1201 5063 1235 5097
rect 1269 5063 1303 5097
rect 1337 5063 1371 5097
rect 1405 5063 1439 5097
rect 1473 5063 1507 5097
rect 1541 5063 1575 5097
rect 1609 5063 1643 5097
rect 1677 5063 1711 5097
rect 1745 5063 1779 5097
rect 1813 5063 1847 5097
rect 1881 5063 1915 5097
rect 1949 5063 1983 5097
rect 2017 5063 2051 5097
rect 2085 5063 2120 5097
rect 520 5000 2120 5063
rect 2440 5097 4040 5120
rect 2440 5063 2475 5097
rect 2509 5063 2543 5097
rect 2577 5063 2611 5097
rect 2645 5063 2679 5097
rect 2713 5063 2747 5097
rect 2781 5063 2815 5097
rect 2849 5063 2883 5097
rect 2917 5063 2951 5097
rect 2985 5063 3019 5097
rect 3053 5063 3087 5097
rect 3121 5063 3155 5097
rect 3189 5063 3223 5097
rect 3257 5063 3291 5097
rect 3325 5063 3359 5097
rect 3393 5063 3427 5097
rect 3461 5063 3495 5097
rect 3529 5063 3563 5097
rect 3597 5063 3631 5097
rect 3665 5063 3699 5097
rect 3733 5063 3767 5097
rect 3801 5063 3835 5097
rect 3869 5063 3903 5097
rect 3937 5063 3971 5097
rect 4005 5063 4040 5097
rect 2440 5000 4040 5063
rect 4360 5097 5960 5120
rect 4360 5063 4395 5097
rect 4429 5063 4463 5097
rect 4497 5063 4531 5097
rect 4565 5063 4599 5097
rect 4633 5063 4667 5097
rect 4701 5063 4735 5097
rect 4769 5063 4803 5097
rect 4837 5063 4871 5097
rect 4905 5063 4939 5097
rect 4973 5063 5007 5097
rect 5041 5063 5075 5097
rect 5109 5063 5143 5097
rect 5177 5063 5211 5097
rect 5245 5063 5279 5097
rect 5313 5063 5347 5097
rect 5381 5063 5415 5097
rect 5449 5063 5483 5097
rect 5517 5063 5551 5097
rect 5585 5063 5619 5097
rect 5653 5063 5687 5097
rect 5721 5063 5755 5097
rect 5789 5063 5823 5097
rect 5857 5063 5891 5097
rect 5925 5063 5960 5097
rect 4360 5000 5960 5063
rect 6280 5097 7880 5120
rect 6280 5063 6315 5097
rect 6349 5063 6383 5097
rect 6417 5063 6451 5097
rect 6485 5063 6519 5097
rect 6553 5063 6587 5097
rect 6621 5063 6655 5097
rect 6689 5063 6723 5097
rect 6757 5063 6791 5097
rect 6825 5063 6859 5097
rect 6893 5063 6927 5097
rect 6961 5063 6995 5097
rect 7029 5063 7063 5097
rect 7097 5063 7131 5097
rect 7165 5063 7199 5097
rect 7233 5063 7267 5097
rect 7301 5063 7335 5097
rect 7369 5063 7403 5097
rect 7437 5063 7471 5097
rect 7505 5063 7539 5097
rect 7573 5063 7607 5097
rect 7641 5063 7675 5097
rect 7709 5063 7743 5097
rect 7777 5063 7811 5097
rect 7845 5063 7880 5097
rect 6280 5000 7880 5063
rect 520 4360 2120 4400
rect 2440 4360 4040 4400
rect 4360 4360 5960 4400
rect 6280 4360 7880 4400
rect 520 3680 2120 3720
rect 2440 3680 4040 3720
rect 4360 3680 5960 3720
rect 6280 3680 7880 3720
rect 520 3017 2120 3080
rect 520 2983 555 3017
rect 589 2983 623 3017
rect 657 2983 691 3017
rect 725 2983 759 3017
rect 793 2983 827 3017
rect 861 2983 895 3017
rect 929 2983 963 3017
rect 997 2983 1031 3017
rect 1065 2983 1099 3017
rect 1133 2983 1167 3017
rect 1201 2983 1235 3017
rect 1269 2983 1303 3017
rect 1337 2983 1371 3017
rect 1405 2983 1439 3017
rect 1473 2983 1507 3017
rect 1541 2983 1575 3017
rect 1609 2983 1643 3017
rect 1677 2983 1711 3017
rect 1745 2983 1779 3017
rect 1813 2983 1847 3017
rect 1881 2983 1915 3017
rect 1949 2983 1983 3017
rect 2017 2983 2051 3017
rect 2085 2983 2120 3017
rect 520 2960 2120 2983
rect 2440 3017 4040 3080
rect 2440 2983 2475 3017
rect 2509 2983 2543 3017
rect 2577 2983 2611 3017
rect 2645 2983 2679 3017
rect 2713 2983 2747 3017
rect 2781 2983 2815 3017
rect 2849 2983 2883 3017
rect 2917 2983 2951 3017
rect 2985 2983 3019 3017
rect 3053 2983 3087 3017
rect 3121 2983 3155 3017
rect 3189 2983 3223 3017
rect 3257 2983 3291 3017
rect 3325 2983 3359 3017
rect 3393 2983 3427 3017
rect 3461 2983 3495 3017
rect 3529 2983 3563 3017
rect 3597 2983 3631 3017
rect 3665 2983 3699 3017
rect 3733 2983 3767 3017
rect 3801 2983 3835 3017
rect 3869 2983 3903 3017
rect 3937 2983 3971 3017
rect 4005 2983 4040 3017
rect 2440 2960 4040 2983
rect 4360 3017 5960 3080
rect 4360 2983 4395 3017
rect 4429 2983 4463 3017
rect 4497 2983 4531 3017
rect 4565 2983 4599 3017
rect 4633 2983 4667 3017
rect 4701 2983 4735 3017
rect 4769 2983 4803 3017
rect 4837 2983 4871 3017
rect 4905 2983 4939 3017
rect 4973 2983 5007 3017
rect 5041 2983 5075 3017
rect 5109 2983 5143 3017
rect 5177 2983 5211 3017
rect 5245 2983 5279 3017
rect 5313 2983 5347 3017
rect 5381 2983 5415 3017
rect 5449 2983 5483 3017
rect 5517 2983 5551 3017
rect 5585 2983 5619 3017
rect 5653 2983 5687 3017
rect 5721 2983 5755 3017
rect 5789 2983 5823 3017
rect 5857 2983 5891 3017
rect 5925 2983 5960 3017
rect 4360 2960 5960 2983
rect 6280 3017 7880 3080
rect 6280 2983 6315 3017
rect 6349 2983 6383 3017
rect 6417 2983 6451 3017
rect 6485 2983 6519 3017
rect 6553 2983 6587 3017
rect 6621 2983 6655 3017
rect 6689 2983 6723 3017
rect 6757 2983 6791 3017
rect 6825 2983 6859 3017
rect 6893 2983 6927 3017
rect 6961 2983 6995 3017
rect 7029 2983 7063 3017
rect 7097 2983 7131 3017
rect 7165 2983 7199 3017
rect 7233 2983 7267 3017
rect 7301 2983 7335 3017
rect 7369 2983 7403 3017
rect 7437 2983 7471 3017
rect 7505 2983 7539 3017
rect 7573 2983 7607 3017
rect 7641 2983 7675 3017
rect 7709 2983 7743 3017
rect 7777 2983 7811 3017
rect 7845 2983 7880 3017
rect 6280 2960 7880 2983
rect 520 2240 2120 2280
rect 2440 2240 4040 2280
rect 4360 2240 5960 2280
rect 6280 2240 7880 2280
rect 520 1577 2120 1640
rect 520 1543 555 1577
rect 589 1543 623 1577
rect 657 1543 691 1577
rect 725 1543 759 1577
rect 793 1543 827 1577
rect 861 1543 895 1577
rect 929 1543 963 1577
rect 997 1543 1031 1577
rect 1065 1543 1099 1577
rect 1133 1543 1167 1577
rect 1201 1543 1235 1577
rect 1269 1543 1303 1577
rect 1337 1543 1371 1577
rect 1405 1543 1439 1577
rect 1473 1543 1507 1577
rect 1541 1543 1575 1577
rect 1609 1543 1643 1577
rect 1677 1543 1711 1577
rect 1745 1543 1779 1577
rect 1813 1543 1847 1577
rect 1881 1543 1915 1577
rect 1949 1543 1983 1577
rect 2017 1543 2051 1577
rect 2085 1543 2120 1577
rect 520 1520 2120 1543
rect 2440 1577 4040 1640
rect 2440 1543 2475 1577
rect 2509 1543 2543 1577
rect 2577 1543 2611 1577
rect 2645 1543 2679 1577
rect 2713 1543 2747 1577
rect 2781 1543 2815 1577
rect 2849 1543 2883 1577
rect 2917 1543 2951 1577
rect 2985 1543 3019 1577
rect 3053 1543 3087 1577
rect 3121 1543 3155 1577
rect 3189 1543 3223 1577
rect 3257 1543 3291 1577
rect 3325 1543 3359 1577
rect 3393 1543 3427 1577
rect 3461 1543 3495 1577
rect 3529 1543 3563 1577
rect 3597 1543 3631 1577
rect 3665 1543 3699 1577
rect 3733 1543 3767 1577
rect 3801 1543 3835 1577
rect 3869 1543 3903 1577
rect 3937 1543 3971 1577
rect 4005 1543 4040 1577
rect 2440 1520 4040 1543
rect 4360 1577 5960 1640
rect 4360 1543 4395 1577
rect 4429 1543 4463 1577
rect 4497 1543 4531 1577
rect 4565 1543 4599 1577
rect 4633 1543 4667 1577
rect 4701 1543 4735 1577
rect 4769 1543 4803 1577
rect 4837 1543 4871 1577
rect 4905 1543 4939 1577
rect 4973 1543 5007 1577
rect 5041 1543 5075 1577
rect 5109 1543 5143 1577
rect 5177 1543 5211 1577
rect 5245 1543 5279 1577
rect 5313 1543 5347 1577
rect 5381 1543 5415 1577
rect 5449 1543 5483 1577
rect 5517 1543 5551 1577
rect 5585 1543 5619 1577
rect 5653 1543 5687 1577
rect 5721 1543 5755 1577
rect 5789 1543 5823 1577
rect 5857 1543 5891 1577
rect 5925 1543 5960 1577
rect 4360 1520 5960 1543
rect 6280 1577 7880 1640
rect 6280 1543 6315 1577
rect 6349 1543 6383 1577
rect 6417 1543 6451 1577
rect 6485 1543 6519 1577
rect 6553 1543 6587 1577
rect 6621 1543 6655 1577
rect 6689 1543 6723 1577
rect 6757 1543 6791 1577
rect 6825 1543 6859 1577
rect 6893 1543 6927 1577
rect 6961 1543 6995 1577
rect 7029 1543 7063 1577
rect 7097 1543 7131 1577
rect 7165 1543 7199 1577
rect 7233 1543 7267 1577
rect 7301 1543 7335 1577
rect 7369 1543 7403 1577
rect 7437 1543 7471 1577
rect 7505 1543 7539 1577
rect 7573 1543 7607 1577
rect 7641 1543 7675 1577
rect 7709 1543 7743 1577
rect 7777 1543 7811 1577
rect 7845 1543 7880 1577
rect 6280 1520 7880 1543
rect 520 457 2120 480
rect 520 423 555 457
rect 589 423 623 457
rect 657 423 691 457
rect 725 423 759 457
rect 793 423 827 457
rect 861 423 895 457
rect 929 423 963 457
rect 997 423 1031 457
rect 1065 423 1099 457
rect 1133 423 1167 457
rect 1201 423 1235 457
rect 1269 423 1303 457
rect 1337 423 1371 457
rect 1405 423 1439 457
rect 1473 423 1507 457
rect 1541 423 1575 457
rect 1609 423 1643 457
rect 1677 423 1711 457
rect 1745 423 1779 457
rect 1813 423 1847 457
rect 1881 423 1915 457
rect 1949 423 1983 457
rect 2017 423 2051 457
rect 2085 423 2120 457
rect 520 360 2120 423
rect 2440 457 4040 480
rect 2440 423 2475 457
rect 2509 423 2543 457
rect 2577 423 2611 457
rect 2645 423 2679 457
rect 2713 423 2747 457
rect 2781 423 2815 457
rect 2849 423 2883 457
rect 2917 423 2951 457
rect 2985 423 3019 457
rect 3053 423 3087 457
rect 3121 423 3155 457
rect 3189 423 3223 457
rect 3257 423 3291 457
rect 3325 423 3359 457
rect 3393 423 3427 457
rect 3461 423 3495 457
rect 3529 423 3563 457
rect 3597 423 3631 457
rect 3665 423 3699 457
rect 3733 423 3767 457
rect 3801 423 3835 457
rect 3869 423 3903 457
rect 3937 423 3971 457
rect 4005 423 4040 457
rect 2440 360 4040 423
rect 4360 457 5960 480
rect 4360 423 4395 457
rect 4429 423 4463 457
rect 4497 423 4531 457
rect 4565 423 4599 457
rect 4633 423 4667 457
rect 4701 423 4735 457
rect 4769 423 4803 457
rect 4837 423 4871 457
rect 4905 423 4939 457
rect 4973 423 5007 457
rect 5041 423 5075 457
rect 5109 423 5143 457
rect 5177 423 5211 457
rect 5245 423 5279 457
rect 5313 423 5347 457
rect 5381 423 5415 457
rect 5449 423 5483 457
rect 5517 423 5551 457
rect 5585 423 5619 457
rect 5653 423 5687 457
rect 5721 423 5755 457
rect 5789 423 5823 457
rect 5857 423 5891 457
rect 5925 423 5960 457
rect 4360 360 5960 423
rect 6280 457 7880 480
rect 6280 423 6315 457
rect 6349 423 6383 457
rect 6417 423 6451 457
rect 6485 423 6519 457
rect 6553 423 6587 457
rect 6621 423 6655 457
rect 6689 423 6723 457
rect 6757 423 6791 457
rect 6825 423 6859 457
rect 6893 423 6927 457
rect 6961 423 6995 457
rect 7029 423 7063 457
rect 7097 423 7131 457
rect 7165 423 7199 457
rect 7233 423 7267 457
rect 7301 423 7335 457
rect 7369 423 7403 457
rect 7437 423 7471 457
rect 7505 423 7539 457
rect 7573 423 7607 457
rect 7641 423 7675 457
rect 7709 423 7743 457
rect 7777 423 7811 457
rect 7845 423 7880 457
rect 6280 360 7880 423
rect 520 120 2120 160
rect 2440 120 4040 160
rect 4360 120 5960 160
rect 6280 120 7880 160
rect 520 -583 2120 -560
rect 520 -617 555 -583
rect 589 -617 623 -583
rect 657 -617 691 -583
rect 725 -617 759 -583
rect 793 -617 827 -583
rect 861 -617 895 -583
rect 929 -617 963 -583
rect 997 -617 1031 -583
rect 1065 -617 1099 -583
rect 1133 -617 1167 -583
rect 1201 -617 1235 -583
rect 1269 -617 1303 -583
rect 1337 -617 1371 -583
rect 1405 -617 1439 -583
rect 1473 -617 1507 -583
rect 1541 -617 1575 -583
rect 1609 -617 1643 -583
rect 1677 -617 1711 -583
rect 1745 -617 1779 -583
rect 1813 -617 1847 -583
rect 1881 -617 1915 -583
rect 1949 -617 1983 -583
rect 2017 -617 2051 -583
rect 2085 -617 2120 -583
rect 520 -680 2120 -617
rect 2440 -583 4040 -560
rect 2440 -617 2475 -583
rect 2509 -617 2543 -583
rect 2577 -617 2611 -583
rect 2645 -617 2679 -583
rect 2713 -617 2747 -583
rect 2781 -617 2815 -583
rect 2849 -617 2883 -583
rect 2917 -617 2951 -583
rect 2985 -617 3019 -583
rect 3053 -617 3087 -583
rect 3121 -617 3155 -583
rect 3189 -617 3223 -583
rect 3257 -617 3291 -583
rect 3325 -617 3359 -583
rect 3393 -617 3427 -583
rect 3461 -617 3495 -583
rect 3529 -617 3563 -583
rect 3597 -617 3631 -583
rect 3665 -617 3699 -583
rect 3733 -617 3767 -583
rect 3801 -617 3835 -583
rect 3869 -617 3903 -583
rect 3937 -617 3971 -583
rect 4005 -617 4040 -583
rect 2440 -680 4040 -617
rect 4360 -583 5960 -560
rect 4360 -617 4395 -583
rect 4429 -617 4463 -583
rect 4497 -617 4531 -583
rect 4565 -617 4599 -583
rect 4633 -617 4667 -583
rect 4701 -617 4735 -583
rect 4769 -617 4803 -583
rect 4837 -617 4871 -583
rect 4905 -617 4939 -583
rect 4973 -617 5007 -583
rect 5041 -617 5075 -583
rect 5109 -617 5143 -583
rect 5177 -617 5211 -583
rect 5245 -617 5279 -583
rect 5313 -617 5347 -583
rect 5381 -617 5415 -583
rect 5449 -617 5483 -583
rect 5517 -617 5551 -583
rect 5585 -617 5619 -583
rect 5653 -617 5687 -583
rect 5721 -617 5755 -583
rect 5789 -617 5823 -583
rect 5857 -617 5891 -583
rect 5925 -617 5960 -583
rect 4360 -680 5960 -617
rect 6280 -583 7880 -560
rect 6280 -617 6315 -583
rect 6349 -617 6383 -583
rect 6417 -617 6451 -583
rect 6485 -617 6519 -583
rect 6553 -617 6587 -583
rect 6621 -617 6655 -583
rect 6689 -617 6723 -583
rect 6757 -617 6791 -583
rect 6825 -617 6859 -583
rect 6893 -617 6927 -583
rect 6961 -617 6995 -583
rect 7029 -617 7063 -583
rect 7097 -617 7131 -583
rect 7165 -617 7199 -583
rect 7233 -617 7267 -583
rect 7301 -617 7335 -583
rect 7369 -617 7403 -583
rect 7437 -617 7471 -583
rect 7505 -617 7539 -583
rect 7573 -617 7607 -583
rect 7641 -617 7675 -583
rect 7709 -617 7743 -583
rect 7777 -617 7811 -583
rect 7845 -617 7880 -583
rect 6280 -680 7880 -617
rect 520 -920 2120 -880
rect 2440 -920 4040 -880
rect 4360 -920 5960 -880
rect 6280 -920 7880 -880
<< polycont >>
rect 555 9063 589 9097
rect 623 9063 657 9097
rect 691 9063 725 9097
rect 759 9063 793 9097
rect 827 9063 861 9097
rect 895 9063 929 9097
rect 963 9063 997 9097
rect 1031 9063 1065 9097
rect 1099 9063 1133 9097
rect 1167 9063 1201 9097
rect 1235 9063 1269 9097
rect 1303 9063 1337 9097
rect 1371 9063 1405 9097
rect 1439 9063 1473 9097
rect 1507 9063 1541 9097
rect 1575 9063 1609 9097
rect 1643 9063 1677 9097
rect 1711 9063 1745 9097
rect 1779 9063 1813 9097
rect 1847 9063 1881 9097
rect 1915 9063 1949 9097
rect 1983 9063 2017 9097
rect 2051 9063 2085 9097
rect 2475 9063 2509 9097
rect 2543 9063 2577 9097
rect 2611 9063 2645 9097
rect 2679 9063 2713 9097
rect 2747 9063 2781 9097
rect 2815 9063 2849 9097
rect 2883 9063 2917 9097
rect 2951 9063 2985 9097
rect 3019 9063 3053 9097
rect 3087 9063 3121 9097
rect 3155 9063 3189 9097
rect 3223 9063 3257 9097
rect 3291 9063 3325 9097
rect 3359 9063 3393 9097
rect 3427 9063 3461 9097
rect 3495 9063 3529 9097
rect 3563 9063 3597 9097
rect 3631 9063 3665 9097
rect 3699 9063 3733 9097
rect 3767 9063 3801 9097
rect 3835 9063 3869 9097
rect 3903 9063 3937 9097
rect 3971 9063 4005 9097
rect 4395 9063 4429 9097
rect 4463 9063 4497 9097
rect 4531 9063 4565 9097
rect 4599 9063 4633 9097
rect 4667 9063 4701 9097
rect 4735 9063 4769 9097
rect 4803 9063 4837 9097
rect 4871 9063 4905 9097
rect 4939 9063 4973 9097
rect 5007 9063 5041 9097
rect 5075 9063 5109 9097
rect 5143 9063 5177 9097
rect 5211 9063 5245 9097
rect 5279 9063 5313 9097
rect 5347 9063 5381 9097
rect 5415 9063 5449 9097
rect 5483 9063 5517 9097
rect 5551 9063 5585 9097
rect 5619 9063 5653 9097
rect 5687 9063 5721 9097
rect 5755 9063 5789 9097
rect 5823 9063 5857 9097
rect 5891 9063 5925 9097
rect 6315 9063 6349 9097
rect 6383 9063 6417 9097
rect 6451 9063 6485 9097
rect 6519 9063 6553 9097
rect 6587 9063 6621 9097
rect 6655 9063 6689 9097
rect 6723 9063 6757 9097
rect 6791 9063 6825 9097
rect 6859 9063 6893 9097
rect 6927 9063 6961 9097
rect 6995 9063 7029 9097
rect 7063 9063 7097 9097
rect 7131 9063 7165 9097
rect 7199 9063 7233 9097
rect 7267 9063 7301 9097
rect 7335 9063 7369 9097
rect 7403 9063 7437 9097
rect 7471 9063 7505 9097
rect 7539 9063 7573 9097
rect 7607 9063 7641 9097
rect 7675 9063 7709 9097
rect 7743 9063 7777 9097
rect 7811 9063 7845 9097
rect 555 7783 589 7817
rect 623 7783 657 7817
rect 691 7783 725 7817
rect 759 7783 793 7817
rect 827 7783 861 7817
rect 895 7783 929 7817
rect 963 7783 997 7817
rect 1031 7783 1065 7817
rect 1099 7783 1133 7817
rect 1167 7783 1201 7817
rect 1235 7783 1269 7817
rect 1303 7783 1337 7817
rect 1371 7783 1405 7817
rect 1439 7783 1473 7817
rect 1507 7783 1541 7817
rect 1575 7783 1609 7817
rect 1643 7783 1677 7817
rect 1711 7783 1745 7817
rect 1779 7783 1813 7817
rect 1847 7783 1881 7817
rect 1915 7783 1949 7817
rect 1983 7783 2017 7817
rect 2051 7783 2085 7817
rect 2475 7783 2509 7817
rect 2543 7783 2577 7817
rect 2611 7783 2645 7817
rect 2679 7783 2713 7817
rect 2747 7783 2781 7817
rect 2815 7783 2849 7817
rect 2883 7783 2917 7817
rect 2951 7783 2985 7817
rect 3019 7783 3053 7817
rect 3087 7783 3121 7817
rect 3155 7783 3189 7817
rect 3223 7783 3257 7817
rect 3291 7783 3325 7817
rect 3359 7783 3393 7817
rect 3427 7783 3461 7817
rect 3495 7783 3529 7817
rect 3563 7783 3597 7817
rect 3631 7783 3665 7817
rect 3699 7783 3733 7817
rect 3767 7783 3801 7817
rect 3835 7783 3869 7817
rect 3903 7783 3937 7817
rect 3971 7783 4005 7817
rect 4395 7783 4429 7817
rect 4463 7783 4497 7817
rect 4531 7783 4565 7817
rect 4599 7783 4633 7817
rect 4667 7783 4701 7817
rect 4735 7783 4769 7817
rect 4803 7783 4837 7817
rect 4871 7783 4905 7817
rect 4939 7783 4973 7817
rect 5007 7783 5041 7817
rect 5075 7783 5109 7817
rect 5143 7783 5177 7817
rect 5211 7783 5245 7817
rect 5279 7783 5313 7817
rect 5347 7783 5381 7817
rect 5415 7783 5449 7817
rect 5483 7783 5517 7817
rect 5551 7783 5585 7817
rect 5619 7783 5653 7817
rect 5687 7783 5721 7817
rect 5755 7783 5789 7817
rect 5823 7783 5857 7817
rect 5891 7783 5925 7817
rect 6315 7783 6349 7817
rect 6383 7783 6417 7817
rect 6451 7783 6485 7817
rect 6519 7783 6553 7817
rect 6587 7783 6621 7817
rect 6655 7783 6689 7817
rect 6723 7783 6757 7817
rect 6791 7783 6825 7817
rect 6859 7783 6893 7817
rect 6927 7783 6961 7817
rect 6995 7783 7029 7817
rect 7063 7783 7097 7817
rect 7131 7783 7165 7817
rect 7199 7783 7233 7817
rect 7267 7783 7301 7817
rect 7335 7783 7369 7817
rect 7403 7783 7437 7817
rect 7471 7783 7505 7817
rect 7539 7783 7573 7817
rect 7607 7783 7641 7817
rect 7675 7783 7709 7817
rect 7743 7783 7777 7817
rect 7811 7783 7845 7817
rect 555 6823 589 6857
rect 623 6823 657 6857
rect 691 6823 725 6857
rect 759 6823 793 6857
rect 827 6823 861 6857
rect 895 6823 929 6857
rect 963 6823 997 6857
rect 1031 6823 1065 6857
rect 1099 6823 1133 6857
rect 1167 6823 1201 6857
rect 1235 6823 1269 6857
rect 1303 6823 1337 6857
rect 1371 6823 1405 6857
rect 1439 6823 1473 6857
rect 1507 6823 1541 6857
rect 1575 6823 1609 6857
rect 1643 6823 1677 6857
rect 1711 6823 1745 6857
rect 1779 6823 1813 6857
rect 1847 6823 1881 6857
rect 1915 6823 1949 6857
rect 1983 6823 2017 6857
rect 2051 6823 2085 6857
rect 2475 6823 2509 6857
rect 2543 6823 2577 6857
rect 2611 6823 2645 6857
rect 2679 6823 2713 6857
rect 2747 6823 2781 6857
rect 2815 6823 2849 6857
rect 2883 6823 2917 6857
rect 2951 6823 2985 6857
rect 3019 6823 3053 6857
rect 3087 6823 3121 6857
rect 3155 6823 3189 6857
rect 3223 6823 3257 6857
rect 3291 6823 3325 6857
rect 3359 6823 3393 6857
rect 3427 6823 3461 6857
rect 3495 6823 3529 6857
rect 3563 6823 3597 6857
rect 3631 6823 3665 6857
rect 3699 6823 3733 6857
rect 3767 6823 3801 6857
rect 3835 6823 3869 6857
rect 3903 6823 3937 6857
rect 3971 6823 4005 6857
rect 4395 6823 4429 6857
rect 4463 6823 4497 6857
rect 4531 6823 4565 6857
rect 4599 6823 4633 6857
rect 4667 6823 4701 6857
rect 4735 6823 4769 6857
rect 4803 6823 4837 6857
rect 4871 6823 4905 6857
rect 4939 6823 4973 6857
rect 5007 6823 5041 6857
rect 5075 6823 5109 6857
rect 5143 6823 5177 6857
rect 5211 6823 5245 6857
rect 5279 6823 5313 6857
rect 5347 6823 5381 6857
rect 5415 6823 5449 6857
rect 5483 6823 5517 6857
rect 5551 6823 5585 6857
rect 5619 6823 5653 6857
rect 5687 6823 5721 6857
rect 5755 6823 5789 6857
rect 5823 6823 5857 6857
rect 5891 6823 5925 6857
rect 6315 6823 6349 6857
rect 6383 6823 6417 6857
rect 6451 6823 6485 6857
rect 6519 6823 6553 6857
rect 6587 6823 6621 6857
rect 6655 6823 6689 6857
rect 6723 6823 6757 6857
rect 6791 6823 6825 6857
rect 6859 6823 6893 6857
rect 6927 6823 6961 6857
rect 6995 6823 7029 6857
rect 7063 6823 7097 6857
rect 7131 6823 7165 6857
rect 7199 6823 7233 6857
rect 7267 6823 7301 6857
rect 7335 6823 7369 6857
rect 7403 6823 7437 6857
rect 7471 6823 7505 6857
rect 7539 6823 7573 6857
rect 7607 6823 7641 6857
rect 7675 6823 7709 6857
rect 7743 6823 7777 6857
rect 7811 6823 7845 6857
rect 555 5063 589 5097
rect 623 5063 657 5097
rect 691 5063 725 5097
rect 759 5063 793 5097
rect 827 5063 861 5097
rect 895 5063 929 5097
rect 963 5063 997 5097
rect 1031 5063 1065 5097
rect 1099 5063 1133 5097
rect 1167 5063 1201 5097
rect 1235 5063 1269 5097
rect 1303 5063 1337 5097
rect 1371 5063 1405 5097
rect 1439 5063 1473 5097
rect 1507 5063 1541 5097
rect 1575 5063 1609 5097
rect 1643 5063 1677 5097
rect 1711 5063 1745 5097
rect 1779 5063 1813 5097
rect 1847 5063 1881 5097
rect 1915 5063 1949 5097
rect 1983 5063 2017 5097
rect 2051 5063 2085 5097
rect 2475 5063 2509 5097
rect 2543 5063 2577 5097
rect 2611 5063 2645 5097
rect 2679 5063 2713 5097
rect 2747 5063 2781 5097
rect 2815 5063 2849 5097
rect 2883 5063 2917 5097
rect 2951 5063 2985 5097
rect 3019 5063 3053 5097
rect 3087 5063 3121 5097
rect 3155 5063 3189 5097
rect 3223 5063 3257 5097
rect 3291 5063 3325 5097
rect 3359 5063 3393 5097
rect 3427 5063 3461 5097
rect 3495 5063 3529 5097
rect 3563 5063 3597 5097
rect 3631 5063 3665 5097
rect 3699 5063 3733 5097
rect 3767 5063 3801 5097
rect 3835 5063 3869 5097
rect 3903 5063 3937 5097
rect 3971 5063 4005 5097
rect 4395 5063 4429 5097
rect 4463 5063 4497 5097
rect 4531 5063 4565 5097
rect 4599 5063 4633 5097
rect 4667 5063 4701 5097
rect 4735 5063 4769 5097
rect 4803 5063 4837 5097
rect 4871 5063 4905 5097
rect 4939 5063 4973 5097
rect 5007 5063 5041 5097
rect 5075 5063 5109 5097
rect 5143 5063 5177 5097
rect 5211 5063 5245 5097
rect 5279 5063 5313 5097
rect 5347 5063 5381 5097
rect 5415 5063 5449 5097
rect 5483 5063 5517 5097
rect 5551 5063 5585 5097
rect 5619 5063 5653 5097
rect 5687 5063 5721 5097
rect 5755 5063 5789 5097
rect 5823 5063 5857 5097
rect 5891 5063 5925 5097
rect 6315 5063 6349 5097
rect 6383 5063 6417 5097
rect 6451 5063 6485 5097
rect 6519 5063 6553 5097
rect 6587 5063 6621 5097
rect 6655 5063 6689 5097
rect 6723 5063 6757 5097
rect 6791 5063 6825 5097
rect 6859 5063 6893 5097
rect 6927 5063 6961 5097
rect 6995 5063 7029 5097
rect 7063 5063 7097 5097
rect 7131 5063 7165 5097
rect 7199 5063 7233 5097
rect 7267 5063 7301 5097
rect 7335 5063 7369 5097
rect 7403 5063 7437 5097
rect 7471 5063 7505 5097
rect 7539 5063 7573 5097
rect 7607 5063 7641 5097
rect 7675 5063 7709 5097
rect 7743 5063 7777 5097
rect 7811 5063 7845 5097
rect 555 2983 589 3017
rect 623 2983 657 3017
rect 691 2983 725 3017
rect 759 2983 793 3017
rect 827 2983 861 3017
rect 895 2983 929 3017
rect 963 2983 997 3017
rect 1031 2983 1065 3017
rect 1099 2983 1133 3017
rect 1167 2983 1201 3017
rect 1235 2983 1269 3017
rect 1303 2983 1337 3017
rect 1371 2983 1405 3017
rect 1439 2983 1473 3017
rect 1507 2983 1541 3017
rect 1575 2983 1609 3017
rect 1643 2983 1677 3017
rect 1711 2983 1745 3017
rect 1779 2983 1813 3017
rect 1847 2983 1881 3017
rect 1915 2983 1949 3017
rect 1983 2983 2017 3017
rect 2051 2983 2085 3017
rect 2475 2983 2509 3017
rect 2543 2983 2577 3017
rect 2611 2983 2645 3017
rect 2679 2983 2713 3017
rect 2747 2983 2781 3017
rect 2815 2983 2849 3017
rect 2883 2983 2917 3017
rect 2951 2983 2985 3017
rect 3019 2983 3053 3017
rect 3087 2983 3121 3017
rect 3155 2983 3189 3017
rect 3223 2983 3257 3017
rect 3291 2983 3325 3017
rect 3359 2983 3393 3017
rect 3427 2983 3461 3017
rect 3495 2983 3529 3017
rect 3563 2983 3597 3017
rect 3631 2983 3665 3017
rect 3699 2983 3733 3017
rect 3767 2983 3801 3017
rect 3835 2983 3869 3017
rect 3903 2983 3937 3017
rect 3971 2983 4005 3017
rect 4395 2983 4429 3017
rect 4463 2983 4497 3017
rect 4531 2983 4565 3017
rect 4599 2983 4633 3017
rect 4667 2983 4701 3017
rect 4735 2983 4769 3017
rect 4803 2983 4837 3017
rect 4871 2983 4905 3017
rect 4939 2983 4973 3017
rect 5007 2983 5041 3017
rect 5075 2983 5109 3017
rect 5143 2983 5177 3017
rect 5211 2983 5245 3017
rect 5279 2983 5313 3017
rect 5347 2983 5381 3017
rect 5415 2983 5449 3017
rect 5483 2983 5517 3017
rect 5551 2983 5585 3017
rect 5619 2983 5653 3017
rect 5687 2983 5721 3017
rect 5755 2983 5789 3017
rect 5823 2983 5857 3017
rect 5891 2983 5925 3017
rect 6315 2983 6349 3017
rect 6383 2983 6417 3017
rect 6451 2983 6485 3017
rect 6519 2983 6553 3017
rect 6587 2983 6621 3017
rect 6655 2983 6689 3017
rect 6723 2983 6757 3017
rect 6791 2983 6825 3017
rect 6859 2983 6893 3017
rect 6927 2983 6961 3017
rect 6995 2983 7029 3017
rect 7063 2983 7097 3017
rect 7131 2983 7165 3017
rect 7199 2983 7233 3017
rect 7267 2983 7301 3017
rect 7335 2983 7369 3017
rect 7403 2983 7437 3017
rect 7471 2983 7505 3017
rect 7539 2983 7573 3017
rect 7607 2983 7641 3017
rect 7675 2983 7709 3017
rect 7743 2983 7777 3017
rect 7811 2983 7845 3017
rect 555 1543 589 1577
rect 623 1543 657 1577
rect 691 1543 725 1577
rect 759 1543 793 1577
rect 827 1543 861 1577
rect 895 1543 929 1577
rect 963 1543 997 1577
rect 1031 1543 1065 1577
rect 1099 1543 1133 1577
rect 1167 1543 1201 1577
rect 1235 1543 1269 1577
rect 1303 1543 1337 1577
rect 1371 1543 1405 1577
rect 1439 1543 1473 1577
rect 1507 1543 1541 1577
rect 1575 1543 1609 1577
rect 1643 1543 1677 1577
rect 1711 1543 1745 1577
rect 1779 1543 1813 1577
rect 1847 1543 1881 1577
rect 1915 1543 1949 1577
rect 1983 1543 2017 1577
rect 2051 1543 2085 1577
rect 2475 1543 2509 1577
rect 2543 1543 2577 1577
rect 2611 1543 2645 1577
rect 2679 1543 2713 1577
rect 2747 1543 2781 1577
rect 2815 1543 2849 1577
rect 2883 1543 2917 1577
rect 2951 1543 2985 1577
rect 3019 1543 3053 1577
rect 3087 1543 3121 1577
rect 3155 1543 3189 1577
rect 3223 1543 3257 1577
rect 3291 1543 3325 1577
rect 3359 1543 3393 1577
rect 3427 1543 3461 1577
rect 3495 1543 3529 1577
rect 3563 1543 3597 1577
rect 3631 1543 3665 1577
rect 3699 1543 3733 1577
rect 3767 1543 3801 1577
rect 3835 1543 3869 1577
rect 3903 1543 3937 1577
rect 3971 1543 4005 1577
rect 4395 1543 4429 1577
rect 4463 1543 4497 1577
rect 4531 1543 4565 1577
rect 4599 1543 4633 1577
rect 4667 1543 4701 1577
rect 4735 1543 4769 1577
rect 4803 1543 4837 1577
rect 4871 1543 4905 1577
rect 4939 1543 4973 1577
rect 5007 1543 5041 1577
rect 5075 1543 5109 1577
rect 5143 1543 5177 1577
rect 5211 1543 5245 1577
rect 5279 1543 5313 1577
rect 5347 1543 5381 1577
rect 5415 1543 5449 1577
rect 5483 1543 5517 1577
rect 5551 1543 5585 1577
rect 5619 1543 5653 1577
rect 5687 1543 5721 1577
rect 5755 1543 5789 1577
rect 5823 1543 5857 1577
rect 5891 1543 5925 1577
rect 6315 1543 6349 1577
rect 6383 1543 6417 1577
rect 6451 1543 6485 1577
rect 6519 1543 6553 1577
rect 6587 1543 6621 1577
rect 6655 1543 6689 1577
rect 6723 1543 6757 1577
rect 6791 1543 6825 1577
rect 6859 1543 6893 1577
rect 6927 1543 6961 1577
rect 6995 1543 7029 1577
rect 7063 1543 7097 1577
rect 7131 1543 7165 1577
rect 7199 1543 7233 1577
rect 7267 1543 7301 1577
rect 7335 1543 7369 1577
rect 7403 1543 7437 1577
rect 7471 1543 7505 1577
rect 7539 1543 7573 1577
rect 7607 1543 7641 1577
rect 7675 1543 7709 1577
rect 7743 1543 7777 1577
rect 7811 1543 7845 1577
rect 555 423 589 457
rect 623 423 657 457
rect 691 423 725 457
rect 759 423 793 457
rect 827 423 861 457
rect 895 423 929 457
rect 963 423 997 457
rect 1031 423 1065 457
rect 1099 423 1133 457
rect 1167 423 1201 457
rect 1235 423 1269 457
rect 1303 423 1337 457
rect 1371 423 1405 457
rect 1439 423 1473 457
rect 1507 423 1541 457
rect 1575 423 1609 457
rect 1643 423 1677 457
rect 1711 423 1745 457
rect 1779 423 1813 457
rect 1847 423 1881 457
rect 1915 423 1949 457
rect 1983 423 2017 457
rect 2051 423 2085 457
rect 2475 423 2509 457
rect 2543 423 2577 457
rect 2611 423 2645 457
rect 2679 423 2713 457
rect 2747 423 2781 457
rect 2815 423 2849 457
rect 2883 423 2917 457
rect 2951 423 2985 457
rect 3019 423 3053 457
rect 3087 423 3121 457
rect 3155 423 3189 457
rect 3223 423 3257 457
rect 3291 423 3325 457
rect 3359 423 3393 457
rect 3427 423 3461 457
rect 3495 423 3529 457
rect 3563 423 3597 457
rect 3631 423 3665 457
rect 3699 423 3733 457
rect 3767 423 3801 457
rect 3835 423 3869 457
rect 3903 423 3937 457
rect 3971 423 4005 457
rect 4395 423 4429 457
rect 4463 423 4497 457
rect 4531 423 4565 457
rect 4599 423 4633 457
rect 4667 423 4701 457
rect 4735 423 4769 457
rect 4803 423 4837 457
rect 4871 423 4905 457
rect 4939 423 4973 457
rect 5007 423 5041 457
rect 5075 423 5109 457
rect 5143 423 5177 457
rect 5211 423 5245 457
rect 5279 423 5313 457
rect 5347 423 5381 457
rect 5415 423 5449 457
rect 5483 423 5517 457
rect 5551 423 5585 457
rect 5619 423 5653 457
rect 5687 423 5721 457
rect 5755 423 5789 457
rect 5823 423 5857 457
rect 5891 423 5925 457
rect 6315 423 6349 457
rect 6383 423 6417 457
rect 6451 423 6485 457
rect 6519 423 6553 457
rect 6587 423 6621 457
rect 6655 423 6689 457
rect 6723 423 6757 457
rect 6791 423 6825 457
rect 6859 423 6893 457
rect 6927 423 6961 457
rect 6995 423 7029 457
rect 7063 423 7097 457
rect 7131 423 7165 457
rect 7199 423 7233 457
rect 7267 423 7301 457
rect 7335 423 7369 457
rect 7403 423 7437 457
rect 7471 423 7505 457
rect 7539 423 7573 457
rect 7607 423 7641 457
rect 7675 423 7709 457
rect 7743 423 7777 457
rect 7811 423 7845 457
rect 555 -617 589 -583
rect 623 -617 657 -583
rect 691 -617 725 -583
rect 759 -617 793 -583
rect 827 -617 861 -583
rect 895 -617 929 -583
rect 963 -617 997 -583
rect 1031 -617 1065 -583
rect 1099 -617 1133 -583
rect 1167 -617 1201 -583
rect 1235 -617 1269 -583
rect 1303 -617 1337 -583
rect 1371 -617 1405 -583
rect 1439 -617 1473 -583
rect 1507 -617 1541 -583
rect 1575 -617 1609 -583
rect 1643 -617 1677 -583
rect 1711 -617 1745 -583
rect 1779 -617 1813 -583
rect 1847 -617 1881 -583
rect 1915 -617 1949 -583
rect 1983 -617 2017 -583
rect 2051 -617 2085 -583
rect 2475 -617 2509 -583
rect 2543 -617 2577 -583
rect 2611 -617 2645 -583
rect 2679 -617 2713 -583
rect 2747 -617 2781 -583
rect 2815 -617 2849 -583
rect 2883 -617 2917 -583
rect 2951 -617 2985 -583
rect 3019 -617 3053 -583
rect 3087 -617 3121 -583
rect 3155 -617 3189 -583
rect 3223 -617 3257 -583
rect 3291 -617 3325 -583
rect 3359 -617 3393 -583
rect 3427 -617 3461 -583
rect 3495 -617 3529 -583
rect 3563 -617 3597 -583
rect 3631 -617 3665 -583
rect 3699 -617 3733 -583
rect 3767 -617 3801 -583
rect 3835 -617 3869 -583
rect 3903 -617 3937 -583
rect 3971 -617 4005 -583
rect 4395 -617 4429 -583
rect 4463 -617 4497 -583
rect 4531 -617 4565 -583
rect 4599 -617 4633 -583
rect 4667 -617 4701 -583
rect 4735 -617 4769 -583
rect 4803 -617 4837 -583
rect 4871 -617 4905 -583
rect 4939 -617 4973 -583
rect 5007 -617 5041 -583
rect 5075 -617 5109 -583
rect 5143 -617 5177 -583
rect 5211 -617 5245 -583
rect 5279 -617 5313 -583
rect 5347 -617 5381 -583
rect 5415 -617 5449 -583
rect 5483 -617 5517 -583
rect 5551 -617 5585 -583
rect 5619 -617 5653 -583
rect 5687 -617 5721 -583
rect 5755 -617 5789 -583
rect 5823 -617 5857 -583
rect 5891 -617 5925 -583
rect 6315 -617 6349 -583
rect 6383 -617 6417 -583
rect 6451 -617 6485 -583
rect 6519 -617 6553 -583
rect 6587 -617 6621 -583
rect 6655 -617 6689 -583
rect 6723 -617 6757 -583
rect 6791 -617 6825 -583
rect 6859 -617 6893 -583
rect 6927 -617 6961 -583
rect 6995 -617 7029 -583
rect 7063 -617 7097 -583
rect 7131 -617 7165 -583
rect 7199 -617 7233 -583
rect 7267 -617 7301 -583
rect 7335 -617 7369 -583
rect 7403 -617 7437 -583
rect 7471 -617 7505 -583
rect 7539 -617 7573 -583
rect 7607 -617 7641 -583
rect 7675 -617 7709 -583
rect 7743 -617 7777 -583
rect 7811 -617 7845 -583
<< locali >>
rect 0 10057 8400 10080
rect 0 10023 137 10057
rect 171 10023 205 10057
rect 239 10023 273 10057
rect 307 10023 341 10057
rect 375 10023 409 10057
rect 443 10023 477 10057
rect 511 10023 545 10057
rect 579 10023 613 10057
rect 647 10023 681 10057
rect 715 10023 749 10057
rect 783 10023 817 10057
rect 851 10023 885 10057
rect 919 10023 953 10057
rect 987 10023 1021 10057
rect 1055 10023 1089 10057
rect 1123 10023 1157 10057
rect 1191 10023 1225 10057
rect 1259 10023 1293 10057
rect 1327 10023 1361 10057
rect 1395 10023 1429 10057
rect 1463 10023 1497 10057
rect 1531 10023 1565 10057
rect 1599 10023 1633 10057
rect 1667 10023 1701 10057
rect 1735 10023 1769 10057
rect 1803 10023 1837 10057
rect 1871 10023 1905 10057
rect 1939 10023 1973 10057
rect 2007 10023 2041 10057
rect 2075 10023 2109 10057
rect 2143 10023 2177 10057
rect 2211 10023 2245 10057
rect 2279 10023 2313 10057
rect 2347 10023 2381 10057
rect 2415 10023 2449 10057
rect 2483 10023 2517 10057
rect 2551 10023 2585 10057
rect 2619 10023 2653 10057
rect 2687 10023 2721 10057
rect 2755 10023 2789 10057
rect 2823 10023 2857 10057
rect 2891 10023 2925 10057
rect 2959 10023 2993 10057
rect 3027 10023 3061 10057
rect 3095 10023 3129 10057
rect 3163 10023 3197 10057
rect 3231 10023 3265 10057
rect 3299 10023 3333 10057
rect 3367 10023 3401 10057
rect 3435 10023 3469 10057
rect 3503 10023 3537 10057
rect 3571 10023 3605 10057
rect 3639 10023 3673 10057
rect 3707 10023 3741 10057
rect 3775 10023 3809 10057
rect 3843 10023 3877 10057
rect 3911 10023 3945 10057
rect 3979 10023 4013 10057
rect 4047 10023 4081 10057
rect 4115 10023 4149 10057
rect 4183 10023 4217 10057
rect 4251 10023 4285 10057
rect 4319 10023 4353 10057
rect 4387 10023 4421 10057
rect 4455 10023 4489 10057
rect 4523 10023 4557 10057
rect 4591 10023 4625 10057
rect 4659 10023 4693 10057
rect 4727 10023 4761 10057
rect 4795 10023 4829 10057
rect 4863 10023 4897 10057
rect 4931 10023 4965 10057
rect 4999 10023 5033 10057
rect 5067 10023 5101 10057
rect 5135 10023 5169 10057
rect 5203 10023 5237 10057
rect 5271 10023 5305 10057
rect 5339 10023 5373 10057
rect 5407 10023 5441 10057
rect 5475 10023 5509 10057
rect 5543 10023 5577 10057
rect 5611 10023 5645 10057
rect 5679 10023 5713 10057
rect 5747 10023 5781 10057
rect 5815 10023 5849 10057
rect 5883 10023 5917 10057
rect 5951 10023 5985 10057
rect 6019 10023 6053 10057
rect 6087 10023 6121 10057
rect 6155 10023 6189 10057
rect 6223 10023 6257 10057
rect 6291 10023 6325 10057
rect 6359 10023 6393 10057
rect 6427 10023 6461 10057
rect 6495 10023 6529 10057
rect 6563 10023 6597 10057
rect 6631 10023 6665 10057
rect 6699 10023 6733 10057
rect 6767 10023 6801 10057
rect 6835 10023 6869 10057
rect 6903 10023 6937 10057
rect 6971 10023 7005 10057
rect 7039 10023 7073 10057
rect 7107 10023 7141 10057
rect 7175 10023 7209 10057
rect 7243 10023 7277 10057
rect 7311 10023 7345 10057
rect 7379 10023 7413 10057
rect 7447 10023 7481 10057
rect 7515 10023 7549 10057
rect 7583 10023 7617 10057
rect 7651 10023 7685 10057
rect 7719 10023 7753 10057
rect 7787 10023 7821 10057
rect 7855 10023 7889 10057
rect 7923 10023 7957 10057
rect 7991 10023 8025 10057
rect 8059 10023 8093 10057
rect 8127 10023 8161 10057
rect 8195 10023 8229 10057
rect 8263 10023 8400 10057
rect 0 10000 8400 10023
rect 0 9927 80 10000
rect 0 9893 23 9927
rect 57 9893 80 9927
rect 8320 9927 8400 10000
rect 0 9859 80 9893
rect 0 9825 23 9859
rect 57 9825 80 9859
rect 0 9791 80 9825
rect 0 9757 23 9791
rect 57 9757 80 9791
rect 0 9723 80 9757
rect 0 9689 23 9723
rect 57 9689 80 9723
rect 0 9655 80 9689
rect 0 9621 23 9655
rect 57 9621 80 9655
rect 0 9587 80 9621
rect 0 9553 23 9587
rect 57 9553 80 9587
rect 0 9519 80 9553
rect 0 9485 23 9519
rect 57 9485 80 9519
rect 0 9451 80 9485
rect 0 9417 23 9451
rect 57 9417 80 9451
rect 0 9383 80 9417
rect 0 9349 23 9383
rect 57 9349 80 9383
rect 0 9315 80 9349
rect 0 9281 23 9315
rect 57 9281 80 9315
rect 0 9247 80 9281
rect 0 9213 23 9247
rect 57 9213 80 9247
rect 0 9179 80 9213
rect 0 9145 23 9179
rect 57 9145 80 9179
rect 0 9111 80 9145
rect 0 9077 23 9111
rect 57 9077 80 9111
rect 0 9043 80 9077
rect 0 9009 23 9043
rect 57 9009 80 9043
rect 0 8975 80 9009
rect 0 8941 23 8975
rect 57 8941 80 8975
rect 0 8907 80 8941
rect 0 8873 23 8907
rect 57 8873 80 8907
rect 160 9897 8240 9920
rect 160 9863 307 9897
rect 341 9863 375 9897
rect 409 9863 443 9897
rect 477 9863 511 9897
rect 545 9863 579 9897
rect 613 9863 647 9897
rect 681 9863 715 9897
rect 749 9863 783 9897
rect 817 9863 851 9897
rect 885 9863 919 9897
rect 953 9863 987 9897
rect 1021 9863 1055 9897
rect 1089 9863 1123 9897
rect 1157 9863 1191 9897
rect 1225 9863 1259 9897
rect 1293 9863 1327 9897
rect 1361 9863 1395 9897
rect 1429 9863 1463 9897
rect 1497 9863 1531 9897
rect 1565 9863 1599 9897
rect 1633 9863 1667 9897
rect 1701 9863 1735 9897
rect 1769 9863 1803 9897
rect 1837 9863 1871 9897
rect 1905 9863 1939 9897
rect 1973 9863 2007 9897
rect 2041 9863 2075 9897
rect 2109 9863 2143 9897
rect 2177 9863 2211 9897
rect 2245 9863 2279 9897
rect 2313 9863 2347 9897
rect 2381 9863 2415 9897
rect 2449 9863 2483 9897
rect 2517 9863 2551 9897
rect 2585 9863 2619 9897
rect 2653 9863 2687 9897
rect 2721 9863 2755 9897
rect 2789 9863 2823 9897
rect 2857 9863 2891 9897
rect 2925 9863 2959 9897
rect 2993 9863 3027 9897
rect 3061 9863 3095 9897
rect 3129 9863 3163 9897
rect 3197 9863 3231 9897
rect 3265 9863 3299 9897
rect 3333 9863 3367 9897
rect 3401 9863 3435 9897
rect 3469 9863 3503 9897
rect 3537 9863 3571 9897
rect 3605 9863 3639 9897
rect 3673 9863 3707 9897
rect 3741 9863 3775 9897
rect 3809 9863 3843 9897
rect 3877 9863 3911 9897
rect 3945 9863 3979 9897
rect 4013 9863 4047 9897
rect 4081 9863 4115 9897
rect 4149 9863 4183 9897
rect 4217 9863 4251 9897
rect 4285 9863 4319 9897
rect 4353 9863 4387 9897
rect 4421 9863 4455 9897
rect 4489 9863 4523 9897
rect 4557 9863 4591 9897
rect 4625 9863 4659 9897
rect 4693 9863 4727 9897
rect 4761 9863 4795 9897
rect 4829 9863 4863 9897
rect 4897 9863 4931 9897
rect 4965 9863 4999 9897
rect 5033 9863 5067 9897
rect 5101 9863 5135 9897
rect 5169 9863 5203 9897
rect 5237 9863 5271 9897
rect 5305 9863 5339 9897
rect 5373 9863 5407 9897
rect 5441 9863 5475 9897
rect 5509 9863 5543 9897
rect 5577 9863 5611 9897
rect 5645 9863 5679 9897
rect 5713 9863 5747 9897
rect 5781 9863 5815 9897
rect 5849 9863 5883 9897
rect 5917 9863 5951 9897
rect 5985 9863 6019 9897
rect 6053 9863 6087 9897
rect 6121 9863 6155 9897
rect 6189 9863 6223 9897
rect 6257 9863 6291 9897
rect 6325 9863 6359 9897
rect 6393 9863 6427 9897
rect 6461 9863 6495 9897
rect 6529 9863 6563 9897
rect 6597 9863 6631 9897
rect 6665 9863 6699 9897
rect 6733 9863 6767 9897
rect 6801 9863 6835 9897
rect 6869 9863 6903 9897
rect 6937 9863 6971 9897
rect 7005 9863 7039 9897
rect 7073 9863 7107 9897
rect 7141 9863 7175 9897
rect 7209 9863 7243 9897
rect 7277 9863 7311 9897
rect 7345 9863 7379 9897
rect 7413 9863 7447 9897
rect 7481 9863 7515 9897
rect 7549 9863 7583 9897
rect 7617 9863 7651 9897
rect 7685 9863 7719 9897
rect 7753 9863 7787 9897
rect 7821 9863 7855 9897
rect 7889 9863 7923 9897
rect 7957 9863 7991 9897
rect 8025 9863 8059 9897
rect 8093 9863 8240 9897
rect 160 9840 8240 9863
rect 160 9791 240 9840
rect 160 9757 183 9791
rect 217 9757 240 9791
rect 160 9723 240 9757
rect 160 9689 183 9723
rect 217 9689 240 9723
rect 160 9655 240 9689
rect 160 9621 183 9655
rect 217 9621 240 9655
rect 160 9587 240 9621
rect 160 9553 183 9587
rect 217 9553 240 9587
rect 160 9519 240 9553
rect 160 9485 183 9519
rect 217 9485 240 9519
rect 160 9451 240 9485
rect 160 9417 183 9451
rect 217 9417 240 9451
rect 160 9383 240 9417
rect 160 9349 183 9383
rect 217 9349 240 9383
rect 160 9315 240 9349
rect 160 9281 183 9315
rect 217 9281 240 9315
rect 160 9247 240 9281
rect 160 9213 183 9247
rect 217 9213 240 9247
rect 160 9179 240 9213
rect 160 9145 183 9179
rect 217 9145 240 9179
rect 320 9729 400 9840
rect 8160 9791 8240 9840
rect 320 9681 343 9729
rect 377 9681 400 9729
rect 320 9657 400 9681
rect 320 9613 343 9657
rect 377 9613 400 9657
rect 320 9585 400 9613
rect 320 9545 343 9585
rect 377 9545 400 9585
rect 320 9513 400 9545
rect 320 9477 343 9513
rect 377 9477 400 9513
rect 320 9443 400 9477
rect 320 9407 343 9443
rect 377 9407 400 9443
rect 320 9375 400 9407
rect 320 9335 343 9375
rect 377 9335 400 9375
rect 320 9307 400 9335
rect 320 9263 343 9307
rect 377 9263 400 9307
rect 320 9239 400 9263
rect 320 9191 343 9239
rect 377 9191 400 9239
rect 320 9160 400 9191
rect 2240 9729 2320 9760
rect 2240 9681 2263 9729
rect 2297 9681 2320 9729
rect 2240 9657 2320 9681
rect 2240 9613 2263 9657
rect 2297 9613 2320 9657
rect 2240 9585 2320 9613
rect 2240 9545 2263 9585
rect 2297 9545 2320 9585
rect 2240 9513 2320 9545
rect 2240 9477 2263 9513
rect 2297 9477 2320 9513
rect 2240 9443 2320 9477
rect 2240 9407 2263 9443
rect 2297 9407 2320 9443
rect 2240 9375 2320 9407
rect 2240 9335 2263 9375
rect 2297 9335 2320 9375
rect 2240 9307 2320 9335
rect 2240 9263 2263 9307
rect 2297 9263 2320 9307
rect 2240 9239 2320 9263
rect 2240 9191 2263 9239
rect 2297 9191 2320 9239
rect 2240 9160 2320 9191
rect 4160 9729 4240 9760
rect 4160 9681 4183 9729
rect 4217 9681 4240 9729
rect 4160 9657 4240 9681
rect 4160 9613 4183 9657
rect 4217 9613 4240 9657
rect 4160 9585 4240 9613
rect 4160 9545 4183 9585
rect 4217 9545 4240 9585
rect 4160 9513 4240 9545
rect 4160 9477 4183 9513
rect 4217 9477 4240 9513
rect 4160 9443 4240 9477
rect 4160 9407 4183 9443
rect 4217 9407 4240 9443
rect 4160 9375 4240 9407
rect 4160 9335 4183 9375
rect 4217 9335 4240 9375
rect 4160 9307 4240 9335
rect 4160 9263 4183 9307
rect 4217 9263 4240 9307
rect 4160 9239 4240 9263
rect 4160 9191 4183 9239
rect 4217 9191 4240 9239
rect 4160 9160 4240 9191
rect 6080 9729 6160 9760
rect 6080 9681 6103 9729
rect 6137 9681 6160 9729
rect 6080 9657 6160 9681
rect 6080 9613 6103 9657
rect 6137 9613 6160 9657
rect 6080 9585 6160 9613
rect 6080 9545 6103 9585
rect 6137 9545 6160 9585
rect 6080 9513 6160 9545
rect 6080 9477 6103 9513
rect 6137 9477 6160 9513
rect 6080 9443 6160 9477
rect 6080 9407 6103 9443
rect 6137 9407 6160 9443
rect 6080 9375 6160 9407
rect 6080 9335 6103 9375
rect 6137 9335 6160 9375
rect 6080 9307 6160 9335
rect 6080 9263 6103 9307
rect 6137 9263 6160 9307
rect 6080 9239 6160 9263
rect 6080 9191 6103 9239
rect 6137 9191 6160 9239
rect 6080 9160 6160 9191
rect 8000 9729 8080 9760
rect 8000 9681 8023 9729
rect 8057 9681 8080 9729
rect 8000 9657 8080 9681
rect 8000 9613 8023 9657
rect 8057 9613 8080 9657
rect 8000 9585 8080 9613
rect 8000 9545 8023 9585
rect 8057 9545 8080 9585
rect 8000 9513 8080 9545
rect 8000 9477 8023 9513
rect 8057 9477 8080 9513
rect 8000 9443 8080 9477
rect 8000 9407 8023 9443
rect 8057 9407 8080 9443
rect 8000 9375 8080 9407
rect 8000 9335 8023 9375
rect 8057 9335 8080 9375
rect 8000 9307 8080 9335
rect 8000 9263 8023 9307
rect 8057 9263 8080 9307
rect 8000 9239 8080 9263
rect 8000 9191 8023 9239
rect 8057 9191 8080 9239
rect 8000 9160 8080 9191
rect 8160 9757 8183 9791
rect 8217 9757 8240 9791
rect 8160 9723 8240 9757
rect 8160 9689 8183 9723
rect 8217 9689 8240 9723
rect 8160 9655 8240 9689
rect 8160 9621 8183 9655
rect 8217 9621 8240 9655
rect 8160 9587 8240 9621
rect 8160 9553 8183 9587
rect 8217 9553 8240 9587
rect 8160 9519 8240 9553
rect 8160 9485 8183 9519
rect 8217 9485 8240 9519
rect 8160 9451 8240 9485
rect 8160 9417 8183 9451
rect 8217 9417 8240 9451
rect 8160 9383 8240 9417
rect 8160 9349 8183 9383
rect 8217 9349 8240 9383
rect 8160 9315 8240 9349
rect 8160 9281 8183 9315
rect 8217 9281 8240 9315
rect 8160 9247 8240 9281
rect 8160 9213 8183 9247
rect 8217 9213 8240 9247
rect 8160 9179 8240 9213
rect 160 9111 240 9145
rect 8160 9145 8183 9179
rect 8217 9145 8240 9179
rect 160 9077 183 9111
rect 217 9077 240 9111
rect 160 9043 240 9077
rect 160 9009 183 9043
rect 217 9009 240 9043
rect 520 9097 2120 9120
rect 520 9063 547 9097
rect 589 9063 619 9097
rect 657 9063 691 9097
rect 725 9063 759 9097
rect 797 9063 827 9097
rect 869 9063 895 9097
rect 941 9063 963 9097
rect 1013 9063 1031 9097
rect 1085 9063 1099 9097
rect 1157 9063 1167 9097
rect 1229 9063 1235 9097
rect 1301 9063 1303 9097
rect 1337 9063 1339 9097
rect 1405 9063 1411 9097
rect 1473 9063 1483 9097
rect 1541 9063 1555 9097
rect 1609 9063 1627 9097
rect 1677 9063 1699 9097
rect 1745 9063 1771 9097
rect 1813 9063 1843 9097
rect 1881 9063 1915 9097
rect 1949 9063 1983 9097
rect 2021 9063 2051 9097
rect 2093 9063 2120 9097
rect 520 9040 2120 9063
rect 2440 9097 4040 9120
rect 2440 9063 2467 9097
rect 2509 9063 2539 9097
rect 2577 9063 2611 9097
rect 2645 9063 2679 9097
rect 2717 9063 2747 9097
rect 2789 9063 2815 9097
rect 2861 9063 2883 9097
rect 2933 9063 2951 9097
rect 3005 9063 3019 9097
rect 3077 9063 3087 9097
rect 3149 9063 3155 9097
rect 3221 9063 3223 9097
rect 3257 9063 3259 9097
rect 3325 9063 3331 9097
rect 3393 9063 3403 9097
rect 3461 9063 3475 9097
rect 3529 9063 3547 9097
rect 3597 9063 3619 9097
rect 3665 9063 3691 9097
rect 3733 9063 3763 9097
rect 3801 9063 3835 9097
rect 3869 9063 3903 9097
rect 3941 9063 3971 9097
rect 4013 9063 4040 9097
rect 2440 9040 4040 9063
rect 4360 9097 5960 9120
rect 4360 9063 4387 9097
rect 4429 9063 4459 9097
rect 4497 9063 4531 9097
rect 4565 9063 4599 9097
rect 4637 9063 4667 9097
rect 4709 9063 4735 9097
rect 4781 9063 4803 9097
rect 4853 9063 4871 9097
rect 4925 9063 4939 9097
rect 4997 9063 5007 9097
rect 5069 9063 5075 9097
rect 5141 9063 5143 9097
rect 5177 9063 5179 9097
rect 5245 9063 5251 9097
rect 5313 9063 5323 9097
rect 5381 9063 5395 9097
rect 5449 9063 5467 9097
rect 5517 9063 5539 9097
rect 5585 9063 5611 9097
rect 5653 9063 5683 9097
rect 5721 9063 5755 9097
rect 5789 9063 5823 9097
rect 5861 9063 5891 9097
rect 5933 9063 5960 9097
rect 4360 9040 5960 9063
rect 6280 9097 7880 9120
rect 6280 9063 6307 9097
rect 6349 9063 6379 9097
rect 6417 9063 6451 9097
rect 6485 9063 6519 9097
rect 6557 9063 6587 9097
rect 6629 9063 6655 9097
rect 6701 9063 6723 9097
rect 6773 9063 6791 9097
rect 6845 9063 6859 9097
rect 6917 9063 6927 9097
rect 6989 9063 6995 9097
rect 7061 9063 7063 9097
rect 7097 9063 7099 9097
rect 7165 9063 7171 9097
rect 7233 9063 7243 9097
rect 7301 9063 7315 9097
rect 7369 9063 7387 9097
rect 7437 9063 7459 9097
rect 7505 9063 7531 9097
rect 7573 9063 7603 9097
rect 7641 9063 7675 9097
rect 7709 9063 7743 9097
rect 7781 9063 7811 9097
rect 7853 9063 7880 9097
rect 6280 9040 7880 9063
rect 8160 9111 8240 9145
rect 8160 9077 8183 9111
rect 8217 9077 8240 9111
rect 8160 9043 8240 9077
rect 160 8960 240 9009
rect 8160 9009 8183 9043
rect 8217 9009 8240 9043
rect 8160 8960 8240 9009
rect 160 8937 8240 8960
rect 160 8903 307 8937
rect 341 8903 375 8937
rect 409 8903 443 8937
rect 477 8903 511 8937
rect 545 8903 579 8937
rect 613 8903 647 8937
rect 681 8903 715 8937
rect 749 8903 783 8937
rect 817 8903 851 8937
rect 885 8903 919 8937
rect 953 8903 987 8937
rect 1021 8903 1055 8937
rect 1089 8903 1123 8937
rect 1157 8903 1191 8937
rect 1225 8903 1259 8937
rect 1293 8903 1327 8937
rect 1361 8903 1395 8937
rect 1429 8903 1463 8937
rect 1497 8903 1531 8937
rect 1565 8903 1599 8937
rect 1633 8903 1667 8937
rect 1701 8903 1735 8937
rect 1769 8903 1803 8937
rect 1837 8903 1871 8937
rect 1905 8903 1939 8937
rect 1973 8903 2007 8937
rect 2041 8903 2075 8937
rect 2109 8903 2143 8937
rect 2177 8903 2211 8937
rect 2245 8903 2279 8937
rect 2313 8903 2347 8937
rect 2381 8903 2415 8937
rect 2449 8903 2483 8937
rect 2517 8903 2551 8937
rect 2585 8903 2619 8937
rect 2653 8903 2687 8937
rect 2721 8903 2755 8937
rect 2789 8903 2823 8937
rect 2857 8903 2891 8937
rect 2925 8903 2959 8937
rect 2993 8903 3027 8937
rect 3061 8903 3095 8937
rect 3129 8903 3163 8937
rect 3197 8903 3231 8937
rect 3265 8903 3299 8937
rect 3333 8903 3367 8937
rect 3401 8903 3435 8937
rect 3469 8903 3503 8937
rect 3537 8903 3571 8937
rect 3605 8903 3639 8937
rect 3673 8903 3707 8937
rect 3741 8903 3775 8937
rect 3809 8903 3843 8937
rect 3877 8903 3911 8937
rect 3945 8903 3979 8937
rect 4013 8903 4047 8937
rect 4081 8903 4115 8937
rect 4149 8903 4183 8937
rect 4217 8903 4251 8937
rect 4285 8903 4319 8937
rect 4353 8903 4387 8937
rect 4421 8903 4455 8937
rect 4489 8903 4523 8937
rect 4557 8903 4591 8937
rect 4625 8903 4659 8937
rect 4693 8903 4727 8937
rect 4761 8903 4795 8937
rect 4829 8903 4863 8937
rect 4897 8903 4931 8937
rect 4965 8903 4999 8937
rect 5033 8903 5067 8937
rect 5101 8903 5135 8937
rect 5169 8903 5203 8937
rect 5237 8903 5271 8937
rect 5305 8903 5339 8937
rect 5373 8903 5407 8937
rect 5441 8903 5475 8937
rect 5509 8903 5543 8937
rect 5577 8903 5611 8937
rect 5645 8903 5679 8937
rect 5713 8903 5747 8937
rect 5781 8903 5815 8937
rect 5849 8903 5883 8937
rect 5917 8903 5951 8937
rect 5985 8903 6019 8937
rect 6053 8903 6087 8937
rect 6121 8903 6155 8937
rect 6189 8903 6223 8937
rect 6257 8903 6291 8937
rect 6325 8903 6359 8937
rect 6393 8903 6427 8937
rect 6461 8903 6495 8937
rect 6529 8903 6563 8937
rect 6597 8903 6631 8937
rect 6665 8903 6699 8937
rect 6733 8903 6767 8937
rect 6801 8903 6835 8937
rect 6869 8903 6903 8937
rect 6937 8903 6971 8937
rect 7005 8903 7039 8937
rect 7073 8903 7107 8937
rect 7141 8903 7175 8937
rect 7209 8903 7243 8937
rect 7277 8903 7311 8937
rect 7345 8903 7379 8937
rect 7413 8903 7447 8937
rect 7481 8903 7515 8937
rect 7549 8903 7583 8937
rect 7617 8903 7651 8937
rect 7685 8903 7719 8937
rect 7753 8903 7787 8937
rect 7821 8903 7855 8937
rect 7889 8903 7923 8937
rect 7957 8903 7991 8937
rect 8025 8903 8059 8937
rect 8093 8903 8240 8937
rect 160 8880 8240 8903
rect 8320 9893 8343 9927
rect 8377 9893 8400 9927
rect 8320 9859 8400 9893
rect 8320 9825 8343 9859
rect 8377 9825 8400 9859
rect 8320 9791 8400 9825
rect 8320 9757 8343 9791
rect 8377 9757 8400 9791
rect 8320 9723 8400 9757
rect 8320 9689 8343 9723
rect 8377 9689 8400 9723
rect 8320 9655 8400 9689
rect 8320 9621 8343 9655
rect 8377 9621 8400 9655
rect 8320 9587 8400 9621
rect 8320 9553 8343 9587
rect 8377 9553 8400 9587
rect 8320 9519 8400 9553
rect 8320 9485 8343 9519
rect 8377 9485 8400 9519
rect 8320 9451 8400 9485
rect 8320 9417 8343 9451
rect 8377 9417 8400 9451
rect 8320 9383 8400 9417
rect 8320 9349 8343 9383
rect 8377 9349 8400 9383
rect 8320 9315 8400 9349
rect 8320 9281 8343 9315
rect 8377 9281 8400 9315
rect 8320 9247 8400 9281
rect 8320 9213 8343 9247
rect 8377 9213 8400 9247
rect 8320 9179 8400 9213
rect 8320 9145 8343 9179
rect 8377 9145 8400 9179
rect 8320 9111 8400 9145
rect 8320 9077 8343 9111
rect 8377 9077 8400 9111
rect 8320 9043 8400 9077
rect 8320 9009 8343 9043
rect 8377 9009 8400 9043
rect 8320 8975 8400 9009
rect 8320 8941 8343 8975
rect 8377 8941 8400 8975
rect 8320 8907 8400 8941
rect 0 8800 80 8873
rect 8320 8873 8343 8907
rect 8377 8873 8400 8907
rect 8320 8800 8400 8873
rect 0 8777 8400 8800
rect 0 8743 137 8777
rect 171 8743 205 8777
rect 239 8743 273 8777
rect 307 8743 341 8777
rect 375 8743 409 8777
rect 443 8743 477 8777
rect 511 8743 545 8777
rect 579 8743 613 8777
rect 647 8743 681 8777
rect 715 8743 749 8777
rect 783 8743 817 8777
rect 851 8743 885 8777
rect 919 8743 953 8777
rect 987 8743 1021 8777
rect 1055 8743 1089 8777
rect 1123 8743 1157 8777
rect 1191 8743 1225 8777
rect 1259 8743 1293 8777
rect 1327 8743 1361 8777
rect 1395 8743 1429 8777
rect 1463 8743 1497 8777
rect 1531 8743 1565 8777
rect 1599 8743 1633 8777
rect 1667 8743 1701 8777
rect 1735 8743 1769 8777
rect 1803 8743 1837 8777
rect 1871 8743 1905 8777
rect 1939 8743 1973 8777
rect 2007 8743 2041 8777
rect 2075 8743 2109 8777
rect 2143 8743 2177 8777
rect 2211 8743 2245 8777
rect 2279 8743 2313 8777
rect 2347 8743 2381 8777
rect 2415 8743 2449 8777
rect 2483 8743 2517 8777
rect 2551 8743 2585 8777
rect 2619 8743 2653 8777
rect 2687 8743 2721 8777
rect 2755 8743 2789 8777
rect 2823 8743 2857 8777
rect 2891 8743 2925 8777
rect 2959 8743 2993 8777
rect 3027 8743 3061 8777
rect 3095 8743 3129 8777
rect 3163 8743 3197 8777
rect 3231 8743 3265 8777
rect 3299 8743 3333 8777
rect 3367 8743 3401 8777
rect 3435 8743 3469 8777
rect 3503 8743 3537 8777
rect 3571 8743 3605 8777
rect 3639 8743 3673 8777
rect 3707 8743 3741 8777
rect 3775 8743 3809 8777
rect 3843 8743 3877 8777
rect 3911 8743 3945 8777
rect 3979 8743 4013 8777
rect 4047 8743 4081 8777
rect 4115 8743 4149 8777
rect 4183 8743 4217 8777
rect 4251 8743 4285 8777
rect 4319 8743 4353 8777
rect 4387 8743 4421 8777
rect 4455 8743 4489 8777
rect 4523 8743 4557 8777
rect 4591 8743 4625 8777
rect 4659 8743 4693 8777
rect 4727 8743 4761 8777
rect 4795 8743 4829 8777
rect 4863 8743 4897 8777
rect 4931 8743 4965 8777
rect 4999 8743 5033 8777
rect 5067 8743 5101 8777
rect 5135 8743 5169 8777
rect 5203 8743 5237 8777
rect 5271 8743 5305 8777
rect 5339 8743 5373 8777
rect 5407 8743 5441 8777
rect 5475 8743 5509 8777
rect 5543 8743 5577 8777
rect 5611 8743 5645 8777
rect 5679 8743 5713 8777
rect 5747 8743 5781 8777
rect 5815 8743 5849 8777
rect 5883 8743 5917 8777
rect 5951 8743 5985 8777
rect 6019 8743 6053 8777
rect 6087 8743 6121 8777
rect 6155 8743 6189 8777
rect 6223 8743 6257 8777
rect 6291 8743 6325 8777
rect 6359 8743 6393 8777
rect 6427 8743 6461 8777
rect 6495 8743 6529 8777
rect 6563 8743 6597 8777
rect 6631 8743 6665 8777
rect 6699 8743 6733 8777
rect 6767 8743 6801 8777
rect 6835 8743 6869 8777
rect 6903 8743 6937 8777
rect 6971 8743 7005 8777
rect 7039 8743 7073 8777
rect 7107 8743 7141 8777
rect 7175 8743 7209 8777
rect 7243 8743 7277 8777
rect 7311 8743 7345 8777
rect 7379 8743 7413 8777
rect 7447 8743 7481 8777
rect 7515 8743 7549 8777
rect 7583 8743 7617 8777
rect 7651 8743 7685 8777
rect 7719 8743 7753 8777
rect 7787 8743 7821 8777
rect 7855 8743 7889 8777
rect 7923 8743 7957 8777
rect 7991 8743 8025 8777
rect 8059 8743 8093 8777
rect 8127 8743 8161 8777
rect 8195 8743 8229 8777
rect 8263 8743 8400 8777
rect 0 8720 8400 8743
rect 0 8000 80 8720
rect 160 8457 8240 8640
rect 160 8423 183 8457
rect 217 8423 8183 8457
rect 8217 8423 8240 8457
rect 160 8400 8240 8423
rect 160 8297 8240 8320
rect 160 8263 183 8297
rect 217 8263 8183 8297
rect 8217 8263 8240 8297
rect 160 8080 8240 8263
rect 8320 8000 8400 8720
rect 0 7977 8400 8000
rect 0 7943 137 7977
rect 171 7943 205 7977
rect 239 7943 273 7977
rect 307 7943 341 7977
rect 375 7943 409 7977
rect 443 7943 477 7977
rect 511 7943 545 7977
rect 579 7943 613 7977
rect 647 7943 681 7977
rect 715 7943 749 7977
rect 783 7943 817 7977
rect 851 7943 885 7977
rect 919 7943 953 7977
rect 987 7943 1021 7977
rect 1055 7943 1089 7977
rect 1123 7943 1157 7977
rect 1191 7943 1225 7977
rect 1259 7943 1293 7977
rect 1327 7943 1361 7977
rect 1395 7943 1429 7977
rect 1463 7943 1497 7977
rect 1531 7943 1565 7977
rect 1599 7943 1633 7977
rect 1667 7943 1701 7977
rect 1735 7943 1769 7977
rect 1803 7943 1837 7977
rect 1871 7943 1905 7977
rect 1939 7943 1973 7977
rect 2007 7943 2041 7977
rect 2075 7943 2109 7977
rect 2143 7943 2177 7977
rect 2211 7943 2245 7977
rect 2279 7943 2313 7977
rect 2347 7943 2381 7977
rect 2415 7943 2449 7977
rect 2483 7943 2517 7977
rect 2551 7943 2585 7977
rect 2619 7943 2653 7977
rect 2687 7943 2721 7977
rect 2755 7943 2789 7977
rect 2823 7943 2857 7977
rect 2891 7943 2925 7977
rect 2959 7943 2993 7977
rect 3027 7943 3061 7977
rect 3095 7943 3129 7977
rect 3163 7943 3197 7977
rect 3231 7943 3265 7977
rect 3299 7943 3333 7977
rect 3367 7943 3401 7977
rect 3435 7943 3469 7977
rect 3503 7943 3537 7977
rect 3571 7943 3605 7977
rect 3639 7943 3673 7977
rect 3707 7943 3741 7977
rect 3775 7943 3809 7977
rect 3843 7943 3877 7977
rect 3911 7943 3945 7977
rect 3979 7943 4013 7977
rect 4047 7943 4081 7977
rect 4115 7943 4149 7977
rect 4183 7943 4217 7977
rect 4251 7943 4285 7977
rect 4319 7943 4353 7977
rect 4387 7943 4421 7977
rect 4455 7943 4489 7977
rect 4523 7943 4557 7977
rect 4591 7943 4625 7977
rect 4659 7943 4693 7977
rect 4727 7943 4761 7977
rect 4795 7943 4829 7977
rect 4863 7943 4897 7977
rect 4931 7943 4965 7977
rect 4999 7943 5033 7977
rect 5067 7943 5101 7977
rect 5135 7943 5169 7977
rect 5203 7943 5237 7977
rect 5271 7943 5305 7977
rect 5339 7943 5373 7977
rect 5407 7943 5441 7977
rect 5475 7943 5509 7977
rect 5543 7943 5577 7977
rect 5611 7943 5645 7977
rect 5679 7943 5713 7977
rect 5747 7943 5781 7977
rect 5815 7943 5849 7977
rect 5883 7943 5917 7977
rect 5951 7943 5985 7977
rect 6019 7943 6053 7977
rect 6087 7943 6121 7977
rect 6155 7943 6189 7977
rect 6223 7943 6257 7977
rect 6291 7943 6325 7977
rect 6359 7943 6393 7977
rect 6427 7943 6461 7977
rect 6495 7943 6529 7977
rect 6563 7943 6597 7977
rect 6631 7943 6665 7977
rect 6699 7943 6733 7977
rect 6767 7943 6801 7977
rect 6835 7943 6869 7977
rect 6903 7943 6937 7977
rect 6971 7943 7005 7977
rect 7039 7943 7073 7977
rect 7107 7943 7141 7977
rect 7175 7943 7209 7977
rect 7243 7943 7277 7977
rect 7311 7943 7345 7977
rect 7379 7943 7413 7977
rect 7447 7943 7481 7977
rect 7515 7943 7549 7977
rect 7583 7943 7617 7977
rect 7651 7943 7685 7977
rect 7719 7943 7753 7977
rect 7787 7943 7821 7977
rect 7855 7943 7889 7977
rect 7923 7943 7957 7977
rect 7991 7943 8025 7977
rect 8059 7943 8093 7977
rect 8127 7943 8161 7977
rect 8195 7943 8229 7977
rect 8263 7943 8400 7977
rect 0 7920 8400 7943
rect 0 7867 80 7920
rect 0 7833 23 7867
rect 57 7833 80 7867
rect 0 7799 80 7833
rect 0 7765 23 7799
rect 57 7765 80 7799
rect 0 7731 80 7765
rect 520 7817 2120 7840
rect 520 7783 547 7817
rect 589 7783 619 7817
rect 657 7783 691 7817
rect 725 7783 759 7817
rect 797 7783 827 7817
rect 869 7783 895 7817
rect 941 7783 963 7817
rect 1013 7783 1031 7817
rect 1085 7783 1099 7817
rect 1157 7783 1167 7817
rect 1229 7783 1235 7817
rect 1301 7783 1303 7817
rect 1337 7783 1339 7817
rect 1405 7783 1411 7817
rect 1473 7783 1483 7817
rect 1541 7783 1555 7817
rect 1609 7783 1627 7817
rect 1677 7783 1699 7817
rect 1745 7783 1771 7817
rect 1813 7783 1843 7817
rect 1881 7783 1915 7817
rect 1949 7783 1983 7817
rect 2021 7783 2051 7817
rect 2093 7783 2120 7817
rect 520 7760 2120 7783
rect 2440 7817 4040 7840
rect 2440 7783 2467 7817
rect 2509 7783 2539 7817
rect 2577 7783 2611 7817
rect 2645 7783 2679 7817
rect 2717 7783 2747 7817
rect 2789 7783 2815 7817
rect 2861 7783 2883 7817
rect 2933 7783 2951 7817
rect 3005 7783 3019 7817
rect 3077 7783 3087 7817
rect 3149 7783 3155 7817
rect 3221 7783 3223 7817
rect 3257 7783 3259 7817
rect 3325 7783 3331 7817
rect 3393 7783 3403 7817
rect 3461 7783 3475 7817
rect 3529 7783 3547 7817
rect 3597 7783 3619 7817
rect 3665 7783 3691 7817
rect 3733 7783 3763 7817
rect 3801 7783 3835 7817
rect 3869 7783 3903 7817
rect 3941 7783 3971 7817
rect 4013 7783 4040 7817
rect 2440 7760 4040 7783
rect 4360 7817 5960 7840
rect 4360 7783 4387 7817
rect 4429 7783 4459 7817
rect 4497 7783 4531 7817
rect 4565 7783 4599 7817
rect 4637 7783 4667 7817
rect 4709 7783 4735 7817
rect 4781 7783 4803 7817
rect 4853 7783 4871 7817
rect 4925 7783 4939 7817
rect 4997 7783 5007 7817
rect 5069 7783 5075 7817
rect 5141 7783 5143 7817
rect 5177 7783 5179 7817
rect 5245 7783 5251 7817
rect 5313 7783 5323 7817
rect 5381 7783 5395 7817
rect 5449 7783 5467 7817
rect 5517 7783 5539 7817
rect 5585 7783 5611 7817
rect 5653 7783 5683 7817
rect 5721 7783 5755 7817
rect 5789 7783 5823 7817
rect 5861 7783 5891 7817
rect 5933 7783 5960 7817
rect 4360 7760 5960 7783
rect 6280 7817 7880 7840
rect 6280 7783 6307 7817
rect 6349 7783 6379 7817
rect 6417 7783 6451 7817
rect 6485 7783 6519 7817
rect 6557 7783 6587 7817
rect 6629 7783 6655 7817
rect 6701 7783 6723 7817
rect 6773 7783 6791 7817
rect 6845 7783 6859 7817
rect 6917 7783 6927 7817
rect 6989 7783 6995 7817
rect 7061 7783 7063 7817
rect 7097 7783 7099 7817
rect 7165 7783 7171 7817
rect 7233 7783 7243 7817
rect 7301 7783 7315 7817
rect 7369 7783 7387 7817
rect 7437 7783 7459 7817
rect 7505 7783 7531 7817
rect 7573 7783 7603 7817
rect 7641 7783 7675 7817
rect 7709 7783 7743 7817
rect 7781 7783 7811 7817
rect 7853 7783 7880 7817
rect 6280 7760 7880 7783
rect 0 7697 23 7731
rect 57 7697 80 7731
rect 0 7663 80 7697
rect 0 7629 23 7663
rect 57 7629 80 7663
rect 0 7595 80 7629
rect 0 7561 23 7595
rect 57 7561 80 7595
rect 0 7527 80 7561
rect 0 7493 23 7527
rect 57 7493 80 7527
rect 0 7440 80 7493
rect 320 7673 400 7720
rect 320 7637 343 7673
rect 377 7637 400 7673
rect 320 7603 400 7637
rect 320 7567 343 7603
rect 377 7567 400 7603
rect 320 7440 400 7567
rect 2240 7673 2320 7720
rect 2240 7637 2263 7673
rect 2297 7637 2320 7673
rect 2240 7603 2320 7637
rect 2240 7567 2263 7603
rect 2297 7567 2320 7603
rect 2240 7520 2320 7567
rect 4160 7673 4240 7720
rect 4160 7637 4183 7673
rect 4217 7637 4240 7673
rect 4160 7603 4240 7637
rect 4160 7567 4183 7603
rect 4217 7567 4240 7603
rect 4160 7520 4240 7567
rect 6080 7673 6160 7720
rect 6080 7637 6103 7673
rect 6137 7637 6160 7673
rect 6080 7603 6160 7637
rect 6080 7567 6103 7603
rect 6137 7567 6160 7603
rect 6080 7520 6160 7567
rect 8000 7673 8080 7720
rect 8000 7637 8023 7673
rect 8057 7637 8080 7673
rect 8000 7603 8080 7637
rect 8000 7567 8023 7603
rect 8057 7567 8080 7603
rect 8000 7520 8080 7567
rect 8320 7440 8400 7920
rect 0 7417 8400 7440
rect 0 7383 137 7417
rect 171 7383 205 7417
rect 239 7383 273 7417
rect 307 7383 341 7417
rect 375 7383 409 7417
rect 443 7383 477 7417
rect 511 7383 545 7417
rect 579 7383 613 7417
rect 647 7383 681 7417
rect 715 7383 749 7417
rect 783 7383 817 7417
rect 851 7383 885 7417
rect 919 7383 953 7417
rect 987 7383 1021 7417
rect 1055 7383 1089 7417
rect 1123 7383 1157 7417
rect 1191 7383 1225 7417
rect 1259 7383 1293 7417
rect 1327 7383 1361 7417
rect 1395 7383 1429 7417
rect 1463 7383 1497 7417
rect 1531 7383 1565 7417
rect 1599 7383 1633 7417
rect 1667 7383 1701 7417
rect 1735 7383 1769 7417
rect 1803 7383 1837 7417
rect 1871 7383 1905 7417
rect 1939 7383 1973 7417
rect 2007 7383 2041 7417
rect 2075 7383 2109 7417
rect 2143 7383 2177 7417
rect 2211 7383 2245 7417
rect 2279 7383 2313 7417
rect 2347 7383 2381 7417
rect 2415 7383 2449 7417
rect 2483 7383 2517 7417
rect 2551 7383 2585 7417
rect 2619 7383 2653 7417
rect 2687 7383 2721 7417
rect 2755 7383 2789 7417
rect 2823 7383 2857 7417
rect 2891 7383 2925 7417
rect 2959 7383 2993 7417
rect 3027 7383 3061 7417
rect 3095 7383 3129 7417
rect 3163 7383 3197 7417
rect 3231 7383 3265 7417
rect 3299 7383 3333 7417
rect 3367 7383 3401 7417
rect 3435 7383 3469 7417
rect 3503 7383 3537 7417
rect 3571 7383 3605 7417
rect 3639 7383 3673 7417
rect 3707 7383 3741 7417
rect 3775 7383 3809 7417
rect 3843 7383 3877 7417
rect 3911 7383 3945 7417
rect 3979 7383 4013 7417
rect 4047 7383 4081 7417
rect 4115 7383 4149 7417
rect 4183 7383 4217 7417
rect 4251 7383 4285 7417
rect 4319 7383 4353 7417
rect 4387 7383 4421 7417
rect 4455 7383 4489 7417
rect 4523 7383 4557 7417
rect 4591 7383 4625 7417
rect 4659 7383 4693 7417
rect 4727 7383 4761 7417
rect 4795 7383 4829 7417
rect 4863 7383 4897 7417
rect 4931 7383 4965 7417
rect 4999 7383 5033 7417
rect 5067 7383 5101 7417
rect 5135 7383 5169 7417
rect 5203 7383 5237 7417
rect 5271 7383 5305 7417
rect 5339 7383 5373 7417
rect 5407 7383 5441 7417
rect 5475 7383 5509 7417
rect 5543 7383 5577 7417
rect 5611 7383 5645 7417
rect 5679 7383 5713 7417
rect 5747 7383 5781 7417
rect 5815 7383 5849 7417
rect 5883 7383 5917 7417
rect 5951 7383 5985 7417
rect 6019 7383 6053 7417
rect 6087 7383 6121 7417
rect 6155 7383 6189 7417
rect 6223 7383 6257 7417
rect 6291 7383 6325 7417
rect 6359 7383 6393 7417
rect 6427 7383 6461 7417
rect 6495 7383 6529 7417
rect 6563 7383 6597 7417
rect 6631 7383 6665 7417
rect 6699 7383 6733 7417
rect 6767 7383 6801 7417
rect 6835 7383 6869 7417
rect 6903 7383 6937 7417
rect 6971 7383 7005 7417
rect 7039 7383 7073 7417
rect 7107 7383 7141 7417
rect 7175 7383 7209 7417
rect 7243 7383 7277 7417
rect 7311 7383 7345 7417
rect 7379 7383 7413 7417
rect 7447 7383 7481 7417
rect 7515 7383 7549 7417
rect 7583 7383 7617 7417
rect 7651 7383 7685 7417
rect 7719 7383 7753 7417
rect 7787 7383 7821 7417
rect 7855 7383 7889 7417
rect 7923 7383 7957 7417
rect 7991 7383 8025 7417
rect 8059 7383 8093 7417
rect 8127 7383 8161 7417
rect 8195 7383 8229 7417
rect 8263 7383 8400 7417
rect 0 7360 8400 7383
rect 0 7280 80 7360
rect 8320 7280 8400 7360
rect 0 7257 8400 7280
rect 0 7223 137 7257
rect 171 7223 205 7257
rect 239 7223 273 7257
rect 307 7223 341 7257
rect 375 7223 409 7257
rect 443 7223 477 7257
rect 511 7223 545 7257
rect 579 7223 613 7257
rect 647 7223 681 7257
rect 715 7223 749 7257
rect 783 7223 817 7257
rect 851 7223 885 7257
rect 919 7223 953 7257
rect 987 7223 1021 7257
rect 1055 7223 1089 7257
rect 1123 7223 1157 7257
rect 1191 7223 1225 7257
rect 1259 7223 1293 7257
rect 1327 7223 1361 7257
rect 1395 7223 1429 7257
rect 1463 7223 1497 7257
rect 1531 7223 1565 7257
rect 1599 7223 1633 7257
rect 1667 7223 1701 7257
rect 1735 7223 1769 7257
rect 1803 7223 1837 7257
rect 1871 7223 1905 7257
rect 1939 7223 1973 7257
rect 2007 7223 2041 7257
rect 2075 7223 2109 7257
rect 2143 7223 2177 7257
rect 2211 7223 2245 7257
rect 2279 7223 2313 7257
rect 2347 7223 2381 7257
rect 2415 7223 2449 7257
rect 2483 7223 2517 7257
rect 2551 7223 2585 7257
rect 2619 7223 2653 7257
rect 2687 7223 2721 7257
rect 2755 7223 2789 7257
rect 2823 7223 2857 7257
rect 2891 7223 2925 7257
rect 2959 7223 2993 7257
rect 3027 7223 3061 7257
rect 3095 7223 3129 7257
rect 3163 7223 3197 7257
rect 3231 7223 3265 7257
rect 3299 7223 3333 7257
rect 3367 7223 3401 7257
rect 3435 7223 3469 7257
rect 3503 7223 3537 7257
rect 3571 7223 3605 7257
rect 3639 7223 3673 7257
rect 3707 7223 3741 7257
rect 3775 7223 3809 7257
rect 3843 7223 3877 7257
rect 3911 7223 3945 7257
rect 3979 7223 4013 7257
rect 4047 7223 4081 7257
rect 4115 7223 4149 7257
rect 4183 7223 4217 7257
rect 4251 7223 4285 7257
rect 4319 7223 4353 7257
rect 4387 7223 4421 7257
rect 4455 7223 4489 7257
rect 4523 7223 4557 7257
rect 4591 7223 4625 7257
rect 4659 7223 4693 7257
rect 4727 7223 4761 7257
rect 4795 7223 4829 7257
rect 4863 7223 4897 7257
rect 4931 7223 4965 7257
rect 4999 7223 5033 7257
rect 5067 7223 5101 7257
rect 5135 7223 5169 7257
rect 5203 7223 5237 7257
rect 5271 7223 5305 7257
rect 5339 7223 5373 7257
rect 5407 7223 5441 7257
rect 5475 7223 5509 7257
rect 5543 7223 5577 7257
rect 5611 7223 5645 7257
rect 5679 7223 5713 7257
rect 5747 7223 5781 7257
rect 5815 7223 5849 7257
rect 5883 7223 5917 7257
rect 5951 7223 5985 7257
rect 6019 7223 6053 7257
rect 6087 7223 6121 7257
rect 6155 7223 6189 7257
rect 6223 7223 6257 7257
rect 6291 7223 6325 7257
rect 6359 7223 6393 7257
rect 6427 7223 6461 7257
rect 6495 7223 6529 7257
rect 6563 7223 6597 7257
rect 6631 7223 6665 7257
rect 6699 7223 6733 7257
rect 6767 7223 6801 7257
rect 6835 7223 6869 7257
rect 6903 7223 6937 7257
rect 6971 7223 7005 7257
rect 7039 7223 7073 7257
rect 7107 7223 7141 7257
rect 7175 7223 7209 7257
rect 7243 7223 7277 7257
rect 7311 7223 7345 7257
rect 7379 7223 7413 7257
rect 7447 7223 7481 7257
rect 7515 7223 7549 7257
rect 7583 7223 7617 7257
rect 7651 7223 7685 7257
rect 7719 7223 7753 7257
rect 7787 7223 7821 7257
rect 7855 7223 7889 7257
rect 7923 7223 7957 7257
rect 7991 7223 8025 7257
rect 8059 7223 8093 7257
rect 8127 7223 8161 7257
rect 8195 7223 8229 7257
rect 8263 7223 8400 7257
rect 0 7200 8400 7223
rect 0 7147 80 7200
rect 0 7113 23 7147
rect 57 7113 80 7147
rect 0 7079 80 7113
rect 0 7045 23 7079
rect 57 7045 80 7079
rect 0 7011 80 7045
rect 0 6977 23 7011
rect 57 6977 80 7011
rect 0 6943 80 6977
rect 0 6909 23 6943
rect 57 6909 80 6943
rect 320 7073 400 7200
rect 320 7037 343 7073
rect 377 7037 400 7073
rect 320 7003 400 7037
rect 320 6967 343 7003
rect 377 6967 400 7003
rect 320 6920 400 6967
rect 2240 7073 2320 7120
rect 2240 7037 2263 7073
rect 2297 7037 2320 7073
rect 2240 7003 2320 7037
rect 2240 6967 2263 7003
rect 2297 6967 2320 7003
rect 2240 6920 2320 6967
rect 4160 7073 4240 7120
rect 4160 7037 4183 7073
rect 4217 7037 4240 7073
rect 4160 7003 4240 7037
rect 4160 6967 4183 7003
rect 4217 6967 4240 7003
rect 4160 6920 4240 6967
rect 6080 7073 6160 7120
rect 6080 7037 6103 7073
rect 6137 7037 6160 7073
rect 6080 7003 6160 7037
rect 6080 6967 6103 7003
rect 6137 6967 6160 7003
rect 6080 6920 6160 6967
rect 8000 7073 8080 7120
rect 8000 7037 8023 7073
rect 8057 7037 8080 7073
rect 8000 7003 8080 7037
rect 8000 6967 8023 7003
rect 8057 6967 8080 7003
rect 8000 6920 8080 6967
rect 0 6875 80 6909
rect 0 6841 23 6875
rect 57 6841 80 6875
rect 0 6807 80 6841
rect 0 6773 23 6807
rect 57 6773 80 6807
rect 520 6857 2120 6880
rect 520 6823 547 6857
rect 589 6823 619 6857
rect 657 6823 691 6857
rect 725 6823 759 6857
rect 797 6823 827 6857
rect 869 6823 895 6857
rect 941 6823 963 6857
rect 1013 6823 1031 6857
rect 1085 6823 1099 6857
rect 1157 6823 1167 6857
rect 1229 6823 1235 6857
rect 1301 6823 1303 6857
rect 1337 6823 1339 6857
rect 1405 6823 1411 6857
rect 1473 6823 1483 6857
rect 1541 6823 1555 6857
rect 1609 6823 1627 6857
rect 1677 6823 1699 6857
rect 1745 6823 1771 6857
rect 1813 6823 1843 6857
rect 1881 6823 1915 6857
rect 1949 6823 1983 6857
rect 2021 6823 2051 6857
rect 2093 6823 2120 6857
rect 520 6800 2120 6823
rect 2440 6857 4040 6880
rect 2440 6823 2467 6857
rect 2509 6823 2539 6857
rect 2577 6823 2611 6857
rect 2645 6823 2679 6857
rect 2717 6823 2747 6857
rect 2789 6823 2815 6857
rect 2861 6823 2883 6857
rect 2933 6823 2951 6857
rect 3005 6823 3019 6857
rect 3077 6823 3087 6857
rect 3149 6823 3155 6857
rect 3221 6823 3223 6857
rect 3257 6823 3259 6857
rect 3325 6823 3331 6857
rect 3393 6823 3403 6857
rect 3461 6823 3475 6857
rect 3529 6823 3547 6857
rect 3597 6823 3619 6857
rect 3665 6823 3691 6857
rect 3733 6823 3763 6857
rect 3801 6823 3835 6857
rect 3869 6823 3903 6857
rect 3941 6823 3971 6857
rect 4013 6823 4040 6857
rect 2440 6800 4040 6823
rect 4360 6857 5960 6880
rect 4360 6823 4387 6857
rect 4429 6823 4459 6857
rect 4497 6823 4531 6857
rect 4565 6823 4599 6857
rect 4637 6823 4667 6857
rect 4709 6823 4735 6857
rect 4781 6823 4803 6857
rect 4853 6823 4871 6857
rect 4925 6823 4939 6857
rect 4997 6823 5007 6857
rect 5069 6823 5075 6857
rect 5141 6823 5143 6857
rect 5177 6823 5179 6857
rect 5245 6823 5251 6857
rect 5313 6823 5323 6857
rect 5381 6823 5395 6857
rect 5449 6823 5467 6857
rect 5517 6823 5539 6857
rect 5585 6823 5611 6857
rect 5653 6823 5683 6857
rect 5721 6823 5755 6857
rect 5789 6823 5823 6857
rect 5861 6823 5891 6857
rect 5933 6823 5960 6857
rect 4360 6800 5960 6823
rect 6280 6857 7880 6880
rect 6280 6823 6307 6857
rect 6349 6823 6379 6857
rect 6417 6823 6451 6857
rect 6485 6823 6519 6857
rect 6557 6823 6587 6857
rect 6629 6823 6655 6857
rect 6701 6823 6723 6857
rect 6773 6823 6791 6857
rect 6845 6823 6859 6857
rect 6917 6823 6927 6857
rect 6989 6823 6995 6857
rect 7061 6823 7063 6857
rect 7097 6823 7099 6857
rect 7165 6823 7171 6857
rect 7233 6823 7243 6857
rect 7301 6823 7315 6857
rect 7369 6823 7387 6857
rect 7437 6823 7459 6857
rect 7505 6823 7531 6857
rect 7573 6823 7603 6857
rect 7641 6823 7675 6857
rect 7709 6823 7743 6857
rect 7781 6823 7811 6857
rect 7853 6823 7880 6857
rect 6280 6800 7880 6823
rect 0 6720 80 6773
rect 8320 6720 8400 7200
rect 0 6697 8400 6720
rect 0 6663 137 6697
rect 171 6663 205 6697
rect 239 6663 273 6697
rect 307 6663 341 6697
rect 375 6663 409 6697
rect 443 6663 477 6697
rect 511 6663 545 6697
rect 579 6663 613 6697
rect 647 6663 681 6697
rect 715 6663 749 6697
rect 783 6663 817 6697
rect 851 6663 885 6697
rect 919 6663 953 6697
rect 987 6663 1021 6697
rect 1055 6663 1089 6697
rect 1123 6663 1157 6697
rect 1191 6663 1225 6697
rect 1259 6663 1293 6697
rect 1327 6663 1361 6697
rect 1395 6663 1429 6697
rect 1463 6663 1497 6697
rect 1531 6663 1565 6697
rect 1599 6663 1633 6697
rect 1667 6663 1701 6697
rect 1735 6663 1769 6697
rect 1803 6663 1837 6697
rect 1871 6663 1905 6697
rect 1939 6663 1973 6697
rect 2007 6663 2041 6697
rect 2075 6663 2109 6697
rect 2143 6663 2177 6697
rect 2211 6663 2245 6697
rect 2279 6663 2313 6697
rect 2347 6663 2381 6697
rect 2415 6663 2449 6697
rect 2483 6663 2517 6697
rect 2551 6663 2585 6697
rect 2619 6663 2653 6697
rect 2687 6663 2721 6697
rect 2755 6663 2789 6697
rect 2823 6663 2857 6697
rect 2891 6663 2925 6697
rect 2959 6663 2993 6697
rect 3027 6663 3061 6697
rect 3095 6663 3129 6697
rect 3163 6663 3197 6697
rect 3231 6663 3265 6697
rect 3299 6663 3333 6697
rect 3367 6663 3401 6697
rect 3435 6663 3469 6697
rect 3503 6663 3537 6697
rect 3571 6663 3605 6697
rect 3639 6663 3673 6697
rect 3707 6663 3741 6697
rect 3775 6663 3809 6697
rect 3843 6663 3877 6697
rect 3911 6663 3945 6697
rect 3979 6663 4013 6697
rect 4047 6663 4081 6697
rect 4115 6663 4149 6697
rect 4183 6663 4217 6697
rect 4251 6663 4285 6697
rect 4319 6663 4353 6697
rect 4387 6663 4421 6697
rect 4455 6663 4489 6697
rect 4523 6663 4557 6697
rect 4591 6663 4625 6697
rect 4659 6663 4693 6697
rect 4727 6663 4761 6697
rect 4795 6663 4829 6697
rect 4863 6663 4897 6697
rect 4931 6663 4965 6697
rect 4999 6663 5033 6697
rect 5067 6663 5101 6697
rect 5135 6663 5169 6697
rect 5203 6663 5237 6697
rect 5271 6663 5305 6697
rect 5339 6663 5373 6697
rect 5407 6663 5441 6697
rect 5475 6663 5509 6697
rect 5543 6663 5577 6697
rect 5611 6663 5645 6697
rect 5679 6663 5713 6697
rect 5747 6663 5781 6697
rect 5815 6663 5849 6697
rect 5883 6663 5917 6697
rect 5951 6663 5985 6697
rect 6019 6663 6053 6697
rect 6087 6663 6121 6697
rect 6155 6663 6189 6697
rect 6223 6663 6257 6697
rect 6291 6663 6325 6697
rect 6359 6663 6393 6697
rect 6427 6663 6461 6697
rect 6495 6663 6529 6697
rect 6563 6663 6597 6697
rect 6631 6663 6665 6697
rect 6699 6663 6733 6697
rect 6767 6663 6801 6697
rect 6835 6663 6869 6697
rect 6903 6663 6937 6697
rect 6971 6663 7005 6697
rect 7039 6663 7073 6697
rect 7107 6663 7141 6697
rect 7175 6663 7209 6697
rect 7243 6663 7277 6697
rect 7311 6663 7345 6697
rect 7379 6663 7413 6697
rect 7447 6663 7481 6697
rect 7515 6663 7549 6697
rect 7583 6663 7617 6697
rect 7651 6663 7685 6697
rect 7719 6663 7753 6697
rect 7787 6663 7821 6697
rect 7855 6663 7889 6697
rect 7923 6663 7957 6697
rect 7991 6663 8025 6697
rect 8059 6663 8093 6697
rect 8127 6663 8161 6697
rect 8195 6663 8229 6697
rect 8263 6663 8400 6697
rect 0 6640 8400 6663
rect 0 5440 80 6640
rect 160 6377 8240 6560
rect 160 6343 183 6377
rect 217 6343 8183 6377
rect 8217 6343 8240 6377
rect 160 6320 8240 6343
rect 160 6217 8240 6240
rect 160 6183 183 6217
rect 217 6183 8183 6217
rect 8217 6183 8240 6217
rect 160 5897 8240 6183
rect 160 5863 183 5897
rect 217 5863 8183 5897
rect 8217 5863 8240 5897
rect 160 5840 8240 5863
rect 160 5737 8240 5760
rect 160 5703 183 5737
rect 217 5703 8183 5737
rect 8217 5703 8240 5737
rect 160 5520 8240 5703
rect 8320 5440 8400 6640
rect 0 5417 8400 5440
rect 0 5383 137 5417
rect 171 5383 205 5417
rect 239 5383 273 5417
rect 307 5383 341 5417
rect 375 5383 409 5417
rect 443 5383 477 5417
rect 511 5383 545 5417
rect 579 5383 613 5417
rect 647 5383 681 5417
rect 715 5383 749 5417
rect 783 5383 817 5417
rect 851 5383 885 5417
rect 919 5383 953 5417
rect 987 5383 1021 5417
rect 1055 5383 1089 5417
rect 1123 5383 1157 5417
rect 1191 5383 1225 5417
rect 1259 5383 1293 5417
rect 1327 5383 1361 5417
rect 1395 5383 1429 5417
rect 1463 5383 1497 5417
rect 1531 5383 1565 5417
rect 1599 5383 1633 5417
rect 1667 5383 1701 5417
rect 1735 5383 1769 5417
rect 1803 5383 1837 5417
rect 1871 5383 1905 5417
rect 1939 5383 1973 5417
rect 2007 5383 2041 5417
rect 2075 5383 2109 5417
rect 2143 5383 2177 5417
rect 2211 5383 2245 5417
rect 2279 5383 2313 5417
rect 2347 5383 2381 5417
rect 2415 5383 2449 5417
rect 2483 5383 2517 5417
rect 2551 5383 2585 5417
rect 2619 5383 2653 5417
rect 2687 5383 2721 5417
rect 2755 5383 2789 5417
rect 2823 5383 2857 5417
rect 2891 5383 2925 5417
rect 2959 5383 2993 5417
rect 3027 5383 3061 5417
rect 3095 5383 3129 5417
rect 3163 5383 3197 5417
rect 3231 5383 3265 5417
rect 3299 5383 3333 5417
rect 3367 5383 3401 5417
rect 3435 5383 3469 5417
rect 3503 5383 3537 5417
rect 3571 5383 3605 5417
rect 3639 5383 3673 5417
rect 3707 5383 3741 5417
rect 3775 5383 3809 5417
rect 3843 5383 3877 5417
rect 3911 5383 3945 5417
rect 3979 5383 4013 5417
rect 4047 5383 4081 5417
rect 4115 5383 4149 5417
rect 4183 5383 4217 5417
rect 4251 5383 4285 5417
rect 4319 5383 4353 5417
rect 4387 5383 4421 5417
rect 4455 5383 4489 5417
rect 4523 5383 4557 5417
rect 4591 5383 4625 5417
rect 4659 5383 4693 5417
rect 4727 5383 4761 5417
rect 4795 5383 4829 5417
rect 4863 5383 4897 5417
rect 4931 5383 4965 5417
rect 4999 5383 5033 5417
rect 5067 5383 5101 5417
rect 5135 5383 5169 5417
rect 5203 5383 5237 5417
rect 5271 5383 5305 5417
rect 5339 5383 5373 5417
rect 5407 5383 5441 5417
rect 5475 5383 5509 5417
rect 5543 5383 5577 5417
rect 5611 5383 5645 5417
rect 5679 5383 5713 5417
rect 5747 5383 5781 5417
rect 5815 5383 5849 5417
rect 5883 5383 5917 5417
rect 5951 5383 5985 5417
rect 6019 5383 6053 5417
rect 6087 5383 6121 5417
rect 6155 5383 6189 5417
rect 6223 5383 6257 5417
rect 6291 5383 6325 5417
rect 6359 5383 6393 5417
rect 6427 5383 6461 5417
rect 6495 5383 6529 5417
rect 6563 5383 6597 5417
rect 6631 5383 6665 5417
rect 6699 5383 6733 5417
rect 6767 5383 6801 5417
rect 6835 5383 6869 5417
rect 6903 5383 6937 5417
rect 6971 5383 7005 5417
rect 7039 5383 7073 5417
rect 7107 5383 7141 5417
rect 7175 5383 7209 5417
rect 7243 5383 7277 5417
rect 7311 5383 7345 5417
rect 7379 5383 7413 5417
rect 7447 5383 7481 5417
rect 7515 5383 7549 5417
rect 7583 5383 7617 5417
rect 7651 5383 7685 5417
rect 7719 5383 7753 5417
rect 7787 5383 7821 5417
rect 7855 5383 7889 5417
rect 7923 5383 7957 5417
rect 7991 5383 8025 5417
rect 8059 5383 8093 5417
rect 8127 5383 8161 5417
rect 8195 5383 8229 5417
rect 8263 5383 8400 5417
rect 0 5360 8400 5383
rect 0 5287 80 5360
rect 0 5253 23 5287
rect 57 5253 80 5287
rect 8320 5287 8400 5360
rect 0 5219 80 5253
rect 0 5185 23 5219
rect 57 5185 80 5219
rect 0 5151 80 5185
rect 0 5117 23 5151
rect 57 5117 80 5151
rect 0 5083 80 5117
rect 0 5049 23 5083
rect 57 5049 80 5083
rect 0 5015 80 5049
rect 0 4981 23 5015
rect 57 4981 80 5015
rect 0 4947 80 4981
rect 0 4913 23 4947
rect 57 4913 80 4947
rect 0 4879 80 4913
rect 0 4845 23 4879
rect 57 4845 80 4879
rect 0 4811 80 4845
rect 0 4777 23 4811
rect 57 4777 80 4811
rect 0 4743 80 4777
rect 0 4709 23 4743
rect 57 4709 80 4743
rect 0 4675 80 4709
rect 0 4641 23 4675
rect 57 4641 80 4675
rect 0 4607 80 4641
rect 0 4573 23 4607
rect 57 4573 80 4607
rect 0 4539 80 4573
rect 0 4505 23 4539
rect 57 4505 80 4539
rect 0 4471 80 4505
rect 0 4437 23 4471
rect 57 4437 80 4471
rect 0 4403 80 4437
rect 0 4369 23 4403
rect 57 4369 80 4403
rect 0 4335 80 4369
rect 0 4301 23 4335
rect 57 4301 80 4335
rect 0 4267 80 4301
rect 0 4233 23 4267
rect 57 4233 80 4267
rect 160 5257 8240 5280
rect 160 5223 307 5257
rect 341 5223 375 5257
rect 409 5223 443 5257
rect 477 5223 511 5257
rect 545 5223 579 5257
rect 613 5223 647 5257
rect 681 5223 715 5257
rect 749 5223 783 5257
rect 817 5223 851 5257
rect 885 5223 919 5257
rect 953 5223 987 5257
rect 1021 5223 1055 5257
rect 1089 5223 1123 5257
rect 1157 5223 1191 5257
rect 1225 5223 1259 5257
rect 1293 5223 1327 5257
rect 1361 5223 1395 5257
rect 1429 5223 1463 5257
rect 1497 5223 1531 5257
rect 1565 5223 1599 5257
rect 1633 5223 1667 5257
rect 1701 5223 1735 5257
rect 1769 5223 1803 5257
rect 1837 5223 1871 5257
rect 1905 5223 1939 5257
rect 1973 5223 2007 5257
rect 2041 5223 2075 5257
rect 2109 5223 2143 5257
rect 2177 5223 2211 5257
rect 2245 5223 2279 5257
rect 2313 5223 2347 5257
rect 2381 5223 2415 5257
rect 2449 5223 2483 5257
rect 2517 5223 2551 5257
rect 2585 5223 2619 5257
rect 2653 5223 2687 5257
rect 2721 5223 2755 5257
rect 2789 5223 2823 5257
rect 2857 5223 2891 5257
rect 2925 5223 2959 5257
rect 2993 5223 3027 5257
rect 3061 5223 3095 5257
rect 3129 5223 3163 5257
rect 3197 5223 3231 5257
rect 3265 5223 3299 5257
rect 3333 5223 3367 5257
rect 3401 5223 3435 5257
rect 3469 5223 3503 5257
rect 3537 5223 3571 5257
rect 3605 5223 3639 5257
rect 3673 5223 3707 5257
rect 3741 5223 3775 5257
rect 3809 5223 3843 5257
rect 3877 5223 3911 5257
rect 3945 5223 3979 5257
rect 4013 5223 4047 5257
rect 4081 5223 4115 5257
rect 4149 5223 4183 5257
rect 4217 5223 4251 5257
rect 4285 5223 4319 5257
rect 4353 5223 4387 5257
rect 4421 5223 4455 5257
rect 4489 5223 4523 5257
rect 4557 5223 4591 5257
rect 4625 5223 4659 5257
rect 4693 5223 4727 5257
rect 4761 5223 4795 5257
rect 4829 5223 4863 5257
rect 4897 5223 4931 5257
rect 4965 5223 4999 5257
rect 5033 5223 5067 5257
rect 5101 5223 5135 5257
rect 5169 5223 5203 5257
rect 5237 5223 5271 5257
rect 5305 5223 5339 5257
rect 5373 5223 5407 5257
rect 5441 5223 5475 5257
rect 5509 5223 5543 5257
rect 5577 5223 5611 5257
rect 5645 5223 5679 5257
rect 5713 5223 5747 5257
rect 5781 5223 5815 5257
rect 5849 5223 5883 5257
rect 5917 5223 5951 5257
rect 5985 5223 6019 5257
rect 6053 5223 6087 5257
rect 6121 5223 6155 5257
rect 6189 5223 6223 5257
rect 6257 5223 6291 5257
rect 6325 5223 6359 5257
rect 6393 5223 6427 5257
rect 6461 5223 6495 5257
rect 6529 5223 6563 5257
rect 6597 5223 6631 5257
rect 6665 5223 6699 5257
rect 6733 5223 6767 5257
rect 6801 5223 6835 5257
rect 6869 5223 6903 5257
rect 6937 5223 6971 5257
rect 7005 5223 7039 5257
rect 7073 5223 7107 5257
rect 7141 5223 7175 5257
rect 7209 5223 7243 5257
rect 7277 5223 7311 5257
rect 7345 5223 7379 5257
rect 7413 5223 7447 5257
rect 7481 5223 7515 5257
rect 7549 5223 7583 5257
rect 7617 5223 7651 5257
rect 7685 5223 7719 5257
rect 7753 5223 7787 5257
rect 7821 5223 7855 5257
rect 7889 5223 7923 5257
rect 7957 5223 7991 5257
rect 8025 5223 8059 5257
rect 8093 5223 8240 5257
rect 160 5200 8240 5223
rect 160 5151 240 5200
rect 160 5117 183 5151
rect 217 5117 240 5151
rect 8160 5151 8240 5200
rect 160 5083 240 5117
rect 160 5049 183 5083
rect 217 5049 240 5083
rect 160 5015 240 5049
rect 520 5097 2120 5120
rect 520 5063 547 5097
rect 589 5063 619 5097
rect 657 5063 691 5097
rect 725 5063 759 5097
rect 797 5063 827 5097
rect 869 5063 895 5097
rect 941 5063 963 5097
rect 1013 5063 1031 5097
rect 1085 5063 1099 5097
rect 1157 5063 1167 5097
rect 1229 5063 1235 5097
rect 1301 5063 1303 5097
rect 1337 5063 1339 5097
rect 1405 5063 1411 5097
rect 1473 5063 1483 5097
rect 1541 5063 1555 5097
rect 1609 5063 1627 5097
rect 1677 5063 1699 5097
rect 1745 5063 1771 5097
rect 1813 5063 1843 5097
rect 1881 5063 1915 5097
rect 1949 5063 1983 5097
rect 2021 5063 2051 5097
rect 2093 5063 2120 5097
rect 520 5040 2120 5063
rect 2440 5097 4040 5120
rect 2440 5063 2467 5097
rect 2509 5063 2539 5097
rect 2577 5063 2611 5097
rect 2645 5063 2679 5097
rect 2717 5063 2747 5097
rect 2789 5063 2815 5097
rect 2861 5063 2883 5097
rect 2933 5063 2951 5097
rect 3005 5063 3019 5097
rect 3077 5063 3087 5097
rect 3149 5063 3155 5097
rect 3221 5063 3223 5097
rect 3257 5063 3259 5097
rect 3325 5063 3331 5097
rect 3393 5063 3403 5097
rect 3461 5063 3475 5097
rect 3529 5063 3547 5097
rect 3597 5063 3619 5097
rect 3665 5063 3691 5097
rect 3733 5063 3763 5097
rect 3801 5063 3835 5097
rect 3869 5063 3903 5097
rect 3941 5063 3971 5097
rect 4013 5063 4040 5097
rect 2440 5040 4040 5063
rect 4360 5097 5960 5120
rect 4360 5063 4387 5097
rect 4429 5063 4459 5097
rect 4497 5063 4531 5097
rect 4565 5063 4599 5097
rect 4637 5063 4667 5097
rect 4709 5063 4735 5097
rect 4781 5063 4803 5097
rect 4853 5063 4871 5097
rect 4925 5063 4939 5097
rect 4997 5063 5007 5097
rect 5069 5063 5075 5097
rect 5141 5063 5143 5097
rect 5177 5063 5179 5097
rect 5245 5063 5251 5097
rect 5313 5063 5323 5097
rect 5381 5063 5395 5097
rect 5449 5063 5467 5097
rect 5517 5063 5539 5097
rect 5585 5063 5611 5097
rect 5653 5063 5683 5097
rect 5721 5063 5755 5097
rect 5789 5063 5823 5097
rect 5861 5063 5891 5097
rect 5933 5063 5960 5097
rect 4360 5040 5960 5063
rect 6280 5097 7880 5120
rect 6280 5063 6307 5097
rect 6349 5063 6379 5097
rect 6417 5063 6451 5097
rect 6485 5063 6519 5097
rect 6557 5063 6587 5097
rect 6629 5063 6655 5097
rect 6701 5063 6723 5097
rect 6773 5063 6791 5097
rect 6845 5063 6859 5097
rect 6917 5063 6927 5097
rect 6989 5063 6995 5097
rect 7061 5063 7063 5097
rect 7097 5063 7099 5097
rect 7165 5063 7171 5097
rect 7233 5063 7243 5097
rect 7301 5063 7315 5097
rect 7369 5063 7387 5097
rect 7437 5063 7459 5097
rect 7505 5063 7531 5097
rect 7573 5063 7603 5097
rect 7641 5063 7675 5097
rect 7709 5063 7743 5097
rect 7781 5063 7811 5097
rect 7853 5063 7880 5097
rect 6280 5040 7880 5063
rect 8160 5117 8183 5151
rect 8217 5117 8240 5151
rect 8160 5083 8240 5117
rect 8160 5049 8183 5083
rect 8217 5049 8240 5083
rect 160 4981 183 5015
rect 217 4981 240 5015
rect 8160 5015 8240 5049
rect 160 4947 240 4981
rect 160 4913 183 4947
rect 217 4913 240 4947
rect 160 4879 240 4913
rect 160 4845 183 4879
rect 217 4845 240 4879
rect 160 4811 240 4845
rect 160 4777 183 4811
rect 217 4777 240 4811
rect 160 4743 240 4777
rect 160 4709 183 4743
rect 217 4709 240 4743
rect 160 4675 240 4709
rect 160 4641 183 4675
rect 217 4641 240 4675
rect 160 4607 240 4641
rect 160 4573 183 4607
rect 217 4573 240 4607
rect 160 4539 240 4573
rect 160 4505 183 4539
rect 217 4505 240 4539
rect 160 4471 240 4505
rect 160 4437 183 4471
rect 217 4437 240 4471
rect 160 4403 240 4437
rect 160 4369 183 4403
rect 217 4369 240 4403
rect 160 4320 240 4369
rect 320 4969 400 5000
rect 320 4921 343 4969
rect 377 4921 400 4969
rect 320 4897 400 4921
rect 320 4853 343 4897
rect 377 4853 400 4897
rect 320 4825 400 4853
rect 320 4785 343 4825
rect 377 4785 400 4825
rect 320 4753 400 4785
rect 320 4717 343 4753
rect 377 4717 400 4753
rect 320 4683 400 4717
rect 320 4647 343 4683
rect 377 4647 400 4683
rect 320 4615 400 4647
rect 320 4575 343 4615
rect 377 4575 400 4615
rect 320 4547 400 4575
rect 320 4503 343 4547
rect 377 4503 400 4547
rect 320 4479 400 4503
rect 320 4431 343 4479
rect 377 4431 400 4479
rect 320 4320 400 4431
rect 2240 4969 2320 5000
rect 2240 4921 2263 4969
rect 2297 4921 2320 4969
rect 2240 4897 2320 4921
rect 2240 4853 2263 4897
rect 2297 4853 2320 4897
rect 2240 4825 2320 4853
rect 2240 4785 2263 4825
rect 2297 4785 2320 4825
rect 2240 4753 2320 4785
rect 2240 4717 2263 4753
rect 2297 4717 2320 4753
rect 2240 4683 2320 4717
rect 2240 4647 2263 4683
rect 2297 4647 2320 4683
rect 2240 4615 2320 4647
rect 2240 4575 2263 4615
rect 2297 4575 2320 4615
rect 2240 4547 2320 4575
rect 2240 4503 2263 4547
rect 2297 4503 2320 4547
rect 2240 4479 2320 4503
rect 2240 4431 2263 4479
rect 2297 4431 2320 4479
rect 2240 4400 2320 4431
rect 4160 4969 4240 5000
rect 4160 4921 4183 4969
rect 4217 4921 4240 4969
rect 4160 4897 4240 4921
rect 4160 4853 4183 4897
rect 4217 4853 4240 4897
rect 4160 4825 4240 4853
rect 4160 4785 4183 4825
rect 4217 4785 4240 4825
rect 4160 4753 4240 4785
rect 4160 4717 4183 4753
rect 4217 4717 4240 4753
rect 4160 4683 4240 4717
rect 4160 4647 4183 4683
rect 4217 4647 4240 4683
rect 4160 4615 4240 4647
rect 4160 4575 4183 4615
rect 4217 4575 4240 4615
rect 4160 4547 4240 4575
rect 4160 4503 4183 4547
rect 4217 4503 4240 4547
rect 4160 4479 4240 4503
rect 4160 4431 4183 4479
rect 4217 4431 4240 4479
rect 4160 4400 4240 4431
rect 6080 4969 6160 5000
rect 6080 4921 6103 4969
rect 6137 4921 6160 4969
rect 6080 4897 6160 4921
rect 6080 4853 6103 4897
rect 6137 4853 6160 4897
rect 6080 4825 6160 4853
rect 6080 4785 6103 4825
rect 6137 4785 6160 4825
rect 6080 4753 6160 4785
rect 6080 4717 6103 4753
rect 6137 4717 6160 4753
rect 6080 4683 6160 4717
rect 6080 4647 6103 4683
rect 6137 4647 6160 4683
rect 6080 4615 6160 4647
rect 6080 4575 6103 4615
rect 6137 4575 6160 4615
rect 6080 4547 6160 4575
rect 6080 4503 6103 4547
rect 6137 4503 6160 4547
rect 6080 4479 6160 4503
rect 6080 4431 6103 4479
rect 6137 4431 6160 4479
rect 6080 4400 6160 4431
rect 8000 4969 8080 5000
rect 8000 4921 8023 4969
rect 8057 4921 8080 4969
rect 8000 4897 8080 4921
rect 8000 4853 8023 4897
rect 8057 4853 8080 4897
rect 8000 4825 8080 4853
rect 8000 4785 8023 4825
rect 8057 4785 8080 4825
rect 8000 4753 8080 4785
rect 8000 4717 8023 4753
rect 8057 4717 8080 4753
rect 8000 4683 8080 4717
rect 8000 4647 8023 4683
rect 8057 4647 8080 4683
rect 8000 4615 8080 4647
rect 8000 4575 8023 4615
rect 8057 4575 8080 4615
rect 8000 4547 8080 4575
rect 8000 4503 8023 4547
rect 8057 4503 8080 4547
rect 8000 4479 8080 4503
rect 8000 4431 8023 4479
rect 8057 4431 8080 4479
rect 8000 4400 8080 4431
rect 8160 4981 8183 5015
rect 8217 4981 8240 5015
rect 8160 4947 8240 4981
rect 8160 4913 8183 4947
rect 8217 4913 8240 4947
rect 8160 4879 8240 4913
rect 8160 4845 8183 4879
rect 8217 4845 8240 4879
rect 8160 4811 8240 4845
rect 8160 4777 8183 4811
rect 8217 4777 8240 4811
rect 8160 4743 8240 4777
rect 8160 4709 8183 4743
rect 8217 4709 8240 4743
rect 8160 4675 8240 4709
rect 8160 4641 8183 4675
rect 8217 4641 8240 4675
rect 8160 4607 8240 4641
rect 8160 4573 8183 4607
rect 8217 4573 8240 4607
rect 8160 4539 8240 4573
rect 8160 4505 8183 4539
rect 8217 4505 8240 4539
rect 8160 4471 8240 4505
rect 8160 4437 8183 4471
rect 8217 4437 8240 4471
rect 8160 4403 8240 4437
rect 8160 4369 8183 4403
rect 8217 4369 8240 4403
rect 8160 4320 8240 4369
rect 160 4297 8240 4320
rect 160 4263 307 4297
rect 341 4263 375 4297
rect 409 4263 443 4297
rect 477 4263 511 4297
rect 545 4263 579 4297
rect 613 4263 647 4297
rect 681 4263 715 4297
rect 749 4263 783 4297
rect 817 4263 851 4297
rect 885 4263 919 4297
rect 953 4263 987 4297
rect 1021 4263 1055 4297
rect 1089 4263 1123 4297
rect 1157 4263 1191 4297
rect 1225 4263 1259 4297
rect 1293 4263 1327 4297
rect 1361 4263 1395 4297
rect 1429 4263 1463 4297
rect 1497 4263 1531 4297
rect 1565 4263 1599 4297
rect 1633 4263 1667 4297
rect 1701 4263 1735 4297
rect 1769 4263 1803 4297
rect 1837 4263 1871 4297
rect 1905 4263 1939 4297
rect 1973 4263 2007 4297
rect 2041 4263 2075 4297
rect 2109 4263 2143 4297
rect 2177 4263 2211 4297
rect 2245 4263 2279 4297
rect 2313 4263 2347 4297
rect 2381 4263 2415 4297
rect 2449 4263 2483 4297
rect 2517 4263 2551 4297
rect 2585 4263 2619 4297
rect 2653 4263 2687 4297
rect 2721 4263 2755 4297
rect 2789 4263 2823 4297
rect 2857 4263 2891 4297
rect 2925 4263 2959 4297
rect 2993 4263 3027 4297
rect 3061 4263 3095 4297
rect 3129 4263 3163 4297
rect 3197 4263 3231 4297
rect 3265 4263 3299 4297
rect 3333 4263 3367 4297
rect 3401 4263 3435 4297
rect 3469 4263 3503 4297
rect 3537 4263 3571 4297
rect 3605 4263 3639 4297
rect 3673 4263 3707 4297
rect 3741 4263 3775 4297
rect 3809 4263 3843 4297
rect 3877 4263 3911 4297
rect 3945 4263 3979 4297
rect 4013 4263 4047 4297
rect 4081 4263 4115 4297
rect 4149 4263 4183 4297
rect 4217 4263 4251 4297
rect 4285 4263 4319 4297
rect 4353 4263 4387 4297
rect 4421 4263 4455 4297
rect 4489 4263 4523 4297
rect 4557 4263 4591 4297
rect 4625 4263 4659 4297
rect 4693 4263 4727 4297
rect 4761 4263 4795 4297
rect 4829 4263 4863 4297
rect 4897 4263 4931 4297
rect 4965 4263 4999 4297
rect 5033 4263 5067 4297
rect 5101 4263 5135 4297
rect 5169 4263 5203 4297
rect 5237 4263 5271 4297
rect 5305 4263 5339 4297
rect 5373 4263 5407 4297
rect 5441 4263 5475 4297
rect 5509 4263 5543 4297
rect 5577 4263 5611 4297
rect 5645 4263 5679 4297
rect 5713 4263 5747 4297
rect 5781 4263 5815 4297
rect 5849 4263 5883 4297
rect 5917 4263 5951 4297
rect 5985 4263 6019 4297
rect 6053 4263 6087 4297
rect 6121 4263 6155 4297
rect 6189 4263 6223 4297
rect 6257 4263 6291 4297
rect 6325 4263 6359 4297
rect 6393 4263 6427 4297
rect 6461 4263 6495 4297
rect 6529 4263 6563 4297
rect 6597 4263 6631 4297
rect 6665 4263 6699 4297
rect 6733 4263 6767 4297
rect 6801 4263 6835 4297
rect 6869 4263 6903 4297
rect 6937 4263 6971 4297
rect 7005 4263 7039 4297
rect 7073 4263 7107 4297
rect 7141 4263 7175 4297
rect 7209 4263 7243 4297
rect 7277 4263 7311 4297
rect 7345 4263 7379 4297
rect 7413 4263 7447 4297
rect 7481 4263 7515 4297
rect 7549 4263 7583 4297
rect 7617 4263 7651 4297
rect 7685 4263 7719 4297
rect 7753 4263 7787 4297
rect 7821 4263 7855 4297
rect 7889 4263 7923 4297
rect 7957 4263 7991 4297
rect 8025 4263 8059 4297
rect 8093 4263 8240 4297
rect 160 4240 8240 4263
rect 8320 5253 8343 5287
rect 8377 5253 8400 5287
rect 8320 5219 8400 5253
rect 8320 5185 8343 5219
rect 8377 5185 8400 5219
rect 8320 5151 8400 5185
rect 8320 5117 8343 5151
rect 8377 5117 8400 5151
rect 8320 5083 8400 5117
rect 8320 5049 8343 5083
rect 8377 5049 8400 5083
rect 8320 5015 8400 5049
rect 8320 4981 8343 5015
rect 8377 4981 8400 5015
rect 8320 4947 8400 4981
rect 8320 4913 8343 4947
rect 8377 4913 8400 4947
rect 8320 4879 8400 4913
rect 8320 4845 8343 4879
rect 8377 4845 8400 4879
rect 8320 4811 8400 4845
rect 8320 4777 8343 4811
rect 8377 4777 8400 4811
rect 8320 4743 8400 4777
rect 8320 4709 8343 4743
rect 8377 4709 8400 4743
rect 8320 4675 8400 4709
rect 8320 4641 8343 4675
rect 8377 4641 8400 4675
rect 8320 4607 8400 4641
rect 8320 4573 8343 4607
rect 8377 4573 8400 4607
rect 8320 4539 8400 4573
rect 8320 4505 8343 4539
rect 8377 4505 8400 4539
rect 8320 4471 8400 4505
rect 8320 4437 8343 4471
rect 8377 4437 8400 4471
rect 8320 4403 8400 4437
rect 8320 4369 8343 4403
rect 8377 4369 8400 4403
rect 8320 4335 8400 4369
rect 8320 4301 8343 4335
rect 8377 4301 8400 4335
rect 8320 4267 8400 4301
rect 0 4160 80 4233
rect 8320 4233 8343 4267
rect 8377 4233 8400 4267
rect 8320 4160 8400 4233
rect 0 4137 8400 4160
rect 0 4103 137 4137
rect 171 4103 205 4137
rect 239 4103 273 4137
rect 307 4103 341 4137
rect 375 4103 409 4137
rect 443 4103 477 4137
rect 511 4103 545 4137
rect 579 4103 613 4137
rect 647 4103 681 4137
rect 715 4103 749 4137
rect 783 4103 817 4137
rect 851 4103 885 4137
rect 919 4103 953 4137
rect 987 4103 1021 4137
rect 1055 4103 1089 4137
rect 1123 4103 1157 4137
rect 1191 4103 1225 4137
rect 1259 4103 1293 4137
rect 1327 4103 1361 4137
rect 1395 4103 1429 4137
rect 1463 4103 1497 4137
rect 1531 4103 1565 4137
rect 1599 4103 1633 4137
rect 1667 4103 1701 4137
rect 1735 4103 1769 4137
rect 1803 4103 1837 4137
rect 1871 4103 1905 4137
rect 1939 4103 1973 4137
rect 2007 4103 2041 4137
rect 2075 4103 2109 4137
rect 2143 4103 2177 4137
rect 2211 4103 2245 4137
rect 2279 4103 2313 4137
rect 2347 4103 2381 4137
rect 2415 4103 2449 4137
rect 2483 4103 2517 4137
rect 2551 4103 2585 4137
rect 2619 4103 2653 4137
rect 2687 4103 2721 4137
rect 2755 4103 2789 4137
rect 2823 4103 2857 4137
rect 2891 4103 2925 4137
rect 2959 4103 2993 4137
rect 3027 4103 3061 4137
rect 3095 4103 3129 4137
rect 3163 4103 3197 4137
rect 3231 4103 3265 4137
rect 3299 4103 3333 4137
rect 3367 4103 3401 4137
rect 3435 4103 3469 4137
rect 3503 4103 3537 4137
rect 3571 4103 3605 4137
rect 3639 4103 3673 4137
rect 3707 4103 3741 4137
rect 3775 4103 3809 4137
rect 3843 4103 3877 4137
rect 3911 4103 3945 4137
rect 3979 4103 4013 4137
rect 4047 4103 4081 4137
rect 4115 4103 4149 4137
rect 4183 4103 4217 4137
rect 4251 4103 4285 4137
rect 4319 4103 4353 4137
rect 4387 4103 4421 4137
rect 4455 4103 4489 4137
rect 4523 4103 4557 4137
rect 4591 4103 4625 4137
rect 4659 4103 4693 4137
rect 4727 4103 4761 4137
rect 4795 4103 4829 4137
rect 4863 4103 4897 4137
rect 4931 4103 4965 4137
rect 4999 4103 5033 4137
rect 5067 4103 5101 4137
rect 5135 4103 5169 4137
rect 5203 4103 5237 4137
rect 5271 4103 5305 4137
rect 5339 4103 5373 4137
rect 5407 4103 5441 4137
rect 5475 4103 5509 4137
rect 5543 4103 5577 4137
rect 5611 4103 5645 4137
rect 5679 4103 5713 4137
rect 5747 4103 5781 4137
rect 5815 4103 5849 4137
rect 5883 4103 5917 4137
rect 5951 4103 5985 4137
rect 6019 4103 6053 4137
rect 6087 4103 6121 4137
rect 6155 4103 6189 4137
rect 6223 4103 6257 4137
rect 6291 4103 6325 4137
rect 6359 4103 6393 4137
rect 6427 4103 6461 4137
rect 6495 4103 6529 4137
rect 6563 4103 6597 4137
rect 6631 4103 6665 4137
rect 6699 4103 6733 4137
rect 6767 4103 6801 4137
rect 6835 4103 6869 4137
rect 6903 4103 6937 4137
rect 6971 4103 7005 4137
rect 7039 4103 7073 4137
rect 7107 4103 7141 4137
rect 7175 4103 7209 4137
rect 7243 4103 7277 4137
rect 7311 4103 7345 4137
rect 7379 4103 7413 4137
rect 7447 4103 7481 4137
rect 7515 4103 7549 4137
rect 7583 4103 7617 4137
rect 7651 4103 7685 4137
rect 7719 4103 7753 4137
rect 7787 4103 7821 4137
rect 7855 4103 7889 4137
rect 7923 4103 7957 4137
rect 7991 4103 8025 4137
rect 8059 4103 8093 4137
rect 8127 4103 8161 4137
rect 8195 4103 8229 4137
rect 8263 4103 8400 4137
rect 0 4080 8400 4103
rect 0 4000 80 4080
rect 8320 4000 8400 4080
rect 0 3977 8400 4000
rect 0 3943 137 3977
rect 171 3943 205 3977
rect 239 3943 273 3977
rect 307 3943 341 3977
rect 375 3943 409 3977
rect 443 3943 477 3977
rect 511 3943 545 3977
rect 579 3943 613 3977
rect 647 3943 681 3977
rect 715 3943 749 3977
rect 783 3943 817 3977
rect 851 3943 885 3977
rect 919 3943 953 3977
rect 987 3943 1021 3977
rect 1055 3943 1089 3977
rect 1123 3943 1157 3977
rect 1191 3943 1225 3977
rect 1259 3943 1293 3977
rect 1327 3943 1361 3977
rect 1395 3943 1429 3977
rect 1463 3943 1497 3977
rect 1531 3943 1565 3977
rect 1599 3943 1633 3977
rect 1667 3943 1701 3977
rect 1735 3943 1769 3977
rect 1803 3943 1837 3977
rect 1871 3943 1905 3977
rect 1939 3943 1973 3977
rect 2007 3943 2041 3977
rect 2075 3943 2109 3977
rect 2143 3943 2177 3977
rect 2211 3943 2245 3977
rect 2279 3943 2313 3977
rect 2347 3943 2381 3977
rect 2415 3943 2449 3977
rect 2483 3943 2517 3977
rect 2551 3943 2585 3977
rect 2619 3943 2653 3977
rect 2687 3943 2721 3977
rect 2755 3943 2789 3977
rect 2823 3943 2857 3977
rect 2891 3943 2925 3977
rect 2959 3943 2993 3977
rect 3027 3943 3061 3977
rect 3095 3943 3129 3977
rect 3163 3943 3197 3977
rect 3231 3943 3265 3977
rect 3299 3943 3333 3977
rect 3367 3943 3401 3977
rect 3435 3943 3469 3977
rect 3503 3943 3537 3977
rect 3571 3943 3605 3977
rect 3639 3943 3673 3977
rect 3707 3943 3741 3977
rect 3775 3943 3809 3977
rect 3843 3943 3877 3977
rect 3911 3943 3945 3977
rect 3979 3943 4013 3977
rect 4047 3943 4081 3977
rect 4115 3943 4149 3977
rect 4183 3943 4217 3977
rect 4251 3943 4285 3977
rect 4319 3943 4353 3977
rect 4387 3943 4421 3977
rect 4455 3943 4489 3977
rect 4523 3943 4557 3977
rect 4591 3943 4625 3977
rect 4659 3943 4693 3977
rect 4727 3943 4761 3977
rect 4795 3943 4829 3977
rect 4863 3943 4897 3977
rect 4931 3943 4965 3977
rect 4999 3943 5033 3977
rect 5067 3943 5101 3977
rect 5135 3943 5169 3977
rect 5203 3943 5237 3977
rect 5271 3943 5305 3977
rect 5339 3943 5373 3977
rect 5407 3943 5441 3977
rect 5475 3943 5509 3977
rect 5543 3943 5577 3977
rect 5611 3943 5645 3977
rect 5679 3943 5713 3977
rect 5747 3943 5781 3977
rect 5815 3943 5849 3977
rect 5883 3943 5917 3977
rect 5951 3943 5985 3977
rect 6019 3943 6053 3977
rect 6087 3943 6121 3977
rect 6155 3943 6189 3977
rect 6223 3943 6257 3977
rect 6291 3943 6325 3977
rect 6359 3943 6393 3977
rect 6427 3943 6461 3977
rect 6495 3943 6529 3977
rect 6563 3943 6597 3977
rect 6631 3943 6665 3977
rect 6699 3943 6733 3977
rect 6767 3943 6801 3977
rect 6835 3943 6869 3977
rect 6903 3943 6937 3977
rect 6971 3943 7005 3977
rect 7039 3943 7073 3977
rect 7107 3943 7141 3977
rect 7175 3943 7209 3977
rect 7243 3943 7277 3977
rect 7311 3943 7345 3977
rect 7379 3943 7413 3977
rect 7447 3943 7481 3977
rect 7515 3943 7549 3977
rect 7583 3943 7617 3977
rect 7651 3943 7685 3977
rect 7719 3943 7753 3977
rect 7787 3943 7821 3977
rect 7855 3943 7889 3977
rect 7923 3943 7957 3977
rect 7991 3943 8025 3977
rect 8059 3943 8093 3977
rect 8127 3943 8161 3977
rect 8195 3943 8229 3977
rect 8263 3943 8400 3977
rect 0 3920 8400 3943
rect 0 3847 80 3920
rect 0 3813 23 3847
rect 57 3813 80 3847
rect 8320 3847 8400 3920
rect 0 3779 80 3813
rect 0 3745 23 3779
rect 57 3745 80 3779
rect 0 3711 80 3745
rect 0 3677 23 3711
rect 57 3677 80 3711
rect 0 3643 80 3677
rect 0 3609 23 3643
rect 57 3609 80 3643
rect 0 3575 80 3609
rect 0 3541 23 3575
rect 57 3541 80 3575
rect 0 3507 80 3541
rect 0 3473 23 3507
rect 57 3473 80 3507
rect 0 3439 80 3473
rect 0 3405 23 3439
rect 57 3405 80 3439
rect 0 3371 80 3405
rect 0 3337 23 3371
rect 57 3337 80 3371
rect 0 3303 80 3337
rect 0 3269 23 3303
rect 57 3269 80 3303
rect 0 3235 80 3269
rect 0 3201 23 3235
rect 57 3201 80 3235
rect 0 3167 80 3201
rect 0 3133 23 3167
rect 57 3133 80 3167
rect 0 3099 80 3133
rect 0 3065 23 3099
rect 57 3065 80 3099
rect 0 3031 80 3065
rect 0 2997 23 3031
rect 57 2997 80 3031
rect 0 2963 80 2997
rect 0 2929 23 2963
rect 57 2929 80 2963
rect 0 2895 80 2929
rect 0 2861 23 2895
rect 57 2861 80 2895
rect 0 2827 80 2861
rect 0 2793 23 2827
rect 57 2793 80 2827
rect 160 3817 8240 3840
rect 160 3783 307 3817
rect 341 3783 375 3817
rect 409 3783 443 3817
rect 477 3783 511 3817
rect 545 3783 579 3817
rect 613 3783 647 3817
rect 681 3783 715 3817
rect 749 3783 783 3817
rect 817 3783 851 3817
rect 885 3783 919 3817
rect 953 3783 987 3817
rect 1021 3783 1055 3817
rect 1089 3783 1123 3817
rect 1157 3783 1191 3817
rect 1225 3783 1259 3817
rect 1293 3783 1327 3817
rect 1361 3783 1395 3817
rect 1429 3783 1463 3817
rect 1497 3783 1531 3817
rect 1565 3783 1599 3817
rect 1633 3783 1667 3817
rect 1701 3783 1735 3817
rect 1769 3783 1803 3817
rect 1837 3783 1871 3817
rect 1905 3783 1939 3817
rect 1973 3783 2007 3817
rect 2041 3783 2075 3817
rect 2109 3783 2143 3817
rect 2177 3783 2211 3817
rect 2245 3783 2279 3817
rect 2313 3783 2347 3817
rect 2381 3783 2415 3817
rect 2449 3783 2483 3817
rect 2517 3783 2551 3817
rect 2585 3783 2619 3817
rect 2653 3783 2687 3817
rect 2721 3783 2755 3817
rect 2789 3783 2823 3817
rect 2857 3783 2891 3817
rect 2925 3783 2959 3817
rect 2993 3783 3027 3817
rect 3061 3783 3095 3817
rect 3129 3783 3163 3817
rect 3197 3783 3231 3817
rect 3265 3783 3299 3817
rect 3333 3783 3367 3817
rect 3401 3783 3435 3817
rect 3469 3783 3503 3817
rect 3537 3783 3571 3817
rect 3605 3783 3639 3817
rect 3673 3783 3707 3817
rect 3741 3783 3775 3817
rect 3809 3783 3843 3817
rect 3877 3783 3911 3817
rect 3945 3783 3979 3817
rect 4013 3783 4047 3817
rect 4081 3783 4115 3817
rect 4149 3783 4183 3817
rect 4217 3783 4251 3817
rect 4285 3783 4319 3817
rect 4353 3783 4387 3817
rect 4421 3783 4455 3817
rect 4489 3783 4523 3817
rect 4557 3783 4591 3817
rect 4625 3783 4659 3817
rect 4693 3783 4727 3817
rect 4761 3783 4795 3817
rect 4829 3783 4863 3817
rect 4897 3783 4931 3817
rect 4965 3783 4999 3817
rect 5033 3783 5067 3817
rect 5101 3783 5135 3817
rect 5169 3783 5203 3817
rect 5237 3783 5271 3817
rect 5305 3783 5339 3817
rect 5373 3783 5407 3817
rect 5441 3783 5475 3817
rect 5509 3783 5543 3817
rect 5577 3783 5611 3817
rect 5645 3783 5679 3817
rect 5713 3783 5747 3817
rect 5781 3783 5815 3817
rect 5849 3783 5883 3817
rect 5917 3783 5951 3817
rect 5985 3783 6019 3817
rect 6053 3783 6087 3817
rect 6121 3783 6155 3817
rect 6189 3783 6223 3817
rect 6257 3783 6291 3817
rect 6325 3783 6359 3817
rect 6393 3783 6427 3817
rect 6461 3783 6495 3817
rect 6529 3783 6563 3817
rect 6597 3783 6631 3817
rect 6665 3783 6699 3817
rect 6733 3783 6767 3817
rect 6801 3783 6835 3817
rect 6869 3783 6903 3817
rect 6937 3783 6971 3817
rect 7005 3783 7039 3817
rect 7073 3783 7107 3817
rect 7141 3783 7175 3817
rect 7209 3783 7243 3817
rect 7277 3783 7311 3817
rect 7345 3783 7379 3817
rect 7413 3783 7447 3817
rect 7481 3783 7515 3817
rect 7549 3783 7583 3817
rect 7617 3783 7651 3817
rect 7685 3783 7719 3817
rect 7753 3783 7787 3817
rect 7821 3783 7855 3817
rect 7889 3783 7923 3817
rect 7957 3783 7991 3817
rect 8025 3783 8059 3817
rect 8093 3783 8240 3817
rect 160 3760 8240 3783
rect 160 3711 240 3760
rect 160 3677 183 3711
rect 217 3677 240 3711
rect 160 3643 240 3677
rect 160 3609 183 3643
rect 217 3609 240 3643
rect 160 3575 240 3609
rect 160 3541 183 3575
rect 217 3541 240 3575
rect 160 3507 240 3541
rect 160 3473 183 3507
rect 217 3473 240 3507
rect 160 3439 240 3473
rect 160 3405 183 3439
rect 217 3405 240 3439
rect 160 3371 240 3405
rect 160 3337 183 3371
rect 217 3337 240 3371
rect 160 3303 240 3337
rect 160 3269 183 3303
rect 217 3269 240 3303
rect 160 3235 240 3269
rect 160 3201 183 3235
rect 217 3201 240 3235
rect 160 3167 240 3201
rect 160 3133 183 3167
rect 217 3133 240 3167
rect 160 3099 240 3133
rect 160 3065 183 3099
rect 217 3065 240 3099
rect 320 3649 400 3680
rect 320 3601 343 3649
rect 377 3601 400 3649
rect 320 3577 400 3601
rect 320 3533 343 3577
rect 377 3533 400 3577
rect 320 3505 400 3533
rect 320 3465 343 3505
rect 377 3465 400 3505
rect 320 3433 400 3465
rect 320 3397 343 3433
rect 377 3397 400 3433
rect 320 3363 400 3397
rect 320 3327 343 3363
rect 377 3327 400 3363
rect 320 3295 400 3327
rect 320 3255 343 3295
rect 377 3255 400 3295
rect 320 3227 400 3255
rect 320 3183 343 3227
rect 377 3183 400 3227
rect 320 3159 400 3183
rect 320 3111 343 3159
rect 377 3111 400 3159
rect 320 3080 400 3111
rect 2240 3649 2320 3680
rect 2240 3601 2263 3649
rect 2297 3601 2320 3649
rect 2240 3577 2320 3601
rect 2240 3533 2263 3577
rect 2297 3533 2320 3577
rect 2240 3505 2320 3533
rect 2240 3465 2263 3505
rect 2297 3465 2320 3505
rect 2240 3433 2320 3465
rect 2240 3397 2263 3433
rect 2297 3397 2320 3433
rect 2240 3363 2320 3397
rect 2240 3327 2263 3363
rect 2297 3327 2320 3363
rect 2240 3295 2320 3327
rect 2240 3255 2263 3295
rect 2297 3255 2320 3295
rect 2240 3227 2320 3255
rect 2240 3183 2263 3227
rect 2297 3183 2320 3227
rect 2240 3159 2320 3183
rect 2240 3111 2263 3159
rect 2297 3111 2320 3159
rect 2240 3080 2320 3111
rect 4160 3649 4240 3680
rect 4160 3601 4183 3649
rect 4217 3601 4240 3649
rect 4160 3577 4240 3601
rect 4160 3533 4183 3577
rect 4217 3533 4240 3577
rect 4160 3505 4240 3533
rect 4160 3465 4183 3505
rect 4217 3465 4240 3505
rect 4160 3433 4240 3465
rect 4160 3397 4183 3433
rect 4217 3397 4240 3433
rect 4160 3363 4240 3397
rect 4160 3327 4183 3363
rect 4217 3327 4240 3363
rect 4160 3295 4240 3327
rect 4160 3255 4183 3295
rect 4217 3255 4240 3295
rect 4160 3227 4240 3255
rect 4160 3183 4183 3227
rect 4217 3183 4240 3227
rect 4160 3159 4240 3183
rect 4160 3111 4183 3159
rect 4217 3111 4240 3159
rect 4160 3080 4240 3111
rect 6080 3649 6160 3680
rect 6080 3601 6103 3649
rect 6137 3601 6160 3649
rect 6080 3577 6160 3601
rect 6080 3533 6103 3577
rect 6137 3533 6160 3577
rect 6080 3505 6160 3533
rect 6080 3465 6103 3505
rect 6137 3465 6160 3505
rect 6080 3433 6160 3465
rect 6080 3397 6103 3433
rect 6137 3397 6160 3433
rect 6080 3363 6160 3397
rect 6080 3327 6103 3363
rect 6137 3327 6160 3363
rect 6080 3295 6160 3327
rect 6080 3255 6103 3295
rect 6137 3255 6160 3295
rect 6080 3227 6160 3255
rect 6080 3183 6103 3227
rect 6137 3183 6160 3227
rect 6080 3159 6160 3183
rect 6080 3111 6103 3159
rect 6137 3111 6160 3159
rect 6080 3080 6160 3111
rect 8000 3649 8080 3760
rect 8000 3601 8023 3649
rect 8057 3601 8080 3649
rect 8000 3577 8080 3601
rect 8000 3533 8023 3577
rect 8057 3533 8080 3577
rect 8000 3505 8080 3533
rect 8000 3465 8023 3505
rect 8057 3465 8080 3505
rect 8000 3433 8080 3465
rect 8000 3397 8023 3433
rect 8057 3397 8080 3433
rect 8000 3363 8080 3397
rect 8000 3327 8023 3363
rect 8057 3327 8080 3363
rect 8000 3295 8080 3327
rect 8000 3255 8023 3295
rect 8057 3255 8080 3295
rect 8000 3227 8080 3255
rect 8000 3183 8023 3227
rect 8057 3183 8080 3227
rect 8000 3159 8080 3183
rect 8000 3111 8023 3159
rect 8057 3111 8080 3159
rect 8000 3080 8080 3111
rect 8160 3711 8240 3760
rect 8160 3677 8183 3711
rect 8217 3677 8240 3711
rect 8160 3643 8240 3677
rect 8160 3609 8183 3643
rect 8217 3609 8240 3643
rect 8160 3575 8240 3609
rect 8160 3541 8183 3575
rect 8217 3541 8240 3575
rect 8160 3507 8240 3541
rect 8160 3473 8183 3507
rect 8217 3473 8240 3507
rect 8160 3439 8240 3473
rect 8160 3405 8183 3439
rect 8217 3405 8240 3439
rect 8160 3371 8240 3405
rect 8160 3337 8183 3371
rect 8217 3337 8240 3371
rect 8160 3303 8240 3337
rect 8160 3269 8183 3303
rect 8217 3269 8240 3303
rect 8160 3235 8240 3269
rect 8160 3201 8183 3235
rect 8217 3201 8240 3235
rect 8160 3167 8240 3201
rect 8160 3133 8183 3167
rect 8217 3133 8240 3167
rect 8160 3099 8240 3133
rect 160 3031 240 3065
rect 8160 3065 8183 3099
rect 8217 3065 8240 3099
rect 160 2997 183 3031
rect 217 2997 240 3031
rect 160 2963 240 2997
rect 160 2929 183 2963
rect 217 2929 240 2963
rect 520 3017 2120 3040
rect 520 2983 547 3017
rect 589 2983 619 3017
rect 657 2983 691 3017
rect 725 2983 759 3017
rect 797 2983 827 3017
rect 869 2983 895 3017
rect 941 2983 963 3017
rect 1013 2983 1031 3017
rect 1085 2983 1099 3017
rect 1157 2983 1167 3017
rect 1229 2983 1235 3017
rect 1301 2983 1303 3017
rect 1337 2983 1339 3017
rect 1405 2983 1411 3017
rect 1473 2983 1483 3017
rect 1541 2983 1555 3017
rect 1609 2983 1627 3017
rect 1677 2983 1699 3017
rect 1745 2983 1771 3017
rect 1813 2983 1843 3017
rect 1881 2983 1915 3017
rect 1949 2983 1983 3017
rect 2021 2983 2051 3017
rect 2093 2983 2120 3017
rect 520 2960 2120 2983
rect 2440 3017 4040 3040
rect 2440 2983 2467 3017
rect 2509 2983 2539 3017
rect 2577 2983 2611 3017
rect 2645 2983 2679 3017
rect 2717 2983 2747 3017
rect 2789 2983 2815 3017
rect 2861 2983 2883 3017
rect 2933 2983 2951 3017
rect 3005 2983 3019 3017
rect 3077 2983 3087 3017
rect 3149 2983 3155 3017
rect 3221 2983 3223 3017
rect 3257 2983 3259 3017
rect 3325 2983 3331 3017
rect 3393 2983 3403 3017
rect 3461 2983 3475 3017
rect 3529 2983 3547 3017
rect 3597 2983 3619 3017
rect 3665 2983 3691 3017
rect 3733 2983 3763 3017
rect 3801 2983 3835 3017
rect 3869 2983 3903 3017
rect 3941 2983 3971 3017
rect 4013 2983 4040 3017
rect 2440 2960 4040 2983
rect 4360 3017 5960 3040
rect 4360 2983 4387 3017
rect 4429 2983 4459 3017
rect 4497 2983 4531 3017
rect 4565 2983 4599 3017
rect 4637 2983 4667 3017
rect 4709 2983 4735 3017
rect 4781 2983 4803 3017
rect 4853 2983 4871 3017
rect 4925 2983 4939 3017
rect 4997 2983 5007 3017
rect 5069 2983 5075 3017
rect 5141 2983 5143 3017
rect 5177 2983 5179 3017
rect 5245 2983 5251 3017
rect 5313 2983 5323 3017
rect 5381 2983 5395 3017
rect 5449 2983 5467 3017
rect 5517 2983 5539 3017
rect 5585 2983 5611 3017
rect 5653 2983 5683 3017
rect 5721 2983 5755 3017
rect 5789 2983 5823 3017
rect 5861 2983 5891 3017
rect 5933 2983 5960 3017
rect 4360 2960 5960 2983
rect 6280 3017 7880 3040
rect 6280 2983 6307 3017
rect 6349 2983 6379 3017
rect 6417 2983 6451 3017
rect 6485 2983 6519 3017
rect 6557 2983 6587 3017
rect 6629 2983 6655 3017
rect 6701 2983 6723 3017
rect 6773 2983 6791 3017
rect 6845 2983 6859 3017
rect 6917 2983 6927 3017
rect 6989 2983 6995 3017
rect 7061 2983 7063 3017
rect 7097 2983 7099 3017
rect 7165 2983 7171 3017
rect 7233 2983 7243 3017
rect 7301 2983 7315 3017
rect 7369 2983 7387 3017
rect 7437 2983 7459 3017
rect 7505 2983 7531 3017
rect 7573 2983 7603 3017
rect 7641 2983 7675 3017
rect 7709 2983 7743 3017
rect 7781 2983 7811 3017
rect 7853 2983 7880 3017
rect 6280 2960 7880 2983
rect 8160 3031 8240 3065
rect 8160 2997 8183 3031
rect 8217 2997 8240 3031
rect 8160 2963 8240 2997
rect 160 2880 240 2929
rect 8160 2929 8183 2963
rect 8217 2929 8240 2963
rect 8160 2880 8240 2929
rect 160 2857 8240 2880
rect 160 2823 307 2857
rect 341 2823 375 2857
rect 409 2823 443 2857
rect 477 2823 511 2857
rect 545 2823 579 2857
rect 613 2823 647 2857
rect 681 2823 715 2857
rect 749 2823 783 2857
rect 817 2823 851 2857
rect 885 2823 919 2857
rect 953 2823 987 2857
rect 1021 2823 1055 2857
rect 1089 2823 1123 2857
rect 1157 2823 1191 2857
rect 1225 2823 1259 2857
rect 1293 2823 1327 2857
rect 1361 2823 1395 2857
rect 1429 2823 1463 2857
rect 1497 2823 1531 2857
rect 1565 2823 1599 2857
rect 1633 2823 1667 2857
rect 1701 2823 1735 2857
rect 1769 2823 1803 2857
rect 1837 2823 1871 2857
rect 1905 2823 1939 2857
rect 1973 2823 2007 2857
rect 2041 2823 2075 2857
rect 2109 2823 2143 2857
rect 2177 2823 2211 2857
rect 2245 2823 2279 2857
rect 2313 2823 2347 2857
rect 2381 2823 2415 2857
rect 2449 2823 2483 2857
rect 2517 2823 2551 2857
rect 2585 2823 2619 2857
rect 2653 2823 2687 2857
rect 2721 2823 2755 2857
rect 2789 2823 2823 2857
rect 2857 2823 2891 2857
rect 2925 2823 2959 2857
rect 2993 2823 3027 2857
rect 3061 2823 3095 2857
rect 3129 2823 3163 2857
rect 3197 2823 3231 2857
rect 3265 2823 3299 2857
rect 3333 2823 3367 2857
rect 3401 2823 3435 2857
rect 3469 2823 3503 2857
rect 3537 2823 3571 2857
rect 3605 2823 3639 2857
rect 3673 2823 3707 2857
rect 3741 2823 3775 2857
rect 3809 2823 3843 2857
rect 3877 2823 3911 2857
rect 3945 2823 3979 2857
rect 4013 2823 4047 2857
rect 4081 2823 4115 2857
rect 4149 2823 4183 2857
rect 4217 2823 4251 2857
rect 4285 2823 4319 2857
rect 4353 2823 4387 2857
rect 4421 2823 4455 2857
rect 4489 2823 4523 2857
rect 4557 2823 4591 2857
rect 4625 2823 4659 2857
rect 4693 2823 4727 2857
rect 4761 2823 4795 2857
rect 4829 2823 4863 2857
rect 4897 2823 4931 2857
rect 4965 2823 4999 2857
rect 5033 2823 5067 2857
rect 5101 2823 5135 2857
rect 5169 2823 5203 2857
rect 5237 2823 5271 2857
rect 5305 2823 5339 2857
rect 5373 2823 5407 2857
rect 5441 2823 5475 2857
rect 5509 2823 5543 2857
rect 5577 2823 5611 2857
rect 5645 2823 5679 2857
rect 5713 2823 5747 2857
rect 5781 2823 5815 2857
rect 5849 2823 5883 2857
rect 5917 2823 5951 2857
rect 5985 2823 6019 2857
rect 6053 2823 6087 2857
rect 6121 2823 6155 2857
rect 6189 2823 6223 2857
rect 6257 2823 6291 2857
rect 6325 2823 6359 2857
rect 6393 2823 6427 2857
rect 6461 2823 6495 2857
rect 6529 2823 6563 2857
rect 6597 2823 6631 2857
rect 6665 2823 6699 2857
rect 6733 2823 6767 2857
rect 6801 2823 6835 2857
rect 6869 2823 6903 2857
rect 6937 2823 6971 2857
rect 7005 2823 7039 2857
rect 7073 2823 7107 2857
rect 7141 2823 7175 2857
rect 7209 2823 7243 2857
rect 7277 2823 7311 2857
rect 7345 2823 7379 2857
rect 7413 2823 7447 2857
rect 7481 2823 7515 2857
rect 7549 2823 7583 2857
rect 7617 2823 7651 2857
rect 7685 2823 7719 2857
rect 7753 2823 7787 2857
rect 7821 2823 7855 2857
rect 7889 2823 7923 2857
rect 7957 2823 7991 2857
rect 8025 2823 8059 2857
rect 8093 2823 8240 2857
rect 160 2800 8240 2823
rect 8320 3813 8343 3847
rect 8377 3813 8400 3847
rect 8320 3779 8400 3813
rect 8320 3745 8343 3779
rect 8377 3745 8400 3779
rect 8320 3711 8400 3745
rect 8320 3677 8343 3711
rect 8377 3677 8400 3711
rect 8320 3643 8400 3677
rect 8320 3609 8343 3643
rect 8377 3609 8400 3643
rect 8320 3575 8400 3609
rect 8320 3541 8343 3575
rect 8377 3541 8400 3575
rect 8320 3507 8400 3541
rect 8320 3473 8343 3507
rect 8377 3473 8400 3507
rect 8320 3439 8400 3473
rect 8320 3405 8343 3439
rect 8377 3405 8400 3439
rect 8320 3371 8400 3405
rect 8320 3337 8343 3371
rect 8377 3337 8400 3371
rect 8320 3303 8400 3337
rect 8320 3269 8343 3303
rect 8377 3269 8400 3303
rect 8320 3235 8400 3269
rect 8320 3201 8343 3235
rect 8377 3201 8400 3235
rect 8320 3167 8400 3201
rect 8320 3133 8343 3167
rect 8377 3133 8400 3167
rect 8320 3099 8400 3133
rect 8320 3065 8343 3099
rect 8377 3065 8400 3099
rect 8320 3031 8400 3065
rect 8320 2997 8343 3031
rect 8377 2997 8400 3031
rect 8320 2963 8400 2997
rect 8320 2929 8343 2963
rect 8377 2929 8400 2963
rect 8320 2895 8400 2929
rect 8320 2861 8343 2895
rect 8377 2861 8400 2895
rect 8320 2827 8400 2861
rect 0 2720 80 2793
rect 8320 2793 8343 2827
rect 8377 2793 8400 2827
rect 8320 2720 8400 2793
rect 0 2697 8400 2720
rect 0 2663 151 2697
rect 185 2663 219 2697
rect 253 2663 287 2697
rect 321 2663 355 2697
rect 389 2663 423 2697
rect 457 2663 491 2697
rect 525 2663 559 2697
rect 593 2663 627 2697
rect 661 2663 695 2697
rect 729 2663 763 2697
rect 797 2663 831 2697
rect 865 2663 899 2697
rect 933 2663 967 2697
rect 1001 2663 1035 2697
rect 1069 2663 1103 2697
rect 1137 2663 1171 2697
rect 1205 2663 1239 2697
rect 1273 2663 1307 2697
rect 1341 2663 1375 2697
rect 1409 2663 1443 2697
rect 1477 2663 1511 2697
rect 1545 2663 1579 2697
rect 1613 2663 1647 2697
rect 1681 2663 1715 2697
rect 1749 2663 1783 2697
rect 1817 2663 1851 2697
rect 1885 2663 1919 2697
rect 1953 2663 1987 2697
rect 2021 2663 2055 2697
rect 2089 2663 2123 2697
rect 2157 2663 2191 2697
rect 2225 2663 2259 2697
rect 2293 2663 2327 2697
rect 2361 2663 2395 2697
rect 2429 2663 2463 2697
rect 2497 2663 2531 2697
rect 2565 2663 2599 2697
rect 2633 2663 2667 2697
rect 2701 2663 2735 2697
rect 2769 2663 2803 2697
rect 2837 2663 2871 2697
rect 2905 2663 2939 2697
rect 2973 2663 3007 2697
rect 3041 2663 3075 2697
rect 3109 2663 3143 2697
rect 3177 2663 3211 2697
rect 3245 2663 3279 2697
rect 3313 2663 3347 2697
rect 3381 2663 3415 2697
rect 3449 2663 3483 2697
rect 3517 2663 3551 2697
rect 3585 2663 3619 2697
rect 3653 2663 3687 2697
rect 3721 2663 3755 2697
rect 3789 2663 3823 2697
rect 3857 2663 3891 2697
rect 3925 2663 3959 2697
rect 3993 2663 4027 2697
rect 4061 2663 4095 2697
rect 4129 2663 4163 2697
rect 4197 2663 4231 2697
rect 4265 2663 4299 2697
rect 4333 2663 4367 2697
rect 4401 2663 4435 2697
rect 4469 2663 4503 2697
rect 4537 2663 4571 2697
rect 4605 2663 4639 2697
rect 4673 2663 4707 2697
rect 4741 2663 4775 2697
rect 4809 2663 4843 2697
rect 4877 2663 4911 2697
rect 4945 2663 4979 2697
rect 5013 2663 5047 2697
rect 5081 2663 5115 2697
rect 5149 2663 5183 2697
rect 5217 2663 5251 2697
rect 5285 2663 5319 2697
rect 5353 2663 5387 2697
rect 5421 2663 5455 2697
rect 5489 2663 5523 2697
rect 5557 2663 5591 2697
rect 5625 2663 5659 2697
rect 5693 2663 5727 2697
rect 5761 2663 5795 2697
rect 5829 2663 5863 2697
rect 5897 2663 5931 2697
rect 5965 2663 5999 2697
rect 6033 2663 6067 2697
rect 6101 2663 6135 2697
rect 6169 2663 6203 2697
rect 6237 2663 6271 2697
rect 6305 2663 6339 2697
rect 6373 2663 6407 2697
rect 6441 2663 6475 2697
rect 6509 2663 6543 2697
rect 6577 2663 6611 2697
rect 6645 2663 6679 2697
rect 6713 2663 6747 2697
rect 6781 2663 6815 2697
rect 6849 2663 6883 2697
rect 6917 2663 6951 2697
rect 6985 2663 7019 2697
rect 7053 2663 7087 2697
rect 7121 2663 7155 2697
rect 7189 2663 7223 2697
rect 7257 2663 7291 2697
rect 7325 2663 7359 2697
rect 7393 2663 7427 2697
rect 7461 2663 7495 2697
rect 7529 2663 7563 2697
rect 7597 2663 7631 2697
rect 7665 2663 7699 2697
rect 7733 2663 7767 2697
rect 7801 2663 7835 2697
rect 7869 2663 7903 2697
rect 7937 2663 7971 2697
rect 8005 2663 8039 2697
rect 8073 2663 8107 2697
rect 8141 2663 8175 2697
rect 8209 2663 8400 2697
rect 0 2640 8400 2663
rect 0 2560 80 2640
rect 8320 2560 8400 2640
rect 0 2537 8400 2560
rect 0 2503 151 2537
rect 185 2503 219 2537
rect 253 2503 287 2537
rect 321 2503 355 2537
rect 389 2503 423 2537
rect 457 2503 491 2537
rect 525 2503 559 2537
rect 593 2503 627 2537
rect 661 2503 695 2537
rect 729 2503 763 2537
rect 797 2503 831 2537
rect 865 2503 899 2537
rect 933 2503 967 2537
rect 1001 2503 1035 2537
rect 1069 2503 1103 2537
rect 1137 2503 1171 2537
rect 1205 2503 1239 2537
rect 1273 2503 1307 2537
rect 1341 2503 1375 2537
rect 1409 2503 1443 2537
rect 1477 2503 1511 2537
rect 1545 2503 1579 2537
rect 1613 2503 1647 2537
rect 1681 2503 1715 2537
rect 1749 2503 1783 2537
rect 1817 2503 1851 2537
rect 1885 2503 1919 2537
rect 1953 2503 1987 2537
rect 2021 2503 2055 2537
rect 2089 2503 2123 2537
rect 2157 2503 2191 2537
rect 2225 2503 2259 2537
rect 2293 2503 2327 2537
rect 2361 2503 2395 2537
rect 2429 2503 2463 2537
rect 2497 2503 2531 2537
rect 2565 2503 2599 2537
rect 2633 2503 2667 2537
rect 2701 2503 2735 2537
rect 2769 2503 2803 2537
rect 2837 2503 2871 2537
rect 2905 2503 2939 2537
rect 2973 2503 3007 2537
rect 3041 2503 3075 2537
rect 3109 2503 3143 2537
rect 3177 2503 3211 2537
rect 3245 2503 3279 2537
rect 3313 2503 3347 2537
rect 3381 2503 3415 2537
rect 3449 2503 3483 2537
rect 3517 2503 3551 2537
rect 3585 2503 3619 2537
rect 3653 2503 3687 2537
rect 3721 2503 3755 2537
rect 3789 2503 3823 2537
rect 3857 2503 3891 2537
rect 3925 2503 3959 2537
rect 3993 2503 4027 2537
rect 4061 2503 4095 2537
rect 4129 2503 4163 2537
rect 4197 2503 4231 2537
rect 4265 2503 4299 2537
rect 4333 2503 4367 2537
rect 4401 2503 4435 2537
rect 4469 2503 4503 2537
rect 4537 2503 4571 2537
rect 4605 2503 4639 2537
rect 4673 2503 4707 2537
rect 4741 2503 4775 2537
rect 4809 2503 4843 2537
rect 4877 2503 4911 2537
rect 4945 2503 4979 2537
rect 5013 2503 5047 2537
rect 5081 2503 5115 2537
rect 5149 2503 5183 2537
rect 5217 2503 5251 2537
rect 5285 2503 5319 2537
rect 5353 2503 5387 2537
rect 5421 2503 5455 2537
rect 5489 2503 5523 2537
rect 5557 2503 5591 2537
rect 5625 2503 5659 2537
rect 5693 2503 5727 2537
rect 5761 2503 5795 2537
rect 5829 2503 5863 2537
rect 5897 2503 5931 2537
rect 5965 2503 5999 2537
rect 6033 2503 6067 2537
rect 6101 2503 6135 2537
rect 6169 2503 6203 2537
rect 6237 2503 6271 2537
rect 6305 2503 6339 2537
rect 6373 2503 6407 2537
rect 6441 2503 6475 2537
rect 6509 2503 6543 2537
rect 6577 2503 6611 2537
rect 6645 2503 6679 2537
rect 6713 2503 6747 2537
rect 6781 2503 6815 2537
rect 6849 2503 6883 2537
rect 6917 2503 6951 2537
rect 6985 2503 7019 2537
rect 7053 2503 7087 2537
rect 7121 2503 7155 2537
rect 7189 2503 7223 2537
rect 7257 2503 7291 2537
rect 7325 2503 7359 2537
rect 7393 2503 7427 2537
rect 7461 2503 7495 2537
rect 7529 2503 7563 2537
rect 7597 2503 7631 2537
rect 7665 2503 7699 2537
rect 7733 2503 7767 2537
rect 7801 2503 7835 2537
rect 7869 2503 7903 2537
rect 7937 2503 7971 2537
rect 8005 2503 8039 2537
rect 8073 2503 8107 2537
rect 8141 2503 8175 2537
rect 8209 2503 8400 2537
rect 0 2480 8400 2503
rect 0 2407 80 2480
rect 0 2373 23 2407
rect 57 2373 80 2407
rect 8320 2419 8400 2480
rect 0 2339 80 2373
rect 0 2305 23 2339
rect 57 2305 80 2339
rect 0 2271 80 2305
rect 0 2237 23 2271
rect 57 2237 80 2271
rect 0 2203 80 2237
rect 0 2169 23 2203
rect 57 2169 80 2203
rect 0 2135 80 2169
rect 0 2101 23 2135
rect 57 2101 80 2135
rect 0 2067 80 2101
rect 0 2033 23 2067
rect 57 2033 80 2067
rect 0 1999 80 2033
rect 0 1965 23 1999
rect 57 1965 80 1999
rect 0 1931 80 1965
rect 0 1897 23 1931
rect 57 1897 80 1931
rect 0 1863 80 1897
rect 0 1829 23 1863
rect 57 1829 80 1863
rect 0 1795 80 1829
rect 0 1761 23 1795
rect 57 1761 80 1795
rect 0 1727 80 1761
rect 0 1693 23 1727
rect 57 1693 80 1727
rect 0 1659 80 1693
rect 0 1625 23 1659
rect 57 1625 80 1659
rect 0 1591 80 1625
rect 0 1557 23 1591
rect 57 1557 80 1591
rect 0 1523 80 1557
rect 0 1489 23 1523
rect 57 1489 80 1523
rect 0 1455 80 1489
rect 0 1421 23 1455
rect 57 1421 80 1455
rect 0 1387 80 1421
rect 0 1353 23 1387
rect 57 1353 80 1387
rect 160 2377 8240 2400
rect 160 2343 307 2377
rect 341 2343 375 2377
rect 409 2343 443 2377
rect 477 2343 511 2377
rect 545 2343 579 2377
rect 613 2343 647 2377
rect 681 2343 715 2377
rect 749 2343 783 2377
rect 817 2343 851 2377
rect 885 2343 919 2377
rect 953 2343 987 2377
rect 1021 2343 1055 2377
rect 1089 2343 1123 2377
rect 1157 2343 1191 2377
rect 1225 2343 1259 2377
rect 1293 2343 1327 2377
rect 1361 2343 1395 2377
rect 1429 2343 1463 2377
rect 1497 2343 1531 2377
rect 1565 2343 1599 2377
rect 1633 2343 1667 2377
rect 1701 2343 1735 2377
rect 1769 2343 1803 2377
rect 1837 2343 1871 2377
rect 1905 2343 1939 2377
rect 1973 2343 2007 2377
rect 2041 2343 2075 2377
rect 2109 2343 2143 2377
rect 2177 2343 2211 2377
rect 2245 2343 2279 2377
rect 2313 2343 2347 2377
rect 2381 2343 2415 2377
rect 2449 2343 2483 2377
rect 2517 2343 2551 2377
rect 2585 2343 2619 2377
rect 2653 2343 2687 2377
rect 2721 2343 2755 2377
rect 2789 2343 2823 2377
rect 2857 2343 2891 2377
rect 2925 2343 2959 2377
rect 2993 2343 3027 2377
rect 3061 2343 3095 2377
rect 3129 2343 3163 2377
rect 3197 2343 3231 2377
rect 3265 2343 3299 2377
rect 3333 2343 3367 2377
rect 3401 2343 3435 2377
rect 3469 2343 3503 2377
rect 3537 2343 3571 2377
rect 3605 2343 3639 2377
rect 3673 2343 3707 2377
rect 3741 2343 3775 2377
rect 3809 2343 3843 2377
rect 3877 2343 3911 2377
rect 3945 2343 3979 2377
rect 4013 2343 4047 2377
rect 4081 2343 4115 2377
rect 4149 2343 4183 2377
rect 4217 2343 4251 2377
rect 4285 2343 4319 2377
rect 4353 2343 4387 2377
rect 4421 2343 4455 2377
rect 4489 2343 4523 2377
rect 4557 2343 4591 2377
rect 4625 2343 4659 2377
rect 4693 2343 4727 2377
rect 4761 2343 4795 2377
rect 4829 2343 4863 2377
rect 4897 2343 4931 2377
rect 4965 2343 4999 2377
rect 5033 2343 5067 2377
rect 5101 2343 5135 2377
rect 5169 2343 5203 2377
rect 5237 2343 5271 2377
rect 5305 2343 5339 2377
rect 5373 2343 5407 2377
rect 5441 2343 5475 2377
rect 5509 2343 5543 2377
rect 5577 2343 5611 2377
rect 5645 2343 5679 2377
rect 5713 2343 5747 2377
rect 5781 2343 5815 2377
rect 5849 2343 5883 2377
rect 5917 2343 5951 2377
rect 5985 2343 6019 2377
rect 6053 2343 6087 2377
rect 6121 2343 6155 2377
rect 6189 2343 6223 2377
rect 6257 2343 6291 2377
rect 6325 2343 6359 2377
rect 6393 2343 6427 2377
rect 6461 2343 6495 2377
rect 6529 2343 6563 2377
rect 6597 2343 6631 2377
rect 6665 2343 6699 2377
rect 6733 2343 6767 2377
rect 6801 2343 6835 2377
rect 6869 2343 6903 2377
rect 6937 2343 6971 2377
rect 7005 2343 7039 2377
rect 7073 2343 7107 2377
rect 7141 2343 7175 2377
rect 7209 2343 7243 2377
rect 7277 2343 7311 2377
rect 7345 2343 7379 2377
rect 7413 2343 7447 2377
rect 7481 2343 7515 2377
rect 7549 2343 7583 2377
rect 7617 2343 7651 2377
rect 7685 2343 7719 2377
rect 7753 2343 7787 2377
rect 7821 2343 7855 2377
rect 7889 2343 7923 2377
rect 7957 2343 7991 2377
rect 8025 2343 8059 2377
rect 8093 2343 8240 2377
rect 160 2320 8240 2343
rect 160 2271 240 2320
rect 160 2237 183 2271
rect 217 2237 240 2271
rect 160 2203 240 2237
rect 160 2169 183 2203
rect 217 2169 240 2203
rect 160 2135 240 2169
rect 160 2101 183 2135
rect 217 2101 240 2135
rect 160 2067 240 2101
rect 160 2033 183 2067
rect 217 2033 240 2067
rect 160 1999 240 2033
rect 160 1965 183 1999
rect 217 1965 240 1999
rect 160 1931 240 1965
rect 160 1897 183 1931
rect 217 1897 240 1931
rect 160 1863 240 1897
rect 160 1829 183 1863
rect 217 1829 240 1863
rect 160 1795 240 1829
rect 160 1761 183 1795
rect 217 1761 240 1795
rect 160 1727 240 1761
rect 160 1693 183 1727
rect 217 1693 240 1727
rect 160 1659 240 1693
rect 160 1625 183 1659
rect 217 1625 240 1659
rect 320 2209 400 2320
rect 8160 2271 8240 2320
rect 320 2161 343 2209
rect 377 2161 400 2209
rect 320 2137 400 2161
rect 320 2093 343 2137
rect 377 2093 400 2137
rect 320 2065 400 2093
rect 320 2025 343 2065
rect 377 2025 400 2065
rect 320 1993 400 2025
rect 320 1957 343 1993
rect 377 1957 400 1993
rect 320 1923 400 1957
rect 320 1887 343 1923
rect 377 1887 400 1923
rect 320 1855 400 1887
rect 320 1815 343 1855
rect 377 1815 400 1855
rect 320 1787 400 1815
rect 320 1743 343 1787
rect 377 1743 400 1787
rect 320 1719 400 1743
rect 320 1671 343 1719
rect 377 1671 400 1719
rect 320 1640 400 1671
rect 2240 2209 2320 2240
rect 2240 2161 2263 2209
rect 2297 2161 2320 2209
rect 2240 2137 2320 2161
rect 2240 2093 2263 2137
rect 2297 2093 2320 2137
rect 2240 2065 2320 2093
rect 2240 2025 2263 2065
rect 2297 2025 2320 2065
rect 2240 1993 2320 2025
rect 2240 1957 2263 1993
rect 2297 1957 2320 1993
rect 2240 1923 2320 1957
rect 2240 1887 2263 1923
rect 2297 1887 2320 1923
rect 2240 1855 2320 1887
rect 2240 1815 2263 1855
rect 2297 1815 2320 1855
rect 2240 1787 2320 1815
rect 2240 1743 2263 1787
rect 2297 1743 2320 1787
rect 2240 1719 2320 1743
rect 2240 1671 2263 1719
rect 2297 1671 2320 1719
rect 2240 1640 2320 1671
rect 4160 2209 4240 2240
rect 4160 2161 4183 2209
rect 4217 2161 4240 2209
rect 4160 2137 4240 2161
rect 4160 2093 4183 2137
rect 4217 2093 4240 2137
rect 4160 2065 4240 2093
rect 4160 2025 4183 2065
rect 4217 2025 4240 2065
rect 4160 1993 4240 2025
rect 4160 1957 4183 1993
rect 4217 1957 4240 1993
rect 4160 1923 4240 1957
rect 4160 1887 4183 1923
rect 4217 1887 4240 1923
rect 4160 1855 4240 1887
rect 4160 1815 4183 1855
rect 4217 1815 4240 1855
rect 4160 1787 4240 1815
rect 4160 1743 4183 1787
rect 4217 1743 4240 1787
rect 4160 1719 4240 1743
rect 4160 1671 4183 1719
rect 4217 1671 4240 1719
rect 4160 1640 4240 1671
rect 6080 2209 6160 2240
rect 6080 2161 6103 2209
rect 6137 2161 6160 2209
rect 6080 2137 6160 2161
rect 6080 2093 6103 2137
rect 6137 2093 6160 2137
rect 6080 2065 6160 2093
rect 6080 2025 6103 2065
rect 6137 2025 6160 2065
rect 6080 1993 6160 2025
rect 6080 1957 6103 1993
rect 6137 1957 6160 1993
rect 6080 1923 6160 1957
rect 6080 1887 6103 1923
rect 6137 1887 6160 1923
rect 6080 1855 6160 1887
rect 6080 1815 6103 1855
rect 6137 1815 6160 1855
rect 6080 1787 6160 1815
rect 6080 1743 6103 1787
rect 6137 1743 6160 1787
rect 6080 1719 6160 1743
rect 6080 1671 6103 1719
rect 6137 1671 6160 1719
rect 6080 1640 6160 1671
rect 8000 2209 8080 2240
rect 8000 2161 8023 2209
rect 8057 2161 8080 2209
rect 8000 2137 8080 2161
rect 8000 2093 8023 2137
rect 8057 2093 8080 2137
rect 8000 2065 8080 2093
rect 8000 2025 8023 2065
rect 8057 2025 8080 2065
rect 8000 1993 8080 2025
rect 8000 1957 8023 1993
rect 8057 1957 8080 1993
rect 8000 1923 8080 1957
rect 8000 1887 8023 1923
rect 8057 1887 8080 1923
rect 8000 1855 8080 1887
rect 8000 1815 8023 1855
rect 8057 1815 8080 1855
rect 8000 1787 8080 1815
rect 8000 1743 8023 1787
rect 8057 1743 8080 1787
rect 8000 1719 8080 1743
rect 8000 1671 8023 1719
rect 8057 1671 8080 1719
rect 8000 1640 8080 1671
rect 8160 2237 8183 2271
rect 8217 2237 8240 2271
rect 8160 2203 8240 2237
rect 8160 2169 8183 2203
rect 8217 2169 8240 2203
rect 8160 2135 8240 2169
rect 8160 2101 8183 2135
rect 8217 2101 8240 2135
rect 8160 2067 8240 2101
rect 8160 2033 8183 2067
rect 8217 2033 8240 2067
rect 8160 1999 8240 2033
rect 8160 1965 8183 1999
rect 8217 1965 8240 1999
rect 8160 1931 8240 1965
rect 8160 1897 8183 1931
rect 8217 1897 8240 1931
rect 8160 1863 8240 1897
rect 8160 1829 8183 1863
rect 8217 1829 8240 1863
rect 8160 1795 8240 1829
rect 8160 1761 8183 1795
rect 8217 1761 8240 1795
rect 8160 1727 8240 1761
rect 8160 1693 8183 1727
rect 8217 1693 8240 1727
rect 8160 1659 8240 1693
rect 160 1591 240 1625
rect 8160 1625 8183 1659
rect 8217 1625 8240 1659
rect 160 1557 183 1591
rect 217 1557 240 1591
rect 160 1523 240 1557
rect 160 1489 183 1523
rect 217 1489 240 1523
rect 520 1577 2120 1600
rect 520 1543 547 1577
rect 589 1543 619 1577
rect 657 1543 691 1577
rect 725 1543 759 1577
rect 797 1543 827 1577
rect 869 1543 895 1577
rect 941 1543 963 1577
rect 1013 1543 1031 1577
rect 1085 1543 1099 1577
rect 1157 1543 1167 1577
rect 1229 1543 1235 1577
rect 1301 1543 1303 1577
rect 1337 1543 1339 1577
rect 1405 1543 1411 1577
rect 1473 1543 1483 1577
rect 1541 1543 1555 1577
rect 1609 1543 1627 1577
rect 1677 1543 1699 1577
rect 1745 1543 1771 1577
rect 1813 1543 1843 1577
rect 1881 1543 1915 1577
rect 1949 1543 1983 1577
rect 2021 1543 2051 1577
rect 2093 1543 2120 1577
rect 520 1520 2120 1543
rect 2440 1577 4040 1600
rect 2440 1543 2467 1577
rect 2509 1543 2539 1577
rect 2577 1543 2611 1577
rect 2645 1543 2679 1577
rect 2717 1543 2747 1577
rect 2789 1543 2815 1577
rect 2861 1543 2883 1577
rect 2933 1543 2951 1577
rect 3005 1543 3019 1577
rect 3077 1543 3087 1577
rect 3149 1543 3155 1577
rect 3221 1543 3223 1577
rect 3257 1543 3259 1577
rect 3325 1543 3331 1577
rect 3393 1543 3403 1577
rect 3461 1543 3475 1577
rect 3529 1543 3547 1577
rect 3597 1543 3619 1577
rect 3665 1543 3691 1577
rect 3733 1543 3763 1577
rect 3801 1543 3835 1577
rect 3869 1543 3903 1577
rect 3941 1543 3971 1577
rect 4013 1543 4040 1577
rect 2440 1520 4040 1543
rect 4360 1577 5960 1600
rect 4360 1543 4387 1577
rect 4429 1543 4459 1577
rect 4497 1543 4531 1577
rect 4565 1543 4599 1577
rect 4637 1543 4667 1577
rect 4709 1543 4735 1577
rect 4781 1543 4803 1577
rect 4853 1543 4871 1577
rect 4925 1543 4939 1577
rect 4997 1543 5007 1577
rect 5069 1543 5075 1577
rect 5141 1543 5143 1577
rect 5177 1543 5179 1577
rect 5245 1543 5251 1577
rect 5313 1543 5323 1577
rect 5381 1543 5395 1577
rect 5449 1543 5467 1577
rect 5517 1543 5539 1577
rect 5585 1543 5611 1577
rect 5653 1543 5683 1577
rect 5721 1543 5755 1577
rect 5789 1543 5823 1577
rect 5861 1543 5891 1577
rect 5933 1543 5960 1577
rect 4360 1520 5960 1543
rect 6280 1577 7880 1600
rect 6280 1543 6307 1577
rect 6349 1543 6379 1577
rect 6417 1543 6451 1577
rect 6485 1543 6519 1577
rect 6557 1543 6587 1577
rect 6629 1543 6655 1577
rect 6701 1543 6723 1577
rect 6773 1543 6791 1577
rect 6845 1543 6859 1577
rect 6917 1543 6927 1577
rect 6989 1543 6995 1577
rect 7061 1543 7063 1577
rect 7097 1543 7099 1577
rect 7165 1543 7171 1577
rect 7233 1543 7243 1577
rect 7301 1543 7315 1577
rect 7369 1543 7387 1577
rect 7437 1543 7459 1577
rect 7505 1543 7531 1577
rect 7573 1543 7603 1577
rect 7641 1543 7675 1577
rect 7709 1543 7743 1577
rect 7781 1543 7811 1577
rect 7853 1543 7880 1577
rect 6280 1520 7880 1543
rect 8160 1591 8240 1625
rect 8160 1557 8183 1591
rect 8217 1557 8240 1591
rect 8160 1523 8240 1557
rect 160 1440 240 1489
rect 8160 1489 8183 1523
rect 8217 1489 8240 1523
rect 8160 1440 8240 1489
rect 160 1417 8240 1440
rect 160 1383 307 1417
rect 341 1383 375 1417
rect 409 1383 443 1417
rect 477 1383 511 1417
rect 545 1383 579 1417
rect 613 1383 647 1417
rect 681 1383 715 1417
rect 749 1383 783 1417
rect 817 1383 851 1417
rect 885 1383 919 1417
rect 953 1383 987 1417
rect 1021 1383 1055 1417
rect 1089 1383 1123 1417
rect 1157 1383 1191 1417
rect 1225 1383 1259 1417
rect 1293 1383 1327 1417
rect 1361 1383 1395 1417
rect 1429 1383 1463 1417
rect 1497 1383 1531 1417
rect 1565 1383 1599 1417
rect 1633 1383 1667 1417
rect 1701 1383 1735 1417
rect 1769 1383 1803 1417
rect 1837 1383 1871 1417
rect 1905 1383 1939 1417
rect 1973 1383 2007 1417
rect 2041 1383 2075 1417
rect 2109 1383 2143 1417
rect 2177 1383 2211 1417
rect 2245 1383 2279 1417
rect 2313 1383 2347 1417
rect 2381 1383 2415 1417
rect 2449 1383 2483 1417
rect 2517 1383 2551 1417
rect 2585 1383 2619 1417
rect 2653 1383 2687 1417
rect 2721 1383 2755 1417
rect 2789 1383 2823 1417
rect 2857 1383 2891 1417
rect 2925 1383 2959 1417
rect 2993 1383 3027 1417
rect 3061 1383 3095 1417
rect 3129 1383 3163 1417
rect 3197 1383 3231 1417
rect 3265 1383 3299 1417
rect 3333 1383 3367 1417
rect 3401 1383 3435 1417
rect 3469 1383 3503 1417
rect 3537 1383 3571 1417
rect 3605 1383 3639 1417
rect 3673 1383 3707 1417
rect 3741 1383 3775 1417
rect 3809 1383 3843 1417
rect 3877 1383 3911 1417
rect 3945 1383 3979 1417
rect 4013 1383 4047 1417
rect 4081 1383 4115 1417
rect 4149 1383 4183 1417
rect 4217 1383 4251 1417
rect 4285 1383 4319 1417
rect 4353 1383 4387 1417
rect 4421 1383 4455 1417
rect 4489 1383 4523 1417
rect 4557 1383 4591 1417
rect 4625 1383 4659 1417
rect 4693 1383 4727 1417
rect 4761 1383 4795 1417
rect 4829 1383 4863 1417
rect 4897 1383 4931 1417
rect 4965 1383 4999 1417
rect 5033 1383 5067 1417
rect 5101 1383 5135 1417
rect 5169 1383 5203 1417
rect 5237 1383 5271 1417
rect 5305 1383 5339 1417
rect 5373 1383 5407 1417
rect 5441 1383 5475 1417
rect 5509 1383 5543 1417
rect 5577 1383 5611 1417
rect 5645 1383 5679 1417
rect 5713 1383 5747 1417
rect 5781 1383 5815 1417
rect 5849 1383 5883 1417
rect 5917 1383 5951 1417
rect 5985 1383 6019 1417
rect 6053 1383 6087 1417
rect 6121 1383 6155 1417
rect 6189 1383 6223 1417
rect 6257 1383 6291 1417
rect 6325 1383 6359 1417
rect 6393 1383 6427 1417
rect 6461 1383 6495 1417
rect 6529 1383 6563 1417
rect 6597 1383 6631 1417
rect 6665 1383 6699 1417
rect 6733 1383 6767 1417
rect 6801 1383 6835 1417
rect 6869 1383 6903 1417
rect 6937 1383 6971 1417
rect 7005 1383 7039 1417
rect 7073 1383 7107 1417
rect 7141 1383 7175 1417
rect 7209 1383 7243 1417
rect 7277 1383 7311 1417
rect 7345 1383 7379 1417
rect 7413 1383 7447 1417
rect 7481 1383 7515 1417
rect 7549 1383 7583 1417
rect 7617 1383 7651 1417
rect 7685 1383 7719 1417
rect 7753 1383 7787 1417
rect 7821 1383 7855 1417
rect 7889 1383 7923 1417
rect 7957 1383 7991 1417
rect 8025 1383 8059 1417
rect 8093 1383 8240 1417
rect 160 1360 8240 1383
rect 8320 2385 8343 2419
rect 8377 2385 8400 2419
rect 8320 2351 8400 2385
rect 8320 2317 8343 2351
rect 8377 2317 8400 2351
rect 8320 2283 8400 2317
rect 8320 2249 8343 2283
rect 8377 2249 8400 2283
rect 8320 2215 8400 2249
rect 8320 2181 8343 2215
rect 8377 2181 8400 2215
rect 8320 2147 8400 2181
rect 8320 2113 8343 2147
rect 8377 2113 8400 2147
rect 8320 2079 8400 2113
rect 8320 2045 8343 2079
rect 8377 2045 8400 2079
rect 8320 2011 8400 2045
rect 8320 1977 8343 2011
rect 8377 1977 8400 2011
rect 8320 1943 8400 1977
rect 8320 1909 8343 1943
rect 8377 1909 8400 1943
rect 8320 1875 8400 1909
rect 8320 1841 8343 1875
rect 8377 1841 8400 1875
rect 8320 1807 8400 1841
rect 8320 1773 8343 1807
rect 8377 1773 8400 1807
rect 8320 1739 8400 1773
rect 8320 1705 8343 1739
rect 8377 1705 8400 1739
rect 8320 1671 8400 1705
rect 8320 1637 8343 1671
rect 8377 1637 8400 1671
rect 8320 1603 8400 1637
rect 8320 1569 8343 1603
rect 8377 1569 8400 1603
rect 8320 1535 8400 1569
rect 8320 1501 8343 1535
rect 8377 1501 8400 1535
rect 8320 1467 8400 1501
rect 8320 1433 8343 1467
rect 8377 1433 8400 1467
rect 8320 1399 8400 1433
rect 8320 1365 8343 1399
rect 8377 1365 8400 1399
rect 0 1280 80 1353
rect 8320 1331 8400 1365
rect 8320 1297 8343 1331
rect 8377 1297 8400 1331
rect 8320 1280 8400 1297
rect 0 1263 8400 1280
rect 0 1257 8343 1263
rect 0 1223 137 1257
rect 171 1223 205 1257
rect 239 1223 273 1257
rect 307 1223 341 1257
rect 375 1223 409 1257
rect 443 1223 477 1257
rect 511 1223 545 1257
rect 579 1223 613 1257
rect 647 1223 681 1257
rect 715 1223 749 1257
rect 783 1223 817 1257
rect 851 1223 885 1257
rect 919 1223 953 1257
rect 987 1223 1021 1257
rect 1055 1223 1089 1257
rect 1123 1223 1157 1257
rect 1191 1223 1225 1257
rect 1259 1223 1293 1257
rect 1327 1223 1361 1257
rect 1395 1223 1429 1257
rect 1463 1223 1497 1257
rect 1531 1223 1565 1257
rect 1599 1223 1633 1257
rect 1667 1223 1701 1257
rect 1735 1223 1769 1257
rect 1803 1223 1837 1257
rect 1871 1223 1905 1257
rect 1939 1223 1973 1257
rect 2007 1223 2041 1257
rect 2075 1223 2109 1257
rect 2143 1223 2177 1257
rect 2211 1223 2245 1257
rect 2279 1223 2313 1257
rect 2347 1223 2381 1257
rect 2415 1223 2449 1257
rect 2483 1223 2517 1257
rect 2551 1223 2585 1257
rect 2619 1223 2653 1257
rect 2687 1223 2721 1257
rect 2755 1223 2789 1257
rect 2823 1223 2857 1257
rect 2891 1223 2925 1257
rect 2959 1223 2993 1257
rect 3027 1223 3061 1257
rect 3095 1223 3129 1257
rect 3163 1223 3197 1257
rect 3231 1223 3265 1257
rect 3299 1223 3333 1257
rect 3367 1223 3401 1257
rect 3435 1223 3469 1257
rect 3503 1223 3537 1257
rect 3571 1223 3605 1257
rect 3639 1223 3673 1257
rect 3707 1223 3741 1257
rect 3775 1223 3809 1257
rect 3843 1223 3877 1257
rect 3911 1223 3945 1257
rect 3979 1223 4013 1257
rect 4047 1223 4081 1257
rect 4115 1223 4149 1257
rect 4183 1223 4217 1257
rect 4251 1223 4285 1257
rect 4319 1223 4353 1257
rect 4387 1223 4421 1257
rect 4455 1223 4489 1257
rect 4523 1223 4557 1257
rect 4591 1223 4625 1257
rect 4659 1223 4693 1257
rect 4727 1223 4761 1257
rect 4795 1223 4829 1257
rect 4863 1223 4897 1257
rect 4931 1223 4965 1257
rect 4999 1223 5033 1257
rect 5067 1223 5101 1257
rect 5135 1223 5169 1257
rect 5203 1223 5237 1257
rect 5271 1223 5305 1257
rect 5339 1223 5373 1257
rect 5407 1223 5441 1257
rect 5475 1223 5509 1257
rect 5543 1223 5577 1257
rect 5611 1223 5645 1257
rect 5679 1223 5713 1257
rect 5747 1223 5781 1257
rect 5815 1223 5849 1257
rect 5883 1223 5917 1257
rect 5951 1223 5985 1257
rect 6019 1223 6053 1257
rect 6087 1223 6121 1257
rect 6155 1223 6189 1257
rect 6223 1223 6257 1257
rect 6291 1223 6325 1257
rect 6359 1223 6393 1257
rect 6427 1223 6461 1257
rect 6495 1223 6529 1257
rect 6563 1223 6597 1257
rect 6631 1223 6665 1257
rect 6699 1223 6733 1257
rect 6767 1223 6801 1257
rect 6835 1223 6869 1257
rect 6903 1223 6937 1257
rect 6971 1223 7005 1257
rect 7039 1223 7073 1257
rect 7107 1223 7141 1257
rect 7175 1223 7209 1257
rect 7243 1223 7277 1257
rect 7311 1223 7345 1257
rect 7379 1223 7413 1257
rect 7447 1223 7481 1257
rect 7515 1223 7549 1257
rect 7583 1223 7617 1257
rect 7651 1223 7685 1257
rect 7719 1223 7753 1257
rect 7787 1223 7821 1257
rect 7855 1223 7889 1257
rect 7923 1223 7957 1257
rect 7991 1223 8025 1257
rect 8059 1223 8093 1257
rect 8127 1223 8161 1257
rect 8195 1223 8229 1257
rect 8263 1229 8343 1257
rect 8377 1229 8400 1263
rect 8263 1223 8400 1229
rect 0 1200 8400 1223
rect 0 640 80 1200
rect 8320 1195 8400 1200
rect 8320 1161 8343 1195
rect 8377 1161 8400 1195
rect 8320 1127 8400 1161
rect 160 937 8240 1120
rect 160 903 183 937
rect 217 903 343 937
rect 377 903 503 937
rect 537 903 663 937
rect 697 903 823 937
rect 857 903 983 937
rect 1017 903 1143 937
rect 1177 903 1463 937
rect 1497 903 1623 937
rect 1657 903 1783 937
rect 1817 903 1943 937
rect 1977 903 2103 937
rect 2137 903 2263 937
rect 2297 903 2423 937
rect 2457 903 2583 937
rect 2617 903 2743 937
rect 2777 903 2903 937
rect 2937 903 3063 937
rect 3097 903 3383 937
rect 3417 903 3543 937
rect 3577 903 3703 937
rect 3737 903 3863 937
rect 3897 903 4023 937
rect 4057 903 4183 937
rect 4217 903 4343 937
rect 4377 903 4503 937
rect 4537 903 4663 937
rect 4697 903 4823 937
rect 4857 903 4983 937
rect 5017 903 5303 937
rect 5337 903 5463 937
rect 5497 903 5623 937
rect 5657 903 5783 937
rect 5817 903 5943 937
rect 5977 903 6103 937
rect 6137 903 6263 937
rect 6297 903 6423 937
rect 6457 903 6583 937
rect 6617 903 6743 937
rect 6777 903 6903 937
rect 6937 903 7223 937
rect 7257 903 7383 937
rect 7417 903 7543 937
rect 7577 903 7703 937
rect 7737 903 7863 937
rect 7897 903 8183 937
rect 8217 903 8240 937
rect 160 720 8240 903
rect 8320 1093 8343 1127
rect 8377 1093 8400 1127
rect 8320 1059 8400 1093
rect 8320 1025 8343 1059
rect 8377 1025 8400 1059
rect 8320 991 8400 1025
rect 8320 957 8343 991
rect 8377 957 8400 991
rect 8320 923 8400 957
rect 8320 889 8343 923
rect 8377 889 8400 923
rect 8320 855 8400 889
rect 8320 821 8343 855
rect 8377 821 8400 855
rect 8320 787 8400 821
rect 8320 753 8343 787
rect 8377 753 8400 787
rect 8320 719 8400 753
rect 8320 685 8343 719
rect 8377 685 8400 719
rect 8320 651 8400 685
rect 8320 640 8343 651
rect 0 617 8343 640
rect 8377 617 8400 651
rect 0 583 137 617
rect 171 583 205 617
rect 239 583 273 617
rect 307 583 341 617
rect 375 583 409 617
rect 443 583 477 617
rect 511 583 545 617
rect 579 583 613 617
rect 647 583 681 617
rect 715 583 749 617
rect 783 583 817 617
rect 851 583 885 617
rect 919 583 953 617
rect 987 583 1021 617
rect 1055 583 1089 617
rect 1123 583 1157 617
rect 1191 583 1225 617
rect 1259 583 1293 617
rect 1327 583 1361 617
rect 1395 583 1429 617
rect 1463 583 1497 617
rect 1531 583 1565 617
rect 1599 583 1633 617
rect 1667 583 1701 617
rect 1735 583 1769 617
rect 1803 583 1837 617
rect 1871 583 1905 617
rect 1939 583 1973 617
rect 2007 583 2041 617
rect 2075 583 2109 617
rect 2143 583 2177 617
rect 2211 583 2245 617
rect 2279 583 2313 617
rect 2347 583 2381 617
rect 2415 583 2449 617
rect 2483 583 2517 617
rect 2551 583 2585 617
rect 2619 583 2653 617
rect 2687 583 2721 617
rect 2755 583 2789 617
rect 2823 583 2857 617
rect 2891 583 2925 617
rect 2959 583 2993 617
rect 3027 583 3061 617
rect 3095 583 3129 617
rect 3163 583 3197 617
rect 3231 583 3265 617
rect 3299 583 3333 617
rect 3367 583 3401 617
rect 3435 583 3469 617
rect 3503 583 3537 617
rect 3571 583 3605 617
rect 3639 583 3673 617
rect 3707 583 3741 617
rect 3775 583 3809 617
rect 3843 583 3877 617
rect 3911 583 3945 617
rect 3979 583 4013 617
rect 4047 583 4081 617
rect 4115 583 4149 617
rect 4183 583 4217 617
rect 4251 583 4285 617
rect 4319 583 4353 617
rect 4387 583 4421 617
rect 4455 583 4489 617
rect 4523 583 4557 617
rect 4591 583 4625 617
rect 4659 583 4693 617
rect 4727 583 4761 617
rect 4795 583 4829 617
rect 4863 583 4897 617
rect 4931 583 4965 617
rect 4999 583 5033 617
rect 5067 583 5101 617
rect 5135 583 5169 617
rect 5203 583 5237 617
rect 5271 583 5305 617
rect 5339 583 5373 617
rect 5407 583 5441 617
rect 5475 583 5509 617
rect 5543 583 5577 617
rect 5611 583 5645 617
rect 5679 583 5713 617
rect 5747 583 5781 617
rect 5815 583 5849 617
rect 5883 583 5917 617
rect 5951 583 5985 617
rect 6019 583 6053 617
rect 6087 583 6121 617
rect 6155 583 6189 617
rect 6223 583 6257 617
rect 6291 583 6325 617
rect 6359 583 6393 617
rect 6427 583 6461 617
rect 6495 583 6529 617
rect 6563 583 6597 617
rect 6631 583 6665 617
rect 6699 583 6733 617
rect 6767 583 6801 617
rect 6835 583 6869 617
rect 6903 583 6937 617
rect 6971 583 7005 617
rect 7039 583 7073 617
rect 7107 583 7141 617
rect 7175 583 7209 617
rect 7243 583 7277 617
rect 7311 583 7345 617
rect 7379 583 7413 617
rect 7447 583 7481 617
rect 7515 583 7549 617
rect 7583 583 7617 617
rect 7651 583 7685 617
rect 7719 583 7753 617
rect 7787 583 7821 617
rect 7855 583 7889 617
rect 7923 583 7957 617
rect 7991 583 8025 617
rect 8059 583 8093 617
rect 8127 583 8161 617
rect 8195 583 8229 617
rect 8263 583 8400 617
rect 0 560 8343 583
rect 0 507 80 560
rect 0 473 23 507
rect 57 473 80 507
rect 8320 549 8343 560
rect 8377 549 8400 583
rect 8320 515 8400 549
rect 8320 481 8343 515
rect 8377 481 8400 515
rect 0 439 80 473
rect 0 405 23 439
rect 57 405 80 439
rect 0 371 80 405
rect 520 457 2120 480
rect 520 423 547 457
rect 589 423 619 457
rect 657 423 691 457
rect 725 423 759 457
rect 797 423 827 457
rect 869 423 895 457
rect 941 423 963 457
rect 1013 423 1031 457
rect 1085 423 1099 457
rect 1157 423 1167 457
rect 1229 423 1235 457
rect 1301 423 1303 457
rect 1337 423 1339 457
rect 1405 423 1411 457
rect 1473 423 1483 457
rect 1541 423 1555 457
rect 1609 423 1627 457
rect 1677 423 1699 457
rect 1745 423 1771 457
rect 1813 423 1843 457
rect 1881 423 1915 457
rect 1949 423 1983 457
rect 2021 423 2051 457
rect 2093 423 2120 457
rect 520 400 2120 423
rect 2440 457 4040 480
rect 2440 423 2467 457
rect 2509 423 2539 457
rect 2577 423 2611 457
rect 2645 423 2679 457
rect 2717 423 2747 457
rect 2789 423 2815 457
rect 2861 423 2883 457
rect 2933 423 2951 457
rect 3005 423 3019 457
rect 3077 423 3087 457
rect 3149 423 3155 457
rect 3221 423 3223 457
rect 3257 423 3259 457
rect 3325 423 3331 457
rect 3393 423 3403 457
rect 3461 423 3475 457
rect 3529 423 3547 457
rect 3597 423 3619 457
rect 3665 423 3691 457
rect 3733 423 3763 457
rect 3801 423 3835 457
rect 3869 423 3903 457
rect 3941 423 3971 457
rect 4013 423 4040 457
rect 2440 400 4040 423
rect 4360 457 5960 480
rect 4360 423 4387 457
rect 4429 423 4459 457
rect 4497 423 4531 457
rect 4565 423 4599 457
rect 4637 423 4667 457
rect 4709 423 4735 457
rect 4781 423 4803 457
rect 4853 423 4871 457
rect 4925 423 4939 457
rect 4997 423 5007 457
rect 5069 423 5075 457
rect 5141 423 5143 457
rect 5177 423 5179 457
rect 5245 423 5251 457
rect 5313 423 5323 457
rect 5381 423 5395 457
rect 5449 423 5467 457
rect 5517 423 5539 457
rect 5585 423 5611 457
rect 5653 423 5683 457
rect 5721 423 5755 457
rect 5789 423 5823 457
rect 5861 423 5891 457
rect 5933 423 5960 457
rect 4360 400 5960 423
rect 6280 457 7880 480
rect 6280 423 6307 457
rect 6349 423 6379 457
rect 6417 423 6451 457
rect 6485 423 6519 457
rect 6557 423 6587 457
rect 6629 423 6655 457
rect 6701 423 6723 457
rect 6773 423 6791 457
rect 6845 423 6859 457
rect 6917 423 6927 457
rect 6989 423 6995 457
rect 7061 423 7063 457
rect 7097 423 7099 457
rect 7165 423 7171 457
rect 7233 423 7243 457
rect 7301 423 7315 457
rect 7369 423 7387 457
rect 7437 423 7459 457
rect 7505 423 7531 457
rect 7573 423 7603 457
rect 7641 423 7675 457
rect 7709 423 7743 457
rect 7781 423 7811 457
rect 7853 423 7880 457
rect 6280 400 7880 423
rect 8320 447 8400 481
rect 8320 413 8343 447
rect 8377 413 8400 447
rect 0 337 23 371
rect 57 337 80 371
rect 8320 379 8400 413
rect 0 303 80 337
rect 0 269 23 303
rect 57 269 80 303
rect 0 235 80 269
rect 0 201 23 235
rect 57 201 80 235
rect 0 167 80 201
rect 0 133 23 167
rect 57 133 80 167
rect 0 80 80 133
rect 320 313 400 360
rect 320 277 343 313
rect 377 277 400 313
rect 320 243 400 277
rect 320 207 343 243
rect 377 207 400 243
rect 320 80 400 207
rect 2240 313 2320 360
rect 2240 277 2263 313
rect 2297 277 2320 313
rect 2240 243 2320 277
rect 2240 207 2263 243
rect 2297 207 2320 243
rect 2240 160 2320 207
rect 4160 313 4240 360
rect 4160 277 4183 313
rect 4217 277 4240 313
rect 4160 243 4240 277
rect 4160 207 4183 243
rect 4217 207 4240 243
rect 4160 160 4240 207
rect 6080 313 6160 360
rect 6080 277 6103 313
rect 6137 277 6160 313
rect 6080 243 6160 277
rect 6080 207 6103 243
rect 6137 207 6160 243
rect 6080 160 6160 207
rect 8000 313 8080 360
rect 8000 277 8023 313
rect 8057 277 8080 313
rect 8000 243 8080 277
rect 8000 207 8023 243
rect 8057 207 8080 243
rect 8000 160 8080 207
rect 8320 345 8343 379
rect 8377 345 8400 379
rect 8320 311 8400 345
rect 8320 277 8343 311
rect 8377 277 8400 311
rect 8320 243 8400 277
rect 8320 209 8343 243
rect 8377 209 8400 243
rect 8320 175 8400 209
rect 8320 141 8343 175
rect 8377 141 8400 175
rect 8320 80 8400 141
rect 0 57 8400 80
rect 0 23 137 57
rect 171 23 205 57
rect 239 23 273 57
rect 307 23 341 57
rect 375 23 409 57
rect 443 23 477 57
rect 511 23 545 57
rect 579 23 613 57
rect 647 23 681 57
rect 715 23 749 57
rect 783 23 817 57
rect 851 23 885 57
rect 919 23 953 57
rect 987 23 1021 57
rect 1055 23 1089 57
rect 1123 23 1157 57
rect 1191 23 1225 57
rect 1259 23 1293 57
rect 1327 23 1361 57
rect 1395 23 1429 57
rect 1463 23 1497 57
rect 1531 23 1565 57
rect 1599 23 1633 57
rect 1667 23 1701 57
rect 1735 23 1769 57
rect 1803 23 1837 57
rect 1871 23 1905 57
rect 1939 23 1973 57
rect 2007 23 2041 57
rect 2075 23 2109 57
rect 2143 23 2177 57
rect 2211 23 2245 57
rect 2279 23 2313 57
rect 2347 23 2381 57
rect 2415 23 2449 57
rect 2483 23 2517 57
rect 2551 23 2585 57
rect 2619 23 2653 57
rect 2687 23 2721 57
rect 2755 23 2789 57
rect 2823 23 2857 57
rect 2891 23 2925 57
rect 2959 23 2993 57
rect 3027 23 3061 57
rect 3095 23 3129 57
rect 3163 23 3197 57
rect 3231 23 3265 57
rect 3299 23 3333 57
rect 3367 23 3401 57
rect 3435 23 3469 57
rect 3503 23 3537 57
rect 3571 23 3605 57
rect 3639 23 3673 57
rect 3707 23 3741 57
rect 3775 23 3809 57
rect 3843 23 3877 57
rect 3911 23 3945 57
rect 3979 23 4013 57
rect 4047 23 4081 57
rect 4115 23 4149 57
rect 4183 23 4217 57
rect 4251 23 4285 57
rect 4319 23 4353 57
rect 4387 23 4421 57
rect 4455 23 4489 57
rect 4523 23 4557 57
rect 4591 23 4625 57
rect 4659 23 4693 57
rect 4727 23 4761 57
rect 4795 23 4829 57
rect 4863 23 4897 57
rect 4931 23 4965 57
rect 4999 23 5033 57
rect 5067 23 5101 57
rect 5135 23 5169 57
rect 5203 23 5237 57
rect 5271 23 5305 57
rect 5339 23 5373 57
rect 5407 23 5441 57
rect 5475 23 5509 57
rect 5543 23 5577 57
rect 5611 23 5645 57
rect 5679 23 5713 57
rect 5747 23 5781 57
rect 5815 23 5849 57
rect 5883 23 5917 57
rect 5951 23 5985 57
rect 6019 23 6053 57
rect 6087 23 6121 57
rect 6155 23 6189 57
rect 6223 23 6257 57
rect 6291 23 6325 57
rect 6359 23 6393 57
rect 6427 23 6461 57
rect 6495 23 6529 57
rect 6563 23 6597 57
rect 6631 23 6665 57
rect 6699 23 6733 57
rect 6767 23 6801 57
rect 6835 23 6869 57
rect 6903 23 6937 57
rect 6971 23 7005 57
rect 7039 23 7073 57
rect 7107 23 7141 57
rect 7175 23 7209 57
rect 7243 23 7277 57
rect 7311 23 7345 57
rect 7379 23 7413 57
rect 7447 23 7481 57
rect 7515 23 7549 57
rect 7583 23 7617 57
rect 7651 23 7685 57
rect 7719 23 7753 57
rect 7787 23 7821 57
rect 7855 23 7889 57
rect 7923 23 7957 57
rect 7991 23 8025 57
rect 8059 23 8093 57
rect 8127 23 8161 57
rect 8195 23 8229 57
rect 8263 23 8400 57
rect 0 0 8400 23
rect 0 -400 80 0
rect 160 -103 8240 -80
rect 160 -137 183 -103
rect 217 -137 343 -103
rect 377 -137 503 -103
rect 537 -137 663 -103
rect 697 -137 823 -103
rect 857 -137 983 -103
rect 1017 -137 1143 -103
rect 1177 -137 1463 -103
rect 1497 -137 1623 -103
rect 1657 -137 1783 -103
rect 1817 -137 1943 -103
rect 1977 -137 2103 -103
rect 2137 -137 2263 -103
rect 2297 -137 2423 -103
rect 2457 -137 2583 -103
rect 2617 -137 2743 -103
rect 2777 -137 2903 -103
rect 2937 -137 3063 -103
rect 3097 -137 3383 -103
rect 3417 -137 3543 -103
rect 3577 -137 3703 -103
rect 3737 -137 3863 -103
rect 3897 -137 4023 -103
rect 4057 -137 4183 -103
rect 4217 -137 4343 -103
rect 4377 -137 4503 -103
rect 4537 -137 4663 -103
rect 4697 -137 4823 -103
rect 4857 -137 4983 -103
rect 5017 -137 5303 -103
rect 5337 -137 5463 -103
rect 5497 -137 5623 -103
rect 5657 -137 5783 -103
rect 5817 -137 5943 -103
rect 5977 -137 6103 -103
rect 6137 -137 6263 -103
rect 6297 -137 6423 -103
rect 6457 -137 6583 -103
rect 6617 -137 6743 -103
rect 6777 -137 6903 -103
rect 6937 -137 7223 -103
rect 7257 -137 7383 -103
rect 7417 -137 7543 -103
rect 7577 -137 7703 -103
rect 7737 -137 7863 -103
rect 7897 -137 8183 -103
rect 8217 -137 8240 -103
rect 160 -320 8240 -137
rect 8320 -400 8400 0
rect 0 -423 8400 -400
rect 0 -457 137 -423
rect 171 -457 205 -423
rect 239 -457 273 -423
rect 307 -457 341 -423
rect 375 -457 409 -423
rect 443 -457 477 -423
rect 511 -457 545 -423
rect 579 -457 613 -423
rect 647 -457 681 -423
rect 715 -457 749 -423
rect 783 -457 817 -423
rect 851 -457 885 -423
rect 919 -457 953 -423
rect 987 -457 1021 -423
rect 1055 -457 1089 -423
rect 1123 -457 1157 -423
rect 1191 -457 1225 -423
rect 1259 -457 1293 -423
rect 1327 -457 1361 -423
rect 1395 -457 1429 -423
rect 1463 -457 1497 -423
rect 1531 -457 1565 -423
rect 1599 -457 1633 -423
rect 1667 -457 1701 -423
rect 1735 -457 1769 -423
rect 1803 -457 1837 -423
rect 1871 -457 1905 -423
rect 1939 -457 1973 -423
rect 2007 -457 2041 -423
rect 2075 -457 2109 -423
rect 2143 -457 2177 -423
rect 2211 -457 2245 -423
rect 2279 -457 2313 -423
rect 2347 -457 2381 -423
rect 2415 -457 2449 -423
rect 2483 -457 2517 -423
rect 2551 -457 2585 -423
rect 2619 -457 2653 -423
rect 2687 -457 2721 -423
rect 2755 -457 2789 -423
rect 2823 -457 2857 -423
rect 2891 -457 2925 -423
rect 2959 -457 2993 -423
rect 3027 -457 3061 -423
rect 3095 -457 3129 -423
rect 3163 -457 3197 -423
rect 3231 -457 3265 -423
rect 3299 -457 3333 -423
rect 3367 -457 3401 -423
rect 3435 -457 3469 -423
rect 3503 -457 3537 -423
rect 3571 -457 3605 -423
rect 3639 -457 3673 -423
rect 3707 -457 3741 -423
rect 3775 -457 3809 -423
rect 3843 -457 3877 -423
rect 3911 -457 3945 -423
rect 3979 -457 4013 -423
rect 4047 -457 4081 -423
rect 4115 -457 4149 -423
rect 4183 -457 4217 -423
rect 4251 -457 4285 -423
rect 4319 -457 4353 -423
rect 4387 -457 4421 -423
rect 4455 -457 4489 -423
rect 4523 -457 4557 -423
rect 4591 -457 4625 -423
rect 4659 -457 4693 -423
rect 4727 -457 4761 -423
rect 4795 -457 4829 -423
rect 4863 -457 4897 -423
rect 4931 -457 4965 -423
rect 4999 -457 5033 -423
rect 5067 -457 5101 -423
rect 5135 -457 5169 -423
rect 5203 -457 5237 -423
rect 5271 -457 5305 -423
rect 5339 -457 5373 -423
rect 5407 -457 5441 -423
rect 5475 -457 5509 -423
rect 5543 -457 5577 -423
rect 5611 -457 5645 -423
rect 5679 -457 5713 -423
rect 5747 -457 5781 -423
rect 5815 -457 5849 -423
rect 5883 -457 5917 -423
rect 5951 -457 5985 -423
rect 6019 -457 6053 -423
rect 6087 -457 6121 -423
rect 6155 -457 6189 -423
rect 6223 -457 6257 -423
rect 6291 -457 6325 -423
rect 6359 -457 6393 -423
rect 6427 -457 6461 -423
rect 6495 -457 6529 -423
rect 6563 -457 6597 -423
rect 6631 -457 6665 -423
rect 6699 -457 6733 -423
rect 6767 -457 6801 -423
rect 6835 -457 6869 -423
rect 6903 -457 6937 -423
rect 6971 -457 7005 -423
rect 7039 -457 7073 -423
rect 7107 -457 7141 -423
rect 7175 -457 7209 -423
rect 7243 -457 7277 -423
rect 7311 -457 7345 -423
rect 7379 -457 7413 -423
rect 7447 -457 7481 -423
rect 7515 -457 7549 -423
rect 7583 -457 7617 -423
rect 7651 -457 7685 -423
rect 7719 -457 7753 -423
rect 7787 -457 7821 -423
rect 7855 -457 7889 -423
rect 7923 -457 7957 -423
rect 7991 -457 8025 -423
rect 8059 -457 8093 -423
rect 8127 -457 8161 -423
rect 8195 -457 8229 -423
rect 8263 -457 8400 -423
rect 0 -480 8400 -457
rect 0 -533 80 -480
rect 0 -567 23 -533
rect 57 -567 80 -533
rect 8320 -533 8400 -480
rect 0 -601 80 -567
rect 0 -635 23 -601
rect 57 -635 80 -601
rect 0 -669 80 -635
rect 520 -583 2120 -560
rect 520 -617 547 -583
rect 589 -617 619 -583
rect 657 -617 691 -583
rect 725 -617 759 -583
rect 797 -617 827 -583
rect 869 -617 895 -583
rect 941 -617 963 -583
rect 1013 -617 1031 -583
rect 1085 -617 1099 -583
rect 1157 -617 1167 -583
rect 1229 -617 1235 -583
rect 1301 -617 1303 -583
rect 1337 -617 1339 -583
rect 1405 -617 1411 -583
rect 1473 -617 1483 -583
rect 1541 -617 1555 -583
rect 1609 -617 1627 -583
rect 1677 -617 1699 -583
rect 1745 -617 1771 -583
rect 1813 -617 1843 -583
rect 1881 -617 1915 -583
rect 1949 -617 1983 -583
rect 2021 -617 2051 -583
rect 2093 -617 2120 -583
rect 520 -640 2120 -617
rect 2440 -583 4040 -560
rect 2440 -617 2467 -583
rect 2509 -617 2539 -583
rect 2577 -617 2611 -583
rect 2645 -617 2679 -583
rect 2717 -617 2747 -583
rect 2789 -617 2815 -583
rect 2861 -617 2883 -583
rect 2933 -617 2951 -583
rect 3005 -617 3019 -583
rect 3077 -617 3087 -583
rect 3149 -617 3155 -583
rect 3221 -617 3223 -583
rect 3257 -617 3259 -583
rect 3325 -617 3331 -583
rect 3393 -617 3403 -583
rect 3461 -617 3475 -583
rect 3529 -617 3547 -583
rect 3597 -617 3619 -583
rect 3665 -617 3691 -583
rect 3733 -617 3763 -583
rect 3801 -617 3835 -583
rect 3869 -617 3903 -583
rect 3941 -617 3971 -583
rect 4013 -617 4040 -583
rect 2440 -640 4040 -617
rect 4360 -583 5960 -560
rect 4360 -617 4387 -583
rect 4429 -617 4459 -583
rect 4497 -617 4531 -583
rect 4565 -617 4599 -583
rect 4637 -617 4667 -583
rect 4709 -617 4735 -583
rect 4781 -617 4803 -583
rect 4853 -617 4871 -583
rect 4925 -617 4939 -583
rect 4997 -617 5007 -583
rect 5069 -617 5075 -583
rect 5141 -617 5143 -583
rect 5177 -617 5179 -583
rect 5245 -617 5251 -583
rect 5313 -617 5323 -583
rect 5381 -617 5395 -583
rect 5449 -617 5467 -583
rect 5517 -617 5539 -583
rect 5585 -617 5611 -583
rect 5653 -617 5683 -583
rect 5721 -617 5755 -583
rect 5789 -617 5823 -583
rect 5861 -617 5891 -583
rect 5933 -617 5960 -583
rect 4360 -640 5960 -617
rect 6280 -583 7880 -560
rect 6280 -617 6307 -583
rect 6349 -617 6379 -583
rect 6417 -617 6451 -583
rect 6485 -617 6519 -583
rect 6557 -617 6587 -583
rect 6629 -617 6655 -583
rect 6701 -617 6723 -583
rect 6773 -617 6791 -583
rect 6845 -617 6859 -583
rect 6917 -617 6927 -583
rect 6989 -617 6995 -583
rect 7061 -617 7063 -583
rect 7097 -617 7099 -583
rect 7165 -617 7171 -583
rect 7233 -617 7243 -583
rect 7301 -617 7315 -583
rect 7369 -617 7387 -583
rect 7437 -617 7459 -583
rect 7505 -617 7531 -583
rect 7573 -617 7603 -583
rect 7641 -617 7675 -583
rect 7709 -617 7743 -583
rect 7781 -617 7811 -583
rect 7853 -617 7880 -583
rect 6280 -640 7880 -617
rect 8320 -567 8343 -533
rect 8377 -567 8400 -533
rect 8320 -601 8400 -567
rect 8320 -635 8343 -601
rect 8377 -635 8400 -601
rect 0 -703 23 -669
rect 57 -703 80 -669
rect 8320 -669 8400 -635
rect 0 -737 80 -703
rect 0 -771 23 -737
rect 57 -771 80 -737
rect 0 -805 80 -771
rect 0 -839 23 -805
rect 57 -839 80 -805
rect 0 -873 80 -839
rect 0 -907 23 -873
rect 57 -907 80 -873
rect 0 -960 80 -907
rect 320 -727 400 -680
rect 320 -763 343 -727
rect 377 -763 400 -727
rect 320 -797 400 -763
rect 320 -833 343 -797
rect 377 -833 400 -797
rect 320 -960 400 -833
rect 2240 -727 2320 -680
rect 2240 -763 2263 -727
rect 2297 -763 2320 -727
rect 2240 -797 2320 -763
rect 2240 -833 2263 -797
rect 2297 -833 2320 -797
rect 2240 -880 2320 -833
rect 4160 -727 4240 -680
rect 4160 -763 4183 -727
rect 4217 -763 4240 -727
rect 4160 -797 4240 -763
rect 4160 -833 4183 -797
rect 4217 -833 4240 -797
rect 4160 -880 4240 -833
rect 6080 -727 6160 -680
rect 6080 -763 6103 -727
rect 6137 -763 6160 -727
rect 6080 -797 6160 -763
rect 6080 -833 6103 -797
rect 6137 -833 6160 -797
rect 6080 -880 6160 -833
rect 8000 -727 8080 -680
rect 8000 -763 8023 -727
rect 8057 -763 8080 -727
rect 8000 -797 8080 -763
rect 8000 -833 8023 -797
rect 8057 -833 8080 -797
rect 8000 -880 8080 -833
rect 8320 -703 8343 -669
rect 8377 -703 8400 -669
rect 8320 -737 8400 -703
rect 8320 -771 8343 -737
rect 8377 -771 8400 -737
rect 8320 -805 8400 -771
rect 8320 -839 8343 -805
rect 8377 -839 8400 -805
rect 8320 -873 8400 -839
rect 8320 -907 8343 -873
rect 8377 -907 8400 -873
rect 8320 -960 8400 -907
rect 0 -983 8400 -960
rect 0 -1017 137 -983
rect 171 -1017 205 -983
rect 239 -1017 273 -983
rect 307 -1017 341 -983
rect 375 -1017 409 -983
rect 443 -1017 477 -983
rect 511 -1017 545 -983
rect 579 -1017 613 -983
rect 647 -1017 681 -983
rect 715 -1017 749 -983
rect 783 -1017 817 -983
rect 851 -1017 885 -983
rect 919 -1017 953 -983
rect 987 -1017 1021 -983
rect 1055 -1017 1089 -983
rect 1123 -1017 1157 -983
rect 1191 -1017 1225 -983
rect 1259 -1017 1293 -983
rect 1327 -1017 1361 -983
rect 1395 -1017 1429 -983
rect 1463 -1017 1497 -983
rect 1531 -1017 1565 -983
rect 1599 -1017 1633 -983
rect 1667 -1017 1701 -983
rect 1735 -1017 1769 -983
rect 1803 -1017 1837 -983
rect 1871 -1017 1905 -983
rect 1939 -1017 1973 -983
rect 2007 -1017 2041 -983
rect 2075 -1017 2109 -983
rect 2143 -1017 2177 -983
rect 2211 -1017 2245 -983
rect 2279 -1017 2313 -983
rect 2347 -1017 2381 -983
rect 2415 -1017 2449 -983
rect 2483 -1017 2517 -983
rect 2551 -1017 2585 -983
rect 2619 -1017 2653 -983
rect 2687 -1017 2721 -983
rect 2755 -1017 2789 -983
rect 2823 -1017 2857 -983
rect 2891 -1017 2925 -983
rect 2959 -1017 2993 -983
rect 3027 -1017 3061 -983
rect 3095 -1017 3129 -983
rect 3163 -1017 3197 -983
rect 3231 -1017 3265 -983
rect 3299 -1017 3333 -983
rect 3367 -1017 3401 -983
rect 3435 -1017 3469 -983
rect 3503 -1017 3537 -983
rect 3571 -1017 3605 -983
rect 3639 -1017 3673 -983
rect 3707 -1017 3741 -983
rect 3775 -1017 3809 -983
rect 3843 -1017 3877 -983
rect 3911 -1017 3945 -983
rect 3979 -1017 4013 -983
rect 4047 -1017 4081 -983
rect 4115 -1017 4149 -983
rect 4183 -1017 4217 -983
rect 4251 -1017 4285 -983
rect 4319 -1017 4353 -983
rect 4387 -1017 4421 -983
rect 4455 -1017 4489 -983
rect 4523 -1017 4557 -983
rect 4591 -1017 4625 -983
rect 4659 -1017 4693 -983
rect 4727 -1017 4761 -983
rect 4795 -1017 4829 -983
rect 4863 -1017 4897 -983
rect 4931 -1017 4965 -983
rect 4999 -1017 5033 -983
rect 5067 -1017 5101 -983
rect 5135 -1017 5169 -983
rect 5203 -1017 5237 -983
rect 5271 -1017 5305 -983
rect 5339 -1017 5373 -983
rect 5407 -1017 5441 -983
rect 5475 -1017 5509 -983
rect 5543 -1017 5577 -983
rect 5611 -1017 5645 -983
rect 5679 -1017 5713 -983
rect 5747 -1017 5781 -983
rect 5815 -1017 5849 -983
rect 5883 -1017 5917 -983
rect 5951 -1017 5985 -983
rect 6019 -1017 6053 -983
rect 6087 -1017 6121 -983
rect 6155 -1017 6189 -983
rect 6223 -1017 6257 -983
rect 6291 -1017 6325 -983
rect 6359 -1017 6393 -983
rect 6427 -1017 6461 -983
rect 6495 -1017 6529 -983
rect 6563 -1017 6597 -983
rect 6631 -1017 6665 -983
rect 6699 -1017 6733 -983
rect 6767 -1017 6801 -983
rect 6835 -1017 6869 -983
rect 6903 -1017 6937 -983
rect 6971 -1017 7005 -983
rect 7039 -1017 7073 -983
rect 7107 -1017 7141 -983
rect 7175 -1017 7209 -983
rect 7243 -1017 7277 -983
rect 7311 -1017 7345 -983
rect 7379 -1017 7413 -983
rect 7447 -1017 7481 -983
rect 7515 -1017 7549 -983
rect 7583 -1017 7617 -983
rect 7651 -1017 7685 -983
rect 7719 -1017 7753 -983
rect 7787 -1017 7821 -983
rect 7855 -1017 7889 -983
rect 7923 -1017 7957 -983
rect 7991 -1017 8025 -983
rect 8059 -1017 8093 -983
rect 8127 -1017 8161 -983
rect 8195 -1017 8229 -983
rect 8263 -1017 8400 -983
rect 0 -1040 8400 -1017
<< viali >>
rect 343 9715 377 9729
rect 343 9695 377 9715
rect 343 9647 377 9657
rect 343 9623 377 9647
rect 343 9579 377 9585
rect 343 9551 377 9579
rect 343 9511 377 9513
rect 343 9479 377 9511
rect 343 9409 377 9441
rect 343 9407 377 9409
rect 343 9341 377 9369
rect 343 9335 377 9341
rect 343 9273 377 9297
rect 343 9263 377 9273
rect 343 9205 377 9225
rect 343 9191 377 9205
rect 2263 9715 2297 9729
rect 2263 9695 2297 9715
rect 2263 9647 2297 9657
rect 2263 9623 2297 9647
rect 2263 9579 2297 9585
rect 2263 9551 2297 9579
rect 2263 9511 2297 9513
rect 2263 9479 2297 9511
rect 2263 9409 2297 9441
rect 2263 9407 2297 9409
rect 2263 9341 2297 9369
rect 2263 9335 2297 9341
rect 2263 9273 2297 9297
rect 2263 9263 2297 9273
rect 2263 9205 2297 9225
rect 2263 9191 2297 9205
rect 4183 9715 4217 9729
rect 4183 9695 4217 9715
rect 4183 9647 4217 9657
rect 4183 9623 4217 9647
rect 4183 9579 4217 9585
rect 4183 9551 4217 9579
rect 4183 9511 4217 9513
rect 4183 9479 4217 9511
rect 4183 9409 4217 9441
rect 4183 9407 4217 9409
rect 4183 9341 4217 9369
rect 4183 9335 4217 9341
rect 4183 9273 4217 9297
rect 4183 9263 4217 9273
rect 4183 9205 4217 9225
rect 4183 9191 4217 9205
rect 6103 9715 6137 9729
rect 6103 9695 6137 9715
rect 6103 9647 6137 9657
rect 6103 9623 6137 9647
rect 6103 9579 6137 9585
rect 6103 9551 6137 9579
rect 6103 9511 6137 9513
rect 6103 9479 6137 9511
rect 6103 9409 6137 9441
rect 6103 9407 6137 9409
rect 6103 9341 6137 9369
rect 6103 9335 6137 9341
rect 6103 9273 6137 9297
rect 6103 9263 6137 9273
rect 6103 9205 6137 9225
rect 6103 9191 6137 9205
rect 8023 9715 8057 9729
rect 8023 9695 8057 9715
rect 8023 9647 8057 9657
rect 8023 9623 8057 9647
rect 8023 9579 8057 9585
rect 8023 9551 8057 9579
rect 8023 9511 8057 9513
rect 8023 9479 8057 9511
rect 8023 9409 8057 9441
rect 8023 9407 8057 9409
rect 8023 9341 8057 9369
rect 8023 9335 8057 9341
rect 8023 9273 8057 9297
rect 8023 9263 8057 9273
rect 8023 9205 8057 9225
rect 8023 9191 8057 9205
rect 547 9063 555 9097
rect 555 9063 581 9097
rect 619 9063 623 9097
rect 623 9063 653 9097
rect 691 9063 725 9097
rect 763 9063 793 9097
rect 793 9063 797 9097
rect 835 9063 861 9097
rect 861 9063 869 9097
rect 907 9063 929 9097
rect 929 9063 941 9097
rect 979 9063 997 9097
rect 997 9063 1013 9097
rect 1051 9063 1065 9097
rect 1065 9063 1085 9097
rect 1123 9063 1133 9097
rect 1133 9063 1157 9097
rect 1195 9063 1201 9097
rect 1201 9063 1229 9097
rect 1267 9063 1269 9097
rect 1269 9063 1301 9097
rect 1339 9063 1371 9097
rect 1371 9063 1373 9097
rect 1411 9063 1439 9097
rect 1439 9063 1445 9097
rect 1483 9063 1507 9097
rect 1507 9063 1517 9097
rect 1555 9063 1575 9097
rect 1575 9063 1589 9097
rect 1627 9063 1643 9097
rect 1643 9063 1661 9097
rect 1699 9063 1711 9097
rect 1711 9063 1733 9097
rect 1771 9063 1779 9097
rect 1779 9063 1805 9097
rect 1843 9063 1847 9097
rect 1847 9063 1877 9097
rect 1915 9063 1949 9097
rect 1987 9063 2017 9097
rect 2017 9063 2021 9097
rect 2059 9063 2085 9097
rect 2085 9063 2093 9097
rect 2467 9063 2475 9097
rect 2475 9063 2501 9097
rect 2539 9063 2543 9097
rect 2543 9063 2573 9097
rect 2611 9063 2645 9097
rect 2683 9063 2713 9097
rect 2713 9063 2717 9097
rect 2755 9063 2781 9097
rect 2781 9063 2789 9097
rect 2827 9063 2849 9097
rect 2849 9063 2861 9097
rect 2899 9063 2917 9097
rect 2917 9063 2933 9097
rect 2971 9063 2985 9097
rect 2985 9063 3005 9097
rect 3043 9063 3053 9097
rect 3053 9063 3077 9097
rect 3115 9063 3121 9097
rect 3121 9063 3149 9097
rect 3187 9063 3189 9097
rect 3189 9063 3221 9097
rect 3259 9063 3291 9097
rect 3291 9063 3293 9097
rect 3331 9063 3359 9097
rect 3359 9063 3365 9097
rect 3403 9063 3427 9097
rect 3427 9063 3437 9097
rect 3475 9063 3495 9097
rect 3495 9063 3509 9097
rect 3547 9063 3563 9097
rect 3563 9063 3581 9097
rect 3619 9063 3631 9097
rect 3631 9063 3653 9097
rect 3691 9063 3699 9097
rect 3699 9063 3725 9097
rect 3763 9063 3767 9097
rect 3767 9063 3797 9097
rect 3835 9063 3869 9097
rect 3907 9063 3937 9097
rect 3937 9063 3941 9097
rect 3979 9063 4005 9097
rect 4005 9063 4013 9097
rect 4387 9063 4395 9097
rect 4395 9063 4421 9097
rect 4459 9063 4463 9097
rect 4463 9063 4493 9097
rect 4531 9063 4565 9097
rect 4603 9063 4633 9097
rect 4633 9063 4637 9097
rect 4675 9063 4701 9097
rect 4701 9063 4709 9097
rect 4747 9063 4769 9097
rect 4769 9063 4781 9097
rect 4819 9063 4837 9097
rect 4837 9063 4853 9097
rect 4891 9063 4905 9097
rect 4905 9063 4925 9097
rect 4963 9063 4973 9097
rect 4973 9063 4997 9097
rect 5035 9063 5041 9097
rect 5041 9063 5069 9097
rect 5107 9063 5109 9097
rect 5109 9063 5141 9097
rect 5179 9063 5211 9097
rect 5211 9063 5213 9097
rect 5251 9063 5279 9097
rect 5279 9063 5285 9097
rect 5323 9063 5347 9097
rect 5347 9063 5357 9097
rect 5395 9063 5415 9097
rect 5415 9063 5429 9097
rect 5467 9063 5483 9097
rect 5483 9063 5501 9097
rect 5539 9063 5551 9097
rect 5551 9063 5573 9097
rect 5611 9063 5619 9097
rect 5619 9063 5645 9097
rect 5683 9063 5687 9097
rect 5687 9063 5717 9097
rect 5755 9063 5789 9097
rect 5827 9063 5857 9097
rect 5857 9063 5861 9097
rect 5899 9063 5925 9097
rect 5925 9063 5933 9097
rect 6307 9063 6315 9097
rect 6315 9063 6341 9097
rect 6379 9063 6383 9097
rect 6383 9063 6413 9097
rect 6451 9063 6485 9097
rect 6523 9063 6553 9097
rect 6553 9063 6557 9097
rect 6595 9063 6621 9097
rect 6621 9063 6629 9097
rect 6667 9063 6689 9097
rect 6689 9063 6701 9097
rect 6739 9063 6757 9097
rect 6757 9063 6773 9097
rect 6811 9063 6825 9097
rect 6825 9063 6845 9097
rect 6883 9063 6893 9097
rect 6893 9063 6917 9097
rect 6955 9063 6961 9097
rect 6961 9063 6989 9097
rect 7027 9063 7029 9097
rect 7029 9063 7061 9097
rect 7099 9063 7131 9097
rect 7131 9063 7133 9097
rect 7171 9063 7199 9097
rect 7199 9063 7205 9097
rect 7243 9063 7267 9097
rect 7267 9063 7277 9097
rect 7315 9063 7335 9097
rect 7335 9063 7349 9097
rect 7387 9063 7403 9097
rect 7403 9063 7421 9097
rect 7459 9063 7471 9097
rect 7471 9063 7493 9097
rect 7531 9063 7539 9097
rect 7539 9063 7565 9097
rect 7603 9063 7607 9097
rect 7607 9063 7637 9097
rect 7675 9063 7709 9097
rect 7747 9063 7777 9097
rect 7777 9063 7781 9097
rect 7819 9063 7845 9097
rect 7845 9063 7853 9097
rect 183 8423 217 8457
rect 8183 8423 8217 8457
rect 183 8263 217 8297
rect 8183 8263 8217 8297
rect 547 7783 555 7817
rect 555 7783 581 7817
rect 619 7783 623 7817
rect 623 7783 653 7817
rect 691 7783 725 7817
rect 763 7783 793 7817
rect 793 7783 797 7817
rect 835 7783 861 7817
rect 861 7783 869 7817
rect 907 7783 929 7817
rect 929 7783 941 7817
rect 979 7783 997 7817
rect 997 7783 1013 7817
rect 1051 7783 1065 7817
rect 1065 7783 1085 7817
rect 1123 7783 1133 7817
rect 1133 7783 1157 7817
rect 1195 7783 1201 7817
rect 1201 7783 1229 7817
rect 1267 7783 1269 7817
rect 1269 7783 1301 7817
rect 1339 7783 1371 7817
rect 1371 7783 1373 7817
rect 1411 7783 1439 7817
rect 1439 7783 1445 7817
rect 1483 7783 1507 7817
rect 1507 7783 1517 7817
rect 1555 7783 1575 7817
rect 1575 7783 1589 7817
rect 1627 7783 1643 7817
rect 1643 7783 1661 7817
rect 1699 7783 1711 7817
rect 1711 7783 1733 7817
rect 1771 7783 1779 7817
rect 1779 7783 1805 7817
rect 1843 7783 1847 7817
rect 1847 7783 1877 7817
rect 1915 7783 1949 7817
rect 1987 7783 2017 7817
rect 2017 7783 2021 7817
rect 2059 7783 2085 7817
rect 2085 7783 2093 7817
rect 2467 7783 2475 7817
rect 2475 7783 2501 7817
rect 2539 7783 2543 7817
rect 2543 7783 2573 7817
rect 2611 7783 2645 7817
rect 2683 7783 2713 7817
rect 2713 7783 2717 7817
rect 2755 7783 2781 7817
rect 2781 7783 2789 7817
rect 2827 7783 2849 7817
rect 2849 7783 2861 7817
rect 2899 7783 2917 7817
rect 2917 7783 2933 7817
rect 2971 7783 2985 7817
rect 2985 7783 3005 7817
rect 3043 7783 3053 7817
rect 3053 7783 3077 7817
rect 3115 7783 3121 7817
rect 3121 7783 3149 7817
rect 3187 7783 3189 7817
rect 3189 7783 3221 7817
rect 3259 7783 3291 7817
rect 3291 7783 3293 7817
rect 3331 7783 3359 7817
rect 3359 7783 3365 7817
rect 3403 7783 3427 7817
rect 3427 7783 3437 7817
rect 3475 7783 3495 7817
rect 3495 7783 3509 7817
rect 3547 7783 3563 7817
rect 3563 7783 3581 7817
rect 3619 7783 3631 7817
rect 3631 7783 3653 7817
rect 3691 7783 3699 7817
rect 3699 7783 3725 7817
rect 3763 7783 3767 7817
rect 3767 7783 3797 7817
rect 3835 7783 3869 7817
rect 3907 7783 3937 7817
rect 3937 7783 3941 7817
rect 3979 7783 4005 7817
rect 4005 7783 4013 7817
rect 4387 7783 4395 7817
rect 4395 7783 4421 7817
rect 4459 7783 4463 7817
rect 4463 7783 4493 7817
rect 4531 7783 4565 7817
rect 4603 7783 4633 7817
rect 4633 7783 4637 7817
rect 4675 7783 4701 7817
rect 4701 7783 4709 7817
rect 4747 7783 4769 7817
rect 4769 7783 4781 7817
rect 4819 7783 4837 7817
rect 4837 7783 4853 7817
rect 4891 7783 4905 7817
rect 4905 7783 4925 7817
rect 4963 7783 4973 7817
rect 4973 7783 4997 7817
rect 5035 7783 5041 7817
rect 5041 7783 5069 7817
rect 5107 7783 5109 7817
rect 5109 7783 5141 7817
rect 5179 7783 5211 7817
rect 5211 7783 5213 7817
rect 5251 7783 5279 7817
rect 5279 7783 5285 7817
rect 5323 7783 5347 7817
rect 5347 7783 5357 7817
rect 5395 7783 5415 7817
rect 5415 7783 5429 7817
rect 5467 7783 5483 7817
rect 5483 7783 5501 7817
rect 5539 7783 5551 7817
rect 5551 7783 5573 7817
rect 5611 7783 5619 7817
rect 5619 7783 5645 7817
rect 5683 7783 5687 7817
rect 5687 7783 5717 7817
rect 5755 7783 5789 7817
rect 5827 7783 5857 7817
rect 5857 7783 5861 7817
rect 5899 7783 5925 7817
rect 5925 7783 5933 7817
rect 6307 7783 6315 7817
rect 6315 7783 6341 7817
rect 6379 7783 6383 7817
rect 6383 7783 6413 7817
rect 6451 7783 6485 7817
rect 6523 7783 6553 7817
rect 6553 7783 6557 7817
rect 6595 7783 6621 7817
rect 6621 7783 6629 7817
rect 6667 7783 6689 7817
rect 6689 7783 6701 7817
rect 6739 7783 6757 7817
rect 6757 7783 6773 7817
rect 6811 7783 6825 7817
rect 6825 7783 6845 7817
rect 6883 7783 6893 7817
rect 6893 7783 6917 7817
rect 6955 7783 6961 7817
rect 6961 7783 6989 7817
rect 7027 7783 7029 7817
rect 7029 7783 7061 7817
rect 7099 7783 7131 7817
rect 7131 7783 7133 7817
rect 7171 7783 7199 7817
rect 7199 7783 7205 7817
rect 7243 7783 7267 7817
rect 7267 7783 7277 7817
rect 7315 7783 7335 7817
rect 7335 7783 7349 7817
rect 7387 7783 7403 7817
rect 7403 7783 7421 7817
rect 7459 7783 7471 7817
rect 7471 7783 7493 7817
rect 7531 7783 7539 7817
rect 7539 7783 7565 7817
rect 7603 7783 7607 7817
rect 7607 7783 7637 7817
rect 7675 7783 7709 7817
rect 7747 7783 7777 7817
rect 7777 7783 7781 7817
rect 7819 7783 7845 7817
rect 7845 7783 7853 7817
rect 343 7671 377 7673
rect 343 7639 377 7671
rect 343 7569 377 7601
rect 343 7567 377 7569
rect 2263 7671 2297 7673
rect 2263 7639 2297 7671
rect 2263 7569 2297 7601
rect 2263 7567 2297 7569
rect 4183 7671 4217 7673
rect 4183 7639 4217 7671
rect 4183 7569 4217 7601
rect 4183 7567 4217 7569
rect 6103 7671 6137 7673
rect 6103 7639 6137 7671
rect 6103 7569 6137 7601
rect 6103 7567 6137 7569
rect 8023 7671 8057 7673
rect 8023 7639 8057 7671
rect 8023 7569 8057 7601
rect 8023 7567 8057 7569
rect 343 7071 377 7073
rect 343 7039 377 7071
rect 343 6969 377 7001
rect 343 6967 377 6969
rect 2263 7071 2297 7073
rect 2263 7039 2297 7071
rect 2263 6969 2297 7001
rect 2263 6967 2297 6969
rect 4183 7071 4217 7073
rect 4183 7039 4217 7071
rect 4183 6969 4217 7001
rect 4183 6967 4217 6969
rect 6103 7071 6137 7073
rect 6103 7039 6137 7071
rect 6103 6969 6137 7001
rect 6103 6967 6137 6969
rect 8023 7071 8057 7073
rect 8023 7039 8057 7071
rect 8023 6969 8057 7001
rect 8023 6967 8057 6969
rect 547 6823 555 6857
rect 555 6823 581 6857
rect 619 6823 623 6857
rect 623 6823 653 6857
rect 691 6823 725 6857
rect 763 6823 793 6857
rect 793 6823 797 6857
rect 835 6823 861 6857
rect 861 6823 869 6857
rect 907 6823 929 6857
rect 929 6823 941 6857
rect 979 6823 997 6857
rect 997 6823 1013 6857
rect 1051 6823 1065 6857
rect 1065 6823 1085 6857
rect 1123 6823 1133 6857
rect 1133 6823 1157 6857
rect 1195 6823 1201 6857
rect 1201 6823 1229 6857
rect 1267 6823 1269 6857
rect 1269 6823 1301 6857
rect 1339 6823 1371 6857
rect 1371 6823 1373 6857
rect 1411 6823 1439 6857
rect 1439 6823 1445 6857
rect 1483 6823 1507 6857
rect 1507 6823 1517 6857
rect 1555 6823 1575 6857
rect 1575 6823 1589 6857
rect 1627 6823 1643 6857
rect 1643 6823 1661 6857
rect 1699 6823 1711 6857
rect 1711 6823 1733 6857
rect 1771 6823 1779 6857
rect 1779 6823 1805 6857
rect 1843 6823 1847 6857
rect 1847 6823 1877 6857
rect 1915 6823 1949 6857
rect 1987 6823 2017 6857
rect 2017 6823 2021 6857
rect 2059 6823 2085 6857
rect 2085 6823 2093 6857
rect 2467 6823 2475 6857
rect 2475 6823 2501 6857
rect 2539 6823 2543 6857
rect 2543 6823 2573 6857
rect 2611 6823 2645 6857
rect 2683 6823 2713 6857
rect 2713 6823 2717 6857
rect 2755 6823 2781 6857
rect 2781 6823 2789 6857
rect 2827 6823 2849 6857
rect 2849 6823 2861 6857
rect 2899 6823 2917 6857
rect 2917 6823 2933 6857
rect 2971 6823 2985 6857
rect 2985 6823 3005 6857
rect 3043 6823 3053 6857
rect 3053 6823 3077 6857
rect 3115 6823 3121 6857
rect 3121 6823 3149 6857
rect 3187 6823 3189 6857
rect 3189 6823 3221 6857
rect 3259 6823 3291 6857
rect 3291 6823 3293 6857
rect 3331 6823 3359 6857
rect 3359 6823 3365 6857
rect 3403 6823 3427 6857
rect 3427 6823 3437 6857
rect 3475 6823 3495 6857
rect 3495 6823 3509 6857
rect 3547 6823 3563 6857
rect 3563 6823 3581 6857
rect 3619 6823 3631 6857
rect 3631 6823 3653 6857
rect 3691 6823 3699 6857
rect 3699 6823 3725 6857
rect 3763 6823 3767 6857
rect 3767 6823 3797 6857
rect 3835 6823 3869 6857
rect 3907 6823 3937 6857
rect 3937 6823 3941 6857
rect 3979 6823 4005 6857
rect 4005 6823 4013 6857
rect 4387 6823 4395 6857
rect 4395 6823 4421 6857
rect 4459 6823 4463 6857
rect 4463 6823 4493 6857
rect 4531 6823 4565 6857
rect 4603 6823 4633 6857
rect 4633 6823 4637 6857
rect 4675 6823 4701 6857
rect 4701 6823 4709 6857
rect 4747 6823 4769 6857
rect 4769 6823 4781 6857
rect 4819 6823 4837 6857
rect 4837 6823 4853 6857
rect 4891 6823 4905 6857
rect 4905 6823 4925 6857
rect 4963 6823 4973 6857
rect 4973 6823 4997 6857
rect 5035 6823 5041 6857
rect 5041 6823 5069 6857
rect 5107 6823 5109 6857
rect 5109 6823 5141 6857
rect 5179 6823 5211 6857
rect 5211 6823 5213 6857
rect 5251 6823 5279 6857
rect 5279 6823 5285 6857
rect 5323 6823 5347 6857
rect 5347 6823 5357 6857
rect 5395 6823 5415 6857
rect 5415 6823 5429 6857
rect 5467 6823 5483 6857
rect 5483 6823 5501 6857
rect 5539 6823 5551 6857
rect 5551 6823 5573 6857
rect 5611 6823 5619 6857
rect 5619 6823 5645 6857
rect 5683 6823 5687 6857
rect 5687 6823 5717 6857
rect 5755 6823 5789 6857
rect 5827 6823 5857 6857
rect 5857 6823 5861 6857
rect 5899 6823 5925 6857
rect 5925 6823 5933 6857
rect 6307 6823 6315 6857
rect 6315 6823 6341 6857
rect 6379 6823 6383 6857
rect 6383 6823 6413 6857
rect 6451 6823 6485 6857
rect 6523 6823 6553 6857
rect 6553 6823 6557 6857
rect 6595 6823 6621 6857
rect 6621 6823 6629 6857
rect 6667 6823 6689 6857
rect 6689 6823 6701 6857
rect 6739 6823 6757 6857
rect 6757 6823 6773 6857
rect 6811 6823 6825 6857
rect 6825 6823 6845 6857
rect 6883 6823 6893 6857
rect 6893 6823 6917 6857
rect 6955 6823 6961 6857
rect 6961 6823 6989 6857
rect 7027 6823 7029 6857
rect 7029 6823 7061 6857
rect 7099 6823 7131 6857
rect 7131 6823 7133 6857
rect 7171 6823 7199 6857
rect 7199 6823 7205 6857
rect 7243 6823 7267 6857
rect 7267 6823 7277 6857
rect 7315 6823 7335 6857
rect 7335 6823 7349 6857
rect 7387 6823 7403 6857
rect 7403 6823 7421 6857
rect 7459 6823 7471 6857
rect 7471 6823 7493 6857
rect 7531 6823 7539 6857
rect 7539 6823 7565 6857
rect 7603 6823 7607 6857
rect 7607 6823 7637 6857
rect 7675 6823 7709 6857
rect 7747 6823 7777 6857
rect 7777 6823 7781 6857
rect 7819 6823 7845 6857
rect 7845 6823 7853 6857
rect 183 6343 217 6377
rect 8183 6343 8217 6377
rect 183 6183 217 6217
rect 8183 6183 8217 6217
rect 183 5863 217 5897
rect 8183 5863 8217 5897
rect 183 5703 217 5737
rect 8183 5703 8217 5737
rect 547 5063 555 5097
rect 555 5063 581 5097
rect 619 5063 623 5097
rect 623 5063 653 5097
rect 691 5063 725 5097
rect 763 5063 793 5097
rect 793 5063 797 5097
rect 835 5063 861 5097
rect 861 5063 869 5097
rect 907 5063 929 5097
rect 929 5063 941 5097
rect 979 5063 997 5097
rect 997 5063 1013 5097
rect 1051 5063 1065 5097
rect 1065 5063 1085 5097
rect 1123 5063 1133 5097
rect 1133 5063 1157 5097
rect 1195 5063 1201 5097
rect 1201 5063 1229 5097
rect 1267 5063 1269 5097
rect 1269 5063 1301 5097
rect 1339 5063 1371 5097
rect 1371 5063 1373 5097
rect 1411 5063 1439 5097
rect 1439 5063 1445 5097
rect 1483 5063 1507 5097
rect 1507 5063 1517 5097
rect 1555 5063 1575 5097
rect 1575 5063 1589 5097
rect 1627 5063 1643 5097
rect 1643 5063 1661 5097
rect 1699 5063 1711 5097
rect 1711 5063 1733 5097
rect 1771 5063 1779 5097
rect 1779 5063 1805 5097
rect 1843 5063 1847 5097
rect 1847 5063 1877 5097
rect 1915 5063 1949 5097
rect 1987 5063 2017 5097
rect 2017 5063 2021 5097
rect 2059 5063 2085 5097
rect 2085 5063 2093 5097
rect 2467 5063 2475 5097
rect 2475 5063 2501 5097
rect 2539 5063 2543 5097
rect 2543 5063 2573 5097
rect 2611 5063 2645 5097
rect 2683 5063 2713 5097
rect 2713 5063 2717 5097
rect 2755 5063 2781 5097
rect 2781 5063 2789 5097
rect 2827 5063 2849 5097
rect 2849 5063 2861 5097
rect 2899 5063 2917 5097
rect 2917 5063 2933 5097
rect 2971 5063 2985 5097
rect 2985 5063 3005 5097
rect 3043 5063 3053 5097
rect 3053 5063 3077 5097
rect 3115 5063 3121 5097
rect 3121 5063 3149 5097
rect 3187 5063 3189 5097
rect 3189 5063 3221 5097
rect 3259 5063 3291 5097
rect 3291 5063 3293 5097
rect 3331 5063 3359 5097
rect 3359 5063 3365 5097
rect 3403 5063 3427 5097
rect 3427 5063 3437 5097
rect 3475 5063 3495 5097
rect 3495 5063 3509 5097
rect 3547 5063 3563 5097
rect 3563 5063 3581 5097
rect 3619 5063 3631 5097
rect 3631 5063 3653 5097
rect 3691 5063 3699 5097
rect 3699 5063 3725 5097
rect 3763 5063 3767 5097
rect 3767 5063 3797 5097
rect 3835 5063 3869 5097
rect 3907 5063 3937 5097
rect 3937 5063 3941 5097
rect 3979 5063 4005 5097
rect 4005 5063 4013 5097
rect 4387 5063 4395 5097
rect 4395 5063 4421 5097
rect 4459 5063 4463 5097
rect 4463 5063 4493 5097
rect 4531 5063 4565 5097
rect 4603 5063 4633 5097
rect 4633 5063 4637 5097
rect 4675 5063 4701 5097
rect 4701 5063 4709 5097
rect 4747 5063 4769 5097
rect 4769 5063 4781 5097
rect 4819 5063 4837 5097
rect 4837 5063 4853 5097
rect 4891 5063 4905 5097
rect 4905 5063 4925 5097
rect 4963 5063 4973 5097
rect 4973 5063 4997 5097
rect 5035 5063 5041 5097
rect 5041 5063 5069 5097
rect 5107 5063 5109 5097
rect 5109 5063 5141 5097
rect 5179 5063 5211 5097
rect 5211 5063 5213 5097
rect 5251 5063 5279 5097
rect 5279 5063 5285 5097
rect 5323 5063 5347 5097
rect 5347 5063 5357 5097
rect 5395 5063 5415 5097
rect 5415 5063 5429 5097
rect 5467 5063 5483 5097
rect 5483 5063 5501 5097
rect 5539 5063 5551 5097
rect 5551 5063 5573 5097
rect 5611 5063 5619 5097
rect 5619 5063 5645 5097
rect 5683 5063 5687 5097
rect 5687 5063 5717 5097
rect 5755 5063 5789 5097
rect 5827 5063 5857 5097
rect 5857 5063 5861 5097
rect 5899 5063 5925 5097
rect 5925 5063 5933 5097
rect 6307 5063 6315 5097
rect 6315 5063 6341 5097
rect 6379 5063 6383 5097
rect 6383 5063 6413 5097
rect 6451 5063 6485 5097
rect 6523 5063 6553 5097
rect 6553 5063 6557 5097
rect 6595 5063 6621 5097
rect 6621 5063 6629 5097
rect 6667 5063 6689 5097
rect 6689 5063 6701 5097
rect 6739 5063 6757 5097
rect 6757 5063 6773 5097
rect 6811 5063 6825 5097
rect 6825 5063 6845 5097
rect 6883 5063 6893 5097
rect 6893 5063 6917 5097
rect 6955 5063 6961 5097
rect 6961 5063 6989 5097
rect 7027 5063 7029 5097
rect 7029 5063 7061 5097
rect 7099 5063 7131 5097
rect 7131 5063 7133 5097
rect 7171 5063 7199 5097
rect 7199 5063 7205 5097
rect 7243 5063 7267 5097
rect 7267 5063 7277 5097
rect 7315 5063 7335 5097
rect 7335 5063 7349 5097
rect 7387 5063 7403 5097
rect 7403 5063 7421 5097
rect 7459 5063 7471 5097
rect 7471 5063 7493 5097
rect 7531 5063 7539 5097
rect 7539 5063 7565 5097
rect 7603 5063 7607 5097
rect 7607 5063 7637 5097
rect 7675 5063 7709 5097
rect 7747 5063 7777 5097
rect 7777 5063 7781 5097
rect 7819 5063 7845 5097
rect 7845 5063 7853 5097
rect 343 4955 377 4969
rect 343 4935 377 4955
rect 343 4887 377 4897
rect 343 4863 377 4887
rect 343 4819 377 4825
rect 343 4791 377 4819
rect 343 4751 377 4753
rect 343 4719 377 4751
rect 343 4649 377 4681
rect 343 4647 377 4649
rect 343 4581 377 4609
rect 343 4575 377 4581
rect 343 4513 377 4537
rect 343 4503 377 4513
rect 343 4445 377 4465
rect 343 4431 377 4445
rect 2263 4955 2297 4969
rect 2263 4935 2297 4955
rect 2263 4887 2297 4897
rect 2263 4863 2297 4887
rect 2263 4819 2297 4825
rect 2263 4791 2297 4819
rect 2263 4751 2297 4753
rect 2263 4719 2297 4751
rect 2263 4649 2297 4681
rect 2263 4647 2297 4649
rect 2263 4581 2297 4609
rect 2263 4575 2297 4581
rect 2263 4513 2297 4537
rect 2263 4503 2297 4513
rect 2263 4445 2297 4465
rect 2263 4431 2297 4445
rect 4183 4955 4217 4969
rect 4183 4935 4217 4955
rect 4183 4887 4217 4897
rect 4183 4863 4217 4887
rect 4183 4819 4217 4825
rect 4183 4791 4217 4819
rect 4183 4751 4217 4753
rect 4183 4719 4217 4751
rect 4183 4649 4217 4681
rect 4183 4647 4217 4649
rect 4183 4581 4217 4609
rect 4183 4575 4217 4581
rect 4183 4513 4217 4537
rect 4183 4503 4217 4513
rect 4183 4445 4217 4465
rect 4183 4431 4217 4445
rect 6103 4955 6137 4969
rect 6103 4935 6137 4955
rect 6103 4887 6137 4897
rect 6103 4863 6137 4887
rect 6103 4819 6137 4825
rect 6103 4791 6137 4819
rect 6103 4751 6137 4753
rect 6103 4719 6137 4751
rect 6103 4649 6137 4681
rect 6103 4647 6137 4649
rect 6103 4581 6137 4609
rect 6103 4575 6137 4581
rect 6103 4513 6137 4537
rect 6103 4503 6137 4513
rect 6103 4445 6137 4465
rect 6103 4431 6137 4445
rect 8023 4955 8057 4969
rect 8023 4935 8057 4955
rect 8023 4887 8057 4897
rect 8023 4863 8057 4887
rect 8023 4819 8057 4825
rect 8023 4791 8057 4819
rect 8023 4751 8057 4753
rect 8023 4719 8057 4751
rect 8023 4649 8057 4681
rect 8023 4647 8057 4649
rect 8023 4581 8057 4609
rect 8023 4575 8057 4581
rect 8023 4513 8057 4537
rect 8023 4503 8057 4513
rect 8023 4445 8057 4465
rect 8023 4431 8057 4445
rect 343 3635 377 3649
rect 343 3615 377 3635
rect 343 3567 377 3577
rect 343 3543 377 3567
rect 343 3499 377 3505
rect 343 3471 377 3499
rect 343 3431 377 3433
rect 343 3399 377 3431
rect 343 3329 377 3361
rect 343 3327 377 3329
rect 343 3261 377 3289
rect 343 3255 377 3261
rect 343 3193 377 3217
rect 343 3183 377 3193
rect 343 3125 377 3145
rect 343 3111 377 3125
rect 2263 3635 2297 3649
rect 2263 3615 2297 3635
rect 2263 3567 2297 3577
rect 2263 3543 2297 3567
rect 2263 3499 2297 3505
rect 2263 3471 2297 3499
rect 2263 3431 2297 3433
rect 2263 3399 2297 3431
rect 2263 3329 2297 3361
rect 2263 3327 2297 3329
rect 2263 3261 2297 3289
rect 2263 3255 2297 3261
rect 2263 3193 2297 3217
rect 2263 3183 2297 3193
rect 2263 3125 2297 3145
rect 2263 3111 2297 3125
rect 4183 3635 4217 3649
rect 4183 3615 4217 3635
rect 4183 3567 4217 3577
rect 4183 3543 4217 3567
rect 4183 3499 4217 3505
rect 4183 3471 4217 3499
rect 4183 3431 4217 3433
rect 4183 3399 4217 3431
rect 4183 3329 4217 3361
rect 4183 3327 4217 3329
rect 4183 3261 4217 3289
rect 4183 3255 4217 3261
rect 4183 3193 4217 3217
rect 4183 3183 4217 3193
rect 4183 3125 4217 3145
rect 4183 3111 4217 3125
rect 6103 3635 6137 3649
rect 6103 3615 6137 3635
rect 6103 3567 6137 3577
rect 6103 3543 6137 3567
rect 6103 3499 6137 3505
rect 6103 3471 6137 3499
rect 6103 3431 6137 3433
rect 6103 3399 6137 3431
rect 6103 3329 6137 3361
rect 6103 3327 6137 3329
rect 6103 3261 6137 3289
rect 6103 3255 6137 3261
rect 6103 3193 6137 3217
rect 6103 3183 6137 3193
rect 6103 3125 6137 3145
rect 6103 3111 6137 3125
rect 8023 3635 8057 3649
rect 8023 3615 8057 3635
rect 8023 3567 8057 3577
rect 8023 3543 8057 3567
rect 8023 3499 8057 3505
rect 8023 3471 8057 3499
rect 8023 3431 8057 3433
rect 8023 3399 8057 3431
rect 8023 3329 8057 3361
rect 8023 3327 8057 3329
rect 8023 3261 8057 3289
rect 8023 3255 8057 3261
rect 8023 3193 8057 3217
rect 8023 3183 8057 3193
rect 8023 3125 8057 3145
rect 8023 3111 8057 3125
rect 547 2983 555 3017
rect 555 2983 581 3017
rect 619 2983 623 3017
rect 623 2983 653 3017
rect 691 2983 725 3017
rect 763 2983 793 3017
rect 793 2983 797 3017
rect 835 2983 861 3017
rect 861 2983 869 3017
rect 907 2983 929 3017
rect 929 2983 941 3017
rect 979 2983 997 3017
rect 997 2983 1013 3017
rect 1051 2983 1065 3017
rect 1065 2983 1085 3017
rect 1123 2983 1133 3017
rect 1133 2983 1157 3017
rect 1195 2983 1201 3017
rect 1201 2983 1229 3017
rect 1267 2983 1269 3017
rect 1269 2983 1301 3017
rect 1339 2983 1371 3017
rect 1371 2983 1373 3017
rect 1411 2983 1439 3017
rect 1439 2983 1445 3017
rect 1483 2983 1507 3017
rect 1507 2983 1517 3017
rect 1555 2983 1575 3017
rect 1575 2983 1589 3017
rect 1627 2983 1643 3017
rect 1643 2983 1661 3017
rect 1699 2983 1711 3017
rect 1711 2983 1733 3017
rect 1771 2983 1779 3017
rect 1779 2983 1805 3017
rect 1843 2983 1847 3017
rect 1847 2983 1877 3017
rect 1915 2983 1949 3017
rect 1987 2983 2017 3017
rect 2017 2983 2021 3017
rect 2059 2983 2085 3017
rect 2085 2983 2093 3017
rect 2467 2983 2475 3017
rect 2475 2983 2501 3017
rect 2539 2983 2543 3017
rect 2543 2983 2573 3017
rect 2611 2983 2645 3017
rect 2683 2983 2713 3017
rect 2713 2983 2717 3017
rect 2755 2983 2781 3017
rect 2781 2983 2789 3017
rect 2827 2983 2849 3017
rect 2849 2983 2861 3017
rect 2899 2983 2917 3017
rect 2917 2983 2933 3017
rect 2971 2983 2985 3017
rect 2985 2983 3005 3017
rect 3043 2983 3053 3017
rect 3053 2983 3077 3017
rect 3115 2983 3121 3017
rect 3121 2983 3149 3017
rect 3187 2983 3189 3017
rect 3189 2983 3221 3017
rect 3259 2983 3291 3017
rect 3291 2983 3293 3017
rect 3331 2983 3359 3017
rect 3359 2983 3365 3017
rect 3403 2983 3427 3017
rect 3427 2983 3437 3017
rect 3475 2983 3495 3017
rect 3495 2983 3509 3017
rect 3547 2983 3563 3017
rect 3563 2983 3581 3017
rect 3619 2983 3631 3017
rect 3631 2983 3653 3017
rect 3691 2983 3699 3017
rect 3699 2983 3725 3017
rect 3763 2983 3767 3017
rect 3767 2983 3797 3017
rect 3835 2983 3869 3017
rect 3907 2983 3937 3017
rect 3937 2983 3941 3017
rect 3979 2983 4005 3017
rect 4005 2983 4013 3017
rect 4387 2983 4395 3017
rect 4395 2983 4421 3017
rect 4459 2983 4463 3017
rect 4463 2983 4493 3017
rect 4531 2983 4565 3017
rect 4603 2983 4633 3017
rect 4633 2983 4637 3017
rect 4675 2983 4701 3017
rect 4701 2983 4709 3017
rect 4747 2983 4769 3017
rect 4769 2983 4781 3017
rect 4819 2983 4837 3017
rect 4837 2983 4853 3017
rect 4891 2983 4905 3017
rect 4905 2983 4925 3017
rect 4963 2983 4973 3017
rect 4973 2983 4997 3017
rect 5035 2983 5041 3017
rect 5041 2983 5069 3017
rect 5107 2983 5109 3017
rect 5109 2983 5141 3017
rect 5179 2983 5211 3017
rect 5211 2983 5213 3017
rect 5251 2983 5279 3017
rect 5279 2983 5285 3017
rect 5323 2983 5347 3017
rect 5347 2983 5357 3017
rect 5395 2983 5415 3017
rect 5415 2983 5429 3017
rect 5467 2983 5483 3017
rect 5483 2983 5501 3017
rect 5539 2983 5551 3017
rect 5551 2983 5573 3017
rect 5611 2983 5619 3017
rect 5619 2983 5645 3017
rect 5683 2983 5687 3017
rect 5687 2983 5717 3017
rect 5755 2983 5789 3017
rect 5827 2983 5857 3017
rect 5857 2983 5861 3017
rect 5899 2983 5925 3017
rect 5925 2983 5933 3017
rect 6307 2983 6315 3017
rect 6315 2983 6341 3017
rect 6379 2983 6383 3017
rect 6383 2983 6413 3017
rect 6451 2983 6485 3017
rect 6523 2983 6553 3017
rect 6553 2983 6557 3017
rect 6595 2983 6621 3017
rect 6621 2983 6629 3017
rect 6667 2983 6689 3017
rect 6689 2983 6701 3017
rect 6739 2983 6757 3017
rect 6757 2983 6773 3017
rect 6811 2983 6825 3017
rect 6825 2983 6845 3017
rect 6883 2983 6893 3017
rect 6893 2983 6917 3017
rect 6955 2983 6961 3017
rect 6961 2983 6989 3017
rect 7027 2983 7029 3017
rect 7029 2983 7061 3017
rect 7099 2983 7131 3017
rect 7131 2983 7133 3017
rect 7171 2983 7199 3017
rect 7199 2983 7205 3017
rect 7243 2983 7267 3017
rect 7267 2983 7277 3017
rect 7315 2983 7335 3017
rect 7335 2983 7349 3017
rect 7387 2983 7403 3017
rect 7403 2983 7421 3017
rect 7459 2983 7471 3017
rect 7471 2983 7493 3017
rect 7531 2983 7539 3017
rect 7539 2983 7565 3017
rect 7603 2983 7607 3017
rect 7607 2983 7637 3017
rect 7675 2983 7709 3017
rect 7747 2983 7777 3017
rect 7777 2983 7781 3017
rect 7819 2983 7845 3017
rect 7845 2983 7853 3017
rect 343 2195 377 2209
rect 343 2175 377 2195
rect 343 2127 377 2137
rect 343 2103 377 2127
rect 343 2059 377 2065
rect 343 2031 377 2059
rect 343 1991 377 1993
rect 343 1959 377 1991
rect 343 1889 377 1921
rect 343 1887 377 1889
rect 343 1821 377 1849
rect 343 1815 377 1821
rect 343 1753 377 1777
rect 343 1743 377 1753
rect 343 1685 377 1705
rect 343 1671 377 1685
rect 2263 2195 2297 2209
rect 2263 2175 2297 2195
rect 2263 2127 2297 2137
rect 2263 2103 2297 2127
rect 2263 2059 2297 2065
rect 2263 2031 2297 2059
rect 2263 1991 2297 1993
rect 2263 1959 2297 1991
rect 2263 1889 2297 1921
rect 2263 1887 2297 1889
rect 2263 1821 2297 1849
rect 2263 1815 2297 1821
rect 2263 1753 2297 1777
rect 2263 1743 2297 1753
rect 2263 1685 2297 1705
rect 2263 1671 2297 1685
rect 4183 2195 4217 2209
rect 4183 2175 4217 2195
rect 4183 2127 4217 2137
rect 4183 2103 4217 2127
rect 4183 2059 4217 2065
rect 4183 2031 4217 2059
rect 4183 1991 4217 1993
rect 4183 1959 4217 1991
rect 4183 1889 4217 1921
rect 4183 1887 4217 1889
rect 4183 1821 4217 1849
rect 4183 1815 4217 1821
rect 4183 1753 4217 1777
rect 4183 1743 4217 1753
rect 4183 1685 4217 1705
rect 4183 1671 4217 1685
rect 6103 2195 6137 2209
rect 6103 2175 6137 2195
rect 6103 2127 6137 2137
rect 6103 2103 6137 2127
rect 6103 2059 6137 2065
rect 6103 2031 6137 2059
rect 6103 1991 6137 1993
rect 6103 1959 6137 1991
rect 6103 1889 6137 1921
rect 6103 1887 6137 1889
rect 6103 1821 6137 1849
rect 6103 1815 6137 1821
rect 6103 1753 6137 1777
rect 6103 1743 6137 1753
rect 6103 1685 6137 1705
rect 6103 1671 6137 1685
rect 8023 2195 8057 2209
rect 8023 2175 8057 2195
rect 8023 2127 8057 2137
rect 8023 2103 8057 2127
rect 8023 2059 8057 2065
rect 8023 2031 8057 2059
rect 8023 1991 8057 1993
rect 8023 1959 8057 1991
rect 8023 1889 8057 1921
rect 8023 1887 8057 1889
rect 8023 1821 8057 1849
rect 8023 1815 8057 1821
rect 8023 1753 8057 1777
rect 8023 1743 8057 1753
rect 8023 1685 8057 1705
rect 8023 1671 8057 1685
rect 547 1543 555 1577
rect 555 1543 581 1577
rect 619 1543 623 1577
rect 623 1543 653 1577
rect 691 1543 725 1577
rect 763 1543 793 1577
rect 793 1543 797 1577
rect 835 1543 861 1577
rect 861 1543 869 1577
rect 907 1543 929 1577
rect 929 1543 941 1577
rect 979 1543 997 1577
rect 997 1543 1013 1577
rect 1051 1543 1065 1577
rect 1065 1543 1085 1577
rect 1123 1543 1133 1577
rect 1133 1543 1157 1577
rect 1195 1543 1201 1577
rect 1201 1543 1229 1577
rect 1267 1543 1269 1577
rect 1269 1543 1301 1577
rect 1339 1543 1371 1577
rect 1371 1543 1373 1577
rect 1411 1543 1439 1577
rect 1439 1543 1445 1577
rect 1483 1543 1507 1577
rect 1507 1543 1517 1577
rect 1555 1543 1575 1577
rect 1575 1543 1589 1577
rect 1627 1543 1643 1577
rect 1643 1543 1661 1577
rect 1699 1543 1711 1577
rect 1711 1543 1733 1577
rect 1771 1543 1779 1577
rect 1779 1543 1805 1577
rect 1843 1543 1847 1577
rect 1847 1543 1877 1577
rect 1915 1543 1949 1577
rect 1987 1543 2017 1577
rect 2017 1543 2021 1577
rect 2059 1543 2085 1577
rect 2085 1543 2093 1577
rect 2467 1543 2475 1577
rect 2475 1543 2501 1577
rect 2539 1543 2543 1577
rect 2543 1543 2573 1577
rect 2611 1543 2645 1577
rect 2683 1543 2713 1577
rect 2713 1543 2717 1577
rect 2755 1543 2781 1577
rect 2781 1543 2789 1577
rect 2827 1543 2849 1577
rect 2849 1543 2861 1577
rect 2899 1543 2917 1577
rect 2917 1543 2933 1577
rect 2971 1543 2985 1577
rect 2985 1543 3005 1577
rect 3043 1543 3053 1577
rect 3053 1543 3077 1577
rect 3115 1543 3121 1577
rect 3121 1543 3149 1577
rect 3187 1543 3189 1577
rect 3189 1543 3221 1577
rect 3259 1543 3291 1577
rect 3291 1543 3293 1577
rect 3331 1543 3359 1577
rect 3359 1543 3365 1577
rect 3403 1543 3427 1577
rect 3427 1543 3437 1577
rect 3475 1543 3495 1577
rect 3495 1543 3509 1577
rect 3547 1543 3563 1577
rect 3563 1543 3581 1577
rect 3619 1543 3631 1577
rect 3631 1543 3653 1577
rect 3691 1543 3699 1577
rect 3699 1543 3725 1577
rect 3763 1543 3767 1577
rect 3767 1543 3797 1577
rect 3835 1543 3869 1577
rect 3907 1543 3937 1577
rect 3937 1543 3941 1577
rect 3979 1543 4005 1577
rect 4005 1543 4013 1577
rect 4387 1543 4395 1577
rect 4395 1543 4421 1577
rect 4459 1543 4463 1577
rect 4463 1543 4493 1577
rect 4531 1543 4565 1577
rect 4603 1543 4633 1577
rect 4633 1543 4637 1577
rect 4675 1543 4701 1577
rect 4701 1543 4709 1577
rect 4747 1543 4769 1577
rect 4769 1543 4781 1577
rect 4819 1543 4837 1577
rect 4837 1543 4853 1577
rect 4891 1543 4905 1577
rect 4905 1543 4925 1577
rect 4963 1543 4973 1577
rect 4973 1543 4997 1577
rect 5035 1543 5041 1577
rect 5041 1543 5069 1577
rect 5107 1543 5109 1577
rect 5109 1543 5141 1577
rect 5179 1543 5211 1577
rect 5211 1543 5213 1577
rect 5251 1543 5279 1577
rect 5279 1543 5285 1577
rect 5323 1543 5347 1577
rect 5347 1543 5357 1577
rect 5395 1543 5415 1577
rect 5415 1543 5429 1577
rect 5467 1543 5483 1577
rect 5483 1543 5501 1577
rect 5539 1543 5551 1577
rect 5551 1543 5573 1577
rect 5611 1543 5619 1577
rect 5619 1543 5645 1577
rect 5683 1543 5687 1577
rect 5687 1543 5717 1577
rect 5755 1543 5789 1577
rect 5827 1543 5857 1577
rect 5857 1543 5861 1577
rect 5899 1543 5925 1577
rect 5925 1543 5933 1577
rect 6307 1543 6315 1577
rect 6315 1543 6341 1577
rect 6379 1543 6383 1577
rect 6383 1543 6413 1577
rect 6451 1543 6485 1577
rect 6523 1543 6553 1577
rect 6553 1543 6557 1577
rect 6595 1543 6621 1577
rect 6621 1543 6629 1577
rect 6667 1543 6689 1577
rect 6689 1543 6701 1577
rect 6739 1543 6757 1577
rect 6757 1543 6773 1577
rect 6811 1543 6825 1577
rect 6825 1543 6845 1577
rect 6883 1543 6893 1577
rect 6893 1543 6917 1577
rect 6955 1543 6961 1577
rect 6961 1543 6989 1577
rect 7027 1543 7029 1577
rect 7029 1543 7061 1577
rect 7099 1543 7131 1577
rect 7131 1543 7133 1577
rect 7171 1543 7199 1577
rect 7199 1543 7205 1577
rect 7243 1543 7267 1577
rect 7267 1543 7277 1577
rect 7315 1543 7335 1577
rect 7335 1543 7349 1577
rect 7387 1543 7403 1577
rect 7403 1543 7421 1577
rect 7459 1543 7471 1577
rect 7471 1543 7493 1577
rect 7531 1543 7539 1577
rect 7539 1543 7565 1577
rect 7603 1543 7607 1577
rect 7607 1543 7637 1577
rect 7675 1543 7709 1577
rect 7747 1543 7777 1577
rect 7777 1543 7781 1577
rect 7819 1543 7845 1577
rect 7845 1543 7853 1577
rect 183 903 217 937
rect 343 903 377 937
rect 503 903 537 937
rect 663 903 697 937
rect 823 903 857 937
rect 983 903 1017 937
rect 1143 903 1177 937
rect 1463 903 1497 937
rect 1623 903 1657 937
rect 1783 903 1817 937
rect 1943 903 1977 937
rect 2103 903 2137 937
rect 2263 903 2297 937
rect 2423 903 2457 937
rect 2583 903 2617 937
rect 2743 903 2777 937
rect 2903 903 2937 937
rect 3063 903 3097 937
rect 3383 903 3417 937
rect 3543 903 3577 937
rect 3703 903 3737 937
rect 3863 903 3897 937
rect 4023 903 4057 937
rect 4183 903 4217 937
rect 4343 903 4377 937
rect 4503 903 4537 937
rect 4663 903 4697 937
rect 4823 903 4857 937
rect 4983 903 5017 937
rect 5303 903 5337 937
rect 5463 903 5497 937
rect 5623 903 5657 937
rect 5783 903 5817 937
rect 5943 903 5977 937
rect 6103 903 6137 937
rect 6263 903 6297 937
rect 6423 903 6457 937
rect 6583 903 6617 937
rect 6743 903 6777 937
rect 6903 903 6937 937
rect 7223 903 7257 937
rect 7383 903 7417 937
rect 7543 903 7577 937
rect 7703 903 7737 937
rect 7863 903 7897 937
rect 8183 903 8217 937
rect 547 423 555 457
rect 555 423 581 457
rect 619 423 623 457
rect 623 423 653 457
rect 691 423 725 457
rect 763 423 793 457
rect 793 423 797 457
rect 835 423 861 457
rect 861 423 869 457
rect 907 423 929 457
rect 929 423 941 457
rect 979 423 997 457
rect 997 423 1013 457
rect 1051 423 1065 457
rect 1065 423 1085 457
rect 1123 423 1133 457
rect 1133 423 1157 457
rect 1195 423 1201 457
rect 1201 423 1229 457
rect 1267 423 1269 457
rect 1269 423 1301 457
rect 1339 423 1371 457
rect 1371 423 1373 457
rect 1411 423 1439 457
rect 1439 423 1445 457
rect 1483 423 1507 457
rect 1507 423 1517 457
rect 1555 423 1575 457
rect 1575 423 1589 457
rect 1627 423 1643 457
rect 1643 423 1661 457
rect 1699 423 1711 457
rect 1711 423 1733 457
rect 1771 423 1779 457
rect 1779 423 1805 457
rect 1843 423 1847 457
rect 1847 423 1877 457
rect 1915 423 1949 457
rect 1987 423 2017 457
rect 2017 423 2021 457
rect 2059 423 2085 457
rect 2085 423 2093 457
rect 2467 423 2475 457
rect 2475 423 2501 457
rect 2539 423 2543 457
rect 2543 423 2573 457
rect 2611 423 2645 457
rect 2683 423 2713 457
rect 2713 423 2717 457
rect 2755 423 2781 457
rect 2781 423 2789 457
rect 2827 423 2849 457
rect 2849 423 2861 457
rect 2899 423 2917 457
rect 2917 423 2933 457
rect 2971 423 2985 457
rect 2985 423 3005 457
rect 3043 423 3053 457
rect 3053 423 3077 457
rect 3115 423 3121 457
rect 3121 423 3149 457
rect 3187 423 3189 457
rect 3189 423 3221 457
rect 3259 423 3291 457
rect 3291 423 3293 457
rect 3331 423 3359 457
rect 3359 423 3365 457
rect 3403 423 3427 457
rect 3427 423 3437 457
rect 3475 423 3495 457
rect 3495 423 3509 457
rect 3547 423 3563 457
rect 3563 423 3581 457
rect 3619 423 3631 457
rect 3631 423 3653 457
rect 3691 423 3699 457
rect 3699 423 3725 457
rect 3763 423 3767 457
rect 3767 423 3797 457
rect 3835 423 3869 457
rect 3907 423 3937 457
rect 3937 423 3941 457
rect 3979 423 4005 457
rect 4005 423 4013 457
rect 4387 423 4395 457
rect 4395 423 4421 457
rect 4459 423 4463 457
rect 4463 423 4493 457
rect 4531 423 4565 457
rect 4603 423 4633 457
rect 4633 423 4637 457
rect 4675 423 4701 457
rect 4701 423 4709 457
rect 4747 423 4769 457
rect 4769 423 4781 457
rect 4819 423 4837 457
rect 4837 423 4853 457
rect 4891 423 4905 457
rect 4905 423 4925 457
rect 4963 423 4973 457
rect 4973 423 4997 457
rect 5035 423 5041 457
rect 5041 423 5069 457
rect 5107 423 5109 457
rect 5109 423 5141 457
rect 5179 423 5211 457
rect 5211 423 5213 457
rect 5251 423 5279 457
rect 5279 423 5285 457
rect 5323 423 5347 457
rect 5347 423 5357 457
rect 5395 423 5415 457
rect 5415 423 5429 457
rect 5467 423 5483 457
rect 5483 423 5501 457
rect 5539 423 5551 457
rect 5551 423 5573 457
rect 5611 423 5619 457
rect 5619 423 5645 457
rect 5683 423 5687 457
rect 5687 423 5717 457
rect 5755 423 5789 457
rect 5827 423 5857 457
rect 5857 423 5861 457
rect 5899 423 5925 457
rect 5925 423 5933 457
rect 6307 423 6315 457
rect 6315 423 6341 457
rect 6379 423 6383 457
rect 6383 423 6413 457
rect 6451 423 6485 457
rect 6523 423 6553 457
rect 6553 423 6557 457
rect 6595 423 6621 457
rect 6621 423 6629 457
rect 6667 423 6689 457
rect 6689 423 6701 457
rect 6739 423 6757 457
rect 6757 423 6773 457
rect 6811 423 6825 457
rect 6825 423 6845 457
rect 6883 423 6893 457
rect 6893 423 6917 457
rect 6955 423 6961 457
rect 6961 423 6989 457
rect 7027 423 7029 457
rect 7029 423 7061 457
rect 7099 423 7131 457
rect 7131 423 7133 457
rect 7171 423 7199 457
rect 7199 423 7205 457
rect 7243 423 7267 457
rect 7267 423 7277 457
rect 7315 423 7335 457
rect 7335 423 7349 457
rect 7387 423 7403 457
rect 7403 423 7421 457
rect 7459 423 7471 457
rect 7471 423 7493 457
rect 7531 423 7539 457
rect 7539 423 7565 457
rect 7603 423 7607 457
rect 7607 423 7637 457
rect 7675 423 7709 457
rect 7747 423 7777 457
rect 7777 423 7781 457
rect 7819 423 7845 457
rect 7845 423 7853 457
rect 343 311 377 313
rect 343 279 377 311
rect 343 209 377 241
rect 343 207 377 209
rect 2263 311 2297 313
rect 2263 279 2297 311
rect 2263 209 2297 241
rect 2263 207 2297 209
rect 4183 311 4217 313
rect 4183 279 4217 311
rect 4183 209 4217 241
rect 4183 207 4217 209
rect 6103 311 6137 313
rect 6103 279 6137 311
rect 6103 209 6137 241
rect 6103 207 6137 209
rect 8023 311 8057 313
rect 8023 279 8057 311
rect 8023 209 8057 241
rect 8023 207 8057 209
rect 183 -137 217 -103
rect 343 -137 377 -103
rect 503 -137 537 -103
rect 663 -137 697 -103
rect 823 -137 857 -103
rect 983 -137 1017 -103
rect 1143 -137 1177 -103
rect 1463 -137 1497 -103
rect 1623 -137 1657 -103
rect 1783 -137 1817 -103
rect 1943 -137 1977 -103
rect 2103 -137 2137 -103
rect 2263 -137 2297 -103
rect 2423 -137 2457 -103
rect 2583 -137 2617 -103
rect 2743 -137 2777 -103
rect 2903 -137 2937 -103
rect 3063 -137 3097 -103
rect 3383 -137 3417 -103
rect 3543 -137 3577 -103
rect 3703 -137 3737 -103
rect 3863 -137 3897 -103
rect 4023 -137 4057 -103
rect 4183 -137 4217 -103
rect 4343 -137 4377 -103
rect 4503 -137 4537 -103
rect 4663 -137 4697 -103
rect 4823 -137 4857 -103
rect 4983 -137 5017 -103
rect 5303 -137 5337 -103
rect 5463 -137 5497 -103
rect 5623 -137 5657 -103
rect 5783 -137 5817 -103
rect 5943 -137 5977 -103
rect 6103 -137 6137 -103
rect 6263 -137 6297 -103
rect 6423 -137 6457 -103
rect 6583 -137 6617 -103
rect 6743 -137 6777 -103
rect 6903 -137 6937 -103
rect 7223 -137 7257 -103
rect 7383 -137 7417 -103
rect 7543 -137 7577 -103
rect 7703 -137 7737 -103
rect 7863 -137 7897 -103
rect 8183 -137 8217 -103
rect 547 -617 555 -583
rect 555 -617 581 -583
rect 619 -617 623 -583
rect 623 -617 653 -583
rect 691 -617 725 -583
rect 763 -617 793 -583
rect 793 -617 797 -583
rect 835 -617 861 -583
rect 861 -617 869 -583
rect 907 -617 929 -583
rect 929 -617 941 -583
rect 979 -617 997 -583
rect 997 -617 1013 -583
rect 1051 -617 1065 -583
rect 1065 -617 1085 -583
rect 1123 -617 1133 -583
rect 1133 -617 1157 -583
rect 1195 -617 1201 -583
rect 1201 -617 1229 -583
rect 1267 -617 1269 -583
rect 1269 -617 1301 -583
rect 1339 -617 1371 -583
rect 1371 -617 1373 -583
rect 1411 -617 1439 -583
rect 1439 -617 1445 -583
rect 1483 -617 1507 -583
rect 1507 -617 1517 -583
rect 1555 -617 1575 -583
rect 1575 -617 1589 -583
rect 1627 -617 1643 -583
rect 1643 -617 1661 -583
rect 1699 -617 1711 -583
rect 1711 -617 1733 -583
rect 1771 -617 1779 -583
rect 1779 -617 1805 -583
rect 1843 -617 1847 -583
rect 1847 -617 1877 -583
rect 1915 -617 1949 -583
rect 1987 -617 2017 -583
rect 2017 -617 2021 -583
rect 2059 -617 2085 -583
rect 2085 -617 2093 -583
rect 2467 -617 2475 -583
rect 2475 -617 2501 -583
rect 2539 -617 2543 -583
rect 2543 -617 2573 -583
rect 2611 -617 2645 -583
rect 2683 -617 2713 -583
rect 2713 -617 2717 -583
rect 2755 -617 2781 -583
rect 2781 -617 2789 -583
rect 2827 -617 2849 -583
rect 2849 -617 2861 -583
rect 2899 -617 2917 -583
rect 2917 -617 2933 -583
rect 2971 -617 2985 -583
rect 2985 -617 3005 -583
rect 3043 -617 3053 -583
rect 3053 -617 3077 -583
rect 3115 -617 3121 -583
rect 3121 -617 3149 -583
rect 3187 -617 3189 -583
rect 3189 -617 3221 -583
rect 3259 -617 3291 -583
rect 3291 -617 3293 -583
rect 3331 -617 3359 -583
rect 3359 -617 3365 -583
rect 3403 -617 3427 -583
rect 3427 -617 3437 -583
rect 3475 -617 3495 -583
rect 3495 -617 3509 -583
rect 3547 -617 3563 -583
rect 3563 -617 3581 -583
rect 3619 -617 3631 -583
rect 3631 -617 3653 -583
rect 3691 -617 3699 -583
rect 3699 -617 3725 -583
rect 3763 -617 3767 -583
rect 3767 -617 3797 -583
rect 3835 -617 3869 -583
rect 3907 -617 3937 -583
rect 3937 -617 3941 -583
rect 3979 -617 4005 -583
rect 4005 -617 4013 -583
rect 4387 -617 4395 -583
rect 4395 -617 4421 -583
rect 4459 -617 4463 -583
rect 4463 -617 4493 -583
rect 4531 -617 4565 -583
rect 4603 -617 4633 -583
rect 4633 -617 4637 -583
rect 4675 -617 4701 -583
rect 4701 -617 4709 -583
rect 4747 -617 4769 -583
rect 4769 -617 4781 -583
rect 4819 -617 4837 -583
rect 4837 -617 4853 -583
rect 4891 -617 4905 -583
rect 4905 -617 4925 -583
rect 4963 -617 4973 -583
rect 4973 -617 4997 -583
rect 5035 -617 5041 -583
rect 5041 -617 5069 -583
rect 5107 -617 5109 -583
rect 5109 -617 5141 -583
rect 5179 -617 5211 -583
rect 5211 -617 5213 -583
rect 5251 -617 5279 -583
rect 5279 -617 5285 -583
rect 5323 -617 5347 -583
rect 5347 -617 5357 -583
rect 5395 -617 5415 -583
rect 5415 -617 5429 -583
rect 5467 -617 5483 -583
rect 5483 -617 5501 -583
rect 5539 -617 5551 -583
rect 5551 -617 5573 -583
rect 5611 -617 5619 -583
rect 5619 -617 5645 -583
rect 5683 -617 5687 -583
rect 5687 -617 5717 -583
rect 5755 -617 5789 -583
rect 5827 -617 5857 -583
rect 5857 -617 5861 -583
rect 5899 -617 5925 -583
rect 5925 -617 5933 -583
rect 6307 -617 6315 -583
rect 6315 -617 6341 -583
rect 6379 -617 6383 -583
rect 6383 -617 6413 -583
rect 6451 -617 6485 -583
rect 6523 -617 6553 -583
rect 6553 -617 6557 -583
rect 6595 -617 6621 -583
rect 6621 -617 6629 -583
rect 6667 -617 6689 -583
rect 6689 -617 6701 -583
rect 6739 -617 6757 -583
rect 6757 -617 6773 -583
rect 6811 -617 6825 -583
rect 6825 -617 6845 -583
rect 6883 -617 6893 -583
rect 6893 -617 6917 -583
rect 6955 -617 6961 -583
rect 6961 -617 6989 -583
rect 7027 -617 7029 -583
rect 7029 -617 7061 -583
rect 7099 -617 7131 -583
rect 7131 -617 7133 -583
rect 7171 -617 7199 -583
rect 7199 -617 7205 -583
rect 7243 -617 7267 -583
rect 7267 -617 7277 -583
rect 7315 -617 7335 -583
rect 7335 -617 7349 -583
rect 7387 -617 7403 -583
rect 7403 -617 7421 -583
rect 7459 -617 7471 -583
rect 7471 -617 7493 -583
rect 7531 -617 7539 -583
rect 7539 -617 7565 -583
rect 7603 -617 7607 -583
rect 7607 -617 7637 -583
rect 7675 -617 7709 -583
rect 7747 -617 7777 -583
rect 7777 -617 7781 -583
rect 7819 -617 7845 -583
rect 7845 -617 7853 -583
rect 343 -729 377 -727
rect 343 -761 377 -729
rect 343 -831 377 -799
rect 343 -833 377 -831
rect 2263 -729 2297 -727
rect 2263 -761 2297 -729
rect 2263 -831 2297 -799
rect 2263 -833 2297 -831
rect 4183 -729 4217 -727
rect 4183 -761 4217 -729
rect 4183 -831 4217 -799
rect 4183 -833 4217 -831
rect 6103 -729 6137 -727
rect 6103 -761 6137 -729
rect 6103 -831 6137 -799
rect 6103 -833 6137 -831
rect 8023 -729 8057 -727
rect 8023 -761 8057 -729
rect 8023 -831 8057 -799
rect 8023 -833 8057 -831
<< metal1 >>
rect 320 9729 400 9760
rect 320 9714 343 9729
rect 377 9714 400 9729
rect 320 9662 334 9714
rect 386 9662 400 9714
rect 320 9657 400 9662
rect 320 9650 343 9657
rect 377 9650 400 9657
rect 320 9598 334 9650
rect 386 9598 400 9650
rect 320 9586 400 9598
rect 320 9534 334 9586
rect 386 9534 400 9586
rect 320 9522 400 9534
rect 320 9470 334 9522
rect 386 9470 400 9522
rect 320 9458 400 9470
rect 320 9406 334 9458
rect 386 9406 400 9458
rect 320 9369 400 9406
rect 320 9335 343 9369
rect 377 9335 400 9369
rect 320 9297 400 9335
rect 320 9263 343 9297
rect 377 9263 400 9297
rect 320 9225 400 9263
rect 320 9191 343 9225
rect 377 9191 400 9225
rect 320 9160 400 9191
rect 2240 9729 2320 9760
rect 2240 9695 2263 9729
rect 2297 9695 2320 9729
rect 2240 9657 2320 9695
rect 2240 9623 2263 9657
rect 2297 9623 2320 9657
rect 2240 9585 2320 9623
rect 2240 9551 2263 9585
rect 2297 9551 2320 9585
rect 2240 9513 2320 9551
rect 2240 9479 2263 9513
rect 2297 9479 2320 9513
rect 2240 9441 2320 9479
rect 2240 9407 2263 9441
rect 2297 9407 2320 9441
rect 2240 9369 2320 9407
rect 2240 9335 2263 9369
rect 2297 9335 2320 9369
rect 2240 9297 2320 9335
rect 2240 9263 2263 9297
rect 2297 9263 2320 9297
rect 2240 9225 2320 9263
rect 2240 9191 2263 9225
rect 2297 9191 2320 9225
rect 2240 9160 2320 9191
rect 4160 9729 4240 9760
rect 4160 9695 4183 9729
rect 4217 9695 4240 9729
rect 4160 9657 4240 9695
rect 4160 9623 4183 9657
rect 4217 9623 4240 9657
rect 4160 9585 4240 9623
rect 4160 9551 4183 9585
rect 4217 9551 4240 9585
rect 4160 9513 4240 9551
rect 4160 9479 4183 9513
rect 4217 9479 4240 9513
rect 4160 9441 4240 9479
rect 4160 9407 4183 9441
rect 4217 9407 4240 9441
rect 4160 9369 4240 9407
rect 4160 9335 4183 9369
rect 4217 9335 4240 9369
rect 4160 9297 4240 9335
rect 4160 9263 4183 9297
rect 4217 9263 4240 9297
rect 4160 9225 4240 9263
rect 4160 9191 4183 9225
rect 4217 9191 4240 9225
rect 4160 9160 4240 9191
rect 6080 9729 6160 9760
rect 6080 9695 6103 9729
rect 6137 9695 6160 9729
rect 6080 9657 6160 9695
rect 6080 9623 6103 9657
rect 6137 9623 6160 9657
rect 6080 9585 6160 9623
rect 6080 9551 6103 9585
rect 6137 9551 6160 9585
rect 6080 9513 6160 9551
rect 6080 9479 6103 9513
rect 6137 9479 6160 9513
rect 6080 9441 6160 9479
rect 6080 9407 6103 9441
rect 6137 9407 6160 9441
rect 6080 9369 6160 9407
rect 6080 9335 6103 9369
rect 6137 9335 6160 9369
rect 6080 9297 6160 9335
rect 6080 9263 6103 9297
rect 6137 9263 6160 9297
rect 6080 9225 6160 9263
rect 6080 9191 6103 9225
rect 6137 9191 6160 9225
rect 6080 9160 6160 9191
rect 8000 9729 8080 9760
rect 8000 9695 8023 9729
rect 8057 9695 8080 9729
rect 8000 9657 8080 9695
rect 8000 9623 8023 9657
rect 8057 9623 8080 9657
rect 8000 9585 8080 9623
rect 8000 9551 8023 9585
rect 8057 9551 8080 9585
rect 8000 9513 8080 9551
rect 8000 9479 8023 9513
rect 8057 9479 8080 9513
rect 8000 9441 8080 9479
rect 8000 9407 8023 9441
rect 8057 9407 8080 9441
rect 8000 9369 8080 9407
rect 8000 9335 8023 9369
rect 8057 9335 8080 9369
rect 8000 9297 8080 9335
rect 8000 9263 8023 9297
rect 8057 9263 8080 9297
rect 8000 9225 8080 9263
rect 8000 9191 8023 9225
rect 8057 9191 8080 9225
rect 520 9097 2120 9120
rect 520 9063 547 9097
rect 581 9063 619 9097
rect 653 9063 691 9097
rect 725 9063 763 9097
rect 797 9063 835 9097
rect 869 9063 907 9097
rect 941 9063 979 9097
rect 1013 9063 1051 9097
rect 1085 9063 1123 9097
rect 1157 9063 1195 9097
rect 1229 9063 1267 9097
rect 1301 9063 1339 9097
rect 1373 9063 1411 9097
rect 1445 9063 1483 9097
rect 1517 9063 1555 9097
rect 1589 9063 1627 9097
rect 1661 9063 1699 9097
rect 1733 9063 1771 9097
rect 1805 9063 1843 9097
rect 1877 9063 1915 9097
rect 1949 9063 1987 9097
rect 2021 9063 2059 9097
rect 2093 9063 2120 9097
rect 520 9040 2120 9063
rect 2440 9097 4040 9120
rect 2440 9063 2467 9097
rect 2501 9063 2539 9097
rect 2573 9063 2611 9097
rect 2645 9063 2683 9097
rect 2717 9063 2755 9097
rect 2789 9063 2827 9097
rect 2861 9063 2899 9097
rect 2933 9063 2971 9097
rect 3005 9063 3043 9097
rect 3077 9063 3115 9097
rect 3149 9063 3187 9097
rect 3221 9063 3259 9097
rect 3293 9063 3331 9097
rect 3365 9063 3403 9097
rect 3437 9063 3475 9097
rect 3509 9063 3547 9097
rect 3581 9063 3619 9097
rect 3653 9063 3691 9097
rect 3725 9063 3763 9097
rect 3797 9063 3835 9097
rect 3869 9063 3907 9097
rect 3941 9063 3979 9097
rect 4013 9063 4040 9097
rect 2440 9040 4040 9063
rect 4360 9097 5960 9120
rect 4360 9063 4387 9097
rect 4421 9063 4459 9097
rect 4493 9063 4531 9097
rect 4565 9063 4603 9097
rect 4637 9063 4675 9097
rect 4709 9063 4747 9097
rect 4781 9063 4819 9097
rect 4853 9063 4891 9097
rect 4925 9063 4963 9097
rect 4997 9063 5035 9097
rect 5069 9063 5107 9097
rect 5141 9063 5179 9097
rect 5213 9063 5251 9097
rect 5285 9063 5323 9097
rect 5357 9063 5395 9097
rect 5429 9063 5467 9097
rect 5501 9063 5539 9097
rect 5573 9063 5611 9097
rect 5645 9063 5683 9097
rect 5717 9063 5755 9097
rect 5789 9063 5827 9097
rect 5861 9063 5899 9097
rect 5933 9063 5960 9097
rect 4360 9040 5960 9063
rect 6280 9097 7880 9120
rect 6280 9063 6307 9097
rect 6341 9063 6379 9097
rect 6413 9063 6451 9097
rect 6485 9063 6523 9097
rect 6557 9063 6595 9097
rect 6629 9063 6667 9097
rect 6701 9063 6739 9097
rect 6773 9063 6811 9097
rect 6845 9063 6883 9097
rect 6917 9063 6955 9097
rect 6989 9063 7027 9097
rect 7061 9063 7099 9097
rect 7133 9063 7171 9097
rect 7205 9063 7243 9097
rect 7277 9063 7315 9097
rect 7349 9063 7387 9097
rect 7421 9063 7459 9097
rect 7493 9063 7531 9097
rect 7565 9063 7603 9097
rect 7637 9063 7675 9097
rect 7709 9063 7747 9097
rect 7781 9063 7819 9097
rect 7853 9063 7880 9097
rect 6280 9040 7880 9063
rect 1280 8626 1360 9040
rect 1280 8574 1294 8626
rect 1346 8574 1360 8626
rect 1280 8560 1360 8574
rect 3200 8626 3280 9040
rect 3200 8574 3214 8626
rect 3266 8574 3280 8626
rect 3200 8560 3280 8574
rect 5120 8626 5200 9040
rect 5120 8574 5134 8626
rect 5186 8574 5200 8626
rect 5120 8560 5200 8574
rect 7040 8626 7120 9040
rect 7040 8574 7054 8626
rect 7106 8574 7120 8626
rect 7040 8560 7120 8574
rect 8000 8626 8080 9191
rect 8000 8574 8014 8626
rect 8066 8574 8080 8626
rect 160 8466 240 8480
rect 160 8414 174 8466
rect 226 8414 240 8466
rect 160 8400 240 8414
rect 160 8306 240 8320
rect 160 8254 174 8306
rect 226 8254 240 8306
rect 160 8240 240 8254
rect 1280 8146 1360 8160
rect 1280 8094 1294 8146
rect 1346 8094 1360 8146
rect 1280 7840 1360 8094
rect 3200 8146 3280 8160
rect 3200 8094 3214 8146
rect 3266 8094 3280 8146
rect 3200 7840 3280 8094
rect 5120 8146 5200 8160
rect 5120 8094 5134 8146
rect 5186 8094 5200 8146
rect 5120 7840 5200 8094
rect 7040 8146 7120 8160
rect 7040 8094 7054 8146
rect 7106 8094 7120 8146
rect 7040 7840 7120 8094
rect 520 7817 2120 7840
rect 520 7783 547 7817
rect 581 7783 619 7817
rect 653 7783 691 7817
rect 725 7783 763 7817
rect 797 7783 835 7817
rect 869 7783 907 7817
rect 941 7783 979 7817
rect 1013 7783 1051 7817
rect 1085 7783 1123 7817
rect 1157 7783 1195 7817
rect 1229 7783 1267 7817
rect 1301 7783 1339 7817
rect 1373 7783 1411 7817
rect 1445 7783 1483 7817
rect 1517 7783 1555 7817
rect 1589 7783 1627 7817
rect 1661 7783 1699 7817
rect 1733 7783 1771 7817
rect 1805 7783 1843 7817
rect 1877 7783 1915 7817
rect 1949 7783 1987 7817
rect 2021 7783 2059 7817
rect 2093 7783 2120 7817
rect 520 7760 2120 7783
rect 2440 7817 4040 7840
rect 2440 7783 2467 7817
rect 2501 7783 2539 7817
rect 2573 7783 2611 7817
rect 2645 7783 2683 7817
rect 2717 7783 2755 7817
rect 2789 7783 2827 7817
rect 2861 7783 2899 7817
rect 2933 7783 2971 7817
rect 3005 7783 3043 7817
rect 3077 7783 3115 7817
rect 3149 7783 3187 7817
rect 3221 7783 3259 7817
rect 3293 7783 3331 7817
rect 3365 7783 3403 7817
rect 3437 7783 3475 7817
rect 3509 7783 3547 7817
rect 3581 7783 3619 7817
rect 3653 7783 3691 7817
rect 3725 7783 3763 7817
rect 3797 7783 3835 7817
rect 3869 7783 3907 7817
rect 3941 7783 3979 7817
rect 4013 7783 4040 7817
rect 2440 7760 4040 7783
rect 4360 7817 5960 7840
rect 4360 7783 4387 7817
rect 4421 7783 4459 7817
rect 4493 7783 4531 7817
rect 4565 7783 4603 7817
rect 4637 7783 4675 7817
rect 4709 7783 4747 7817
rect 4781 7783 4819 7817
rect 4853 7783 4891 7817
rect 4925 7783 4963 7817
rect 4997 7783 5035 7817
rect 5069 7783 5107 7817
rect 5141 7783 5179 7817
rect 5213 7783 5251 7817
rect 5285 7783 5323 7817
rect 5357 7783 5395 7817
rect 5429 7783 5467 7817
rect 5501 7783 5539 7817
rect 5573 7783 5611 7817
rect 5645 7783 5683 7817
rect 5717 7783 5755 7817
rect 5789 7783 5827 7817
rect 5861 7783 5899 7817
rect 5933 7783 5960 7817
rect 4360 7760 5960 7783
rect 6280 7817 7880 7840
rect 6280 7783 6307 7817
rect 6341 7783 6379 7817
rect 6413 7783 6451 7817
rect 6485 7783 6523 7817
rect 6557 7783 6595 7817
rect 6629 7783 6667 7817
rect 6701 7783 6739 7817
rect 6773 7783 6811 7817
rect 6845 7783 6883 7817
rect 6917 7783 6955 7817
rect 6989 7783 7027 7817
rect 7061 7783 7099 7817
rect 7133 7783 7171 7817
rect 7205 7783 7243 7817
rect 7277 7783 7315 7817
rect 7349 7783 7387 7817
rect 7421 7783 7459 7817
rect 7493 7783 7531 7817
rect 7565 7783 7603 7817
rect 7637 7783 7675 7817
rect 7709 7783 7747 7817
rect 7781 7783 7819 7817
rect 7853 7783 7880 7817
rect 6280 7760 7880 7783
rect 320 7678 400 7720
rect 320 7626 334 7678
rect 386 7626 400 7678
rect 320 7614 400 7626
rect 320 7562 334 7614
rect 386 7562 400 7614
rect 320 7520 400 7562
rect 2240 7673 2320 7720
rect 2240 7639 2263 7673
rect 2297 7639 2320 7673
rect 2240 7601 2320 7639
rect 2240 7567 2263 7601
rect 2297 7567 2320 7601
rect 2240 7520 2320 7567
rect 4160 7673 4240 7720
rect 4160 7639 4183 7673
rect 4217 7639 4240 7673
rect 4160 7601 4240 7639
rect 4160 7567 4183 7601
rect 4217 7567 4240 7601
rect 4160 7520 4240 7567
rect 6080 7673 6160 7720
rect 6080 7639 6103 7673
rect 6137 7639 6160 7673
rect 6080 7601 6160 7639
rect 6080 7567 6103 7601
rect 6137 7567 6160 7601
rect 6080 7520 6160 7567
rect 8000 7673 8080 8574
rect 8160 8466 8240 8480
rect 8160 8414 8174 8466
rect 8226 8414 8240 8466
rect 8160 8400 8240 8414
rect 8160 8306 8240 8320
rect 8160 8254 8174 8306
rect 8226 8254 8240 8306
rect 8160 8240 8240 8254
rect 8000 7639 8023 7673
rect 8057 7639 8080 7673
rect 8000 7601 8080 7639
rect 8000 7567 8023 7601
rect 8057 7567 8080 7601
rect 8000 7520 8080 7567
rect 320 7078 400 7120
rect 320 7026 334 7078
rect 386 7026 400 7078
rect 320 7014 400 7026
rect 320 6962 334 7014
rect 386 6962 400 7014
rect 320 6920 400 6962
rect 2240 7073 2320 7120
rect 2240 7039 2263 7073
rect 2297 7039 2320 7073
rect 2240 7001 2320 7039
rect 2240 6967 2263 7001
rect 2297 6967 2320 7001
rect 2240 6920 2320 6967
rect 4160 7073 4240 7120
rect 4160 7039 4183 7073
rect 4217 7039 4240 7073
rect 4160 7001 4240 7039
rect 4160 6967 4183 7001
rect 4217 6967 4240 7001
rect 4160 6920 4240 6967
rect 6080 7073 6160 7120
rect 6080 7039 6103 7073
rect 6137 7039 6160 7073
rect 6080 7001 6160 7039
rect 6080 6967 6103 7001
rect 6137 6967 6160 7001
rect 6080 6920 6160 6967
rect 8000 7073 8080 7120
rect 8000 7039 8023 7073
rect 8057 7039 8080 7073
rect 8000 7001 8080 7039
rect 8000 6967 8023 7001
rect 8057 6967 8080 7001
rect 520 6857 2120 6880
rect 520 6823 547 6857
rect 581 6823 619 6857
rect 653 6823 691 6857
rect 725 6823 763 6857
rect 797 6823 835 6857
rect 869 6823 907 6857
rect 941 6823 979 6857
rect 1013 6823 1051 6857
rect 1085 6823 1123 6857
rect 1157 6823 1195 6857
rect 1229 6823 1267 6857
rect 1301 6823 1339 6857
rect 1373 6823 1411 6857
rect 1445 6823 1483 6857
rect 1517 6823 1555 6857
rect 1589 6823 1627 6857
rect 1661 6823 1699 6857
rect 1733 6823 1771 6857
rect 1805 6823 1843 6857
rect 1877 6823 1915 6857
rect 1949 6823 1987 6857
rect 2021 6823 2059 6857
rect 2093 6823 2120 6857
rect 520 6800 2120 6823
rect 2440 6857 4040 6880
rect 2440 6823 2467 6857
rect 2501 6823 2539 6857
rect 2573 6823 2611 6857
rect 2645 6823 2683 6857
rect 2717 6823 2755 6857
rect 2789 6823 2827 6857
rect 2861 6823 2899 6857
rect 2933 6823 2971 6857
rect 3005 6823 3043 6857
rect 3077 6823 3115 6857
rect 3149 6823 3187 6857
rect 3221 6823 3259 6857
rect 3293 6823 3331 6857
rect 3365 6823 3403 6857
rect 3437 6823 3475 6857
rect 3509 6823 3547 6857
rect 3581 6823 3619 6857
rect 3653 6823 3691 6857
rect 3725 6823 3763 6857
rect 3797 6823 3835 6857
rect 3869 6823 3907 6857
rect 3941 6823 3979 6857
rect 4013 6823 4040 6857
rect 2440 6800 4040 6823
rect 4360 6857 5960 6880
rect 4360 6823 4387 6857
rect 4421 6823 4459 6857
rect 4493 6823 4531 6857
rect 4565 6823 4603 6857
rect 4637 6823 4675 6857
rect 4709 6823 4747 6857
rect 4781 6823 4819 6857
rect 4853 6823 4891 6857
rect 4925 6823 4963 6857
rect 4997 6823 5035 6857
rect 5069 6823 5107 6857
rect 5141 6823 5179 6857
rect 5213 6823 5251 6857
rect 5285 6823 5323 6857
rect 5357 6823 5395 6857
rect 5429 6823 5467 6857
rect 5501 6823 5539 6857
rect 5573 6823 5611 6857
rect 5645 6823 5683 6857
rect 5717 6823 5755 6857
rect 5789 6823 5827 6857
rect 5861 6823 5899 6857
rect 5933 6823 5960 6857
rect 4360 6800 5960 6823
rect 6280 6857 7880 6880
rect 6280 6823 6307 6857
rect 6341 6823 6379 6857
rect 6413 6823 6451 6857
rect 6485 6823 6523 6857
rect 6557 6823 6595 6857
rect 6629 6823 6667 6857
rect 6701 6823 6739 6857
rect 6773 6823 6811 6857
rect 6845 6823 6883 6857
rect 6917 6823 6955 6857
rect 6989 6823 7027 6857
rect 7061 6823 7099 6857
rect 7133 6823 7171 6857
rect 7205 6823 7243 6857
rect 7277 6823 7315 6857
rect 7349 6823 7387 6857
rect 7421 6823 7459 6857
rect 7493 6823 7531 6857
rect 7565 6823 7603 6857
rect 7637 6823 7675 6857
rect 7709 6823 7747 6857
rect 7781 6823 7819 6857
rect 7853 6823 7880 6857
rect 6280 6800 7880 6823
rect 1280 6546 1360 6800
rect 1280 6494 1294 6546
rect 1346 6494 1360 6546
rect 1280 6480 1360 6494
rect 3200 6546 3280 6800
rect 3200 6494 3214 6546
rect 3266 6494 3280 6546
rect 3200 6480 3280 6494
rect 5120 6546 5200 6800
rect 5120 6494 5134 6546
rect 5186 6494 5200 6546
rect 5120 6480 5200 6494
rect 7040 6546 7120 6800
rect 7040 6494 7054 6546
rect 7106 6494 7120 6546
rect 7040 6480 7120 6494
rect 160 6386 240 6400
rect 160 6334 174 6386
rect 226 6334 240 6386
rect 160 6320 240 6334
rect 160 6226 240 6240
rect 160 6174 174 6226
rect 226 6174 240 6226
rect 160 6160 240 6174
rect 8000 6066 8080 6967
rect 8160 6386 8240 6400
rect 8160 6334 8174 6386
rect 8226 6334 8240 6386
rect 8160 6320 8240 6334
rect 8160 6226 8240 6240
rect 8160 6174 8174 6226
rect 8226 6174 8240 6226
rect 8160 6160 8240 6174
rect 8000 6014 8014 6066
rect 8066 6014 8080 6066
rect 160 5906 240 5920
rect 160 5854 174 5906
rect 226 5854 240 5906
rect 160 5840 240 5854
rect 160 5746 240 5760
rect 160 5694 174 5746
rect 226 5694 240 5746
rect 160 5680 240 5694
rect 1280 5586 1360 5600
rect 1280 5534 1294 5586
rect 1346 5534 1360 5586
rect 1280 5120 1360 5534
rect 3200 5586 3280 5600
rect 3200 5534 3214 5586
rect 3266 5534 3280 5586
rect 3200 5120 3280 5534
rect 5120 5586 5200 5600
rect 5120 5534 5134 5586
rect 5186 5534 5200 5586
rect 5120 5120 5200 5534
rect 7040 5586 7120 5600
rect 7040 5534 7054 5586
rect 7106 5534 7120 5586
rect 7040 5120 7120 5534
rect 520 5097 2120 5120
rect 520 5063 547 5097
rect 581 5063 619 5097
rect 653 5063 691 5097
rect 725 5063 763 5097
rect 797 5063 835 5097
rect 869 5063 907 5097
rect 941 5063 979 5097
rect 1013 5063 1051 5097
rect 1085 5063 1123 5097
rect 1157 5063 1195 5097
rect 1229 5063 1267 5097
rect 1301 5063 1339 5097
rect 1373 5063 1411 5097
rect 1445 5063 1483 5097
rect 1517 5063 1555 5097
rect 1589 5063 1627 5097
rect 1661 5063 1699 5097
rect 1733 5063 1771 5097
rect 1805 5063 1843 5097
rect 1877 5063 1915 5097
rect 1949 5063 1987 5097
rect 2021 5063 2059 5097
rect 2093 5063 2120 5097
rect 520 5040 2120 5063
rect 2440 5097 4040 5120
rect 2440 5063 2467 5097
rect 2501 5063 2539 5097
rect 2573 5063 2611 5097
rect 2645 5063 2683 5097
rect 2717 5063 2755 5097
rect 2789 5063 2827 5097
rect 2861 5063 2899 5097
rect 2933 5063 2971 5097
rect 3005 5063 3043 5097
rect 3077 5063 3115 5097
rect 3149 5063 3187 5097
rect 3221 5063 3259 5097
rect 3293 5063 3331 5097
rect 3365 5063 3403 5097
rect 3437 5063 3475 5097
rect 3509 5063 3547 5097
rect 3581 5063 3619 5097
rect 3653 5063 3691 5097
rect 3725 5063 3763 5097
rect 3797 5063 3835 5097
rect 3869 5063 3907 5097
rect 3941 5063 3979 5097
rect 4013 5063 4040 5097
rect 2440 5040 4040 5063
rect 4360 5097 5960 5120
rect 4360 5063 4387 5097
rect 4421 5063 4459 5097
rect 4493 5063 4531 5097
rect 4565 5063 4603 5097
rect 4637 5063 4675 5097
rect 4709 5063 4747 5097
rect 4781 5063 4819 5097
rect 4853 5063 4891 5097
rect 4925 5063 4963 5097
rect 4997 5063 5035 5097
rect 5069 5063 5107 5097
rect 5141 5063 5179 5097
rect 5213 5063 5251 5097
rect 5285 5063 5323 5097
rect 5357 5063 5395 5097
rect 5429 5063 5467 5097
rect 5501 5063 5539 5097
rect 5573 5063 5611 5097
rect 5645 5063 5683 5097
rect 5717 5063 5755 5097
rect 5789 5063 5827 5097
rect 5861 5063 5899 5097
rect 5933 5063 5960 5097
rect 4360 5040 5960 5063
rect 6280 5097 7880 5120
rect 6280 5063 6307 5097
rect 6341 5063 6379 5097
rect 6413 5063 6451 5097
rect 6485 5063 6523 5097
rect 6557 5063 6595 5097
rect 6629 5063 6667 5097
rect 6701 5063 6739 5097
rect 6773 5063 6811 5097
rect 6845 5063 6883 5097
rect 6917 5063 6955 5097
rect 6989 5063 7027 5097
rect 7061 5063 7099 5097
rect 7133 5063 7171 5097
rect 7205 5063 7243 5097
rect 7277 5063 7315 5097
rect 7349 5063 7387 5097
rect 7421 5063 7459 5097
rect 7493 5063 7531 5097
rect 7565 5063 7603 5097
rect 7637 5063 7675 5097
rect 7709 5063 7747 5097
rect 7781 5063 7819 5097
rect 7853 5063 7880 5097
rect 6280 5040 7880 5063
rect 320 4969 400 5000
rect 320 4935 343 4969
rect 377 4935 400 4969
rect 320 4897 400 4935
rect 320 4863 343 4897
rect 377 4863 400 4897
rect 320 4825 400 4863
rect 320 4791 343 4825
rect 377 4791 400 4825
rect 320 4754 400 4791
rect 320 4702 334 4754
rect 386 4702 400 4754
rect 320 4690 400 4702
rect 320 4638 334 4690
rect 386 4638 400 4690
rect 320 4626 400 4638
rect 320 4574 334 4626
rect 386 4574 400 4626
rect 320 4562 400 4574
rect 320 4510 334 4562
rect 386 4510 400 4562
rect 320 4503 343 4510
rect 377 4503 400 4510
rect 320 4498 400 4503
rect 320 4446 334 4498
rect 386 4446 400 4498
rect 320 4431 343 4446
rect 377 4431 400 4446
rect 320 4400 400 4431
rect 2240 4969 2320 5000
rect 2240 4935 2263 4969
rect 2297 4935 2320 4969
rect 2240 4897 2320 4935
rect 2240 4863 2263 4897
rect 2297 4863 2320 4897
rect 2240 4825 2320 4863
rect 2240 4791 2263 4825
rect 2297 4791 2320 4825
rect 2240 4753 2320 4791
rect 2240 4719 2263 4753
rect 2297 4719 2320 4753
rect 2240 4681 2320 4719
rect 2240 4647 2263 4681
rect 2297 4647 2320 4681
rect 2240 4609 2320 4647
rect 2240 4575 2263 4609
rect 2297 4575 2320 4609
rect 2240 4537 2320 4575
rect 2240 4503 2263 4537
rect 2297 4503 2320 4537
rect 2240 4465 2320 4503
rect 2240 4431 2263 4465
rect 2297 4431 2320 4465
rect 2240 4400 2320 4431
rect 4160 4969 4240 5000
rect 4160 4935 4183 4969
rect 4217 4935 4240 4969
rect 4160 4897 4240 4935
rect 4160 4863 4183 4897
rect 4217 4863 4240 4897
rect 4160 4825 4240 4863
rect 4160 4791 4183 4825
rect 4217 4791 4240 4825
rect 4160 4753 4240 4791
rect 4160 4719 4183 4753
rect 4217 4719 4240 4753
rect 4160 4681 4240 4719
rect 4160 4647 4183 4681
rect 4217 4647 4240 4681
rect 4160 4609 4240 4647
rect 4160 4575 4183 4609
rect 4217 4575 4240 4609
rect 4160 4537 4240 4575
rect 4160 4503 4183 4537
rect 4217 4503 4240 4537
rect 4160 4465 4240 4503
rect 4160 4431 4183 4465
rect 4217 4431 4240 4465
rect 4160 4400 4240 4431
rect 6080 4969 6160 5000
rect 6080 4935 6103 4969
rect 6137 4935 6160 4969
rect 6080 4897 6160 4935
rect 6080 4863 6103 4897
rect 6137 4863 6160 4897
rect 6080 4825 6160 4863
rect 6080 4791 6103 4825
rect 6137 4791 6160 4825
rect 6080 4753 6160 4791
rect 6080 4719 6103 4753
rect 6137 4719 6160 4753
rect 6080 4681 6160 4719
rect 6080 4647 6103 4681
rect 6137 4647 6160 4681
rect 6080 4609 6160 4647
rect 6080 4575 6103 4609
rect 6137 4575 6160 4609
rect 6080 4537 6160 4575
rect 6080 4503 6103 4537
rect 6137 4503 6160 4537
rect 6080 4465 6160 4503
rect 6080 4431 6103 4465
rect 6137 4431 6160 4465
rect 6080 4400 6160 4431
rect 8000 4969 8080 6014
rect 8160 5906 8240 5920
rect 8160 5854 8174 5906
rect 8226 5854 8240 5906
rect 8160 5840 8240 5854
rect 8160 5746 8240 5760
rect 8160 5694 8174 5746
rect 8226 5694 8240 5746
rect 8160 5680 8240 5694
rect 8000 4935 8023 4969
rect 8057 4935 8080 4969
rect 8000 4897 8080 4935
rect 8000 4863 8023 4897
rect 8057 4863 8080 4897
rect 8000 4825 8080 4863
rect 8000 4791 8023 4825
rect 8057 4791 8080 4825
rect 8000 4753 8080 4791
rect 8000 4719 8023 4753
rect 8057 4719 8080 4753
rect 8000 4681 8080 4719
rect 8000 4647 8023 4681
rect 8057 4647 8080 4681
rect 8000 4609 8080 4647
rect 8000 4575 8023 4609
rect 8057 4575 8080 4609
rect 8000 4537 8080 4575
rect 8000 4503 8023 4537
rect 8057 4503 8080 4537
rect 8000 4465 8080 4503
rect 8000 4431 8023 4465
rect 8057 4431 8080 4465
rect 8000 4400 8080 4431
rect 320 3649 400 3680
rect 320 3615 343 3649
rect 377 3615 400 3649
rect 320 3577 400 3615
rect 320 3543 343 3577
rect 377 3543 400 3577
rect 320 3505 400 3543
rect 320 3471 343 3505
rect 377 3471 400 3505
rect 320 3433 400 3471
rect 320 3399 343 3433
rect 377 3399 400 3433
rect 320 3361 400 3399
rect 320 3327 343 3361
rect 377 3327 400 3361
rect 320 3289 400 3327
rect 320 3255 343 3289
rect 377 3255 400 3289
rect 320 3217 400 3255
rect 320 3183 343 3217
rect 377 3183 400 3217
rect 320 3145 400 3183
rect 320 3111 343 3145
rect 377 3111 400 3145
rect 0 2786 80 2800
rect 0 2734 14 2786
rect 66 2734 80 2786
rect 0 2466 80 2734
rect 0 2414 14 2466
rect 66 2414 80 2466
rect 0 2400 80 2414
rect 160 2786 240 2800
rect 160 2734 174 2786
rect 226 2734 240 2786
rect 160 2466 240 2734
rect 160 2414 174 2466
rect 226 2414 240 2466
rect 160 2400 240 2414
rect 320 2786 400 3111
rect 2240 3649 2320 3680
rect 2240 3615 2263 3649
rect 2297 3615 2320 3649
rect 2240 3577 2320 3615
rect 2240 3543 2263 3577
rect 2297 3543 2320 3577
rect 2240 3505 2320 3543
rect 2240 3471 2263 3505
rect 2297 3471 2320 3505
rect 2240 3433 2320 3471
rect 2240 3399 2263 3433
rect 2297 3399 2320 3433
rect 2240 3361 2320 3399
rect 2240 3327 2263 3361
rect 2297 3327 2320 3361
rect 2240 3289 2320 3327
rect 2240 3255 2263 3289
rect 2297 3255 2320 3289
rect 2240 3217 2320 3255
rect 2240 3183 2263 3217
rect 2297 3183 2320 3217
rect 2240 3145 2320 3183
rect 2240 3111 2263 3145
rect 2297 3111 2320 3145
rect 2240 3080 2320 3111
rect 4160 3649 4240 3680
rect 4160 3615 4183 3649
rect 4217 3615 4240 3649
rect 4160 3577 4240 3615
rect 4160 3543 4183 3577
rect 4217 3543 4240 3577
rect 4160 3505 4240 3543
rect 4160 3471 4183 3505
rect 4217 3471 4240 3505
rect 4160 3433 4240 3471
rect 4160 3399 4183 3433
rect 4217 3399 4240 3433
rect 4160 3361 4240 3399
rect 4160 3327 4183 3361
rect 4217 3327 4240 3361
rect 4160 3289 4240 3327
rect 4160 3255 4183 3289
rect 4217 3255 4240 3289
rect 4160 3217 4240 3255
rect 4160 3183 4183 3217
rect 4217 3183 4240 3217
rect 4160 3145 4240 3183
rect 4160 3111 4183 3145
rect 4217 3111 4240 3145
rect 4160 3080 4240 3111
rect 6080 3649 6160 3680
rect 6080 3615 6103 3649
rect 6137 3615 6160 3649
rect 6080 3577 6160 3615
rect 6080 3543 6103 3577
rect 6137 3543 6160 3577
rect 6080 3505 6160 3543
rect 6080 3471 6103 3505
rect 6137 3471 6160 3505
rect 6080 3433 6160 3471
rect 6080 3399 6103 3433
rect 6137 3399 6160 3433
rect 6080 3361 6160 3399
rect 6080 3327 6103 3361
rect 6137 3327 6160 3361
rect 6080 3289 6160 3327
rect 6080 3255 6103 3289
rect 6137 3255 6160 3289
rect 6080 3217 6160 3255
rect 6080 3183 6103 3217
rect 6137 3183 6160 3217
rect 6080 3145 6160 3183
rect 6080 3111 6103 3145
rect 6137 3111 6160 3145
rect 6080 3080 6160 3111
rect 8000 3649 8080 3680
rect 8000 3634 8023 3649
rect 8057 3634 8080 3649
rect 8000 3582 8014 3634
rect 8066 3582 8080 3634
rect 8000 3577 8080 3582
rect 8000 3570 8023 3577
rect 8057 3570 8080 3577
rect 8000 3518 8014 3570
rect 8066 3518 8080 3570
rect 8000 3506 8080 3518
rect 8000 3454 8014 3506
rect 8066 3454 8080 3506
rect 8000 3442 8080 3454
rect 8000 3390 8014 3442
rect 8066 3390 8080 3442
rect 8000 3378 8080 3390
rect 8000 3326 8014 3378
rect 8066 3326 8080 3378
rect 8000 3289 8080 3326
rect 8000 3255 8023 3289
rect 8057 3255 8080 3289
rect 8000 3217 8080 3255
rect 8000 3183 8023 3217
rect 8057 3183 8080 3217
rect 8000 3145 8080 3183
rect 8000 3111 8023 3145
rect 8057 3111 8080 3145
rect 8000 3080 8080 3111
rect 520 3017 2120 3040
rect 520 2983 547 3017
rect 581 2983 619 3017
rect 653 2983 691 3017
rect 725 2983 763 3017
rect 797 2983 835 3017
rect 869 2983 907 3017
rect 941 2983 979 3017
rect 1013 2983 1051 3017
rect 1085 2983 1123 3017
rect 1157 2983 1195 3017
rect 1229 2983 1267 3017
rect 1301 2983 1339 3017
rect 1373 2983 1411 3017
rect 1445 2983 1483 3017
rect 1517 2983 1555 3017
rect 1589 2983 1627 3017
rect 1661 2983 1699 3017
rect 1733 2983 1771 3017
rect 1805 2983 1843 3017
rect 1877 2983 1915 3017
rect 1949 2983 1987 3017
rect 2021 2983 2059 3017
rect 2093 2983 2120 3017
rect 520 2960 2120 2983
rect 2440 3017 4040 3040
rect 2440 2983 2467 3017
rect 2501 2983 2539 3017
rect 2573 2983 2611 3017
rect 2645 2983 2683 3017
rect 2717 2983 2755 3017
rect 2789 2983 2827 3017
rect 2861 2983 2899 3017
rect 2933 2983 2971 3017
rect 3005 2983 3043 3017
rect 3077 2983 3115 3017
rect 3149 2983 3187 3017
rect 3221 2983 3259 3017
rect 3293 2983 3331 3017
rect 3365 2983 3403 3017
rect 3437 2983 3475 3017
rect 3509 2983 3547 3017
rect 3581 2983 3619 3017
rect 3653 2983 3691 3017
rect 3725 2983 3763 3017
rect 3797 2983 3835 3017
rect 3869 2983 3907 3017
rect 3941 2983 3979 3017
rect 4013 2983 4040 3017
rect 2440 2960 4040 2983
rect 4360 3017 5960 3040
rect 4360 2983 4387 3017
rect 4421 2983 4459 3017
rect 4493 2983 4531 3017
rect 4565 2983 4603 3017
rect 4637 2983 4675 3017
rect 4709 2983 4747 3017
rect 4781 2983 4819 3017
rect 4853 2983 4891 3017
rect 4925 2983 4963 3017
rect 4997 2983 5035 3017
rect 5069 2983 5107 3017
rect 5141 2983 5179 3017
rect 5213 2983 5251 3017
rect 5285 2983 5323 3017
rect 5357 2983 5395 3017
rect 5429 2983 5467 3017
rect 5501 2983 5539 3017
rect 5573 2983 5611 3017
rect 5645 2983 5683 3017
rect 5717 2983 5755 3017
rect 5789 2983 5827 3017
rect 5861 2983 5899 3017
rect 5933 2983 5960 3017
rect 4360 2960 5960 2983
rect 6280 3017 7880 3040
rect 6280 2983 6307 3017
rect 6341 2983 6379 3017
rect 6413 2983 6451 3017
rect 6485 2983 6523 3017
rect 6557 2983 6595 3017
rect 6629 2983 6667 3017
rect 6701 2983 6739 3017
rect 6773 2983 6811 3017
rect 6845 2983 6883 3017
rect 6917 2983 6955 3017
rect 6989 2983 7027 3017
rect 7061 2983 7099 3017
rect 7133 2983 7171 3017
rect 7205 2983 7243 3017
rect 7277 2983 7315 3017
rect 7349 2983 7387 3017
rect 7421 2983 7459 3017
rect 7493 2983 7531 3017
rect 7565 2983 7603 3017
rect 7637 2983 7675 3017
rect 7709 2983 7747 3017
rect 7781 2983 7819 3017
rect 7853 2983 7880 3017
rect 6280 2960 7880 2983
rect 320 2734 334 2786
rect 386 2734 400 2786
rect 320 2466 400 2734
rect 320 2414 334 2466
rect 386 2414 400 2466
rect 320 2209 400 2414
rect 480 2786 560 2800
rect 480 2734 494 2786
rect 546 2734 560 2786
rect 480 2466 560 2734
rect 480 2414 494 2466
rect 546 2414 560 2466
rect 480 2400 560 2414
rect 640 2786 720 2800
rect 640 2734 654 2786
rect 706 2734 720 2786
rect 640 2466 720 2734
rect 640 2414 654 2466
rect 706 2414 720 2466
rect 640 2400 720 2414
rect 800 2786 880 2800
rect 800 2734 814 2786
rect 866 2734 880 2786
rect 800 2466 880 2734
rect 800 2414 814 2466
rect 866 2414 880 2466
rect 800 2400 880 2414
rect 960 2786 1040 2800
rect 960 2734 974 2786
rect 1026 2734 1040 2786
rect 960 2466 1040 2734
rect 960 2414 974 2466
rect 1026 2414 1040 2466
rect 960 2400 1040 2414
rect 1120 2786 1200 2800
rect 1120 2734 1134 2786
rect 1186 2734 1200 2786
rect 1120 2466 1200 2734
rect 1280 2626 1360 2960
rect 1280 2574 1294 2626
rect 1346 2574 1360 2626
rect 1280 2560 1360 2574
rect 1440 2786 1520 2800
rect 1440 2734 1454 2786
rect 1506 2734 1520 2786
rect 1120 2414 1134 2466
rect 1186 2414 1200 2466
rect 1120 2400 1200 2414
rect 1440 2466 1520 2734
rect 1440 2414 1454 2466
rect 1506 2414 1520 2466
rect 1440 2400 1520 2414
rect 1600 2786 1680 2800
rect 1600 2734 1614 2786
rect 1666 2734 1680 2786
rect 1600 2466 1680 2734
rect 1600 2414 1614 2466
rect 1666 2414 1680 2466
rect 1600 2400 1680 2414
rect 1760 2786 1840 2800
rect 1760 2734 1774 2786
rect 1826 2734 1840 2786
rect 1760 2466 1840 2734
rect 1760 2414 1774 2466
rect 1826 2414 1840 2466
rect 1760 2400 1840 2414
rect 1920 2786 2000 2800
rect 1920 2734 1934 2786
rect 1986 2734 2000 2786
rect 1920 2466 2000 2734
rect 1920 2414 1934 2466
rect 1986 2414 2000 2466
rect 1920 2400 2000 2414
rect 2080 2786 2160 2800
rect 2080 2734 2094 2786
rect 2146 2734 2160 2786
rect 2080 2466 2160 2734
rect 2080 2414 2094 2466
rect 2146 2414 2160 2466
rect 2080 2400 2160 2414
rect 2240 2786 2320 2800
rect 2240 2734 2254 2786
rect 2306 2734 2320 2786
rect 2240 2466 2320 2734
rect 2240 2414 2254 2466
rect 2306 2414 2320 2466
rect 2240 2400 2320 2414
rect 2400 2786 2480 2800
rect 2400 2734 2414 2786
rect 2466 2734 2480 2786
rect 2400 2466 2480 2734
rect 2400 2414 2414 2466
rect 2466 2414 2480 2466
rect 2400 2400 2480 2414
rect 2560 2786 2640 2800
rect 2560 2734 2574 2786
rect 2626 2734 2640 2786
rect 2560 2466 2640 2734
rect 2560 2414 2574 2466
rect 2626 2414 2640 2466
rect 2560 2400 2640 2414
rect 2720 2786 2800 2800
rect 2720 2734 2734 2786
rect 2786 2734 2800 2786
rect 2720 2466 2800 2734
rect 2720 2414 2734 2466
rect 2786 2414 2800 2466
rect 2720 2400 2800 2414
rect 2880 2786 2960 2800
rect 2880 2734 2894 2786
rect 2946 2734 2960 2786
rect 2880 2466 2960 2734
rect 2880 2414 2894 2466
rect 2946 2414 2960 2466
rect 2880 2400 2960 2414
rect 3040 2786 3120 2800
rect 3040 2734 3054 2786
rect 3106 2734 3120 2786
rect 3040 2466 3120 2734
rect 3200 2626 3280 2960
rect 3200 2574 3214 2626
rect 3266 2574 3280 2626
rect 3200 2560 3280 2574
rect 3360 2786 3440 2800
rect 3360 2734 3374 2786
rect 3426 2734 3440 2786
rect 3040 2414 3054 2466
rect 3106 2414 3120 2466
rect 3040 2400 3120 2414
rect 3360 2466 3440 2734
rect 3360 2414 3374 2466
rect 3426 2414 3440 2466
rect 3360 2400 3440 2414
rect 3520 2786 3600 2800
rect 3520 2734 3534 2786
rect 3586 2734 3600 2786
rect 3520 2466 3600 2734
rect 3520 2414 3534 2466
rect 3586 2414 3600 2466
rect 3520 2400 3600 2414
rect 3680 2786 3760 2800
rect 3680 2734 3694 2786
rect 3746 2734 3760 2786
rect 3680 2466 3760 2734
rect 3680 2414 3694 2466
rect 3746 2414 3760 2466
rect 3680 2400 3760 2414
rect 3840 2786 3920 2800
rect 3840 2734 3854 2786
rect 3906 2734 3920 2786
rect 3840 2466 3920 2734
rect 3840 2414 3854 2466
rect 3906 2414 3920 2466
rect 3840 2400 3920 2414
rect 4000 2786 4080 2800
rect 4000 2734 4014 2786
rect 4066 2734 4080 2786
rect 4000 2466 4080 2734
rect 4000 2414 4014 2466
rect 4066 2414 4080 2466
rect 4000 2400 4080 2414
rect 4160 2786 4240 2800
rect 4160 2734 4174 2786
rect 4226 2734 4240 2786
rect 4160 2466 4240 2734
rect 4160 2414 4174 2466
rect 4226 2414 4240 2466
rect 4160 2400 4240 2414
rect 4320 2786 4400 2800
rect 4320 2734 4334 2786
rect 4386 2734 4400 2786
rect 4320 2466 4400 2734
rect 4320 2414 4334 2466
rect 4386 2414 4400 2466
rect 4320 2400 4400 2414
rect 4480 2786 4560 2800
rect 4480 2734 4494 2786
rect 4546 2734 4560 2786
rect 4480 2466 4560 2734
rect 4480 2414 4494 2466
rect 4546 2414 4560 2466
rect 4480 2400 4560 2414
rect 4640 2786 4720 2800
rect 4640 2734 4654 2786
rect 4706 2734 4720 2786
rect 4640 2466 4720 2734
rect 4640 2414 4654 2466
rect 4706 2414 4720 2466
rect 4640 2400 4720 2414
rect 4800 2786 4880 2800
rect 4800 2734 4814 2786
rect 4866 2734 4880 2786
rect 4800 2466 4880 2734
rect 4800 2414 4814 2466
rect 4866 2414 4880 2466
rect 4800 2400 4880 2414
rect 4960 2786 5040 2800
rect 4960 2734 4974 2786
rect 5026 2734 5040 2786
rect 4960 2466 5040 2734
rect 5120 2626 5200 2960
rect 5120 2574 5134 2626
rect 5186 2574 5200 2626
rect 5120 2560 5200 2574
rect 5280 2786 5360 2800
rect 5280 2734 5294 2786
rect 5346 2734 5360 2786
rect 4960 2414 4974 2466
rect 5026 2414 5040 2466
rect 4960 2400 5040 2414
rect 5280 2466 5360 2734
rect 5280 2414 5294 2466
rect 5346 2414 5360 2466
rect 5280 2400 5360 2414
rect 5440 2786 5520 2800
rect 5440 2734 5454 2786
rect 5506 2734 5520 2786
rect 5440 2466 5520 2734
rect 5440 2414 5454 2466
rect 5506 2414 5520 2466
rect 5440 2400 5520 2414
rect 5600 2786 5680 2800
rect 5600 2734 5614 2786
rect 5666 2734 5680 2786
rect 5600 2466 5680 2734
rect 5600 2414 5614 2466
rect 5666 2414 5680 2466
rect 5600 2400 5680 2414
rect 5760 2786 5840 2800
rect 5760 2734 5774 2786
rect 5826 2734 5840 2786
rect 5760 2466 5840 2734
rect 5760 2414 5774 2466
rect 5826 2414 5840 2466
rect 5760 2400 5840 2414
rect 5920 2786 6000 2800
rect 5920 2734 5934 2786
rect 5986 2734 6000 2786
rect 5920 2466 6000 2734
rect 5920 2414 5934 2466
rect 5986 2414 6000 2466
rect 5920 2400 6000 2414
rect 6080 2786 6160 2800
rect 6080 2734 6094 2786
rect 6146 2734 6160 2786
rect 6080 2466 6160 2734
rect 6080 2414 6094 2466
rect 6146 2414 6160 2466
rect 6080 2400 6160 2414
rect 6240 2786 6320 2800
rect 6240 2734 6254 2786
rect 6306 2734 6320 2786
rect 6240 2466 6320 2734
rect 6240 2414 6254 2466
rect 6306 2414 6320 2466
rect 6240 2400 6320 2414
rect 6400 2786 6480 2800
rect 6400 2734 6414 2786
rect 6466 2734 6480 2786
rect 6400 2466 6480 2734
rect 6400 2414 6414 2466
rect 6466 2414 6480 2466
rect 6400 2400 6480 2414
rect 6560 2786 6640 2800
rect 6560 2734 6574 2786
rect 6626 2734 6640 2786
rect 6560 2466 6640 2734
rect 6560 2414 6574 2466
rect 6626 2414 6640 2466
rect 6560 2400 6640 2414
rect 6720 2786 6800 2800
rect 6720 2734 6734 2786
rect 6786 2734 6800 2786
rect 6720 2466 6800 2734
rect 6720 2414 6734 2466
rect 6786 2414 6800 2466
rect 6720 2400 6800 2414
rect 6880 2786 6960 2800
rect 6880 2734 6894 2786
rect 6946 2734 6960 2786
rect 6880 2466 6960 2734
rect 7040 2626 7120 2960
rect 7040 2574 7054 2626
rect 7106 2574 7120 2626
rect 7040 2560 7120 2574
rect 7200 2786 7280 2800
rect 7200 2734 7214 2786
rect 7266 2734 7280 2786
rect 6880 2414 6894 2466
rect 6946 2414 6960 2466
rect 6880 2400 6960 2414
rect 7200 2466 7280 2734
rect 7200 2414 7214 2466
rect 7266 2414 7280 2466
rect 7200 2400 7280 2414
rect 7360 2786 7440 2800
rect 7360 2734 7374 2786
rect 7426 2734 7440 2786
rect 7360 2466 7440 2734
rect 7360 2414 7374 2466
rect 7426 2414 7440 2466
rect 7360 2400 7440 2414
rect 7520 2786 7600 2800
rect 7520 2734 7534 2786
rect 7586 2734 7600 2786
rect 7520 2466 7600 2734
rect 7520 2414 7534 2466
rect 7586 2414 7600 2466
rect 7520 2400 7600 2414
rect 7680 2786 7760 2800
rect 7680 2734 7694 2786
rect 7746 2734 7760 2786
rect 7680 2466 7760 2734
rect 7680 2414 7694 2466
rect 7746 2414 7760 2466
rect 7680 2400 7760 2414
rect 7840 2786 7920 2800
rect 7840 2734 7854 2786
rect 7906 2734 7920 2786
rect 7840 2466 7920 2734
rect 7840 2414 7854 2466
rect 7906 2414 7920 2466
rect 7840 2400 7920 2414
rect 8000 2786 8080 2800
rect 8000 2734 8014 2786
rect 8066 2734 8080 2786
rect 8000 2466 8080 2734
rect 8000 2414 8014 2466
rect 8066 2414 8080 2466
rect 8000 2400 8080 2414
rect 8160 2786 8240 2800
rect 8160 2734 8174 2786
rect 8226 2734 8240 2786
rect 8160 2466 8240 2734
rect 8160 2414 8174 2466
rect 8226 2414 8240 2466
rect 8160 2400 8240 2414
rect 8320 2786 8400 2800
rect 8320 2734 8334 2786
rect 8386 2734 8400 2786
rect 8320 2466 8400 2734
rect 8320 2414 8334 2466
rect 8386 2414 8400 2466
rect 8320 2400 8400 2414
rect 320 2175 343 2209
rect 377 2175 400 2209
rect 320 2137 400 2175
rect 320 2103 343 2137
rect 377 2103 400 2137
rect 320 2065 400 2103
rect 320 2031 343 2065
rect 377 2031 400 2065
rect 320 1993 400 2031
rect 320 1959 343 1993
rect 377 1959 400 1993
rect 320 1921 400 1959
rect 320 1887 343 1921
rect 377 1887 400 1921
rect 320 1849 400 1887
rect 320 1815 343 1849
rect 377 1815 400 1849
rect 320 1777 400 1815
rect 320 1743 343 1777
rect 377 1743 400 1777
rect 320 1705 400 1743
rect 320 1671 343 1705
rect 377 1671 400 1705
rect 320 1640 400 1671
rect 2240 2209 2320 2240
rect 2240 2175 2263 2209
rect 2297 2175 2320 2209
rect 2240 2137 2320 2175
rect 2240 2103 2263 2137
rect 2297 2103 2320 2137
rect 2240 2065 2320 2103
rect 2240 2031 2263 2065
rect 2297 2031 2320 2065
rect 2240 1993 2320 2031
rect 2240 1959 2263 1993
rect 2297 1959 2320 1993
rect 2240 1921 2320 1959
rect 2240 1887 2263 1921
rect 2297 1887 2320 1921
rect 2240 1849 2320 1887
rect 2240 1815 2263 1849
rect 2297 1815 2320 1849
rect 2240 1777 2320 1815
rect 2240 1743 2263 1777
rect 2297 1743 2320 1777
rect 2240 1705 2320 1743
rect 2240 1671 2263 1705
rect 2297 1671 2320 1705
rect 2240 1640 2320 1671
rect 4160 2209 4240 2240
rect 4160 2175 4183 2209
rect 4217 2175 4240 2209
rect 4160 2137 4240 2175
rect 4160 2103 4183 2137
rect 4217 2103 4240 2137
rect 4160 2065 4240 2103
rect 4160 2031 4183 2065
rect 4217 2031 4240 2065
rect 4160 1993 4240 2031
rect 4160 1959 4183 1993
rect 4217 1959 4240 1993
rect 4160 1921 4240 1959
rect 4160 1887 4183 1921
rect 4217 1887 4240 1921
rect 4160 1849 4240 1887
rect 4160 1815 4183 1849
rect 4217 1815 4240 1849
rect 4160 1777 4240 1815
rect 4160 1743 4183 1777
rect 4217 1743 4240 1777
rect 4160 1705 4240 1743
rect 4160 1671 4183 1705
rect 4217 1671 4240 1705
rect 4160 1640 4240 1671
rect 6080 2209 6160 2240
rect 6080 2175 6103 2209
rect 6137 2175 6160 2209
rect 6080 2137 6160 2175
rect 6080 2103 6103 2137
rect 6137 2103 6160 2137
rect 6080 2065 6160 2103
rect 6080 2031 6103 2065
rect 6137 2031 6160 2065
rect 6080 1993 6160 2031
rect 6080 1959 6103 1993
rect 6137 1959 6160 1993
rect 6080 1921 6160 1959
rect 6080 1887 6103 1921
rect 6137 1887 6160 1921
rect 6080 1849 6160 1887
rect 6080 1815 6103 1849
rect 6137 1815 6160 1849
rect 6080 1777 6160 1815
rect 6080 1743 6103 1777
rect 6137 1743 6160 1777
rect 6080 1705 6160 1743
rect 6080 1671 6103 1705
rect 6137 1671 6160 1705
rect 6080 1640 6160 1671
rect 8000 2209 8080 2240
rect 8000 2175 8023 2209
rect 8057 2175 8080 2209
rect 8000 2137 8080 2175
rect 8000 2103 8023 2137
rect 8057 2103 8080 2137
rect 8000 2065 8080 2103
rect 8000 2031 8023 2065
rect 8057 2031 8080 2065
rect 8000 1993 8080 2031
rect 8000 1959 8023 1993
rect 8057 1959 8080 1993
rect 8000 1921 8080 1959
rect 8000 1887 8023 1921
rect 8057 1887 8080 1921
rect 8000 1849 8080 1887
rect 8000 1815 8023 1849
rect 8057 1815 8080 1849
rect 8000 1777 8080 1815
rect 8000 1743 8023 1777
rect 8057 1743 8080 1777
rect 8000 1705 8080 1743
rect 8000 1671 8023 1705
rect 8057 1671 8080 1705
rect 520 1577 2120 1600
rect 520 1543 547 1577
rect 581 1543 619 1577
rect 653 1543 691 1577
rect 725 1543 763 1577
rect 797 1543 835 1577
rect 869 1543 907 1577
rect 941 1543 979 1577
rect 1013 1543 1051 1577
rect 1085 1543 1123 1577
rect 1157 1543 1195 1577
rect 1229 1543 1267 1577
rect 1301 1543 1339 1577
rect 1373 1543 1411 1577
rect 1445 1543 1483 1577
rect 1517 1543 1555 1577
rect 1589 1543 1627 1577
rect 1661 1543 1699 1577
rect 1733 1543 1771 1577
rect 1805 1543 1843 1577
rect 1877 1543 1915 1577
rect 1949 1543 1987 1577
rect 2021 1543 2059 1577
rect 2093 1543 2120 1577
rect 520 1520 2120 1543
rect 2440 1577 4040 1600
rect 2440 1543 2467 1577
rect 2501 1543 2539 1577
rect 2573 1543 2611 1577
rect 2645 1543 2683 1577
rect 2717 1543 2755 1577
rect 2789 1543 2827 1577
rect 2861 1543 2899 1577
rect 2933 1543 2971 1577
rect 3005 1543 3043 1577
rect 3077 1543 3115 1577
rect 3149 1543 3187 1577
rect 3221 1543 3259 1577
rect 3293 1543 3331 1577
rect 3365 1543 3403 1577
rect 3437 1543 3475 1577
rect 3509 1543 3547 1577
rect 3581 1543 3619 1577
rect 3653 1543 3691 1577
rect 3725 1543 3763 1577
rect 3797 1543 3835 1577
rect 3869 1543 3907 1577
rect 3941 1543 3979 1577
rect 4013 1543 4040 1577
rect 2440 1520 4040 1543
rect 4360 1577 5960 1600
rect 4360 1543 4387 1577
rect 4421 1543 4459 1577
rect 4493 1543 4531 1577
rect 4565 1543 4603 1577
rect 4637 1543 4675 1577
rect 4709 1543 4747 1577
rect 4781 1543 4819 1577
rect 4853 1543 4891 1577
rect 4925 1543 4963 1577
rect 4997 1543 5035 1577
rect 5069 1543 5107 1577
rect 5141 1543 5179 1577
rect 5213 1543 5251 1577
rect 5285 1543 5323 1577
rect 5357 1543 5395 1577
rect 5429 1543 5467 1577
rect 5501 1543 5539 1577
rect 5573 1543 5611 1577
rect 5645 1543 5683 1577
rect 5717 1543 5755 1577
rect 5789 1543 5827 1577
rect 5861 1543 5899 1577
rect 5933 1543 5960 1577
rect 4360 1520 5960 1543
rect 6280 1577 7880 1600
rect 6280 1543 6307 1577
rect 6341 1543 6379 1577
rect 6413 1543 6451 1577
rect 6485 1543 6523 1577
rect 6557 1543 6595 1577
rect 6629 1543 6667 1577
rect 6701 1543 6739 1577
rect 6773 1543 6811 1577
rect 6845 1543 6883 1577
rect 6917 1543 6955 1577
rect 6989 1543 7027 1577
rect 7061 1543 7099 1577
rect 7133 1543 7171 1577
rect 7205 1543 7243 1577
rect 7277 1543 7315 1577
rect 7349 1543 7387 1577
rect 7421 1543 7459 1577
rect 7493 1543 7531 1577
rect 7565 1543 7603 1577
rect 7637 1543 7675 1577
rect 7709 1543 7747 1577
rect 7781 1543 7819 1577
rect 7853 1543 7880 1577
rect 6280 1520 7880 1543
rect 1280 1106 1360 1520
rect 1280 1054 1294 1106
rect 1346 1054 1360 1106
rect 160 946 240 960
rect 160 894 174 946
rect 226 894 240 946
rect 160 880 240 894
rect 320 937 400 960
rect 320 903 343 937
rect 377 903 400 937
rect 320 880 400 903
rect 480 937 560 960
rect 480 903 503 937
rect 537 903 560 937
rect 480 880 560 903
rect 640 937 720 960
rect 640 903 663 937
rect 697 903 720 937
rect 640 880 720 903
rect 800 937 880 960
rect 800 903 823 937
rect 857 903 880 937
rect 800 880 880 903
rect 960 937 1040 960
rect 960 903 983 937
rect 1017 903 1040 937
rect 960 880 1040 903
rect 1120 937 1200 960
rect 1120 903 1143 937
rect 1177 903 1200 937
rect 1120 880 1200 903
rect 1280 480 1360 1054
rect 3200 1106 3280 1520
rect 3200 1054 3214 1106
rect 3266 1054 3280 1106
rect 1440 937 1520 960
rect 1440 903 1463 937
rect 1497 903 1520 937
rect 1440 880 1520 903
rect 1600 937 1680 960
rect 1600 903 1623 937
rect 1657 903 1680 937
rect 1600 880 1680 903
rect 1760 937 1840 960
rect 1760 903 1783 937
rect 1817 903 1840 937
rect 1760 880 1840 903
rect 1920 937 2000 960
rect 1920 903 1943 937
rect 1977 903 2000 937
rect 1920 880 2000 903
rect 2080 937 2160 960
rect 2080 903 2103 937
rect 2137 903 2160 937
rect 2080 880 2160 903
rect 2240 937 2320 960
rect 2240 903 2263 937
rect 2297 903 2320 937
rect 2240 880 2320 903
rect 2400 937 2480 960
rect 2400 903 2423 937
rect 2457 903 2480 937
rect 2400 880 2480 903
rect 2560 937 2640 960
rect 2560 903 2583 937
rect 2617 903 2640 937
rect 2560 880 2640 903
rect 2720 937 2800 960
rect 2720 903 2743 937
rect 2777 903 2800 937
rect 2720 880 2800 903
rect 2880 937 2960 960
rect 2880 903 2903 937
rect 2937 903 2960 937
rect 2880 880 2960 903
rect 3040 937 3120 960
rect 3040 903 3063 937
rect 3097 903 3120 937
rect 3040 880 3120 903
rect 3200 480 3280 1054
rect 5120 1106 5200 1520
rect 5120 1054 5134 1106
rect 5186 1054 5200 1106
rect 3360 937 3440 960
rect 3360 903 3383 937
rect 3417 903 3440 937
rect 3360 880 3440 903
rect 3520 937 3600 960
rect 3520 903 3543 937
rect 3577 903 3600 937
rect 3520 880 3600 903
rect 3680 937 3760 960
rect 3680 903 3703 937
rect 3737 903 3760 937
rect 3680 880 3760 903
rect 3840 937 3920 960
rect 3840 903 3863 937
rect 3897 903 3920 937
rect 3840 880 3920 903
rect 4000 937 4080 960
rect 4000 903 4023 937
rect 4057 903 4080 937
rect 4000 880 4080 903
rect 4160 937 4240 960
rect 4160 903 4183 937
rect 4217 903 4240 937
rect 4160 880 4240 903
rect 4320 937 4400 960
rect 4320 903 4343 937
rect 4377 903 4400 937
rect 4320 880 4400 903
rect 4480 937 4560 960
rect 4480 903 4503 937
rect 4537 903 4560 937
rect 4480 880 4560 903
rect 4640 937 4720 960
rect 4640 903 4663 937
rect 4697 903 4720 937
rect 4640 880 4720 903
rect 4800 937 4880 960
rect 4800 903 4823 937
rect 4857 903 4880 937
rect 4800 880 4880 903
rect 4960 937 5040 960
rect 4960 903 4983 937
rect 5017 903 5040 937
rect 4960 880 5040 903
rect 5120 480 5200 1054
rect 7040 1106 7120 1520
rect 7040 1054 7054 1106
rect 7106 1054 7120 1106
rect 5280 937 5360 960
rect 5280 903 5303 937
rect 5337 903 5360 937
rect 5280 880 5360 903
rect 5440 937 5520 960
rect 5440 903 5463 937
rect 5497 903 5520 937
rect 5440 880 5520 903
rect 5600 937 5680 960
rect 5600 903 5623 937
rect 5657 903 5680 937
rect 5600 880 5680 903
rect 5760 937 5840 960
rect 5760 903 5783 937
rect 5817 903 5840 937
rect 5760 880 5840 903
rect 5920 937 6000 960
rect 5920 903 5943 937
rect 5977 903 6000 937
rect 5920 880 6000 903
rect 6080 937 6160 960
rect 6080 903 6103 937
rect 6137 903 6160 937
rect 6080 880 6160 903
rect 6240 937 6320 960
rect 6240 903 6263 937
rect 6297 903 6320 937
rect 6240 880 6320 903
rect 6400 937 6480 960
rect 6400 903 6423 937
rect 6457 903 6480 937
rect 6400 880 6480 903
rect 6560 937 6640 960
rect 6560 903 6583 937
rect 6617 903 6640 937
rect 6560 880 6640 903
rect 6720 937 6800 960
rect 6720 903 6743 937
rect 6777 903 6800 937
rect 6720 880 6800 903
rect 6880 937 6960 960
rect 6880 903 6903 937
rect 6937 903 6960 937
rect 6880 880 6960 903
rect 7040 480 7120 1054
rect 8000 1106 8080 1671
rect 8000 1054 8014 1106
rect 8066 1054 8080 1106
rect 7200 937 7280 960
rect 7200 903 7223 937
rect 7257 903 7280 937
rect 7200 880 7280 903
rect 7360 937 7440 960
rect 7360 903 7383 937
rect 7417 903 7440 937
rect 7360 880 7440 903
rect 7520 937 7600 960
rect 7520 903 7543 937
rect 7577 903 7600 937
rect 7520 880 7600 903
rect 7680 937 7760 960
rect 7680 903 7703 937
rect 7737 903 7760 937
rect 7680 880 7760 903
rect 7840 937 7920 960
rect 7840 903 7863 937
rect 7897 903 7920 937
rect 7840 880 7920 903
rect 8000 786 8080 1054
rect 8160 937 8240 960
rect 8160 903 8183 937
rect 8217 903 8240 937
rect 8160 880 8240 903
rect 8000 734 8014 786
rect 8066 734 8080 786
rect 520 457 2120 480
rect 520 423 547 457
rect 581 423 619 457
rect 653 423 691 457
rect 725 423 763 457
rect 797 423 835 457
rect 869 423 907 457
rect 941 423 979 457
rect 1013 423 1051 457
rect 1085 423 1123 457
rect 1157 423 1195 457
rect 1229 423 1267 457
rect 1301 423 1339 457
rect 1373 423 1411 457
rect 1445 423 1483 457
rect 1517 423 1555 457
rect 1589 423 1627 457
rect 1661 423 1699 457
rect 1733 423 1771 457
rect 1805 423 1843 457
rect 1877 423 1915 457
rect 1949 423 1987 457
rect 2021 423 2059 457
rect 2093 423 2120 457
rect 520 400 2120 423
rect 2440 457 4040 480
rect 2440 423 2467 457
rect 2501 423 2539 457
rect 2573 423 2611 457
rect 2645 423 2683 457
rect 2717 423 2755 457
rect 2789 423 2827 457
rect 2861 423 2899 457
rect 2933 423 2971 457
rect 3005 423 3043 457
rect 3077 423 3115 457
rect 3149 423 3187 457
rect 3221 423 3259 457
rect 3293 423 3331 457
rect 3365 423 3403 457
rect 3437 423 3475 457
rect 3509 423 3547 457
rect 3581 423 3619 457
rect 3653 423 3691 457
rect 3725 423 3763 457
rect 3797 423 3835 457
rect 3869 423 3907 457
rect 3941 423 3979 457
rect 4013 423 4040 457
rect 2440 400 4040 423
rect 4360 457 5960 480
rect 4360 423 4387 457
rect 4421 423 4459 457
rect 4493 423 4531 457
rect 4565 423 4603 457
rect 4637 423 4675 457
rect 4709 423 4747 457
rect 4781 423 4819 457
rect 4853 423 4891 457
rect 4925 423 4963 457
rect 4997 423 5035 457
rect 5069 423 5107 457
rect 5141 423 5179 457
rect 5213 423 5251 457
rect 5285 423 5323 457
rect 5357 423 5395 457
rect 5429 423 5467 457
rect 5501 423 5539 457
rect 5573 423 5611 457
rect 5645 423 5683 457
rect 5717 423 5755 457
rect 5789 423 5827 457
rect 5861 423 5899 457
rect 5933 423 5960 457
rect 4360 400 5960 423
rect 6280 457 7880 480
rect 6280 423 6307 457
rect 6341 423 6379 457
rect 6413 423 6451 457
rect 6485 423 6523 457
rect 6557 423 6595 457
rect 6629 423 6667 457
rect 6701 423 6739 457
rect 6773 423 6811 457
rect 6845 423 6883 457
rect 6917 423 6955 457
rect 6989 423 7027 457
rect 7061 423 7099 457
rect 7133 423 7171 457
rect 7205 423 7243 457
rect 7277 423 7315 457
rect 7349 423 7387 457
rect 7421 423 7459 457
rect 7493 423 7531 457
rect 7565 423 7603 457
rect 7637 423 7675 457
rect 7709 423 7747 457
rect 7781 423 7819 457
rect 7853 423 7880 457
rect 6280 400 7880 423
rect 320 318 400 360
rect 320 266 334 318
rect 386 266 400 318
rect 320 254 400 266
rect 320 202 334 254
rect 386 202 400 254
rect 320 160 400 202
rect 2240 313 2320 360
rect 2240 279 2263 313
rect 2297 279 2320 313
rect 2240 241 2320 279
rect 2240 207 2263 241
rect 2297 207 2320 241
rect 2240 160 2320 207
rect 4160 313 4240 360
rect 4160 279 4183 313
rect 4217 279 4240 313
rect 4160 241 4240 279
rect 4160 207 4183 241
rect 4217 207 4240 241
rect 4160 160 4240 207
rect 6080 313 6160 360
rect 6080 279 6103 313
rect 6137 279 6160 313
rect 6080 241 6160 279
rect 6080 207 6103 241
rect 6137 207 6160 241
rect 6080 160 6160 207
rect 8000 313 8080 734
rect 8000 279 8023 313
rect 8057 279 8080 313
rect 8000 241 8080 279
rect 8000 207 8023 241
rect 8057 207 8080 241
rect 8000 160 8080 207
rect 160 -94 240 -80
rect 160 -146 174 -94
rect 226 -146 240 -94
rect 160 -160 240 -146
rect 320 -94 400 -80
rect 320 -146 334 -94
rect 386 -146 400 -94
rect 320 -160 400 -146
rect 480 -94 560 -80
rect 480 -146 494 -94
rect 546 -146 560 -94
rect 480 -160 560 -146
rect 640 -94 720 -80
rect 640 -146 654 -94
rect 706 -146 720 -94
rect 640 -160 720 -146
rect 800 -94 880 -80
rect 800 -146 814 -94
rect 866 -146 880 -94
rect 800 -160 880 -146
rect 960 -94 1040 -80
rect 960 -146 974 -94
rect 1026 -146 1040 -94
rect 960 -160 1040 -146
rect 1120 -94 1200 -80
rect 1120 -146 1134 -94
rect 1186 -146 1200 -94
rect 1120 -160 1200 -146
rect 1440 -94 1520 -80
rect 1440 -146 1454 -94
rect 1506 -146 1520 -94
rect 1440 -160 1520 -146
rect 1600 -94 1680 -80
rect 1600 -146 1614 -94
rect 1666 -146 1680 -94
rect 1600 -160 1680 -146
rect 1760 -94 1840 -80
rect 1760 -146 1774 -94
rect 1826 -146 1840 -94
rect 1760 -160 1840 -146
rect 1920 -94 2000 -80
rect 1920 -146 1934 -94
rect 1986 -146 2000 -94
rect 1920 -160 2000 -146
rect 2080 -94 2160 -80
rect 2080 -146 2094 -94
rect 2146 -146 2160 -94
rect 2080 -160 2160 -146
rect 2240 -94 2320 -80
rect 2240 -146 2254 -94
rect 2306 -146 2320 -94
rect 2240 -160 2320 -146
rect 2400 -94 2480 -80
rect 2400 -146 2414 -94
rect 2466 -146 2480 -94
rect 2400 -160 2480 -146
rect 2560 -94 2640 -80
rect 2560 -146 2574 -94
rect 2626 -146 2640 -94
rect 2560 -160 2640 -146
rect 2720 -94 2800 -80
rect 2720 -146 2734 -94
rect 2786 -146 2800 -94
rect 2720 -160 2800 -146
rect 2880 -94 2960 -80
rect 2880 -146 2894 -94
rect 2946 -146 2960 -94
rect 2880 -160 2960 -146
rect 3040 -94 3120 -80
rect 3040 -146 3054 -94
rect 3106 -146 3120 -94
rect 3040 -160 3120 -146
rect 3360 -94 3440 -80
rect 3360 -146 3374 -94
rect 3426 -146 3440 -94
rect 3360 -160 3440 -146
rect 3520 -94 3600 -80
rect 3520 -146 3534 -94
rect 3586 -146 3600 -94
rect 3520 -160 3600 -146
rect 3680 -94 3760 -80
rect 3680 -146 3694 -94
rect 3746 -146 3760 -94
rect 3680 -160 3760 -146
rect 3840 -94 3920 -80
rect 3840 -146 3854 -94
rect 3906 -146 3920 -94
rect 3840 -160 3920 -146
rect 4000 -94 4080 -80
rect 4000 -146 4014 -94
rect 4066 -146 4080 -94
rect 4000 -160 4080 -146
rect 4160 -94 4240 -80
rect 4160 -146 4174 -94
rect 4226 -146 4240 -94
rect 4160 -160 4240 -146
rect 4320 -94 4400 -80
rect 4320 -146 4334 -94
rect 4386 -146 4400 -94
rect 4320 -160 4400 -146
rect 4480 -94 4560 -80
rect 4480 -146 4494 -94
rect 4546 -146 4560 -94
rect 4480 -160 4560 -146
rect 4640 -94 4720 -80
rect 4640 -146 4654 -94
rect 4706 -146 4720 -94
rect 4640 -160 4720 -146
rect 4800 -94 4880 -80
rect 4800 -146 4814 -94
rect 4866 -146 4880 -94
rect 4800 -160 4880 -146
rect 4960 -94 5040 -80
rect 4960 -146 4974 -94
rect 5026 -146 5040 -94
rect 4960 -160 5040 -146
rect 5280 -94 5360 -80
rect 5280 -146 5294 -94
rect 5346 -146 5360 -94
rect 5280 -160 5360 -146
rect 5440 -94 5520 -80
rect 5440 -146 5454 -94
rect 5506 -146 5520 -94
rect 5440 -160 5520 -146
rect 5600 -94 5680 -80
rect 5600 -146 5614 -94
rect 5666 -146 5680 -94
rect 5600 -160 5680 -146
rect 5760 -94 5840 -80
rect 5760 -146 5774 -94
rect 5826 -146 5840 -94
rect 5760 -160 5840 -146
rect 5920 -94 6000 -80
rect 5920 -146 5934 -94
rect 5986 -146 6000 -94
rect 5920 -160 6000 -146
rect 6080 -94 6160 -80
rect 6080 -146 6094 -94
rect 6146 -146 6160 -94
rect 6080 -160 6160 -146
rect 6240 -94 6320 -80
rect 6240 -146 6254 -94
rect 6306 -146 6320 -94
rect 6240 -160 6320 -146
rect 6400 -94 6480 -80
rect 6400 -146 6414 -94
rect 6466 -146 6480 -94
rect 6400 -160 6480 -146
rect 6560 -94 6640 -80
rect 6560 -146 6574 -94
rect 6626 -146 6640 -94
rect 6560 -160 6640 -146
rect 6720 -94 6800 -80
rect 6720 -146 6734 -94
rect 6786 -146 6800 -94
rect 6720 -160 6800 -146
rect 6880 -94 6960 -80
rect 6880 -146 6894 -94
rect 6946 -146 6960 -94
rect 6880 -160 6960 -146
rect 7200 -94 7280 -80
rect 7200 -146 7214 -94
rect 7266 -146 7280 -94
rect 7200 -160 7280 -146
rect 7360 -94 7440 -80
rect 7360 -146 7374 -94
rect 7426 -146 7440 -94
rect 7360 -160 7440 -146
rect 7520 -94 7600 -80
rect 7520 -146 7534 -94
rect 7586 -146 7600 -94
rect 7520 -160 7600 -146
rect 7680 -94 7760 -80
rect 7680 -146 7694 -94
rect 7746 -146 7760 -94
rect 7680 -160 7760 -146
rect 7840 -94 7920 -80
rect 7840 -146 7854 -94
rect 7906 -146 7920 -94
rect 7840 -160 7920 -146
rect 8160 -94 8240 -80
rect 8160 -146 8174 -94
rect 8226 -146 8240 -94
rect 8160 -160 8240 -146
rect 1280 -254 1360 -240
rect 1280 -306 1294 -254
rect 1346 -306 1360 -254
rect 1280 -560 1360 -306
rect 3200 -254 3280 -240
rect 3200 -306 3214 -254
rect 3266 -306 3280 -254
rect 3200 -560 3280 -306
rect 5120 -254 5200 -240
rect 5120 -306 5134 -254
rect 5186 -306 5200 -254
rect 5120 -560 5200 -306
rect 7040 -254 7120 -240
rect 7040 -306 7054 -254
rect 7106 -306 7120 -254
rect 7040 -560 7120 -306
rect 8000 -254 8080 -240
rect 8000 -306 8014 -254
rect 8066 -306 8080 -254
rect 520 -583 2120 -560
rect 520 -617 547 -583
rect 581 -617 619 -583
rect 653 -617 691 -583
rect 725 -617 763 -583
rect 797 -617 835 -583
rect 869 -617 907 -583
rect 941 -617 979 -583
rect 1013 -617 1051 -583
rect 1085 -617 1123 -583
rect 1157 -617 1195 -583
rect 1229 -617 1267 -583
rect 1301 -617 1339 -583
rect 1373 -617 1411 -583
rect 1445 -617 1483 -583
rect 1517 -617 1555 -583
rect 1589 -617 1627 -583
rect 1661 -617 1699 -583
rect 1733 -617 1771 -583
rect 1805 -617 1843 -583
rect 1877 -617 1915 -583
rect 1949 -617 1987 -583
rect 2021 -617 2059 -583
rect 2093 -617 2120 -583
rect 520 -640 2120 -617
rect 2440 -583 4040 -560
rect 2440 -617 2467 -583
rect 2501 -617 2539 -583
rect 2573 -617 2611 -583
rect 2645 -617 2683 -583
rect 2717 -617 2755 -583
rect 2789 -617 2827 -583
rect 2861 -617 2899 -583
rect 2933 -617 2971 -583
rect 3005 -617 3043 -583
rect 3077 -617 3115 -583
rect 3149 -617 3187 -583
rect 3221 -617 3259 -583
rect 3293 -617 3331 -583
rect 3365 -617 3403 -583
rect 3437 -617 3475 -583
rect 3509 -617 3547 -583
rect 3581 -617 3619 -583
rect 3653 -617 3691 -583
rect 3725 -617 3763 -583
rect 3797 -617 3835 -583
rect 3869 -617 3907 -583
rect 3941 -617 3979 -583
rect 4013 -617 4040 -583
rect 2440 -640 4040 -617
rect 4360 -583 5960 -560
rect 4360 -617 4387 -583
rect 4421 -617 4459 -583
rect 4493 -617 4531 -583
rect 4565 -617 4603 -583
rect 4637 -617 4675 -583
rect 4709 -617 4747 -583
rect 4781 -617 4819 -583
rect 4853 -617 4891 -583
rect 4925 -617 4963 -583
rect 4997 -617 5035 -583
rect 5069 -617 5107 -583
rect 5141 -617 5179 -583
rect 5213 -617 5251 -583
rect 5285 -617 5323 -583
rect 5357 -617 5395 -583
rect 5429 -617 5467 -583
rect 5501 -617 5539 -583
rect 5573 -617 5611 -583
rect 5645 -617 5683 -583
rect 5717 -617 5755 -583
rect 5789 -617 5827 -583
rect 5861 -617 5899 -583
rect 5933 -617 5960 -583
rect 4360 -640 5960 -617
rect 6280 -583 7880 -560
rect 6280 -617 6307 -583
rect 6341 -617 6379 -583
rect 6413 -617 6451 -583
rect 6485 -617 6523 -583
rect 6557 -617 6595 -583
rect 6629 -617 6667 -583
rect 6701 -617 6739 -583
rect 6773 -617 6811 -583
rect 6845 -617 6883 -583
rect 6917 -617 6955 -583
rect 6989 -617 7027 -583
rect 7061 -617 7099 -583
rect 7133 -617 7171 -583
rect 7205 -617 7243 -583
rect 7277 -617 7315 -583
rect 7349 -617 7387 -583
rect 7421 -617 7459 -583
rect 7493 -617 7531 -583
rect 7565 -617 7603 -583
rect 7637 -617 7675 -583
rect 7709 -617 7747 -583
rect 7781 -617 7819 -583
rect 7853 -617 7880 -583
rect 6280 -640 7880 -617
rect 320 -722 400 -680
rect 320 -774 334 -722
rect 386 -774 400 -722
rect 320 -786 400 -774
rect 320 -838 334 -786
rect 386 -838 400 -786
rect 320 -880 400 -838
rect 2240 -727 2320 -680
rect 2240 -761 2263 -727
rect 2297 -761 2320 -727
rect 2240 -799 2320 -761
rect 2240 -833 2263 -799
rect 2297 -833 2320 -799
rect 2240 -880 2320 -833
rect 4160 -727 4240 -680
rect 4160 -761 4183 -727
rect 4217 -761 4240 -727
rect 4160 -799 4240 -761
rect 4160 -833 4183 -799
rect 4217 -833 4240 -799
rect 4160 -880 4240 -833
rect 6080 -727 6160 -680
rect 6080 -761 6103 -727
rect 6137 -761 6160 -727
rect 6080 -799 6160 -761
rect 6080 -833 6103 -799
rect 6137 -833 6160 -799
rect 6080 -880 6160 -833
rect 8000 -727 8080 -306
rect 8000 -761 8023 -727
rect 8057 -761 8080 -727
rect 8000 -799 8080 -761
rect 8000 -833 8023 -799
rect 8057 -833 8080 -799
rect 8000 -880 8080 -833
<< via1 >>
rect 334 9695 343 9714
rect 343 9695 377 9714
rect 377 9695 386 9714
rect 334 9662 386 9695
rect 334 9623 343 9650
rect 343 9623 377 9650
rect 377 9623 386 9650
rect 334 9598 386 9623
rect 334 9585 386 9586
rect 334 9551 343 9585
rect 343 9551 377 9585
rect 377 9551 386 9585
rect 334 9534 386 9551
rect 334 9513 386 9522
rect 334 9479 343 9513
rect 343 9479 377 9513
rect 377 9479 386 9513
rect 334 9470 386 9479
rect 334 9441 386 9458
rect 334 9407 343 9441
rect 343 9407 377 9441
rect 377 9407 386 9441
rect 334 9406 386 9407
rect 1294 8574 1346 8626
rect 3214 8574 3266 8626
rect 5134 8574 5186 8626
rect 7054 8574 7106 8626
rect 8014 8574 8066 8626
rect 174 8457 226 8466
rect 174 8423 183 8457
rect 183 8423 217 8457
rect 217 8423 226 8457
rect 174 8414 226 8423
rect 174 8297 226 8306
rect 174 8263 183 8297
rect 183 8263 217 8297
rect 217 8263 226 8297
rect 174 8254 226 8263
rect 1294 8094 1346 8146
rect 3214 8094 3266 8146
rect 5134 8094 5186 8146
rect 7054 8094 7106 8146
rect 334 7673 386 7678
rect 334 7639 343 7673
rect 343 7639 377 7673
rect 377 7639 386 7673
rect 334 7626 386 7639
rect 334 7601 386 7614
rect 334 7567 343 7601
rect 343 7567 377 7601
rect 377 7567 386 7601
rect 334 7562 386 7567
rect 8174 8457 8226 8466
rect 8174 8423 8183 8457
rect 8183 8423 8217 8457
rect 8217 8423 8226 8457
rect 8174 8414 8226 8423
rect 8174 8297 8226 8306
rect 8174 8263 8183 8297
rect 8183 8263 8217 8297
rect 8217 8263 8226 8297
rect 8174 8254 8226 8263
rect 334 7073 386 7078
rect 334 7039 343 7073
rect 343 7039 377 7073
rect 377 7039 386 7073
rect 334 7026 386 7039
rect 334 7001 386 7014
rect 334 6967 343 7001
rect 343 6967 377 7001
rect 377 6967 386 7001
rect 334 6962 386 6967
rect 1294 6494 1346 6546
rect 3214 6494 3266 6546
rect 5134 6494 5186 6546
rect 7054 6494 7106 6546
rect 174 6377 226 6386
rect 174 6343 183 6377
rect 183 6343 217 6377
rect 217 6343 226 6377
rect 174 6334 226 6343
rect 174 6217 226 6226
rect 174 6183 183 6217
rect 183 6183 217 6217
rect 217 6183 226 6217
rect 174 6174 226 6183
rect 8174 6377 8226 6386
rect 8174 6343 8183 6377
rect 8183 6343 8217 6377
rect 8217 6343 8226 6377
rect 8174 6334 8226 6343
rect 8174 6217 8226 6226
rect 8174 6183 8183 6217
rect 8183 6183 8217 6217
rect 8217 6183 8226 6217
rect 8174 6174 8226 6183
rect 8014 6014 8066 6066
rect 174 5897 226 5906
rect 174 5863 183 5897
rect 183 5863 217 5897
rect 217 5863 226 5897
rect 174 5854 226 5863
rect 174 5737 226 5746
rect 174 5703 183 5737
rect 183 5703 217 5737
rect 217 5703 226 5737
rect 174 5694 226 5703
rect 1294 5534 1346 5586
rect 3214 5534 3266 5586
rect 5134 5534 5186 5586
rect 7054 5534 7106 5586
rect 334 4753 386 4754
rect 334 4719 343 4753
rect 343 4719 377 4753
rect 377 4719 386 4753
rect 334 4702 386 4719
rect 334 4681 386 4690
rect 334 4647 343 4681
rect 343 4647 377 4681
rect 377 4647 386 4681
rect 334 4638 386 4647
rect 334 4609 386 4626
rect 334 4575 343 4609
rect 343 4575 377 4609
rect 377 4575 386 4609
rect 334 4574 386 4575
rect 334 4537 386 4562
rect 334 4510 343 4537
rect 343 4510 377 4537
rect 377 4510 386 4537
rect 334 4465 386 4498
rect 334 4446 343 4465
rect 343 4446 377 4465
rect 377 4446 386 4465
rect 8174 5897 8226 5906
rect 8174 5863 8183 5897
rect 8183 5863 8217 5897
rect 8217 5863 8226 5897
rect 8174 5854 8226 5863
rect 8174 5737 8226 5746
rect 8174 5703 8183 5737
rect 8183 5703 8217 5737
rect 8217 5703 8226 5737
rect 8174 5694 8226 5703
rect 14 2734 66 2786
rect 14 2414 66 2466
rect 174 2734 226 2786
rect 174 2414 226 2466
rect 8014 3615 8023 3634
rect 8023 3615 8057 3634
rect 8057 3615 8066 3634
rect 8014 3582 8066 3615
rect 8014 3543 8023 3570
rect 8023 3543 8057 3570
rect 8057 3543 8066 3570
rect 8014 3518 8066 3543
rect 8014 3505 8066 3506
rect 8014 3471 8023 3505
rect 8023 3471 8057 3505
rect 8057 3471 8066 3505
rect 8014 3454 8066 3471
rect 8014 3433 8066 3442
rect 8014 3399 8023 3433
rect 8023 3399 8057 3433
rect 8057 3399 8066 3433
rect 8014 3390 8066 3399
rect 8014 3361 8066 3378
rect 8014 3327 8023 3361
rect 8023 3327 8057 3361
rect 8057 3327 8066 3361
rect 8014 3326 8066 3327
rect 334 2734 386 2786
rect 334 2414 386 2466
rect 494 2734 546 2786
rect 494 2414 546 2466
rect 654 2734 706 2786
rect 654 2414 706 2466
rect 814 2734 866 2786
rect 814 2414 866 2466
rect 974 2734 1026 2786
rect 974 2414 1026 2466
rect 1134 2734 1186 2786
rect 1294 2574 1346 2626
rect 1454 2734 1506 2786
rect 1134 2414 1186 2466
rect 1454 2414 1506 2466
rect 1614 2734 1666 2786
rect 1614 2414 1666 2466
rect 1774 2734 1826 2786
rect 1774 2414 1826 2466
rect 1934 2734 1986 2786
rect 1934 2414 1986 2466
rect 2094 2734 2146 2786
rect 2094 2414 2146 2466
rect 2254 2734 2306 2786
rect 2254 2414 2306 2466
rect 2414 2734 2466 2786
rect 2414 2414 2466 2466
rect 2574 2734 2626 2786
rect 2574 2414 2626 2466
rect 2734 2734 2786 2786
rect 2734 2414 2786 2466
rect 2894 2734 2946 2786
rect 2894 2414 2946 2466
rect 3054 2734 3106 2786
rect 3214 2574 3266 2626
rect 3374 2734 3426 2786
rect 3054 2414 3106 2466
rect 3374 2414 3426 2466
rect 3534 2734 3586 2786
rect 3534 2414 3586 2466
rect 3694 2734 3746 2786
rect 3694 2414 3746 2466
rect 3854 2734 3906 2786
rect 3854 2414 3906 2466
rect 4014 2734 4066 2786
rect 4014 2414 4066 2466
rect 4174 2734 4226 2786
rect 4174 2414 4226 2466
rect 4334 2734 4386 2786
rect 4334 2414 4386 2466
rect 4494 2734 4546 2786
rect 4494 2414 4546 2466
rect 4654 2734 4706 2786
rect 4654 2414 4706 2466
rect 4814 2734 4866 2786
rect 4814 2414 4866 2466
rect 4974 2734 5026 2786
rect 5134 2574 5186 2626
rect 5294 2734 5346 2786
rect 4974 2414 5026 2466
rect 5294 2414 5346 2466
rect 5454 2734 5506 2786
rect 5454 2414 5506 2466
rect 5614 2734 5666 2786
rect 5614 2414 5666 2466
rect 5774 2734 5826 2786
rect 5774 2414 5826 2466
rect 5934 2734 5986 2786
rect 5934 2414 5986 2466
rect 6094 2734 6146 2786
rect 6094 2414 6146 2466
rect 6254 2734 6306 2786
rect 6254 2414 6306 2466
rect 6414 2734 6466 2786
rect 6414 2414 6466 2466
rect 6574 2734 6626 2786
rect 6574 2414 6626 2466
rect 6734 2734 6786 2786
rect 6734 2414 6786 2466
rect 6894 2734 6946 2786
rect 7054 2574 7106 2626
rect 7214 2734 7266 2786
rect 6894 2414 6946 2466
rect 7214 2414 7266 2466
rect 7374 2734 7426 2786
rect 7374 2414 7426 2466
rect 7534 2734 7586 2786
rect 7534 2414 7586 2466
rect 7694 2734 7746 2786
rect 7694 2414 7746 2466
rect 7854 2734 7906 2786
rect 7854 2414 7906 2466
rect 8014 2734 8066 2786
rect 8014 2414 8066 2466
rect 8174 2734 8226 2786
rect 8174 2414 8226 2466
rect 8334 2734 8386 2786
rect 8334 2414 8386 2466
rect 1294 1054 1346 1106
rect 174 937 226 946
rect 174 903 183 937
rect 183 903 217 937
rect 217 903 226 937
rect 174 894 226 903
rect 3214 1054 3266 1106
rect 5134 1054 5186 1106
rect 7054 1054 7106 1106
rect 8014 1054 8066 1106
rect 8014 734 8066 786
rect 334 313 386 318
rect 334 279 343 313
rect 343 279 377 313
rect 377 279 386 313
rect 334 266 386 279
rect 334 241 386 254
rect 334 207 343 241
rect 343 207 377 241
rect 377 207 386 241
rect 334 202 386 207
rect 174 -103 226 -94
rect 174 -137 183 -103
rect 183 -137 217 -103
rect 217 -137 226 -103
rect 174 -146 226 -137
rect 334 -103 386 -94
rect 334 -137 343 -103
rect 343 -137 377 -103
rect 377 -137 386 -103
rect 334 -146 386 -137
rect 494 -103 546 -94
rect 494 -137 503 -103
rect 503 -137 537 -103
rect 537 -137 546 -103
rect 494 -146 546 -137
rect 654 -103 706 -94
rect 654 -137 663 -103
rect 663 -137 697 -103
rect 697 -137 706 -103
rect 654 -146 706 -137
rect 814 -103 866 -94
rect 814 -137 823 -103
rect 823 -137 857 -103
rect 857 -137 866 -103
rect 814 -146 866 -137
rect 974 -103 1026 -94
rect 974 -137 983 -103
rect 983 -137 1017 -103
rect 1017 -137 1026 -103
rect 974 -146 1026 -137
rect 1134 -103 1186 -94
rect 1134 -137 1143 -103
rect 1143 -137 1177 -103
rect 1177 -137 1186 -103
rect 1134 -146 1186 -137
rect 1454 -103 1506 -94
rect 1454 -137 1463 -103
rect 1463 -137 1497 -103
rect 1497 -137 1506 -103
rect 1454 -146 1506 -137
rect 1614 -103 1666 -94
rect 1614 -137 1623 -103
rect 1623 -137 1657 -103
rect 1657 -137 1666 -103
rect 1614 -146 1666 -137
rect 1774 -103 1826 -94
rect 1774 -137 1783 -103
rect 1783 -137 1817 -103
rect 1817 -137 1826 -103
rect 1774 -146 1826 -137
rect 1934 -103 1986 -94
rect 1934 -137 1943 -103
rect 1943 -137 1977 -103
rect 1977 -137 1986 -103
rect 1934 -146 1986 -137
rect 2094 -103 2146 -94
rect 2094 -137 2103 -103
rect 2103 -137 2137 -103
rect 2137 -137 2146 -103
rect 2094 -146 2146 -137
rect 2254 -103 2306 -94
rect 2254 -137 2263 -103
rect 2263 -137 2297 -103
rect 2297 -137 2306 -103
rect 2254 -146 2306 -137
rect 2414 -103 2466 -94
rect 2414 -137 2423 -103
rect 2423 -137 2457 -103
rect 2457 -137 2466 -103
rect 2414 -146 2466 -137
rect 2574 -103 2626 -94
rect 2574 -137 2583 -103
rect 2583 -137 2617 -103
rect 2617 -137 2626 -103
rect 2574 -146 2626 -137
rect 2734 -103 2786 -94
rect 2734 -137 2743 -103
rect 2743 -137 2777 -103
rect 2777 -137 2786 -103
rect 2734 -146 2786 -137
rect 2894 -103 2946 -94
rect 2894 -137 2903 -103
rect 2903 -137 2937 -103
rect 2937 -137 2946 -103
rect 2894 -146 2946 -137
rect 3054 -103 3106 -94
rect 3054 -137 3063 -103
rect 3063 -137 3097 -103
rect 3097 -137 3106 -103
rect 3054 -146 3106 -137
rect 3374 -103 3426 -94
rect 3374 -137 3383 -103
rect 3383 -137 3417 -103
rect 3417 -137 3426 -103
rect 3374 -146 3426 -137
rect 3534 -103 3586 -94
rect 3534 -137 3543 -103
rect 3543 -137 3577 -103
rect 3577 -137 3586 -103
rect 3534 -146 3586 -137
rect 3694 -103 3746 -94
rect 3694 -137 3703 -103
rect 3703 -137 3737 -103
rect 3737 -137 3746 -103
rect 3694 -146 3746 -137
rect 3854 -103 3906 -94
rect 3854 -137 3863 -103
rect 3863 -137 3897 -103
rect 3897 -137 3906 -103
rect 3854 -146 3906 -137
rect 4014 -103 4066 -94
rect 4014 -137 4023 -103
rect 4023 -137 4057 -103
rect 4057 -137 4066 -103
rect 4014 -146 4066 -137
rect 4174 -103 4226 -94
rect 4174 -137 4183 -103
rect 4183 -137 4217 -103
rect 4217 -137 4226 -103
rect 4174 -146 4226 -137
rect 4334 -103 4386 -94
rect 4334 -137 4343 -103
rect 4343 -137 4377 -103
rect 4377 -137 4386 -103
rect 4334 -146 4386 -137
rect 4494 -103 4546 -94
rect 4494 -137 4503 -103
rect 4503 -137 4537 -103
rect 4537 -137 4546 -103
rect 4494 -146 4546 -137
rect 4654 -103 4706 -94
rect 4654 -137 4663 -103
rect 4663 -137 4697 -103
rect 4697 -137 4706 -103
rect 4654 -146 4706 -137
rect 4814 -103 4866 -94
rect 4814 -137 4823 -103
rect 4823 -137 4857 -103
rect 4857 -137 4866 -103
rect 4814 -146 4866 -137
rect 4974 -103 5026 -94
rect 4974 -137 4983 -103
rect 4983 -137 5017 -103
rect 5017 -137 5026 -103
rect 4974 -146 5026 -137
rect 5294 -103 5346 -94
rect 5294 -137 5303 -103
rect 5303 -137 5337 -103
rect 5337 -137 5346 -103
rect 5294 -146 5346 -137
rect 5454 -103 5506 -94
rect 5454 -137 5463 -103
rect 5463 -137 5497 -103
rect 5497 -137 5506 -103
rect 5454 -146 5506 -137
rect 5614 -103 5666 -94
rect 5614 -137 5623 -103
rect 5623 -137 5657 -103
rect 5657 -137 5666 -103
rect 5614 -146 5666 -137
rect 5774 -103 5826 -94
rect 5774 -137 5783 -103
rect 5783 -137 5817 -103
rect 5817 -137 5826 -103
rect 5774 -146 5826 -137
rect 5934 -103 5986 -94
rect 5934 -137 5943 -103
rect 5943 -137 5977 -103
rect 5977 -137 5986 -103
rect 5934 -146 5986 -137
rect 6094 -103 6146 -94
rect 6094 -137 6103 -103
rect 6103 -137 6137 -103
rect 6137 -137 6146 -103
rect 6094 -146 6146 -137
rect 6254 -103 6306 -94
rect 6254 -137 6263 -103
rect 6263 -137 6297 -103
rect 6297 -137 6306 -103
rect 6254 -146 6306 -137
rect 6414 -103 6466 -94
rect 6414 -137 6423 -103
rect 6423 -137 6457 -103
rect 6457 -137 6466 -103
rect 6414 -146 6466 -137
rect 6574 -103 6626 -94
rect 6574 -137 6583 -103
rect 6583 -137 6617 -103
rect 6617 -137 6626 -103
rect 6574 -146 6626 -137
rect 6734 -103 6786 -94
rect 6734 -137 6743 -103
rect 6743 -137 6777 -103
rect 6777 -137 6786 -103
rect 6734 -146 6786 -137
rect 6894 -103 6946 -94
rect 6894 -137 6903 -103
rect 6903 -137 6937 -103
rect 6937 -137 6946 -103
rect 6894 -146 6946 -137
rect 7214 -103 7266 -94
rect 7214 -137 7223 -103
rect 7223 -137 7257 -103
rect 7257 -137 7266 -103
rect 7214 -146 7266 -137
rect 7374 -103 7426 -94
rect 7374 -137 7383 -103
rect 7383 -137 7417 -103
rect 7417 -137 7426 -103
rect 7374 -146 7426 -137
rect 7534 -103 7586 -94
rect 7534 -137 7543 -103
rect 7543 -137 7577 -103
rect 7577 -137 7586 -103
rect 7534 -146 7586 -137
rect 7694 -103 7746 -94
rect 7694 -137 7703 -103
rect 7703 -137 7737 -103
rect 7737 -137 7746 -103
rect 7694 -146 7746 -137
rect 7854 -103 7906 -94
rect 7854 -137 7863 -103
rect 7863 -137 7897 -103
rect 7897 -137 7906 -103
rect 7854 -146 7906 -137
rect 8174 -103 8226 -94
rect 8174 -137 8183 -103
rect 8183 -137 8217 -103
rect 8217 -137 8226 -103
rect 8174 -146 8226 -137
rect 1294 -306 1346 -254
rect 3214 -306 3266 -254
rect 5134 -306 5186 -254
rect 7054 -306 7106 -254
rect 8014 -306 8066 -254
rect 334 -727 386 -722
rect 334 -761 343 -727
rect 343 -761 377 -727
rect 377 -761 386 -727
rect 334 -774 386 -761
rect 334 -799 386 -786
rect 334 -833 343 -799
rect 343 -833 377 -799
rect 377 -833 386 -799
rect 334 -838 386 -833
<< metal2 >>
rect 320 9714 400 9760
rect 320 9708 334 9714
rect 386 9708 400 9714
rect 320 9652 332 9708
rect 388 9652 400 9708
rect 320 9650 400 9652
rect 320 9628 334 9650
rect 386 9628 400 9650
rect 320 9572 332 9628
rect 388 9572 400 9628
rect 320 9548 334 9572
rect 386 9548 400 9572
rect 320 9492 332 9548
rect 388 9492 400 9548
rect 320 9470 334 9492
rect 386 9470 400 9492
rect 320 9468 400 9470
rect 320 9412 332 9468
rect 388 9412 400 9468
rect 320 9406 334 9412
rect 386 9406 400 9412
rect 320 9360 400 9406
rect 0 8788 8400 8800
rect 0 8732 172 8788
rect 228 8732 332 8788
rect 388 8732 492 8788
rect 548 8732 652 8788
rect 708 8732 812 8788
rect 868 8732 972 8788
rect 1028 8732 1132 8788
rect 1188 8732 1452 8788
rect 1508 8732 1612 8788
rect 1668 8732 1772 8788
rect 1828 8732 1932 8788
rect 1988 8732 2092 8788
rect 2148 8732 2252 8788
rect 2308 8732 2412 8788
rect 2468 8732 2572 8788
rect 2628 8732 2732 8788
rect 2788 8732 2892 8788
rect 2948 8732 3052 8788
rect 3108 8732 3372 8788
rect 3428 8732 3532 8788
rect 3588 8732 3692 8788
rect 3748 8732 3852 8788
rect 3908 8732 4012 8788
rect 4068 8732 4172 8788
rect 4228 8732 4332 8788
rect 4388 8732 4492 8788
rect 4548 8732 4652 8788
rect 4708 8732 4812 8788
rect 4868 8732 4972 8788
rect 5028 8732 5292 8788
rect 5348 8732 5452 8788
rect 5508 8732 5612 8788
rect 5668 8732 5772 8788
rect 5828 8732 5932 8788
rect 5988 8732 6092 8788
rect 6148 8732 6252 8788
rect 6308 8732 6412 8788
rect 6468 8732 6572 8788
rect 6628 8732 6732 8788
rect 6788 8732 6892 8788
rect 6948 8732 7212 8788
rect 7268 8732 7372 8788
rect 7428 8732 7532 8788
rect 7588 8732 7692 8788
rect 7748 8732 7852 8788
rect 7908 8732 8012 8788
rect 8068 8732 8172 8788
rect 8228 8732 8400 8788
rect 0 8720 8400 8732
rect 0 8626 8400 8640
rect 0 8574 1294 8626
rect 1346 8574 3214 8626
rect 3266 8574 5134 8626
rect 5186 8574 7054 8626
rect 7106 8574 8014 8626
rect 8066 8574 8400 8626
rect 0 8560 8400 8574
rect 0 8468 8400 8480
rect 0 8412 172 8468
rect 228 8412 332 8468
rect 388 8412 492 8468
rect 548 8412 652 8468
rect 708 8412 812 8468
rect 868 8412 972 8468
rect 1028 8412 1132 8468
rect 1188 8412 1452 8468
rect 1508 8412 1612 8468
rect 1668 8412 1772 8468
rect 1828 8412 1932 8468
rect 1988 8412 2092 8468
rect 2148 8412 2252 8468
rect 2308 8412 2412 8468
rect 2468 8412 2572 8468
rect 2628 8412 2732 8468
rect 2788 8412 2892 8468
rect 2948 8412 3052 8468
rect 3108 8412 3372 8468
rect 3428 8412 3532 8468
rect 3588 8412 3692 8468
rect 3748 8412 3852 8468
rect 3908 8412 4012 8468
rect 4068 8412 4172 8468
rect 4228 8412 4332 8468
rect 4388 8412 4492 8468
rect 4548 8412 4652 8468
rect 4708 8412 4812 8468
rect 4868 8412 4972 8468
rect 5028 8412 5292 8468
rect 5348 8412 5452 8468
rect 5508 8412 5612 8468
rect 5668 8412 5772 8468
rect 5828 8412 5932 8468
rect 5988 8412 6092 8468
rect 6148 8412 6252 8468
rect 6308 8412 6412 8468
rect 6468 8412 6572 8468
rect 6628 8412 6732 8468
rect 6788 8412 6892 8468
rect 6948 8412 7212 8468
rect 7268 8412 7372 8468
rect 7428 8412 7532 8468
rect 7588 8412 7692 8468
rect 7748 8412 7852 8468
rect 7908 8412 8012 8468
rect 8068 8412 8172 8468
rect 8228 8412 8400 8468
rect 0 8400 8400 8412
rect 0 8308 8400 8320
rect 0 8252 172 8308
rect 228 8252 332 8308
rect 388 8252 492 8308
rect 548 8252 652 8308
rect 708 8252 812 8308
rect 868 8252 972 8308
rect 1028 8252 1132 8308
rect 1188 8252 1452 8308
rect 1508 8252 1612 8308
rect 1668 8252 1772 8308
rect 1828 8252 1932 8308
rect 1988 8252 2092 8308
rect 2148 8252 2252 8308
rect 2308 8252 2412 8308
rect 2468 8252 2572 8308
rect 2628 8252 2732 8308
rect 2788 8252 2892 8308
rect 2948 8252 3052 8308
rect 3108 8252 3372 8308
rect 3428 8252 3532 8308
rect 3588 8252 3692 8308
rect 3748 8252 3852 8308
rect 3908 8252 4012 8308
rect 4068 8252 4172 8308
rect 4228 8252 4332 8308
rect 4388 8252 4492 8308
rect 4548 8252 4652 8308
rect 4708 8252 4812 8308
rect 4868 8252 4972 8308
rect 5028 8252 5292 8308
rect 5348 8252 5452 8308
rect 5508 8252 5612 8308
rect 5668 8252 5772 8308
rect 5828 8252 5932 8308
rect 5988 8252 6092 8308
rect 6148 8252 6252 8308
rect 6308 8252 6412 8308
rect 6468 8252 6572 8308
rect 6628 8252 6732 8308
rect 6788 8252 6892 8308
rect 6948 8252 7212 8308
rect 7268 8252 7372 8308
rect 7428 8252 7532 8308
rect 7588 8252 7692 8308
rect 7748 8252 7852 8308
rect 7908 8252 8012 8308
rect 8068 8252 8172 8308
rect 8228 8252 8400 8308
rect 0 8240 8400 8252
rect 0 8146 8400 8160
rect 0 8094 1294 8146
rect 1346 8094 3214 8146
rect 3266 8094 5134 8146
rect 5186 8094 7054 8146
rect 7106 8094 8400 8146
rect 0 8080 8400 8094
rect 0 7988 8400 8000
rect 0 7932 172 7988
rect 228 7932 332 7988
rect 388 7932 492 7988
rect 548 7932 652 7988
rect 708 7932 812 7988
rect 868 7932 972 7988
rect 1028 7932 1132 7988
rect 1188 7932 1452 7988
rect 1508 7932 1612 7988
rect 1668 7932 1772 7988
rect 1828 7932 1932 7988
rect 1988 7932 2092 7988
rect 2148 7932 2252 7988
rect 2308 7932 2412 7988
rect 2468 7932 2572 7988
rect 2628 7932 2732 7988
rect 2788 7932 2892 7988
rect 2948 7932 3052 7988
rect 3108 7932 3372 7988
rect 3428 7932 3532 7988
rect 3588 7932 3692 7988
rect 3748 7932 3852 7988
rect 3908 7932 4012 7988
rect 4068 7932 4172 7988
rect 4228 7932 4332 7988
rect 4388 7932 4492 7988
rect 4548 7932 4652 7988
rect 4708 7932 4812 7988
rect 4868 7932 4972 7988
rect 5028 7932 5292 7988
rect 5348 7932 5452 7988
rect 5508 7932 5612 7988
rect 5668 7932 5772 7988
rect 5828 7932 5932 7988
rect 5988 7932 6092 7988
rect 6148 7932 6252 7988
rect 6308 7932 6412 7988
rect 6468 7932 6572 7988
rect 6628 7932 6732 7988
rect 6788 7932 6892 7988
rect 6948 7932 7212 7988
rect 7268 7932 7372 7988
rect 7428 7932 7532 7988
rect 7588 7932 7692 7988
rect 7748 7932 7852 7988
rect 7908 7932 8012 7988
rect 8068 7932 8172 7988
rect 8228 7932 8400 7988
rect 0 7920 8400 7932
rect 320 7688 400 7720
rect 320 7632 332 7688
rect 388 7632 400 7688
rect 320 7626 334 7632
rect 386 7626 400 7632
rect 320 7614 400 7626
rect 320 7608 334 7614
rect 386 7608 400 7614
rect 320 7552 332 7608
rect 388 7552 400 7608
rect 320 7520 400 7552
rect 320 7088 400 7120
rect 320 7032 332 7088
rect 388 7032 400 7088
rect 320 7026 334 7032
rect 386 7026 400 7032
rect 320 7014 400 7026
rect 320 7008 334 7014
rect 386 7008 400 7014
rect 320 6952 332 7008
rect 388 6952 400 7008
rect 320 6920 400 6952
rect 0 6708 8400 6720
rect 0 6652 172 6708
rect 228 6652 332 6708
rect 388 6652 492 6708
rect 548 6652 652 6708
rect 708 6652 812 6708
rect 868 6652 972 6708
rect 1028 6652 1132 6708
rect 1188 6652 1452 6708
rect 1508 6652 1612 6708
rect 1668 6652 1772 6708
rect 1828 6652 1932 6708
rect 1988 6652 2092 6708
rect 2148 6652 2252 6708
rect 2308 6652 2412 6708
rect 2468 6652 2572 6708
rect 2628 6652 2732 6708
rect 2788 6652 2892 6708
rect 2948 6652 3052 6708
rect 3108 6652 3372 6708
rect 3428 6652 3532 6708
rect 3588 6652 3692 6708
rect 3748 6652 3852 6708
rect 3908 6652 4012 6708
rect 4068 6652 4172 6708
rect 4228 6652 4332 6708
rect 4388 6652 4492 6708
rect 4548 6652 4652 6708
rect 4708 6652 4812 6708
rect 4868 6652 4972 6708
rect 5028 6652 5292 6708
rect 5348 6652 5452 6708
rect 5508 6652 5612 6708
rect 5668 6652 5772 6708
rect 5828 6652 5932 6708
rect 5988 6652 6092 6708
rect 6148 6652 6252 6708
rect 6308 6652 6412 6708
rect 6468 6652 6572 6708
rect 6628 6652 6732 6708
rect 6788 6652 6892 6708
rect 6948 6652 7212 6708
rect 7268 6652 7372 6708
rect 7428 6652 7532 6708
rect 7588 6652 7692 6708
rect 7748 6652 7852 6708
rect 7908 6652 8172 6708
rect 8228 6652 8400 6708
rect 0 6640 8400 6652
rect 0 6546 8400 6560
rect 0 6494 1294 6546
rect 1346 6494 3214 6546
rect 3266 6494 5134 6546
rect 5186 6494 7054 6546
rect 7106 6494 8400 6546
rect 0 6480 8400 6494
rect 0 6388 8400 6400
rect 0 6332 172 6388
rect 228 6332 332 6388
rect 388 6332 492 6388
rect 548 6332 652 6388
rect 708 6332 812 6388
rect 868 6332 972 6388
rect 1028 6332 1132 6388
rect 1188 6332 1452 6388
rect 1508 6332 1612 6388
rect 1668 6332 1772 6388
rect 1828 6332 1932 6388
rect 1988 6332 2092 6388
rect 2148 6332 2252 6388
rect 2308 6332 2412 6388
rect 2468 6332 2572 6388
rect 2628 6332 2732 6388
rect 2788 6332 2892 6388
rect 2948 6332 3052 6388
rect 3108 6332 3372 6388
rect 3428 6332 3532 6388
rect 3588 6332 3692 6388
rect 3748 6332 3852 6388
rect 3908 6332 4012 6388
rect 4068 6332 4172 6388
rect 4228 6332 4332 6388
rect 4388 6332 4492 6388
rect 4548 6332 4652 6388
rect 4708 6332 4812 6388
rect 4868 6332 4972 6388
rect 5028 6332 5292 6388
rect 5348 6332 5452 6388
rect 5508 6332 5612 6388
rect 5668 6332 5772 6388
rect 5828 6332 5932 6388
rect 5988 6332 6092 6388
rect 6148 6332 6252 6388
rect 6308 6332 6412 6388
rect 6468 6332 6572 6388
rect 6628 6332 6732 6388
rect 6788 6332 6892 6388
rect 6948 6332 7212 6388
rect 7268 6332 7372 6388
rect 7428 6332 7532 6388
rect 7588 6332 7692 6388
rect 7748 6332 7852 6388
rect 7908 6332 8172 6388
rect 8228 6332 8400 6388
rect 0 6320 8400 6332
rect 0 6228 8400 6240
rect 0 6172 172 6228
rect 228 6172 332 6228
rect 388 6172 492 6228
rect 548 6172 652 6228
rect 708 6172 812 6228
rect 868 6172 972 6228
rect 1028 6172 1132 6228
rect 1188 6172 1292 6228
rect 1348 6172 1452 6228
rect 1508 6172 1612 6228
rect 1668 6172 1772 6228
rect 1828 6172 1932 6228
rect 1988 6172 2092 6228
rect 2148 6172 2252 6228
rect 2308 6172 2412 6228
rect 2468 6172 2572 6228
rect 2628 6172 2732 6228
rect 2788 6172 2892 6228
rect 2948 6172 3052 6228
rect 3108 6172 3212 6228
rect 3268 6172 3372 6228
rect 3428 6172 3532 6228
rect 3588 6172 3692 6228
rect 3748 6172 3852 6228
rect 3908 6172 4012 6228
rect 4068 6172 4172 6228
rect 4228 6172 4332 6228
rect 4388 6172 4492 6228
rect 4548 6172 4652 6228
rect 4708 6172 4812 6228
rect 4868 6172 4972 6228
rect 5028 6172 5132 6228
rect 5188 6172 5292 6228
rect 5348 6172 5452 6228
rect 5508 6172 5612 6228
rect 5668 6172 5772 6228
rect 5828 6172 5932 6228
rect 5988 6172 6092 6228
rect 6148 6172 6252 6228
rect 6308 6172 6412 6228
rect 6468 6172 6572 6228
rect 6628 6172 6732 6228
rect 6788 6172 6892 6228
rect 6948 6172 7052 6228
rect 7108 6172 7212 6228
rect 7268 6172 7372 6228
rect 7428 6172 7532 6228
rect 7588 6172 7692 6228
rect 7748 6172 7852 6228
rect 7908 6172 8172 6228
rect 8228 6172 8400 6228
rect 0 6160 8400 6172
rect 0 6066 8400 6080
rect 0 6014 8014 6066
rect 8066 6014 8400 6066
rect 0 6000 8400 6014
rect 0 5908 8400 5920
rect 0 5852 172 5908
rect 228 5852 332 5908
rect 388 5852 492 5908
rect 548 5852 652 5908
rect 708 5852 812 5908
rect 868 5852 972 5908
rect 1028 5852 1132 5908
rect 1188 5852 1292 5908
rect 1348 5852 1452 5908
rect 1508 5852 1612 5908
rect 1668 5852 1772 5908
rect 1828 5852 1932 5908
rect 1988 5852 2092 5908
rect 2148 5852 2252 5908
rect 2308 5852 2412 5908
rect 2468 5852 2572 5908
rect 2628 5852 2732 5908
rect 2788 5852 2892 5908
rect 2948 5852 3052 5908
rect 3108 5852 3212 5908
rect 3268 5852 3372 5908
rect 3428 5852 3532 5908
rect 3588 5852 3692 5908
rect 3748 5852 3852 5908
rect 3908 5852 4012 5908
rect 4068 5852 4172 5908
rect 4228 5852 4332 5908
rect 4388 5852 4492 5908
rect 4548 5852 4652 5908
rect 4708 5852 4812 5908
rect 4868 5852 4972 5908
rect 5028 5852 5132 5908
rect 5188 5852 5292 5908
rect 5348 5852 5452 5908
rect 5508 5852 5612 5908
rect 5668 5852 5772 5908
rect 5828 5852 5932 5908
rect 5988 5852 6092 5908
rect 6148 5852 6252 5908
rect 6308 5852 6412 5908
rect 6468 5852 6572 5908
rect 6628 5852 6732 5908
rect 6788 5852 6892 5908
rect 6948 5852 7052 5908
rect 7108 5852 7212 5908
rect 7268 5852 7372 5908
rect 7428 5852 7532 5908
rect 7588 5852 7692 5908
rect 7748 5852 7852 5908
rect 7908 5852 8172 5908
rect 8228 5852 8400 5908
rect 0 5840 8400 5852
rect 0 5748 8400 5760
rect 0 5692 172 5748
rect 228 5692 332 5748
rect 388 5692 492 5748
rect 548 5692 652 5748
rect 708 5692 812 5748
rect 868 5692 972 5748
rect 1028 5692 1132 5748
rect 1188 5692 1452 5748
rect 1508 5692 1612 5748
rect 1668 5692 1772 5748
rect 1828 5692 1932 5748
rect 1988 5692 2092 5748
rect 2148 5692 2252 5748
rect 2308 5692 2412 5748
rect 2468 5692 2572 5748
rect 2628 5692 2732 5748
rect 2788 5692 2892 5748
rect 2948 5692 3052 5748
rect 3108 5692 3372 5748
rect 3428 5692 3532 5748
rect 3588 5692 3692 5748
rect 3748 5692 3852 5748
rect 3908 5692 4012 5748
rect 4068 5692 4172 5748
rect 4228 5692 4332 5748
rect 4388 5692 4492 5748
rect 4548 5692 4652 5748
rect 4708 5692 4812 5748
rect 4868 5692 4972 5748
rect 5028 5692 5292 5748
rect 5348 5692 5452 5748
rect 5508 5692 5612 5748
rect 5668 5692 5772 5748
rect 5828 5692 5932 5748
rect 5988 5692 6092 5748
rect 6148 5692 6252 5748
rect 6308 5692 6412 5748
rect 6468 5692 6572 5748
rect 6628 5692 6732 5748
rect 6788 5692 6892 5748
rect 6948 5692 7212 5748
rect 7268 5692 7372 5748
rect 7428 5692 7532 5748
rect 7588 5692 7692 5748
rect 7748 5692 7852 5748
rect 7908 5692 8172 5748
rect 8228 5692 8400 5748
rect 0 5680 8400 5692
rect 0 5586 8400 5600
rect 0 5534 1294 5586
rect 1346 5534 3214 5586
rect 3266 5534 5134 5586
rect 5186 5534 7054 5586
rect 7106 5534 8400 5586
rect 0 5520 8400 5534
rect 0 5428 8400 5440
rect 0 5372 172 5428
rect 228 5372 332 5428
rect 388 5372 492 5428
rect 548 5372 652 5428
rect 708 5372 812 5428
rect 868 5372 972 5428
rect 1028 5372 1132 5428
rect 1188 5372 1452 5428
rect 1508 5372 1612 5428
rect 1668 5372 1772 5428
rect 1828 5372 1932 5428
rect 1988 5372 2092 5428
rect 2148 5372 2252 5428
rect 2308 5372 2412 5428
rect 2468 5372 2572 5428
rect 2628 5372 2732 5428
rect 2788 5372 2892 5428
rect 2948 5372 3052 5428
rect 3108 5372 3372 5428
rect 3428 5372 3532 5428
rect 3588 5372 3692 5428
rect 3748 5372 3852 5428
rect 3908 5372 4012 5428
rect 4068 5372 4172 5428
rect 4228 5372 4332 5428
rect 4388 5372 4492 5428
rect 4548 5372 4652 5428
rect 4708 5372 4812 5428
rect 4868 5372 4972 5428
rect 5028 5372 5292 5428
rect 5348 5372 5452 5428
rect 5508 5372 5612 5428
rect 5668 5372 5772 5428
rect 5828 5372 5932 5428
rect 5988 5372 6092 5428
rect 6148 5372 6252 5428
rect 6308 5372 6412 5428
rect 6468 5372 6572 5428
rect 6628 5372 6732 5428
rect 6788 5372 6892 5428
rect 6948 5372 7212 5428
rect 7268 5372 7372 5428
rect 7428 5372 7532 5428
rect 7588 5372 7692 5428
rect 7748 5372 7852 5428
rect 7908 5372 8172 5428
rect 8228 5372 8400 5428
rect 0 5360 8400 5372
rect 320 4754 400 4800
rect 320 4748 334 4754
rect 386 4748 400 4754
rect 320 4692 332 4748
rect 388 4692 400 4748
rect 320 4690 400 4692
rect 320 4668 334 4690
rect 386 4668 400 4690
rect 320 4612 332 4668
rect 388 4612 400 4668
rect 320 4588 334 4612
rect 386 4588 400 4612
rect 320 4532 332 4588
rect 388 4532 400 4588
rect 320 4510 334 4532
rect 386 4510 400 4532
rect 320 4508 400 4510
rect 320 4452 332 4508
rect 388 4452 400 4508
rect 320 4446 334 4452
rect 386 4446 400 4452
rect 320 4400 400 4446
rect 8000 3634 8080 3680
rect 8000 3628 8014 3634
rect 8066 3628 8080 3634
rect 8000 3572 8012 3628
rect 8068 3572 8080 3628
rect 8000 3570 8080 3572
rect 8000 3548 8014 3570
rect 8066 3548 8080 3570
rect 8000 3492 8012 3548
rect 8068 3492 8080 3548
rect 8000 3468 8014 3492
rect 8066 3468 8080 3492
rect 8000 3412 8012 3468
rect 8068 3412 8080 3468
rect 8000 3390 8014 3412
rect 8066 3390 8080 3412
rect 8000 3388 8080 3390
rect 8000 3332 8012 3388
rect 8068 3332 8080 3388
rect 8000 3326 8014 3332
rect 8066 3326 8080 3332
rect 8000 3280 8080 3326
rect 0 2788 8400 2800
rect 0 2732 12 2788
rect 68 2732 172 2788
rect 228 2732 332 2788
rect 388 2732 492 2788
rect 548 2732 652 2788
rect 708 2732 812 2788
rect 868 2732 972 2788
rect 1028 2732 1132 2788
rect 1188 2732 1452 2788
rect 1508 2732 1612 2788
rect 1668 2732 1772 2788
rect 1828 2732 1932 2788
rect 1988 2732 2092 2788
rect 2148 2732 2252 2788
rect 2308 2732 2412 2788
rect 2468 2732 2572 2788
rect 2628 2732 2732 2788
rect 2788 2732 2892 2788
rect 2948 2732 3052 2788
rect 3108 2732 3372 2788
rect 3428 2732 3532 2788
rect 3588 2732 3692 2788
rect 3748 2732 3852 2788
rect 3908 2732 4012 2788
rect 4068 2732 4172 2788
rect 4228 2732 4332 2788
rect 4388 2732 4492 2788
rect 4548 2732 4652 2788
rect 4708 2732 4812 2788
rect 4868 2732 4972 2788
rect 5028 2732 5292 2788
rect 5348 2732 5452 2788
rect 5508 2732 5612 2788
rect 5668 2732 5772 2788
rect 5828 2732 5932 2788
rect 5988 2732 6092 2788
rect 6148 2732 6252 2788
rect 6308 2732 6412 2788
rect 6468 2732 6572 2788
rect 6628 2732 6732 2788
rect 6788 2732 6892 2788
rect 6948 2732 7212 2788
rect 7268 2732 7372 2788
rect 7428 2732 7532 2788
rect 7588 2732 7692 2788
rect 7748 2732 7852 2788
rect 7908 2732 8012 2788
rect 8068 2732 8172 2788
rect 8228 2732 8332 2788
rect 8388 2732 8400 2788
rect 0 2720 8400 2732
rect 0 2626 8400 2640
rect 0 2574 1294 2626
rect 1346 2574 3214 2626
rect 3266 2574 5134 2626
rect 5186 2574 7054 2626
rect 7106 2574 8400 2626
rect 0 2560 8400 2574
rect 0 2468 8400 2480
rect 0 2412 12 2468
rect 68 2412 172 2468
rect 228 2412 332 2468
rect 388 2412 492 2468
rect 548 2412 652 2468
rect 708 2412 812 2468
rect 868 2412 972 2468
rect 1028 2412 1132 2468
rect 1188 2412 1452 2468
rect 1508 2412 1612 2468
rect 1668 2412 1772 2468
rect 1828 2412 1932 2468
rect 1988 2412 2092 2468
rect 2148 2412 2252 2468
rect 2308 2412 2412 2468
rect 2468 2412 2572 2468
rect 2628 2412 2732 2468
rect 2788 2412 2892 2468
rect 2948 2412 3052 2468
rect 3108 2412 3372 2468
rect 3428 2412 3532 2468
rect 3588 2412 3692 2468
rect 3748 2412 3852 2468
rect 3908 2412 4012 2468
rect 4068 2412 4172 2468
rect 4228 2412 4332 2468
rect 4388 2412 4492 2468
rect 4548 2412 4652 2468
rect 4708 2412 4812 2468
rect 4868 2412 4972 2468
rect 5028 2412 5292 2468
rect 5348 2412 5452 2468
rect 5508 2412 5612 2468
rect 5668 2412 5772 2468
rect 5828 2412 5932 2468
rect 5988 2412 6092 2468
rect 6148 2412 6252 2468
rect 6308 2412 6412 2468
rect 6468 2412 6572 2468
rect 6628 2412 6732 2468
rect 6788 2412 6892 2468
rect 6948 2412 7212 2468
rect 7268 2412 7372 2468
rect 7428 2412 7532 2468
rect 7588 2412 7692 2468
rect 7748 2412 7852 2468
rect 7908 2412 8012 2468
rect 8068 2412 8172 2468
rect 8228 2412 8332 2468
rect 8388 2412 8400 2468
rect 0 2400 8400 2412
rect 0 1268 8400 1280
rect 0 1212 172 1268
rect 228 1212 332 1268
rect 388 1212 492 1268
rect 548 1212 652 1268
rect 708 1212 812 1268
rect 868 1212 972 1268
rect 1028 1212 1132 1268
rect 1188 1212 1452 1268
rect 1508 1212 1612 1268
rect 1668 1212 1772 1268
rect 1828 1212 1932 1268
rect 1988 1212 2092 1268
rect 2148 1212 2252 1268
rect 2308 1212 2412 1268
rect 2468 1212 2572 1268
rect 2628 1212 2732 1268
rect 2788 1212 2892 1268
rect 2948 1212 3052 1268
rect 3108 1212 3372 1268
rect 3428 1212 3532 1268
rect 3588 1212 3692 1268
rect 3748 1212 3852 1268
rect 3908 1212 4012 1268
rect 4068 1212 4172 1268
rect 4228 1212 4332 1268
rect 4388 1212 4492 1268
rect 4548 1212 4652 1268
rect 4708 1212 4812 1268
rect 4868 1212 4972 1268
rect 5028 1212 5292 1268
rect 5348 1212 5452 1268
rect 5508 1212 5612 1268
rect 5668 1212 5772 1268
rect 5828 1212 5932 1268
rect 5988 1212 6092 1268
rect 6148 1212 6252 1268
rect 6308 1212 6412 1268
rect 6468 1212 6572 1268
rect 6628 1212 6732 1268
rect 6788 1212 6892 1268
rect 6948 1212 7212 1268
rect 7268 1212 7372 1268
rect 7428 1212 7532 1268
rect 7588 1212 7692 1268
rect 7748 1212 7852 1268
rect 7908 1212 8012 1268
rect 8068 1212 8172 1268
rect 8228 1212 8400 1268
rect 0 1200 8400 1212
rect 0 1106 8400 1120
rect 0 1054 1294 1106
rect 1346 1054 3214 1106
rect 3266 1054 5134 1106
rect 5186 1054 7054 1106
rect 7106 1054 8014 1106
rect 8066 1054 8400 1106
rect 0 1040 8400 1054
rect 0 948 8400 960
rect 0 892 172 948
rect 228 892 332 948
rect 388 892 492 948
rect 548 892 652 948
rect 708 892 812 948
rect 868 892 972 948
rect 1028 892 1132 948
rect 1188 892 1452 948
rect 1508 892 1612 948
rect 1668 892 1772 948
rect 1828 892 1932 948
rect 1988 892 2092 948
rect 2148 892 2252 948
rect 2308 892 2412 948
rect 2468 892 2572 948
rect 2628 892 2732 948
rect 2788 892 2892 948
rect 2948 892 3052 948
rect 3108 892 3372 948
rect 3428 892 3532 948
rect 3588 892 3692 948
rect 3748 892 3852 948
rect 3908 892 4012 948
rect 4068 892 4172 948
rect 4228 892 4332 948
rect 4388 892 4492 948
rect 4548 892 4652 948
rect 4708 892 4812 948
rect 4868 892 4972 948
rect 5028 892 5292 948
rect 5348 892 5452 948
rect 5508 892 5612 948
rect 5668 892 5772 948
rect 5828 892 5932 948
rect 5988 892 6092 948
rect 6148 892 6252 948
rect 6308 892 6412 948
rect 6468 892 6572 948
rect 6628 892 6732 948
rect 6788 892 6892 948
rect 6948 892 7212 948
rect 7268 892 7372 948
rect 7428 892 7532 948
rect 7588 892 7692 948
rect 7748 892 7852 948
rect 7908 892 8172 948
rect 8228 892 8400 948
rect 0 880 8400 892
rect 0 786 8400 800
rect 0 734 8014 786
rect 8066 734 8400 786
rect 0 720 8400 734
rect 0 628 8400 640
rect 0 572 172 628
rect 228 572 332 628
rect 388 572 492 628
rect 548 572 652 628
rect 708 572 812 628
rect 868 572 972 628
rect 1028 572 1132 628
rect 1188 572 1452 628
rect 1508 572 1612 628
rect 1668 572 1772 628
rect 1828 572 1932 628
rect 1988 572 2092 628
rect 2148 572 2252 628
rect 2308 572 2412 628
rect 2468 572 2572 628
rect 2628 572 2732 628
rect 2788 572 2892 628
rect 2948 572 3052 628
rect 3108 572 3372 628
rect 3428 572 3532 628
rect 3588 572 3692 628
rect 3748 572 3852 628
rect 3908 572 4012 628
rect 4068 572 4172 628
rect 4228 572 4332 628
rect 4388 572 4492 628
rect 4548 572 4652 628
rect 4708 572 4812 628
rect 4868 572 4972 628
rect 5028 572 5292 628
rect 5348 572 5452 628
rect 5508 572 5612 628
rect 5668 572 5772 628
rect 5828 572 5932 628
rect 5988 572 6092 628
rect 6148 572 6252 628
rect 6308 572 6412 628
rect 6468 572 6572 628
rect 6628 572 6732 628
rect 6788 572 6892 628
rect 6948 572 7212 628
rect 7268 572 7372 628
rect 7428 572 7532 628
rect 7588 572 7692 628
rect 7748 572 7852 628
rect 7908 572 8012 628
rect 8068 572 8172 628
rect 8228 572 8400 628
rect 0 560 8400 572
rect 320 328 400 360
rect 320 272 332 328
rect 388 272 400 328
rect 320 266 334 272
rect 386 266 400 272
rect 320 254 400 266
rect 320 248 334 254
rect 386 248 400 254
rect 320 192 332 248
rect 388 192 400 248
rect 320 160 400 192
rect 0 -92 8400 -80
rect 0 -148 172 -92
rect 228 -148 332 -92
rect 388 -148 492 -92
rect 548 -148 652 -92
rect 708 -148 812 -92
rect 868 -148 972 -92
rect 1028 -148 1132 -92
rect 1188 -148 1452 -92
rect 1508 -148 1612 -92
rect 1668 -148 1772 -92
rect 1828 -148 1932 -92
rect 1988 -148 2092 -92
rect 2148 -148 2252 -92
rect 2308 -148 2412 -92
rect 2468 -148 2572 -92
rect 2628 -148 2732 -92
rect 2788 -148 2892 -92
rect 2948 -148 3052 -92
rect 3108 -148 3372 -92
rect 3428 -148 3532 -92
rect 3588 -148 3692 -92
rect 3748 -148 3852 -92
rect 3908 -148 4012 -92
rect 4068 -148 4172 -92
rect 4228 -148 4332 -92
rect 4388 -148 4492 -92
rect 4548 -148 4652 -92
rect 4708 -148 4812 -92
rect 4868 -148 4972 -92
rect 5028 -148 5292 -92
rect 5348 -148 5452 -92
rect 5508 -148 5612 -92
rect 5668 -148 5772 -92
rect 5828 -148 5932 -92
rect 5988 -148 6092 -92
rect 6148 -148 6252 -92
rect 6308 -148 6412 -92
rect 6468 -148 6572 -92
rect 6628 -148 6732 -92
rect 6788 -148 6892 -92
rect 6948 -148 7212 -92
rect 7268 -148 7372 -92
rect 7428 -148 7532 -92
rect 7588 -148 7692 -92
rect 7748 -148 7852 -92
rect 7908 -148 8172 -92
rect 8228 -148 8400 -92
rect 0 -160 8400 -148
rect 0 -254 8400 -240
rect 0 -306 1294 -254
rect 1346 -306 3214 -254
rect 3266 -306 5134 -254
rect 5186 -306 7054 -254
rect 7106 -306 8014 -254
rect 8066 -306 8400 -254
rect 0 -320 8400 -306
rect 0 -412 8400 -400
rect 0 -468 172 -412
rect 228 -468 332 -412
rect 388 -468 492 -412
rect 548 -468 652 -412
rect 708 -468 812 -412
rect 868 -468 972 -412
rect 1028 -468 1132 -412
rect 1188 -468 1452 -412
rect 1508 -468 1612 -412
rect 1668 -468 1772 -412
rect 1828 -468 1932 -412
rect 1988 -468 2092 -412
rect 2148 -468 2252 -412
rect 2308 -468 2412 -412
rect 2468 -468 2572 -412
rect 2628 -468 2732 -412
rect 2788 -468 2892 -412
rect 2948 -468 3052 -412
rect 3108 -468 3372 -412
rect 3428 -468 3532 -412
rect 3588 -468 3692 -412
rect 3748 -468 3852 -412
rect 3908 -468 4012 -412
rect 4068 -468 4172 -412
rect 4228 -468 4332 -412
rect 4388 -468 4492 -412
rect 4548 -468 4652 -412
rect 4708 -468 4812 -412
rect 4868 -468 4972 -412
rect 5028 -468 5292 -412
rect 5348 -468 5452 -412
rect 5508 -468 5612 -412
rect 5668 -468 5772 -412
rect 5828 -468 5932 -412
rect 5988 -468 6092 -412
rect 6148 -468 6252 -412
rect 6308 -468 6412 -412
rect 6468 -468 6572 -412
rect 6628 -468 6732 -412
rect 6788 -468 6892 -412
rect 6948 -468 7212 -412
rect 7268 -468 7372 -412
rect 7428 -468 7532 -412
rect 7588 -468 7692 -412
rect 7748 -468 7852 -412
rect 7908 -468 8172 -412
rect 8228 -468 8400 -412
rect 0 -480 8400 -468
rect 320 -712 400 -680
rect 320 -768 332 -712
rect 388 -768 400 -712
rect 320 -774 334 -768
rect 386 -774 400 -768
rect 320 -786 400 -774
rect 320 -792 334 -786
rect 386 -792 400 -786
rect 320 -848 332 -792
rect 388 -848 400 -792
rect 320 -880 400 -848
<< via2 >>
rect 332 9662 334 9708
rect 334 9662 386 9708
rect 386 9662 388 9708
rect 332 9652 388 9662
rect 332 9598 334 9628
rect 334 9598 386 9628
rect 386 9598 388 9628
rect 332 9586 388 9598
rect 332 9572 334 9586
rect 334 9572 386 9586
rect 386 9572 388 9586
rect 332 9534 334 9548
rect 334 9534 386 9548
rect 386 9534 388 9548
rect 332 9522 388 9534
rect 332 9492 334 9522
rect 334 9492 386 9522
rect 386 9492 388 9522
rect 332 9458 388 9468
rect 332 9412 334 9458
rect 334 9412 386 9458
rect 386 9412 388 9458
rect 172 8732 228 8788
rect 332 8732 388 8788
rect 492 8732 548 8788
rect 652 8732 708 8788
rect 812 8732 868 8788
rect 972 8732 1028 8788
rect 1132 8732 1188 8788
rect 1452 8732 1508 8788
rect 1612 8732 1668 8788
rect 1772 8732 1828 8788
rect 1932 8732 1988 8788
rect 2092 8732 2148 8788
rect 2252 8732 2308 8788
rect 2412 8732 2468 8788
rect 2572 8732 2628 8788
rect 2732 8732 2788 8788
rect 2892 8732 2948 8788
rect 3052 8732 3108 8788
rect 3372 8732 3428 8788
rect 3532 8732 3588 8788
rect 3692 8732 3748 8788
rect 3852 8732 3908 8788
rect 4012 8732 4068 8788
rect 4172 8732 4228 8788
rect 4332 8732 4388 8788
rect 4492 8732 4548 8788
rect 4652 8732 4708 8788
rect 4812 8732 4868 8788
rect 4972 8732 5028 8788
rect 5292 8732 5348 8788
rect 5452 8732 5508 8788
rect 5612 8732 5668 8788
rect 5772 8732 5828 8788
rect 5932 8732 5988 8788
rect 6092 8732 6148 8788
rect 6252 8732 6308 8788
rect 6412 8732 6468 8788
rect 6572 8732 6628 8788
rect 6732 8732 6788 8788
rect 6892 8732 6948 8788
rect 7212 8732 7268 8788
rect 7372 8732 7428 8788
rect 7532 8732 7588 8788
rect 7692 8732 7748 8788
rect 7852 8732 7908 8788
rect 8012 8732 8068 8788
rect 8172 8732 8228 8788
rect 172 8466 228 8468
rect 172 8414 174 8466
rect 174 8414 226 8466
rect 226 8414 228 8466
rect 172 8412 228 8414
rect 332 8412 388 8468
rect 492 8412 548 8468
rect 652 8412 708 8468
rect 812 8412 868 8468
rect 972 8412 1028 8468
rect 1132 8412 1188 8468
rect 1452 8412 1508 8468
rect 1612 8412 1668 8468
rect 1772 8412 1828 8468
rect 1932 8412 1988 8468
rect 2092 8412 2148 8468
rect 2252 8412 2308 8468
rect 2412 8412 2468 8468
rect 2572 8412 2628 8468
rect 2732 8412 2788 8468
rect 2892 8412 2948 8468
rect 3052 8412 3108 8468
rect 3372 8412 3428 8468
rect 3532 8412 3588 8468
rect 3692 8412 3748 8468
rect 3852 8412 3908 8468
rect 4012 8412 4068 8468
rect 4172 8412 4228 8468
rect 4332 8412 4388 8468
rect 4492 8412 4548 8468
rect 4652 8412 4708 8468
rect 4812 8412 4868 8468
rect 4972 8412 5028 8468
rect 5292 8412 5348 8468
rect 5452 8412 5508 8468
rect 5612 8412 5668 8468
rect 5772 8412 5828 8468
rect 5932 8412 5988 8468
rect 6092 8412 6148 8468
rect 6252 8412 6308 8468
rect 6412 8412 6468 8468
rect 6572 8412 6628 8468
rect 6732 8412 6788 8468
rect 6892 8412 6948 8468
rect 7212 8412 7268 8468
rect 7372 8412 7428 8468
rect 7532 8412 7588 8468
rect 7692 8412 7748 8468
rect 7852 8412 7908 8468
rect 8012 8412 8068 8468
rect 8172 8466 8228 8468
rect 8172 8414 8174 8466
rect 8174 8414 8226 8466
rect 8226 8414 8228 8466
rect 8172 8412 8228 8414
rect 172 8306 228 8308
rect 172 8254 174 8306
rect 174 8254 226 8306
rect 226 8254 228 8306
rect 172 8252 228 8254
rect 332 8252 388 8308
rect 492 8252 548 8308
rect 652 8252 708 8308
rect 812 8252 868 8308
rect 972 8252 1028 8308
rect 1132 8252 1188 8308
rect 1452 8252 1508 8308
rect 1612 8252 1668 8308
rect 1772 8252 1828 8308
rect 1932 8252 1988 8308
rect 2092 8252 2148 8308
rect 2252 8252 2308 8308
rect 2412 8252 2468 8308
rect 2572 8252 2628 8308
rect 2732 8252 2788 8308
rect 2892 8252 2948 8308
rect 3052 8252 3108 8308
rect 3372 8252 3428 8308
rect 3532 8252 3588 8308
rect 3692 8252 3748 8308
rect 3852 8252 3908 8308
rect 4012 8252 4068 8308
rect 4172 8252 4228 8308
rect 4332 8252 4388 8308
rect 4492 8252 4548 8308
rect 4652 8252 4708 8308
rect 4812 8252 4868 8308
rect 4972 8252 5028 8308
rect 5292 8252 5348 8308
rect 5452 8252 5508 8308
rect 5612 8252 5668 8308
rect 5772 8252 5828 8308
rect 5932 8252 5988 8308
rect 6092 8252 6148 8308
rect 6252 8252 6308 8308
rect 6412 8252 6468 8308
rect 6572 8252 6628 8308
rect 6732 8252 6788 8308
rect 6892 8252 6948 8308
rect 7212 8252 7268 8308
rect 7372 8252 7428 8308
rect 7532 8252 7588 8308
rect 7692 8252 7748 8308
rect 7852 8252 7908 8308
rect 8012 8252 8068 8308
rect 8172 8306 8228 8308
rect 8172 8254 8174 8306
rect 8174 8254 8226 8306
rect 8226 8254 8228 8306
rect 8172 8252 8228 8254
rect 172 7932 228 7988
rect 332 7932 388 7988
rect 492 7932 548 7988
rect 652 7932 708 7988
rect 812 7932 868 7988
rect 972 7932 1028 7988
rect 1132 7932 1188 7988
rect 1452 7932 1508 7988
rect 1612 7932 1668 7988
rect 1772 7932 1828 7988
rect 1932 7932 1988 7988
rect 2092 7932 2148 7988
rect 2252 7932 2308 7988
rect 2412 7932 2468 7988
rect 2572 7932 2628 7988
rect 2732 7932 2788 7988
rect 2892 7932 2948 7988
rect 3052 7932 3108 7988
rect 3372 7932 3428 7988
rect 3532 7932 3588 7988
rect 3692 7932 3748 7988
rect 3852 7932 3908 7988
rect 4012 7932 4068 7988
rect 4172 7932 4228 7988
rect 4332 7932 4388 7988
rect 4492 7932 4548 7988
rect 4652 7932 4708 7988
rect 4812 7932 4868 7988
rect 4972 7932 5028 7988
rect 5292 7932 5348 7988
rect 5452 7932 5508 7988
rect 5612 7932 5668 7988
rect 5772 7932 5828 7988
rect 5932 7932 5988 7988
rect 6092 7932 6148 7988
rect 6252 7932 6308 7988
rect 6412 7932 6468 7988
rect 6572 7932 6628 7988
rect 6732 7932 6788 7988
rect 6892 7932 6948 7988
rect 7212 7932 7268 7988
rect 7372 7932 7428 7988
rect 7532 7932 7588 7988
rect 7692 7932 7748 7988
rect 7852 7932 7908 7988
rect 8012 7932 8068 7988
rect 8172 7932 8228 7988
rect 332 7678 388 7688
rect 332 7632 334 7678
rect 334 7632 386 7678
rect 386 7632 388 7678
rect 332 7562 334 7608
rect 334 7562 386 7608
rect 386 7562 388 7608
rect 332 7552 388 7562
rect 332 7078 388 7088
rect 332 7032 334 7078
rect 334 7032 386 7078
rect 386 7032 388 7078
rect 332 6962 334 7008
rect 334 6962 386 7008
rect 386 6962 388 7008
rect 332 6952 388 6962
rect 172 6652 228 6708
rect 332 6652 388 6708
rect 492 6652 548 6708
rect 652 6652 708 6708
rect 812 6652 868 6708
rect 972 6652 1028 6708
rect 1132 6652 1188 6708
rect 1452 6652 1508 6708
rect 1612 6652 1668 6708
rect 1772 6652 1828 6708
rect 1932 6652 1988 6708
rect 2092 6652 2148 6708
rect 2252 6652 2308 6708
rect 2412 6652 2468 6708
rect 2572 6652 2628 6708
rect 2732 6652 2788 6708
rect 2892 6652 2948 6708
rect 3052 6652 3108 6708
rect 3372 6652 3428 6708
rect 3532 6652 3588 6708
rect 3692 6652 3748 6708
rect 3852 6652 3908 6708
rect 4012 6652 4068 6708
rect 4172 6652 4228 6708
rect 4332 6652 4388 6708
rect 4492 6652 4548 6708
rect 4652 6652 4708 6708
rect 4812 6652 4868 6708
rect 4972 6652 5028 6708
rect 5292 6652 5348 6708
rect 5452 6652 5508 6708
rect 5612 6652 5668 6708
rect 5772 6652 5828 6708
rect 5932 6652 5988 6708
rect 6092 6652 6148 6708
rect 6252 6652 6308 6708
rect 6412 6652 6468 6708
rect 6572 6652 6628 6708
rect 6732 6652 6788 6708
rect 6892 6652 6948 6708
rect 7212 6652 7268 6708
rect 7372 6652 7428 6708
rect 7532 6652 7588 6708
rect 7692 6652 7748 6708
rect 7852 6652 7908 6708
rect 8172 6652 8228 6708
rect 172 6386 228 6388
rect 172 6334 174 6386
rect 174 6334 226 6386
rect 226 6334 228 6386
rect 172 6332 228 6334
rect 332 6332 388 6388
rect 492 6332 548 6388
rect 652 6332 708 6388
rect 812 6332 868 6388
rect 972 6332 1028 6388
rect 1132 6332 1188 6388
rect 1452 6332 1508 6388
rect 1612 6332 1668 6388
rect 1772 6332 1828 6388
rect 1932 6332 1988 6388
rect 2092 6332 2148 6388
rect 2252 6332 2308 6388
rect 2412 6332 2468 6388
rect 2572 6332 2628 6388
rect 2732 6332 2788 6388
rect 2892 6332 2948 6388
rect 3052 6332 3108 6388
rect 3372 6332 3428 6388
rect 3532 6332 3588 6388
rect 3692 6332 3748 6388
rect 3852 6332 3908 6388
rect 4012 6332 4068 6388
rect 4172 6332 4228 6388
rect 4332 6332 4388 6388
rect 4492 6332 4548 6388
rect 4652 6332 4708 6388
rect 4812 6332 4868 6388
rect 4972 6332 5028 6388
rect 5292 6332 5348 6388
rect 5452 6332 5508 6388
rect 5612 6332 5668 6388
rect 5772 6332 5828 6388
rect 5932 6332 5988 6388
rect 6092 6332 6148 6388
rect 6252 6332 6308 6388
rect 6412 6332 6468 6388
rect 6572 6332 6628 6388
rect 6732 6332 6788 6388
rect 6892 6332 6948 6388
rect 7212 6332 7268 6388
rect 7372 6332 7428 6388
rect 7532 6332 7588 6388
rect 7692 6332 7748 6388
rect 7852 6332 7908 6388
rect 8172 6386 8228 6388
rect 8172 6334 8174 6386
rect 8174 6334 8226 6386
rect 8226 6334 8228 6386
rect 8172 6332 8228 6334
rect 172 6226 228 6228
rect 172 6174 174 6226
rect 174 6174 226 6226
rect 226 6174 228 6226
rect 172 6172 228 6174
rect 332 6172 388 6228
rect 492 6172 548 6228
rect 652 6172 708 6228
rect 812 6172 868 6228
rect 972 6172 1028 6228
rect 1132 6172 1188 6228
rect 1292 6172 1348 6228
rect 1452 6172 1508 6228
rect 1612 6172 1668 6228
rect 1772 6172 1828 6228
rect 1932 6172 1988 6228
rect 2092 6172 2148 6228
rect 2252 6172 2308 6228
rect 2412 6172 2468 6228
rect 2572 6172 2628 6228
rect 2732 6172 2788 6228
rect 2892 6172 2948 6228
rect 3052 6172 3108 6228
rect 3212 6172 3268 6228
rect 3372 6172 3428 6228
rect 3532 6172 3588 6228
rect 3692 6172 3748 6228
rect 3852 6172 3908 6228
rect 4012 6172 4068 6228
rect 4172 6172 4228 6228
rect 4332 6172 4388 6228
rect 4492 6172 4548 6228
rect 4652 6172 4708 6228
rect 4812 6172 4868 6228
rect 4972 6172 5028 6228
rect 5132 6172 5188 6228
rect 5292 6172 5348 6228
rect 5452 6172 5508 6228
rect 5612 6172 5668 6228
rect 5772 6172 5828 6228
rect 5932 6172 5988 6228
rect 6092 6172 6148 6228
rect 6252 6172 6308 6228
rect 6412 6172 6468 6228
rect 6572 6172 6628 6228
rect 6732 6172 6788 6228
rect 6892 6172 6948 6228
rect 7052 6172 7108 6228
rect 7212 6172 7268 6228
rect 7372 6172 7428 6228
rect 7532 6172 7588 6228
rect 7692 6172 7748 6228
rect 7852 6172 7908 6228
rect 8172 6226 8228 6228
rect 8172 6174 8174 6226
rect 8174 6174 8226 6226
rect 8226 6174 8228 6226
rect 8172 6172 8228 6174
rect 172 5906 228 5908
rect 172 5854 174 5906
rect 174 5854 226 5906
rect 226 5854 228 5906
rect 172 5852 228 5854
rect 332 5852 388 5908
rect 492 5852 548 5908
rect 652 5852 708 5908
rect 812 5852 868 5908
rect 972 5852 1028 5908
rect 1132 5852 1188 5908
rect 1292 5852 1348 5908
rect 1452 5852 1508 5908
rect 1612 5852 1668 5908
rect 1772 5852 1828 5908
rect 1932 5852 1988 5908
rect 2092 5852 2148 5908
rect 2252 5852 2308 5908
rect 2412 5852 2468 5908
rect 2572 5852 2628 5908
rect 2732 5852 2788 5908
rect 2892 5852 2948 5908
rect 3052 5852 3108 5908
rect 3212 5852 3268 5908
rect 3372 5852 3428 5908
rect 3532 5852 3588 5908
rect 3692 5852 3748 5908
rect 3852 5852 3908 5908
rect 4012 5852 4068 5908
rect 4172 5852 4228 5908
rect 4332 5852 4388 5908
rect 4492 5852 4548 5908
rect 4652 5852 4708 5908
rect 4812 5852 4868 5908
rect 4972 5852 5028 5908
rect 5132 5852 5188 5908
rect 5292 5852 5348 5908
rect 5452 5852 5508 5908
rect 5612 5852 5668 5908
rect 5772 5852 5828 5908
rect 5932 5852 5988 5908
rect 6092 5852 6148 5908
rect 6252 5852 6308 5908
rect 6412 5852 6468 5908
rect 6572 5852 6628 5908
rect 6732 5852 6788 5908
rect 6892 5852 6948 5908
rect 7052 5852 7108 5908
rect 7212 5852 7268 5908
rect 7372 5852 7428 5908
rect 7532 5852 7588 5908
rect 7692 5852 7748 5908
rect 7852 5852 7908 5908
rect 8172 5906 8228 5908
rect 8172 5854 8174 5906
rect 8174 5854 8226 5906
rect 8226 5854 8228 5906
rect 8172 5852 8228 5854
rect 172 5746 228 5748
rect 172 5694 174 5746
rect 174 5694 226 5746
rect 226 5694 228 5746
rect 172 5692 228 5694
rect 332 5692 388 5748
rect 492 5692 548 5748
rect 652 5692 708 5748
rect 812 5692 868 5748
rect 972 5692 1028 5748
rect 1132 5692 1188 5748
rect 1452 5692 1508 5748
rect 1612 5692 1668 5748
rect 1772 5692 1828 5748
rect 1932 5692 1988 5748
rect 2092 5692 2148 5748
rect 2252 5692 2308 5748
rect 2412 5692 2468 5748
rect 2572 5692 2628 5748
rect 2732 5692 2788 5748
rect 2892 5692 2948 5748
rect 3052 5692 3108 5748
rect 3372 5692 3428 5748
rect 3532 5692 3588 5748
rect 3692 5692 3748 5748
rect 3852 5692 3908 5748
rect 4012 5692 4068 5748
rect 4172 5692 4228 5748
rect 4332 5692 4388 5748
rect 4492 5692 4548 5748
rect 4652 5692 4708 5748
rect 4812 5692 4868 5748
rect 4972 5692 5028 5748
rect 5292 5692 5348 5748
rect 5452 5692 5508 5748
rect 5612 5692 5668 5748
rect 5772 5692 5828 5748
rect 5932 5692 5988 5748
rect 6092 5692 6148 5748
rect 6252 5692 6308 5748
rect 6412 5692 6468 5748
rect 6572 5692 6628 5748
rect 6732 5692 6788 5748
rect 6892 5692 6948 5748
rect 7212 5692 7268 5748
rect 7372 5692 7428 5748
rect 7532 5692 7588 5748
rect 7692 5692 7748 5748
rect 7852 5692 7908 5748
rect 8172 5746 8228 5748
rect 8172 5694 8174 5746
rect 8174 5694 8226 5746
rect 8226 5694 8228 5746
rect 8172 5692 8228 5694
rect 172 5372 228 5428
rect 332 5372 388 5428
rect 492 5372 548 5428
rect 652 5372 708 5428
rect 812 5372 868 5428
rect 972 5372 1028 5428
rect 1132 5372 1188 5428
rect 1452 5372 1508 5428
rect 1612 5372 1668 5428
rect 1772 5372 1828 5428
rect 1932 5372 1988 5428
rect 2092 5372 2148 5428
rect 2252 5372 2308 5428
rect 2412 5372 2468 5428
rect 2572 5372 2628 5428
rect 2732 5372 2788 5428
rect 2892 5372 2948 5428
rect 3052 5372 3108 5428
rect 3372 5372 3428 5428
rect 3532 5372 3588 5428
rect 3692 5372 3748 5428
rect 3852 5372 3908 5428
rect 4012 5372 4068 5428
rect 4172 5372 4228 5428
rect 4332 5372 4388 5428
rect 4492 5372 4548 5428
rect 4652 5372 4708 5428
rect 4812 5372 4868 5428
rect 4972 5372 5028 5428
rect 5292 5372 5348 5428
rect 5452 5372 5508 5428
rect 5612 5372 5668 5428
rect 5772 5372 5828 5428
rect 5932 5372 5988 5428
rect 6092 5372 6148 5428
rect 6252 5372 6308 5428
rect 6412 5372 6468 5428
rect 6572 5372 6628 5428
rect 6732 5372 6788 5428
rect 6892 5372 6948 5428
rect 7212 5372 7268 5428
rect 7372 5372 7428 5428
rect 7532 5372 7588 5428
rect 7692 5372 7748 5428
rect 7852 5372 7908 5428
rect 8172 5372 8228 5428
rect 332 4702 334 4748
rect 334 4702 386 4748
rect 386 4702 388 4748
rect 332 4692 388 4702
rect 332 4638 334 4668
rect 334 4638 386 4668
rect 386 4638 388 4668
rect 332 4626 388 4638
rect 332 4612 334 4626
rect 334 4612 386 4626
rect 386 4612 388 4626
rect 332 4574 334 4588
rect 334 4574 386 4588
rect 386 4574 388 4588
rect 332 4562 388 4574
rect 332 4532 334 4562
rect 334 4532 386 4562
rect 386 4532 388 4562
rect 332 4498 388 4508
rect 332 4452 334 4498
rect 334 4452 386 4498
rect 386 4452 388 4498
rect 8012 3582 8014 3628
rect 8014 3582 8066 3628
rect 8066 3582 8068 3628
rect 8012 3572 8068 3582
rect 8012 3518 8014 3548
rect 8014 3518 8066 3548
rect 8066 3518 8068 3548
rect 8012 3506 8068 3518
rect 8012 3492 8014 3506
rect 8014 3492 8066 3506
rect 8066 3492 8068 3506
rect 8012 3454 8014 3468
rect 8014 3454 8066 3468
rect 8066 3454 8068 3468
rect 8012 3442 8068 3454
rect 8012 3412 8014 3442
rect 8014 3412 8066 3442
rect 8066 3412 8068 3442
rect 8012 3378 8068 3388
rect 8012 3332 8014 3378
rect 8014 3332 8066 3378
rect 8066 3332 8068 3378
rect 12 2786 68 2788
rect 12 2734 14 2786
rect 14 2734 66 2786
rect 66 2734 68 2786
rect 12 2732 68 2734
rect 172 2786 228 2788
rect 172 2734 174 2786
rect 174 2734 226 2786
rect 226 2734 228 2786
rect 172 2732 228 2734
rect 332 2786 388 2788
rect 332 2734 334 2786
rect 334 2734 386 2786
rect 386 2734 388 2786
rect 332 2732 388 2734
rect 492 2786 548 2788
rect 492 2734 494 2786
rect 494 2734 546 2786
rect 546 2734 548 2786
rect 492 2732 548 2734
rect 652 2786 708 2788
rect 652 2734 654 2786
rect 654 2734 706 2786
rect 706 2734 708 2786
rect 652 2732 708 2734
rect 812 2786 868 2788
rect 812 2734 814 2786
rect 814 2734 866 2786
rect 866 2734 868 2786
rect 812 2732 868 2734
rect 972 2786 1028 2788
rect 972 2734 974 2786
rect 974 2734 1026 2786
rect 1026 2734 1028 2786
rect 972 2732 1028 2734
rect 1132 2786 1188 2788
rect 1132 2734 1134 2786
rect 1134 2734 1186 2786
rect 1186 2734 1188 2786
rect 1132 2732 1188 2734
rect 1452 2786 1508 2788
rect 1452 2734 1454 2786
rect 1454 2734 1506 2786
rect 1506 2734 1508 2786
rect 1452 2732 1508 2734
rect 1612 2786 1668 2788
rect 1612 2734 1614 2786
rect 1614 2734 1666 2786
rect 1666 2734 1668 2786
rect 1612 2732 1668 2734
rect 1772 2786 1828 2788
rect 1772 2734 1774 2786
rect 1774 2734 1826 2786
rect 1826 2734 1828 2786
rect 1772 2732 1828 2734
rect 1932 2786 1988 2788
rect 1932 2734 1934 2786
rect 1934 2734 1986 2786
rect 1986 2734 1988 2786
rect 1932 2732 1988 2734
rect 2092 2786 2148 2788
rect 2092 2734 2094 2786
rect 2094 2734 2146 2786
rect 2146 2734 2148 2786
rect 2092 2732 2148 2734
rect 2252 2786 2308 2788
rect 2252 2734 2254 2786
rect 2254 2734 2306 2786
rect 2306 2734 2308 2786
rect 2252 2732 2308 2734
rect 2412 2786 2468 2788
rect 2412 2734 2414 2786
rect 2414 2734 2466 2786
rect 2466 2734 2468 2786
rect 2412 2732 2468 2734
rect 2572 2786 2628 2788
rect 2572 2734 2574 2786
rect 2574 2734 2626 2786
rect 2626 2734 2628 2786
rect 2572 2732 2628 2734
rect 2732 2786 2788 2788
rect 2732 2734 2734 2786
rect 2734 2734 2786 2786
rect 2786 2734 2788 2786
rect 2732 2732 2788 2734
rect 2892 2786 2948 2788
rect 2892 2734 2894 2786
rect 2894 2734 2946 2786
rect 2946 2734 2948 2786
rect 2892 2732 2948 2734
rect 3052 2786 3108 2788
rect 3052 2734 3054 2786
rect 3054 2734 3106 2786
rect 3106 2734 3108 2786
rect 3052 2732 3108 2734
rect 3372 2786 3428 2788
rect 3372 2734 3374 2786
rect 3374 2734 3426 2786
rect 3426 2734 3428 2786
rect 3372 2732 3428 2734
rect 3532 2786 3588 2788
rect 3532 2734 3534 2786
rect 3534 2734 3586 2786
rect 3586 2734 3588 2786
rect 3532 2732 3588 2734
rect 3692 2786 3748 2788
rect 3692 2734 3694 2786
rect 3694 2734 3746 2786
rect 3746 2734 3748 2786
rect 3692 2732 3748 2734
rect 3852 2786 3908 2788
rect 3852 2734 3854 2786
rect 3854 2734 3906 2786
rect 3906 2734 3908 2786
rect 3852 2732 3908 2734
rect 4012 2786 4068 2788
rect 4012 2734 4014 2786
rect 4014 2734 4066 2786
rect 4066 2734 4068 2786
rect 4012 2732 4068 2734
rect 4172 2786 4228 2788
rect 4172 2734 4174 2786
rect 4174 2734 4226 2786
rect 4226 2734 4228 2786
rect 4172 2732 4228 2734
rect 4332 2786 4388 2788
rect 4332 2734 4334 2786
rect 4334 2734 4386 2786
rect 4386 2734 4388 2786
rect 4332 2732 4388 2734
rect 4492 2786 4548 2788
rect 4492 2734 4494 2786
rect 4494 2734 4546 2786
rect 4546 2734 4548 2786
rect 4492 2732 4548 2734
rect 4652 2786 4708 2788
rect 4652 2734 4654 2786
rect 4654 2734 4706 2786
rect 4706 2734 4708 2786
rect 4652 2732 4708 2734
rect 4812 2786 4868 2788
rect 4812 2734 4814 2786
rect 4814 2734 4866 2786
rect 4866 2734 4868 2786
rect 4812 2732 4868 2734
rect 4972 2786 5028 2788
rect 4972 2734 4974 2786
rect 4974 2734 5026 2786
rect 5026 2734 5028 2786
rect 4972 2732 5028 2734
rect 5292 2786 5348 2788
rect 5292 2734 5294 2786
rect 5294 2734 5346 2786
rect 5346 2734 5348 2786
rect 5292 2732 5348 2734
rect 5452 2786 5508 2788
rect 5452 2734 5454 2786
rect 5454 2734 5506 2786
rect 5506 2734 5508 2786
rect 5452 2732 5508 2734
rect 5612 2786 5668 2788
rect 5612 2734 5614 2786
rect 5614 2734 5666 2786
rect 5666 2734 5668 2786
rect 5612 2732 5668 2734
rect 5772 2786 5828 2788
rect 5772 2734 5774 2786
rect 5774 2734 5826 2786
rect 5826 2734 5828 2786
rect 5772 2732 5828 2734
rect 5932 2786 5988 2788
rect 5932 2734 5934 2786
rect 5934 2734 5986 2786
rect 5986 2734 5988 2786
rect 5932 2732 5988 2734
rect 6092 2786 6148 2788
rect 6092 2734 6094 2786
rect 6094 2734 6146 2786
rect 6146 2734 6148 2786
rect 6092 2732 6148 2734
rect 6252 2786 6308 2788
rect 6252 2734 6254 2786
rect 6254 2734 6306 2786
rect 6306 2734 6308 2786
rect 6252 2732 6308 2734
rect 6412 2786 6468 2788
rect 6412 2734 6414 2786
rect 6414 2734 6466 2786
rect 6466 2734 6468 2786
rect 6412 2732 6468 2734
rect 6572 2786 6628 2788
rect 6572 2734 6574 2786
rect 6574 2734 6626 2786
rect 6626 2734 6628 2786
rect 6572 2732 6628 2734
rect 6732 2786 6788 2788
rect 6732 2734 6734 2786
rect 6734 2734 6786 2786
rect 6786 2734 6788 2786
rect 6732 2732 6788 2734
rect 6892 2786 6948 2788
rect 6892 2734 6894 2786
rect 6894 2734 6946 2786
rect 6946 2734 6948 2786
rect 6892 2732 6948 2734
rect 7212 2786 7268 2788
rect 7212 2734 7214 2786
rect 7214 2734 7266 2786
rect 7266 2734 7268 2786
rect 7212 2732 7268 2734
rect 7372 2786 7428 2788
rect 7372 2734 7374 2786
rect 7374 2734 7426 2786
rect 7426 2734 7428 2786
rect 7372 2732 7428 2734
rect 7532 2786 7588 2788
rect 7532 2734 7534 2786
rect 7534 2734 7586 2786
rect 7586 2734 7588 2786
rect 7532 2732 7588 2734
rect 7692 2786 7748 2788
rect 7692 2734 7694 2786
rect 7694 2734 7746 2786
rect 7746 2734 7748 2786
rect 7692 2732 7748 2734
rect 7852 2786 7908 2788
rect 7852 2734 7854 2786
rect 7854 2734 7906 2786
rect 7906 2734 7908 2786
rect 7852 2732 7908 2734
rect 8012 2786 8068 2788
rect 8012 2734 8014 2786
rect 8014 2734 8066 2786
rect 8066 2734 8068 2786
rect 8012 2732 8068 2734
rect 8172 2786 8228 2788
rect 8172 2734 8174 2786
rect 8174 2734 8226 2786
rect 8226 2734 8228 2786
rect 8172 2732 8228 2734
rect 8332 2786 8388 2788
rect 8332 2734 8334 2786
rect 8334 2734 8386 2786
rect 8386 2734 8388 2786
rect 8332 2732 8388 2734
rect 12 2466 68 2468
rect 12 2414 14 2466
rect 14 2414 66 2466
rect 66 2414 68 2466
rect 12 2412 68 2414
rect 172 2466 228 2468
rect 172 2414 174 2466
rect 174 2414 226 2466
rect 226 2414 228 2466
rect 172 2412 228 2414
rect 332 2466 388 2468
rect 332 2414 334 2466
rect 334 2414 386 2466
rect 386 2414 388 2466
rect 332 2412 388 2414
rect 492 2466 548 2468
rect 492 2414 494 2466
rect 494 2414 546 2466
rect 546 2414 548 2466
rect 492 2412 548 2414
rect 652 2466 708 2468
rect 652 2414 654 2466
rect 654 2414 706 2466
rect 706 2414 708 2466
rect 652 2412 708 2414
rect 812 2466 868 2468
rect 812 2414 814 2466
rect 814 2414 866 2466
rect 866 2414 868 2466
rect 812 2412 868 2414
rect 972 2466 1028 2468
rect 972 2414 974 2466
rect 974 2414 1026 2466
rect 1026 2414 1028 2466
rect 972 2412 1028 2414
rect 1132 2466 1188 2468
rect 1132 2414 1134 2466
rect 1134 2414 1186 2466
rect 1186 2414 1188 2466
rect 1132 2412 1188 2414
rect 1452 2466 1508 2468
rect 1452 2414 1454 2466
rect 1454 2414 1506 2466
rect 1506 2414 1508 2466
rect 1452 2412 1508 2414
rect 1612 2466 1668 2468
rect 1612 2414 1614 2466
rect 1614 2414 1666 2466
rect 1666 2414 1668 2466
rect 1612 2412 1668 2414
rect 1772 2466 1828 2468
rect 1772 2414 1774 2466
rect 1774 2414 1826 2466
rect 1826 2414 1828 2466
rect 1772 2412 1828 2414
rect 1932 2466 1988 2468
rect 1932 2414 1934 2466
rect 1934 2414 1986 2466
rect 1986 2414 1988 2466
rect 1932 2412 1988 2414
rect 2092 2466 2148 2468
rect 2092 2414 2094 2466
rect 2094 2414 2146 2466
rect 2146 2414 2148 2466
rect 2092 2412 2148 2414
rect 2252 2466 2308 2468
rect 2252 2414 2254 2466
rect 2254 2414 2306 2466
rect 2306 2414 2308 2466
rect 2252 2412 2308 2414
rect 2412 2466 2468 2468
rect 2412 2414 2414 2466
rect 2414 2414 2466 2466
rect 2466 2414 2468 2466
rect 2412 2412 2468 2414
rect 2572 2466 2628 2468
rect 2572 2414 2574 2466
rect 2574 2414 2626 2466
rect 2626 2414 2628 2466
rect 2572 2412 2628 2414
rect 2732 2466 2788 2468
rect 2732 2414 2734 2466
rect 2734 2414 2786 2466
rect 2786 2414 2788 2466
rect 2732 2412 2788 2414
rect 2892 2466 2948 2468
rect 2892 2414 2894 2466
rect 2894 2414 2946 2466
rect 2946 2414 2948 2466
rect 2892 2412 2948 2414
rect 3052 2466 3108 2468
rect 3052 2414 3054 2466
rect 3054 2414 3106 2466
rect 3106 2414 3108 2466
rect 3052 2412 3108 2414
rect 3372 2466 3428 2468
rect 3372 2414 3374 2466
rect 3374 2414 3426 2466
rect 3426 2414 3428 2466
rect 3372 2412 3428 2414
rect 3532 2466 3588 2468
rect 3532 2414 3534 2466
rect 3534 2414 3586 2466
rect 3586 2414 3588 2466
rect 3532 2412 3588 2414
rect 3692 2466 3748 2468
rect 3692 2414 3694 2466
rect 3694 2414 3746 2466
rect 3746 2414 3748 2466
rect 3692 2412 3748 2414
rect 3852 2466 3908 2468
rect 3852 2414 3854 2466
rect 3854 2414 3906 2466
rect 3906 2414 3908 2466
rect 3852 2412 3908 2414
rect 4012 2466 4068 2468
rect 4012 2414 4014 2466
rect 4014 2414 4066 2466
rect 4066 2414 4068 2466
rect 4012 2412 4068 2414
rect 4172 2466 4228 2468
rect 4172 2414 4174 2466
rect 4174 2414 4226 2466
rect 4226 2414 4228 2466
rect 4172 2412 4228 2414
rect 4332 2466 4388 2468
rect 4332 2414 4334 2466
rect 4334 2414 4386 2466
rect 4386 2414 4388 2466
rect 4332 2412 4388 2414
rect 4492 2466 4548 2468
rect 4492 2414 4494 2466
rect 4494 2414 4546 2466
rect 4546 2414 4548 2466
rect 4492 2412 4548 2414
rect 4652 2466 4708 2468
rect 4652 2414 4654 2466
rect 4654 2414 4706 2466
rect 4706 2414 4708 2466
rect 4652 2412 4708 2414
rect 4812 2466 4868 2468
rect 4812 2414 4814 2466
rect 4814 2414 4866 2466
rect 4866 2414 4868 2466
rect 4812 2412 4868 2414
rect 4972 2466 5028 2468
rect 4972 2414 4974 2466
rect 4974 2414 5026 2466
rect 5026 2414 5028 2466
rect 4972 2412 5028 2414
rect 5292 2466 5348 2468
rect 5292 2414 5294 2466
rect 5294 2414 5346 2466
rect 5346 2414 5348 2466
rect 5292 2412 5348 2414
rect 5452 2466 5508 2468
rect 5452 2414 5454 2466
rect 5454 2414 5506 2466
rect 5506 2414 5508 2466
rect 5452 2412 5508 2414
rect 5612 2466 5668 2468
rect 5612 2414 5614 2466
rect 5614 2414 5666 2466
rect 5666 2414 5668 2466
rect 5612 2412 5668 2414
rect 5772 2466 5828 2468
rect 5772 2414 5774 2466
rect 5774 2414 5826 2466
rect 5826 2414 5828 2466
rect 5772 2412 5828 2414
rect 5932 2466 5988 2468
rect 5932 2414 5934 2466
rect 5934 2414 5986 2466
rect 5986 2414 5988 2466
rect 5932 2412 5988 2414
rect 6092 2466 6148 2468
rect 6092 2414 6094 2466
rect 6094 2414 6146 2466
rect 6146 2414 6148 2466
rect 6092 2412 6148 2414
rect 6252 2466 6308 2468
rect 6252 2414 6254 2466
rect 6254 2414 6306 2466
rect 6306 2414 6308 2466
rect 6252 2412 6308 2414
rect 6412 2466 6468 2468
rect 6412 2414 6414 2466
rect 6414 2414 6466 2466
rect 6466 2414 6468 2466
rect 6412 2412 6468 2414
rect 6572 2466 6628 2468
rect 6572 2414 6574 2466
rect 6574 2414 6626 2466
rect 6626 2414 6628 2466
rect 6572 2412 6628 2414
rect 6732 2466 6788 2468
rect 6732 2414 6734 2466
rect 6734 2414 6786 2466
rect 6786 2414 6788 2466
rect 6732 2412 6788 2414
rect 6892 2466 6948 2468
rect 6892 2414 6894 2466
rect 6894 2414 6946 2466
rect 6946 2414 6948 2466
rect 6892 2412 6948 2414
rect 7212 2466 7268 2468
rect 7212 2414 7214 2466
rect 7214 2414 7266 2466
rect 7266 2414 7268 2466
rect 7212 2412 7268 2414
rect 7372 2466 7428 2468
rect 7372 2414 7374 2466
rect 7374 2414 7426 2466
rect 7426 2414 7428 2466
rect 7372 2412 7428 2414
rect 7532 2466 7588 2468
rect 7532 2414 7534 2466
rect 7534 2414 7586 2466
rect 7586 2414 7588 2466
rect 7532 2412 7588 2414
rect 7692 2466 7748 2468
rect 7692 2414 7694 2466
rect 7694 2414 7746 2466
rect 7746 2414 7748 2466
rect 7692 2412 7748 2414
rect 7852 2466 7908 2468
rect 7852 2414 7854 2466
rect 7854 2414 7906 2466
rect 7906 2414 7908 2466
rect 7852 2412 7908 2414
rect 8012 2466 8068 2468
rect 8012 2414 8014 2466
rect 8014 2414 8066 2466
rect 8066 2414 8068 2466
rect 8012 2412 8068 2414
rect 8172 2466 8228 2468
rect 8172 2414 8174 2466
rect 8174 2414 8226 2466
rect 8226 2414 8228 2466
rect 8172 2412 8228 2414
rect 8332 2466 8388 2468
rect 8332 2414 8334 2466
rect 8334 2414 8386 2466
rect 8386 2414 8388 2466
rect 8332 2412 8388 2414
rect 172 1212 228 1268
rect 332 1212 388 1268
rect 492 1212 548 1268
rect 652 1212 708 1268
rect 812 1212 868 1268
rect 972 1212 1028 1268
rect 1132 1212 1188 1268
rect 1452 1212 1508 1268
rect 1612 1212 1668 1268
rect 1772 1212 1828 1268
rect 1932 1212 1988 1268
rect 2092 1212 2148 1268
rect 2252 1212 2308 1268
rect 2412 1212 2468 1268
rect 2572 1212 2628 1268
rect 2732 1212 2788 1268
rect 2892 1212 2948 1268
rect 3052 1212 3108 1268
rect 3372 1212 3428 1268
rect 3532 1212 3588 1268
rect 3692 1212 3748 1268
rect 3852 1212 3908 1268
rect 4012 1212 4068 1268
rect 4172 1212 4228 1268
rect 4332 1212 4388 1268
rect 4492 1212 4548 1268
rect 4652 1212 4708 1268
rect 4812 1212 4868 1268
rect 4972 1212 5028 1268
rect 5292 1212 5348 1268
rect 5452 1212 5508 1268
rect 5612 1212 5668 1268
rect 5772 1212 5828 1268
rect 5932 1212 5988 1268
rect 6092 1212 6148 1268
rect 6252 1212 6308 1268
rect 6412 1212 6468 1268
rect 6572 1212 6628 1268
rect 6732 1212 6788 1268
rect 6892 1212 6948 1268
rect 7212 1212 7268 1268
rect 7372 1212 7428 1268
rect 7532 1212 7588 1268
rect 7692 1212 7748 1268
rect 7852 1212 7908 1268
rect 8012 1212 8068 1268
rect 8172 1212 8228 1268
rect 172 946 228 948
rect 172 894 174 946
rect 174 894 226 946
rect 226 894 228 946
rect 172 892 228 894
rect 332 892 388 948
rect 492 892 548 948
rect 652 892 708 948
rect 812 892 868 948
rect 972 892 1028 948
rect 1132 892 1188 948
rect 1452 892 1508 948
rect 1612 892 1668 948
rect 1772 892 1828 948
rect 1932 892 1988 948
rect 2092 892 2148 948
rect 2252 892 2308 948
rect 2412 892 2468 948
rect 2572 892 2628 948
rect 2732 892 2788 948
rect 2892 892 2948 948
rect 3052 892 3108 948
rect 3372 892 3428 948
rect 3532 892 3588 948
rect 3692 892 3748 948
rect 3852 892 3908 948
rect 4012 892 4068 948
rect 4172 892 4228 948
rect 4332 892 4388 948
rect 4492 892 4548 948
rect 4652 892 4708 948
rect 4812 892 4868 948
rect 4972 892 5028 948
rect 5292 892 5348 948
rect 5452 892 5508 948
rect 5612 892 5668 948
rect 5772 892 5828 948
rect 5932 892 5988 948
rect 6092 892 6148 948
rect 6252 892 6308 948
rect 6412 892 6468 948
rect 6572 892 6628 948
rect 6732 892 6788 948
rect 6892 892 6948 948
rect 7212 892 7268 948
rect 7372 892 7428 948
rect 7532 892 7588 948
rect 7692 892 7748 948
rect 7852 892 7908 948
rect 8172 892 8228 948
rect 172 572 228 628
rect 332 572 388 628
rect 492 572 548 628
rect 652 572 708 628
rect 812 572 868 628
rect 972 572 1028 628
rect 1132 572 1188 628
rect 1452 572 1508 628
rect 1612 572 1668 628
rect 1772 572 1828 628
rect 1932 572 1988 628
rect 2092 572 2148 628
rect 2252 572 2308 628
rect 2412 572 2468 628
rect 2572 572 2628 628
rect 2732 572 2788 628
rect 2892 572 2948 628
rect 3052 572 3108 628
rect 3372 572 3428 628
rect 3532 572 3588 628
rect 3692 572 3748 628
rect 3852 572 3908 628
rect 4012 572 4068 628
rect 4172 572 4228 628
rect 4332 572 4388 628
rect 4492 572 4548 628
rect 4652 572 4708 628
rect 4812 572 4868 628
rect 4972 572 5028 628
rect 5292 572 5348 628
rect 5452 572 5508 628
rect 5612 572 5668 628
rect 5772 572 5828 628
rect 5932 572 5988 628
rect 6092 572 6148 628
rect 6252 572 6308 628
rect 6412 572 6468 628
rect 6572 572 6628 628
rect 6732 572 6788 628
rect 6892 572 6948 628
rect 7212 572 7268 628
rect 7372 572 7428 628
rect 7532 572 7588 628
rect 7692 572 7748 628
rect 7852 572 7908 628
rect 8012 572 8068 628
rect 8172 572 8228 628
rect 332 318 388 328
rect 332 272 334 318
rect 334 272 386 318
rect 386 272 388 318
rect 332 202 334 248
rect 334 202 386 248
rect 386 202 388 248
rect 332 192 388 202
rect 172 -94 228 -92
rect 172 -146 174 -94
rect 174 -146 226 -94
rect 226 -146 228 -94
rect 172 -148 228 -146
rect 332 -94 388 -92
rect 332 -146 334 -94
rect 334 -146 386 -94
rect 386 -146 388 -94
rect 332 -148 388 -146
rect 492 -94 548 -92
rect 492 -146 494 -94
rect 494 -146 546 -94
rect 546 -146 548 -94
rect 492 -148 548 -146
rect 652 -94 708 -92
rect 652 -146 654 -94
rect 654 -146 706 -94
rect 706 -146 708 -94
rect 652 -148 708 -146
rect 812 -94 868 -92
rect 812 -146 814 -94
rect 814 -146 866 -94
rect 866 -146 868 -94
rect 812 -148 868 -146
rect 972 -94 1028 -92
rect 972 -146 974 -94
rect 974 -146 1026 -94
rect 1026 -146 1028 -94
rect 972 -148 1028 -146
rect 1132 -94 1188 -92
rect 1132 -146 1134 -94
rect 1134 -146 1186 -94
rect 1186 -146 1188 -94
rect 1132 -148 1188 -146
rect 1452 -94 1508 -92
rect 1452 -146 1454 -94
rect 1454 -146 1506 -94
rect 1506 -146 1508 -94
rect 1452 -148 1508 -146
rect 1612 -94 1668 -92
rect 1612 -146 1614 -94
rect 1614 -146 1666 -94
rect 1666 -146 1668 -94
rect 1612 -148 1668 -146
rect 1772 -94 1828 -92
rect 1772 -146 1774 -94
rect 1774 -146 1826 -94
rect 1826 -146 1828 -94
rect 1772 -148 1828 -146
rect 1932 -94 1988 -92
rect 1932 -146 1934 -94
rect 1934 -146 1986 -94
rect 1986 -146 1988 -94
rect 1932 -148 1988 -146
rect 2092 -94 2148 -92
rect 2092 -146 2094 -94
rect 2094 -146 2146 -94
rect 2146 -146 2148 -94
rect 2092 -148 2148 -146
rect 2252 -94 2308 -92
rect 2252 -146 2254 -94
rect 2254 -146 2306 -94
rect 2306 -146 2308 -94
rect 2252 -148 2308 -146
rect 2412 -94 2468 -92
rect 2412 -146 2414 -94
rect 2414 -146 2466 -94
rect 2466 -146 2468 -94
rect 2412 -148 2468 -146
rect 2572 -94 2628 -92
rect 2572 -146 2574 -94
rect 2574 -146 2626 -94
rect 2626 -146 2628 -94
rect 2572 -148 2628 -146
rect 2732 -94 2788 -92
rect 2732 -146 2734 -94
rect 2734 -146 2786 -94
rect 2786 -146 2788 -94
rect 2732 -148 2788 -146
rect 2892 -94 2948 -92
rect 2892 -146 2894 -94
rect 2894 -146 2946 -94
rect 2946 -146 2948 -94
rect 2892 -148 2948 -146
rect 3052 -94 3108 -92
rect 3052 -146 3054 -94
rect 3054 -146 3106 -94
rect 3106 -146 3108 -94
rect 3052 -148 3108 -146
rect 3372 -94 3428 -92
rect 3372 -146 3374 -94
rect 3374 -146 3426 -94
rect 3426 -146 3428 -94
rect 3372 -148 3428 -146
rect 3532 -94 3588 -92
rect 3532 -146 3534 -94
rect 3534 -146 3586 -94
rect 3586 -146 3588 -94
rect 3532 -148 3588 -146
rect 3692 -94 3748 -92
rect 3692 -146 3694 -94
rect 3694 -146 3746 -94
rect 3746 -146 3748 -94
rect 3692 -148 3748 -146
rect 3852 -94 3908 -92
rect 3852 -146 3854 -94
rect 3854 -146 3906 -94
rect 3906 -146 3908 -94
rect 3852 -148 3908 -146
rect 4012 -94 4068 -92
rect 4012 -146 4014 -94
rect 4014 -146 4066 -94
rect 4066 -146 4068 -94
rect 4012 -148 4068 -146
rect 4172 -94 4228 -92
rect 4172 -146 4174 -94
rect 4174 -146 4226 -94
rect 4226 -146 4228 -94
rect 4172 -148 4228 -146
rect 4332 -94 4388 -92
rect 4332 -146 4334 -94
rect 4334 -146 4386 -94
rect 4386 -146 4388 -94
rect 4332 -148 4388 -146
rect 4492 -94 4548 -92
rect 4492 -146 4494 -94
rect 4494 -146 4546 -94
rect 4546 -146 4548 -94
rect 4492 -148 4548 -146
rect 4652 -94 4708 -92
rect 4652 -146 4654 -94
rect 4654 -146 4706 -94
rect 4706 -146 4708 -94
rect 4652 -148 4708 -146
rect 4812 -94 4868 -92
rect 4812 -146 4814 -94
rect 4814 -146 4866 -94
rect 4866 -146 4868 -94
rect 4812 -148 4868 -146
rect 4972 -94 5028 -92
rect 4972 -146 4974 -94
rect 4974 -146 5026 -94
rect 5026 -146 5028 -94
rect 4972 -148 5028 -146
rect 5292 -94 5348 -92
rect 5292 -146 5294 -94
rect 5294 -146 5346 -94
rect 5346 -146 5348 -94
rect 5292 -148 5348 -146
rect 5452 -94 5508 -92
rect 5452 -146 5454 -94
rect 5454 -146 5506 -94
rect 5506 -146 5508 -94
rect 5452 -148 5508 -146
rect 5612 -94 5668 -92
rect 5612 -146 5614 -94
rect 5614 -146 5666 -94
rect 5666 -146 5668 -94
rect 5612 -148 5668 -146
rect 5772 -94 5828 -92
rect 5772 -146 5774 -94
rect 5774 -146 5826 -94
rect 5826 -146 5828 -94
rect 5772 -148 5828 -146
rect 5932 -94 5988 -92
rect 5932 -146 5934 -94
rect 5934 -146 5986 -94
rect 5986 -146 5988 -94
rect 5932 -148 5988 -146
rect 6092 -94 6148 -92
rect 6092 -146 6094 -94
rect 6094 -146 6146 -94
rect 6146 -146 6148 -94
rect 6092 -148 6148 -146
rect 6252 -94 6308 -92
rect 6252 -146 6254 -94
rect 6254 -146 6306 -94
rect 6306 -146 6308 -94
rect 6252 -148 6308 -146
rect 6412 -94 6468 -92
rect 6412 -146 6414 -94
rect 6414 -146 6466 -94
rect 6466 -146 6468 -94
rect 6412 -148 6468 -146
rect 6572 -94 6628 -92
rect 6572 -146 6574 -94
rect 6574 -146 6626 -94
rect 6626 -146 6628 -94
rect 6572 -148 6628 -146
rect 6732 -94 6788 -92
rect 6732 -146 6734 -94
rect 6734 -146 6786 -94
rect 6786 -146 6788 -94
rect 6732 -148 6788 -146
rect 6892 -94 6948 -92
rect 6892 -146 6894 -94
rect 6894 -146 6946 -94
rect 6946 -146 6948 -94
rect 6892 -148 6948 -146
rect 7212 -94 7268 -92
rect 7212 -146 7214 -94
rect 7214 -146 7266 -94
rect 7266 -146 7268 -94
rect 7212 -148 7268 -146
rect 7372 -94 7428 -92
rect 7372 -146 7374 -94
rect 7374 -146 7426 -94
rect 7426 -146 7428 -94
rect 7372 -148 7428 -146
rect 7532 -94 7588 -92
rect 7532 -146 7534 -94
rect 7534 -146 7586 -94
rect 7586 -146 7588 -94
rect 7532 -148 7588 -146
rect 7692 -94 7748 -92
rect 7692 -146 7694 -94
rect 7694 -146 7746 -94
rect 7746 -146 7748 -94
rect 7692 -148 7748 -146
rect 7852 -94 7908 -92
rect 7852 -146 7854 -94
rect 7854 -146 7906 -94
rect 7906 -146 7908 -94
rect 7852 -148 7908 -146
rect 8172 -94 8228 -92
rect 8172 -146 8174 -94
rect 8174 -146 8226 -94
rect 8226 -146 8228 -94
rect 8172 -148 8228 -146
rect 172 -468 228 -412
rect 332 -468 388 -412
rect 492 -468 548 -412
rect 652 -468 708 -412
rect 812 -468 868 -412
rect 972 -468 1028 -412
rect 1132 -468 1188 -412
rect 1452 -468 1508 -412
rect 1612 -468 1668 -412
rect 1772 -468 1828 -412
rect 1932 -468 1988 -412
rect 2092 -468 2148 -412
rect 2252 -468 2308 -412
rect 2412 -468 2468 -412
rect 2572 -468 2628 -412
rect 2732 -468 2788 -412
rect 2892 -468 2948 -412
rect 3052 -468 3108 -412
rect 3372 -468 3428 -412
rect 3532 -468 3588 -412
rect 3692 -468 3748 -412
rect 3852 -468 3908 -412
rect 4012 -468 4068 -412
rect 4172 -468 4228 -412
rect 4332 -468 4388 -412
rect 4492 -468 4548 -412
rect 4652 -468 4708 -412
rect 4812 -468 4868 -412
rect 4972 -468 5028 -412
rect 5292 -468 5348 -412
rect 5452 -468 5508 -412
rect 5612 -468 5668 -412
rect 5772 -468 5828 -412
rect 5932 -468 5988 -412
rect 6092 -468 6148 -412
rect 6252 -468 6308 -412
rect 6412 -468 6468 -412
rect 6572 -468 6628 -412
rect 6732 -468 6788 -412
rect 6892 -468 6948 -412
rect 7212 -468 7268 -412
rect 7372 -468 7428 -412
rect 7532 -468 7588 -412
rect 7692 -468 7748 -412
rect 7852 -468 7908 -412
rect 8172 -468 8228 -412
rect 332 -722 388 -712
rect 332 -768 334 -722
rect 334 -768 386 -722
rect 386 -768 388 -722
rect 332 -838 334 -792
rect 334 -838 386 -792
rect 386 -838 388 -792
rect 332 -848 388 -838
<< metal3 >>
rect 320 9712 400 9760
rect 320 9648 328 9712
rect 392 9648 400 9712
rect 320 9632 400 9648
rect 320 9568 328 9632
rect 392 9568 400 9632
rect 320 9552 400 9568
rect 320 9488 328 9552
rect 392 9488 400 9552
rect 320 9472 400 9488
rect 320 9408 328 9472
rect 392 9408 400 9472
rect 320 9360 400 9408
rect 160 8792 240 8800
rect 160 8728 168 8792
rect 232 8728 240 8792
rect 160 8632 240 8728
rect 160 8568 168 8632
rect 232 8568 240 8632
rect 160 8472 240 8568
rect 160 8408 168 8472
rect 232 8408 240 8472
rect 160 8400 240 8408
rect 320 8792 400 8800
rect 320 8728 328 8792
rect 392 8728 400 8792
rect 320 8632 400 8728
rect 320 8568 328 8632
rect 392 8568 400 8632
rect 320 8472 400 8568
rect 320 8408 328 8472
rect 392 8408 400 8472
rect 320 8400 400 8408
rect 480 8792 560 8800
rect 480 8728 488 8792
rect 552 8728 560 8792
rect 480 8632 560 8728
rect 480 8568 488 8632
rect 552 8568 560 8632
rect 480 8472 560 8568
rect 480 8408 488 8472
rect 552 8408 560 8472
rect 480 8400 560 8408
rect 640 8792 720 8800
rect 640 8728 648 8792
rect 712 8728 720 8792
rect 640 8632 720 8728
rect 640 8568 648 8632
rect 712 8568 720 8632
rect 640 8472 720 8568
rect 640 8408 648 8472
rect 712 8408 720 8472
rect 640 8400 720 8408
rect 800 8792 880 8800
rect 800 8728 808 8792
rect 872 8728 880 8792
rect 800 8632 880 8728
rect 800 8568 808 8632
rect 872 8568 880 8632
rect 800 8472 880 8568
rect 800 8408 808 8472
rect 872 8408 880 8472
rect 800 8400 880 8408
rect 960 8792 1040 8800
rect 960 8728 968 8792
rect 1032 8728 1040 8792
rect 960 8632 1040 8728
rect 960 8568 968 8632
rect 1032 8568 1040 8632
rect 960 8472 1040 8568
rect 960 8408 968 8472
rect 1032 8408 1040 8472
rect 960 8400 1040 8408
rect 1120 8792 1200 8800
rect 1120 8728 1128 8792
rect 1192 8728 1200 8792
rect 1120 8632 1200 8728
rect 1120 8568 1128 8632
rect 1192 8568 1200 8632
rect 1120 8472 1200 8568
rect 1120 8408 1128 8472
rect 1192 8408 1200 8472
rect 1120 8400 1200 8408
rect 1440 8792 1520 8800
rect 1440 8728 1448 8792
rect 1512 8728 1520 8792
rect 1440 8632 1520 8728
rect 1440 8568 1448 8632
rect 1512 8568 1520 8632
rect 1440 8472 1520 8568
rect 1440 8408 1448 8472
rect 1512 8408 1520 8472
rect 1440 8400 1520 8408
rect 1600 8792 1680 8800
rect 1600 8728 1608 8792
rect 1672 8728 1680 8792
rect 1600 8632 1680 8728
rect 1600 8568 1608 8632
rect 1672 8568 1680 8632
rect 1600 8472 1680 8568
rect 1600 8408 1608 8472
rect 1672 8408 1680 8472
rect 1600 8400 1680 8408
rect 1760 8792 1840 8800
rect 1760 8728 1768 8792
rect 1832 8728 1840 8792
rect 1760 8632 1840 8728
rect 1760 8568 1768 8632
rect 1832 8568 1840 8632
rect 1760 8472 1840 8568
rect 1760 8408 1768 8472
rect 1832 8408 1840 8472
rect 1760 8400 1840 8408
rect 1920 8792 2000 8800
rect 1920 8728 1928 8792
rect 1992 8728 2000 8792
rect 1920 8632 2000 8728
rect 1920 8568 1928 8632
rect 1992 8568 2000 8632
rect 1920 8472 2000 8568
rect 1920 8408 1928 8472
rect 1992 8408 2000 8472
rect 1920 8400 2000 8408
rect 2080 8792 2160 8800
rect 2080 8728 2088 8792
rect 2152 8728 2160 8792
rect 2080 8632 2160 8728
rect 2080 8568 2088 8632
rect 2152 8568 2160 8632
rect 2080 8472 2160 8568
rect 2080 8408 2088 8472
rect 2152 8408 2160 8472
rect 2080 8400 2160 8408
rect 2240 8792 2320 8800
rect 2240 8728 2248 8792
rect 2312 8728 2320 8792
rect 2240 8632 2320 8728
rect 2240 8568 2248 8632
rect 2312 8568 2320 8632
rect 2240 8472 2320 8568
rect 2240 8408 2248 8472
rect 2312 8408 2320 8472
rect 2240 8400 2320 8408
rect 2400 8792 2480 8800
rect 2400 8728 2408 8792
rect 2472 8728 2480 8792
rect 2400 8632 2480 8728
rect 2400 8568 2408 8632
rect 2472 8568 2480 8632
rect 2400 8472 2480 8568
rect 2400 8408 2408 8472
rect 2472 8408 2480 8472
rect 2400 8400 2480 8408
rect 2560 8792 2640 8800
rect 2560 8728 2568 8792
rect 2632 8728 2640 8792
rect 2560 8632 2640 8728
rect 2560 8568 2568 8632
rect 2632 8568 2640 8632
rect 2560 8472 2640 8568
rect 2560 8408 2568 8472
rect 2632 8408 2640 8472
rect 2560 8400 2640 8408
rect 2720 8792 2800 8800
rect 2720 8728 2728 8792
rect 2792 8728 2800 8792
rect 2720 8632 2800 8728
rect 2720 8568 2728 8632
rect 2792 8568 2800 8632
rect 2720 8472 2800 8568
rect 2720 8408 2728 8472
rect 2792 8408 2800 8472
rect 2720 8400 2800 8408
rect 2880 8792 2960 8800
rect 2880 8728 2888 8792
rect 2952 8728 2960 8792
rect 2880 8632 2960 8728
rect 2880 8568 2888 8632
rect 2952 8568 2960 8632
rect 2880 8472 2960 8568
rect 2880 8408 2888 8472
rect 2952 8408 2960 8472
rect 2880 8400 2960 8408
rect 3040 8792 3120 8800
rect 3040 8728 3048 8792
rect 3112 8728 3120 8792
rect 3040 8632 3120 8728
rect 3040 8568 3048 8632
rect 3112 8568 3120 8632
rect 3040 8472 3120 8568
rect 3040 8408 3048 8472
rect 3112 8408 3120 8472
rect 3040 8400 3120 8408
rect 3360 8792 3440 8800
rect 3360 8728 3368 8792
rect 3432 8728 3440 8792
rect 3360 8632 3440 8728
rect 3360 8568 3368 8632
rect 3432 8568 3440 8632
rect 3360 8472 3440 8568
rect 3360 8408 3368 8472
rect 3432 8408 3440 8472
rect 3360 8400 3440 8408
rect 3520 8792 3600 8800
rect 3520 8728 3528 8792
rect 3592 8728 3600 8792
rect 3520 8632 3600 8728
rect 3520 8568 3528 8632
rect 3592 8568 3600 8632
rect 3520 8472 3600 8568
rect 3520 8408 3528 8472
rect 3592 8408 3600 8472
rect 3520 8400 3600 8408
rect 3680 8792 3760 8800
rect 3680 8728 3688 8792
rect 3752 8728 3760 8792
rect 3680 8632 3760 8728
rect 3680 8568 3688 8632
rect 3752 8568 3760 8632
rect 3680 8472 3760 8568
rect 3680 8408 3688 8472
rect 3752 8408 3760 8472
rect 3680 8400 3760 8408
rect 3840 8792 3920 8800
rect 3840 8728 3848 8792
rect 3912 8728 3920 8792
rect 3840 8632 3920 8728
rect 3840 8568 3848 8632
rect 3912 8568 3920 8632
rect 3840 8472 3920 8568
rect 3840 8408 3848 8472
rect 3912 8408 3920 8472
rect 3840 8400 3920 8408
rect 4000 8792 4080 8800
rect 4000 8728 4008 8792
rect 4072 8728 4080 8792
rect 4000 8632 4080 8728
rect 4000 8568 4008 8632
rect 4072 8568 4080 8632
rect 4000 8472 4080 8568
rect 4000 8408 4008 8472
rect 4072 8408 4080 8472
rect 4000 8400 4080 8408
rect 4160 8792 4240 8800
rect 4160 8728 4168 8792
rect 4232 8728 4240 8792
rect 4160 8632 4240 8728
rect 4160 8568 4168 8632
rect 4232 8568 4240 8632
rect 4160 8472 4240 8568
rect 4160 8408 4168 8472
rect 4232 8408 4240 8472
rect 4160 8400 4240 8408
rect 4320 8792 4400 8800
rect 4320 8728 4328 8792
rect 4392 8728 4400 8792
rect 4320 8632 4400 8728
rect 4320 8568 4328 8632
rect 4392 8568 4400 8632
rect 4320 8472 4400 8568
rect 4320 8408 4328 8472
rect 4392 8408 4400 8472
rect 4320 8400 4400 8408
rect 4480 8792 4560 8800
rect 4480 8728 4488 8792
rect 4552 8728 4560 8792
rect 4480 8632 4560 8728
rect 4480 8568 4488 8632
rect 4552 8568 4560 8632
rect 4480 8472 4560 8568
rect 4480 8408 4488 8472
rect 4552 8408 4560 8472
rect 4480 8400 4560 8408
rect 4640 8792 4720 8800
rect 4640 8728 4648 8792
rect 4712 8728 4720 8792
rect 4640 8632 4720 8728
rect 4640 8568 4648 8632
rect 4712 8568 4720 8632
rect 4640 8472 4720 8568
rect 4640 8408 4648 8472
rect 4712 8408 4720 8472
rect 4640 8400 4720 8408
rect 4800 8792 4880 8800
rect 4800 8728 4808 8792
rect 4872 8728 4880 8792
rect 4800 8632 4880 8728
rect 4800 8568 4808 8632
rect 4872 8568 4880 8632
rect 4800 8472 4880 8568
rect 4800 8408 4808 8472
rect 4872 8408 4880 8472
rect 4800 8400 4880 8408
rect 4960 8792 5040 8800
rect 4960 8728 4968 8792
rect 5032 8728 5040 8792
rect 4960 8632 5040 8728
rect 4960 8568 4968 8632
rect 5032 8568 5040 8632
rect 4960 8472 5040 8568
rect 4960 8408 4968 8472
rect 5032 8408 5040 8472
rect 4960 8400 5040 8408
rect 5280 8792 5360 8800
rect 5280 8728 5288 8792
rect 5352 8728 5360 8792
rect 5280 8632 5360 8728
rect 5280 8568 5288 8632
rect 5352 8568 5360 8632
rect 5280 8472 5360 8568
rect 5280 8408 5288 8472
rect 5352 8408 5360 8472
rect 5280 8400 5360 8408
rect 5440 8792 5520 8800
rect 5440 8728 5448 8792
rect 5512 8728 5520 8792
rect 5440 8632 5520 8728
rect 5440 8568 5448 8632
rect 5512 8568 5520 8632
rect 5440 8472 5520 8568
rect 5440 8408 5448 8472
rect 5512 8408 5520 8472
rect 5440 8400 5520 8408
rect 5600 8792 5680 8800
rect 5600 8728 5608 8792
rect 5672 8728 5680 8792
rect 5600 8632 5680 8728
rect 5600 8568 5608 8632
rect 5672 8568 5680 8632
rect 5600 8472 5680 8568
rect 5600 8408 5608 8472
rect 5672 8408 5680 8472
rect 5600 8400 5680 8408
rect 5760 8792 5840 8800
rect 5760 8728 5768 8792
rect 5832 8728 5840 8792
rect 5760 8632 5840 8728
rect 5760 8568 5768 8632
rect 5832 8568 5840 8632
rect 5760 8472 5840 8568
rect 5760 8408 5768 8472
rect 5832 8408 5840 8472
rect 5760 8400 5840 8408
rect 5920 8792 6000 8800
rect 5920 8728 5928 8792
rect 5992 8728 6000 8792
rect 5920 8632 6000 8728
rect 5920 8568 5928 8632
rect 5992 8568 6000 8632
rect 5920 8472 6000 8568
rect 5920 8408 5928 8472
rect 5992 8408 6000 8472
rect 5920 8400 6000 8408
rect 6080 8792 6160 8800
rect 6080 8728 6088 8792
rect 6152 8728 6160 8792
rect 6080 8632 6160 8728
rect 6080 8568 6088 8632
rect 6152 8568 6160 8632
rect 6080 8472 6160 8568
rect 6080 8408 6088 8472
rect 6152 8408 6160 8472
rect 6080 8400 6160 8408
rect 6240 8792 6320 8800
rect 6240 8728 6248 8792
rect 6312 8728 6320 8792
rect 6240 8632 6320 8728
rect 6240 8568 6248 8632
rect 6312 8568 6320 8632
rect 6240 8472 6320 8568
rect 6240 8408 6248 8472
rect 6312 8408 6320 8472
rect 6240 8400 6320 8408
rect 6400 8792 6480 8800
rect 6400 8728 6408 8792
rect 6472 8728 6480 8792
rect 6400 8632 6480 8728
rect 6400 8568 6408 8632
rect 6472 8568 6480 8632
rect 6400 8472 6480 8568
rect 6400 8408 6408 8472
rect 6472 8408 6480 8472
rect 6400 8400 6480 8408
rect 6560 8792 6640 8800
rect 6560 8728 6568 8792
rect 6632 8728 6640 8792
rect 6560 8632 6640 8728
rect 6560 8568 6568 8632
rect 6632 8568 6640 8632
rect 6560 8472 6640 8568
rect 6560 8408 6568 8472
rect 6632 8408 6640 8472
rect 6560 8400 6640 8408
rect 6720 8792 6800 8800
rect 6720 8728 6728 8792
rect 6792 8728 6800 8792
rect 6720 8632 6800 8728
rect 6720 8568 6728 8632
rect 6792 8568 6800 8632
rect 6720 8472 6800 8568
rect 6720 8408 6728 8472
rect 6792 8408 6800 8472
rect 6720 8400 6800 8408
rect 6880 8792 6960 8800
rect 6880 8728 6888 8792
rect 6952 8728 6960 8792
rect 6880 8632 6960 8728
rect 6880 8568 6888 8632
rect 6952 8568 6960 8632
rect 6880 8472 6960 8568
rect 6880 8408 6888 8472
rect 6952 8408 6960 8472
rect 6880 8400 6960 8408
rect 7200 8792 7280 8800
rect 7200 8728 7208 8792
rect 7272 8728 7280 8792
rect 7200 8632 7280 8728
rect 7200 8568 7208 8632
rect 7272 8568 7280 8632
rect 7200 8472 7280 8568
rect 7200 8408 7208 8472
rect 7272 8408 7280 8472
rect 7200 8400 7280 8408
rect 7360 8792 7440 8800
rect 7360 8728 7368 8792
rect 7432 8728 7440 8792
rect 7360 8632 7440 8728
rect 7360 8568 7368 8632
rect 7432 8568 7440 8632
rect 7360 8472 7440 8568
rect 7360 8408 7368 8472
rect 7432 8408 7440 8472
rect 7360 8400 7440 8408
rect 7520 8792 7600 8800
rect 7520 8728 7528 8792
rect 7592 8728 7600 8792
rect 7520 8632 7600 8728
rect 7520 8568 7528 8632
rect 7592 8568 7600 8632
rect 7520 8472 7600 8568
rect 7520 8408 7528 8472
rect 7592 8408 7600 8472
rect 7520 8400 7600 8408
rect 7680 8792 7760 8800
rect 7680 8728 7688 8792
rect 7752 8728 7760 8792
rect 7680 8632 7760 8728
rect 7680 8568 7688 8632
rect 7752 8568 7760 8632
rect 7680 8472 7760 8568
rect 7680 8408 7688 8472
rect 7752 8408 7760 8472
rect 7680 8400 7760 8408
rect 7840 8792 7920 8800
rect 7840 8728 7848 8792
rect 7912 8728 7920 8792
rect 7840 8632 7920 8728
rect 7840 8568 7848 8632
rect 7912 8568 7920 8632
rect 7840 8472 7920 8568
rect 7840 8408 7848 8472
rect 7912 8408 7920 8472
rect 7840 8400 7920 8408
rect 8000 8792 8080 8800
rect 8000 8728 8008 8792
rect 8072 8728 8080 8792
rect 8000 8632 8080 8728
rect 8000 8568 8008 8632
rect 8072 8568 8080 8632
rect 8000 8472 8080 8568
rect 8000 8408 8008 8472
rect 8072 8408 8080 8472
rect 8000 8400 8080 8408
rect 8160 8792 8240 8800
rect 8160 8728 8168 8792
rect 8232 8728 8240 8792
rect 8160 8632 8240 8728
rect 8160 8568 8168 8632
rect 8232 8568 8240 8632
rect 8160 8472 8240 8568
rect 8160 8408 8168 8472
rect 8232 8408 8240 8472
rect 8160 8400 8240 8408
rect 160 8312 240 8320
rect 160 8248 168 8312
rect 232 8248 240 8312
rect 160 8152 240 8248
rect 160 8088 168 8152
rect 232 8088 240 8152
rect 160 7992 240 8088
rect 160 7928 168 7992
rect 232 7928 240 7992
rect 160 7920 240 7928
rect 320 8312 400 8320
rect 320 8248 328 8312
rect 392 8248 400 8312
rect 320 8152 400 8248
rect 320 8088 328 8152
rect 392 8088 400 8152
rect 320 7992 400 8088
rect 320 7928 328 7992
rect 392 7928 400 7992
rect 320 7920 400 7928
rect 480 8312 560 8320
rect 480 8248 488 8312
rect 552 8248 560 8312
rect 480 8152 560 8248
rect 480 8088 488 8152
rect 552 8088 560 8152
rect 480 7992 560 8088
rect 480 7928 488 7992
rect 552 7928 560 7992
rect 480 7920 560 7928
rect 640 8312 720 8320
rect 640 8248 648 8312
rect 712 8248 720 8312
rect 640 8152 720 8248
rect 640 8088 648 8152
rect 712 8088 720 8152
rect 640 7992 720 8088
rect 640 7928 648 7992
rect 712 7928 720 7992
rect 640 7920 720 7928
rect 800 8312 880 8320
rect 800 8248 808 8312
rect 872 8248 880 8312
rect 800 8152 880 8248
rect 800 8088 808 8152
rect 872 8088 880 8152
rect 800 7992 880 8088
rect 800 7928 808 7992
rect 872 7928 880 7992
rect 800 7920 880 7928
rect 960 8312 1040 8320
rect 960 8248 968 8312
rect 1032 8248 1040 8312
rect 960 8152 1040 8248
rect 960 8088 968 8152
rect 1032 8088 1040 8152
rect 960 7992 1040 8088
rect 960 7928 968 7992
rect 1032 7928 1040 7992
rect 960 7920 1040 7928
rect 1120 8312 1200 8320
rect 1120 8248 1128 8312
rect 1192 8248 1200 8312
rect 1120 8152 1200 8248
rect 1120 8088 1128 8152
rect 1192 8088 1200 8152
rect 1120 7992 1200 8088
rect 1120 7928 1128 7992
rect 1192 7928 1200 7992
rect 1120 7920 1200 7928
rect 1440 8312 1520 8320
rect 1440 8248 1448 8312
rect 1512 8248 1520 8312
rect 1440 8152 1520 8248
rect 1440 8088 1448 8152
rect 1512 8088 1520 8152
rect 1440 7992 1520 8088
rect 1440 7928 1448 7992
rect 1512 7928 1520 7992
rect 1440 7920 1520 7928
rect 1600 8312 1680 8320
rect 1600 8248 1608 8312
rect 1672 8248 1680 8312
rect 1600 8152 1680 8248
rect 1600 8088 1608 8152
rect 1672 8088 1680 8152
rect 1600 7992 1680 8088
rect 1600 7928 1608 7992
rect 1672 7928 1680 7992
rect 1600 7920 1680 7928
rect 1760 8312 1840 8320
rect 1760 8248 1768 8312
rect 1832 8248 1840 8312
rect 1760 8152 1840 8248
rect 1760 8088 1768 8152
rect 1832 8088 1840 8152
rect 1760 7992 1840 8088
rect 1760 7928 1768 7992
rect 1832 7928 1840 7992
rect 1760 7920 1840 7928
rect 1920 8312 2000 8320
rect 1920 8248 1928 8312
rect 1992 8248 2000 8312
rect 1920 8152 2000 8248
rect 1920 8088 1928 8152
rect 1992 8088 2000 8152
rect 1920 7992 2000 8088
rect 1920 7928 1928 7992
rect 1992 7928 2000 7992
rect 1920 7920 2000 7928
rect 2080 8312 2160 8320
rect 2080 8248 2088 8312
rect 2152 8248 2160 8312
rect 2080 8152 2160 8248
rect 2080 8088 2088 8152
rect 2152 8088 2160 8152
rect 2080 7992 2160 8088
rect 2080 7928 2088 7992
rect 2152 7928 2160 7992
rect 2080 7920 2160 7928
rect 2240 8312 2320 8320
rect 2240 8248 2248 8312
rect 2312 8248 2320 8312
rect 2240 8152 2320 8248
rect 2240 8088 2248 8152
rect 2312 8088 2320 8152
rect 2240 7992 2320 8088
rect 2240 7928 2248 7992
rect 2312 7928 2320 7992
rect 2240 7920 2320 7928
rect 2400 8312 2480 8320
rect 2400 8248 2408 8312
rect 2472 8248 2480 8312
rect 2400 8152 2480 8248
rect 2400 8088 2408 8152
rect 2472 8088 2480 8152
rect 2400 7992 2480 8088
rect 2400 7928 2408 7992
rect 2472 7928 2480 7992
rect 2400 7920 2480 7928
rect 2560 8312 2640 8320
rect 2560 8248 2568 8312
rect 2632 8248 2640 8312
rect 2560 8152 2640 8248
rect 2560 8088 2568 8152
rect 2632 8088 2640 8152
rect 2560 7992 2640 8088
rect 2560 7928 2568 7992
rect 2632 7928 2640 7992
rect 2560 7920 2640 7928
rect 2720 8312 2800 8320
rect 2720 8248 2728 8312
rect 2792 8248 2800 8312
rect 2720 8152 2800 8248
rect 2720 8088 2728 8152
rect 2792 8088 2800 8152
rect 2720 7992 2800 8088
rect 2720 7928 2728 7992
rect 2792 7928 2800 7992
rect 2720 7920 2800 7928
rect 2880 8312 2960 8320
rect 2880 8248 2888 8312
rect 2952 8248 2960 8312
rect 2880 8152 2960 8248
rect 2880 8088 2888 8152
rect 2952 8088 2960 8152
rect 2880 7992 2960 8088
rect 2880 7928 2888 7992
rect 2952 7928 2960 7992
rect 2880 7920 2960 7928
rect 3040 8312 3120 8320
rect 3040 8248 3048 8312
rect 3112 8248 3120 8312
rect 3040 8152 3120 8248
rect 3040 8088 3048 8152
rect 3112 8088 3120 8152
rect 3040 7992 3120 8088
rect 3040 7928 3048 7992
rect 3112 7928 3120 7992
rect 3040 7920 3120 7928
rect 3360 8312 3440 8320
rect 3360 8248 3368 8312
rect 3432 8248 3440 8312
rect 3360 8152 3440 8248
rect 3360 8088 3368 8152
rect 3432 8088 3440 8152
rect 3360 7992 3440 8088
rect 3360 7928 3368 7992
rect 3432 7928 3440 7992
rect 3360 7920 3440 7928
rect 3520 8312 3600 8320
rect 3520 8248 3528 8312
rect 3592 8248 3600 8312
rect 3520 8152 3600 8248
rect 3520 8088 3528 8152
rect 3592 8088 3600 8152
rect 3520 7992 3600 8088
rect 3520 7928 3528 7992
rect 3592 7928 3600 7992
rect 3520 7920 3600 7928
rect 3680 8312 3760 8320
rect 3680 8248 3688 8312
rect 3752 8248 3760 8312
rect 3680 8152 3760 8248
rect 3680 8088 3688 8152
rect 3752 8088 3760 8152
rect 3680 7992 3760 8088
rect 3680 7928 3688 7992
rect 3752 7928 3760 7992
rect 3680 7920 3760 7928
rect 3840 8312 3920 8320
rect 3840 8248 3848 8312
rect 3912 8248 3920 8312
rect 3840 8152 3920 8248
rect 3840 8088 3848 8152
rect 3912 8088 3920 8152
rect 3840 7992 3920 8088
rect 3840 7928 3848 7992
rect 3912 7928 3920 7992
rect 3840 7920 3920 7928
rect 4000 8312 4080 8320
rect 4000 8248 4008 8312
rect 4072 8248 4080 8312
rect 4000 8152 4080 8248
rect 4000 8088 4008 8152
rect 4072 8088 4080 8152
rect 4000 7992 4080 8088
rect 4000 7928 4008 7992
rect 4072 7928 4080 7992
rect 4000 7920 4080 7928
rect 4160 8312 4240 8320
rect 4160 8248 4168 8312
rect 4232 8248 4240 8312
rect 4160 8152 4240 8248
rect 4160 8088 4168 8152
rect 4232 8088 4240 8152
rect 4160 7992 4240 8088
rect 4160 7928 4168 7992
rect 4232 7928 4240 7992
rect 4160 7920 4240 7928
rect 4320 8312 4400 8320
rect 4320 8248 4328 8312
rect 4392 8248 4400 8312
rect 4320 8152 4400 8248
rect 4320 8088 4328 8152
rect 4392 8088 4400 8152
rect 4320 7992 4400 8088
rect 4320 7928 4328 7992
rect 4392 7928 4400 7992
rect 4320 7920 4400 7928
rect 4480 8312 4560 8320
rect 4480 8248 4488 8312
rect 4552 8248 4560 8312
rect 4480 8152 4560 8248
rect 4480 8088 4488 8152
rect 4552 8088 4560 8152
rect 4480 7992 4560 8088
rect 4480 7928 4488 7992
rect 4552 7928 4560 7992
rect 4480 7920 4560 7928
rect 4640 8312 4720 8320
rect 4640 8248 4648 8312
rect 4712 8248 4720 8312
rect 4640 8152 4720 8248
rect 4640 8088 4648 8152
rect 4712 8088 4720 8152
rect 4640 7992 4720 8088
rect 4640 7928 4648 7992
rect 4712 7928 4720 7992
rect 4640 7920 4720 7928
rect 4800 8312 4880 8320
rect 4800 8248 4808 8312
rect 4872 8248 4880 8312
rect 4800 8152 4880 8248
rect 4800 8088 4808 8152
rect 4872 8088 4880 8152
rect 4800 7992 4880 8088
rect 4800 7928 4808 7992
rect 4872 7928 4880 7992
rect 4800 7920 4880 7928
rect 4960 8312 5040 8320
rect 4960 8248 4968 8312
rect 5032 8248 5040 8312
rect 4960 8152 5040 8248
rect 4960 8088 4968 8152
rect 5032 8088 5040 8152
rect 4960 7992 5040 8088
rect 4960 7928 4968 7992
rect 5032 7928 5040 7992
rect 4960 7920 5040 7928
rect 5280 8312 5360 8320
rect 5280 8248 5288 8312
rect 5352 8248 5360 8312
rect 5280 8152 5360 8248
rect 5280 8088 5288 8152
rect 5352 8088 5360 8152
rect 5280 7992 5360 8088
rect 5280 7928 5288 7992
rect 5352 7928 5360 7992
rect 5280 7920 5360 7928
rect 5440 8312 5520 8320
rect 5440 8248 5448 8312
rect 5512 8248 5520 8312
rect 5440 8152 5520 8248
rect 5440 8088 5448 8152
rect 5512 8088 5520 8152
rect 5440 7992 5520 8088
rect 5440 7928 5448 7992
rect 5512 7928 5520 7992
rect 5440 7920 5520 7928
rect 5600 8312 5680 8320
rect 5600 8248 5608 8312
rect 5672 8248 5680 8312
rect 5600 8152 5680 8248
rect 5600 8088 5608 8152
rect 5672 8088 5680 8152
rect 5600 7992 5680 8088
rect 5600 7928 5608 7992
rect 5672 7928 5680 7992
rect 5600 7920 5680 7928
rect 5760 8312 5840 8320
rect 5760 8248 5768 8312
rect 5832 8248 5840 8312
rect 5760 8152 5840 8248
rect 5760 8088 5768 8152
rect 5832 8088 5840 8152
rect 5760 7992 5840 8088
rect 5760 7928 5768 7992
rect 5832 7928 5840 7992
rect 5760 7920 5840 7928
rect 5920 8312 6000 8320
rect 5920 8248 5928 8312
rect 5992 8248 6000 8312
rect 5920 8152 6000 8248
rect 5920 8088 5928 8152
rect 5992 8088 6000 8152
rect 5920 7992 6000 8088
rect 5920 7928 5928 7992
rect 5992 7928 6000 7992
rect 5920 7920 6000 7928
rect 6080 8312 6160 8320
rect 6080 8248 6088 8312
rect 6152 8248 6160 8312
rect 6080 8152 6160 8248
rect 6080 8088 6088 8152
rect 6152 8088 6160 8152
rect 6080 7992 6160 8088
rect 6080 7928 6088 7992
rect 6152 7928 6160 7992
rect 6080 7920 6160 7928
rect 6240 8312 6320 8320
rect 6240 8248 6248 8312
rect 6312 8248 6320 8312
rect 6240 8152 6320 8248
rect 6240 8088 6248 8152
rect 6312 8088 6320 8152
rect 6240 7992 6320 8088
rect 6240 7928 6248 7992
rect 6312 7928 6320 7992
rect 6240 7920 6320 7928
rect 6400 8312 6480 8320
rect 6400 8248 6408 8312
rect 6472 8248 6480 8312
rect 6400 8152 6480 8248
rect 6400 8088 6408 8152
rect 6472 8088 6480 8152
rect 6400 7992 6480 8088
rect 6400 7928 6408 7992
rect 6472 7928 6480 7992
rect 6400 7920 6480 7928
rect 6560 8312 6640 8320
rect 6560 8248 6568 8312
rect 6632 8248 6640 8312
rect 6560 8152 6640 8248
rect 6560 8088 6568 8152
rect 6632 8088 6640 8152
rect 6560 7992 6640 8088
rect 6560 7928 6568 7992
rect 6632 7928 6640 7992
rect 6560 7920 6640 7928
rect 6720 8312 6800 8320
rect 6720 8248 6728 8312
rect 6792 8248 6800 8312
rect 6720 8152 6800 8248
rect 6720 8088 6728 8152
rect 6792 8088 6800 8152
rect 6720 7992 6800 8088
rect 6720 7928 6728 7992
rect 6792 7928 6800 7992
rect 6720 7920 6800 7928
rect 6880 8312 6960 8320
rect 6880 8248 6888 8312
rect 6952 8248 6960 8312
rect 6880 8152 6960 8248
rect 6880 8088 6888 8152
rect 6952 8088 6960 8152
rect 6880 7992 6960 8088
rect 6880 7928 6888 7992
rect 6952 7928 6960 7992
rect 6880 7920 6960 7928
rect 7200 8312 7280 8320
rect 7200 8248 7208 8312
rect 7272 8248 7280 8312
rect 7200 8152 7280 8248
rect 7200 8088 7208 8152
rect 7272 8088 7280 8152
rect 7200 7992 7280 8088
rect 7200 7928 7208 7992
rect 7272 7928 7280 7992
rect 7200 7920 7280 7928
rect 7360 8312 7440 8320
rect 7360 8248 7368 8312
rect 7432 8248 7440 8312
rect 7360 8152 7440 8248
rect 7360 8088 7368 8152
rect 7432 8088 7440 8152
rect 7360 7992 7440 8088
rect 7360 7928 7368 7992
rect 7432 7928 7440 7992
rect 7360 7920 7440 7928
rect 7520 8312 7600 8320
rect 7520 8248 7528 8312
rect 7592 8248 7600 8312
rect 7520 8152 7600 8248
rect 7520 8088 7528 8152
rect 7592 8088 7600 8152
rect 7520 7992 7600 8088
rect 7520 7928 7528 7992
rect 7592 7928 7600 7992
rect 7520 7920 7600 7928
rect 7680 8312 7760 8320
rect 7680 8248 7688 8312
rect 7752 8248 7760 8312
rect 7680 8152 7760 8248
rect 7680 8088 7688 8152
rect 7752 8088 7760 8152
rect 7680 7992 7760 8088
rect 7680 7928 7688 7992
rect 7752 7928 7760 7992
rect 7680 7920 7760 7928
rect 7840 8312 7920 8320
rect 7840 8248 7848 8312
rect 7912 8248 7920 8312
rect 7840 8152 7920 8248
rect 7840 8088 7848 8152
rect 7912 8088 7920 8152
rect 7840 7992 7920 8088
rect 7840 7928 7848 7992
rect 7912 7928 7920 7992
rect 7840 7920 7920 7928
rect 8000 8312 8080 8320
rect 8000 8248 8008 8312
rect 8072 8248 8080 8312
rect 8000 8152 8080 8248
rect 8000 8088 8008 8152
rect 8072 8088 8080 8152
rect 8000 7992 8080 8088
rect 8000 7928 8008 7992
rect 8072 7928 8080 7992
rect 8000 7920 8080 7928
rect 8160 8312 8240 8320
rect 8160 8248 8168 8312
rect 8232 8248 8240 8312
rect 8160 8152 8240 8248
rect 8160 8088 8168 8152
rect 8232 8088 8240 8152
rect 8160 7992 8240 8088
rect 8160 7928 8168 7992
rect 8232 7928 8240 7992
rect 8160 7920 8240 7928
rect 320 7692 400 7720
rect 320 7628 328 7692
rect 392 7628 400 7692
rect 320 7612 400 7628
rect 320 7548 328 7612
rect 392 7548 400 7612
rect 320 7520 400 7548
rect 320 7092 400 7120
rect 320 7028 328 7092
rect 392 7028 400 7092
rect 320 7012 400 7028
rect 320 6948 328 7012
rect 392 6948 400 7012
rect 320 6920 400 6948
rect 160 6712 240 6720
rect 160 6648 168 6712
rect 232 6648 240 6712
rect 160 6552 240 6648
rect 160 6488 168 6552
rect 232 6488 240 6552
rect 160 6392 240 6488
rect 160 6328 168 6392
rect 232 6328 240 6392
rect 160 6320 240 6328
rect 320 6712 400 6720
rect 320 6648 328 6712
rect 392 6648 400 6712
rect 320 6552 400 6648
rect 320 6488 328 6552
rect 392 6488 400 6552
rect 320 6392 400 6488
rect 320 6328 328 6392
rect 392 6328 400 6392
rect 320 6320 400 6328
rect 480 6712 560 6720
rect 480 6648 488 6712
rect 552 6648 560 6712
rect 480 6552 560 6648
rect 480 6488 488 6552
rect 552 6488 560 6552
rect 480 6392 560 6488
rect 480 6328 488 6392
rect 552 6328 560 6392
rect 480 6320 560 6328
rect 640 6712 720 6720
rect 640 6648 648 6712
rect 712 6648 720 6712
rect 640 6552 720 6648
rect 640 6488 648 6552
rect 712 6488 720 6552
rect 640 6392 720 6488
rect 640 6328 648 6392
rect 712 6328 720 6392
rect 640 6320 720 6328
rect 800 6712 880 6720
rect 800 6648 808 6712
rect 872 6648 880 6712
rect 800 6552 880 6648
rect 800 6488 808 6552
rect 872 6488 880 6552
rect 800 6392 880 6488
rect 800 6328 808 6392
rect 872 6328 880 6392
rect 800 6320 880 6328
rect 960 6712 1040 6720
rect 960 6648 968 6712
rect 1032 6648 1040 6712
rect 960 6552 1040 6648
rect 960 6488 968 6552
rect 1032 6488 1040 6552
rect 960 6392 1040 6488
rect 960 6328 968 6392
rect 1032 6328 1040 6392
rect 960 6320 1040 6328
rect 1120 6712 1200 6720
rect 1120 6648 1128 6712
rect 1192 6648 1200 6712
rect 1120 6552 1200 6648
rect 1120 6488 1128 6552
rect 1192 6488 1200 6552
rect 1120 6392 1200 6488
rect 1120 6328 1128 6392
rect 1192 6328 1200 6392
rect 1120 6320 1200 6328
rect 1440 6712 1520 6720
rect 1440 6648 1448 6712
rect 1512 6648 1520 6712
rect 1440 6552 1520 6648
rect 1440 6488 1448 6552
rect 1512 6488 1520 6552
rect 1440 6392 1520 6488
rect 1440 6328 1448 6392
rect 1512 6328 1520 6392
rect 1440 6320 1520 6328
rect 1600 6712 1680 6720
rect 1600 6648 1608 6712
rect 1672 6648 1680 6712
rect 1600 6552 1680 6648
rect 1600 6488 1608 6552
rect 1672 6488 1680 6552
rect 1600 6392 1680 6488
rect 1600 6328 1608 6392
rect 1672 6328 1680 6392
rect 1600 6320 1680 6328
rect 1760 6712 1840 6720
rect 1760 6648 1768 6712
rect 1832 6648 1840 6712
rect 1760 6552 1840 6648
rect 1760 6488 1768 6552
rect 1832 6488 1840 6552
rect 1760 6392 1840 6488
rect 1760 6328 1768 6392
rect 1832 6328 1840 6392
rect 1760 6320 1840 6328
rect 1920 6712 2000 6720
rect 1920 6648 1928 6712
rect 1992 6648 2000 6712
rect 1920 6552 2000 6648
rect 1920 6488 1928 6552
rect 1992 6488 2000 6552
rect 1920 6392 2000 6488
rect 1920 6328 1928 6392
rect 1992 6328 2000 6392
rect 1920 6320 2000 6328
rect 2080 6712 2160 6720
rect 2080 6648 2088 6712
rect 2152 6648 2160 6712
rect 2080 6552 2160 6648
rect 2080 6488 2088 6552
rect 2152 6488 2160 6552
rect 2080 6392 2160 6488
rect 2080 6328 2088 6392
rect 2152 6328 2160 6392
rect 2080 6320 2160 6328
rect 2240 6712 2320 6720
rect 2240 6648 2248 6712
rect 2312 6648 2320 6712
rect 2240 6552 2320 6648
rect 2240 6488 2248 6552
rect 2312 6488 2320 6552
rect 2240 6392 2320 6488
rect 2240 6328 2248 6392
rect 2312 6328 2320 6392
rect 2240 6320 2320 6328
rect 2400 6712 2480 6720
rect 2400 6648 2408 6712
rect 2472 6648 2480 6712
rect 2400 6552 2480 6648
rect 2400 6488 2408 6552
rect 2472 6488 2480 6552
rect 2400 6392 2480 6488
rect 2400 6328 2408 6392
rect 2472 6328 2480 6392
rect 2400 6320 2480 6328
rect 2560 6712 2640 6720
rect 2560 6648 2568 6712
rect 2632 6648 2640 6712
rect 2560 6552 2640 6648
rect 2560 6488 2568 6552
rect 2632 6488 2640 6552
rect 2560 6392 2640 6488
rect 2560 6328 2568 6392
rect 2632 6328 2640 6392
rect 2560 6320 2640 6328
rect 2720 6712 2800 6720
rect 2720 6648 2728 6712
rect 2792 6648 2800 6712
rect 2720 6552 2800 6648
rect 2720 6488 2728 6552
rect 2792 6488 2800 6552
rect 2720 6392 2800 6488
rect 2720 6328 2728 6392
rect 2792 6328 2800 6392
rect 2720 6320 2800 6328
rect 2880 6712 2960 6720
rect 2880 6648 2888 6712
rect 2952 6648 2960 6712
rect 2880 6552 2960 6648
rect 2880 6488 2888 6552
rect 2952 6488 2960 6552
rect 2880 6392 2960 6488
rect 2880 6328 2888 6392
rect 2952 6328 2960 6392
rect 2880 6320 2960 6328
rect 3040 6712 3120 6720
rect 3040 6648 3048 6712
rect 3112 6648 3120 6712
rect 3040 6552 3120 6648
rect 3040 6488 3048 6552
rect 3112 6488 3120 6552
rect 3040 6392 3120 6488
rect 3040 6328 3048 6392
rect 3112 6328 3120 6392
rect 3040 6320 3120 6328
rect 3360 6712 3440 6720
rect 3360 6648 3368 6712
rect 3432 6648 3440 6712
rect 3360 6552 3440 6648
rect 3360 6488 3368 6552
rect 3432 6488 3440 6552
rect 3360 6392 3440 6488
rect 3360 6328 3368 6392
rect 3432 6328 3440 6392
rect 3360 6320 3440 6328
rect 3520 6712 3600 6720
rect 3520 6648 3528 6712
rect 3592 6648 3600 6712
rect 3520 6552 3600 6648
rect 3520 6488 3528 6552
rect 3592 6488 3600 6552
rect 3520 6392 3600 6488
rect 3520 6328 3528 6392
rect 3592 6328 3600 6392
rect 3520 6320 3600 6328
rect 3680 6712 3760 6720
rect 3680 6648 3688 6712
rect 3752 6648 3760 6712
rect 3680 6552 3760 6648
rect 3680 6488 3688 6552
rect 3752 6488 3760 6552
rect 3680 6392 3760 6488
rect 3680 6328 3688 6392
rect 3752 6328 3760 6392
rect 3680 6320 3760 6328
rect 3840 6712 3920 6720
rect 3840 6648 3848 6712
rect 3912 6648 3920 6712
rect 3840 6552 3920 6648
rect 3840 6488 3848 6552
rect 3912 6488 3920 6552
rect 3840 6392 3920 6488
rect 3840 6328 3848 6392
rect 3912 6328 3920 6392
rect 3840 6320 3920 6328
rect 4000 6712 4080 6720
rect 4000 6648 4008 6712
rect 4072 6648 4080 6712
rect 4000 6552 4080 6648
rect 4000 6488 4008 6552
rect 4072 6488 4080 6552
rect 4000 6392 4080 6488
rect 4000 6328 4008 6392
rect 4072 6328 4080 6392
rect 4000 6320 4080 6328
rect 4160 6712 4240 6720
rect 4160 6648 4168 6712
rect 4232 6648 4240 6712
rect 4160 6552 4240 6648
rect 4160 6488 4168 6552
rect 4232 6488 4240 6552
rect 4160 6392 4240 6488
rect 4160 6328 4168 6392
rect 4232 6328 4240 6392
rect 4160 6320 4240 6328
rect 4320 6712 4400 6720
rect 4320 6648 4328 6712
rect 4392 6648 4400 6712
rect 4320 6552 4400 6648
rect 4320 6488 4328 6552
rect 4392 6488 4400 6552
rect 4320 6392 4400 6488
rect 4320 6328 4328 6392
rect 4392 6328 4400 6392
rect 4320 6320 4400 6328
rect 4480 6712 4560 6720
rect 4480 6648 4488 6712
rect 4552 6648 4560 6712
rect 4480 6552 4560 6648
rect 4480 6488 4488 6552
rect 4552 6488 4560 6552
rect 4480 6392 4560 6488
rect 4480 6328 4488 6392
rect 4552 6328 4560 6392
rect 4480 6320 4560 6328
rect 4640 6712 4720 6720
rect 4640 6648 4648 6712
rect 4712 6648 4720 6712
rect 4640 6552 4720 6648
rect 4640 6488 4648 6552
rect 4712 6488 4720 6552
rect 4640 6392 4720 6488
rect 4640 6328 4648 6392
rect 4712 6328 4720 6392
rect 4640 6320 4720 6328
rect 4800 6712 4880 6720
rect 4800 6648 4808 6712
rect 4872 6648 4880 6712
rect 4800 6552 4880 6648
rect 4800 6488 4808 6552
rect 4872 6488 4880 6552
rect 4800 6392 4880 6488
rect 4800 6328 4808 6392
rect 4872 6328 4880 6392
rect 4800 6320 4880 6328
rect 4960 6712 5040 6720
rect 4960 6648 4968 6712
rect 5032 6648 5040 6712
rect 4960 6552 5040 6648
rect 4960 6488 4968 6552
rect 5032 6488 5040 6552
rect 4960 6392 5040 6488
rect 4960 6328 4968 6392
rect 5032 6328 5040 6392
rect 4960 6320 5040 6328
rect 5280 6712 5360 6720
rect 5280 6648 5288 6712
rect 5352 6648 5360 6712
rect 5280 6552 5360 6648
rect 5280 6488 5288 6552
rect 5352 6488 5360 6552
rect 5280 6392 5360 6488
rect 5280 6328 5288 6392
rect 5352 6328 5360 6392
rect 5280 6320 5360 6328
rect 5440 6712 5520 6720
rect 5440 6648 5448 6712
rect 5512 6648 5520 6712
rect 5440 6552 5520 6648
rect 5440 6488 5448 6552
rect 5512 6488 5520 6552
rect 5440 6392 5520 6488
rect 5440 6328 5448 6392
rect 5512 6328 5520 6392
rect 5440 6320 5520 6328
rect 5600 6712 5680 6720
rect 5600 6648 5608 6712
rect 5672 6648 5680 6712
rect 5600 6552 5680 6648
rect 5600 6488 5608 6552
rect 5672 6488 5680 6552
rect 5600 6392 5680 6488
rect 5600 6328 5608 6392
rect 5672 6328 5680 6392
rect 5600 6320 5680 6328
rect 5760 6712 5840 6720
rect 5760 6648 5768 6712
rect 5832 6648 5840 6712
rect 5760 6552 5840 6648
rect 5760 6488 5768 6552
rect 5832 6488 5840 6552
rect 5760 6392 5840 6488
rect 5760 6328 5768 6392
rect 5832 6328 5840 6392
rect 5760 6320 5840 6328
rect 5920 6712 6000 6720
rect 5920 6648 5928 6712
rect 5992 6648 6000 6712
rect 5920 6552 6000 6648
rect 5920 6488 5928 6552
rect 5992 6488 6000 6552
rect 5920 6392 6000 6488
rect 5920 6328 5928 6392
rect 5992 6328 6000 6392
rect 5920 6320 6000 6328
rect 6080 6712 6160 6720
rect 6080 6648 6088 6712
rect 6152 6648 6160 6712
rect 6080 6552 6160 6648
rect 6080 6488 6088 6552
rect 6152 6488 6160 6552
rect 6080 6392 6160 6488
rect 6080 6328 6088 6392
rect 6152 6328 6160 6392
rect 6080 6320 6160 6328
rect 6240 6712 6320 6720
rect 6240 6648 6248 6712
rect 6312 6648 6320 6712
rect 6240 6552 6320 6648
rect 6240 6488 6248 6552
rect 6312 6488 6320 6552
rect 6240 6392 6320 6488
rect 6240 6328 6248 6392
rect 6312 6328 6320 6392
rect 6240 6320 6320 6328
rect 6400 6712 6480 6720
rect 6400 6648 6408 6712
rect 6472 6648 6480 6712
rect 6400 6552 6480 6648
rect 6400 6488 6408 6552
rect 6472 6488 6480 6552
rect 6400 6392 6480 6488
rect 6400 6328 6408 6392
rect 6472 6328 6480 6392
rect 6400 6320 6480 6328
rect 6560 6712 6640 6720
rect 6560 6648 6568 6712
rect 6632 6648 6640 6712
rect 6560 6552 6640 6648
rect 6560 6488 6568 6552
rect 6632 6488 6640 6552
rect 6560 6392 6640 6488
rect 6560 6328 6568 6392
rect 6632 6328 6640 6392
rect 6560 6320 6640 6328
rect 6720 6712 6800 6720
rect 6720 6648 6728 6712
rect 6792 6648 6800 6712
rect 6720 6552 6800 6648
rect 6720 6488 6728 6552
rect 6792 6488 6800 6552
rect 6720 6392 6800 6488
rect 6720 6328 6728 6392
rect 6792 6328 6800 6392
rect 6720 6320 6800 6328
rect 6880 6712 6960 6720
rect 6880 6648 6888 6712
rect 6952 6648 6960 6712
rect 6880 6552 6960 6648
rect 6880 6488 6888 6552
rect 6952 6488 6960 6552
rect 6880 6392 6960 6488
rect 6880 6328 6888 6392
rect 6952 6328 6960 6392
rect 6880 6320 6960 6328
rect 7200 6712 7280 6720
rect 7200 6648 7208 6712
rect 7272 6648 7280 6712
rect 7200 6552 7280 6648
rect 7200 6488 7208 6552
rect 7272 6488 7280 6552
rect 7200 6392 7280 6488
rect 7200 6328 7208 6392
rect 7272 6328 7280 6392
rect 7200 6320 7280 6328
rect 7360 6712 7440 6720
rect 7360 6648 7368 6712
rect 7432 6648 7440 6712
rect 7360 6552 7440 6648
rect 7360 6488 7368 6552
rect 7432 6488 7440 6552
rect 7360 6392 7440 6488
rect 7360 6328 7368 6392
rect 7432 6328 7440 6392
rect 7360 6320 7440 6328
rect 7520 6712 7600 6720
rect 7520 6648 7528 6712
rect 7592 6648 7600 6712
rect 7520 6552 7600 6648
rect 7520 6488 7528 6552
rect 7592 6488 7600 6552
rect 7520 6392 7600 6488
rect 7520 6328 7528 6392
rect 7592 6328 7600 6392
rect 7520 6320 7600 6328
rect 7680 6712 7760 6720
rect 7680 6648 7688 6712
rect 7752 6648 7760 6712
rect 7680 6552 7760 6648
rect 7680 6488 7688 6552
rect 7752 6488 7760 6552
rect 7680 6392 7760 6488
rect 7680 6328 7688 6392
rect 7752 6328 7760 6392
rect 7680 6320 7760 6328
rect 7840 6712 7920 6720
rect 7840 6648 7848 6712
rect 7912 6648 7920 6712
rect 7840 6552 7920 6648
rect 7840 6488 7848 6552
rect 7912 6488 7920 6552
rect 7840 6392 7920 6488
rect 7840 6328 7848 6392
rect 7912 6328 7920 6392
rect 7840 6320 7920 6328
rect 8160 6712 8240 6720
rect 8160 6648 8168 6712
rect 8232 6648 8240 6712
rect 8160 6552 8240 6648
rect 8160 6488 8168 6552
rect 8232 6488 8240 6552
rect 8160 6392 8240 6488
rect 8160 6328 8168 6392
rect 8232 6328 8240 6392
rect 8160 6320 8240 6328
rect 160 6232 240 6240
rect 160 6168 168 6232
rect 232 6168 240 6232
rect 160 6072 240 6168
rect 160 6008 168 6072
rect 232 6008 240 6072
rect 160 5912 240 6008
rect 160 5848 168 5912
rect 232 5848 240 5912
rect 160 5840 240 5848
rect 320 6232 400 6240
rect 320 6168 328 6232
rect 392 6168 400 6232
rect 320 6072 400 6168
rect 320 6008 328 6072
rect 392 6008 400 6072
rect 320 5912 400 6008
rect 320 5848 328 5912
rect 392 5848 400 5912
rect 320 5840 400 5848
rect 480 6232 560 6240
rect 480 6168 488 6232
rect 552 6168 560 6232
rect 480 6072 560 6168
rect 480 6008 488 6072
rect 552 6008 560 6072
rect 480 5912 560 6008
rect 480 5848 488 5912
rect 552 5848 560 5912
rect 480 5840 560 5848
rect 640 6232 720 6240
rect 640 6168 648 6232
rect 712 6168 720 6232
rect 640 6072 720 6168
rect 640 6008 648 6072
rect 712 6008 720 6072
rect 640 5912 720 6008
rect 640 5848 648 5912
rect 712 5848 720 5912
rect 640 5840 720 5848
rect 800 6232 880 6240
rect 800 6168 808 6232
rect 872 6168 880 6232
rect 800 6072 880 6168
rect 800 6008 808 6072
rect 872 6008 880 6072
rect 800 5912 880 6008
rect 800 5848 808 5912
rect 872 5848 880 5912
rect 800 5840 880 5848
rect 960 6232 1040 6240
rect 960 6168 968 6232
rect 1032 6168 1040 6232
rect 960 6072 1040 6168
rect 960 6008 968 6072
rect 1032 6008 1040 6072
rect 960 5912 1040 6008
rect 960 5848 968 5912
rect 1032 5848 1040 5912
rect 960 5840 1040 5848
rect 1120 6232 1200 6240
rect 1120 6168 1128 6232
rect 1192 6168 1200 6232
rect 1120 6072 1200 6168
rect 1120 6008 1128 6072
rect 1192 6008 1200 6072
rect 1120 5912 1200 6008
rect 1120 5848 1128 5912
rect 1192 5848 1200 5912
rect 1120 5840 1200 5848
rect 1280 6232 1360 6240
rect 1280 6168 1288 6232
rect 1352 6168 1360 6232
rect 1280 6072 1360 6168
rect 1280 6008 1288 6072
rect 1352 6008 1360 6072
rect 1280 5912 1360 6008
rect 1280 5848 1288 5912
rect 1352 5848 1360 5912
rect 1280 5840 1360 5848
rect 1440 6232 1520 6240
rect 1440 6168 1448 6232
rect 1512 6168 1520 6232
rect 1440 6072 1520 6168
rect 1440 6008 1448 6072
rect 1512 6008 1520 6072
rect 1440 5912 1520 6008
rect 1440 5848 1448 5912
rect 1512 5848 1520 5912
rect 1440 5840 1520 5848
rect 1600 6232 1680 6240
rect 1600 6168 1608 6232
rect 1672 6168 1680 6232
rect 1600 6072 1680 6168
rect 1600 6008 1608 6072
rect 1672 6008 1680 6072
rect 1600 5912 1680 6008
rect 1600 5848 1608 5912
rect 1672 5848 1680 5912
rect 1600 5840 1680 5848
rect 1760 6232 1840 6240
rect 1760 6168 1768 6232
rect 1832 6168 1840 6232
rect 1760 6072 1840 6168
rect 1760 6008 1768 6072
rect 1832 6008 1840 6072
rect 1760 5912 1840 6008
rect 1760 5848 1768 5912
rect 1832 5848 1840 5912
rect 1760 5840 1840 5848
rect 1920 6232 2000 6240
rect 1920 6168 1928 6232
rect 1992 6168 2000 6232
rect 1920 6072 2000 6168
rect 1920 6008 1928 6072
rect 1992 6008 2000 6072
rect 1920 5912 2000 6008
rect 1920 5848 1928 5912
rect 1992 5848 2000 5912
rect 1920 5840 2000 5848
rect 2080 6232 2160 6240
rect 2080 6168 2088 6232
rect 2152 6168 2160 6232
rect 2080 6072 2160 6168
rect 2080 6008 2088 6072
rect 2152 6008 2160 6072
rect 2080 5912 2160 6008
rect 2080 5848 2088 5912
rect 2152 5848 2160 5912
rect 2080 5840 2160 5848
rect 2240 6232 2320 6240
rect 2240 6168 2248 6232
rect 2312 6168 2320 6232
rect 2240 6072 2320 6168
rect 2240 6008 2248 6072
rect 2312 6008 2320 6072
rect 2240 5912 2320 6008
rect 2240 5848 2248 5912
rect 2312 5848 2320 5912
rect 2240 5840 2320 5848
rect 2400 6232 2480 6240
rect 2400 6168 2408 6232
rect 2472 6168 2480 6232
rect 2400 6072 2480 6168
rect 2400 6008 2408 6072
rect 2472 6008 2480 6072
rect 2400 5912 2480 6008
rect 2400 5848 2408 5912
rect 2472 5848 2480 5912
rect 2400 5840 2480 5848
rect 2560 6232 2640 6240
rect 2560 6168 2568 6232
rect 2632 6168 2640 6232
rect 2560 6072 2640 6168
rect 2560 6008 2568 6072
rect 2632 6008 2640 6072
rect 2560 5912 2640 6008
rect 2560 5848 2568 5912
rect 2632 5848 2640 5912
rect 2560 5840 2640 5848
rect 2720 6232 2800 6240
rect 2720 6168 2728 6232
rect 2792 6168 2800 6232
rect 2720 6072 2800 6168
rect 2720 6008 2728 6072
rect 2792 6008 2800 6072
rect 2720 5912 2800 6008
rect 2720 5848 2728 5912
rect 2792 5848 2800 5912
rect 2720 5840 2800 5848
rect 2880 6232 2960 6240
rect 2880 6168 2888 6232
rect 2952 6168 2960 6232
rect 2880 6072 2960 6168
rect 2880 6008 2888 6072
rect 2952 6008 2960 6072
rect 2880 5912 2960 6008
rect 2880 5848 2888 5912
rect 2952 5848 2960 5912
rect 2880 5840 2960 5848
rect 3040 6232 3120 6240
rect 3040 6168 3048 6232
rect 3112 6168 3120 6232
rect 3040 6072 3120 6168
rect 3040 6008 3048 6072
rect 3112 6008 3120 6072
rect 3040 5912 3120 6008
rect 3040 5848 3048 5912
rect 3112 5848 3120 5912
rect 3040 5840 3120 5848
rect 3200 6232 3280 6240
rect 3200 6168 3208 6232
rect 3272 6168 3280 6232
rect 3200 6072 3280 6168
rect 3200 6008 3208 6072
rect 3272 6008 3280 6072
rect 3200 5912 3280 6008
rect 3200 5848 3208 5912
rect 3272 5848 3280 5912
rect 3200 5840 3280 5848
rect 3360 6232 3440 6240
rect 3360 6168 3368 6232
rect 3432 6168 3440 6232
rect 3360 6072 3440 6168
rect 3360 6008 3368 6072
rect 3432 6008 3440 6072
rect 3360 5912 3440 6008
rect 3360 5848 3368 5912
rect 3432 5848 3440 5912
rect 3360 5840 3440 5848
rect 3520 6232 3600 6240
rect 3520 6168 3528 6232
rect 3592 6168 3600 6232
rect 3520 6072 3600 6168
rect 3520 6008 3528 6072
rect 3592 6008 3600 6072
rect 3520 5912 3600 6008
rect 3520 5848 3528 5912
rect 3592 5848 3600 5912
rect 3520 5840 3600 5848
rect 3680 6232 3760 6240
rect 3680 6168 3688 6232
rect 3752 6168 3760 6232
rect 3680 6072 3760 6168
rect 3680 6008 3688 6072
rect 3752 6008 3760 6072
rect 3680 5912 3760 6008
rect 3680 5848 3688 5912
rect 3752 5848 3760 5912
rect 3680 5840 3760 5848
rect 3840 6232 3920 6240
rect 3840 6168 3848 6232
rect 3912 6168 3920 6232
rect 3840 6072 3920 6168
rect 3840 6008 3848 6072
rect 3912 6008 3920 6072
rect 3840 5912 3920 6008
rect 3840 5848 3848 5912
rect 3912 5848 3920 5912
rect 3840 5840 3920 5848
rect 4000 6232 4080 6240
rect 4000 6168 4008 6232
rect 4072 6168 4080 6232
rect 4000 6072 4080 6168
rect 4000 6008 4008 6072
rect 4072 6008 4080 6072
rect 4000 5912 4080 6008
rect 4000 5848 4008 5912
rect 4072 5848 4080 5912
rect 4000 5840 4080 5848
rect 4160 6232 4240 6240
rect 4160 6168 4168 6232
rect 4232 6168 4240 6232
rect 4160 6072 4240 6168
rect 4160 6008 4168 6072
rect 4232 6008 4240 6072
rect 4160 5912 4240 6008
rect 4160 5848 4168 5912
rect 4232 5848 4240 5912
rect 4160 5840 4240 5848
rect 4320 6232 4400 6240
rect 4320 6168 4328 6232
rect 4392 6168 4400 6232
rect 4320 6072 4400 6168
rect 4320 6008 4328 6072
rect 4392 6008 4400 6072
rect 4320 5912 4400 6008
rect 4320 5848 4328 5912
rect 4392 5848 4400 5912
rect 4320 5840 4400 5848
rect 4480 6232 4560 6240
rect 4480 6168 4488 6232
rect 4552 6168 4560 6232
rect 4480 6072 4560 6168
rect 4480 6008 4488 6072
rect 4552 6008 4560 6072
rect 4480 5912 4560 6008
rect 4480 5848 4488 5912
rect 4552 5848 4560 5912
rect 4480 5840 4560 5848
rect 4640 6232 4720 6240
rect 4640 6168 4648 6232
rect 4712 6168 4720 6232
rect 4640 6072 4720 6168
rect 4640 6008 4648 6072
rect 4712 6008 4720 6072
rect 4640 5912 4720 6008
rect 4640 5848 4648 5912
rect 4712 5848 4720 5912
rect 4640 5840 4720 5848
rect 4800 6232 4880 6240
rect 4800 6168 4808 6232
rect 4872 6168 4880 6232
rect 4800 6072 4880 6168
rect 4800 6008 4808 6072
rect 4872 6008 4880 6072
rect 4800 5912 4880 6008
rect 4800 5848 4808 5912
rect 4872 5848 4880 5912
rect 4800 5840 4880 5848
rect 4960 6232 5040 6240
rect 4960 6168 4968 6232
rect 5032 6168 5040 6232
rect 4960 6072 5040 6168
rect 4960 6008 4968 6072
rect 5032 6008 5040 6072
rect 4960 5912 5040 6008
rect 4960 5848 4968 5912
rect 5032 5848 5040 5912
rect 4960 5840 5040 5848
rect 5120 6232 5200 6240
rect 5120 6168 5128 6232
rect 5192 6168 5200 6232
rect 5120 6072 5200 6168
rect 5120 6008 5128 6072
rect 5192 6008 5200 6072
rect 5120 5912 5200 6008
rect 5120 5848 5128 5912
rect 5192 5848 5200 5912
rect 5120 5840 5200 5848
rect 5280 6232 5360 6240
rect 5280 6168 5288 6232
rect 5352 6168 5360 6232
rect 5280 6072 5360 6168
rect 5280 6008 5288 6072
rect 5352 6008 5360 6072
rect 5280 5912 5360 6008
rect 5280 5848 5288 5912
rect 5352 5848 5360 5912
rect 5280 5840 5360 5848
rect 5440 6232 5520 6240
rect 5440 6168 5448 6232
rect 5512 6168 5520 6232
rect 5440 6072 5520 6168
rect 5440 6008 5448 6072
rect 5512 6008 5520 6072
rect 5440 5912 5520 6008
rect 5440 5848 5448 5912
rect 5512 5848 5520 5912
rect 5440 5840 5520 5848
rect 5600 6232 5680 6240
rect 5600 6168 5608 6232
rect 5672 6168 5680 6232
rect 5600 6072 5680 6168
rect 5600 6008 5608 6072
rect 5672 6008 5680 6072
rect 5600 5912 5680 6008
rect 5600 5848 5608 5912
rect 5672 5848 5680 5912
rect 5600 5840 5680 5848
rect 5760 6232 5840 6240
rect 5760 6168 5768 6232
rect 5832 6168 5840 6232
rect 5760 6072 5840 6168
rect 5760 6008 5768 6072
rect 5832 6008 5840 6072
rect 5760 5912 5840 6008
rect 5760 5848 5768 5912
rect 5832 5848 5840 5912
rect 5760 5840 5840 5848
rect 5920 6232 6000 6240
rect 5920 6168 5928 6232
rect 5992 6168 6000 6232
rect 5920 6072 6000 6168
rect 5920 6008 5928 6072
rect 5992 6008 6000 6072
rect 5920 5912 6000 6008
rect 5920 5848 5928 5912
rect 5992 5848 6000 5912
rect 5920 5840 6000 5848
rect 6080 6232 6160 6240
rect 6080 6168 6088 6232
rect 6152 6168 6160 6232
rect 6080 6072 6160 6168
rect 6080 6008 6088 6072
rect 6152 6008 6160 6072
rect 6080 5912 6160 6008
rect 6080 5848 6088 5912
rect 6152 5848 6160 5912
rect 6080 5840 6160 5848
rect 6240 6232 6320 6240
rect 6240 6168 6248 6232
rect 6312 6168 6320 6232
rect 6240 6072 6320 6168
rect 6240 6008 6248 6072
rect 6312 6008 6320 6072
rect 6240 5912 6320 6008
rect 6240 5848 6248 5912
rect 6312 5848 6320 5912
rect 6240 5840 6320 5848
rect 6400 6232 6480 6240
rect 6400 6168 6408 6232
rect 6472 6168 6480 6232
rect 6400 6072 6480 6168
rect 6400 6008 6408 6072
rect 6472 6008 6480 6072
rect 6400 5912 6480 6008
rect 6400 5848 6408 5912
rect 6472 5848 6480 5912
rect 6400 5840 6480 5848
rect 6560 6232 6640 6240
rect 6560 6168 6568 6232
rect 6632 6168 6640 6232
rect 6560 6072 6640 6168
rect 6560 6008 6568 6072
rect 6632 6008 6640 6072
rect 6560 5912 6640 6008
rect 6560 5848 6568 5912
rect 6632 5848 6640 5912
rect 6560 5840 6640 5848
rect 6720 6232 6800 6240
rect 6720 6168 6728 6232
rect 6792 6168 6800 6232
rect 6720 6072 6800 6168
rect 6720 6008 6728 6072
rect 6792 6008 6800 6072
rect 6720 5912 6800 6008
rect 6720 5848 6728 5912
rect 6792 5848 6800 5912
rect 6720 5840 6800 5848
rect 6880 6232 6960 6240
rect 6880 6168 6888 6232
rect 6952 6168 6960 6232
rect 6880 6072 6960 6168
rect 6880 6008 6888 6072
rect 6952 6008 6960 6072
rect 6880 5912 6960 6008
rect 6880 5848 6888 5912
rect 6952 5848 6960 5912
rect 6880 5840 6960 5848
rect 7040 6232 7120 6240
rect 7040 6168 7048 6232
rect 7112 6168 7120 6232
rect 7040 6072 7120 6168
rect 7040 6008 7048 6072
rect 7112 6008 7120 6072
rect 7040 5912 7120 6008
rect 7040 5848 7048 5912
rect 7112 5848 7120 5912
rect 7040 5840 7120 5848
rect 7200 6232 7280 6240
rect 7200 6168 7208 6232
rect 7272 6168 7280 6232
rect 7200 6072 7280 6168
rect 7200 6008 7208 6072
rect 7272 6008 7280 6072
rect 7200 5912 7280 6008
rect 7200 5848 7208 5912
rect 7272 5848 7280 5912
rect 7200 5840 7280 5848
rect 7360 6232 7440 6240
rect 7360 6168 7368 6232
rect 7432 6168 7440 6232
rect 7360 6072 7440 6168
rect 7360 6008 7368 6072
rect 7432 6008 7440 6072
rect 7360 5912 7440 6008
rect 7360 5848 7368 5912
rect 7432 5848 7440 5912
rect 7360 5840 7440 5848
rect 7520 6232 7600 6240
rect 7520 6168 7528 6232
rect 7592 6168 7600 6232
rect 7520 6072 7600 6168
rect 7520 6008 7528 6072
rect 7592 6008 7600 6072
rect 7520 5912 7600 6008
rect 7520 5848 7528 5912
rect 7592 5848 7600 5912
rect 7520 5840 7600 5848
rect 7680 6232 7760 6240
rect 7680 6168 7688 6232
rect 7752 6168 7760 6232
rect 7680 6072 7760 6168
rect 7680 6008 7688 6072
rect 7752 6008 7760 6072
rect 7680 5912 7760 6008
rect 7680 5848 7688 5912
rect 7752 5848 7760 5912
rect 7680 5840 7760 5848
rect 7840 6232 7920 6240
rect 7840 6168 7848 6232
rect 7912 6168 7920 6232
rect 7840 6072 7920 6168
rect 7840 6008 7848 6072
rect 7912 6008 7920 6072
rect 7840 5912 7920 6008
rect 7840 5848 7848 5912
rect 7912 5848 7920 5912
rect 7840 5840 7920 5848
rect 8160 6232 8240 6240
rect 8160 6168 8168 6232
rect 8232 6168 8240 6232
rect 8160 6072 8240 6168
rect 8160 6008 8168 6072
rect 8232 6008 8240 6072
rect 8160 5912 8240 6008
rect 8160 5848 8168 5912
rect 8232 5848 8240 5912
rect 8160 5840 8240 5848
rect 160 5752 240 5760
rect 160 5688 168 5752
rect 232 5688 240 5752
rect 160 5592 240 5688
rect 160 5528 168 5592
rect 232 5528 240 5592
rect 160 5432 240 5528
rect 160 5368 168 5432
rect 232 5368 240 5432
rect 160 5360 240 5368
rect 320 5752 400 5760
rect 320 5688 328 5752
rect 392 5688 400 5752
rect 320 5592 400 5688
rect 320 5528 328 5592
rect 392 5528 400 5592
rect 320 5432 400 5528
rect 320 5368 328 5432
rect 392 5368 400 5432
rect 320 5360 400 5368
rect 480 5752 560 5760
rect 480 5688 488 5752
rect 552 5688 560 5752
rect 480 5592 560 5688
rect 480 5528 488 5592
rect 552 5528 560 5592
rect 480 5432 560 5528
rect 480 5368 488 5432
rect 552 5368 560 5432
rect 480 5360 560 5368
rect 640 5752 720 5760
rect 640 5688 648 5752
rect 712 5688 720 5752
rect 640 5592 720 5688
rect 640 5528 648 5592
rect 712 5528 720 5592
rect 640 5432 720 5528
rect 640 5368 648 5432
rect 712 5368 720 5432
rect 640 5360 720 5368
rect 800 5752 880 5760
rect 800 5688 808 5752
rect 872 5688 880 5752
rect 800 5592 880 5688
rect 800 5528 808 5592
rect 872 5528 880 5592
rect 800 5432 880 5528
rect 800 5368 808 5432
rect 872 5368 880 5432
rect 800 5360 880 5368
rect 960 5752 1040 5760
rect 960 5688 968 5752
rect 1032 5688 1040 5752
rect 960 5592 1040 5688
rect 960 5528 968 5592
rect 1032 5528 1040 5592
rect 960 5432 1040 5528
rect 960 5368 968 5432
rect 1032 5368 1040 5432
rect 960 5360 1040 5368
rect 1120 5752 1200 5760
rect 1120 5688 1128 5752
rect 1192 5688 1200 5752
rect 1120 5592 1200 5688
rect 1120 5528 1128 5592
rect 1192 5528 1200 5592
rect 1120 5432 1200 5528
rect 1120 5368 1128 5432
rect 1192 5368 1200 5432
rect 1120 5360 1200 5368
rect 1440 5752 1520 5760
rect 1440 5688 1448 5752
rect 1512 5688 1520 5752
rect 1440 5592 1520 5688
rect 1440 5528 1448 5592
rect 1512 5528 1520 5592
rect 1440 5432 1520 5528
rect 1440 5368 1448 5432
rect 1512 5368 1520 5432
rect 1440 5360 1520 5368
rect 1600 5752 1680 5760
rect 1600 5688 1608 5752
rect 1672 5688 1680 5752
rect 1600 5592 1680 5688
rect 1600 5528 1608 5592
rect 1672 5528 1680 5592
rect 1600 5432 1680 5528
rect 1600 5368 1608 5432
rect 1672 5368 1680 5432
rect 1600 5360 1680 5368
rect 1760 5752 1840 5760
rect 1760 5688 1768 5752
rect 1832 5688 1840 5752
rect 1760 5592 1840 5688
rect 1760 5528 1768 5592
rect 1832 5528 1840 5592
rect 1760 5432 1840 5528
rect 1760 5368 1768 5432
rect 1832 5368 1840 5432
rect 1760 5360 1840 5368
rect 1920 5752 2000 5760
rect 1920 5688 1928 5752
rect 1992 5688 2000 5752
rect 1920 5592 2000 5688
rect 1920 5528 1928 5592
rect 1992 5528 2000 5592
rect 1920 5432 2000 5528
rect 1920 5368 1928 5432
rect 1992 5368 2000 5432
rect 1920 5360 2000 5368
rect 2080 5752 2160 5760
rect 2080 5688 2088 5752
rect 2152 5688 2160 5752
rect 2080 5592 2160 5688
rect 2080 5528 2088 5592
rect 2152 5528 2160 5592
rect 2080 5432 2160 5528
rect 2080 5368 2088 5432
rect 2152 5368 2160 5432
rect 2080 5360 2160 5368
rect 2240 5752 2320 5760
rect 2240 5688 2248 5752
rect 2312 5688 2320 5752
rect 2240 5592 2320 5688
rect 2240 5528 2248 5592
rect 2312 5528 2320 5592
rect 2240 5432 2320 5528
rect 2240 5368 2248 5432
rect 2312 5368 2320 5432
rect 2240 5360 2320 5368
rect 2400 5752 2480 5760
rect 2400 5688 2408 5752
rect 2472 5688 2480 5752
rect 2400 5592 2480 5688
rect 2400 5528 2408 5592
rect 2472 5528 2480 5592
rect 2400 5432 2480 5528
rect 2400 5368 2408 5432
rect 2472 5368 2480 5432
rect 2400 5360 2480 5368
rect 2560 5752 2640 5760
rect 2560 5688 2568 5752
rect 2632 5688 2640 5752
rect 2560 5592 2640 5688
rect 2560 5528 2568 5592
rect 2632 5528 2640 5592
rect 2560 5432 2640 5528
rect 2560 5368 2568 5432
rect 2632 5368 2640 5432
rect 2560 5360 2640 5368
rect 2720 5752 2800 5760
rect 2720 5688 2728 5752
rect 2792 5688 2800 5752
rect 2720 5592 2800 5688
rect 2720 5528 2728 5592
rect 2792 5528 2800 5592
rect 2720 5432 2800 5528
rect 2720 5368 2728 5432
rect 2792 5368 2800 5432
rect 2720 5360 2800 5368
rect 2880 5752 2960 5760
rect 2880 5688 2888 5752
rect 2952 5688 2960 5752
rect 2880 5592 2960 5688
rect 2880 5528 2888 5592
rect 2952 5528 2960 5592
rect 2880 5432 2960 5528
rect 2880 5368 2888 5432
rect 2952 5368 2960 5432
rect 2880 5360 2960 5368
rect 3040 5752 3120 5760
rect 3040 5688 3048 5752
rect 3112 5688 3120 5752
rect 3040 5592 3120 5688
rect 3040 5528 3048 5592
rect 3112 5528 3120 5592
rect 3040 5432 3120 5528
rect 3040 5368 3048 5432
rect 3112 5368 3120 5432
rect 3040 5360 3120 5368
rect 3360 5752 3440 5760
rect 3360 5688 3368 5752
rect 3432 5688 3440 5752
rect 3360 5592 3440 5688
rect 3360 5528 3368 5592
rect 3432 5528 3440 5592
rect 3360 5432 3440 5528
rect 3360 5368 3368 5432
rect 3432 5368 3440 5432
rect 3360 5360 3440 5368
rect 3520 5752 3600 5760
rect 3520 5688 3528 5752
rect 3592 5688 3600 5752
rect 3520 5592 3600 5688
rect 3520 5528 3528 5592
rect 3592 5528 3600 5592
rect 3520 5432 3600 5528
rect 3520 5368 3528 5432
rect 3592 5368 3600 5432
rect 3520 5360 3600 5368
rect 3680 5752 3760 5760
rect 3680 5688 3688 5752
rect 3752 5688 3760 5752
rect 3680 5592 3760 5688
rect 3680 5528 3688 5592
rect 3752 5528 3760 5592
rect 3680 5432 3760 5528
rect 3680 5368 3688 5432
rect 3752 5368 3760 5432
rect 3680 5360 3760 5368
rect 3840 5752 3920 5760
rect 3840 5688 3848 5752
rect 3912 5688 3920 5752
rect 3840 5592 3920 5688
rect 3840 5528 3848 5592
rect 3912 5528 3920 5592
rect 3840 5432 3920 5528
rect 3840 5368 3848 5432
rect 3912 5368 3920 5432
rect 3840 5360 3920 5368
rect 4000 5752 4080 5760
rect 4000 5688 4008 5752
rect 4072 5688 4080 5752
rect 4000 5592 4080 5688
rect 4000 5528 4008 5592
rect 4072 5528 4080 5592
rect 4000 5432 4080 5528
rect 4000 5368 4008 5432
rect 4072 5368 4080 5432
rect 4000 5360 4080 5368
rect 4160 5752 4240 5760
rect 4160 5688 4168 5752
rect 4232 5688 4240 5752
rect 4160 5592 4240 5688
rect 4160 5528 4168 5592
rect 4232 5528 4240 5592
rect 4160 5432 4240 5528
rect 4160 5368 4168 5432
rect 4232 5368 4240 5432
rect 4160 5360 4240 5368
rect 4320 5752 4400 5760
rect 4320 5688 4328 5752
rect 4392 5688 4400 5752
rect 4320 5592 4400 5688
rect 4320 5528 4328 5592
rect 4392 5528 4400 5592
rect 4320 5432 4400 5528
rect 4320 5368 4328 5432
rect 4392 5368 4400 5432
rect 4320 5360 4400 5368
rect 4480 5752 4560 5760
rect 4480 5688 4488 5752
rect 4552 5688 4560 5752
rect 4480 5592 4560 5688
rect 4480 5528 4488 5592
rect 4552 5528 4560 5592
rect 4480 5432 4560 5528
rect 4480 5368 4488 5432
rect 4552 5368 4560 5432
rect 4480 5360 4560 5368
rect 4640 5752 4720 5760
rect 4640 5688 4648 5752
rect 4712 5688 4720 5752
rect 4640 5592 4720 5688
rect 4640 5528 4648 5592
rect 4712 5528 4720 5592
rect 4640 5432 4720 5528
rect 4640 5368 4648 5432
rect 4712 5368 4720 5432
rect 4640 5360 4720 5368
rect 4800 5752 4880 5760
rect 4800 5688 4808 5752
rect 4872 5688 4880 5752
rect 4800 5592 4880 5688
rect 4800 5528 4808 5592
rect 4872 5528 4880 5592
rect 4800 5432 4880 5528
rect 4800 5368 4808 5432
rect 4872 5368 4880 5432
rect 4800 5360 4880 5368
rect 4960 5752 5040 5760
rect 4960 5688 4968 5752
rect 5032 5688 5040 5752
rect 4960 5592 5040 5688
rect 4960 5528 4968 5592
rect 5032 5528 5040 5592
rect 4960 5432 5040 5528
rect 4960 5368 4968 5432
rect 5032 5368 5040 5432
rect 4960 5360 5040 5368
rect 5280 5752 5360 5760
rect 5280 5688 5288 5752
rect 5352 5688 5360 5752
rect 5280 5592 5360 5688
rect 5280 5528 5288 5592
rect 5352 5528 5360 5592
rect 5280 5432 5360 5528
rect 5280 5368 5288 5432
rect 5352 5368 5360 5432
rect 5280 5360 5360 5368
rect 5440 5752 5520 5760
rect 5440 5688 5448 5752
rect 5512 5688 5520 5752
rect 5440 5592 5520 5688
rect 5440 5528 5448 5592
rect 5512 5528 5520 5592
rect 5440 5432 5520 5528
rect 5440 5368 5448 5432
rect 5512 5368 5520 5432
rect 5440 5360 5520 5368
rect 5600 5752 5680 5760
rect 5600 5688 5608 5752
rect 5672 5688 5680 5752
rect 5600 5592 5680 5688
rect 5600 5528 5608 5592
rect 5672 5528 5680 5592
rect 5600 5432 5680 5528
rect 5600 5368 5608 5432
rect 5672 5368 5680 5432
rect 5600 5360 5680 5368
rect 5760 5752 5840 5760
rect 5760 5688 5768 5752
rect 5832 5688 5840 5752
rect 5760 5592 5840 5688
rect 5760 5528 5768 5592
rect 5832 5528 5840 5592
rect 5760 5432 5840 5528
rect 5760 5368 5768 5432
rect 5832 5368 5840 5432
rect 5760 5360 5840 5368
rect 5920 5752 6000 5760
rect 5920 5688 5928 5752
rect 5992 5688 6000 5752
rect 5920 5592 6000 5688
rect 5920 5528 5928 5592
rect 5992 5528 6000 5592
rect 5920 5432 6000 5528
rect 5920 5368 5928 5432
rect 5992 5368 6000 5432
rect 5920 5360 6000 5368
rect 6080 5752 6160 5760
rect 6080 5688 6088 5752
rect 6152 5688 6160 5752
rect 6080 5592 6160 5688
rect 6080 5528 6088 5592
rect 6152 5528 6160 5592
rect 6080 5432 6160 5528
rect 6080 5368 6088 5432
rect 6152 5368 6160 5432
rect 6080 5360 6160 5368
rect 6240 5752 6320 5760
rect 6240 5688 6248 5752
rect 6312 5688 6320 5752
rect 6240 5592 6320 5688
rect 6240 5528 6248 5592
rect 6312 5528 6320 5592
rect 6240 5432 6320 5528
rect 6240 5368 6248 5432
rect 6312 5368 6320 5432
rect 6240 5360 6320 5368
rect 6400 5752 6480 5760
rect 6400 5688 6408 5752
rect 6472 5688 6480 5752
rect 6400 5592 6480 5688
rect 6400 5528 6408 5592
rect 6472 5528 6480 5592
rect 6400 5432 6480 5528
rect 6400 5368 6408 5432
rect 6472 5368 6480 5432
rect 6400 5360 6480 5368
rect 6560 5752 6640 5760
rect 6560 5688 6568 5752
rect 6632 5688 6640 5752
rect 6560 5592 6640 5688
rect 6560 5528 6568 5592
rect 6632 5528 6640 5592
rect 6560 5432 6640 5528
rect 6560 5368 6568 5432
rect 6632 5368 6640 5432
rect 6560 5360 6640 5368
rect 6720 5752 6800 5760
rect 6720 5688 6728 5752
rect 6792 5688 6800 5752
rect 6720 5592 6800 5688
rect 6720 5528 6728 5592
rect 6792 5528 6800 5592
rect 6720 5432 6800 5528
rect 6720 5368 6728 5432
rect 6792 5368 6800 5432
rect 6720 5360 6800 5368
rect 6880 5752 6960 5760
rect 6880 5688 6888 5752
rect 6952 5688 6960 5752
rect 6880 5592 6960 5688
rect 6880 5528 6888 5592
rect 6952 5528 6960 5592
rect 6880 5432 6960 5528
rect 6880 5368 6888 5432
rect 6952 5368 6960 5432
rect 6880 5360 6960 5368
rect 7200 5752 7280 5760
rect 7200 5688 7208 5752
rect 7272 5688 7280 5752
rect 7200 5592 7280 5688
rect 7200 5528 7208 5592
rect 7272 5528 7280 5592
rect 7200 5432 7280 5528
rect 7200 5368 7208 5432
rect 7272 5368 7280 5432
rect 7200 5360 7280 5368
rect 7360 5752 7440 5760
rect 7360 5688 7368 5752
rect 7432 5688 7440 5752
rect 7360 5592 7440 5688
rect 7360 5528 7368 5592
rect 7432 5528 7440 5592
rect 7360 5432 7440 5528
rect 7360 5368 7368 5432
rect 7432 5368 7440 5432
rect 7360 5360 7440 5368
rect 7520 5752 7600 5760
rect 7520 5688 7528 5752
rect 7592 5688 7600 5752
rect 7520 5592 7600 5688
rect 7520 5528 7528 5592
rect 7592 5528 7600 5592
rect 7520 5432 7600 5528
rect 7520 5368 7528 5432
rect 7592 5368 7600 5432
rect 7520 5360 7600 5368
rect 7680 5752 7760 5760
rect 7680 5688 7688 5752
rect 7752 5688 7760 5752
rect 7680 5592 7760 5688
rect 7680 5528 7688 5592
rect 7752 5528 7760 5592
rect 7680 5432 7760 5528
rect 7680 5368 7688 5432
rect 7752 5368 7760 5432
rect 7680 5360 7760 5368
rect 7840 5752 7920 5760
rect 7840 5688 7848 5752
rect 7912 5688 7920 5752
rect 7840 5592 7920 5688
rect 7840 5528 7848 5592
rect 7912 5528 7920 5592
rect 7840 5432 7920 5528
rect 7840 5368 7848 5432
rect 7912 5368 7920 5432
rect 7840 5360 7920 5368
rect 8160 5752 8240 5760
rect 8160 5688 8168 5752
rect 8232 5688 8240 5752
rect 8160 5592 8240 5688
rect 8160 5528 8168 5592
rect 8232 5528 8240 5592
rect 8160 5432 8240 5528
rect 8160 5368 8168 5432
rect 8232 5368 8240 5432
rect 8160 5360 8240 5368
rect 320 4752 400 4800
rect 320 4688 328 4752
rect 392 4688 400 4752
rect 320 4672 400 4688
rect 320 4608 328 4672
rect 392 4608 400 4672
rect 320 4592 400 4608
rect 320 4528 328 4592
rect 392 4528 400 4592
rect 320 4512 400 4528
rect 320 4448 328 4512
rect 392 4448 400 4512
rect 320 4400 400 4448
rect 8000 3632 8080 3680
rect 8000 3568 8008 3632
rect 8072 3568 8080 3632
rect 8000 3552 8080 3568
rect 8000 3488 8008 3552
rect 8072 3488 8080 3552
rect 8000 3472 8080 3488
rect 8000 3408 8008 3472
rect 8072 3408 8080 3472
rect 8000 3392 8080 3408
rect 8000 3328 8008 3392
rect 8072 3328 8080 3392
rect 8000 3280 8080 3328
rect 0 2792 80 2800
rect 0 2728 8 2792
rect 72 2728 80 2792
rect 0 2472 80 2728
rect 0 2408 8 2472
rect 72 2408 80 2472
rect 0 2400 80 2408
rect 160 2792 240 2800
rect 160 2728 168 2792
rect 232 2728 240 2792
rect 160 2472 240 2728
rect 160 2408 168 2472
rect 232 2408 240 2472
rect 160 2400 240 2408
rect 320 2792 400 2800
rect 320 2728 328 2792
rect 392 2728 400 2792
rect 320 2472 400 2728
rect 320 2408 328 2472
rect 392 2408 400 2472
rect 320 2400 400 2408
rect 480 2792 560 2800
rect 480 2728 488 2792
rect 552 2728 560 2792
rect 480 2472 560 2728
rect 480 2408 488 2472
rect 552 2408 560 2472
rect 480 2400 560 2408
rect 640 2792 720 2800
rect 640 2728 648 2792
rect 712 2728 720 2792
rect 640 2472 720 2728
rect 640 2408 648 2472
rect 712 2408 720 2472
rect 640 2400 720 2408
rect 800 2792 880 2800
rect 800 2728 808 2792
rect 872 2728 880 2792
rect 800 2472 880 2728
rect 800 2408 808 2472
rect 872 2408 880 2472
rect 800 2400 880 2408
rect 960 2792 1040 2800
rect 960 2728 968 2792
rect 1032 2728 1040 2792
rect 960 2472 1040 2728
rect 960 2408 968 2472
rect 1032 2408 1040 2472
rect 960 2400 1040 2408
rect 1120 2792 1200 2800
rect 1120 2728 1128 2792
rect 1192 2728 1200 2792
rect 1120 2472 1200 2728
rect 1120 2408 1128 2472
rect 1192 2408 1200 2472
rect 1120 2400 1200 2408
rect 1440 2792 1520 2800
rect 1440 2728 1448 2792
rect 1512 2728 1520 2792
rect 1440 2472 1520 2728
rect 1440 2408 1448 2472
rect 1512 2408 1520 2472
rect 1440 2400 1520 2408
rect 1600 2792 1680 2800
rect 1600 2728 1608 2792
rect 1672 2728 1680 2792
rect 1600 2472 1680 2728
rect 1600 2408 1608 2472
rect 1672 2408 1680 2472
rect 1600 2400 1680 2408
rect 1760 2792 1840 2800
rect 1760 2728 1768 2792
rect 1832 2728 1840 2792
rect 1760 2472 1840 2728
rect 1760 2408 1768 2472
rect 1832 2408 1840 2472
rect 1760 2400 1840 2408
rect 1920 2792 2000 2800
rect 1920 2728 1928 2792
rect 1992 2728 2000 2792
rect 1920 2472 2000 2728
rect 1920 2408 1928 2472
rect 1992 2408 2000 2472
rect 1920 2400 2000 2408
rect 2080 2792 2160 2800
rect 2080 2728 2088 2792
rect 2152 2728 2160 2792
rect 2080 2472 2160 2728
rect 2080 2408 2088 2472
rect 2152 2408 2160 2472
rect 2080 2400 2160 2408
rect 2240 2792 2320 2800
rect 2240 2728 2248 2792
rect 2312 2728 2320 2792
rect 2240 2472 2320 2728
rect 2240 2408 2248 2472
rect 2312 2408 2320 2472
rect 2240 2400 2320 2408
rect 2400 2792 2480 2800
rect 2400 2728 2408 2792
rect 2472 2728 2480 2792
rect 2400 2472 2480 2728
rect 2400 2408 2408 2472
rect 2472 2408 2480 2472
rect 2400 2400 2480 2408
rect 2560 2792 2640 2800
rect 2560 2728 2568 2792
rect 2632 2728 2640 2792
rect 2560 2472 2640 2728
rect 2560 2408 2568 2472
rect 2632 2408 2640 2472
rect 2560 2400 2640 2408
rect 2720 2792 2800 2800
rect 2720 2728 2728 2792
rect 2792 2728 2800 2792
rect 2720 2472 2800 2728
rect 2720 2408 2728 2472
rect 2792 2408 2800 2472
rect 2720 2400 2800 2408
rect 2880 2792 2960 2800
rect 2880 2728 2888 2792
rect 2952 2728 2960 2792
rect 2880 2472 2960 2728
rect 2880 2408 2888 2472
rect 2952 2408 2960 2472
rect 2880 2400 2960 2408
rect 3040 2792 3120 2800
rect 3040 2728 3048 2792
rect 3112 2728 3120 2792
rect 3040 2472 3120 2728
rect 3040 2408 3048 2472
rect 3112 2408 3120 2472
rect 3040 2400 3120 2408
rect 3360 2792 3440 2800
rect 3360 2728 3368 2792
rect 3432 2728 3440 2792
rect 3360 2472 3440 2728
rect 3360 2408 3368 2472
rect 3432 2408 3440 2472
rect 3360 2400 3440 2408
rect 3520 2792 3600 2800
rect 3520 2728 3528 2792
rect 3592 2728 3600 2792
rect 3520 2472 3600 2728
rect 3520 2408 3528 2472
rect 3592 2408 3600 2472
rect 3520 2400 3600 2408
rect 3680 2792 3760 2800
rect 3680 2728 3688 2792
rect 3752 2728 3760 2792
rect 3680 2472 3760 2728
rect 3680 2408 3688 2472
rect 3752 2408 3760 2472
rect 3680 2400 3760 2408
rect 3840 2792 3920 2800
rect 3840 2728 3848 2792
rect 3912 2728 3920 2792
rect 3840 2472 3920 2728
rect 3840 2408 3848 2472
rect 3912 2408 3920 2472
rect 3840 2400 3920 2408
rect 4000 2792 4080 2800
rect 4000 2728 4008 2792
rect 4072 2728 4080 2792
rect 4000 2472 4080 2728
rect 4000 2408 4008 2472
rect 4072 2408 4080 2472
rect 4000 2400 4080 2408
rect 4160 2792 4240 2800
rect 4160 2728 4168 2792
rect 4232 2728 4240 2792
rect 4160 2472 4240 2728
rect 4160 2408 4168 2472
rect 4232 2408 4240 2472
rect 4160 2400 4240 2408
rect 4320 2792 4400 2800
rect 4320 2728 4328 2792
rect 4392 2728 4400 2792
rect 4320 2472 4400 2728
rect 4320 2408 4328 2472
rect 4392 2408 4400 2472
rect 4320 2400 4400 2408
rect 4480 2792 4560 2800
rect 4480 2728 4488 2792
rect 4552 2728 4560 2792
rect 4480 2472 4560 2728
rect 4480 2408 4488 2472
rect 4552 2408 4560 2472
rect 4480 2400 4560 2408
rect 4640 2792 4720 2800
rect 4640 2728 4648 2792
rect 4712 2728 4720 2792
rect 4640 2472 4720 2728
rect 4640 2408 4648 2472
rect 4712 2408 4720 2472
rect 4640 2400 4720 2408
rect 4800 2792 4880 2800
rect 4800 2728 4808 2792
rect 4872 2728 4880 2792
rect 4800 2472 4880 2728
rect 4800 2408 4808 2472
rect 4872 2408 4880 2472
rect 4800 2400 4880 2408
rect 4960 2792 5040 2800
rect 4960 2728 4968 2792
rect 5032 2728 5040 2792
rect 4960 2472 5040 2728
rect 4960 2408 4968 2472
rect 5032 2408 5040 2472
rect 4960 2400 5040 2408
rect 5280 2792 5360 2800
rect 5280 2728 5288 2792
rect 5352 2728 5360 2792
rect 5280 2472 5360 2728
rect 5280 2408 5288 2472
rect 5352 2408 5360 2472
rect 5280 2400 5360 2408
rect 5440 2792 5520 2800
rect 5440 2728 5448 2792
rect 5512 2728 5520 2792
rect 5440 2472 5520 2728
rect 5440 2408 5448 2472
rect 5512 2408 5520 2472
rect 5440 2400 5520 2408
rect 5600 2792 5680 2800
rect 5600 2728 5608 2792
rect 5672 2728 5680 2792
rect 5600 2472 5680 2728
rect 5600 2408 5608 2472
rect 5672 2408 5680 2472
rect 5600 2400 5680 2408
rect 5760 2792 5840 2800
rect 5760 2728 5768 2792
rect 5832 2728 5840 2792
rect 5760 2472 5840 2728
rect 5760 2408 5768 2472
rect 5832 2408 5840 2472
rect 5760 2400 5840 2408
rect 5920 2792 6000 2800
rect 5920 2728 5928 2792
rect 5992 2728 6000 2792
rect 5920 2472 6000 2728
rect 5920 2408 5928 2472
rect 5992 2408 6000 2472
rect 5920 2400 6000 2408
rect 6080 2792 6160 2800
rect 6080 2728 6088 2792
rect 6152 2728 6160 2792
rect 6080 2472 6160 2728
rect 6080 2408 6088 2472
rect 6152 2408 6160 2472
rect 6080 2400 6160 2408
rect 6240 2792 6320 2800
rect 6240 2728 6248 2792
rect 6312 2728 6320 2792
rect 6240 2472 6320 2728
rect 6240 2408 6248 2472
rect 6312 2408 6320 2472
rect 6240 2400 6320 2408
rect 6400 2792 6480 2800
rect 6400 2728 6408 2792
rect 6472 2728 6480 2792
rect 6400 2472 6480 2728
rect 6400 2408 6408 2472
rect 6472 2408 6480 2472
rect 6400 2400 6480 2408
rect 6560 2792 6640 2800
rect 6560 2728 6568 2792
rect 6632 2728 6640 2792
rect 6560 2472 6640 2728
rect 6560 2408 6568 2472
rect 6632 2408 6640 2472
rect 6560 2400 6640 2408
rect 6720 2792 6800 2800
rect 6720 2728 6728 2792
rect 6792 2728 6800 2792
rect 6720 2472 6800 2728
rect 6720 2408 6728 2472
rect 6792 2408 6800 2472
rect 6720 2400 6800 2408
rect 6880 2792 6960 2800
rect 6880 2728 6888 2792
rect 6952 2728 6960 2792
rect 6880 2472 6960 2728
rect 6880 2408 6888 2472
rect 6952 2408 6960 2472
rect 6880 2400 6960 2408
rect 7200 2792 7280 2800
rect 7200 2728 7208 2792
rect 7272 2728 7280 2792
rect 7200 2472 7280 2728
rect 7200 2408 7208 2472
rect 7272 2408 7280 2472
rect 7200 2400 7280 2408
rect 7360 2792 7440 2800
rect 7360 2728 7368 2792
rect 7432 2728 7440 2792
rect 7360 2472 7440 2728
rect 7360 2408 7368 2472
rect 7432 2408 7440 2472
rect 7360 2400 7440 2408
rect 7520 2792 7600 2800
rect 7520 2728 7528 2792
rect 7592 2728 7600 2792
rect 7520 2472 7600 2728
rect 7520 2408 7528 2472
rect 7592 2408 7600 2472
rect 7520 2400 7600 2408
rect 7680 2792 7760 2800
rect 7680 2728 7688 2792
rect 7752 2728 7760 2792
rect 7680 2472 7760 2728
rect 7680 2408 7688 2472
rect 7752 2408 7760 2472
rect 7680 2400 7760 2408
rect 7840 2792 7920 2800
rect 7840 2728 7848 2792
rect 7912 2728 7920 2792
rect 7840 2472 7920 2728
rect 7840 2408 7848 2472
rect 7912 2408 7920 2472
rect 7840 2400 7920 2408
rect 8000 2792 8080 2800
rect 8000 2728 8008 2792
rect 8072 2728 8080 2792
rect 8000 2472 8080 2728
rect 8000 2408 8008 2472
rect 8072 2408 8080 2472
rect 8000 2400 8080 2408
rect 8160 2792 8240 2800
rect 8160 2728 8168 2792
rect 8232 2728 8240 2792
rect 8160 2472 8240 2728
rect 8160 2408 8168 2472
rect 8232 2408 8240 2472
rect 8160 2400 8240 2408
rect 8320 2792 8400 2800
rect 8320 2728 8328 2792
rect 8392 2728 8400 2792
rect 8320 2472 8400 2728
rect 8320 2408 8328 2472
rect 8392 2408 8400 2472
rect 8320 2400 8400 2408
rect 160 1268 240 1280
rect 160 1212 172 1268
rect 228 1212 240 1268
rect 160 1112 240 1212
rect 160 1048 168 1112
rect 232 1048 240 1112
rect 160 952 240 1048
rect 160 888 168 952
rect 232 888 240 952
rect 160 792 240 888
rect 160 728 168 792
rect 232 728 240 792
rect 160 628 240 728
rect 160 572 172 628
rect 228 572 240 628
rect 160 560 240 572
rect 320 1268 400 1280
rect 320 1212 332 1268
rect 388 1212 400 1268
rect 320 1112 400 1212
rect 320 1048 328 1112
rect 392 1048 400 1112
rect 320 952 400 1048
rect 320 888 328 952
rect 392 888 400 952
rect 320 792 400 888
rect 320 728 328 792
rect 392 728 400 792
rect 320 628 400 728
rect 320 572 332 628
rect 388 572 400 628
rect 320 560 400 572
rect 480 1268 560 1280
rect 480 1212 492 1268
rect 548 1212 560 1268
rect 480 1112 560 1212
rect 480 1048 488 1112
rect 552 1048 560 1112
rect 480 952 560 1048
rect 480 888 488 952
rect 552 888 560 952
rect 480 792 560 888
rect 480 728 488 792
rect 552 728 560 792
rect 480 628 560 728
rect 480 572 492 628
rect 548 572 560 628
rect 480 560 560 572
rect 640 1268 720 1280
rect 640 1212 652 1268
rect 708 1212 720 1268
rect 640 1112 720 1212
rect 640 1048 648 1112
rect 712 1048 720 1112
rect 640 952 720 1048
rect 640 888 648 952
rect 712 888 720 952
rect 640 792 720 888
rect 640 728 648 792
rect 712 728 720 792
rect 640 628 720 728
rect 640 572 652 628
rect 708 572 720 628
rect 640 560 720 572
rect 800 1268 880 1280
rect 800 1212 812 1268
rect 868 1212 880 1268
rect 800 1112 880 1212
rect 800 1048 808 1112
rect 872 1048 880 1112
rect 800 952 880 1048
rect 800 888 808 952
rect 872 888 880 952
rect 800 792 880 888
rect 800 728 808 792
rect 872 728 880 792
rect 800 628 880 728
rect 800 572 812 628
rect 868 572 880 628
rect 800 560 880 572
rect 960 1268 1040 1280
rect 960 1212 972 1268
rect 1028 1212 1040 1268
rect 960 1112 1040 1212
rect 960 1048 968 1112
rect 1032 1048 1040 1112
rect 960 952 1040 1048
rect 960 888 968 952
rect 1032 888 1040 952
rect 960 792 1040 888
rect 960 728 968 792
rect 1032 728 1040 792
rect 960 628 1040 728
rect 960 572 972 628
rect 1028 572 1040 628
rect 960 560 1040 572
rect 1120 1268 1200 1280
rect 1120 1212 1132 1268
rect 1188 1212 1200 1268
rect 1120 1112 1200 1212
rect 1120 1048 1128 1112
rect 1192 1048 1200 1112
rect 1120 952 1200 1048
rect 1120 888 1128 952
rect 1192 888 1200 952
rect 1120 792 1200 888
rect 1120 728 1128 792
rect 1192 728 1200 792
rect 1120 628 1200 728
rect 1120 572 1132 628
rect 1188 572 1200 628
rect 1120 560 1200 572
rect 1440 1268 1520 1280
rect 1440 1212 1452 1268
rect 1508 1212 1520 1268
rect 1440 1112 1520 1212
rect 1440 1048 1448 1112
rect 1512 1048 1520 1112
rect 1440 952 1520 1048
rect 1440 888 1448 952
rect 1512 888 1520 952
rect 1440 792 1520 888
rect 1440 728 1448 792
rect 1512 728 1520 792
rect 1440 628 1520 728
rect 1440 572 1452 628
rect 1508 572 1520 628
rect 1440 560 1520 572
rect 1600 1268 1680 1280
rect 1600 1212 1612 1268
rect 1668 1212 1680 1268
rect 1600 1112 1680 1212
rect 1600 1048 1608 1112
rect 1672 1048 1680 1112
rect 1600 952 1680 1048
rect 1600 888 1608 952
rect 1672 888 1680 952
rect 1600 792 1680 888
rect 1600 728 1608 792
rect 1672 728 1680 792
rect 1600 628 1680 728
rect 1600 572 1612 628
rect 1668 572 1680 628
rect 1600 560 1680 572
rect 1760 1268 1840 1280
rect 1760 1212 1772 1268
rect 1828 1212 1840 1268
rect 1760 1112 1840 1212
rect 1760 1048 1768 1112
rect 1832 1048 1840 1112
rect 1760 952 1840 1048
rect 1760 888 1768 952
rect 1832 888 1840 952
rect 1760 792 1840 888
rect 1760 728 1768 792
rect 1832 728 1840 792
rect 1760 628 1840 728
rect 1760 572 1772 628
rect 1828 572 1840 628
rect 1760 560 1840 572
rect 1920 1268 2000 1280
rect 1920 1212 1932 1268
rect 1988 1212 2000 1268
rect 1920 1112 2000 1212
rect 1920 1048 1928 1112
rect 1992 1048 2000 1112
rect 1920 952 2000 1048
rect 1920 888 1928 952
rect 1992 888 2000 952
rect 1920 792 2000 888
rect 1920 728 1928 792
rect 1992 728 2000 792
rect 1920 628 2000 728
rect 1920 572 1932 628
rect 1988 572 2000 628
rect 1920 560 2000 572
rect 2080 1268 2160 1280
rect 2080 1212 2092 1268
rect 2148 1212 2160 1268
rect 2080 1112 2160 1212
rect 2080 1048 2088 1112
rect 2152 1048 2160 1112
rect 2080 952 2160 1048
rect 2080 888 2088 952
rect 2152 888 2160 952
rect 2080 792 2160 888
rect 2080 728 2088 792
rect 2152 728 2160 792
rect 2080 628 2160 728
rect 2080 572 2092 628
rect 2148 572 2160 628
rect 2080 560 2160 572
rect 2240 1268 2320 1280
rect 2240 1212 2252 1268
rect 2308 1212 2320 1268
rect 2240 1112 2320 1212
rect 2240 1048 2248 1112
rect 2312 1048 2320 1112
rect 2240 952 2320 1048
rect 2240 888 2248 952
rect 2312 888 2320 952
rect 2240 792 2320 888
rect 2240 728 2248 792
rect 2312 728 2320 792
rect 2240 628 2320 728
rect 2240 572 2252 628
rect 2308 572 2320 628
rect 2240 560 2320 572
rect 2400 1268 2480 1280
rect 2400 1212 2412 1268
rect 2468 1212 2480 1268
rect 2400 1112 2480 1212
rect 2400 1048 2408 1112
rect 2472 1048 2480 1112
rect 2400 952 2480 1048
rect 2400 888 2408 952
rect 2472 888 2480 952
rect 2400 792 2480 888
rect 2400 728 2408 792
rect 2472 728 2480 792
rect 2400 628 2480 728
rect 2400 572 2412 628
rect 2468 572 2480 628
rect 2400 560 2480 572
rect 2560 1268 2640 1280
rect 2560 1212 2572 1268
rect 2628 1212 2640 1268
rect 2560 1112 2640 1212
rect 2560 1048 2568 1112
rect 2632 1048 2640 1112
rect 2560 952 2640 1048
rect 2560 888 2568 952
rect 2632 888 2640 952
rect 2560 792 2640 888
rect 2560 728 2568 792
rect 2632 728 2640 792
rect 2560 628 2640 728
rect 2560 572 2572 628
rect 2628 572 2640 628
rect 2560 560 2640 572
rect 2720 1268 2800 1280
rect 2720 1212 2732 1268
rect 2788 1212 2800 1268
rect 2720 1112 2800 1212
rect 2720 1048 2728 1112
rect 2792 1048 2800 1112
rect 2720 952 2800 1048
rect 2720 888 2728 952
rect 2792 888 2800 952
rect 2720 792 2800 888
rect 2720 728 2728 792
rect 2792 728 2800 792
rect 2720 628 2800 728
rect 2720 572 2732 628
rect 2788 572 2800 628
rect 2720 560 2800 572
rect 2880 1268 2960 1280
rect 2880 1212 2892 1268
rect 2948 1212 2960 1268
rect 2880 1112 2960 1212
rect 2880 1048 2888 1112
rect 2952 1048 2960 1112
rect 2880 952 2960 1048
rect 2880 888 2888 952
rect 2952 888 2960 952
rect 2880 792 2960 888
rect 2880 728 2888 792
rect 2952 728 2960 792
rect 2880 628 2960 728
rect 2880 572 2892 628
rect 2948 572 2960 628
rect 2880 560 2960 572
rect 3040 1268 3120 1280
rect 3040 1212 3052 1268
rect 3108 1212 3120 1268
rect 3040 1112 3120 1212
rect 3040 1048 3048 1112
rect 3112 1048 3120 1112
rect 3040 952 3120 1048
rect 3040 888 3048 952
rect 3112 888 3120 952
rect 3040 792 3120 888
rect 3040 728 3048 792
rect 3112 728 3120 792
rect 3040 628 3120 728
rect 3040 572 3052 628
rect 3108 572 3120 628
rect 3040 560 3120 572
rect 3360 1268 3440 1280
rect 3360 1212 3372 1268
rect 3428 1212 3440 1268
rect 3360 1112 3440 1212
rect 3360 1048 3368 1112
rect 3432 1048 3440 1112
rect 3360 952 3440 1048
rect 3360 888 3368 952
rect 3432 888 3440 952
rect 3360 792 3440 888
rect 3360 728 3368 792
rect 3432 728 3440 792
rect 3360 628 3440 728
rect 3360 572 3372 628
rect 3428 572 3440 628
rect 3360 560 3440 572
rect 3520 1268 3600 1280
rect 3520 1212 3532 1268
rect 3588 1212 3600 1268
rect 3520 1112 3600 1212
rect 3520 1048 3528 1112
rect 3592 1048 3600 1112
rect 3520 952 3600 1048
rect 3520 888 3528 952
rect 3592 888 3600 952
rect 3520 792 3600 888
rect 3520 728 3528 792
rect 3592 728 3600 792
rect 3520 628 3600 728
rect 3520 572 3532 628
rect 3588 572 3600 628
rect 3520 560 3600 572
rect 3680 1268 3760 1280
rect 3680 1212 3692 1268
rect 3748 1212 3760 1268
rect 3680 1112 3760 1212
rect 3680 1048 3688 1112
rect 3752 1048 3760 1112
rect 3680 952 3760 1048
rect 3680 888 3688 952
rect 3752 888 3760 952
rect 3680 792 3760 888
rect 3680 728 3688 792
rect 3752 728 3760 792
rect 3680 628 3760 728
rect 3680 572 3692 628
rect 3748 572 3760 628
rect 3680 560 3760 572
rect 3840 1268 3920 1280
rect 3840 1212 3852 1268
rect 3908 1212 3920 1268
rect 3840 1112 3920 1212
rect 3840 1048 3848 1112
rect 3912 1048 3920 1112
rect 3840 952 3920 1048
rect 3840 888 3848 952
rect 3912 888 3920 952
rect 3840 792 3920 888
rect 3840 728 3848 792
rect 3912 728 3920 792
rect 3840 628 3920 728
rect 3840 572 3852 628
rect 3908 572 3920 628
rect 3840 560 3920 572
rect 4000 1268 4080 1280
rect 4000 1212 4012 1268
rect 4068 1212 4080 1268
rect 4000 1112 4080 1212
rect 4000 1048 4008 1112
rect 4072 1048 4080 1112
rect 4000 952 4080 1048
rect 4000 888 4008 952
rect 4072 888 4080 952
rect 4000 792 4080 888
rect 4000 728 4008 792
rect 4072 728 4080 792
rect 4000 628 4080 728
rect 4000 572 4012 628
rect 4068 572 4080 628
rect 4000 560 4080 572
rect 4160 1268 4240 1280
rect 4160 1212 4172 1268
rect 4228 1212 4240 1268
rect 4160 1112 4240 1212
rect 4160 1048 4168 1112
rect 4232 1048 4240 1112
rect 4160 952 4240 1048
rect 4160 888 4168 952
rect 4232 888 4240 952
rect 4160 792 4240 888
rect 4160 728 4168 792
rect 4232 728 4240 792
rect 4160 628 4240 728
rect 4160 572 4172 628
rect 4228 572 4240 628
rect 4160 560 4240 572
rect 4320 1268 4400 1280
rect 4320 1212 4332 1268
rect 4388 1212 4400 1268
rect 4320 1112 4400 1212
rect 4320 1048 4328 1112
rect 4392 1048 4400 1112
rect 4320 952 4400 1048
rect 4320 888 4328 952
rect 4392 888 4400 952
rect 4320 792 4400 888
rect 4320 728 4328 792
rect 4392 728 4400 792
rect 4320 628 4400 728
rect 4320 572 4332 628
rect 4388 572 4400 628
rect 4320 560 4400 572
rect 4480 1268 4560 1280
rect 4480 1212 4492 1268
rect 4548 1212 4560 1268
rect 4480 1112 4560 1212
rect 4480 1048 4488 1112
rect 4552 1048 4560 1112
rect 4480 952 4560 1048
rect 4480 888 4488 952
rect 4552 888 4560 952
rect 4480 792 4560 888
rect 4480 728 4488 792
rect 4552 728 4560 792
rect 4480 628 4560 728
rect 4480 572 4492 628
rect 4548 572 4560 628
rect 4480 560 4560 572
rect 4640 1268 4720 1280
rect 4640 1212 4652 1268
rect 4708 1212 4720 1268
rect 4640 1112 4720 1212
rect 4640 1048 4648 1112
rect 4712 1048 4720 1112
rect 4640 952 4720 1048
rect 4640 888 4648 952
rect 4712 888 4720 952
rect 4640 792 4720 888
rect 4640 728 4648 792
rect 4712 728 4720 792
rect 4640 628 4720 728
rect 4640 572 4652 628
rect 4708 572 4720 628
rect 4640 560 4720 572
rect 4800 1268 4880 1280
rect 4800 1212 4812 1268
rect 4868 1212 4880 1268
rect 4800 1112 4880 1212
rect 4800 1048 4808 1112
rect 4872 1048 4880 1112
rect 4800 952 4880 1048
rect 4800 888 4808 952
rect 4872 888 4880 952
rect 4800 792 4880 888
rect 4800 728 4808 792
rect 4872 728 4880 792
rect 4800 628 4880 728
rect 4800 572 4812 628
rect 4868 572 4880 628
rect 4800 560 4880 572
rect 4960 1268 5040 1280
rect 4960 1212 4972 1268
rect 5028 1212 5040 1268
rect 4960 1112 5040 1212
rect 4960 1048 4968 1112
rect 5032 1048 5040 1112
rect 4960 952 5040 1048
rect 4960 888 4968 952
rect 5032 888 5040 952
rect 4960 792 5040 888
rect 4960 728 4968 792
rect 5032 728 5040 792
rect 4960 628 5040 728
rect 4960 572 4972 628
rect 5028 572 5040 628
rect 4960 560 5040 572
rect 5280 1268 5360 1280
rect 5280 1212 5292 1268
rect 5348 1212 5360 1268
rect 5280 1112 5360 1212
rect 5280 1048 5288 1112
rect 5352 1048 5360 1112
rect 5280 952 5360 1048
rect 5280 888 5288 952
rect 5352 888 5360 952
rect 5280 792 5360 888
rect 5280 728 5288 792
rect 5352 728 5360 792
rect 5280 628 5360 728
rect 5280 572 5292 628
rect 5348 572 5360 628
rect 5280 560 5360 572
rect 5440 1268 5520 1280
rect 5440 1212 5452 1268
rect 5508 1212 5520 1268
rect 5440 1112 5520 1212
rect 5440 1048 5448 1112
rect 5512 1048 5520 1112
rect 5440 952 5520 1048
rect 5440 888 5448 952
rect 5512 888 5520 952
rect 5440 792 5520 888
rect 5440 728 5448 792
rect 5512 728 5520 792
rect 5440 628 5520 728
rect 5440 572 5452 628
rect 5508 572 5520 628
rect 5440 560 5520 572
rect 5600 1268 5680 1280
rect 5600 1212 5612 1268
rect 5668 1212 5680 1268
rect 5600 1112 5680 1212
rect 5600 1048 5608 1112
rect 5672 1048 5680 1112
rect 5600 952 5680 1048
rect 5600 888 5608 952
rect 5672 888 5680 952
rect 5600 792 5680 888
rect 5600 728 5608 792
rect 5672 728 5680 792
rect 5600 628 5680 728
rect 5600 572 5612 628
rect 5668 572 5680 628
rect 5600 560 5680 572
rect 5760 1268 5840 1280
rect 5760 1212 5772 1268
rect 5828 1212 5840 1268
rect 5760 1112 5840 1212
rect 5760 1048 5768 1112
rect 5832 1048 5840 1112
rect 5760 952 5840 1048
rect 5760 888 5768 952
rect 5832 888 5840 952
rect 5760 792 5840 888
rect 5760 728 5768 792
rect 5832 728 5840 792
rect 5760 628 5840 728
rect 5760 572 5772 628
rect 5828 572 5840 628
rect 5760 560 5840 572
rect 5920 1268 6000 1280
rect 5920 1212 5932 1268
rect 5988 1212 6000 1268
rect 5920 1112 6000 1212
rect 5920 1048 5928 1112
rect 5992 1048 6000 1112
rect 5920 952 6000 1048
rect 5920 888 5928 952
rect 5992 888 6000 952
rect 5920 792 6000 888
rect 5920 728 5928 792
rect 5992 728 6000 792
rect 5920 628 6000 728
rect 5920 572 5932 628
rect 5988 572 6000 628
rect 5920 560 6000 572
rect 6080 1268 6160 1280
rect 6080 1212 6092 1268
rect 6148 1212 6160 1268
rect 6080 1112 6160 1212
rect 6080 1048 6088 1112
rect 6152 1048 6160 1112
rect 6080 952 6160 1048
rect 6080 888 6088 952
rect 6152 888 6160 952
rect 6080 792 6160 888
rect 6080 728 6088 792
rect 6152 728 6160 792
rect 6080 628 6160 728
rect 6080 572 6092 628
rect 6148 572 6160 628
rect 6080 560 6160 572
rect 6240 1268 6320 1280
rect 6240 1212 6252 1268
rect 6308 1212 6320 1268
rect 6240 1112 6320 1212
rect 6240 1048 6248 1112
rect 6312 1048 6320 1112
rect 6240 952 6320 1048
rect 6240 888 6248 952
rect 6312 888 6320 952
rect 6240 792 6320 888
rect 6240 728 6248 792
rect 6312 728 6320 792
rect 6240 628 6320 728
rect 6240 572 6252 628
rect 6308 572 6320 628
rect 6240 560 6320 572
rect 6400 1268 6480 1280
rect 6400 1212 6412 1268
rect 6468 1212 6480 1268
rect 6400 1112 6480 1212
rect 6400 1048 6408 1112
rect 6472 1048 6480 1112
rect 6400 952 6480 1048
rect 6400 888 6408 952
rect 6472 888 6480 952
rect 6400 792 6480 888
rect 6400 728 6408 792
rect 6472 728 6480 792
rect 6400 628 6480 728
rect 6400 572 6412 628
rect 6468 572 6480 628
rect 6400 560 6480 572
rect 6560 1268 6640 1280
rect 6560 1212 6572 1268
rect 6628 1212 6640 1268
rect 6560 1112 6640 1212
rect 6560 1048 6568 1112
rect 6632 1048 6640 1112
rect 6560 952 6640 1048
rect 6560 888 6568 952
rect 6632 888 6640 952
rect 6560 792 6640 888
rect 6560 728 6568 792
rect 6632 728 6640 792
rect 6560 628 6640 728
rect 6560 572 6572 628
rect 6628 572 6640 628
rect 6560 560 6640 572
rect 6720 1268 6800 1280
rect 6720 1212 6732 1268
rect 6788 1212 6800 1268
rect 6720 1112 6800 1212
rect 6720 1048 6728 1112
rect 6792 1048 6800 1112
rect 6720 952 6800 1048
rect 6720 888 6728 952
rect 6792 888 6800 952
rect 6720 792 6800 888
rect 6720 728 6728 792
rect 6792 728 6800 792
rect 6720 628 6800 728
rect 6720 572 6732 628
rect 6788 572 6800 628
rect 6720 560 6800 572
rect 6880 1268 6960 1280
rect 6880 1212 6892 1268
rect 6948 1212 6960 1268
rect 6880 1112 6960 1212
rect 6880 1048 6888 1112
rect 6952 1048 6960 1112
rect 6880 952 6960 1048
rect 6880 888 6888 952
rect 6952 888 6960 952
rect 6880 792 6960 888
rect 6880 728 6888 792
rect 6952 728 6960 792
rect 6880 628 6960 728
rect 6880 572 6892 628
rect 6948 572 6960 628
rect 6880 560 6960 572
rect 7200 1268 7280 1280
rect 7200 1212 7212 1268
rect 7268 1212 7280 1268
rect 7200 1112 7280 1212
rect 7200 1048 7208 1112
rect 7272 1048 7280 1112
rect 7200 952 7280 1048
rect 7200 888 7208 952
rect 7272 888 7280 952
rect 7200 792 7280 888
rect 7200 728 7208 792
rect 7272 728 7280 792
rect 7200 628 7280 728
rect 7200 572 7212 628
rect 7268 572 7280 628
rect 7200 560 7280 572
rect 7360 1268 7440 1280
rect 7360 1212 7372 1268
rect 7428 1212 7440 1268
rect 7360 1112 7440 1212
rect 7360 1048 7368 1112
rect 7432 1048 7440 1112
rect 7360 952 7440 1048
rect 7360 888 7368 952
rect 7432 888 7440 952
rect 7360 792 7440 888
rect 7360 728 7368 792
rect 7432 728 7440 792
rect 7360 628 7440 728
rect 7360 572 7372 628
rect 7428 572 7440 628
rect 7360 560 7440 572
rect 7520 1268 7600 1280
rect 7520 1212 7532 1268
rect 7588 1212 7600 1268
rect 7520 1112 7600 1212
rect 7520 1048 7528 1112
rect 7592 1048 7600 1112
rect 7520 952 7600 1048
rect 7520 888 7528 952
rect 7592 888 7600 952
rect 7520 792 7600 888
rect 7520 728 7528 792
rect 7592 728 7600 792
rect 7520 628 7600 728
rect 7520 572 7532 628
rect 7588 572 7600 628
rect 7520 560 7600 572
rect 7680 1268 7760 1280
rect 7680 1212 7692 1268
rect 7748 1212 7760 1268
rect 7680 1112 7760 1212
rect 7680 1048 7688 1112
rect 7752 1048 7760 1112
rect 7680 952 7760 1048
rect 7680 888 7688 952
rect 7752 888 7760 952
rect 7680 792 7760 888
rect 7680 728 7688 792
rect 7752 728 7760 792
rect 7680 628 7760 728
rect 7680 572 7692 628
rect 7748 572 7760 628
rect 7680 560 7760 572
rect 7840 1268 7920 1280
rect 7840 1212 7852 1268
rect 7908 1212 7920 1268
rect 7840 1112 7920 1212
rect 8000 1268 8080 1280
rect 8000 1212 8012 1268
rect 8068 1212 8080 1268
rect 8000 1120 8080 1212
rect 8160 1268 8240 1280
rect 8160 1212 8172 1268
rect 8228 1212 8240 1268
rect 7840 1048 7848 1112
rect 7912 1048 7920 1112
rect 7840 952 7920 1048
rect 7840 888 7848 952
rect 7912 888 7920 952
rect 7840 792 7920 888
rect 7840 728 7848 792
rect 7912 728 7920 792
rect 7840 628 7920 728
rect 8160 1112 8240 1212
rect 8160 1048 8168 1112
rect 8232 1048 8240 1112
rect 8160 952 8240 1048
rect 8160 888 8168 952
rect 8232 888 8240 952
rect 8160 792 8240 888
rect 8160 728 8168 792
rect 8232 728 8240 792
rect 7840 572 7852 628
rect 7908 572 7920 628
rect 7840 560 7920 572
rect 8000 628 8080 720
rect 8000 572 8012 628
rect 8068 572 8080 628
rect 8000 560 8080 572
rect 8160 628 8240 728
rect 8160 572 8172 628
rect 8228 572 8240 628
rect 8160 560 8240 572
rect 320 332 400 360
rect 320 268 328 332
rect 392 268 400 332
rect 320 252 400 268
rect 320 188 328 252
rect 392 188 400 252
rect 320 160 400 188
rect 160 -88 240 -80
rect 160 -152 168 -88
rect 232 -152 240 -88
rect 160 -248 240 -152
rect 160 -312 168 -248
rect 232 -312 240 -248
rect 160 -408 240 -312
rect 160 -472 168 -408
rect 232 -472 240 -408
rect 160 -480 240 -472
rect 320 -88 400 -80
rect 320 -152 328 -88
rect 392 -152 400 -88
rect 320 -248 400 -152
rect 320 -312 328 -248
rect 392 -312 400 -248
rect 320 -408 400 -312
rect 320 -472 328 -408
rect 392 -472 400 -408
rect 320 -480 400 -472
rect 480 -88 560 -80
rect 480 -152 488 -88
rect 552 -152 560 -88
rect 480 -248 560 -152
rect 480 -312 488 -248
rect 552 -312 560 -248
rect 480 -408 560 -312
rect 480 -472 488 -408
rect 552 -472 560 -408
rect 480 -480 560 -472
rect 640 -88 720 -80
rect 640 -152 648 -88
rect 712 -152 720 -88
rect 640 -248 720 -152
rect 640 -312 648 -248
rect 712 -312 720 -248
rect 640 -408 720 -312
rect 640 -472 648 -408
rect 712 -472 720 -408
rect 640 -480 720 -472
rect 800 -88 880 -80
rect 800 -152 808 -88
rect 872 -152 880 -88
rect 800 -248 880 -152
rect 800 -312 808 -248
rect 872 -312 880 -248
rect 800 -408 880 -312
rect 800 -472 808 -408
rect 872 -472 880 -408
rect 800 -480 880 -472
rect 960 -88 1040 -80
rect 960 -152 968 -88
rect 1032 -152 1040 -88
rect 960 -248 1040 -152
rect 960 -312 968 -248
rect 1032 -312 1040 -248
rect 960 -408 1040 -312
rect 960 -472 968 -408
rect 1032 -472 1040 -408
rect 960 -480 1040 -472
rect 1120 -88 1200 -80
rect 1120 -152 1128 -88
rect 1192 -152 1200 -88
rect 1120 -248 1200 -152
rect 1120 -312 1128 -248
rect 1192 -312 1200 -248
rect 1120 -408 1200 -312
rect 1120 -472 1128 -408
rect 1192 -472 1200 -408
rect 1120 -480 1200 -472
rect 1440 -88 1520 -80
rect 1440 -152 1448 -88
rect 1512 -152 1520 -88
rect 1440 -248 1520 -152
rect 1440 -312 1448 -248
rect 1512 -312 1520 -248
rect 1440 -408 1520 -312
rect 1440 -472 1448 -408
rect 1512 -472 1520 -408
rect 1440 -480 1520 -472
rect 1600 -88 1680 -80
rect 1600 -152 1608 -88
rect 1672 -152 1680 -88
rect 1600 -248 1680 -152
rect 1600 -312 1608 -248
rect 1672 -312 1680 -248
rect 1600 -408 1680 -312
rect 1600 -472 1608 -408
rect 1672 -472 1680 -408
rect 1600 -480 1680 -472
rect 1760 -88 1840 -80
rect 1760 -152 1768 -88
rect 1832 -152 1840 -88
rect 1760 -248 1840 -152
rect 1760 -312 1768 -248
rect 1832 -312 1840 -248
rect 1760 -408 1840 -312
rect 1760 -472 1768 -408
rect 1832 -472 1840 -408
rect 1760 -480 1840 -472
rect 1920 -88 2000 -80
rect 1920 -152 1928 -88
rect 1992 -152 2000 -88
rect 1920 -248 2000 -152
rect 1920 -312 1928 -248
rect 1992 -312 2000 -248
rect 1920 -408 2000 -312
rect 1920 -472 1928 -408
rect 1992 -472 2000 -408
rect 1920 -480 2000 -472
rect 2080 -88 2160 -80
rect 2080 -152 2088 -88
rect 2152 -152 2160 -88
rect 2080 -248 2160 -152
rect 2080 -312 2088 -248
rect 2152 -312 2160 -248
rect 2080 -408 2160 -312
rect 2080 -472 2088 -408
rect 2152 -472 2160 -408
rect 2080 -480 2160 -472
rect 2240 -88 2320 -80
rect 2240 -152 2248 -88
rect 2312 -152 2320 -88
rect 2240 -248 2320 -152
rect 2240 -312 2248 -248
rect 2312 -312 2320 -248
rect 2240 -408 2320 -312
rect 2240 -472 2248 -408
rect 2312 -472 2320 -408
rect 2240 -480 2320 -472
rect 2400 -88 2480 -80
rect 2400 -152 2408 -88
rect 2472 -152 2480 -88
rect 2400 -248 2480 -152
rect 2400 -312 2408 -248
rect 2472 -312 2480 -248
rect 2400 -408 2480 -312
rect 2400 -472 2408 -408
rect 2472 -472 2480 -408
rect 2400 -480 2480 -472
rect 2560 -88 2640 -80
rect 2560 -152 2568 -88
rect 2632 -152 2640 -88
rect 2560 -248 2640 -152
rect 2560 -312 2568 -248
rect 2632 -312 2640 -248
rect 2560 -408 2640 -312
rect 2560 -472 2568 -408
rect 2632 -472 2640 -408
rect 2560 -480 2640 -472
rect 2720 -88 2800 -80
rect 2720 -152 2728 -88
rect 2792 -152 2800 -88
rect 2720 -248 2800 -152
rect 2720 -312 2728 -248
rect 2792 -312 2800 -248
rect 2720 -408 2800 -312
rect 2720 -472 2728 -408
rect 2792 -472 2800 -408
rect 2720 -480 2800 -472
rect 2880 -88 2960 -80
rect 2880 -152 2888 -88
rect 2952 -152 2960 -88
rect 2880 -248 2960 -152
rect 2880 -312 2888 -248
rect 2952 -312 2960 -248
rect 2880 -408 2960 -312
rect 2880 -472 2888 -408
rect 2952 -472 2960 -408
rect 2880 -480 2960 -472
rect 3040 -88 3120 -80
rect 3040 -152 3048 -88
rect 3112 -152 3120 -88
rect 3040 -248 3120 -152
rect 3040 -312 3048 -248
rect 3112 -312 3120 -248
rect 3040 -408 3120 -312
rect 3040 -472 3048 -408
rect 3112 -472 3120 -408
rect 3040 -480 3120 -472
rect 3360 -88 3440 -80
rect 3360 -152 3368 -88
rect 3432 -152 3440 -88
rect 3360 -248 3440 -152
rect 3360 -312 3368 -248
rect 3432 -312 3440 -248
rect 3360 -408 3440 -312
rect 3360 -472 3368 -408
rect 3432 -472 3440 -408
rect 3360 -480 3440 -472
rect 3520 -88 3600 -80
rect 3520 -152 3528 -88
rect 3592 -152 3600 -88
rect 3520 -248 3600 -152
rect 3520 -312 3528 -248
rect 3592 -312 3600 -248
rect 3520 -408 3600 -312
rect 3520 -472 3528 -408
rect 3592 -472 3600 -408
rect 3520 -480 3600 -472
rect 3680 -88 3760 -80
rect 3680 -152 3688 -88
rect 3752 -152 3760 -88
rect 3680 -248 3760 -152
rect 3680 -312 3688 -248
rect 3752 -312 3760 -248
rect 3680 -408 3760 -312
rect 3680 -472 3688 -408
rect 3752 -472 3760 -408
rect 3680 -480 3760 -472
rect 3840 -88 3920 -80
rect 3840 -152 3848 -88
rect 3912 -152 3920 -88
rect 3840 -248 3920 -152
rect 3840 -312 3848 -248
rect 3912 -312 3920 -248
rect 3840 -408 3920 -312
rect 3840 -472 3848 -408
rect 3912 -472 3920 -408
rect 3840 -480 3920 -472
rect 4000 -88 4080 -80
rect 4000 -152 4008 -88
rect 4072 -152 4080 -88
rect 4000 -248 4080 -152
rect 4000 -312 4008 -248
rect 4072 -312 4080 -248
rect 4000 -408 4080 -312
rect 4000 -472 4008 -408
rect 4072 -472 4080 -408
rect 4000 -480 4080 -472
rect 4160 -88 4240 -80
rect 4160 -152 4168 -88
rect 4232 -152 4240 -88
rect 4160 -248 4240 -152
rect 4160 -312 4168 -248
rect 4232 -312 4240 -248
rect 4160 -408 4240 -312
rect 4160 -472 4168 -408
rect 4232 -472 4240 -408
rect 4160 -480 4240 -472
rect 4320 -88 4400 -80
rect 4320 -152 4328 -88
rect 4392 -152 4400 -88
rect 4320 -248 4400 -152
rect 4320 -312 4328 -248
rect 4392 -312 4400 -248
rect 4320 -408 4400 -312
rect 4320 -472 4328 -408
rect 4392 -472 4400 -408
rect 4320 -480 4400 -472
rect 4480 -88 4560 -80
rect 4480 -152 4488 -88
rect 4552 -152 4560 -88
rect 4480 -248 4560 -152
rect 4480 -312 4488 -248
rect 4552 -312 4560 -248
rect 4480 -408 4560 -312
rect 4480 -472 4488 -408
rect 4552 -472 4560 -408
rect 4480 -480 4560 -472
rect 4640 -88 4720 -80
rect 4640 -152 4648 -88
rect 4712 -152 4720 -88
rect 4640 -248 4720 -152
rect 4640 -312 4648 -248
rect 4712 -312 4720 -248
rect 4640 -408 4720 -312
rect 4640 -472 4648 -408
rect 4712 -472 4720 -408
rect 4640 -480 4720 -472
rect 4800 -88 4880 -80
rect 4800 -152 4808 -88
rect 4872 -152 4880 -88
rect 4800 -248 4880 -152
rect 4800 -312 4808 -248
rect 4872 -312 4880 -248
rect 4800 -408 4880 -312
rect 4800 -472 4808 -408
rect 4872 -472 4880 -408
rect 4800 -480 4880 -472
rect 4960 -88 5040 -80
rect 4960 -152 4968 -88
rect 5032 -152 5040 -88
rect 4960 -248 5040 -152
rect 4960 -312 4968 -248
rect 5032 -312 5040 -248
rect 4960 -408 5040 -312
rect 4960 -472 4968 -408
rect 5032 -472 5040 -408
rect 4960 -480 5040 -472
rect 5280 -88 5360 -80
rect 5280 -152 5288 -88
rect 5352 -152 5360 -88
rect 5280 -248 5360 -152
rect 5280 -312 5288 -248
rect 5352 -312 5360 -248
rect 5280 -408 5360 -312
rect 5280 -472 5288 -408
rect 5352 -472 5360 -408
rect 5280 -480 5360 -472
rect 5440 -88 5520 -80
rect 5440 -152 5448 -88
rect 5512 -152 5520 -88
rect 5440 -248 5520 -152
rect 5440 -312 5448 -248
rect 5512 -312 5520 -248
rect 5440 -408 5520 -312
rect 5440 -472 5448 -408
rect 5512 -472 5520 -408
rect 5440 -480 5520 -472
rect 5600 -88 5680 -80
rect 5600 -152 5608 -88
rect 5672 -152 5680 -88
rect 5600 -248 5680 -152
rect 5600 -312 5608 -248
rect 5672 -312 5680 -248
rect 5600 -408 5680 -312
rect 5600 -472 5608 -408
rect 5672 -472 5680 -408
rect 5600 -480 5680 -472
rect 5760 -88 5840 -80
rect 5760 -152 5768 -88
rect 5832 -152 5840 -88
rect 5760 -248 5840 -152
rect 5760 -312 5768 -248
rect 5832 -312 5840 -248
rect 5760 -408 5840 -312
rect 5760 -472 5768 -408
rect 5832 -472 5840 -408
rect 5760 -480 5840 -472
rect 5920 -88 6000 -80
rect 5920 -152 5928 -88
rect 5992 -152 6000 -88
rect 5920 -248 6000 -152
rect 5920 -312 5928 -248
rect 5992 -312 6000 -248
rect 5920 -408 6000 -312
rect 5920 -472 5928 -408
rect 5992 -472 6000 -408
rect 5920 -480 6000 -472
rect 6080 -88 6160 -80
rect 6080 -152 6088 -88
rect 6152 -152 6160 -88
rect 6080 -248 6160 -152
rect 6080 -312 6088 -248
rect 6152 -312 6160 -248
rect 6080 -408 6160 -312
rect 6080 -472 6088 -408
rect 6152 -472 6160 -408
rect 6080 -480 6160 -472
rect 6240 -88 6320 -80
rect 6240 -152 6248 -88
rect 6312 -152 6320 -88
rect 6240 -248 6320 -152
rect 6240 -312 6248 -248
rect 6312 -312 6320 -248
rect 6240 -408 6320 -312
rect 6240 -472 6248 -408
rect 6312 -472 6320 -408
rect 6240 -480 6320 -472
rect 6400 -88 6480 -80
rect 6400 -152 6408 -88
rect 6472 -152 6480 -88
rect 6400 -248 6480 -152
rect 6400 -312 6408 -248
rect 6472 -312 6480 -248
rect 6400 -408 6480 -312
rect 6400 -472 6408 -408
rect 6472 -472 6480 -408
rect 6400 -480 6480 -472
rect 6560 -88 6640 -80
rect 6560 -152 6568 -88
rect 6632 -152 6640 -88
rect 6560 -248 6640 -152
rect 6560 -312 6568 -248
rect 6632 -312 6640 -248
rect 6560 -408 6640 -312
rect 6560 -472 6568 -408
rect 6632 -472 6640 -408
rect 6560 -480 6640 -472
rect 6720 -88 6800 -80
rect 6720 -152 6728 -88
rect 6792 -152 6800 -88
rect 6720 -248 6800 -152
rect 6720 -312 6728 -248
rect 6792 -312 6800 -248
rect 6720 -408 6800 -312
rect 6720 -472 6728 -408
rect 6792 -472 6800 -408
rect 6720 -480 6800 -472
rect 6880 -88 6960 -80
rect 6880 -152 6888 -88
rect 6952 -152 6960 -88
rect 6880 -248 6960 -152
rect 6880 -312 6888 -248
rect 6952 -312 6960 -248
rect 6880 -408 6960 -312
rect 6880 -472 6888 -408
rect 6952 -472 6960 -408
rect 6880 -480 6960 -472
rect 7200 -88 7280 -80
rect 7200 -152 7208 -88
rect 7272 -152 7280 -88
rect 7200 -248 7280 -152
rect 7200 -312 7208 -248
rect 7272 -312 7280 -248
rect 7200 -408 7280 -312
rect 7200 -472 7208 -408
rect 7272 -472 7280 -408
rect 7200 -480 7280 -472
rect 7360 -88 7440 -80
rect 7360 -152 7368 -88
rect 7432 -152 7440 -88
rect 7360 -248 7440 -152
rect 7360 -312 7368 -248
rect 7432 -312 7440 -248
rect 7360 -408 7440 -312
rect 7360 -472 7368 -408
rect 7432 -472 7440 -408
rect 7360 -480 7440 -472
rect 7520 -88 7600 -80
rect 7520 -152 7528 -88
rect 7592 -152 7600 -88
rect 7520 -248 7600 -152
rect 7520 -312 7528 -248
rect 7592 -312 7600 -248
rect 7520 -408 7600 -312
rect 7520 -472 7528 -408
rect 7592 -472 7600 -408
rect 7520 -480 7600 -472
rect 7680 -88 7760 -80
rect 7680 -152 7688 -88
rect 7752 -152 7760 -88
rect 7680 -248 7760 -152
rect 7680 -312 7688 -248
rect 7752 -312 7760 -248
rect 7680 -408 7760 -312
rect 7680 -472 7688 -408
rect 7752 -472 7760 -408
rect 7680 -480 7760 -472
rect 7840 -88 7920 -80
rect 7840 -152 7848 -88
rect 7912 -152 7920 -88
rect 7840 -248 7920 -152
rect 7840 -312 7848 -248
rect 7912 -312 7920 -248
rect 7840 -408 7920 -312
rect 7840 -472 7848 -408
rect 7912 -472 7920 -408
rect 7840 -480 7920 -472
rect 8160 -88 8240 -80
rect 8160 -152 8168 -88
rect 8232 -152 8240 -88
rect 8160 -248 8240 -152
rect 8160 -312 8168 -248
rect 8232 -312 8240 -248
rect 8160 -408 8240 -312
rect 8160 -472 8168 -408
rect 8232 -472 8240 -408
rect 8160 -480 8240 -472
rect 320 -708 400 -680
rect 320 -772 328 -708
rect 392 -772 400 -708
rect 320 -788 400 -772
rect 320 -852 328 -788
rect 392 -852 400 -788
rect 320 -880 400 -852
<< via3 >>
rect 328 9708 392 9712
rect 328 9652 332 9708
rect 332 9652 388 9708
rect 388 9652 392 9708
rect 328 9648 392 9652
rect 328 9628 392 9632
rect 328 9572 332 9628
rect 332 9572 388 9628
rect 388 9572 392 9628
rect 328 9568 392 9572
rect 328 9548 392 9552
rect 328 9492 332 9548
rect 332 9492 388 9548
rect 388 9492 392 9548
rect 328 9488 392 9492
rect 328 9468 392 9472
rect 328 9412 332 9468
rect 332 9412 388 9468
rect 388 9412 392 9468
rect 328 9408 392 9412
rect 168 8788 232 8792
rect 168 8732 172 8788
rect 172 8732 228 8788
rect 228 8732 232 8788
rect 168 8728 232 8732
rect 168 8568 232 8632
rect 168 8468 232 8472
rect 168 8412 172 8468
rect 172 8412 228 8468
rect 228 8412 232 8468
rect 168 8408 232 8412
rect 328 8788 392 8792
rect 328 8732 332 8788
rect 332 8732 388 8788
rect 388 8732 392 8788
rect 328 8728 392 8732
rect 328 8568 392 8632
rect 328 8468 392 8472
rect 328 8412 332 8468
rect 332 8412 388 8468
rect 388 8412 392 8468
rect 328 8408 392 8412
rect 488 8788 552 8792
rect 488 8732 492 8788
rect 492 8732 548 8788
rect 548 8732 552 8788
rect 488 8728 552 8732
rect 488 8568 552 8632
rect 488 8468 552 8472
rect 488 8412 492 8468
rect 492 8412 548 8468
rect 548 8412 552 8468
rect 488 8408 552 8412
rect 648 8788 712 8792
rect 648 8732 652 8788
rect 652 8732 708 8788
rect 708 8732 712 8788
rect 648 8728 712 8732
rect 648 8568 712 8632
rect 648 8468 712 8472
rect 648 8412 652 8468
rect 652 8412 708 8468
rect 708 8412 712 8468
rect 648 8408 712 8412
rect 808 8788 872 8792
rect 808 8732 812 8788
rect 812 8732 868 8788
rect 868 8732 872 8788
rect 808 8728 872 8732
rect 808 8568 872 8632
rect 808 8468 872 8472
rect 808 8412 812 8468
rect 812 8412 868 8468
rect 868 8412 872 8468
rect 808 8408 872 8412
rect 968 8788 1032 8792
rect 968 8732 972 8788
rect 972 8732 1028 8788
rect 1028 8732 1032 8788
rect 968 8728 1032 8732
rect 968 8568 1032 8632
rect 968 8468 1032 8472
rect 968 8412 972 8468
rect 972 8412 1028 8468
rect 1028 8412 1032 8468
rect 968 8408 1032 8412
rect 1128 8788 1192 8792
rect 1128 8732 1132 8788
rect 1132 8732 1188 8788
rect 1188 8732 1192 8788
rect 1128 8728 1192 8732
rect 1128 8568 1192 8632
rect 1128 8468 1192 8472
rect 1128 8412 1132 8468
rect 1132 8412 1188 8468
rect 1188 8412 1192 8468
rect 1128 8408 1192 8412
rect 1448 8788 1512 8792
rect 1448 8732 1452 8788
rect 1452 8732 1508 8788
rect 1508 8732 1512 8788
rect 1448 8728 1512 8732
rect 1448 8568 1512 8632
rect 1448 8468 1512 8472
rect 1448 8412 1452 8468
rect 1452 8412 1508 8468
rect 1508 8412 1512 8468
rect 1448 8408 1512 8412
rect 1608 8788 1672 8792
rect 1608 8732 1612 8788
rect 1612 8732 1668 8788
rect 1668 8732 1672 8788
rect 1608 8728 1672 8732
rect 1608 8568 1672 8632
rect 1608 8468 1672 8472
rect 1608 8412 1612 8468
rect 1612 8412 1668 8468
rect 1668 8412 1672 8468
rect 1608 8408 1672 8412
rect 1768 8788 1832 8792
rect 1768 8732 1772 8788
rect 1772 8732 1828 8788
rect 1828 8732 1832 8788
rect 1768 8728 1832 8732
rect 1768 8568 1832 8632
rect 1768 8468 1832 8472
rect 1768 8412 1772 8468
rect 1772 8412 1828 8468
rect 1828 8412 1832 8468
rect 1768 8408 1832 8412
rect 1928 8788 1992 8792
rect 1928 8732 1932 8788
rect 1932 8732 1988 8788
rect 1988 8732 1992 8788
rect 1928 8728 1992 8732
rect 1928 8568 1992 8632
rect 1928 8468 1992 8472
rect 1928 8412 1932 8468
rect 1932 8412 1988 8468
rect 1988 8412 1992 8468
rect 1928 8408 1992 8412
rect 2088 8788 2152 8792
rect 2088 8732 2092 8788
rect 2092 8732 2148 8788
rect 2148 8732 2152 8788
rect 2088 8728 2152 8732
rect 2088 8568 2152 8632
rect 2088 8468 2152 8472
rect 2088 8412 2092 8468
rect 2092 8412 2148 8468
rect 2148 8412 2152 8468
rect 2088 8408 2152 8412
rect 2248 8788 2312 8792
rect 2248 8732 2252 8788
rect 2252 8732 2308 8788
rect 2308 8732 2312 8788
rect 2248 8728 2312 8732
rect 2248 8568 2312 8632
rect 2248 8468 2312 8472
rect 2248 8412 2252 8468
rect 2252 8412 2308 8468
rect 2308 8412 2312 8468
rect 2248 8408 2312 8412
rect 2408 8788 2472 8792
rect 2408 8732 2412 8788
rect 2412 8732 2468 8788
rect 2468 8732 2472 8788
rect 2408 8728 2472 8732
rect 2408 8568 2472 8632
rect 2408 8468 2472 8472
rect 2408 8412 2412 8468
rect 2412 8412 2468 8468
rect 2468 8412 2472 8468
rect 2408 8408 2472 8412
rect 2568 8788 2632 8792
rect 2568 8732 2572 8788
rect 2572 8732 2628 8788
rect 2628 8732 2632 8788
rect 2568 8728 2632 8732
rect 2568 8568 2632 8632
rect 2568 8468 2632 8472
rect 2568 8412 2572 8468
rect 2572 8412 2628 8468
rect 2628 8412 2632 8468
rect 2568 8408 2632 8412
rect 2728 8788 2792 8792
rect 2728 8732 2732 8788
rect 2732 8732 2788 8788
rect 2788 8732 2792 8788
rect 2728 8728 2792 8732
rect 2728 8568 2792 8632
rect 2728 8468 2792 8472
rect 2728 8412 2732 8468
rect 2732 8412 2788 8468
rect 2788 8412 2792 8468
rect 2728 8408 2792 8412
rect 2888 8788 2952 8792
rect 2888 8732 2892 8788
rect 2892 8732 2948 8788
rect 2948 8732 2952 8788
rect 2888 8728 2952 8732
rect 2888 8568 2952 8632
rect 2888 8468 2952 8472
rect 2888 8412 2892 8468
rect 2892 8412 2948 8468
rect 2948 8412 2952 8468
rect 2888 8408 2952 8412
rect 3048 8788 3112 8792
rect 3048 8732 3052 8788
rect 3052 8732 3108 8788
rect 3108 8732 3112 8788
rect 3048 8728 3112 8732
rect 3048 8568 3112 8632
rect 3048 8468 3112 8472
rect 3048 8412 3052 8468
rect 3052 8412 3108 8468
rect 3108 8412 3112 8468
rect 3048 8408 3112 8412
rect 3368 8788 3432 8792
rect 3368 8732 3372 8788
rect 3372 8732 3428 8788
rect 3428 8732 3432 8788
rect 3368 8728 3432 8732
rect 3368 8568 3432 8632
rect 3368 8468 3432 8472
rect 3368 8412 3372 8468
rect 3372 8412 3428 8468
rect 3428 8412 3432 8468
rect 3368 8408 3432 8412
rect 3528 8788 3592 8792
rect 3528 8732 3532 8788
rect 3532 8732 3588 8788
rect 3588 8732 3592 8788
rect 3528 8728 3592 8732
rect 3528 8568 3592 8632
rect 3528 8468 3592 8472
rect 3528 8412 3532 8468
rect 3532 8412 3588 8468
rect 3588 8412 3592 8468
rect 3528 8408 3592 8412
rect 3688 8788 3752 8792
rect 3688 8732 3692 8788
rect 3692 8732 3748 8788
rect 3748 8732 3752 8788
rect 3688 8728 3752 8732
rect 3688 8568 3752 8632
rect 3688 8468 3752 8472
rect 3688 8412 3692 8468
rect 3692 8412 3748 8468
rect 3748 8412 3752 8468
rect 3688 8408 3752 8412
rect 3848 8788 3912 8792
rect 3848 8732 3852 8788
rect 3852 8732 3908 8788
rect 3908 8732 3912 8788
rect 3848 8728 3912 8732
rect 3848 8568 3912 8632
rect 3848 8468 3912 8472
rect 3848 8412 3852 8468
rect 3852 8412 3908 8468
rect 3908 8412 3912 8468
rect 3848 8408 3912 8412
rect 4008 8788 4072 8792
rect 4008 8732 4012 8788
rect 4012 8732 4068 8788
rect 4068 8732 4072 8788
rect 4008 8728 4072 8732
rect 4008 8568 4072 8632
rect 4008 8468 4072 8472
rect 4008 8412 4012 8468
rect 4012 8412 4068 8468
rect 4068 8412 4072 8468
rect 4008 8408 4072 8412
rect 4168 8788 4232 8792
rect 4168 8732 4172 8788
rect 4172 8732 4228 8788
rect 4228 8732 4232 8788
rect 4168 8728 4232 8732
rect 4168 8568 4232 8632
rect 4168 8468 4232 8472
rect 4168 8412 4172 8468
rect 4172 8412 4228 8468
rect 4228 8412 4232 8468
rect 4168 8408 4232 8412
rect 4328 8788 4392 8792
rect 4328 8732 4332 8788
rect 4332 8732 4388 8788
rect 4388 8732 4392 8788
rect 4328 8728 4392 8732
rect 4328 8568 4392 8632
rect 4328 8468 4392 8472
rect 4328 8412 4332 8468
rect 4332 8412 4388 8468
rect 4388 8412 4392 8468
rect 4328 8408 4392 8412
rect 4488 8788 4552 8792
rect 4488 8732 4492 8788
rect 4492 8732 4548 8788
rect 4548 8732 4552 8788
rect 4488 8728 4552 8732
rect 4488 8568 4552 8632
rect 4488 8468 4552 8472
rect 4488 8412 4492 8468
rect 4492 8412 4548 8468
rect 4548 8412 4552 8468
rect 4488 8408 4552 8412
rect 4648 8788 4712 8792
rect 4648 8732 4652 8788
rect 4652 8732 4708 8788
rect 4708 8732 4712 8788
rect 4648 8728 4712 8732
rect 4648 8568 4712 8632
rect 4648 8468 4712 8472
rect 4648 8412 4652 8468
rect 4652 8412 4708 8468
rect 4708 8412 4712 8468
rect 4648 8408 4712 8412
rect 4808 8788 4872 8792
rect 4808 8732 4812 8788
rect 4812 8732 4868 8788
rect 4868 8732 4872 8788
rect 4808 8728 4872 8732
rect 4808 8568 4872 8632
rect 4808 8468 4872 8472
rect 4808 8412 4812 8468
rect 4812 8412 4868 8468
rect 4868 8412 4872 8468
rect 4808 8408 4872 8412
rect 4968 8788 5032 8792
rect 4968 8732 4972 8788
rect 4972 8732 5028 8788
rect 5028 8732 5032 8788
rect 4968 8728 5032 8732
rect 4968 8568 5032 8632
rect 4968 8468 5032 8472
rect 4968 8412 4972 8468
rect 4972 8412 5028 8468
rect 5028 8412 5032 8468
rect 4968 8408 5032 8412
rect 5288 8788 5352 8792
rect 5288 8732 5292 8788
rect 5292 8732 5348 8788
rect 5348 8732 5352 8788
rect 5288 8728 5352 8732
rect 5288 8568 5352 8632
rect 5288 8468 5352 8472
rect 5288 8412 5292 8468
rect 5292 8412 5348 8468
rect 5348 8412 5352 8468
rect 5288 8408 5352 8412
rect 5448 8788 5512 8792
rect 5448 8732 5452 8788
rect 5452 8732 5508 8788
rect 5508 8732 5512 8788
rect 5448 8728 5512 8732
rect 5448 8568 5512 8632
rect 5448 8468 5512 8472
rect 5448 8412 5452 8468
rect 5452 8412 5508 8468
rect 5508 8412 5512 8468
rect 5448 8408 5512 8412
rect 5608 8788 5672 8792
rect 5608 8732 5612 8788
rect 5612 8732 5668 8788
rect 5668 8732 5672 8788
rect 5608 8728 5672 8732
rect 5608 8568 5672 8632
rect 5608 8468 5672 8472
rect 5608 8412 5612 8468
rect 5612 8412 5668 8468
rect 5668 8412 5672 8468
rect 5608 8408 5672 8412
rect 5768 8788 5832 8792
rect 5768 8732 5772 8788
rect 5772 8732 5828 8788
rect 5828 8732 5832 8788
rect 5768 8728 5832 8732
rect 5768 8568 5832 8632
rect 5768 8468 5832 8472
rect 5768 8412 5772 8468
rect 5772 8412 5828 8468
rect 5828 8412 5832 8468
rect 5768 8408 5832 8412
rect 5928 8788 5992 8792
rect 5928 8732 5932 8788
rect 5932 8732 5988 8788
rect 5988 8732 5992 8788
rect 5928 8728 5992 8732
rect 5928 8568 5992 8632
rect 5928 8468 5992 8472
rect 5928 8412 5932 8468
rect 5932 8412 5988 8468
rect 5988 8412 5992 8468
rect 5928 8408 5992 8412
rect 6088 8788 6152 8792
rect 6088 8732 6092 8788
rect 6092 8732 6148 8788
rect 6148 8732 6152 8788
rect 6088 8728 6152 8732
rect 6088 8568 6152 8632
rect 6088 8468 6152 8472
rect 6088 8412 6092 8468
rect 6092 8412 6148 8468
rect 6148 8412 6152 8468
rect 6088 8408 6152 8412
rect 6248 8788 6312 8792
rect 6248 8732 6252 8788
rect 6252 8732 6308 8788
rect 6308 8732 6312 8788
rect 6248 8728 6312 8732
rect 6248 8568 6312 8632
rect 6248 8468 6312 8472
rect 6248 8412 6252 8468
rect 6252 8412 6308 8468
rect 6308 8412 6312 8468
rect 6248 8408 6312 8412
rect 6408 8788 6472 8792
rect 6408 8732 6412 8788
rect 6412 8732 6468 8788
rect 6468 8732 6472 8788
rect 6408 8728 6472 8732
rect 6408 8568 6472 8632
rect 6408 8468 6472 8472
rect 6408 8412 6412 8468
rect 6412 8412 6468 8468
rect 6468 8412 6472 8468
rect 6408 8408 6472 8412
rect 6568 8788 6632 8792
rect 6568 8732 6572 8788
rect 6572 8732 6628 8788
rect 6628 8732 6632 8788
rect 6568 8728 6632 8732
rect 6568 8568 6632 8632
rect 6568 8468 6632 8472
rect 6568 8412 6572 8468
rect 6572 8412 6628 8468
rect 6628 8412 6632 8468
rect 6568 8408 6632 8412
rect 6728 8788 6792 8792
rect 6728 8732 6732 8788
rect 6732 8732 6788 8788
rect 6788 8732 6792 8788
rect 6728 8728 6792 8732
rect 6728 8568 6792 8632
rect 6728 8468 6792 8472
rect 6728 8412 6732 8468
rect 6732 8412 6788 8468
rect 6788 8412 6792 8468
rect 6728 8408 6792 8412
rect 6888 8788 6952 8792
rect 6888 8732 6892 8788
rect 6892 8732 6948 8788
rect 6948 8732 6952 8788
rect 6888 8728 6952 8732
rect 6888 8568 6952 8632
rect 6888 8468 6952 8472
rect 6888 8412 6892 8468
rect 6892 8412 6948 8468
rect 6948 8412 6952 8468
rect 6888 8408 6952 8412
rect 7208 8788 7272 8792
rect 7208 8732 7212 8788
rect 7212 8732 7268 8788
rect 7268 8732 7272 8788
rect 7208 8728 7272 8732
rect 7208 8568 7272 8632
rect 7208 8468 7272 8472
rect 7208 8412 7212 8468
rect 7212 8412 7268 8468
rect 7268 8412 7272 8468
rect 7208 8408 7272 8412
rect 7368 8788 7432 8792
rect 7368 8732 7372 8788
rect 7372 8732 7428 8788
rect 7428 8732 7432 8788
rect 7368 8728 7432 8732
rect 7368 8568 7432 8632
rect 7368 8468 7432 8472
rect 7368 8412 7372 8468
rect 7372 8412 7428 8468
rect 7428 8412 7432 8468
rect 7368 8408 7432 8412
rect 7528 8788 7592 8792
rect 7528 8732 7532 8788
rect 7532 8732 7588 8788
rect 7588 8732 7592 8788
rect 7528 8728 7592 8732
rect 7528 8568 7592 8632
rect 7528 8468 7592 8472
rect 7528 8412 7532 8468
rect 7532 8412 7588 8468
rect 7588 8412 7592 8468
rect 7528 8408 7592 8412
rect 7688 8788 7752 8792
rect 7688 8732 7692 8788
rect 7692 8732 7748 8788
rect 7748 8732 7752 8788
rect 7688 8728 7752 8732
rect 7688 8568 7752 8632
rect 7688 8468 7752 8472
rect 7688 8412 7692 8468
rect 7692 8412 7748 8468
rect 7748 8412 7752 8468
rect 7688 8408 7752 8412
rect 7848 8788 7912 8792
rect 7848 8732 7852 8788
rect 7852 8732 7908 8788
rect 7908 8732 7912 8788
rect 7848 8728 7912 8732
rect 7848 8568 7912 8632
rect 7848 8468 7912 8472
rect 7848 8412 7852 8468
rect 7852 8412 7908 8468
rect 7908 8412 7912 8468
rect 7848 8408 7912 8412
rect 8008 8788 8072 8792
rect 8008 8732 8012 8788
rect 8012 8732 8068 8788
rect 8068 8732 8072 8788
rect 8008 8728 8072 8732
rect 8008 8568 8072 8632
rect 8008 8468 8072 8472
rect 8008 8412 8012 8468
rect 8012 8412 8068 8468
rect 8068 8412 8072 8468
rect 8008 8408 8072 8412
rect 8168 8788 8232 8792
rect 8168 8732 8172 8788
rect 8172 8732 8228 8788
rect 8228 8732 8232 8788
rect 8168 8728 8232 8732
rect 8168 8568 8232 8632
rect 8168 8468 8232 8472
rect 8168 8412 8172 8468
rect 8172 8412 8228 8468
rect 8228 8412 8232 8468
rect 8168 8408 8232 8412
rect 168 8308 232 8312
rect 168 8252 172 8308
rect 172 8252 228 8308
rect 228 8252 232 8308
rect 168 8248 232 8252
rect 168 8088 232 8152
rect 168 7988 232 7992
rect 168 7932 172 7988
rect 172 7932 228 7988
rect 228 7932 232 7988
rect 168 7928 232 7932
rect 328 8308 392 8312
rect 328 8252 332 8308
rect 332 8252 388 8308
rect 388 8252 392 8308
rect 328 8248 392 8252
rect 328 8088 392 8152
rect 328 7988 392 7992
rect 328 7932 332 7988
rect 332 7932 388 7988
rect 388 7932 392 7988
rect 328 7928 392 7932
rect 488 8308 552 8312
rect 488 8252 492 8308
rect 492 8252 548 8308
rect 548 8252 552 8308
rect 488 8248 552 8252
rect 488 8088 552 8152
rect 488 7988 552 7992
rect 488 7932 492 7988
rect 492 7932 548 7988
rect 548 7932 552 7988
rect 488 7928 552 7932
rect 648 8308 712 8312
rect 648 8252 652 8308
rect 652 8252 708 8308
rect 708 8252 712 8308
rect 648 8248 712 8252
rect 648 8088 712 8152
rect 648 7988 712 7992
rect 648 7932 652 7988
rect 652 7932 708 7988
rect 708 7932 712 7988
rect 648 7928 712 7932
rect 808 8308 872 8312
rect 808 8252 812 8308
rect 812 8252 868 8308
rect 868 8252 872 8308
rect 808 8248 872 8252
rect 808 8088 872 8152
rect 808 7988 872 7992
rect 808 7932 812 7988
rect 812 7932 868 7988
rect 868 7932 872 7988
rect 808 7928 872 7932
rect 968 8308 1032 8312
rect 968 8252 972 8308
rect 972 8252 1028 8308
rect 1028 8252 1032 8308
rect 968 8248 1032 8252
rect 968 8088 1032 8152
rect 968 7988 1032 7992
rect 968 7932 972 7988
rect 972 7932 1028 7988
rect 1028 7932 1032 7988
rect 968 7928 1032 7932
rect 1128 8308 1192 8312
rect 1128 8252 1132 8308
rect 1132 8252 1188 8308
rect 1188 8252 1192 8308
rect 1128 8248 1192 8252
rect 1128 8088 1192 8152
rect 1128 7988 1192 7992
rect 1128 7932 1132 7988
rect 1132 7932 1188 7988
rect 1188 7932 1192 7988
rect 1128 7928 1192 7932
rect 1448 8308 1512 8312
rect 1448 8252 1452 8308
rect 1452 8252 1508 8308
rect 1508 8252 1512 8308
rect 1448 8248 1512 8252
rect 1448 8088 1512 8152
rect 1448 7988 1512 7992
rect 1448 7932 1452 7988
rect 1452 7932 1508 7988
rect 1508 7932 1512 7988
rect 1448 7928 1512 7932
rect 1608 8308 1672 8312
rect 1608 8252 1612 8308
rect 1612 8252 1668 8308
rect 1668 8252 1672 8308
rect 1608 8248 1672 8252
rect 1608 8088 1672 8152
rect 1608 7988 1672 7992
rect 1608 7932 1612 7988
rect 1612 7932 1668 7988
rect 1668 7932 1672 7988
rect 1608 7928 1672 7932
rect 1768 8308 1832 8312
rect 1768 8252 1772 8308
rect 1772 8252 1828 8308
rect 1828 8252 1832 8308
rect 1768 8248 1832 8252
rect 1768 8088 1832 8152
rect 1768 7988 1832 7992
rect 1768 7932 1772 7988
rect 1772 7932 1828 7988
rect 1828 7932 1832 7988
rect 1768 7928 1832 7932
rect 1928 8308 1992 8312
rect 1928 8252 1932 8308
rect 1932 8252 1988 8308
rect 1988 8252 1992 8308
rect 1928 8248 1992 8252
rect 1928 8088 1992 8152
rect 1928 7988 1992 7992
rect 1928 7932 1932 7988
rect 1932 7932 1988 7988
rect 1988 7932 1992 7988
rect 1928 7928 1992 7932
rect 2088 8308 2152 8312
rect 2088 8252 2092 8308
rect 2092 8252 2148 8308
rect 2148 8252 2152 8308
rect 2088 8248 2152 8252
rect 2088 8088 2152 8152
rect 2088 7988 2152 7992
rect 2088 7932 2092 7988
rect 2092 7932 2148 7988
rect 2148 7932 2152 7988
rect 2088 7928 2152 7932
rect 2248 8308 2312 8312
rect 2248 8252 2252 8308
rect 2252 8252 2308 8308
rect 2308 8252 2312 8308
rect 2248 8248 2312 8252
rect 2248 8088 2312 8152
rect 2248 7988 2312 7992
rect 2248 7932 2252 7988
rect 2252 7932 2308 7988
rect 2308 7932 2312 7988
rect 2248 7928 2312 7932
rect 2408 8308 2472 8312
rect 2408 8252 2412 8308
rect 2412 8252 2468 8308
rect 2468 8252 2472 8308
rect 2408 8248 2472 8252
rect 2408 8088 2472 8152
rect 2408 7988 2472 7992
rect 2408 7932 2412 7988
rect 2412 7932 2468 7988
rect 2468 7932 2472 7988
rect 2408 7928 2472 7932
rect 2568 8308 2632 8312
rect 2568 8252 2572 8308
rect 2572 8252 2628 8308
rect 2628 8252 2632 8308
rect 2568 8248 2632 8252
rect 2568 8088 2632 8152
rect 2568 7988 2632 7992
rect 2568 7932 2572 7988
rect 2572 7932 2628 7988
rect 2628 7932 2632 7988
rect 2568 7928 2632 7932
rect 2728 8308 2792 8312
rect 2728 8252 2732 8308
rect 2732 8252 2788 8308
rect 2788 8252 2792 8308
rect 2728 8248 2792 8252
rect 2728 8088 2792 8152
rect 2728 7988 2792 7992
rect 2728 7932 2732 7988
rect 2732 7932 2788 7988
rect 2788 7932 2792 7988
rect 2728 7928 2792 7932
rect 2888 8308 2952 8312
rect 2888 8252 2892 8308
rect 2892 8252 2948 8308
rect 2948 8252 2952 8308
rect 2888 8248 2952 8252
rect 2888 8088 2952 8152
rect 2888 7988 2952 7992
rect 2888 7932 2892 7988
rect 2892 7932 2948 7988
rect 2948 7932 2952 7988
rect 2888 7928 2952 7932
rect 3048 8308 3112 8312
rect 3048 8252 3052 8308
rect 3052 8252 3108 8308
rect 3108 8252 3112 8308
rect 3048 8248 3112 8252
rect 3048 8088 3112 8152
rect 3048 7988 3112 7992
rect 3048 7932 3052 7988
rect 3052 7932 3108 7988
rect 3108 7932 3112 7988
rect 3048 7928 3112 7932
rect 3368 8308 3432 8312
rect 3368 8252 3372 8308
rect 3372 8252 3428 8308
rect 3428 8252 3432 8308
rect 3368 8248 3432 8252
rect 3368 8088 3432 8152
rect 3368 7988 3432 7992
rect 3368 7932 3372 7988
rect 3372 7932 3428 7988
rect 3428 7932 3432 7988
rect 3368 7928 3432 7932
rect 3528 8308 3592 8312
rect 3528 8252 3532 8308
rect 3532 8252 3588 8308
rect 3588 8252 3592 8308
rect 3528 8248 3592 8252
rect 3528 8088 3592 8152
rect 3528 7988 3592 7992
rect 3528 7932 3532 7988
rect 3532 7932 3588 7988
rect 3588 7932 3592 7988
rect 3528 7928 3592 7932
rect 3688 8308 3752 8312
rect 3688 8252 3692 8308
rect 3692 8252 3748 8308
rect 3748 8252 3752 8308
rect 3688 8248 3752 8252
rect 3688 8088 3752 8152
rect 3688 7988 3752 7992
rect 3688 7932 3692 7988
rect 3692 7932 3748 7988
rect 3748 7932 3752 7988
rect 3688 7928 3752 7932
rect 3848 8308 3912 8312
rect 3848 8252 3852 8308
rect 3852 8252 3908 8308
rect 3908 8252 3912 8308
rect 3848 8248 3912 8252
rect 3848 8088 3912 8152
rect 3848 7988 3912 7992
rect 3848 7932 3852 7988
rect 3852 7932 3908 7988
rect 3908 7932 3912 7988
rect 3848 7928 3912 7932
rect 4008 8308 4072 8312
rect 4008 8252 4012 8308
rect 4012 8252 4068 8308
rect 4068 8252 4072 8308
rect 4008 8248 4072 8252
rect 4008 8088 4072 8152
rect 4008 7988 4072 7992
rect 4008 7932 4012 7988
rect 4012 7932 4068 7988
rect 4068 7932 4072 7988
rect 4008 7928 4072 7932
rect 4168 8308 4232 8312
rect 4168 8252 4172 8308
rect 4172 8252 4228 8308
rect 4228 8252 4232 8308
rect 4168 8248 4232 8252
rect 4168 8088 4232 8152
rect 4168 7988 4232 7992
rect 4168 7932 4172 7988
rect 4172 7932 4228 7988
rect 4228 7932 4232 7988
rect 4168 7928 4232 7932
rect 4328 8308 4392 8312
rect 4328 8252 4332 8308
rect 4332 8252 4388 8308
rect 4388 8252 4392 8308
rect 4328 8248 4392 8252
rect 4328 8088 4392 8152
rect 4328 7988 4392 7992
rect 4328 7932 4332 7988
rect 4332 7932 4388 7988
rect 4388 7932 4392 7988
rect 4328 7928 4392 7932
rect 4488 8308 4552 8312
rect 4488 8252 4492 8308
rect 4492 8252 4548 8308
rect 4548 8252 4552 8308
rect 4488 8248 4552 8252
rect 4488 8088 4552 8152
rect 4488 7988 4552 7992
rect 4488 7932 4492 7988
rect 4492 7932 4548 7988
rect 4548 7932 4552 7988
rect 4488 7928 4552 7932
rect 4648 8308 4712 8312
rect 4648 8252 4652 8308
rect 4652 8252 4708 8308
rect 4708 8252 4712 8308
rect 4648 8248 4712 8252
rect 4648 8088 4712 8152
rect 4648 7988 4712 7992
rect 4648 7932 4652 7988
rect 4652 7932 4708 7988
rect 4708 7932 4712 7988
rect 4648 7928 4712 7932
rect 4808 8308 4872 8312
rect 4808 8252 4812 8308
rect 4812 8252 4868 8308
rect 4868 8252 4872 8308
rect 4808 8248 4872 8252
rect 4808 8088 4872 8152
rect 4808 7988 4872 7992
rect 4808 7932 4812 7988
rect 4812 7932 4868 7988
rect 4868 7932 4872 7988
rect 4808 7928 4872 7932
rect 4968 8308 5032 8312
rect 4968 8252 4972 8308
rect 4972 8252 5028 8308
rect 5028 8252 5032 8308
rect 4968 8248 5032 8252
rect 4968 8088 5032 8152
rect 4968 7988 5032 7992
rect 4968 7932 4972 7988
rect 4972 7932 5028 7988
rect 5028 7932 5032 7988
rect 4968 7928 5032 7932
rect 5288 8308 5352 8312
rect 5288 8252 5292 8308
rect 5292 8252 5348 8308
rect 5348 8252 5352 8308
rect 5288 8248 5352 8252
rect 5288 8088 5352 8152
rect 5288 7988 5352 7992
rect 5288 7932 5292 7988
rect 5292 7932 5348 7988
rect 5348 7932 5352 7988
rect 5288 7928 5352 7932
rect 5448 8308 5512 8312
rect 5448 8252 5452 8308
rect 5452 8252 5508 8308
rect 5508 8252 5512 8308
rect 5448 8248 5512 8252
rect 5448 8088 5512 8152
rect 5448 7988 5512 7992
rect 5448 7932 5452 7988
rect 5452 7932 5508 7988
rect 5508 7932 5512 7988
rect 5448 7928 5512 7932
rect 5608 8308 5672 8312
rect 5608 8252 5612 8308
rect 5612 8252 5668 8308
rect 5668 8252 5672 8308
rect 5608 8248 5672 8252
rect 5608 8088 5672 8152
rect 5608 7988 5672 7992
rect 5608 7932 5612 7988
rect 5612 7932 5668 7988
rect 5668 7932 5672 7988
rect 5608 7928 5672 7932
rect 5768 8308 5832 8312
rect 5768 8252 5772 8308
rect 5772 8252 5828 8308
rect 5828 8252 5832 8308
rect 5768 8248 5832 8252
rect 5768 8088 5832 8152
rect 5768 7988 5832 7992
rect 5768 7932 5772 7988
rect 5772 7932 5828 7988
rect 5828 7932 5832 7988
rect 5768 7928 5832 7932
rect 5928 8308 5992 8312
rect 5928 8252 5932 8308
rect 5932 8252 5988 8308
rect 5988 8252 5992 8308
rect 5928 8248 5992 8252
rect 5928 8088 5992 8152
rect 5928 7988 5992 7992
rect 5928 7932 5932 7988
rect 5932 7932 5988 7988
rect 5988 7932 5992 7988
rect 5928 7928 5992 7932
rect 6088 8308 6152 8312
rect 6088 8252 6092 8308
rect 6092 8252 6148 8308
rect 6148 8252 6152 8308
rect 6088 8248 6152 8252
rect 6088 8088 6152 8152
rect 6088 7988 6152 7992
rect 6088 7932 6092 7988
rect 6092 7932 6148 7988
rect 6148 7932 6152 7988
rect 6088 7928 6152 7932
rect 6248 8308 6312 8312
rect 6248 8252 6252 8308
rect 6252 8252 6308 8308
rect 6308 8252 6312 8308
rect 6248 8248 6312 8252
rect 6248 8088 6312 8152
rect 6248 7988 6312 7992
rect 6248 7932 6252 7988
rect 6252 7932 6308 7988
rect 6308 7932 6312 7988
rect 6248 7928 6312 7932
rect 6408 8308 6472 8312
rect 6408 8252 6412 8308
rect 6412 8252 6468 8308
rect 6468 8252 6472 8308
rect 6408 8248 6472 8252
rect 6408 8088 6472 8152
rect 6408 7988 6472 7992
rect 6408 7932 6412 7988
rect 6412 7932 6468 7988
rect 6468 7932 6472 7988
rect 6408 7928 6472 7932
rect 6568 8308 6632 8312
rect 6568 8252 6572 8308
rect 6572 8252 6628 8308
rect 6628 8252 6632 8308
rect 6568 8248 6632 8252
rect 6568 8088 6632 8152
rect 6568 7988 6632 7992
rect 6568 7932 6572 7988
rect 6572 7932 6628 7988
rect 6628 7932 6632 7988
rect 6568 7928 6632 7932
rect 6728 8308 6792 8312
rect 6728 8252 6732 8308
rect 6732 8252 6788 8308
rect 6788 8252 6792 8308
rect 6728 8248 6792 8252
rect 6728 8088 6792 8152
rect 6728 7988 6792 7992
rect 6728 7932 6732 7988
rect 6732 7932 6788 7988
rect 6788 7932 6792 7988
rect 6728 7928 6792 7932
rect 6888 8308 6952 8312
rect 6888 8252 6892 8308
rect 6892 8252 6948 8308
rect 6948 8252 6952 8308
rect 6888 8248 6952 8252
rect 6888 8088 6952 8152
rect 6888 7988 6952 7992
rect 6888 7932 6892 7988
rect 6892 7932 6948 7988
rect 6948 7932 6952 7988
rect 6888 7928 6952 7932
rect 7208 8308 7272 8312
rect 7208 8252 7212 8308
rect 7212 8252 7268 8308
rect 7268 8252 7272 8308
rect 7208 8248 7272 8252
rect 7208 8088 7272 8152
rect 7208 7988 7272 7992
rect 7208 7932 7212 7988
rect 7212 7932 7268 7988
rect 7268 7932 7272 7988
rect 7208 7928 7272 7932
rect 7368 8308 7432 8312
rect 7368 8252 7372 8308
rect 7372 8252 7428 8308
rect 7428 8252 7432 8308
rect 7368 8248 7432 8252
rect 7368 8088 7432 8152
rect 7368 7988 7432 7992
rect 7368 7932 7372 7988
rect 7372 7932 7428 7988
rect 7428 7932 7432 7988
rect 7368 7928 7432 7932
rect 7528 8308 7592 8312
rect 7528 8252 7532 8308
rect 7532 8252 7588 8308
rect 7588 8252 7592 8308
rect 7528 8248 7592 8252
rect 7528 8088 7592 8152
rect 7528 7988 7592 7992
rect 7528 7932 7532 7988
rect 7532 7932 7588 7988
rect 7588 7932 7592 7988
rect 7528 7928 7592 7932
rect 7688 8308 7752 8312
rect 7688 8252 7692 8308
rect 7692 8252 7748 8308
rect 7748 8252 7752 8308
rect 7688 8248 7752 8252
rect 7688 8088 7752 8152
rect 7688 7988 7752 7992
rect 7688 7932 7692 7988
rect 7692 7932 7748 7988
rect 7748 7932 7752 7988
rect 7688 7928 7752 7932
rect 7848 8308 7912 8312
rect 7848 8252 7852 8308
rect 7852 8252 7908 8308
rect 7908 8252 7912 8308
rect 7848 8248 7912 8252
rect 7848 8088 7912 8152
rect 7848 7988 7912 7992
rect 7848 7932 7852 7988
rect 7852 7932 7908 7988
rect 7908 7932 7912 7988
rect 7848 7928 7912 7932
rect 8008 8308 8072 8312
rect 8008 8252 8012 8308
rect 8012 8252 8068 8308
rect 8068 8252 8072 8308
rect 8008 8248 8072 8252
rect 8008 8088 8072 8152
rect 8008 7988 8072 7992
rect 8008 7932 8012 7988
rect 8012 7932 8068 7988
rect 8068 7932 8072 7988
rect 8008 7928 8072 7932
rect 8168 8308 8232 8312
rect 8168 8252 8172 8308
rect 8172 8252 8228 8308
rect 8228 8252 8232 8308
rect 8168 8248 8232 8252
rect 8168 8088 8232 8152
rect 8168 7988 8232 7992
rect 8168 7932 8172 7988
rect 8172 7932 8228 7988
rect 8228 7932 8232 7988
rect 8168 7928 8232 7932
rect 328 7688 392 7692
rect 328 7632 332 7688
rect 332 7632 388 7688
rect 388 7632 392 7688
rect 328 7628 392 7632
rect 328 7608 392 7612
rect 328 7552 332 7608
rect 332 7552 388 7608
rect 388 7552 392 7608
rect 328 7548 392 7552
rect 328 7088 392 7092
rect 328 7032 332 7088
rect 332 7032 388 7088
rect 388 7032 392 7088
rect 328 7028 392 7032
rect 328 7008 392 7012
rect 328 6952 332 7008
rect 332 6952 388 7008
rect 388 6952 392 7008
rect 328 6948 392 6952
rect 168 6708 232 6712
rect 168 6652 172 6708
rect 172 6652 228 6708
rect 228 6652 232 6708
rect 168 6648 232 6652
rect 168 6488 232 6552
rect 168 6388 232 6392
rect 168 6332 172 6388
rect 172 6332 228 6388
rect 228 6332 232 6388
rect 168 6328 232 6332
rect 328 6708 392 6712
rect 328 6652 332 6708
rect 332 6652 388 6708
rect 388 6652 392 6708
rect 328 6648 392 6652
rect 328 6488 392 6552
rect 328 6388 392 6392
rect 328 6332 332 6388
rect 332 6332 388 6388
rect 388 6332 392 6388
rect 328 6328 392 6332
rect 488 6708 552 6712
rect 488 6652 492 6708
rect 492 6652 548 6708
rect 548 6652 552 6708
rect 488 6648 552 6652
rect 488 6488 552 6552
rect 488 6388 552 6392
rect 488 6332 492 6388
rect 492 6332 548 6388
rect 548 6332 552 6388
rect 488 6328 552 6332
rect 648 6708 712 6712
rect 648 6652 652 6708
rect 652 6652 708 6708
rect 708 6652 712 6708
rect 648 6648 712 6652
rect 648 6488 712 6552
rect 648 6388 712 6392
rect 648 6332 652 6388
rect 652 6332 708 6388
rect 708 6332 712 6388
rect 648 6328 712 6332
rect 808 6708 872 6712
rect 808 6652 812 6708
rect 812 6652 868 6708
rect 868 6652 872 6708
rect 808 6648 872 6652
rect 808 6488 872 6552
rect 808 6388 872 6392
rect 808 6332 812 6388
rect 812 6332 868 6388
rect 868 6332 872 6388
rect 808 6328 872 6332
rect 968 6708 1032 6712
rect 968 6652 972 6708
rect 972 6652 1028 6708
rect 1028 6652 1032 6708
rect 968 6648 1032 6652
rect 968 6488 1032 6552
rect 968 6388 1032 6392
rect 968 6332 972 6388
rect 972 6332 1028 6388
rect 1028 6332 1032 6388
rect 968 6328 1032 6332
rect 1128 6708 1192 6712
rect 1128 6652 1132 6708
rect 1132 6652 1188 6708
rect 1188 6652 1192 6708
rect 1128 6648 1192 6652
rect 1128 6488 1192 6552
rect 1128 6388 1192 6392
rect 1128 6332 1132 6388
rect 1132 6332 1188 6388
rect 1188 6332 1192 6388
rect 1128 6328 1192 6332
rect 1448 6708 1512 6712
rect 1448 6652 1452 6708
rect 1452 6652 1508 6708
rect 1508 6652 1512 6708
rect 1448 6648 1512 6652
rect 1448 6488 1512 6552
rect 1448 6388 1512 6392
rect 1448 6332 1452 6388
rect 1452 6332 1508 6388
rect 1508 6332 1512 6388
rect 1448 6328 1512 6332
rect 1608 6708 1672 6712
rect 1608 6652 1612 6708
rect 1612 6652 1668 6708
rect 1668 6652 1672 6708
rect 1608 6648 1672 6652
rect 1608 6488 1672 6552
rect 1608 6388 1672 6392
rect 1608 6332 1612 6388
rect 1612 6332 1668 6388
rect 1668 6332 1672 6388
rect 1608 6328 1672 6332
rect 1768 6708 1832 6712
rect 1768 6652 1772 6708
rect 1772 6652 1828 6708
rect 1828 6652 1832 6708
rect 1768 6648 1832 6652
rect 1768 6488 1832 6552
rect 1768 6388 1832 6392
rect 1768 6332 1772 6388
rect 1772 6332 1828 6388
rect 1828 6332 1832 6388
rect 1768 6328 1832 6332
rect 1928 6708 1992 6712
rect 1928 6652 1932 6708
rect 1932 6652 1988 6708
rect 1988 6652 1992 6708
rect 1928 6648 1992 6652
rect 1928 6488 1992 6552
rect 1928 6388 1992 6392
rect 1928 6332 1932 6388
rect 1932 6332 1988 6388
rect 1988 6332 1992 6388
rect 1928 6328 1992 6332
rect 2088 6708 2152 6712
rect 2088 6652 2092 6708
rect 2092 6652 2148 6708
rect 2148 6652 2152 6708
rect 2088 6648 2152 6652
rect 2088 6488 2152 6552
rect 2088 6388 2152 6392
rect 2088 6332 2092 6388
rect 2092 6332 2148 6388
rect 2148 6332 2152 6388
rect 2088 6328 2152 6332
rect 2248 6708 2312 6712
rect 2248 6652 2252 6708
rect 2252 6652 2308 6708
rect 2308 6652 2312 6708
rect 2248 6648 2312 6652
rect 2248 6488 2312 6552
rect 2248 6388 2312 6392
rect 2248 6332 2252 6388
rect 2252 6332 2308 6388
rect 2308 6332 2312 6388
rect 2248 6328 2312 6332
rect 2408 6708 2472 6712
rect 2408 6652 2412 6708
rect 2412 6652 2468 6708
rect 2468 6652 2472 6708
rect 2408 6648 2472 6652
rect 2408 6488 2472 6552
rect 2408 6388 2472 6392
rect 2408 6332 2412 6388
rect 2412 6332 2468 6388
rect 2468 6332 2472 6388
rect 2408 6328 2472 6332
rect 2568 6708 2632 6712
rect 2568 6652 2572 6708
rect 2572 6652 2628 6708
rect 2628 6652 2632 6708
rect 2568 6648 2632 6652
rect 2568 6488 2632 6552
rect 2568 6388 2632 6392
rect 2568 6332 2572 6388
rect 2572 6332 2628 6388
rect 2628 6332 2632 6388
rect 2568 6328 2632 6332
rect 2728 6708 2792 6712
rect 2728 6652 2732 6708
rect 2732 6652 2788 6708
rect 2788 6652 2792 6708
rect 2728 6648 2792 6652
rect 2728 6488 2792 6552
rect 2728 6388 2792 6392
rect 2728 6332 2732 6388
rect 2732 6332 2788 6388
rect 2788 6332 2792 6388
rect 2728 6328 2792 6332
rect 2888 6708 2952 6712
rect 2888 6652 2892 6708
rect 2892 6652 2948 6708
rect 2948 6652 2952 6708
rect 2888 6648 2952 6652
rect 2888 6488 2952 6552
rect 2888 6388 2952 6392
rect 2888 6332 2892 6388
rect 2892 6332 2948 6388
rect 2948 6332 2952 6388
rect 2888 6328 2952 6332
rect 3048 6708 3112 6712
rect 3048 6652 3052 6708
rect 3052 6652 3108 6708
rect 3108 6652 3112 6708
rect 3048 6648 3112 6652
rect 3048 6488 3112 6552
rect 3048 6388 3112 6392
rect 3048 6332 3052 6388
rect 3052 6332 3108 6388
rect 3108 6332 3112 6388
rect 3048 6328 3112 6332
rect 3368 6708 3432 6712
rect 3368 6652 3372 6708
rect 3372 6652 3428 6708
rect 3428 6652 3432 6708
rect 3368 6648 3432 6652
rect 3368 6488 3432 6552
rect 3368 6388 3432 6392
rect 3368 6332 3372 6388
rect 3372 6332 3428 6388
rect 3428 6332 3432 6388
rect 3368 6328 3432 6332
rect 3528 6708 3592 6712
rect 3528 6652 3532 6708
rect 3532 6652 3588 6708
rect 3588 6652 3592 6708
rect 3528 6648 3592 6652
rect 3528 6488 3592 6552
rect 3528 6388 3592 6392
rect 3528 6332 3532 6388
rect 3532 6332 3588 6388
rect 3588 6332 3592 6388
rect 3528 6328 3592 6332
rect 3688 6708 3752 6712
rect 3688 6652 3692 6708
rect 3692 6652 3748 6708
rect 3748 6652 3752 6708
rect 3688 6648 3752 6652
rect 3688 6488 3752 6552
rect 3688 6388 3752 6392
rect 3688 6332 3692 6388
rect 3692 6332 3748 6388
rect 3748 6332 3752 6388
rect 3688 6328 3752 6332
rect 3848 6708 3912 6712
rect 3848 6652 3852 6708
rect 3852 6652 3908 6708
rect 3908 6652 3912 6708
rect 3848 6648 3912 6652
rect 3848 6488 3912 6552
rect 3848 6388 3912 6392
rect 3848 6332 3852 6388
rect 3852 6332 3908 6388
rect 3908 6332 3912 6388
rect 3848 6328 3912 6332
rect 4008 6708 4072 6712
rect 4008 6652 4012 6708
rect 4012 6652 4068 6708
rect 4068 6652 4072 6708
rect 4008 6648 4072 6652
rect 4008 6488 4072 6552
rect 4008 6388 4072 6392
rect 4008 6332 4012 6388
rect 4012 6332 4068 6388
rect 4068 6332 4072 6388
rect 4008 6328 4072 6332
rect 4168 6708 4232 6712
rect 4168 6652 4172 6708
rect 4172 6652 4228 6708
rect 4228 6652 4232 6708
rect 4168 6648 4232 6652
rect 4168 6488 4232 6552
rect 4168 6388 4232 6392
rect 4168 6332 4172 6388
rect 4172 6332 4228 6388
rect 4228 6332 4232 6388
rect 4168 6328 4232 6332
rect 4328 6708 4392 6712
rect 4328 6652 4332 6708
rect 4332 6652 4388 6708
rect 4388 6652 4392 6708
rect 4328 6648 4392 6652
rect 4328 6488 4392 6552
rect 4328 6388 4392 6392
rect 4328 6332 4332 6388
rect 4332 6332 4388 6388
rect 4388 6332 4392 6388
rect 4328 6328 4392 6332
rect 4488 6708 4552 6712
rect 4488 6652 4492 6708
rect 4492 6652 4548 6708
rect 4548 6652 4552 6708
rect 4488 6648 4552 6652
rect 4488 6488 4552 6552
rect 4488 6388 4552 6392
rect 4488 6332 4492 6388
rect 4492 6332 4548 6388
rect 4548 6332 4552 6388
rect 4488 6328 4552 6332
rect 4648 6708 4712 6712
rect 4648 6652 4652 6708
rect 4652 6652 4708 6708
rect 4708 6652 4712 6708
rect 4648 6648 4712 6652
rect 4648 6488 4712 6552
rect 4648 6388 4712 6392
rect 4648 6332 4652 6388
rect 4652 6332 4708 6388
rect 4708 6332 4712 6388
rect 4648 6328 4712 6332
rect 4808 6708 4872 6712
rect 4808 6652 4812 6708
rect 4812 6652 4868 6708
rect 4868 6652 4872 6708
rect 4808 6648 4872 6652
rect 4808 6488 4872 6552
rect 4808 6388 4872 6392
rect 4808 6332 4812 6388
rect 4812 6332 4868 6388
rect 4868 6332 4872 6388
rect 4808 6328 4872 6332
rect 4968 6708 5032 6712
rect 4968 6652 4972 6708
rect 4972 6652 5028 6708
rect 5028 6652 5032 6708
rect 4968 6648 5032 6652
rect 4968 6488 5032 6552
rect 4968 6388 5032 6392
rect 4968 6332 4972 6388
rect 4972 6332 5028 6388
rect 5028 6332 5032 6388
rect 4968 6328 5032 6332
rect 5288 6708 5352 6712
rect 5288 6652 5292 6708
rect 5292 6652 5348 6708
rect 5348 6652 5352 6708
rect 5288 6648 5352 6652
rect 5288 6488 5352 6552
rect 5288 6388 5352 6392
rect 5288 6332 5292 6388
rect 5292 6332 5348 6388
rect 5348 6332 5352 6388
rect 5288 6328 5352 6332
rect 5448 6708 5512 6712
rect 5448 6652 5452 6708
rect 5452 6652 5508 6708
rect 5508 6652 5512 6708
rect 5448 6648 5512 6652
rect 5448 6488 5512 6552
rect 5448 6388 5512 6392
rect 5448 6332 5452 6388
rect 5452 6332 5508 6388
rect 5508 6332 5512 6388
rect 5448 6328 5512 6332
rect 5608 6708 5672 6712
rect 5608 6652 5612 6708
rect 5612 6652 5668 6708
rect 5668 6652 5672 6708
rect 5608 6648 5672 6652
rect 5608 6488 5672 6552
rect 5608 6388 5672 6392
rect 5608 6332 5612 6388
rect 5612 6332 5668 6388
rect 5668 6332 5672 6388
rect 5608 6328 5672 6332
rect 5768 6708 5832 6712
rect 5768 6652 5772 6708
rect 5772 6652 5828 6708
rect 5828 6652 5832 6708
rect 5768 6648 5832 6652
rect 5768 6488 5832 6552
rect 5768 6388 5832 6392
rect 5768 6332 5772 6388
rect 5772 6332 5828 6388
rect 5828 6332 5832 6388
rect 5768 6328 5832 6332
rect 5928 6708 5992 6712
rect 5928 6652 5932 6708
rect 5932 6652 5988 6708
rect 5988 6652 5992 6708
rect 5928 6648 5992 6652
rect 5928 6488 5992 6552
rect 5928 6388 5992 6392
rect 5928 6332 5932 6388
rect 5932 6332 5988 6388
rect 5988 6332 5992 6388
rect 5928 6328 5992 6332
rect 6088 6708 6152 6712
rect 6088 6652 6092 6708
rect 6092 6652 6148 6708
rect 6148 6652 6152 6708
rect 6088 6648 6152 6652
rect 6088 6488 6152 6552
rect 6088 6388 6152 6392
rect 6088 6332 6092 6388
rect 6092 6332 6148 6388
rect 6148 6332 6152 6388
rect 6088 6328 6152 6332
rect 6248 6708 6312 6712
rect 6248 6652 6252 6708
rect 6252 6652 6308 6708
rect 6308 6652 6312 6708
rect 6248 6648 6312 6652
rect 6248 6488 6312 6552
rect 6248 6388 6312 6392
rect 6248 6332 6252 6388
rect 6252 6332 6308 6388
rect 6308 6332 6312 6388
rect 6248 6328 6312 6332
rect 6408 6708 6472 6712
rect 6408 6652 6412 6708
rect 6412 6652 6468 6708
rect 6468 6652 6472 6708
rect 6408 6648 6472 6652
rect 6408 6488 6472 6552
rect 6408 6388 6472 6392
rect 6408 6332 6412 6388
rect 6412 6332 6468 6388
rect 6468 6332 6472 6388
rect 6408 6328 6472 6332
rect 6568 6708 6632 6712
rect 6568 6652 6572 6708
rect 6572 6652 6628 6708
rect 6628 6652 6632 6708
rect 6568 6648 6632 6652
rect 6568 6488 6632 6552
rect 6568 6388 6632 6392
rect 6568 6332 6572 6388
rect 6572 6332 6628 6388
rect 6628 6332 6632 6388
rect 6568 6328 6632 6332
rect 6728 6708 6792 6712
rect 6728 6652 6732 6708
rect 6732 6652 6788 6708
rect 6788 6652 6792 6708
rect 6728 6648 6792 6652
rect 6728 6488 6792 6552
rect 6728 6388 6792 6392
rect 6728 6332 6732 6388
rect 6732 6332 6788 6388
rect 6788 6332 6792 6388
rect 6728 6328 6792 6332
rect 6888 6708 6952 6712
rect 6888 6652 6892 6708
rect 6892 6652 6948 6708
rect 6948 6652 6952 6708
rect 6888 6648 6952 6652
rect 6888 6488 6952 6552
rect 6888 6388 6952 6392
rect 6888 6332 6892 6388
rect 6892 6332 6948 6388
rect 6948 6332 6952 6388
rect 6888 6328 6952 6332
rect 7208 6708 7272 6712
rect 7208 6652 7212 6708
rect 7212 6652 7268 6708
rect 7268 6652 7272 6708
rect 7208 6648 7272 6652
rect 7208 6488 7272 6552
rect 7208 6388 7272 6392
rect 7208 6332 7212 6388
rect 7212 6332 7268 6388
rect 7268 6332 7272 6388
rect 7208 6328 7272 6332
rect 7368 6708 7432 6712
rect 7368 6652 7372 6708
rect 7372 6652 7428 6708
rect 7428 6652 7432 6708
rect 7368 6648 7432 6652
rect 7368 6488 7432 6552
rect 7368 6388 7432 6392
rect 7368 6332 7372 6388
rect 7372 6332 7428 6388
rect 7428 6332 7432 6388
rect 7368 6328 7432 6332
rect 7528 6708 7592 6712
rect 7528 6652 7532 6708
rect 7532 6652 7588 6708
rect 7588 6652 7592 6708
rect 7528 6648 7592 6652
rect 7528 6488 7592 6552
rect 7528 6388 7592 6392
rect 7528 6332 7532 6388
rect 7532 6332 7588 6388
rect 7588 6332 7592 6388
rect 7528 6328 7592 6332
rect 7688 6708 7752 6712
rect 7688 6652 7692 6708
rect 7692 6652 7748 6708
rect 7748 6652 7752 6708
rect 7688 6648 7752 6652
rect 7688 6488 7752 6552
rect 7688 6388 7752 6392
rect 7688 6332 7692 6388
rect 7692 6332 7748 6388
rect 7748 6332 7752 6388
rect 7688 6328 7752 6332
rect 7848 6708 7912 6712
rect 7848 6652 7852 6708
rect 7852 6652 7908 6708
rect 7908 6652 7912 6708
rect 7848 6648 7912 6652
rect 7848 6488 7912 6552
rect 7848 6388 7912 6392
rect 7848 6332 7852 6388
rect 7852 6332 7908 6388
rect 7908 6332 7912 6388
rect 7848 6328 7912 6332
rect 8168 6708 8232 6712
rect 8168 6652 8172 6708
rect 8172 6652 8228 6708
rect 8228 6652 8232 6708
rect 8168 6648 8232 6652
rect 8168 6488 8232 6552
rect 8168 6388 8232 6392
rect 8168 6332 8172 6388
rect 8172 6332 8228 6388
rect 8228 6332 8232 6388
rect 8168 6328 8232 6332
rect 168 6228 232 6232
rect 168 6172 172 6228
rect 172 6172 228 6228
rect 228 6172 232 6228
rect 168 6168 232 6172
rect 168 6008 232 6072
rect 168 5908 232 5912
rect 168 5852 172 5908
rect 172 5852 228 5908
rect 228 5852 232 5908
rect 168 5848 232 5852
rect 328 6228 392 6232
rect 328 6172 332 6228
rect 332 6172 388 6228
rect 388 6172 392 6228
rect 328 6168 392 6172
rect 328 6008 392 6072
rect 328 5908 392 5912
rect 328 5852 332 5908
rect 332 5852 388 5908
rect 388 5852 392 5908
rect 328 5848 392 5852
rect 488 6228 552 6232
rect 488 6172 492 6228
rect 492 6172 548 6228
rect 548 6172 552 6228
rect 488 6168 552 6172
rect 488 6008 552 6072
rect 488 5908 552 5912
rect 488 5852 492 5908
rect 492 5852 548 5908
rect 548 5852 552 5908
rect 488 5848 552 5852
rect 648 6228 712 6232
rect 648 6172 652 6228
rect 652 6172 708 6228
rect 708 6172 712 6228
rect 648 6168 712 6172
rect 648 6008 712 6072
rect 648 5908 712 5912
rect 648 5852 652 5908
rect 652 5852 708 5908
rect 708 5852 712 5908
rect 648 5848 712 5852
rect 808 6228 872 6232
rect 808 6172 812 6228
rect 812 6172 868 6228
rect 868 6172 872 6228
rect 808 6168 872 6172
rect 808 6008 872 6072
rect 808 5908 872 5912
rect 808 5852 812 5908
rect 812 5852 868 5908
rect 868 5852 872 5908
rect 808 5848 872 5852
rect 968 6228 1032 6232
rect 968 6172 972 6228
rect 972 6172 1028 6228
rect 1028 6172 1032 6228
rect 968 6168 1032 6172
rect 968 6008 1032 6072
rect 968 5908 1032 5912
rect 968 5852 972 5908
rect 972 5852 1028 5908
rect 1028 5852 1032 5908
rect 968 5848 1032 5852
rect 1128 6228 1192 6232
rect 1128 6172 1132 6228
rect 1132 6172 1188 6228
rect 1188 6172 1192 6228
rect 1128 6168 1192 6172
rect 1128 6008 1192 6072
rect 1128 5908 1192 5912
rect 1128 5852 1132 5908
rect 1132 5852 1188 5908
rect 1188 5852 1192 5908
rect 1128 5848 1192 5852
rect 1288 6228 1352 6232
rect 1288 6172 1292 6228
rect 1292 6172 1348 6228
rect 1348 6172 1352 6228
rect 1288 6168 1352 6172
rect 1288 6008 1352 6072
rect 1288 5908 1352 5912
rect 1288 5852 1292 5908
rect 1292 5852 1348 5908
rect 1348 5852 1352 5908
rect 1288 5848 1352 5852
rect 1448 6228 1512 6232
rect 1448 6172 1452 6228
rect 1452 6172 1508 6228
rect 1508 6172 1512 6228
rect 1448 6168 1512 6172
rect 1448 6008 1512 6072
rect 1448 5908 1512 5912
rect 1448 5852 1452 5908
rect 1452 5852 1508 5908
rect 1508 5852 1512 5908
rect 1448 5848 1512 5852
rect 1608 6228 1672 6232
rect 1608 6172 1612 6228
rect 1612 6172 1668 6228
rect 1668 6172 1672 6228
rect 1608 6168 1672 6172
rect 1608 6008 1672 6072
rect 1608 5908 1672 5912
rect 1608 5852 1612 5908
rect 1612 5852 1668 5908
rect 1668 5852 1672 5908
rect 1608 5848 1672 5852
rect 1768 6228 1832 6232
rect 1768 6172 1772 6228
rect 1772 6172 1828 6228
rect 1828 6172 1832 6228
rect 1768 6168 1832 6172
rect 1768 6008 1832 6072
rect 1768 5908 1832 5912
rect 1768 5852 1772 5908
rect 1772 5852 1828 5908
rect 1828 5852 1832 5908
rect 1768 5848 1832 5852
rect 1928 6228 1992 6232
rect 1928 6172 1932 6228
rect 1932 6172 1988 6228
rect 1988 6172 1992 6228
rect 1928 6168 1992 6172
rect 1928 6008 1992 6072
rect 1928 5908 1992 5912
rect 1928 5852 1932 5908
rect 1932 5852 1988 5908
rect 1988 5852 1992 5908
rect 1928 5848 1992 5852
rect 2088 6228 2152 6232
rect 2088 6172 2092 6228
rect 2092 6172 2148 6228
rect 2148 6172 2152 6228
rect 2088 6168 2152 6172
rect 2088 6008 2152 6072
rect 2088 5908 2152 5912
rect 2088 5852 2092 5908
rect 2092 5852 2148 5908
rect 2148 5852 2152 5908
rect 2088 5848 2152 5852
rect 2248 6228 2312 6232
rect 2248 6172 2252 6228
rect 2252 6172 2308 6228
rect 2308 6172 2312 6228
rect 2248 6168 2312 6172
rect 2248 6008 2312 6072
rect 2248 5908 2312 5912
rect 2248 5852 2252 5908
rect 2252 5852 2308 5908
rect 2308 5852 2312 5908
rect 2248 5848 2312 5852
rect 2408 6228 2472 6232
rect 2408 6172 2412 6228
rect 2412 6172 2468 6228
rect 2468 6172 2472 6228
rect 2408 6168 2472 6172
rect 2408 6008 2472 6072
rect 2408 5908 2472 5912
rect 2408 5852 2412 5908
rect 2412 5852 2468 5908
rect 2468 5852 2472 5908
rect 2408 5848 2472 5852
rect 2568 6228 2632 6232
rect 2568 6172 2572 6228
rect 2572 6172 2628 6228
rect 2628 6172 2632 6228
rect 2568 6168 2632 6172
rect 2568 6008 2632 6072
rect 2568 5908 2632 5912
rect 2568 5852 2572 5908
rect 2572 5852 2628 5908
rect 2628 5852 2632 5908
rect 2568 5848 2632 5852
rect 2728 6228 2792 6232
rect 2728 6172 2732 6228
rect 2732 6172 2788 6228
rect 2788 6172 2792 6228
rect 2728 6168 2792 6172
rect 2728 6008 2792 6072
rect 2728 5908 2792 5912
rect 2728 5852 2732 5908
rect 2732 5852 2788 5908
rect 2788 5852 2792 5908
rect 2728 5848 2792 5852
rect 2888 6228 2952 6232
rect 2888 6172 2892 6228
rect 2892 6172 2948 6228
rect 2948 6172 2952 6228
rect 2888 6168 2952 6172
rect 2888 6008 2952 6072
rect 2888 5908 2952 5912
rect 2888 5852 2892 5908
rect 2892 5852 2948 5908
rect 2948 5852 2952 5908
rect 2888 5848 2952 5852
rect 3048 6228 3112 6232
rect 3048 6172 3052 6228
rect 3052 6172 3108 6228
rect 3108 6172 3112 6228
rect 3048 6168 3112 6172
rect 3048 6008 3112 6072
rect 3048 5908 3112 5912
rect 3048 5852 3052 5908
rect 3052 5852 3108 5908
rect 3108 5852 3112 5908
rect 3048 5848 3112 5852
rect 3208 6228 3272 6232
rect 3208 6172 3212 6228
rect 3212 6172 3268 6228
rect 3268 6172 3272 6228
rect 3208 6168 3272 6172
rect 3208 6008 3272 6072
rect 3208 5908 3272 5912
rect 3208 5852 3212 5908
rect 3212 5852 3268 5908
rect 3268 5852 3272 5908
rect 3208 5848 3272 5852
rect 3368 6228 3432 6232
rect 3368 6172 3372 6228
rect 3372 6172 3428 6228
rect 3428 6172 3432 6228
rect 3368 6168 3432 6172
rect 3368 6008 3432 6072
rect 3368 5908 3432 5912
rect 3368 5852 3372 5908
rect 3372 5852 3428 5908
rect 3428 5852 3432 5908
rect 3368 5848 3432 5852
rect 3528 6228 3592 6232
rect 3528 6172 3532 6228
rect 3532 6172 3588 6228
rect 3588 6172 3592 6228
rect 3528 6168 3592 6172
rect 3528 6008 3592 6072
rect 3528 5908 3592 5912
rect 3528 5852 3532 5908
rect 3532 5852 3588 5908
rect 3588 5852 3592 5908
rect 3528 5848 3592 5852
rect 3688 6228 3752 6232
rect 3688 6172 3692 6228
rect 3692 6172 3748 6228
rect 3748 6172 3752 6228
rect 3688 6168 3752 6172
rect 3688 6008 3752 6072
rect 3688 5908 3752 5912
rect 3688 5852 3692 5908
rect 3692 5852 3748 5908
rect 3748 5852 3752 5908
rect 3688 5848 3752 5852
rect 3848 6228 3912 6232
rect 3848 6172 3852 6228
rect 3852 6172 3908 6228
rect 3908 6172 3912 6228
rect 3848 6168 3912 6172
rect 3848 6008 3912 6072
rect 3848 5908 3912 5912
rect 3848 5852 3852 5908
rect 3852 5852 3908 5908
rect 3908 5852 3912 5908
rect 3848 5848 3912 5852
rect 4008 6228 4072 6232
rect 4008 6172 4012 6228
rect 4012 6172 4068 6228
rect 4068 6172 4072 6228
rect 4008 6168 4072 6172
rect 4008 6008 4072 6072
rect 4008 5908 4072 5912
rect 4008 5852 4012 5908
rect 4012 5852 4068 5908
rect 4068 5852 4072 5908
rect 4008 5848 4072 5852
rect 4168 6228 4232 6232
rect 4168 6172 4172 6228
rect 4172 6172 4228 6228
rect 4228 6172 4232 6228
rect 4168 6168 4232 6172
rect 4168 6008 4232 6072
rect 4168 5908 4232 5912
rect 4168 5852 4172 5908
rect 4172 5852 4228 5908
rect 4228 5852 4232 5908
rect 4168 5848 4232 5852
rect 4328 6228 4392 6232
rect 4328 6172 4332 6228
rect 4332 6172 4388 6228
rect 4388 6172 4392 6228
rect 4328 6168 4392 6172
rect 4328 6008 4392 6072
rect 4328 5908 4392 5912
rect 4328 5852 4332 5908
rect 4332 5852 4388 5908
rect 4388 5852 4392 5908
rect 4328 5848 4392 5852
rect 4488 6228 4552 6232
rect 4488 6172 4492 6228
rect 4492 6172 4548 6228
rect 4548 6172 4552 6228
rect 4488 6168 4552 6172
rect 4488 6008 4552 6072
rect 4488 5908 4552 5912
rect 4488 5852 4492 5908
rect 4492 5852 4548 5908
rect 4548 5852 4552 5908
rect 4488 5848 4552 5852
rect 4648 6228 4712 6232
rect 4648 6172 4652 6228
rect 4652 6172 4708 6228
rect 4708 6172 4712 6228
rect 4648 6168 4712 6172
rect 4648 6008 4712 6072
rect 4648 5908 4712 5912
rect 4648 5852 4652 5908
rect 4652 5852 4708 5908
rect 4708 5852 4712 5908
rect 4648 5848 4712 5852
rect 4808 6228 4872 6232
rect 4808 6172 4812 6228
rect 4812 6172 4868 6228
rect 4868 6172 4872 6228
rect 4808 6168 4872 6172
rect 4808 6008 4872 6072
rect 4808 5908 4872 5912
rect 4808 5852 4812 5908
rect 4812 5852 4868 5908
rect 4868 5852 4872 5908
rect 4808 5848 4872 5852
rect 4968 6228 5032 6232
rect 4968 6172 4972 6228
rect 4972 6172 5028 6228
rect 5028 6172 5032 6228
rect 4968 6168 5032 6172
rect 4968 6008 5032 6072
rect 4968 5908 5032 5912
rect 4968 5852 4972 5908
rect 4972 5852 5028 5908
rect 5028 5852 5032 5908
rect 4968 5848 5032 5852
rect 5128 6228 5192 6232
rect 5128 6172 5132 6228
rect 5132 6172 5188 6228
rect 5188 6172 5192 6228
rect 5128 6168 5192 6172
rect 5128 6008 5192 6072
rect 5128 5908 5192 5912
rect 5128 5852 5132 5908
rect 5132 5852 5188 5908
rect 5188 5852 5192 5908
rect 5128 5848 5192 5852
rect 5288 6228 5352 6232
rect 5288 6172 5292 6228
rect 5292 6172 5348 6228
rect 5348 6172 5352 6228
rect 5288 6168 5352 6172
rect 5288 6008 5352 6072
rect 5288 5908 5352 5912
rect 5288 5852 5292 5908
rect 5292 5852 5348 5908
rect 5348 5852 5352 5908
rect 5288 5848 5352 5852
rect 5448 6228 5512 6232
rect 5448 6172 5452 6228
rect 5452 6172 5508 6228
rect 5508 6172 5512 6228
rect 5448 6168 5512 6172
rect 5448 6008 5512 6072
rect 5448 5908 5512 5912
rect 5448 5852 5452 5908
rect 5452 5852 5508 5908
rect 5508 5852 5512 5908
rect 5448 5848 5512 5852
rect 5608 6228 5672 6232
rect 5608 6172 5612 6228
rect 5612 6172 5668 6228
rect 5668 6172 5672 6228
rect 5608 6168 5672 6172
rect 5608 6008 5672 6072
rect 5608 5908 5672 5912
rect 5608 5852 5612 5908
rect 5612 5852 5668 5908
rect 5668 5852 5672 5908
rect 5608 5848 5672 5852
rect 5768 6228 5832 6232
rect 5768 6172 5772 6228
rect 5772 6172 5828 6228
rect 5828 6172 5832 6228
rect 5768 6168 5832 6172
rect 5768 6008 5832 6072
rect 5768 5908 5832 5912
rect 5768 5852 5772 5908
rect 5772 5852 5828 5908
rect 5828 5852 5832 5908
rect 5768 5848 5832 5852
rect 5928 6228 5992 6232
rect 5928 6172 5932 6228
rect 5932 6172 5988 6228
rect 5988 6172 5992 6228
rect 5928 6168 5992 6172
rect 5928 6008 5992 6072
rect 5928 5908 5992 5912
rect 5928 5852 5932 5908
rect 5932 5852 5988 5908
rect 5988 5852 5992 5908
rect 5928 5848 5992 5852
rect 6088 6228 6152 6232
rect 6088 6172 6092 6228
rect 6092 6172 6148 6228
rect 6148 6172 6152 6228
rect 6088 6168 6152 6172
rect 6088 6008 6152 6072
rect 6088 5908 6152 5912
rect 6088 5852 6092 5908
rect 6092 5852 6148 5908
rect 6148 5852 6152 5908
rect 6088 5848 6152 5852
rect 6248 6228 6312 6232
rect 6248 6172 6252 6228
rect 6252 6172 6308 6228
rect 6308 6172 6312 6228
rect 6248 6168 6312 6172
rect 6248 6008 6312 6072
rect 6248 5908 6312 5912
rect 6248 5852 6252 5908
rect 6252 5852 6308 5908
rect 6308 5852 6312 5908
rect 6248 5848 6312 5852
rect 6408 6228 6472 6232
rect 6408 6172 6412 6228
rect 6412 6172 6468 6228
rect 6468 6172 6472 6228
rect 6408 6168 6472 6172
rect 6408 6008 6472 6072
rect 6408 5908 6472 5912
rect 6408 5852 6412 5908
rect 6412 5852 6468 5908
rect 6468 5852 6472 5908
rect 6408 5848 6472 5852
rect 6568 6228 6632 6232
rect 6568 6172 6572 6228
rect 6572 6172 6628 6228
rect 6628 6172 6632 6228
rect 6568 6168 6632 6172
rect 6568 6008 6632 6072
rect 6568 5908 6632 5912
rect 6568 5852 6572 5908
rect 6572 5852 6628 5908
rect 6628 5852 6632 5908
rect 6568 5848 6632 5852
rect 6728 6228 6792 6232
rect 6728 6172 6732 6228
rect 6732 6172 6788 6228
rect 6788 6172 6792 6228
rect 6728 6168 6792 6172
rect 6728 6008 6792 6072
rect 6728 5908 6792 5912
rect 6728 5852 6732 5908
rect 6732 5852 6788 5908
rect 6788 5852 6792 5908
rect 6728 5848 6792 5852
rect 6888 6228 6952 6232
rect 6888 6172 6892 6228
rect 6892 6172 6948 6228
rect 6948 6172 6952 6228
rect 6888 6168 6952 6172
rect 6888 6008 6952 6072
rect 6888 5908 6952 5912
rect 6888 5852 6892 5908
rect 6892 5852 6948 5908
rect 6948 5852 6952 5908
rect 6888 5848 6952 5852
rect 7048 6228 7112 6232
rect 7048 6172 7052 6228
rect 7052 6172 7108 6228
rect 7108 6172 7112 6228
rect 7048 6168 7112 6172
rect 7048 6008 7112 6072
rect 7048 5908 7112 5912
rect 7048 5852 7052 5908
rect 7052 5852 7108 5908
rect 7108 5852 7112 5908
rect 7048 5848 7112 5852
rect 7208 6228 7272 6232
rect 7208 6172 7212 6228
rect 7212 6172 7268 6228
rect 7268 6172 7272 6228
rect 7208 6168 7272 6172
rect 7208 6008 7272 6072
rect 7208 5908 7272 5912
rect 7208 5852 7212 5908
rect 7212 5852 7268 5908
rect 7268 5852 7272 5908
rect 7208 5848 7272 5852
rect 7368 6228 7432 6232
rect 7368 6172 7372 6228
rect 7372 6172 7428 6228
rect 7428 6172 7432 6228
rect 7368 6168 7432 6172
rect 7368 6008 7432 6072
rect 7368 5908 7432 5912
rect 7368 5852 7372 5908
rect 7372 5852 7428 5908
rect 7428 5852 7432 5908
rect 7368 5848 7432 5852
rect 7528 6228 7592 6232
rect 7528 6172 7532 6228
rect 7532 6172 7588 6228
rect 7588 6172 7592 6228
rect 7528 6168 7592 6172
rect 7528 6008 7592 6072
rect 7528 5908 7592 5912
rect 7528 5852 7532 5908
rect 7532 5852 7588 5908
rect 7588 5852 7592 5908
rect 7528 5848 7592 5852
rect 7688 6228 7752 6232
rect 7688 6172 7692 6228
rect 7692 6172 7748 6228
rect 7748 6172 7752 6228
rect 7688 6168 7752 6172
rect 7688 6008 7752 6072
rect 7688 5908 7752 5912
rect 7688 5852 7692 5908
rect 7692 5852 7748 5908
rect 7748 5852 7752 5908
rect 7688 5848 7752 5852
rect 7848 6228 7912 6232
rect 7848 6172 7852 6228
rect 7852 6172 7908 6228
rect 7908 6172 7912 6228
rect 7848 6168 7912 6172
rect 7848 6008 7912 6072
rect 7848 5908 7912 5912
rect 7848 5852 7852 5908
rect 7852 5852 7908 5908
rect 7908 5852 7912 5908
rect 7848 5848 7912 5852
rect 8168 6228 8232 6232
rect 8168 6172 8172 6228
rect 8172 6172 8228 6228
rect 8228 6172 8232 6228
rect 8168 6168 8232 6172
rect 8168 6008 8232 6072
rect 8168 5908 8232 5912
rect 8168 5852 8172 5908
rect 8172 5852 8228 5908
rect 8228 5852 8232 5908
rect 8168 5848 8232 5852
rect 168 5748 232 5752
rect 168 5692 172 5748
rect 172 5692 228 5748
rect 228 5692 232 5748
rect 168 5688 232 5692
rect 168 5528 232 5592
rect 168 5428 232 5432
rect 168 5372 172 5428
rect 172 5372 228 5428
rect 228 5372 232 5428
rect 168 5368 232 5372
rect 328 5748 392 5752
rect 328 5692 332 5748
rect 332 5692 388 5748
rect 388 5692 392 5748
rect 328 5688 392 5692
rect 328 5528 392 5592
rect 328 5428 392 5432
rect 328 5372 332 5428
rect 332 5372 388 5428
rect 388 5372 392 5428
rect 328 5368 392 5372
rect 488 5748 552 5752
rect 488 5692 492 5748
rect 492 5692 548 5748
rect 548 5692 552 5748
rect 488 5688 552 5692
rect 488 5528 552 5592
rect 488 5428 552 5432
rect 488 5372 492 5428
rect 492 5372 548 5428
rect 548 5372 552 5428
rect 488 5368 552 5372
rect 648 5748 712 5752
rect 648 5692 652 5748
rect 652 5692 708 5748
rect 708 5692 712 5748
rect 648 5688 712 5692
rect 648 5528 712 5592
rect 648 5428 712 5432
rect 648 5372 652 5428
rect 652 5372 708 5428
rect 708 5372 712 5428
rect 648 5368 712 5372
rect 808 5748 872 5752
rect 808 5692 812 5748
rect 812 5692 868 5748
rect 868 5692 872 5748
rect 808 5688 872 5692
rect 808 5528 872 5592
rect 808 5428 872 5432
rect 808 5372 812 5428
rect 812 5372 868 5428
rect 868 5372 872 5428
rect 808 5368 872 5372
rect 968 5748 1032 5752
rect 968 5692 972 5748
rect 972 5692 1028 5748
rect 1028 5692 1032 5748
rect 968 5688 1032 5692
rect 968 5528 1032 5592
rect 968 5428 1032 5432
rect 968 5372 972 5428
rect 972 5372 1028 5428
rect 1028 5372 1032 5428
rect 968 5368 1032 5372
rect 1128 5748 1192 5752
rect 1128 5692 1132 5748
rect 1132 5692 1188 5748
rect 1188 5692 1192 5748
rect 1128 5688 1192 5692
rect 1128 5528 1192 5592
rect 1128 5428 1192 5432
rect 1128 5372 1132 5428
rect 1132 5372 1188 5428
rect 1188 5372 1192 5428
rect 1128 5368 1192 5372
rect 1448 5748 1512 5752
rect 1448 5692 1452 5748
rect 1452 5692 1508 5748
rect 1508 5692 1512 5748
rect 1448 5688 1512 5692
rect 1448 5528 1512 5592
rect 1448 5428 1512 5432
rect 1448 5372 1452 5428
rect 1452 5372 1508 5428
rect 1508 5372 1512 5428
rect 1448 5368 1512 5372
rect 1608 5748 1672 5752
rect 1608 5692 1612 5748
rect 1612 5692 1668 5748
rect 1668 5692 1672 5748
rect 1608 5688 1672 5692
rect 1608 5528 1672 5592
rect 1608 5428 1672 5432
rect 1608 5372 1612 5428
rect 1612 5372 1668 5428
rect 1668 5372 1672 5428
rect 1608 5368 1672 5372
rect 1768 5748 1832 5752
rect 1768 5692 1772 5748
rect 1772 5692 1828 5748
rect 1828 5692 1832 5748
rect 1768 5688 1832 5692
rect 1768 5528 1832 5592
rect 1768 5428 1832 5432
rect 1768 5372 1772 5428
rect 1772 5372 1828 5428
rect 1828 5372 1832 5428
rect 1768 5368 1832 5372
rect 1928 5748 1992 5752
rect 1928 5692 1932 5748
rect 1932 5692 1988 5748
rect 1988 5692 1992 5748
rect 1928 5688 1992 5692
rect 1928 5528 1992 5592
rect 1928 5428 1992 5432
rect 1928 5372 1932 5428
rect 1932 5372 1988 5428
rect 1988 5372 1992 5428
rect 1928 5368 1992 5372
rect 2088 5748 2152 5752
rect 2088 5692 2092 5748
rect 2092 5692 2148 5748
rect 2148 5692 2152 5748
rect 2088 5688 2152 5692
rect 2088 5528 2152 5592
rect 2088 5428 2152 5432
rect 2088 5372 2092 5428
rect 2092 5372 2148 5428
rect 2148 5372 2152 5428
rect 2088 5368 2152 5372
rect 2248 5748 2312 5752
rect 2248 5692 2252 5748
rect 2252 5692 2308 5748
rect 2308 5692 2312 5748
rect 2248 5688 2312 5692
rect 2248 5528 2312 5592
rect 2248 5428 2312 5432
rect 2248 5372 2252 5428
rect 2252 5372 2308 5428
rect 2308 5372 2312 5428
rect 2248 5368 2312 5372
rect 2408 5748 2472 5752
rect 2408 5692 2412 5748
rect 2412 5692 2468 5748
rect 2468 5692 2472 5748
rect 2408 5688 2472 5692
rect 2408 5528 2472 5592
rect 2408 5428 2472 5432
rect 2408 5372 2412 5428
rect 2412 5372 2468 5428
rect 2468 5372 2472 5428
rect 2408 5368 2472 5372
rect 2568 5748 2632 5752
rect 2568 5692 2572 5748
rect 2572 5692 2628 5748
rect 2628 5692 2632 5748
rect 2568 5688 2632 5692
rect 2568 5528 2632 5592
rect 2568 5428 2632 5432
rect 2568 5372 2572 5428
rect 2572 5372 2628 5428
rect 2628 5372 2632 5428
rect 2568 5368 2632 5372
rect 2728 5748 2792 5752
rect 2728 5692 2732 5748
rect 2732 5692 2788 5748
rect 2788 5692 2792 5748
rect 2728 5688 2792 5692
rect 2728 5528 2792 5592
rect 2728 5428 2792 5432
rect 2728 5372 2732 5428
rect 2732 5372 2788 5428
rect 2788 5372 2792 5428
rect 2728 5368 2792 5372
rect 2888 5748 2952 5752
rect 2888 5692 2892 5748
rect 2892 5692 2948 5748
rect 2948 5692 2952 5748
rect 2888 5688 2952 5692
rect 2888 5528 2952 5592
rect 2888 5428 2952 5432
rect 2888 5372 2892 5428
rect 2892 5372 2948 5428
rect 2948 5372 2952 5428
rect 2888 5368 2952 5372
rect 3048 5748 3112 5752
rect 3048 5692 3052 5748
rect 3052 5692 3108 5748
rect 3108 5692 3112 5748
rect 3048 5688 3112 5692
rect 3048 5528 3112 5592
rect 3048 5428 3112 5432
rect 3048 5372 3052 5428
rect 3052 5372 3108 5428
rect 3108 5372 3112 5428
rect 3048 5368 3112 5372
rect 3368 5748 3432 5752
rect 3368 5692 3372 5748
rect 3372 5692 3428 5748
rect 3428 5692 3432 5748
rect 3368 5688 3432 5692
rect 3368 5528 3432 5592
rect 3368 5428 3432 5432
rect 3368 5372 3372 5428
rect 3372 5372 3428 5428
rect 3428 5372 3432 5428
rect 3368 5368 3432 5372
rect 3528 5748 3592 5752
rect 3528 5692 3532 5748
rect 3532 5692 3588 5748
rect 3588 5692 3592 5748
rect 3528 5688 3592 5692
rect 3528 5528 3592 5592
rect 3528 5428 3592 5432
rect 3528 5372 3532 5428
rect 3532 5372 3588 5428
rect 3588 5372 3592 5428
rect 3528 5368 3592 5372
rect 3688 5748 3752 5752
rect 3688 5692 3692 5748
rect 3692 5692 3748 5748
rect 3748 5692 3752 5748
rect 3688 5688 3752 5692
rect 3688 5528 3752 5592
rect 3688 5428 3752 5432
rect 3688 5372 3692 5428
rect 3692 5372 3748 5428
rect 3748 5372 3752 5428
rect 3688 5368 3752 5372
rect 3848 5748 3912 5752
rect 3848 5692 3852 5748
rect 3852 5692 3908 5748
rect 3908 5692 3912 5748
rect 3848 5688 3912 5692
rect 3848 5528 3912 5592
rect 3848 5428 3912 5432
rect 3848 5372 3852 5428
rect 3852 5372 3908 5428
rect 3908 5372 3912 5428
rect 3848 5368 3912 5372
rect 4008 5748 4072 5752
rect 4008 5692 4012 5748
rect 4012 5692 4068 5748
rect 4068 5692 4072 5748
rect 4008 5688 4072 5692
rect 4008 5528 4072 5592
rect 4008 5428 4072 5432
rect 4008 5372 4012 5428
rect 4012 5372 4068 5428
rect 4068 5372 4072 5428
rect 4008 5368 4072 5372
rect 4168 5748 4232 5752
rect 4168 5692 4172 5748
rect 4172 5692 4228 5748
rect 4228 5692 4232 5748
rect 4168 5688 4232 5692
rect 4168 5528 4232 5592
rect 4168 5428 4232 5432
rect 4168 5372 4172 5428
rect 4172 5372 4228 5428
rect 4228 5372 4232 5428
rect 4168 5368 4232 5372
rect 4328 5748 4392 5752
rect 4328 5692 4332 5748
rect 4332 5692 4388 5748
rect 4388 5692 4392 5748
rect 4328 5688 4392 5692
rect 4328 5528 4392 5592
rect 4328 5428 4392 5432
rect 4328 5372 4332 5428
rect 4332 5372 4388 5428
rect 4388 5372 4392 5428
rect 4328 5368 4392 5372
rect 4488 5748 4552 5752
rect 4488 5692 4492 5748
rect 4492 5692 4548 5748
rect 4548 5692 4552 5748
rect 4488 5688 4552 5692
rect 4488 5528 4552 5592
rect 4488 5428 4552 5432
rect 4488 5372 4492 5428
rect 4492 5372 4548 5428
rect 4548 5372 4552 5428
rect 4488 5368 4552 5372
rect 4648 5748 4712 5752
rect 4648 5692 4652 5748
rect 4652 5692 4708 5748
rect 4708 5692 4712 5748
rect 4648 5688 4712 5692
rect 4648 5528 4712 5592
rect 4648 5428 4712 5432
rect 4648 5372 4652 5428
rect 4652 5372 4708 5428
rect 4708 5372 4712 5428
rect 4648 5368 4712 5372
rect 4808 5748 4872 5752
rect 4808 5692 4812 5748
rect 4812 5692 4868 5748
rect 4868 5692 4872 5748
rect 4808 5688 4872 5692
rect 4808 5528 4872 5592
rect 4808 5428 4872 5432
rect 4808 5372 4812 5428
rect 4812 5372 4868 5428
rect 4868 5372 4872 5428
rect 4808 5368 4872 5372
rect 4968 5748 5032 5752
rect 4968 5692 4972 5748
rect 4972 5692 5028 5748
rect 5028 5692 5032 5748
rect 4968 5688 5032 5692
rect 4968 5528 5032 5592
rect 4968 5428 5032 5432
rect 4968 5372 4972 5428
rect 4972 5372 5028 5428
rect 5028 5372 5032 5428
rect 4968 5368 5032 5372
rect 5288 5748 5352 5752
rect 5288 5692 5292 5748
rect 5292 5692 5348 5748
rect 5348 5692 5352 5748
rect 5288 5688 5352 5692
rect 5288 5528 5352 5592
rect 5288 5428 5352 5432
rect 5288 5372 5292 5428
rect 5292 5372 5348 5428
rect 5348 5372 5352 5428
rect 5288 5368 5352 5372
rect 5448 5748 5512 5752
rect 5448 5692 5452 5748
rect 5452 5692 5508 5748
rect 5508 5692 5512 5748
rect 5448 5688 5512 5692
rect 5448 5528 5512 5592
rect 5448 5428 5512 5432
rect 5448 5372 5452 5428
rect 5452 5372 5508 5428
rect 5508 5372 5512 5428
rect 5448 5368 5512 5372
rect 5608 5748 5672 5752
rect 5608 5692 5612 5748
rect 5612 5692 5668 5748
rect 5668 5692 5672 5748
rect 5608 5688 5672 5692
rect 5608 5528 5672 5592
rect 5608 5428 5672 5432
rect 5608 5372 5612 5428
rect 5612 5372 5668 5428
rect 5668 5372 5672 5428
rect 5608 5368 5672 5372
rect 5768 5748 5832 5752
rect 5768 5692 5772 5748
rect 5772 5692 5828 5748
rect 5828 5692 5832 5748
rect 5768 5688 5832 5692
rect 5768 5528 5832 5592
rect 5768 5428 5832 5432
rect 5768 5372 5772 5428
rect 5772 5372 5828 5428
rect 5828 5372 5832 5428
rect 5768 5368 5832 5372
rect 5928 5748 5992 5752
rect 5928 5692 5932 5748
rect 5932 5692 5988 5748
rect 5988 5692 5992 5748
rect 5928 5688 5992 5692
rect 5928 5528 5992 5592
rect 5928 5428 5992 5432
rect 5928 5372 5932 5428
rect 5932 5372 5988 5428
rect 5988 5372 5992 5428
rect 5928 5368 5992 5372
rect 6088 5748 6152 5752
rect 6088 5692 6092 5748
rect 6092 5692 6148 5748
rect 6148 5692 6152 5748
rect 6088 5688 6152 5692
rect 6088 5528 6152 5592
rect 6088 5428 6152 5432
rect 6088 5372 6092 5428
rect 6092 5372 6148 5428
rect 6148 5372 6152 5428
rect 6088 5368 6152 5372
rect 6248 5748 6312 5752
rect 6248 5692 6252 5748
rect 6252 5692 6308 5748
rect 6308 5692 6312 5748
rect 6248 5688 6312 5692
rect 6248 5528 6312 5592
rect 6248 5428 6312 5432
rect 6248 5372 6252 5428
rect 6252 5372 6308 5428
rect 6308 5372 6312 5428
rect 6248 5368 6312 5372
rect 6408 5748 6472 5752
rect 6408 5692 6412 5748
rect 6412 5692 6468 5748
rect 6468 5692 6472 5748
rect 6408 5688 6472 5692
rect 6408 5528 6472 5592
rect 6408 5428 6472 5432
rect 6408 5372 6412 5428
rect 6412 5372 6468 5428
rect 6468 5372 6472 5428
rect 6408 5368 6472 5372
rect 6568 5748 6632 5752
rect 6568 5692 6572 5748
rect 6572 5692 6628 5748
rect 6628 5692 6632 5748
rect 6568 5688 6632 5692
rect 6568 5528 6632 5592
rect 6568 5428 6632 5432
rect 6568 5372 6572 5428
rect 6572 5372 6628 5428
rect 6628 5372 6632 5428
rect 6568 5368 6632 5372
rect 6728 5748 6792 5752
rect 6728 5692 6732 5748
rect 6732 5692 6788 5748
rect 6788 5692 6792 5748
rect 6728 5688 6792 5692
rect 6728 5528 6792 5592
rect 6728 5428 6792 5432
rect 6728 5372 6732 5428
rect 6732 5372 6788 5428
rect 6788 5372 6792 5428
rect 6728 5368 6792 5372
rect 6888 5748 6952 5752
rect 6888 5692 6892 5748
rect 6892 5692 6948 5748
rect 6948 5692 6952 5748
rect 6888 5688 6952 5692
rect 6888 5528 6952 5592
rect 6888 5428 6952 5432
rect 6888 5372 6892 5428
rect 6892 5372 6948 5428
rect 6948 5372 6952 5428
rect 6888 5368 6952 5372
rect 7208 5748 7272 5752
rect 7208 5692 7212 5748
rect 7212 5692 7268 5748
rect 7268 5692 7272 5748
rect 7208 5688 7272 5692
rect 7208 5528 7272 5592
rect 7208 5428 7272 5432
rect 7208 5372 7212 5428
rect 7212 5372 7268 5428
rect 7268 5372 7272 5428
rect 7208 5368 7272 5372
rect 7368 5748 7432 5752
rect 7368 5692 7372 5748
rect 7372 5692 7428 5748
rect 7428 5692 7432 5748
rect 7368 5688 7432 5692
rect 7368 5528 7432 5592
rect 7368 5428 7432 5432
rect 7368 5372 7372 5428
rect 7372 5372 7428 5428
rect 7428 5372 7432 5428
rect 7368 5368 7432 5372
rect 7528 5748 7592 5752
rect 7528 5692 7532 5748
rect 7532 5692 7588 5748
rect 7588 5692 7592 5748
rect 7528 5688 7592 5692
rect 7528 5528 7592 5592
rect 7528 5428 7592 5432
rect 7528 5372 7532 5428
rect 7532 5372 7588 5428
rect 7588 5372 7592 5428
rect 7528 5368 7592 5372
rect 7688 5748 7752 5752
rect 7688 5692 7692 5748
rect 7692 5692 7748 5748
rect 7748 5692 7752 5748
rect 7688 5688 7752 5692
rect 7688 5528 7752 5592
rect 7688 5428 7752 5432
rect 7688 5372 7692 5428
rect 7692 5372 7748 5428
rect 7748 5372 7752 5428
rect 7688 5368 7752 5372
rect 7848 5748 7912 5752
rect 7848 5692 7852 5748
rect 7852 5692 7908 5748
rect 7908 5692 7912 5748
rect 7848 5688 7912 5692
rect 7848 5528 7912 5592
rect 7848 5428 7912 5432
rect 7848 5372 7852 5428
rect 7852 5372 7908 5428
rect 7908 5372 7912 5428
rect 7848 5368 7912 5372
rect 8168 5748 8232 5752
rect 8168 5692 8172 5748
rect 8172 5692 8228 5748
rect 8228 5692 8232 5748
rect 8168 5688 8232 5692
rect 8168 5528 8232 5592
rect 8168 5428 8232 5432
rect 8168 5372 8172 5428
rect 8172 5372 8228 5428
rect 8228 5372 8232 5428
rect 8168 5368 8232 5372
rect 328 4748 392 4752
rect 328 4692 332 4748
rect 332 4692 388 4748
rect 388 4692 392 4748
rect 328 4688 392 4692
rect 328 4668 392 4672
rect 328 4612 332 4668
rect 332 4612 388 4668
rect 388 4612 392 4668
rect 328 4608 392 4612
rect 328 4588 392 4592
rect 328 4532 332 4588
rect 332 4532 388 4588
rect 388 4532 392 4588
rect 328 4528 392 4532
rect 328 4508 392 4512
rect 328 4452 332 4508
rect 332 4452 388 4508
rect 388 4452 392 4508
rect 328 4448 392 4452
rect 8008 3628 8072 3632
rect 8008 3572 8012 3628
rect 8012 3572 8068 3628
rect 8068 3572 8072 3628
rect 8008 3568 8072 3572
rect 8008 3548 8072 3552
rect 8008 3492 8012 3548
rect 8012 3492 8068 3548
rect 8068 3492 8072 3548
rect 8008 3488 8072 3492
rect 8008 3468 8072 3472
rect 8008 3412 8012 3468
rect 8012 3412 8068 3468
rect 8068 3412 8072 3468
rect 8008 3408 8072 3412
rect 8008 3388 8072 3392
rect 8008 3332 8012 3388
rect 8012 3332 8068 3388
rect 8068 3332 8072 3388
rect 8008 3328 8072 3332
rect 8 2788 72 2792
rect 8 2732 12 2788
rect 12 2732 68 2788
rect 68 2732 72 2788
rect 8 2728 72 2732
rect 8 2468 72 2472
rect 8 2412 12 2468
rect 12 2412 68 2468
rect 68 2412 72 2468
rect 8 2408 72 2412
rect 168 2788 232 2792
rect 168 2732 172 2788
rect 172 2732 228 2788
rect 228 2732 232 2788
rect 168 2728 232 2732
rect 168 2468 232 2472
rect 168 2412 172 2468
rect 172 2412 228 2468
rect 228 2412 232 2468
rect 168 2408 232 2412
rect 328 2788 392 2792
rect 328 2732 332 2788
rect 332 2732 388 2788
rect 388 2732 392 2788
rect 328 2728 392 2732
rect 328 2468 392 2472
rect 328 2412 332 2468
rect 332 2412 388 2468
rect 388 2412 392 2468
rect 328 2408 392 2412
rect 488 2788 552 2792
rect 488 2732 492 2788
rect 492 2732 548 2788
rect 548 2732 552 2788
rect 488 2728 552 2732
rect 488 2468 552 2472
rect 488 2412 492 2468
rect 492 2412 548 2468
rect 548 2412 552 2468
rect 488 2408 552 2412
rect 648 2788 712 2792
rect 648 2732 652 2788
rect 652 2732 708 2788
rect 708 2732 712 2788
rect 648 2728 712 2732
rect 648 2468 712 2472
rect 648 2412 652 2468
rect 652 2412 708 2468
rect 708 2412 712 2468
rect 648 2408 712 2412
rect 808 2788 872 2792
rect 808 2732 812 2788
rect 812 2732 868 2788
rect 868 2732 872 2788
rect 808 2728 872 2732
rect 808 2468 872 2472
rect 808 2412 812 2468
rect 812 2412 868 2468
rect 868 2412 872 2468
rect 808 2408 872 2412
rect 968 2788 1032 2792
rect 968 2732 972 2788
rect 972 2732 1028 2788
rect 1028 2732 1032 2788
rect 968 2728 1032 2732
rect 968 2468 1032 2472
rect 968 2412 972 2468
rect 972 2412 1028 2468
rect 1028 2412 1032 2468
rect 968 2408 1032 2412
rect 1128 2788 1192 2792
rect 1128 2732 1132 2788
rect 1132 2732 1188 2788
rect 1188 2732 1192 2788
rect 1128 2728 1192 2732
rect 1128 2468 1192 2472
rect 1128 2412 1132 2468
rect 1132 2412 1188 2468
rect 1188 2412 1192 2468
rect 1128 2408 1192 2412
rect 1448 2788 1512 2792
rect 1448 2732 1452 2788
rect 1452 2732 1508 2788
rect 1508 2732 1512 2788
rect 1448 2728 1512 2732
rect 1448 2468 1512 2472
rect 1448 2412 1452 2468
rect 1452 2412 1508 2468
rect 1508 2412 1512 2468
rect 1448 2408 1512 2412
rect 1608 2788 1672 2792
rect 1608 2732 1612 2788
rect 1612 2732 1668 2788
rect 1668 2732 1672 2788
rect 1608 2728 1672 2732
rect 1608 2468 1672 2472
rect 1608 2412 1612 2468
rect 1612 2412 1668 2468
rect 1668 2412 1672 2468
rect 1608 2408 1672 2412
rect 1768 2788 1832 2792
rect 1768 2732 1772 2788
rect 1772 2732 1828 2788
rect 1828 2732 1832 2788
rect 1768 2728 1832 2732
rect 1768 2468 1832 2472
rect 1768 2412 1772 2468
rect 1772 2412 1828 2468
rect 1828 2412 1832 2468
rect 1768 2408 1832 2412
rect 1928 2788 1992 2792
rect 1928 2732 1932 2788
rect 1932 2732 1988 2788
rect 1988 2732 1992 2788
rect 1928 2728 1992 2732
rect 1928 2468 1992 2472
rect 1928 2412 1932 2468
rect 1932 2412 1988 2468
rect 1988 2412 1992 2468
rect 1928 2408 1992 2412
rect 2088 2788 2152 2792
rect 2088 2732 2092 2788
rect 2092 2732 2148 2788
rect 2148 2732 2152 2788
rect 2088 2728 2152 2732
rect 2088 2468 2152 2472
rect 2088 2412 2092 2468
rect 2092 2412 2148 2468
rect 2148 2412 2152 2468
rect 2088 2408 2152 2412
rect 2248 2788 2312 2792
rect 2248 2732 2252 2788
rect 2252 2732 2308 2788
rect 2308 2732 2312 2788
rect 2248 2728 2312 2732
rect 2248 2468 2312 2472
rect 2248 2412 2252 2468
rect 2252 2412 2308 2468
rect 2308 2412 2312 2468
rect 2248 2408 2312 2412
rect 2408 2788 2472 2792
rect 2408 2732 2412 2788
rect 2412 2732 2468 2788
rect 2468 2732 2472 2788
rect 2408 2728 2472 2732
rect 2408 2468 2472 2472
rect 2408 2412 2412 2468
rect 2412 2412 2468 2468
rect 2468 2412 2472 2468
rect 2408 2408 2472 2412
rect 2568 2788 2632 2792
rect 2568 2732 2572 2788
rect 2572 2732 2628 2788
rect 2628 2732 2632 2788
rect 2568 2728 2632 2732
rect 2568 2468 2632 2472
rect 2568 2412 2572 2468
rect 2572 2412 2628 2468
rect 2628 2412 2632 2468
rect 2568 2408 2632 2412
rect 2728 2788 2792 2792
rect 2728 2732 2732 2788
rect 2732 2732 2788 2788
rect 2788 2732 2792 2788
rect 2728 2728 2792 2732
rect 2728 2468 2792 2472
rect 2728 2412 2732 2468
rect 2732 2412 2788 2468
rect 2788 2412 2792 2468
rect 2728 2408 2792 2412
rect 2888 2788 2952 2792
rect 2888 2732 2892 2788
rect 2892 2732 2948 2788
rect 2948 2732 2952 2788
rect 2888 2728 2952 2732
rect 2888 2468 2952 2472
rect 2888 2412 2892 2468
rect 2892 2412 2948 2468
rect 2948 2412 2952 2468
rect 2888 2408 2952 2412
rect 3048 2788 3112 2792
rect 3048 2732 3052 2788
rect 3052 2732 3108 2788
rect 3108 2732 3112 2788
rect 3048 2728 3112 2732
rect 3048 2468 3112 2472
rect 3048 2412 3052 2468
rect 3052 2412 3108 2468
rect 3108 2412 3112 2468
rect 3048 2408 3112 2412
rect 3368 2788 3432 2792
rect 3368 2732 3372 2788
rect 3372 2732 3428 2788
rect 3428 2732 3432 2788
rect 3368 2728 3432 2732
rect 3368 2468 3432 2472
rect 3368 2412 3372 2468
rect 3372 2412 3428 2468
rect 3428 2412 3432 2468
rect 3368 2408 3432 2412
rect 3528 2788 3592 2792
rect 3528 2732 3532 2788
rect 3532 2732 3588 2788
rect 3588 2732 3592 2788
rect 3528 2728 3592 2732
rect 3528 2468 3592 2472
rect 3528 2412 3532 2468
rect 3532 2412 3588 2468
rect 3588 2412 3592 2468
rect 3528 2408 3592 2412
rect 3688 2788 3752 2792
rect 3688 2732 3692 2788
rect 3692 2732 3748 2788
rect 3748 2732 3752 2788
rect 3688 2728 3752 2732
rect 3688 2468 3752 2472
rect 3688 2412 3692 2468
rect 3692 2412 3748 2468
rect 3748 2412 3752 2468
rect 3688 2408 3752 2412
rect 3848 2788 3912 2792
rect 3848 2732 3852 2788
rect 3852 2732 3908 2788
rect 3908 2732 3912 2788
rect 3848 2728 3912 2732
rect 3848 2468 3912 2472
rect 3848 2412 3852 2468
rect 3852 2412 3908 2468
rect 3908 2412 3912 2468
rect 3848 2408 3912 2412
rect 4008 2788 4072 2792
rect 4008 2732 4012 2788
rect 4012 2732 4068 2788
rect 4068 2732 4072 2788
rect 4008 2728 4072 2732
rect 4008 2468 4072 2472
rect 4008 2412 4012 2468
rect 4012 2412 4068 2468
rect 4068 2412 4072 2468
rect 4008 2408 4072 2412
rect 4168 2788 4232 2792
rect 4168 2732 4172 2788
rect 4172 2732 4228 2788
rect 4228 2732 4232 2788
rect 4168 2728 4232 2732
rect 4168 2468 4232 2472
rect 4168 2412 4172 2468
rect 4172 2412 4228 2468
rect 4228 2412 4232 2468
rect 4168 2408 4232 2412
rect 4328 2788 4392 2792
rect 4328 2732 4332 2788
rect 4332 2732 4388 2788
rect 4388 2732 4392 2788
rect 4328 2728 4392 2732
rect 4328 2468 4392 2472
rect 4328 2412 4332 2468
rect 4332 2412 4388 2468
rect 4388 2412 4392 2468
rect 4328 2408 4392 2412
rect 4488 2788 4552 2792
rect 4488 2732 4492 2788
rect 4492 2732 4548 2788
rect 4548 2732 4552 2788
rect 4488 2728 4552 2732
rect 4488 2468 4552 2472
rect 4488 2412 4492 2468
rect 4492 2412 4548 2468
rect 4548 2412 4552 2468
rect 4488 2408 4552 2412
rect 4648 2788 4712 2792
rect 4648 2732 4652 2788
rect 4652 2732 4708 2788
rect 4708 2732 4712 2788
rect 4648 2728 4712 2732
rect 4648 2468 4712 2472
rect 4648 2412 4652 2468
rect 4652 2412 4708 2468
rect 4708 2412 4712 2468
rect 4648 2408 4712 2412
rect 4808 2788 4872 2792
rect 4808 2732 4812 2788
rect 4812 2732 4868 2788
rect 4868 2732 4872 2788
rect 4808 2728 4872 2732
rect 4808 2468 4872 2472
rect 4808 2412 4812 2468
rect 4812 2412 4868 2468
rect 4868 2412 4872 2468
rect 4808 2408 4872 2412
rect 4968 2788 5032 2792
rect 4968 2732 4972 2788
rect 4972 2732 5028 2788
rect 5028 2732 5032 2788
rect 4968 2728 5032 2732
rect 4968 2468 5032 2472
rect 4968 2412 4972 2468
rect 4972 2412 5028 2468
rect 5028 2412 5032 2468
rect 4968 2408 5032 2412
rect 5288 2788 5352 2792
rect 5288 2732 5292 2788
rect 5292 2732 5348 2788
rect 5348 2732 5352 2788
rect 5288 2728 5352 2732
rect 5288 2468 5352 2472
rect 5288 2412 5292 2468
rect 5292 2412 5348 2468
rect 5348 2412 5352 2468
rect 5288 2408 5352 2412
rect 5448 2788 5512 2792
rect 5448 2732 5452 2788
rect 5452 2732 5508 2788
rect 5508 2732 5512 2788
rect 5448 2728 5512 2732
rect 5448 2468 5512 2472
rect 5448 2412 5452 2468
rect 5452 2412 5508 2468
rect 5508 2412 5512 2468
rect 5448 2408 5512 2412
rect 5608 2788 5672 2792
rect 5608 2732 5612 2788
rect 5612 2732 5668 2788
rect 5668 2732 5672 2788
rect 5608 2728 5672 2732
rect 5608 2468 5672 2472
rect 5608 2412 5612 2468
rect 5612 2412 5668 2468
rect 5668 2412 5672 2468
rect 5608 2408 5672 2412
rect 5768 2788 5832 2792
rect 5768 2732 5772 2788
rect 5772 2732 5828 2788
rect 5828 2732 5832 2788
rect 5768 2728 5832 2732
rect 5768 2468 5832 2472
rect 5768 2412 5772 2468
rect 5772 2412 5828 2468
rect 5828 2412 5832 2468
rect 5768 2408 5832 2412
rect 5928 2788 5992 2792
rect 5928 2732 5932 2788
rect 5932 2732 5988 2788
rect 5988 2732 5992 2788
rect 5928 2728 5992 2732
rect 5928 2468 5992 2472
rect 5928 2412 5932 2468
rect 5932 2412 5988 2468
rect 5988 2412 5992 2468
rect 5928 2408 5992 2412
rect 6088 2788 6152 2792
rect 6088 2732 6092 2788
rect 6092 2732 6148 2788
rect 6148 2732 6152 2788
rect 6088 2728 6152 2732
rect 6088 2468 6152 2472
rect 6088 2412 6092 2468
rect 6092 2412 6148 2468
rect 6148 2412 6152 2468
rect 6088 2408 6152 2412
rect 6248 2788 6312 2792
rect 6248 2732 6252 2788
rect 6252 2732 6308 2788
rect 6308 2732 6312 2788
rect 6248 2728 6312 2732
rect 6248 2468 6312 2472
rect 6248 2412 6252 2468
rect 6252 2412 6308 2468
rect 6308 2412 6312 2468
rect 6248 2408 6312 2412
rect 6408 2788 6472 2792
rect 6408 2732 6412 2788
rect 6412 2732 6468 2788
rect 6468 2732 6472 2788
rect 6408 2728 6472 2732
rect 6408 2468 6472 2472
rect 6408 2412 6412 2468
rect 6412 2412 6468 2468
rect 6468 2412 6472 2468
rect 6408 2408 6472 2412
rect 6568 2788 6632 2792
rect 6568 2732 6572 2788
rect 6572 2732 6628 2788
rect 6628 2732 6632 2788
rect 6568 2728 6632 2732
rect 6568 2468 6632 2472
rect 6568 2412 6572 2468
rect 6572 2412 6628 2468
rect 6628 2412 6632 2468
rect 6568 2408 6632 2412
rect 6728 2788 6792 2792
rect 6728 2732 6732 2788
rect 6732 2732 6788 2788
rect 6788 2732 6792 2788
rect 6728 2728 6792 2732
rect 6728 2468 6792 2472
rect 6728 2412 6732 2468
rect 6732 2412 6788 2468
rect 6788 2412 6792 2468
rect 6728 2408 6792 2412
rect 6888 2788 6952 2792
rect 6888 2732 6892 2788
rect 6892 2732 6948 2788
rect 6948 2732 6952 2788
rect 6888 2728 6952 2732
rect 6888 2468 6952 2472
rect 6888 2412 6892 2468
rect 6892 2412 6948 2468
rect 6948 2412 6952 2468
rect 6888 2408 6952 2412
rect 7208 2788 7272 2792
rect 7208 2732 7212 2788
rect 7212 2732 7268 2788
rect 7268 2732 7272 2788
rect 7208 2728 7272 2732
rect 7208 2468 7272 2472
rect 7208 2412 7212 2468
rect 7212 2412 7268 2468
rect 7268 2412 7272 2468
rect 7208 2408 7272 2412
rect 7368 2788 7432 2792
rect 7368 2732 7372 2788
rect 7372 2732 7428 2788
rect 7428 2732 7432 2788
rect 7368 2728 7432 2732
rect 7368 2468 7432 2472
rect 7368 2412 7372 2468
rect 7372 2412 7428 2468
rect 7428 2412 7432 2468
rect 7368 2408 7432 2412
rect 7528 2788 7592 2792
rect 7528 2732 7532 2788
rect 7532 2732 7588 2788
rect 7588 2732 7592 2788
rect 7528 2728 7592 2732
rect 7528 2468 7592 2472
rect 7528 2412 7532 2468
rect 7532 2412 7588 2468
rect 7588 2412 7592 2468
rect 7528 2408 7592 2412
rect 7688 2788 7752 2792
rect 7688 2732 7692 2788
rect 7692 2732 7748 2788
rect 7748 2732 7752 2788
rect 7688 2728 7752 2732
rect 7688 2468 7752 2472
rect 7688 2412 7692 2468
rect 7692 2412 7748 2468
rect 7748 2412 7752 2468
rect 7688 2408 7752 2412
rect 7848 2788 7912 2792
rect 7848 2732 7852 2788
rect 7852 2732 7908 2788
rect 7908 2732 7912 2788
rect 7848 2728 7912 2732
rect 7848 2468 7912 2472
rect 7848 2412 7852 2468
rect 7852 2412 7908 2468
rect 7908 2412 7912 2468
rect 7848 2408 7912 2412
rect 8008 2788 8072 2792
rect 8008 2732 8012 2788
rect 8012 2732 8068 2788
rect 8068 2732 8072 2788
rect 8008 2728 8072 2732
rect 8008 2468 8072 2472
rect 8008 2412 8012 2468
rect 8012 2412 8068 2468
rect 8068 2412 8072 2468
rect 8008 2408 8072 2412
rect 8168 2788 8232 2792
rect 8168 2732 8172 2788
rect 8172 2732 8228 2788
rect 8228 2732 8232 2788
rect 8168 2728 8232 2732
rect 8168 2468 8232 2472
rect 8168 2412 8172 2468
rect 8172 2412 8228 2468
rect 8228 2412 8232 2468
rect 8168 2408 8232 2412
rect 8328 2788 8392 2792
rect 8328 2732 8332 2788
rect 8332 2732 8388 2788
rect 8388 2732 8392 2788
rect 8328 2728 8392 2732
rect 8328 2468 8392 2472
rect 8328 2412 8332 2468
rect 8332 2412 8388 2468
rect 8388 2412 8392 2468
rect 8328 2408 8392 2412
rect 168 1048 232 1112
rect 168 948 232 952
rect 168 892 172 948
rect 172 892 228 948
rect 228 892 232 948
rect 168 888 232 892
rect 168 728 232 792
rect 328 1048 392 1112
rect 328 948 392 952
rect 328 892 332 948
rect 332 892 388 948
rect 388 892 392 948
rect 328 888 392 892
rect 328 728 392 792
rect 488 1048 552 1112
rect 488 948 552 952
rect 488 892 492 948
rect 492 892 548 948
rect 548 892 552 948
rect 488 888 552 892
rect 488 728 552 792
rect 648 1048 712 1112
rect 648 948 712 952
rect 648 892 652 948
rect 652 892 708 948
rect 708 892 712 948
rect 648 888 712 892
rect 648 728 712 792
rect 808 1048 872 1112
rect 808 948 872 952
rect 808 892 812 948
rect 812 892 868 948
rect 868 892 872 948
rect 808 888 872 892
rect 808 728 872 792
rect 968 1048 1032 1112
rect 968 948 1032 952
rect 968 892 972 948
rect 972 892 1028 948
rect 1028 892 1032 948
rect 968 888 1032 892
rect 968 728 1032 792
rect 1128 1048 1192 1112
rect 1128 948 1192 952
rect 1128 892 1132 948
rect 1132 892 1188 948
rect 1188 892 1192 948
rect 1128 888 1192 892
rect 1128 728 1192 792
rect 1448 1048 1512 1112
rect 1448 948 1512 952
rect 1448 892 1452 948
rect 1452 892 1508 948
rect 1508 892 1512 948
rect 1448 888 1512 892
rect 1448 728 1512 792
rect 1608 1048 1672 1112
rect 1608 948 1672 952
rect 1608 892 1612 948
rect 1612 892 1668 948
rect 1668 892 1672 948
rect 1608 888 1672 892
rect 1608 728 1672 792
rect 1768 1048 1832 1112
rect 1768 948 1832 952
rect 1768 892 1772 948
rect 1772 892 1828 948
rect 1828 892 1832 948
rect 1768 888 1832 892
rect 1768 728 1832 792
rect 1928 1048 1992 1112
rect 1928 948 1992 952
rect 1928 892 1932 948
rect 1932 892 1988 948
rect 1988 892 1992 948
rect 1928 888 1992 892
rect 1928 728 1992 792
rect 2088 1048 2152 1112
rect 2088 948 2152 952
rect 2088 892 2092 948
rect 2092 892 2148 948
rect 2148 892 2152 948
rect 2088 888 2152 892
rect 2088 728 2152 792
rect 2248 1048 2312 1112
rect 2248 948 2312 952
rect 2248 892 2252 948
rect 2252 892 2308 948
rect 2308 892 2312 948
rect 2248 888 2312 892
rect 2248 728 2312 792
rect 2408 1048 2472 1112
rect 2408 948 2472 952
rect 2408 892 2412 948
rect 2412 892 2468 948
rect 2468 892 2472 948
rect 2408 888 2472 892
rect 2408 728 2472 792
rect 2568 1048 2632 1112
rect 2568 948 2632 952
rect 2568 892 2572 948
rect 2572 892 2628 948
rect 2628 892 2632 948
rect 2568 888 2632 892
rect 2568 728 2632 792
rect 2728 1048 2792 1112
rect 2728 948 2792 952
rect 2728 892 2732 948
rect 2732 892 2788 948
rect 2788 892 2792 948
rect 2728 888 2792 892
rect 2728 728 2792 792
rect 2888 1048 2952 1112
rect 2888 948 2952 952
rect 2888 892 2892 948
rect 2892 892 2948 948
rect 2948 892 2952 948
rect 2888 888 2952 892
rect 2888 728 2952 792
rect 3048 1048 3112 1112
rect 3048 948 3112 952
rect 3048 892 3052 948
rect 3052 892 3108 948
rect 3108 892 3112 948
rect 3048 888 3112 892
rect 3048 728 3112 792
rect 3368 1048 3432 1112
rect 3368 948 3432 952
rect 3368 892 3372 948
rect 3372 892 3428 948
rect 3428 892 3432 948
rect 3368 888 3432 892
rect 3368 728 3432 792
rect 3528 1048 3592 1112
rect 3528 948 3592 952
rect 3528 892 3532 948
rect 3532 892 3588 948
rect 3588 892 3592 948
rect 3528 888 3592 892
rect 3528 728 3592 792
rect 3688 1048 3752 1112
rect 3688 948 3752 952
rect 3688 892 3692 948
rect 3692 892 3748 948
rect 3748 892 3752 948
rect 3688 888 3752 892
rect 3688 728 3752 792
rect 3848 1048 3912 1112
rect 3848 948 3912 952
rect 3848 892 3852 948
rect 3852 892 3908 948
rect 3908 892 3912 948
rect 3848 888 3912 892
rect 3848 728 3912 792
rect 4008 1048 4072 1112
rect 4008 948 4072 952
rect 4008 892 4012 948
rect 4012 892 4068 948
rect 4068 892 4072 948
rect 4008 888 4072 892
rect 4008 728 4072 792
rect 4168 1048 4232 1112
rect 4168 948 4232 952
rect 4168 892 4172 948
rect 4172 892 4228 948
rect 4228 892 4232 948
rect 4168 888 4232 892
rect 4168 728 4232 792
rect 4328 1048 4392 1112
rect 4328 948 4392 952
rect 4328 892 4332 948
rect 4332 892 4388 948
rect 4388 892 4392 948
rect 4328 888 4392 892
rect 4328 728 4392 792
rect 4488 1048 4552 1112
rect 4488 948 4552 952
rect 4488 892 4492 948
rect 4492 892 4548 948
rect 4548 892 4552 948
rect 4488 888 4552 892
rect 4488 728 4552 792
rect 4648 1048 4712 1112
rect 4648 948 4712 952
rect 4648 892 4652 948
rect 4652 892 4708 948
rect 4708 892 4712 948
rect 4648 888 4712 892
rect 4648 728 4712 792
rect 4808 1048 4872 1112
rect 4808 948 4872 952
rect 4808 892 4812 948
rect 4812 892 4868 948
rect 4868 892 4872 948
rect 4808 888 4872 892
rect 4808 728 4872 792
rect 4968 1048 5032 1112
rect 4968 948 5032 952
rect 4968 892 4972 948
rect 4972 892 5028 948
rect 5028 892 5032 948
rect 4968 888 5032 892
rect 4968 728 5032 792
rect 5288 1048 5352 1112
rect 5288 948 5352 952
rect 5288 892 5292 948
rect 5292 892 5348 948
rect 5348 892 5352 948
rect 5288 888 5352 892
rect 5288 728 5352 792
rect 5448 1048 5512 1112
rect 5448 948 5512 952
rect 5448 892 5452 948
rect 5452 892 5508 948
rect 5508 892 5512 948
rect 5448 888 5512 892
rect 5448 728 5512 792
rect 5608 1048 5672 1112
rect 5608 948 5672 952
rect 5608 892 5612 948
rect 5612 892 5668 948
rect 5668 892 5672 948
rect 5608 888 5672 892
rect 5608 728 5672 792
rect 5768 1048 5832 1112
rect 5768 948 5832 952
rect 5768 892 5772 948
rect 5772 892 5828 948
rect 5828 892 5832 948
rect 5768 888 5832 892
rect 5768 728 5832 792
rect 5928 1048 5992 1112
rect 5928 948 5992 952
rect 5928 892 5932 948
rect 5932 892 5988 948
rect 5988 892 5992 948
rect 5928 888 5992 892
rect 5928 728 5992 792
rect 6088 1048 6152 1112
rect 6088 948 6152 952
rect 6088 892 6092 948
rect 6092 892 6148 948
rect 6148 892 6152 948
rect 6088 888 6152 892
rect 6088 728 6152 792
rect 6248 1048 6312 1112
rect 6248 948 6312 952
rect 6248 892 6252 948
rect 6252 892 6308 948
rect 6308 892 6312 948
rect 6248 888 6312 892
rect 6248 728 6312 792
rect 6408 1048 6472 1112
rect 6408 948 6472 952
rect 6408 892 6412 948
rect 6412 892 6468 948
rect 6468 892 6472 948
rect 6408 888 6472 892
rect 6408 728 6472 792
rect 6568 1048 6632 1112
rect 6568 948 6632 952
rect 6568 892 6572 948
rect 6572 892 6628 948
rect 6628 892 6632 948
rect 6568 888 6632 892
rect 6568 728 6632 792
rect 6728 1048 6792 1112
rect 6728 948 6792 952
rect 6728 892 6732 948
rect 6732 892 6788 948
rect 6788 892 6792 948
rect 6728 888 6792 892
rect 6728 728 6792 792
rect 6888 1048 6952 1112
rect 6888 948 6952 952
rect 6888 892 6892 948
rect 6892 892 6948 948
rect 6948 892 6952 948
rect 6888 888 6952 892
rect 6888 728 6952 792
rect 7208 1048 7272 1112
rect 7208 948 7272 952
rect 7208 892 7212 948
rect 7212 892 7268 948
rect 7268 892 7272 948
rect 7208 888 7272 892
rect 7208 728 7272 792
rect 7368 1048 7432 1112
rect 7368 948 7432 952
rect 7368 892 7372 948
rect 7372 892 7428 948
rect 7428 892 7432 948
rect 7368 888 7432 892
rect 7368 728 7432 792
rect 7528 1048 7592 1112
rect 7528 948 7592 952
rect 7528 892 7532 948
rect 7532 892 7588 948
rect 7588 892 7592 948
rect 7528 888 7592 892
rect 7528 728 7592 792
rect 7688 1048 7752 1112
rect 7688 948 7752 952
rect 7688 892 7692 948
rect 7692 892 7748 948
rect 7748 892 7752 948
rect 7688 888 7752 892
rect 7688 728 7752 792
rect 7848 1048 7912 1112
rect 7848 948 7912 952
rect 7848 892 7852 948
rect 7852 892 7908 948
rect 7908 892 7912 948
rect 7848 888 7912 892
rect 7848 728 7912 792
rect 8168 1048 8232 1112
rect 8168 948 8232 952
rect 8168 892 8172 948
rect 8172 892 8228 948
rect 8228 892 8232 948
rect 8168 888 8232 892
rect 8168 728 8232 792
rect 328 328 392 332
rect 328 272 332 328
rect 332 272 388 328
rect 388 272 392 328
rect 328 268 392 272
rect 328 248 392 252
rect 328 192 332 248
rect 332 192 388 248
rect 388 192 392 248
rect 328 188 392 192
rect 168 -92 232 -88
rect 168 -148 172 -92
rect 172 -148 228 -92
rect 228 -148 232 -92
rect 168 -152 232 -148
rect 168 -312 232 -248
rect 168 -412 232 -408
rect 168 -468 172 -412
rect 172 -468 228 -412
rect 228 -468 232 -412
rect 168 -472 232 -468
rect 328 -92 392 -88
rect 328 -148 332 -92
rect 332 -148 388 -92
rect 388 -148 392 -92
rect 328 -152 392 -148
rect 328 -312 392 -248
rect 328 -412 392 -408
rect 328 -468 332 -412
rect 332 -468 388 -412
rect 388 -468 392 -412
rect 328 -472 392 -468
rect 488 -92 552 -88
rect 488 -148 492 -92
rect 492 -148 548 -92
rect 548 -148 552 -92
rect 488 -152 552 -148
rect 488 -312 552 -248
rect 488 -412 552 -408
rect 488 -468 492 -412
rect 492 -468 548 -412
rect 548 -468 552 -412
rect 488 -472 552 -468
rect 648 -92 712 -88
rect 648 -148 652 -92
rect 652 -148 708 -92
rect 708 -148 712 -92
rect 648 -152 712 -148
rect 648 -312 712 -248
rect 648 -412 712 -408
rect 648 -468 652 -412
rect 652 -468 708 -412
rect 708 -468 712 -412
rect 648 -472 712 -468
rect 808 -92 872 -88
rect 808 -148 812 -92
rect 812 -148 868 -92
rect 868 -148 872 -92
rect 808 -152 872 -148
rect 808 -312 872 -248
rect 808 -412 872 -408
rect 808 -468 812 -412
rect 812 -468 868 -412
rect 868 -468 872 -412
rect 808 -472 872 -468
rect 968 -92 1032 -88
rect 968 -148 972 -92
rect 972 -148 1028 -92
rect 1028 -148 1032 -92
rect 968 -152 1032 -148
rect 968 -312 1032 -248
rect 968 -412 1032 -408
rect 968 -468 972 -412
rect 972 -468 1028 -412
rect 1028 -468 1032 -412
rect 968 -472 1032 -468
rect 1128 -92 1192 -88
rect 1128 -148 1132 -92
rect 1132 -148 1188 -92
rect 1188 -148 1192 -92
rect 1128 -152 1192 -148
rect 1128 -312 1192 -248
rect 1128 -412 1192 -408
rect 1128 -468 1132 -412
rect 1132 -468 1188 -412
rect 1188 -468 1192 -412
rect 1128 -472 1192 -468
rect 1448 -92 1512 -88
rect 1448 -148 1452 -92
rect 1452 -148 1508 -92
rect 1508 -148 1512 -92
rect 1448 -152 1512 -148
rect 1448 -312 1512 -248
rect 1448 -412 1512 -408
rect 1448 -468 1452 -412
rect 1452 -468 1508 -412
rect 1508 -468 1512 -412
rect 1448 -472 1512 -468
rect 1608 -92 1672 -88
rect 1608 -148 1612 -92
rect 1612 -148 1668 -92
rect 1668 -148 1672 -92
rect 1608 -152 1672 -148
rect 1608 -312 1672 -248
rect 1608 -412 1672 -408
rect 1608 -468 1612 -412
rect 1612 -468 1668 -412
rect 1668 -468 1672 -412
rect 1608 -472 1672 -468
rect 1768 -92 1832 -88
rect 1768 -148 1772 -92
rect 1772 -148 1828 -92
rect 1828 -148 1832 -92
rect 1768 -152 1832 -148
rect 1768 -312 1832 -248
rect 1768 -412 1832 -408
rect 1768 -468 1772 -412
rect 1772 -468 1828 -412
rect 1828 -468 1832 -412
rect 1768 -472 1832 -468
rect 1928 -92 1992 -88
rect 1928 -148 1932 -92
rect 1932 -148 1988 -92
rect 1988 -148 1992 -92
rect 1928 -152 1992 -148
rect 1928 -312 1992 -248
rect 1928 -412 1992 -408
rect 1928 -468 1932 -412
rect 1932 -468 1988 -412
rect 1988 -468 1992 -412
rect 1928 -472 1992 -468
rect 2088 -92 2152 -88
rect 2088 -148 2092 -92
rect 2092 -148 2148 -92
rect 2148 -148 2152 -92
rect 2088 -152 2152 -148
rect 2088 -312 2152 -248
rect 2088 -412 2152 -408
rect 2088 -468 2092 -412
rect 2092 -468 2148 -412
rect 2148 -468 2152 -412
rect 2088 -472 2152 -468
rect 2248 -92 2312 -88
rect 2248 -148 2252 -92
rect 2252 -148 2308 -92
rect 2308 -148 2312 -92
rect 2248 -152 2312 -148
rect 2248 -312 2312 -248
rect 2248 -412 2312 -408
rect 2248 -468 2252 -412
rect 2252 -468 2308 -412
rect 2308 -468 2312 -412
rect 2248 -472 2312 -468
rect 2408 -92 2472 -88
rect 2408 -148 2412 -92
rect 2412 -148 2468 -92
rect 2468 -148 2472 -92
rect 2408 -152 2472 -148
rect 2408 -312 2472 -248
rect 2408 -412 2472 -408
rect 2408 -468 2412 -412
rect 2412 -468 2468 -412
rect 2468 -468 2472 -412
rect 2408 -472 2472 -468
rect 2568 -92 2632 -88
rect 2568 -148 2572 -92
rect 2572 -148 2628 -92
rect 2628 -148 2632 -92
rect 2568 -152 2632 -148
rect 2568 -312 2632 -248
rect 2568 -412 2632 -408
rect 2568 -468 2572 -412
rect 2572 -468 2628 -412
rect 2628 -468 2632 -412
rect 2568 -472 2632 -468
rect 2728 -92 2792 -88
rect 2728 -148 2732 -92
rect 2732 -148 2788 -92
rect 2788 -148 2792 -92
rect 2728 -152 2792 -148
rect 2728 -312 2792 -248
rect 2728 -412 2792 -408
rect 2728 -468 2732 -412
rect 2732 -468 2788 -412
rect 2788 -468 2792 -412
rect 2728 -472 2792 -468
rect 2888 -92 2952 -88
rect 2888 -148 2892 -92
rect 2892 -148 2948 -92
rect 2948 -148 2952 -92
rect 2888 -152 2952 -148
rect 2888 -312 2952 -248
rect 2888 -412 2952 -408
rect 2888 -468 2892 -412
rect 2892 -468 2948 -412
rect 2948 -468 2952 -412
rect 2888 -472 2952 -468
rect 3048 -92 3112 -88
rect 3048 -148 3052 -92
rect 3052 -148 3108 -92
rect 3108 -148 3112 -92
rect 3048 -152 3112 -148
rect 3048 -312 3112 -248
rect 3048 -412 3112 -408
rect 3048 -468 3052 -412
rect 3052 -468 3108 -412
rect 3108 -468 3112 -412
rect 3048 -472 3112 -468
rect 3368 -92 3432 -88
rect 3368 -148 3372 -92
rect 3372 -148 3428 -92
rect 3428 -148 3432 -92
rect 3368 -152 3432 -148
rect 3368 -312 3432 -248
rect 3368 -412 3432 -408
rect 3368 -468 3372 -412
rect 3372 -468 3428 -412
rect 3428 -468 3432 -412
rect 3368 -472 3432 -468
rect 3528 -92 3592 -88
rect 3528 -148 3532 -92
rect 3532 -148 3588 -92
rect 3588 -148 3592 -92
rect 3528 -152 3592 -148
rect 3528 -312 3592 -248
rect 3528 -412 3592 -408
rect 3528 -468 3532 -412
rect 3532 -468 3588 -412
rect 3588 -468 3592 -412
rect 3528 -472 3592 -468
rect 3688 -92 3752 -88
rect 3688 -148 3692 -92
rect 3692 -148 3748 -92
rect 3748 -148 3752 -92
rect 3688 -152 3752 -148
rect 3688 -312 3752 -248
rect 3688 -412 3752 -408
rect 3688 -468 3692 -412
rect 3692 -468 3748 -412
rect 3748 -468 3752 -412
rect 3688 -472 3752 -468
rect 3848 -92 3912 -88
rect 3848 -148 3852 -92
rect 3852 -148 3908 -92
rect 3908 -148 3912 -92
rect 3848 -152 3912 -148
rect 3848 -312 3912 -248
rect 3848 -412 3912 -408
rect 3848 -468 3852 -412
rect 3852 -468 3908 -412
rect 3908 -468 3912 -412
rect 3848 -472 3912 -468
rect 4008 -92 4072 -88
rect 4008 -148 4012 -92
rect 4012 -148 4068 -92
rect 4068 -148 4072 -92
rect 4008 -152 4072 -148
rect 4008 -312 4072 -248
rect 4008 -412 4072 -408
rect 4008 -468 4012 -412
rect 4012 -468 4068 -412
rect 4068 -468 4072 -412
rect 4008 -472 4072 -468
rect 4168 -92 4232 -88
rect 4168 -148 4172 -92
rect 4172 -148 4228 -92
rect 4228 -148 4232 -92
rect 4168 -152 4232 -148
rect 4168 -312 4232 -248
rect 4168 -412 4232 -408
rect 4168 -468 4172 -412
rect 4172 -468 4228 -412
rect 4228 -468 4232 -412
rect 4168 -472 4232 -468
rect 4328 -92 4392 -88
rect 4328 -148 4332 -92
rect 4332 -148 4388 -92
rect 4388 -148 4392 -92
rect 4328 -152 4392 -148
rect 4328 -312 4392 -248
rect 4328 -412 4392 -408
rect 4328 -468 4332 -412
rect 4332 -468 4388 -412
rect 4388 -468 4392 -412
rect 4328 -472 4392 -468
rect 4488 -92 4552 -88
rect 4488 -148 4492 -92
rect 4492 -148 4548 -92
rect 4548 -148 4552 -92
rect 4488 -152 4552 -148
rect 4488 -312 4552 -248
rect 4488 -412 4552 -408
rect 4488 -468 4492 -412
rect 4492 -468 4548 -412
rect 4548 -468 4552 -412
rect 4488 -472 4552 -468
rect 4648 -92 4712 -88
rect 4648 -148 4652 -92
rect 4652 -148 4708 -92
rect 4708 -148 4712 -92
rect 4648 -152 4712 -148
rect 4648 -312 4712 -248
rect 4648 -412 4712 -408
rect 4648 -468 4652 -412
rect 4652 -468 4708 -412
rect 4708 -468 4712 -412
rect 4648 -472 4712 -468
rect 4808 -92 4872 -88
rect 4808 -148 4812 -92
rect 4812 -148 4868 -92
rect 4868 -148 4872 -92
rect 4808 -152 4872 -148
rect 4808 -312 4872 -248
rect 4808 -412 4872 -408
rect 4808 -468 4812 -412
rect 4812 -468 4868 -412
rect 4868 -468 4872 -412
rect 4808 -472 4872 -468
rect 4968 -92 5032 -88
rect 4968 -148 4972 -92
rect 4972 -148 5028 -92
rect 5028 -148 5032 -92
rect 4968 -152 5032 -148
rect 4968 -312 5032 -248
rect 4968 -412 5032 -408
rect 4968 -468 4972 -412
rect 4972 -468 5028 -412
rect 5028 -468 5032 -412
rect 4968 -472 5032 -468
rect 5288 -92 5352 -88
rect 5288 -148 5292 -92
rect 5292 -148 5348 -92
rect 5348 -148 5352 -92
rect 5288 -152 5352 -148
rect 5288 -312 5352 -248
rect 5288 -412 5352 -408
rect 5288 -468 5292 -412
rect 5292 -468 5348 -412
rect 5348 -468 5352 -412
rect 5288 -472 5352 -468
rect 5448 -92 5512 -88
rect 5448 -148 5452 -92
rect 5452 -148 5508 -92
rect 5508 -148 5512 -92
rect 5448 -152 5512 -148
rect 5448 -312 5512 -248
rect 5448 -412 5512 -408
rect 5448 -468 5452 -412
rect 5452 -468 5508 -412
rect 5508 -468 5512 -412
rect 5448 -472 5512 -468
rect 5608 -92 5672 -88
rect 5608 -148 5612 -92
rect 5612 -148 5668 -92
rect 5668 -148 5672 -92
rect 5608 -152 5672 -148
rect 5608 -312 5672 -248
rect 5608 -412 5672 -408
rect 5608 -468 5612 -412
rect 5612 -468 5668 -412
rect 5668 -468 5672 -412
rect 5608 -472 5672 -468
rect 5768 -92 5832 -88
rect 5768 -148 5772 -92
rect 5772 -148 5828 -92
rect 5828 -148 5832 -92
rect 5768 -152 5832 -148
rect 5768 -312 5832 -248
rect 5768 -412 5832 -408
rect 5768 -468 5772 -412
rect 5772 -468 5828 -412
rect 5828 -468 5832 -412
rect 5768 -472 5832 -468
rect 5928 -92 5992 -88
rect 5928 -148 5932 -92
rect 5932 -148 5988 -92
rect 5988 -148 5992 -92
rect 5928 -152 5992 -148
rect 5928 -312 5992 -248
rect 5928 -412 5992 -408
rect 5928 -468 5932 -412
rect 5932 -468 5988 -412
rect 5988 -468 5992 -412
rect 5928 -472 5992 -468
rect 6088 -92 6152 -88
rect 6088 -148 6092 -92
rect 6092 -148 6148 -92
rect 6148 -148 6152 -92
rect 6088 -152 6152 -148
rect 6088 -312 6152 -248
rect 6088 -412 6152 -408
rect 6088 -468 6092 -412
rect 6092 -468 6148 -412
rect 6148 -468 6152 -412
rect 6088 -472 6152 -468
rect 6248 -92 6312 -88
rect 6248 -148 6252 -92
rect 6252 -148 6308 -92
rect 6308 -148 6312 -92
rect 6248 -152 6312 -148
rect 6248 -312 6312 -248
rect 6248 -412 6312 -408
rect 6248 -468 6252 -412
rect 6252 -468 6308 -412
rect 6308 -468 6312 -412
rect 6248 -472 6312 -468
rect 6408 -92 6472 -88
rect 6408 -148 6412 -92
rect 6412 -148 6468 -92
rect 6468 -148 6472 -92
rect 6408 -152 6472 -148
rect 6408 -312 6472 -248
rect 6408 -412 6472 -408
rect 6408 -468 6412 -412
rect 6412 -468 6468 -412
rect 6468 -468 6472 -412
rect 6408 -472 6472 -468
rect 6568 -92 6632 -88
rect 6568 -148 6572 -92
rect 6572 -148 6628 -92
rect 6628 -148 6632 -92
rect 6568 -152 6632 -148
rect 6568 -312 6632 -248
rect 6568 -412 6632 -408
rect 6568 -468 6572 -412
rect 6572 -468 6628 -412
rect 6628 -468 6632 -412
rect 6568 -472 6632 -468
rect 6728 -92 6792 -88
rect 6728 -148 6732 -92
rect 6732 -148 6788 -92
rect 6788 -148 6792 -92
rect 6728 -152 6792 -148
rect 6728 -312 6792 -248
rect 6728 -412 6792 -408
rect 6728 -468 6732 -412
rect 6732 -468 6788 -412
rect 6788 -468 6792 -412
rect 6728 -472 6792 -468
rect 6888 -92 6952 -88
rect 6888 -148 6892 -92
rect 6892 -148 6948 -92
rect 6948 -148 6952 -92
rect 6888 -152 6952 -148
rect 6888 -312 6952 -248
rect 6888 -412 6952 -408
rect 6888 -468 6892 -412
rect 6892 -468 6948 -412
rect 6948 -468 6952 -412
rect 6888 -472 6952 -468
rect 7208 -92 7272 -88
rect 7208 -148 7212 -92
rect 7212 -148 7268 -92
rect 7268 -148 7272 -92
rect 7208 -152 7272 -148
rect 7208 -312 7272 -248
rect 7208 -412 7272 -408
rect 7208 -468 7212 -412
rect 7212 -468 7268 -412
rect 7268 -468 7272 -412
rect 7208 -472 7272 -468
rect 7368 -92 7432 -88
rect 7368 -148 7372 -92
rect 7372 -148 7428 -92
rect 7428 -148 7432 -92
rect 7368 -152 7432 -148
rect 7368 -312 7432 -248
rect 7368 -412 7432 -408
rect 7368 -468 7372 -412
rect 7372 -468 7428 -412
rect 7428 -468 7432 -412
rect 7368 -472 7432 -468
rect 7528 -92 7592 -88
rect 7528 -148 7532 -92
rect 7532 -148 7588 -92
rect 7588 -148 7592 -92
rect 7528 -152 7592 -148
rect 7528 -312 7592 -248
rect 7528 -412 7592 -408
rect 7528 -468 7532 -412
rect 7532 -468 7588 -412
rect 7588 -468 7592 -412
rect 7528 -472 7592 -468
rect 7688 -92 7752 -88
rect 7688 -148 7692 -92
rect 7692 -148 7748 -92
rect 7748 -148 7752 -92
rect 7688 -152 7752 -148
rect 7688 -312 7752 -248
rect 7688 -412 7752 -408
rect 7688 -468 7692 -412
rect 7692 -468 7748 -412
rect 7748 -468 7752 -412
rect 7688 -472 7752 -468
rect 7848 -92 7912 -88
rect 7848 -148 7852 -92
rect 7852 -148 7908 -92
rect 7908 -148 7912 -92
rect 7848 -152 7912 -148
rect 7848 -312 7912 -248
rect 7848 -412 7912 -408
rect 7848 -468 7852 -412
rect 7852 -468 7908 -412
rect 7908 -468 7912 -412
rect 7848 -472 7912 -468
rect 8168 -92 8232 -88
rect 8168 -148 8172 -92
rect 8172 -148 8228 -92
rect 8228 -148 8232 -92
rect 8168 -152 8232 -148
rect 8168 -312 8232 -248
rect 8168 -412 8232 -408
rect 8168 -468 8172 -412
rect 8172 -468 8228 -412
rect 8228 -468 8232 -412
rect 8168 -472 8232 -468
rect 328 -712 392 -708
rect 328 -768 332 -712
rect 332 -768 388 -712
rect 388 -768 392 -712
rect 328 -772 392 -768
rect 328 -792 392 -788
rect 328 -848 332 -792
rect 332 -848 388 -792
rect 388 -848 392 -792
rect 328 -852 392 -848
<< metal4 >>
rect 0 9712 8400 9760
rect 0 9678 328 9712
rect 392 9678 8400 9712
rect 0 9442 242 9678
rect 478 9442 7922 9678
rect 8158 9442 8400 9678
rect 0 9408 328 9442
rect 392 9408 8400 9442
rect 0 9360 8400 9408
rect 0 8792 8400 8800
rect 0 8728 168 8792
rect 232 8728 328 8792
rect 392 8728 488 8792
rect 552 8728 648 8792
rect 712 8728 808 8792
rect 872 8728 968 8792
rect 1032 8728 1128 8792
rect 1192 8728 1448 8792
rect 1512 8728 1608 8792
rect 1672 8728 1768 8792
rect 1832 8728 1928 8792
rect 1992 8728 2088 8792
rect 2152 8728 2248 8792
rect 2312 8728 2408 8792
rect 2472 8728 2568 8792
rect 2632 8728 2728 8792
rect 2792 8728 2888 8792
rect 2952 8728 3048 8792
rect 3112 8728 3368 8792
rect 3432 8728 3528 8792
rect 3592 8728 3688 8792
rect 3752 8728 3848 8792
rect 3912 8728 4008 8792
rect 4072 8728 4168 8792
rect 4232 8728 4328 8792
rect 4392 8728 4488 8792
rect 4552 8728 4648 8792
rect 4712 8728 4808 8792
rect 4872 8728 4968 8792
rect 5032 8728 5288 8792
rect 5352 8728 5448 8792
rect 5512 8728 5608 8792
rect 5672 8728 5768 8792
rect 5832 8728 5928 8792
rect 5992 8728 6088 8792
rect 6152 8728 6248 8792
rect 6312 8728 6408 8792
rect 6472 8728 6568 8792
rect 6632 8728 6728 8792
rect 6792 8728 6888 8792
rect 6952 8728 7208 8792
rect 7272 8728 7368 8792
rect 7432 8728 7528 8792
rect 7592 8728 7688 8792
rect 7752 8728 7848 8792
rect 7912 8728 8008 8792
rect 8072 8728 8168 8792
rect 8232 8728 8400 8792
rect 0 8718 8400 8728
rect 0 8632 242 8718
rect 478 8632 7922 8718
rect 8158 8632 8400 8718
rect 0 8568 168 8632
rect 232 8568 242 8632
rect 478 8568 488 8632
rect 552 8568 648 8632
rect 712 8568 808 8632
rect 872 8568 968 8632
rect 1032 8568 1128 8632
rect 1192 8568 1448 8632
rect 1512 8568 1608 8632
rect 1672 8568 1768 8632
rect 1832 8568 1928 8632
rect 1992 8568 2088 8632
rect 2152 8568 2248 8632
rect 2312 8568 2408 8632
rect 2472 8568 2568 8632
rect 2632 8568 2728 8632
rect 2792 8568 2888 8632
rect 2952 8568 3048 8632
rect 3112 8568 3368 8632
rect 3432 8568 3528 8632
rect 3592 8568 3688 8632
rect 3752 8568 3848 8632
rect 3912 8568 4008 8632
rect 4072 8568 4168 8632
rect 4232 8568 4328 8632
rect 4392 8568 4488 8632
rect 4552 8568 4648 8632
rect 4712 8568 4808 8632
rect 4872 8568 4968 8632
rect 5032 8568 5288 8632
rect 5352 8568 5448 8632
rect 5512 8568 5608 8632
rect 5672 8568 5768 8632
rect 5832 8568 5928 8632
rect 5992 8568 6088 8632
rect 6152 8568 6248 8632
rect 6312 8568 6408 8632
rect 6472 8568 6568 8632
rect 6632 8568 6728 8632
rect 6792 8568 6888 8632
rect 6952 8568 7208 8632
rect 7272 8568 7368 8632
rect 7432 8568 7528 8632
rect 7592 8568 7688 8632
rect 7752 8568 7848 8632
rect 7912 8568 7922 8632
rect 8158 8568 8168 8632
rect 8232 8568 8400 8632
rect 0 8482 242 8568
rect 478 8482 7922 8568
rect 8158 8482 8400 8568
rect 0 8472 8400 8482
rect 0 8408 168 8472
rect 232 8408 328 8472
rect 392 8408 488 8472
rect 552 8408 648 8472
rect 712 8408 808 8472
rect 872 8408 968 8472
rect 1032 8408 1128 8472
rect 1192 8408 1448 8472
rect 1512 8408 1608 8472
rect 1672 8408 1768 8472
rect 1832 8408 1928 8472
rect 1992 8408 2088 8472
rect 2152 8408 2248 8472
rect 2312 8408 2408 8472
rect 2472 8408 2568 8472
rect 2632 8408 2728 8472
rect 2792 8408 2888 8472
rect 2952 8408 3048 8472
rect 3112 8408 3368 8472
rect 3432 8408 3528 8472
rect 3592 8408 3688 8472
rect 3752 8408 3848 8472
rect 3912 8408 4008 8472
rect 4072 8408 4168 8472
rect 4232 8408 4328 8472
rect 4392 8408 4488 8472
rect 4552 8408 4648 8472
rect 4712 8408 4808 8472
rect 4872 8408 4968 8472
rect 5032 8408 5288 8472
rect 5352 8408 5448 8472
rect 5512 8408 5608 8472
rect 5672 8408 5768 8472
rect 5832 8408 5928 8472
rect 5992 8408 6088 8472
rect 6152 8408 6248 8472
rect 6312 8408 6408 8472
rect 6472 8408 6568 8472
rect 6632 8408 6728 8472
rect 6792 8408 6888 8472
rect 6952 8408 7208 8472
rect 7272 8408 7368 8472
rect 7432 8408 7528 8472
rect 7592 8408 7688 8472
rect 7752 8408 7848 8472
rect 7912 8408 8008 8472
rect 8072 8408 8168 8472
rect 8232 8408 8400 8472
rect 0 8400 8400 8408
rect 0 8312 8400 8320
rect 0 8248 168 8312
rect 232 8248 328 8312
rect 392 8248 488 8312
rect 552 8248 648 8312
rect 712 8248 808 8312
rect 872 8248 968 8312
rect 1032 8248 1128 8312
rect 1192 8248 1448 8312
rect 1512 8248 1608 8312
rect 1672 8248 1768 8312
rect 1832 8248 1928 8312
rect 1992 8248 2088 8312
rect 2152 8248 2248 8312
rect 2312 8248 2408 8312
rect 2472 8248 2568 8312
rect 2632 8248 2728 8312
rect 2792 8248 2888 8312
rect 2952 8248 3048 8312
rect 3112 8248 3368 8312
rect 3432 8248 3528 8312
rect 3592 8248 3688 8312
rect 3752 8248 3848 8312
rect 3912 8248 4008 8312
rect 4072 8248 4168 8312
rect 4232 8248 4328 8312
rect 4392 8248 4488 8312
rect 4552 8248 4648 8312
rect 4712 8248 4808 8312
rect 4872 8248 4968 8312
rect 5032 8248 5288 8312
rect 5352 8248 5448 8312
rect 5512 8248 5608 8312
rect 5672 8248 5768 8312
rect 5832 8248 5928 8312
rect 5992 8248 6088 8312
rect 6152 8248 6248 8312
rect 6312 8248 6408 8312
rect 6472 8248 6568 8312
rect 6632 8248 6728 8312
rect 6792 8248 6888 8312
rect 6952 8248 7208 8312
rect 7272 8248 7368 8312
rect 7432 8248 7528 8312
rect 7592 8248 7688 8312
rect 7752 8248 7848 8312
rect 7912 8248 8008 8312
rect 8072 8248 8168 8312
rect 8232 8248 8400 8312
rect 0 8238 8400 8248
rect 0 8152 3122 8238
rect 0 8088 168 8152
rect 232 8088 328 8152
rect 392 8088 488 8152
rect 552 8088 648 8152
rect 712 8088 808 8152
rect 872 8088 968 8152
rect 1032 8088 1128 8152
rect 1192 8088 1448 8152
rect 1512 8088 1608 8152
rect 1672 8088 1768 8152
rect 1832 8088 1928 8152
rect 1992 8088 2088 8152
rect 2152 8088 2248 8152
rect 2312 8088 2408 8152
rect 2472 8088 2568 8152
rect 2632 8088 2728 8152
rect 2792 8088 2888 8152
rect 2952 8088 3048 8152
rect 3112 8088 3122 8152
rect 0 8002 3122 8088
rect 3358 8152 5042 8238
rect 3358 8088 3368 8152
rect 3432 8088 3528 8152
rect 3592 8088 3688 8152
rect 3752 8088 3848 8152
rect 3912 8088 4008 8152
rect 4072 8088 4168 8152
rect 4232 8088 4328 8152
rect 4392 8088 4488 8152
rect 4552 8088 4648 8152
rect 4712 8088 4808 8152
rect 4872 8088 4968 8152
rect 5032 8088 5042 8152
rect 3358 8002 5042 8088
rect 5278 8152 8400 8238
rect 5278 8088 5288 8152
rect 5352 8088 5448 8152
rect 5512 8088 5608 8152
rect 5672 8088 5768 8152
rect 5832 8088 5928 8152
rect 5992 8088 6088 8152
rect 6152 8088 6248 8152
rect 6312 8088 6408 8152
rect 6472 8088 6568 8152
rect 6632 8088 6728 8152
rect 6792 8088 6888 8152
rect 6952 8088 7208 8152
rect 7272 8088 7368 8152
rect 7432 8088 7528 8152
rect 7592 8088 7688 8152
rect 7752 8088 7848 8152
rect 7912 8088 8008 8152
rect 8072 8088 8168 8152
rect 8232 8088 8400 8152
rect 5278 8002 8400 8088
rect 0 7992 8400 8002
rect 0 7928 168 7992
rect 232 7928 328 7992
rect 392 7928 488 7992
rect 552 7928 648 7992
rect 712 7928 808 7992
rect 872 7928 968 7992
rect 1032 7928 1128 7992
rect 1192 7928 1448 7992
rect 1512 7928 1608 7992
rect 1672 7928 1768 7992
rect 1832 7928 1928 7992
rect 1992 7928 2088 7992
rect 2152 7928 2248 7992
rect 2312 7928 2408 7992
rect 2472 7928 2568 7992
rect 2632 7928 2728 7992
rect 2792 7928 2888 7992
rect 2952 7928 3048 7992
rect 3112 7928 3368 7992
rect 3432 7928 3528 7992
rect 3592 7928 3688 7992
rect 3752 7928 3848 7992
rect 3912 7928 4008 7992
rect 4072 7928 4168 7992
rect 4232 7928 4328 7992
rect 4392 7928 4488 7992
rect 4552 7928 4648 7992
rect 4712 7928 4808 7992
rect 4872 7928 4968 7992
rect 5032 7928 5288 7992
rect 5352 7928 5448 7992
rect 5512 7928 5608 7992
rect 5672 7928 5768 7992
rect 5832 7928 5928 7992
rect 5992 7928 6088 7992
rect 6152 7928 6248 7992
rect 6312 7928 6408 7992
rect 6472 7928 6568 7992
rect 6632 7928 6728 7992
rect 6792 7928 6888 7992
rect 6952 7928 7208 7992
rect 7272 7928 7368 7992
rect 7432 7928 7528 7992
rect 7592 7928 7688 7992
rect 7752 7928 7848 7992
rect 7912 7928 8008 7992
rect 8072 7928 8168 7992
rect 8232 7928 8400 7992
rect 0 7920 8400 7928
rect 0 7692 8400 7760
rect 0 7628 328 7692
rect 392 7678 8400 7692
rect 392 7628 3122 7678
rect 0 7612 3122 7628
rect 0 7548 328 7612
rect 392 7548 3122 7612
rect 0 7442 3122 7548
rect 3358 7442 5042 7678
rect 5278 7442 8400 7678
rect 0 7360 8400 7442
rect 0 7198 8400 7280
rect 0 7092 3122 7198
rect 0 7028 328 7092
rect 392 7028 3122 7092
rect 0 7012 3122 7028
rect 0 6948 328 7012
rect 392 6962 3122 7012
rect 3358 6962 5042 7198
rect 5278 6962 8400 7198
rect 392 6948 8400 6962
rect 0 6880 8400 6948
rect 0 6712 8400 6720
rect 0 6648 168 6712
rect 232 6648 328 6712
rect 392 6648 488 6712
rect 552 6648 648 6712
rect 712 6648 808 6712
rect 872 6648 968 6712
rect 1032 6648 1128 6712
rect 1192 6648 1448 6712
rect 1512 6648 1608 6712
rect 1672 6648 1768 6712
rect 1832 6648 1928 6712
rect 1992 6648 2088 6712
rect 2152 6648 2248 6712
rect 2312 6648 2408 6712
rect 2472 6648 2568 6712
rect 2632 6648 2728 6712
rect 2792 6648 2888 6712
rect 2952 6648 3048 6712
rect 3112 6648 3368 6712
rect 3432 6648 3528 6712
rect 3592 6648 3688 6712
rect 3752 6648 3848 6712
rect 3912 6648 4008 6712
rect 4072 6648 4168 6712
rect 4232 6648 4328 6712
rect 4392 6648 4488 6712
rect 4552 6648 4648 6712
rect 4712 6648 4808 6712
rect 4872 6648 4968 6712
rect 5032 6648 5288 6712
rect 5352 6648 5448 6712
rect 5512 6648 5608 6712
rect 5672 6648 5768 6712
rect 5832 6648 5928 6712
rect 5992 6648 6088 6712
rect 6152 6648 6248 6712
rect 6312 6648 6408 6712
rect 6472 6648 6568 6712
rect 6632 6648 6728 6712
rect 6792 6648 6888 6712
rect 6952 6648 7208 6712
rect 7272 6648 7368 6712
rect 7432 6648 7528 6712
rect 7592 6648 7688 6712
rect 7752 6648 7848 6712
rect 7912 6648 8168 6712
rect 8232 6648 8400 6712
rect 0 6638 8400 6648
rect 0 6552 3122 6638
rect 0 6488 168 6552
rect 232 6488 328 6552
rect 392 6488 488 6552
rect 552 6488 648 6552
rect 712 6488 808 6552
rect 872 6488 968 6552
rect 1032 6488 1128 6552
rect 1192 6488 1448 6552
rect 1512 6488 1608 6552
rect 1672 6488 1768 6552
rect 1832 6488 1928 6552
rect 1992 6488 2088 6552
rect 2152 6488 2248 6552
rect 2312 6488 2408 6552
rect 2472 6488 2568 6552
rect 2632 6488 2728 6552
rect 2792 6488 2888 6552
rect 2952 6488 3048 6552
rect 3112 6488 3122 6552
rect 0 6402 3122 6488
rect 3358 6552 5042 6638
rect 3358 6488 3368 6552
rect 3432 6488 3528 6552
rect 3592 6488 3688 6552
rect 3752 6488 3848 6552
rect 3912 6488 4008 6552
rect 4072 6488 4168 6552
rect 4232 6488 4328 6552
rect 4392 6488 4488 6552
rect 4552 6488 4648 6552
rect 4712 6488 4808 6552
rect 4872 6488 4968 6552
rect 5032 6488 5042 6552
rect 3358 6402 5042 6488
rect 5278 6552 8400 6638
rect 5278 6488 5288 6552
rect 5352 6488 5448 6552
rect 5512 6488 5608 6552
rect 5672 6488 5768 6552
rect 5832 6488 5928 6552
rect 5992 6488 6088 6552
rect 6152 6488 6248 6552
rect 6312 6488 6408 6552
rect 6472 6488 6568 6552
rect 6632 6488 6728 6552
rect 6792 6488 6888 6552
rect 6952 6488 7208 6552
rect 7272 6488 7368 6552
rect 7432 6488 7528 6552
rect 7592 6488 7688 6552
rect 7752 6488 7848 6552
rect 7912 6488 8168 6552
rect 8232 6488 8400 6552
rect 5278 6402 8400 6488
rect 0 6392 8400 6402
rect 0 6328 168 6392
rect 232 6328 328 6392
rect 392 6328 488 6392
rect 552 6328 648 6392
rect 712 6328 808 6392
rect 872 6328 968 6392
rect 1032 6328 1128 6392
rect 1192 6328 1448 6392
rect 1512 6328 1608 6392
rect 1672 6328 1768 6392
rect 1832 6328 1928 6392
rect 1992 6328 2088 6392
rect 2152 6328 2248 6392
rect 2312 6328 2408 6392
rect 2472 6328 2568 6392
rect 2632 6328 2728 6392
rect 2792 6328 2888 6392
rect 2952 6328 3048 6392
rect 3112 6328 3368 6392
rect 3432 6328 3528 6392
rect 3592 6328 3688 6392
rect 3752 6328 3848 6392
rect 3912 6328 4008 6392
rect 4072 6328 4168 6392
rect 4232 6328 4328 6392
rect 4392 6328 4488 6392
rect 4552 6328 4648 6392
rect 4712 6328 4808 6392
rect 4872 6328 4968 6392
rect 5032 6328 5288 6392
rect 5352 6328 5448 6392
rect 5512 6328 5608 6392
rect 5672 6328 5768 6392
rect 5832 6328 5928 6392
rect 5992 6328 6088 6392
rect 6152 6328 6248 6392
rect 6312 6328 6408 6392
rect 6472 6328 6568 6392
rect 6632 6328 6728 6392
rect 6792 6328 6888 6392
rect 6952 6328 7208 6392
rect 7272 6328 7368 6392
rect 7432 6328 7528 6392
rect 7592 6328 7688 6392
rect 7752 6328 7848 6392
rect 7912 6328 8168 6392
rect 8232 6328 8400 6392
rect 0 6320 8400 6328
rect 0 6232 8400 6240
rect 0 6168 168 6232
rect 232 6168 328 6232
rect 392 6168 488 6232
rect 552 6168 648 6232
rect 712 6168 808 6232
rect 872 6168 968 6232
rect 1032 6168 1128 6232
rect 1192 6168 1288 6232
rect 1352 6168 1448 6232
rect 1512 6168 1608 6232
rect 1672 6168 1768 6232
rect 1832 6168 1928 6232
rect 1992 6168 2088 6232
rect 2152 6168 2248 6232
rect 2312 6168 2408 6232
rect 2472 6168 2568 6232
rect 2632 6168 2728 6232
rect 2792 6168 2888 6232
rect 2952 6168 3048 6232
rect 3112 6168 3208 6232
rect 3272 6168 3368 6232
rect 3432 6168 3528 6232
rect 3592 6168 3688 6232
rect 3752 6168 3848 6232
rect 3912 6168 4008 6232
rect 4072 6168 4168 6232
rect 4232 6168 4328 6232
rect 4392 6168 4488 6232
rect 4552 6168 4648 6232
rect 4712 6168 4808 6232
rect 4872 6168 4968 6232
rect 5032 6168 5128 6232
rect 5192 6168 5288 6232
rect 5352 6168 5448 6232
rect 5512 6168 5608 6232
rect 5672 6168 5768 6232
rect 5832 6168 5928 6232
rect 5992 6168 6088 6232
rect 6152 6168 6248 6232
rect 6312 6168 6408 6232
rect 6472 6168 6568 6232
rect 6632 6168 6728 6232
rect 6792 6168 6888 6232
rect 6952 6168 7048 6232
rect 7112 6168 7208 6232
rect 7272 6168 7368 6232
rect 7432 6168 7528 6232
rect 7592 6168 7688 6232
rect 7752 6168 7848 6232
rect 7912 6168 8168 6232
rect 8232 6168 8400 6232
rect 0 6158 8400 6168
rect 0 6072 1202 6158
rect 1438 6072 6962 6158
rect 7198 6072 8400 6158
rect 0 6008 168 6072
rect 232 6008 328 6072
rect 392 6008 488 6072
rect 552 6008 648 6072
rect 712 6008 808 6072
rect 872 6008 968 6072
rect 1032 6008 1128 6072
rect 1192 6008 1202 6072
rect 1438 6008 1448 6072
rect 1512 6008 1608 6072
rect 1672 6008 1768 6072
rect 1832 6008 1928 6072
rect 1992 6008 2088 6072
rect 2152 6008 2248 6072
rect 2312 6008 2408 6072
rect 2472 6008 2568 6072
rect 2632 6008 2728 6072
rect 2792 6008 2888 6072
rect 2952 6008 3048 6072
rect 3112 6008 3208 6072
rect 3272 6008 3368 6072
rect 3432 6008 3528 6072
rect 3592 6008 3688 6072
rect 3752 6008 3848 6072
rect 3912 6008 4008 6072
rect 4072 6008 4168 6072
rect 4232 6008 4328 6072
rect 4392 6008 4488 6072
rect 4552 6008 4648 6072
rect 4712 6008 4808 6072
rect 4872 6008 4968 6072
rect 5032 6008 5128 6072
rect 5192 6008 5288 6072
rect 5352 6008 5448 6072
rect 5512 6008 5608 6072
rect 5672 6008 5768 6072
rect 5832 6008 5928 6072
rect 5992 6008 6088 6072
rect 6152 6008 6248 6072
rect 6312 6008 6408 6072
rect 6472 6008 6568 6072
rect 6632 6008 6728 6072
rect 6792 6008 6888 6072
rect 6952 6008 6962 6072
rect 7198 6008 7208 6072
rect 7272 6008 7368 6072
rect 7432 6008 7528 6072
rect 7592 6008 7688 6072
rect 7752 6008 7848 6072
rect 7912 6008 8168 6072
rect 8232 6008 8400 6072
rect 0 5922 1202 6008
rect 1438 5922 6962 6008
rect 7198 5922 8400 6008
rect 0 5912 8400 5922
rect 0 5848 168 5912
rect 232 5848 328 5912
rect 392 5848 488 5912
rect 552 5848 648 5912
rect 712 5848 808 5912
rect 872 5848 968 5912
rect 1032 5848 1128 5912
rect 1192 5848 1288 5912
rect 1352 5848 1448 5912
rect 1512 5848 1608 5912
rect 1672 5848 1768 5912
rect 1832 5848 1928 5912
rect 1992 5848 2088 5912
rect 2152 5848 2248 5912
rect 2312 5848 2408 5912
rect 2472 5848 2568 5912
rect 2632 5848 2728 5912
rect 2792 5848 2888 5912
rect 2952 5848 3048 5912
rect 3112 5848 3208 5912
rect 3272 5848 3368 5912
rect 3432 5848 3528 5912
rect 3592 5848 3688 5912
rect 3752 5848 3848 5912
rect 3912 5848 4008 5912
rect 4072 5848 4168 5912
rect 4232 5848 4328 5912
rect 4392 5848 4488 5912
rect 4552 5848 4648 5912
rect 4712 5848 4808 5912
rect 4872 5848 4968 5912
rect 5032 5848 5128 5912
rect 5192 5848 5288 5912
rect 5352 5848 5448 5912
rect 5512 5848 5608 5912
rect 5672 5848 5768 5912
rect 5832 5848 5928 5912
rect 5992 5848 6088 5912
rect 6152 5848 6248 5912
rect 6312 5848 6408 5912
rect 6472 5848 6568 5912
rect 6632 5848 6728 5912
rect 6792 5848 6888 5912
rect 6952 5848 7048 5912
rect 7112 5848 7208 5912
rect 7272 5848 7368 5912
rect 7432 5848 7528 5912
rect 7592 5848 7688 5912
rect 7752 5848 7848 5912
rect 7912 5848 8168 5912
rect 8232 5848 8400 5912
rect 0 5840 8400 5848
rect 0 5752 8400 5760
rect 0 5688 168 5752
rect 232 5688 328 5752
rect 392 5688 488 5752
rect 552 5688 648 5752
rect 712 5688 808 5752
rect 872 5688 968 5752
rect 1032 5688 1128 5752
rect 1192 5688 1448 5752
rect 1512 5688 1608 5752
rect 1672 5688 1768 5752
rect 1832 5688 1928 5752
rect 1992 5688 2088 5752
rect 2152 5688 2248 5752
rect 2312 5688 2408 5752
rect 2472 5688 2568 5752
rect 2632 5688 2728 5752
rect 2792 5688 2888 5752
rect 2952 5688 3048 5752
rect 3112 5688 3368 5752
rect 3432 5688 3528 5752
rect 3592 5688 3688 5752
rect 3752 5688 3848 5752
rect 3912 5688 4008 5752
rect 4072 5688 4168 5752
rect 4232 5688 4328 5752
rect 4392 5688 4488 5752
rect 4552 5688 4648 5752
rect 4712 5688 4808 5752
rect 4872 5688 4968 5752
rect 5032 5688 5288 5752
rect 5352 5688 5448 5752
rect 5512 5688 5608 5752
rect 5672 5688 5768 5752
rect 5832 5688 5928 5752
rect 5992 5688 6088 5752
rect 6152 5688 6248 5752
rect 6312 5688 6408 5752
rect 6472 5688 6568 5752
rect 6632 5688 6728 5752
rect 6792 5688 6888 5752
rect 6952 5688 7208 5752
rect 7272 5688 7368 5752
rect 7432 5688 7528 5752
rect 7592 5688 7688 5752
rect 7752 5688 7848 5752
rect 7912 5688 8168 5752
rect 8232 5688 8400 5752
rect 0 5678 8400 5688
rect 0 5592 242 5678
rect 478 5592 7922 5678
rect 0 5528 168 5592
rect 232 5528 242 5592
rect 478 5528 488 5592
rect 552 5528 648 5592
rect 712 5528 808 5592
rect 872 5528 968 5592
rect 1032 5528 1128 5592
rect 1192 5528 1448 5592
rect 1512 5528 1608 5592
rect 1672 5528 1768 5592
rect 1832 5528 1928 5592
rect 1992 5528 2088 5592
rect 2152 5528 2248 5592
rect 2312 5528 2408 5592
rect 2472 5528 2568 5592
rect 2632 5528 2728 5592
rect 2792 5528 2888 5592
rect 2952 5528 3048 5592
rect 3112 5528 3368 5592
rect 3432 5528 3528 5592
rect 3592 5528 3688 5592
rect 3752 5528 3848 5592
rect 3912 5528 4008 5592
rect 4072 5528 4168 5592
rect 4232 5528 4328 5592
rect 4392 5528 4488 5592
rect 4552 5528 4648 5592
rect 4712 5528 4808 5592
rect 4872 5528 4968 5592
rect 5032 5528 5288 5592
rect 5352 5528 5448 5592
rect 5512 5528 5608 5592
rect 5672 5528 5768 5592
rect 5832 5528 5928 5592
rect 5992 5528 6088 5592
rect 6152 5528 6248 5592
rect 6312 5528 6408 5592
rect 6472 5528 6568 5592
rect 6632 5528 6728 5592
rect 6792 5528 6888 5592
rect 6952 5528 7208 5592
rect 7272 5528 7368 5592
rect 7432 5528 7528 5592
rect 7592 5528 7688 5592
rect 7752 5528 7848 5592
rect 7912 5528 7922 5592
rect 0 5442 242 5528
rect 478 5442 7922 5528
rect 8158 5592 8400 5678
rect 8158 5528 8168 5592
rect 8232 5528 8400 5592
rect 8158 5442 8400 5528
rect 0 5432 8400 5442
rect 0 5368 168 5432
rect 232 5368 328 5432
rect 392 5368 488 5432
rect 552 5368 648 5432
rect 712 5368 808 5432
rect 872 5368 968 5432
rect 1032 5368 1128 5432
rect 1192 5368 1448 5432
rect 1512 5368 1608 5432
rect 1672 5368 1768 5432
rect 1832 5368 1928 5432
rect 1992 5368 2088 5432
rect 2152 5368 2248 5432
rect 2312 5368 2408 5432
rect 2472 5368 2568 5432
rect 2632 5368 2728 5432
rect 2792 5368 2888 5432
rect 2952 5368 3048 5432
rect 3112 5368 3368 5432
rect 3432 5368 3528 5432
rect 3592 5368 3688 5432
rect 3752 5368 3848 5432
rect 3912 5368 4008 5432
rect 4072 5368 4168 5432
rect 4232 5368 4328 5432
rect 4392 5368 4488 5432
rect 4552 5368 4648 5432
rect 4712 5368 4808 5432
rect 4872 5368 4968 5432
rect 5032 5368 5288 5432
rect 5352 5368 5448 5432
rect 5512 5368 5608 5432
rect 5672 5368 5768 5432
rect 5832 5368 5928 5432
rect 5992 5368 6088 5432
rect 6152 5368 6248 5432
rect 6312 5368 6408 5432
rect 6472 5368 6568 5432
rect 6632 5368 6728 5432
rect 6792 5368 6888 5432
rect 6952 5368 7208 5432
rect 7272 5368 7368 5432
rect 7432 5368 7528 5432
rect 7592 5368 7688 5432
rect 7752 5368 7848 5432
rect 7912 5368 8168 5432
rect 8232 5368 8400 5432
rect 0 5360 8400 5368
rect 0 4752 8400 4800
rect 0 4718 328 4752
rect 392 4718 8400 4752
rect 0 4482 242 4718
rect 478 4482 7922 4718
rect 8158 4482 8400 4718
rect 0 4448 328 4482
rect 392 4448 8400 4482
rect 0 4400 8400 4448
rect 0 3632 8400 3680
rect 0 3598 8008 3632
rect 8072 3598 8400 3632
rect 0 3362 242 3598
rect 478 3362 7922 3598
rect 8158 3362 8400 3598
rect 0 3328 8008 3362
rect 8072 3328 8400 3362
rect 0 3280 8400 3328
rect 0 2792 8400 2800
rect 0 2728 8 2792
rect 72 2728 168 2792
rect 232 2728 328 2792
rect 392 2728 488 2792
rect 552 2728 648 2792
rect 712 2728 808 2792
rect 872 2728 968 2792
rect 1032 2728 1128 2792
rect 1192 2728 1448 2792
rect 1512 2728 1608 2792
rect 1672 2728 1768 2792
rect 1832 2728 1928 2792
rect 1992 2728 2088 2792
rect 2152 2728 2248 2792
rect 2312 2728 2408 2792
rect 2472 2728 2568 2792
rect 2632 2728 2728 2792
rect 2792 2728 2888 2792
rect 2952 2728 3048 2792
rect 3112 2728 3368 2792
rect 3432 2728 3528 2792
rect 3592 2728 3688 2792
rect 3752 2728 3848 2792
rect 3912 2728 4008 2792
rect 4072 2728 4168 2792
rect 4232 2728 4328 2792
rect 4392 2728 4488 2792
rect 4552 2728 4648 2792
rect 4712 2728 4808 2792
rect 4872 2728 4968 2792
rect 5032 2728 5288 2792
rect 5352 2728 5448 2792
rect 5512 2728 5608 2792
rect 5672 2728 5768 2792
rect 5832 2728 5928 2792
rect 5992 2728 6088 2792
rect 6152 2728 6248 2792
rect 6312 2728 6408 2792
rect 6472 2728 6568 2792
rect 6632 2728 6728 2792
rect 6792 2728 6888 2792
rect 6952 2728 7208 2792
rect 7272 2728 7368 2792
rect 7432 2728 7528 2792
rect 7592 2728 7688 2792
rect 7752 2728 7848 2792
rect 7912 2728 8008 2792
rect 8072 2728 8168 2792
rect 8232 2728 8328 2792
rect 8392 2728 8400 2792
rect 0 2718 8400 2728
rect 0 2482 1202 2718
rect 1438 2482 6962 2718
rect 7198 2482 8400 2718
rect 0 2472 8400 2482
rect 0 2408 8 2472
rect 72 2408 168 2472
rect 232 2408 328 2472
rect 392 2408 488 2472
rect 552 2408 648 2472
rect 712 2408 808 2472
rect 872 2408 968 2472
rect 1032 2408 1128 2472
rect 1192 2408 1448 2472
rect 1512 2408 1608 2472
rect 1672 2408 1768 2472
rect 1832 2408 1928 2472
rect 1992 2408 2088 2472
rect 2152 2408 2248 2472
rect 2312 2408 2408 2472
rect 2472 2408 2568 2472
rect 2632 2408 2728 2472
rect 2792 2408 2888 2472
rect 2952 2408 3048 2472
rect 3112 2408 3368 2472
rect 3432 2408 3528 2472
rect 3592 2408 3688 2472
rect 3752 2408 3848 2472
rect 3912 2408 4008 2472
rect 4072 2408 4168 2472
rect 4232 2408 4328 2472
rect 4392 2408 4488 2472
rect 4552 2408 4648 2472
rect 4712 2408 4808 2472
rect 4872 2408 4968 2472
rect 5032 2408 5288 2472
rect 5352 2408 5448 2472
rect 5512 2408 5608 2472
rect 5672 2408 5768 2472
rect 5832 2408 5928 2472
rect 5992 2408 6088 2472
rect 6152 2408 6248 2472
rect 6312 2408 6408 2472
rect 6472 2408 6568 2472
rect 6632 2408 6728 2472
rect 6792 2408 6888 2472
rect 6952 2408 7208 2472
rect 7272 2408 7368 2472
rect 7432 2408 7528 2472
rect 7592 2408 7688 2472
rect 7752 2408 7848 2472
rect 7912 2408 8008 2472
rect 8072 2408 8168 2472
rect 8232 2408 8328 2472
rect 8392 2408 8400 2472
rect 0 2400 8400 2408
rect 0 1112 8400 1120
rect 0 1048 168 1112
rect 232 1048 328 1112
rect 392 1048 488 1112
rect 552 1048 648 1112
rect 712 1048 808 1112
rect 872 1048 968 1112
rect 1032 1048 1128 1112
rect 1192 1048 1448 1112
rect 1512 1048 1608 1112
rect 1672 1048 1768 1112
rect 1832 1048 1928 1112
rect 1992 1048 2088 1112
rect 2152 1048 2248 1112
rect 2312 1048 2408 1112
rect 2472 1048 2568 1112
rect 2632 1048 2728 1112
rect 2792 1048 2888 1112
rect 2952 1048 3048 1112
rect 3112 1048 3368 1112
rect 3432 1048 3528 1112
rect 3592 1048 3688 1112
rect 3752 1048 3848 1112
rect 3912 1048 4008 1112
rect 4072 1048 4168 1112
rect 4232 1048 4328 1112
rect 4392 1048 4488 1112
rect 4552 1048 4648 1112
rect 4712 1048 4808 1112
rect 4872 1048 4968 1112
rect 5032 1048 5288 1112
rect 5352 1048 5448 1112
rect 5512 1048 5608 1112
rect 5672 1048 5768 1112
rect 5832 1048 5928 1112
rect 5992 1048 6088 1112
rect 6152 1048 6248 1112
rect 6312 1048 6408 1112
rect 6472 1048 6568 1112
rect 6632 1048 6728 1112
rect 6792 1048 6888 1112
rect 6952 1048 7208 1112
rect 7272 1048 7368 1112
rect 7432 1048 7528 1112
rect 7592 1048 7688 1112
rect 7752 1048 7848 1112
rect 7912 1048 8168 1112
rect 8232 1048 8400 1112
rect 0 1038 8400 1048
rect 0 952 2162 1038
rect 2398 952 4082 1038
rect 4318 952 6002 1038
rect 6238 952 8400 1038
rect 0 888 168 952
rect 232 888 328 952
rect 392 888 488 952
rect 552 888 648 952
rect 712 888 808 952
rect 872 888 968 952
rect 1032 888 1128 952
rect 1192 888 1448 952
rect 1512 888 1608 952
rect 1672 888 1768 952
rect 1832 888 1928 952
rect 1992 888 2088 952
rect 2152 888 2162 952
rect 2398 888 2408 952
rect 2472 888 2568 952
rect 2632 888 2728 952
rect 2792 888 2888 952
rect 2952 888 3048 952
rect 3112 888 3368 952
rect 3432 888 3528 952
rect 3592 888 3688 952
rect 3752 888 3848 952
rect 3912 888 4008 952
rect 4072 888 4082 952
rect 4318 888 4328 952
rect 4392 888 4488 952
rect 4552 888 4648 952
rect 4712 888 4808 952
rect 4872 888 4968 952
rect 5032 888 5288 952
rect 5352 888 5448 952
rect 5512 888 5608 952
rect 5672 888 5768 952
rect 5832 888 5928 952
rect 5992 888 6002 952
rect 6238 888 6248 952
rect 6312 888 6408 952
rect 6472 888 6568 952
rect 6632 888 6728 952
rect 6792 888 6888 952
rect 6952 888 7208 952
rect 7272 888 7368 952
rect 7432 888 7528 952
rect 7592 888 7688 952
rect 7752 888 7848 952
rect 7912 888 8168 952
rect 8232 888 8400 952
rect 0 802 2162 888
rect 2398 802 4082 888
rect 4318 802 6002 888
rect 6238 802 8400 888
rect 0 792 8400 802
rect 0 728 168 792
rect 232 728 328 792
rect 392 728 488 792
rect 552 728 648 792
rect 712 728 808 792
rect 872 728 968 792
rect 1032 728 1128 792
rect 1192 728 1448 792
rect 1512 728 1608 792
rect 1672 728 1768 792
rect 1832 728 1928 792
rect 1992 728 2088 792
rect 2152 728 2248 792
rect 2312 728 2408 792
rect 2472 728 2568 792
rect 2632 728 2728 792
rect 2792 728 2888 792
rect 2952 728 3048 792
rect 3112 728 3368 792
rect 3432 728 3528 792
rect 3592 728 3688 792
rect 3752 728 3848 792
rect 3912 728 4008 792
rect 4072 728 4168 792
rect 4232 728 4328 792
rect 4392 728 4488 792
rect 4552 728 4648 792
rect 4712 728 4808 792
rect 4872 728 4968 792
rect 5032 728 5288 792
rect 5352 728 5448 792
rect 5512 728 5608 792
rect 5672 728 5768 792
rect 5832 728 5928 792
rect 5992 728 6088 792
rect 6152 728 6248 792
rect 6312 728 6408 792
rect 6472 728 6568 792
rect 6632 728 6728 792
rect 6792 728 6888 792
rect 6952 728 7208 792
rect 7272 728 7368 792
rect 7432 728 7528 792
rect 7592 728 7688 792
rect 7752 728 7848 792
rect 7912 728 8168 792
rect 8232 728 8400 792
rect 0 720 8400 728
rect 0 332 8400 400
rect 0 268 328 332
rect 392 318 8400 332
rect 392 268 3122 318
rect 0 252 3122 268
rect 0 188 328 252
rect 392 188 3122 252
rect 0 82 3122 188
rect 3358 82 5042 318
rect 5278 82 8400 318
rect 0 0 8400 82
rect 0 -88 8400 -80
rect 0 -152 168 -88
rect 232 -152 328 -88
rect 392 -152 488 -88
rect 552 -152 648 -88
rect 712 -152 808 -88
rect 872 -152 968 -88
rect 1032 -152 1128 -88
rect 1192 -152 1448 -88
rect 1512 -152 1608 -88
rect 1672 -152 1768 -88
rect 1832 -152 1928 -88
rect 1992 -152 2088 -88
rect 2152 -152 2248 -88
rect 2312 -152 2408 -88
rect 2472 -152 2568 -88
rect 2632 -152 2728 -88
rect 2792 -152 2888 -88
rect 2952 -152 3048 -88
rect 3112 -152 3368 -88
rect 3432 -152 3528 -88
rect 3592 -152 3688 -88
rect 3752 -152 3848 -88
rect 3912 -152 4008 -88
rect 4072 -152 4168 -88
rect 4232 -152 4328 -88
rect 4392 -152 4488 -88
rect 4552 -152 4648 -88
rect 4712 -152 4808 -88
rect 4872 -152 4968 -88
rect 5032 -152 5288 -88
rect 5352 -152 5448 -88
rect 5512 -152 5608 -88
rect 5672 -152 5768 -88
rect 5832 -152 5928 -88
rect 5992 -152 6088 -88
rect 6152 -152 6248 -88
rect 6312 -152 6408 -88
rect 6472 -152 6568 -88
rect 6632 -152 6728 -88
rect 6792 -152 6888 -88
rect 6952 -152 7208 -88
rect 7272 -152 7368 -88
rect 7432 -152 7528 -88
rect 7592 -152 7688 -88
rect 7752 -152 7848 -88
rect 7912 -152 8168 -88
rect 8232 -152 8400 -88
rect 0 -162 8400 -152
rect 0 -248 3122 -162
rect 0 -312 168 -248
rect 232 -312 328 -248
rect 392 -312 488 -248
rect 552 -312 648 -248
rect 712 -312 808 -248
rect 872 -312 968 -248
rect 1032 -312 1128 -248
rect 1192 -312 1448 -248
rect 1512 -312 1608 -248
rect 1672 -312 1768 -248
rect 1832 -312 1928 -248
rect 1992 -312 2088 -248
rect 2152 -312 2248 -248
rect 2312 -312 2408 -248
rect 2472 -312 2568 -248
rect 2632 -312 2728 -248
rect 2792 -312 2888 -248
rect 2952 -312 3048 -248
rect 3112 -312 3122 -248
rect 0 -398 3122 -312
rect 3358 -248 5042 -162
rect 3358 -312 3368 -248
rect 3432 -312 3528 -248
rect 3592 -312 3688 -248
rect 3752 -312 3848 -248
rect 3912 -312 4008 -248
rect 4072 -312 4168 -248
rect 4232 -312 4328 -248
rect 4392 -312 4488 -248
rect 4552 -312 4648 -248
rect 4712 -312 4808 -248
rect 4872 -312 4968 -248
rect 5032 -312 5042 -248
rect 3358 -398 5042 -312
rect 5278 -248 8400 -162
rect 5278 -312 5288 -248
rect 5352 -312 5448 -248
rect 5512 -312 5608 -248
rect 5672 -312 5768 -248
rect 5832 -312 5928 -248
rect 5992 -312 6088 -248
rect 6152 -312 6248 -248
rect 6312 -312 6408 -248
rect 6472 -312 6568 -248
rect 6632 -312 6728 -248
rect 6792 -312 6888 -248
rect 6952 -312 7208 -248
rect 7272 -312 7368 -248
rect 7432 -312 7528 -248
rect 7592 -312 7688 -248
rect 7752 -312 7848 -248
rect 7912 -312 8168 -248
rect 8232 -312 8400 -248
rect 5278 -398 8400 -312
rect 0 -408 8400 -398
rect 0 -472 168 -408
rect 232 -472 328 -408
rect 392 -472 488 -408
rect 552 -472 648 -408
rect 712 -472 808 -408
rect 872 -472 968 -408
rect 1032 -472 1128 -408
rect 1192 -472 1448 -408
rect 1512 -472 1608 -408
rect 1672 -472 1768 -408
rect 1832 -472 1928 -408
rect 1992 -472 2088 -408
rect 2152 -472 2248 -408
rect 2312 -472 2408 -408
rect 2472 -472 2568 -408
rect 2632 -472 2728 -408
rect 2792 -472 2888 -408
rect 2952 -472 3048 -408
rect 3112 -472 3368 -408
rect 3432 -472 3528 -408
rect 3592 -472 3688 -408
rect 3752 -472 3848 -408
rect 3912 -472 4008 -408
rect 4072 -472 4168 -408
rect 4232 -472 4328 -408
rect 4392 -472 4488 -408
rect 4552 -472 4648 -408
rect 4712 -472 4808 -408
rect 4872 -472 4968 -408
rect 5032 -472 5288 -408
rect 5352 -472 5448 -408
rect 5512 -472 5608 -408
rect 5672 -472 5768 -408
rect 5832 -472 5928 -408
rect 5992 -472 6088 -408
rect 6152 -472 6248 -408
rect 6312 -472 6408 -408
rect 6472 -472 6568 -408
rect 6632 -472 6728 -408
rect 6792 -472 6888 -408
rect 6952 -472 7208 -408
rect 7272 -472 7368 -408
rect 7432 -472 7528 -408
rect 7592 -472 7688 -408
rect 7752 -472 7848 -408
rect 7912 -472 8168 -408
rect 8232 -472 8400 -408
rect 0 -480 8400 -472
rect 0 -708 8400 -640
rect 0 -772 328 -708
rect 392 -722 8400 -708
rect 392 -772 3122 -722
rect 0 -788 3122 -772
rect 0 -852 328 -788
rect 392 -852 3122 -788
rect 0 -958 3122 -852
rect 3358 -958 5042 -722
rect 5278 -958 8400 -722
rect 0 -1040 8400 -958
<< via4 >>
rect 242 9648 328 9678
rect 328 9648 392 9678
rect 392 9648 478 9678
rect 242 9632 478 9648
rect 242 9568 328 9632
rect 328 9568 392 9632
rect 392 9568 478 9632
rect 242 9552 478 9568
rect 242 9488 328 9552
rect 328 9488 392 9552
rect 392 9488 478 9552
rect 242 9472 478 9488
rect 242 9442 328 9472
rect 328 9442 392 9472
rect 392 9442 478 9472
rect 7922 9442 8158 9678
rect 242 8632 478 8718
rect 7922 8632 8158 8718
rect 242 8568 328 8632
rect 328 8568 392 8632
rect 392 8568 478 8632
rect 7922 8568 8008 8632
rect 8008 8568 8072 8632
rect 8072 8568 8158 8632
rect 242 8482 478 8568
rect 7922 8482 8158 8568
rect 3122 8002 3358 8238
rect 5042 8002 5278 8238
rect 3122 7442 3358 7678
rect 5042 7442 5278 7678
rect 3122 6962 3358 7198
rect 5042 6962 5278 7198
rect 3122 6402 3358 6638
rect 5042 6402 5278 6638
rect 1202 6072 1438 6158
rect 6962 6072 7198 6158
rect 1202 6008 1288 6072
rect 1288 6008 1352 6072
rect 1352 6008 1438 6072
rect 6962 6008 7048 6072
rect 7048 6008 7112 6072
rect 7112 6008 7198 6072
rect 1202 5922 1438 6008
rect 6962 5922 7198 6008
rect 242 5592 478 5678
rect 242 5528 328 5592
rect 328 5528 392 5592
rect 392 5528 478 5592
rect 242 5442 478 5528
rect 7922 5442 8158 5678
rect 242 4688 328 4718
rect 328 4688 392 4718
rect 392 4688 478 4718
rect 242 4672 478 4688
rect 242 4608 328 4672
rect 328 4608 392 4672
rect 392 4608 478 4672
rect 242 4592 478 4608
rect 242 4528 328 4592
rect 328 4528 392 4592
rect 392 4528 478 4592
rect 242 4512 478 4528
rect 242 4482 328 4512
rect 328 4482 392 4512
rect 392 4482 478 4512
rect 7922 4482 8158 4718
rect 242 3362 478 3598
rect 7922 3568 8008 3598
rect 8008 3568 8072 3598
rect 8072 3568 8158 3598
rect 7922 3552 8158 3568
rect 7922 3488 8008 3552
rect 8008 3488 8072 3552
rect 8072 3488 8158 3552
rect 7922 3472 8158 3488
rect 7922 3408 8008 3472
rect 8008 3408 8072 3472
rect 8072 3408 8158 3472
rect 7922 3392 8158 3408
rect 7922 3362 8008 3392
rect 8008 3362 8072 3392
rect 8072 3362 8158 3392
rect 1202 2482 1438 2718
rect 6962 2482 7198 2718
rect 2162 952 2398 1038
rect 4082 952 4318 1038
rect 6002 952 6238 1038
rect 2162 888 2248 952
rect 2248 888 2312 952
rect 2312 888 2398 952
rect 4082 888 4168 952
rect 4168 888 4232 952
rect 4232 888 4318 952
rect 6002 888 6088 952
rect 6088 888 6152 952
rect 6152 888 6238 952
rect 2162 802 2398 888
rect 4082 802 4318 888
rect 6002 802 6238 888
rect 3122 82 3358 318
rect 5042 82 5278 318
rect 3122 -398 3358 -162
rect 5042 -398 5278 -162
rect 3122 -958 3358 -722
rect 5042 -958 5278 -722
<< metal5 >>
rect 160 9678 560 10080
rect 160 9442 242 9678
rect 478 9442 560 9678
rect 160 8718 560 9442
rect 160 8482 242 8718
rect 478 8482 560 8718
rect 160 5678 560 8482
rect 160 5442 242 5678
rect 478 5442 560 5678
rect 160 4718 560 5442
rect 160 4482 242 4718
rect 478 4482 560 4718
rect 160 3598 560 4482
rect 160 3362 242 3598
rect 478 3362 560 3598
rect 160 -1040 560 3362
rect 1120 6158 1520 10080
rect 1120 5922 1202 6158
rect 1438 5922 1520 6158
rect 1120 2718 1520 5922
rect 1120 2482 1202 2718
rect 1438 2482 1520 2718
rect 1120 -1040 1520 2482
rect 2080 1038 2480 10080
rect 2080 802 2162 1038
rect 2398 802 2480 1038
rect 2080 -1040 2480 802
rect 3040 8238 3440 10080
rect 3040 8002 3122 8238
rect 3358 8002 3440 8238
rect 3040 7678 3440 8002
rect 3040 7442 3122 7678
rect 3358 7442 3440 7678
rect 3040 7198 3440 7442
rect 3040 6962 3122 7198
rect 3358 6962 3440 7198
rect 3040 6638 3440 6962
rect 3040 6402 3122 6638
rect 3358 6402 3440 6638
rect 3040 318 3440 6402
rect 3040 82 3122 318
rect 3358 82 3440 318
rect 3040 -162 3440 82
rect 3040 -398 3122 -162
rect 3358 -398 3440 -162
rect 3040 -722 3440 -398
rect 3040 -958 3122 -722
rect 3358 -958 3440 -722
rect 3040 -1040 3440 -958
rect 4000 1038 4400 10080
rect 4000 802 4082 1038
rect 4318 802 4400 1038
rect 4000 -1040 4400 802
rect 4960 8238 5360 10080
rect 4960 8002 5042 8238
rect 5278 8002 5360 8238
rect 4960 7678 5360 8002
rect 4960 7442 5042 7678
rect 5278 7442 5360 7678
rect 4960 7198 5360 7442
rect 4960 6962 5042 7198
rect 5278 6962 5360 7198
rect 4960 6638 5360 6962
rect 4960 6402 5042 6638
rect 5278 6402 5360 6638
rect 4960 318 5360 6402
rect 4960 82 5042 318
rect 5278 82 5360 318
rect 4960 -162 5360 82
rect 4960 -398 5042 -162
rect 5278 -398 5360 -162
rect 4960 -722 5360 -398
rect 4960 -958 5042 -722
rect 5278 -958 5360 -722
rect 4960 -1040 5360 -958
rect 5920 1038 6320 10080
rect 5920 802 6002 1038
rect 6238 802 6320 1038
rect 5920 -1040 6320 802
rect 6880 6158 7280 10080
rect 6880 5922 6962 6158
rect 7198 5922 7280 6158
rect 6880 2718 7280 5922
rect 6880 2482 6962 2718
rect 7198 2482 7280 2718
rect 6880 -1040 7280 2482
rect 7840 9678 8240 10080
rect 7840 9442 7922 9678
rect 8158 9442 8240 9678
rect 7840 8718 8240 9442
rect 7840 8482 7922 8718
rect 8158 8482 8240 8718
rect 7840 5678 8240 8482
rect 7840 5442 7922 5678
rect 8158 5442 8240 5678
rect 7840 4718 8240 5442
rect 7840 4482 7922 4718
rect 8158 4482 8240 4718
rect 7840 3598 8240 4482
rect 7840 3362 7922 3598
rect 8158 3362 8240 3598
rect 7840 -1040 8240 3362
<< labels >>
rlabel metal1 s 2240 -880 2320 -680 4 na1
rlabel metal1 s 4160 -880 4240 -680 4 na2
rlabel metal1 s 6080 -880 6160 -680 4 na3
rlabel metal1 s 2240 160 2320 360 4 qa1
rlabel metal1 s 4160 160 4240 360 4 qa2
rlabel metal1 s 6080 160 6160 360 4 qa3
rlabel metal1 s 6080 1640 6160 2240 4 qa4
rlabel metal1 s 4160 1640 4240 2240 4 qa5
rlabel metal1 s 2240 1640 2320 2240 4 qa6
rlabel metal1 s 6080 3080 6160 3680 4 bpa1
rlabel metal1 s 4160 3080 4240 3680 4 bpa2
rlabel metal1 s 2240 3080 2320 3680 4 bpa3
rlabel metal1 s 2240 4400 2320 5000 4 xa1
rlabel metal1 s 4160 4400 4240 5000 4 xa2
rlabel metal1 s 6080 4400 6160 5000 4 xa3
rlabel metal1 s 2240 6920 2320 7120 4 nb1
rlabel metal1 s 4160 6920 4240 7120 4 nb2
rlabel metal1 s 6080 6920 6160 7120 4 nb3
rlabel metal1 s 2240 7520 2320 7720 4 qb1
rlabel metal1 s 4160 7520 4240 7720 4 qb2
rlabel metal1 s 6080 7520 6160 7720 4 qb3
rlabel metal1 s 2240 9160 2320 9760 4 xb1
rlabel metal1 s 4160 9160 4240 9760 4 xb2
rlabel metal1 s 6080 9160 6160 9760 4 xb3
rlabel metal2 s 0 2560 8400 2640 4 bpa
port 1 nsew
rlabel metal2 s 0 6000 8400 6080 4 bpb
port 2 nsew
rlabel metal5 s 2080 -1040 2480 10080 4 gnda
port 3 nsew
rlabel metal2 s 0 -320 8400 -240 4 na
port 4 nsew
rlabel metal2 s 0 6480 8400 6560 4 nb
port 5 nsew
rlabel metal2 s 0 720 8400 800 4 qa
port 6 nsew
rlabel metal2 s 0 8080 8400 8160 4 qb
port 7 nsew
rlabel metal5 s 160 -1040 560 10080 4 vdda
port 8 nsew
rlabel metal5 s 1120 -1040 1520 10080 4 vddx
port 9 nsew
rlabel metal5 s 3040 -1040 3440 10080 4 vssa
port 10 nsew
rlabel metal2 s 0 5520 8400 5600 4 xa
port 11 nsew
rlabel metal2 s 0 8560 8400 8640 4 xb
port 12 nsew
<< end >>
