magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< error_s >>
rect 8 66691 8392 66712
rect 12488 66691 20872 66712
rect 8 66657 8377 66691
rect 12503 66657 20872 66691
rect 8 66640 8392 66657
rect 8 66560 80 66640
rect 94 66600 8306 66626
rect 94 65480 120 66600
rect 160 66534 8240 66560
rect 160 65592 232 66534
rect 8214 65592 8240 66534
rect 160 65520 8240 65592
rect 8280 65480 8306 66600
rect 8320 65520 8392 66640
rect 12488 66640 20872 66657
rect 12488 66560 12560 66640
rect 12574 66600 20786 66626
rect 94 65454 8306 65480
rect 12574 65480 12600 66600
rect 12640 66534 20720 66560
rect 12640 65592 12712 66534
rect 20694 65592 20720 66534
rect 12640 65520 20720 65592
rect 20760 65480 20786 66600
rect 20800 65520 20872 66640
rect 21048 66640 22300 66712
rect 21048 66560 21120 66640
rect 21134 66600 22300 66626
rect 12574 65454 20786 65480
rect 21134 65480 21160 66600
rect 21200 66534 22300 66560
rect 21200 65592 21272 66534
rect 21200 65520 22300 65592
rect 21134 65454 22300 65480
rect 8 65200 8392 65272
rect 8 65120 80 65200
rect 94 65160 8306 65186
rect 94 64040 120 65160
rect 160 65094 8240 65120
rect 160 64152 232 65094
rect 8214 64152 8240 65094
rect 160 64080 8240 64152
rect 8280 64040 8306 65160
rect 8320 64080 8392 65200
rect 12488 65200 20872 65272
rect 12488 65120 12560 65200
rect 12574 65160 20786 65186
rect 94 64014 8306 64040
rect 12574 64040 12600 65160
rect 12640 65094 20720 65120
rect 12640 64152 12712 65094
rect 20694 64152 20720 65094
rect 12640 64080 20720 64152
rect 20760 64040 20786 65160
rect 20800 64080 20872 65200
rect 21048 65200 22300 65272
rect 21048 65120 21120 65200
rect 21134 65160 22300 65186
rect 12574 64014 20786 64040
rect 21134 64040 21160 65160
rect 21200 65094 22300 65120
rect 21200 64152 21272 65094
rect 21200 64080 22300 64152
rect 21134 64014 22300 64040
rect 8 63760 8392 63832
rect 8 63680 80 63760
rect 94 63720 8306 63746
rect 94 62600 120 63720
rect 160 63654 8240 63680
rect 160 62712 232 63654
rect 8214 62712 8240 63654
rect 160 62640 8240 62712
rect 8280 62600 8306 63720
rect 8320 62640 8392 63760
rect 12488 63760 20872 63832
rect 12488 63680 12560 63760
rect 12574 63720 20786 63746
rect 94 62574 8306 62600
rect 12574 62600 12600 63720
rect 12640 63654 20720 63680
rect 12640 62712 12712 63654
rect 20694 62712 20720 63654
rect 12640 62640 20720 62712
rect 20760 62600 20786 63720
rect 20800 62640 20872 63760
rect 21048 63760 22300 63832
rect 21048 63680 21120 63760
rect 21134 63720 22300 63746
rect 12574 62574 20786 62600
rect 21134 62600 21160 63720
rect 21200 63654 22300 63680
rect 21200 62712 21272 63654
rect 21200 62640 22300 62712
rect 21134 62574 22300 62600
rect 19754 59120 20872 59192
rect 19754 59080 20786 59106
rect 19754 59014 20720 59040
rect 20694 58072 20720 59014
rect 19754 58000 20720 58072
rect 20760 57960 20786 59080
rect 20800 58000 20872 59120
rect 21048 59120 22166 59192
rect 21048 59040 21120 59120
rect 21134 59080 22166 59106
rect 19754 57934 20786 57960
rect 21134 57960 21160 59080
rect 21200 59014 22166 59040
rect 21200 58072 21272 59014
rect 21200 58000 22166 58072
rect 21134 57934 22166 57960
rect 19754 56480 20872 56552
rect 19754 56440 20786 56466
rect 19754 56374 20720 56400
rect 20694 55432 20720 56374
rect 19754 55360 20720 55432
rect 20760 55320 20786 56440
rect 20800 55360 20872 56480
rect 21048 56480 22166 56552
rect 21048 56400 21120 56480
rect 21134 56440 22166 56466
rect 19754 55294 20786 55320
rect 21134 55320 21160 56440
rect 21200 56374 22166 56400
rect 21200 55432 21272 56374
rect 21200 55360 22166 55432
rect 21134 55294 22166 55320
rect 19754 55040 20872 55112
rect 19754 55000 20786 55026
rect 19754 54934 20720 54960
rect 20694 53992 20720 54934
rect 19754 53920 20720 53992
rect 20760 53880 20786 55000
rect 20800 53920 20872 55040
rect 21048 55040 22166 55112
rect 21048 54960 21120 55040
rect 21134 55000 22166 55026
rect 19754 53854 20786 53880
rect 21134 53880 21160 55000
rect 21200 54934 22166 54960
rect 21200 53992 21272 54934
rect 21200 53920 22166 53992
rect 21134 53854 22166 53880
rect 19754 53600 20872 53672
rect 19754 53560 20786 53586
rect 19754 53494 20720 53520
rect 20694 52552 20720 53494
rect 19754 52480 20720 52552
rect 20760 52440 20786 53560
rect 20800 52480 20872 53600
rect 21048 53600 22166 53672
rect 21048 53520 21120 53600
rect 21134 53560 22166 53586
rect 19754 52414 20786 52440
rect 21134 52440 21160 53560
rect 21200 53494 22166 53520
rect 21200 52552 21272 53494
rect 21200 52480 22166 52552
rect 21134 52414 22166 52440
rect 19754 52160 20872 52232
rect 19754 52120 20786 52146
rect 19754 52054 20720 52080
rect 20694 51112 20720 52054
rect 19754 51040 20720 51112
rect 20760 51000 20786 52120
rect 20800 51040 20872 52160
rect 21048 52160 22166 52232
rect 21048 52080 21120 52160
rect 21134 52120 22166 52146
rect 19754 50974 20786 51000
rect 21134 51000 21160 52120
rect 21200 52054 22166 52080
rect 21200 51112 21272 52054
rect 21200 51040 22166 51112
rect 21134 50974 22166 51000
rect 19754 48320 20872 48392
rect 19754 48280 20786 48306
rect 19754 48214 20720 48240
rect 20694 47272 20720 48214
rect 19754 47200 20720 47272
rect 20760 47160 20786 48280
rect 20800 47200 20872 48320
rect 21048 48320 22166 48392
rect 21048 48240 21120 48320
rect 21134 48280 22166 48306
rect 19754 47134 20786 47160
rect 21134 47160 21160 48280
rect 21200 48214 22166 48240
rect 21200 47272 21272 48214
rect 21200 47200 22166 47272
rect 21134 47134 22166 47160
rect 19754 46880 20872 46952
rect 19754 46840 20786 46866
rect 19754 46774 20720 46800
rect 20694 45832 20720 46774
rect 19754 45760 20720 45832
rect 20760 45720 20786 46840
rect 20800 45760 20872 46880
rect 21048 46880 22166 46952
rect 21048 46800 21120 46880
rect 21134 46840 22166 46866
rect 19754 45694 20786 45720
rect 21134 45720 21160 46840
rect 21200 46774 22166 46800
rect 21200 45832 21272 46774
rect 21200 45760 22166 45832
rect 21134 45694 22166 45720
rect 19754 45440 20872 45512
rect 19754 45400 20786 45426
rect 19754 45334 20720 45360
rect 20694 44392 20720 45334
rect 19754 44320 20720 44392
rect 20760 44280 20786 45400
rect 20800 44320 20872 45440
rect 21048 45440 22166 45512
rect 21048 45360 21120 45440
rect 21134 45400 22166 45426
rect 19754 44254 20786 44280
rect 21134 44280 21160 45400
rect 21200 45334 22166 45360
rect 21200 44392 21272 45334
rect 21200 44320 22166 44392
rect 21134 44254 22166 44280
rect 19754 44000 20872 44072
rect 19754 43960 20786 43986
rect 19754 43894 20720 43920
rect 20694 42952 20720 43894
rect 19754 42880 20720 42952
rect 20760 42840 20786 43960
rect 20800 42880 20872 44000
rect 21048 44000 22166 44072
rect 21048 43920 21120 44000
rect 21134 43960 22166 43986
rect 19754 42814 20786 42840
rect 21134 42840 21160 43960
rect 21200 43894 22166 43920
rect 21200 42952 21272 43894
rect 21200 42880 22166 42952
rect 21134 42814 22166 42840
rect 8 40160 8392 40232
rect 8 40080 80 40160
rect 94 40120 8306 40146
rect 94 39000 120 40120
rect 160 40054 8240 40080
rect 160 39112 232 40054
rect 8214 39112 8240 40054
rect 160 39040 8240 39112
rect 8280 39000 8306 40120
rect 8320 39040 8392 40160
rect 12488 40160 20872 40232
rect 12488 40080 12560 40160
rect 12574 40120 20786 40146
rect 94 38974 8306 39000
rect 12574 39000 12600 40120
rect 12640 40054 20720 40080
rect 12640 39112 12712 40054
rect 20694 39112 20720 40054
rect 12640 39040 20720 39112
rect 20760 39000 20786 40120
rect 20800 39040 20872 40160
rect 21048 40160 29432 40232
rect 21048 40080 21120 40160
rect 21134 40120 29346 40146
rect 12574 38974 20786 39000
rect 21134 39000 21160 40120
rect 21200 40054 29280 40080
rect 21200 39112 21272 40054
rect 29254 39112 29280 40054
rect 21200 39040 29280 39112
rect 29320 39000 29346 40120
rect 29360 39040 29432 40160
rect 33528 40160 40320 40232
rect 33528 40080 33600 40160
rect 33614 40120 40320 40146
rect 21134 38974 29346 39000
rect 33614 39000 33640 40120
rect 33680 40054 40320 40080
rect 33680 39112 33752 40054
rect 33680 39040 40320 39112
rect 33614 38974 40320 39000
rect 8 38720 8392 38792
rect 8 38640 80 38720
rect 94 38680 8306 38706
rect 94 37560 120 38680
rect 160 38614 8240 38640
rect 160 37672 232 38614
rect 8214 37672 8240 38614
rect 160 37600 8240 37672
rect 8280 37560 8306 38680
rect 8320 37600 8392 38720
rect 12488 38720 20872 38792
rect 12488 38640 12560 38720
rect 12574 38680 20786 38706
rect 94 37534 8306 37560
rect 12574 37560 12600 38680
rect 12640 38614 20720 38640
rect 12640 37672 12712 38614
rect 20694 37672 20720 38614
rect 12640 37600 20720 37672
rect 20760 37560 20786 38680
rect 20800 37600 20872 38720
rect 21048 38720 29432 38792
rect 21048 38640 21120 38720
rect 21134 38680 29346 38706
rect 12574 37534 20786 37560
rect 21134 37560 21160 38680
rect 21200 38614 29280 38640
rect 21200 37672 21272 38614
rect 29254 37672 29280 38614
rect 21200 37600 29280 37672
rect 29320 37560 29346 38680
rect 29360 37600 29432 38720
rect 33528 38720 40320 38792
rect 33528 38640 33600 38720
rect 33614 38680 40320 38706
rect 21134 37534 29346 37560
rect 33614 37560 33640 38680
rect 33680 38620 40320 38640
rect 33680 38614 41760 38620
rect 33680 37672 33752 38614
rect 41734 37672 41760 38614
rect 33680 37600 41760 37672
rect 41800 37560 41826 38620
rect 41840 37600 41912 38620
rect 33614 37534 41826 37560
rect 8 29280 8392 29352
rect 8 29200 80 29280
rect 94 29240 8306 29266
rect 94 28120 120 29240
rect 160 29174 8240 29200
rect 160 28232 232 29174
rect 8214 28232 8240 29174
rect 160 28160 8240 28232
rect 8280 28120 8306 29240
rect 8320 28160 8392 29280
rect 12488 29280 20872 29352
rect 12488 29200 12560 29280
rect 12574 29240 20786 29266
rect 94 28094 8306 28120
rect 12574 28120 12600 29240
rect 12640 29174 20720 29200
rect 12640 28232 12712 29174
rect 20694 28232 20720 29174
rect 12640 28160 20720 28232
rect 20760 28120 20786 29240
rect 20800 28160 20872 29280
rect 21048 29280 29432 29352
rect 21048 29200 21120 29280
rect 21134 29240 29346 29266
rect 12574 28094 20786 28120
rect 21134 28120 21160 29240
rect 21200 29174 29280 29200
rect 21200 28232 21272 29174
rect 29254 28232 29280 29174
rect 21200 28160 29280 28232
rect 29320 28120 29346 29240
rect 29360 28160 29432 29280
rect 33528 29280 41912 29352
rect 33528 29200 33600 29280
rect 33614 29240 41826 29266
rect 21134 28094 29346 28120
rect 33614 28120 33640 29240
rect 33680 29174 41760 29200
rect 33680 28232 33752 29174
rect 41734 28232 41760 29174
rect 33680 28180 41760 28232
rect 41800 28180 41826 29240
rect 41840 28180 41912 29280
rect 33680 28160 40320 28180
rect 33614 28094 40320 28120
rect 8 27840 8392 27912
rect 8 27760 80 27840
rect 94 27800 8306 27826
rect 94 26680 120 27800
rect 160 27734 8240 27760
rect 160 26792 232 27734
rect 8214 26792 8240 27734
rect 160 26720 8240 26792
rect 8280 26680 8306 27800
rect 8320 26720 8392 27840
rect 12488 27840 20872 27912
rect 12488 27760 12560 27840
rect 12574 27800 20786 27826
rect 94 26654 8306 26680
rect 12574 26680 12600 27800
rect 12640 27734 20720 27760
rect 12640 26792 12712 27734
rect 20694 26792 20720 27734
rect 12640 26720 20720 26792
rect 20760 26680 20786 27800
rect 20800 26720 20872 27840
rect 21048 27840 29432 27912
rect 21048 27760 21120 27840
rect 21134 27800 29346 27826
rect 12574 26654 20786 26680
rect 21134 26680 21160 27800
rect 21200 27734 29280 27760
rect 21200 26792 21272 27734
rect 29254 26792 29280 27734
rect 21200 26720 29280 26792
rect 29320 26680 29346 27800
rect 29360 26720 29432 27840
rect 33528 27840 40320 27912
rect 33528 27760 33600 27840
rect 33614 27800 40320 27826
rect 21134 26654 29346 26680
rect 33614 26680 33640 27800
rect 33680 27734 40320 27760
rect 33680 26792 33752 27734
rect 33680 26720 40320 26792
rect 33614 26654 40320 26680
rect 8 24000 8392 24072
rect 8 23920 80 24000
rect 94 23960 8306 23986
rect 94 22840 120 23960
rect 160 23894 8240 23920
rect 160 22952 232 23894
rect 8214 22952 8240 23894
rect 160 22880 8240 22952
rect 8280 22840 8306 23960
rect 8320 22880 8392 24000
rect 12488 24000 20872 24072
rect 12488 23920 12560 24000
rect 12574 23960 20786 23986
rect 94 22814 8306 22840
rect 12574 22840 12600 23960
rect 12640 23894 20720 23920
rect 12640 22952 12712 23894
rect 20694 22952 20720 23894
rect 12640 22880 20720 22952
rect 20760 22840 20786 23960
rect 20800 22880 20872 24000
rect 21048 24000 29432 24072
rect 21048 23920 21120 24000
rect 21134 23960 29346 23986
rect 12574 22814 20786 22840
rect 21134 22840 21160 23960
rect 21200 23894 29280 23920
rect 21200 22952 21272 23894
rect 29254 22952 29280 23894
rect 21200 22880 29280 22952
rect 29320 22840 29346 23960
rect 29360 22880 29432 24000
rect 33528 24000 40320 24072
rect 33528 23920 33600 24000
rect 33614 23960 40320 23986
rect 21134 22814 29346 22840
rect 33614 22840 33640 23960
rect 33680 23894 40320 23920
rect 33680 22952 33752 23894
rect 33680 22880 40320 22952
rect 33614 22814 40320 22840
rect 8 22560 8392 22632
rect 8 22480 80 22560
rect 94 22520 8306 22546
rect 94 21400 120 22520
rect 160 22454 8240 22480
rect 160 21512 232 22454
rect 8214 21512 8240 22454
rect 160 21440 8240 21512
rect 8280 21400 8306 22520
rect 8320 21440 8392 22560
rect 12488 22560 20872 22632
rect 12488 22480 12560 22560
rect 12574 22520 20786 22546
rect 94 21374 8306 21400
rect 12574 21400 12600 22520
rect 12640 22454 20720 22480
rect 12640 21512 12712 22454
rect 20694 21512 20720 22454
rect 12640 21440 20720 21512
rect 20760 21400 20786 22520
rect 20800 21440 20872 22560
rect 21048 22560 29432 22632
rect 21048 22480 21120 22560
rect 21134 22520 29346 22546
rect 12574 21374 20786 21400
rect 21134 21400 21160 22520
rect 21200 22454 29280 22480
rect 21200 21512 21272 22454
rect 29254 21512 29280 22454
rect 21200 21440 29280 21512
rect 29320 21400 29346 22520
rect 29360 21440 29432 22560
rect 33528 22560 40320 22632
rect 33528 22480 33600 22560
rect 33614 22520 40320 22546
rect 21134 21374 29346 21400
rect 33614 21400 33640 22520
rect 33680 22454 40320 22480
rect 33680 21512 33752 22454
rect 33680 21440 40320 21512
rect 33614 21374 40320 21400
rect 8 21120 8392 21192
rect 8 21040 80 21120
rect 94 21080 8306 21106
rect 94 20160 120 21080
rect 160 21014 8240 21040
rect 160 20160 232 21014
rect 8214 20160 8240 21014
rect 8280 20160 8306 21080
rect 8320 20160 8392 21120
rect 12488 21120 20872 21192
rect 12488 21040 12560 21120
rect 12574 21080 20786 21106
rect 12574 20160 12600 21080
rect 12640 21014 20720 21040
rect 12640 20160 12712 21014
rect 20694 20072 20720 21014
rect 19754 20000 20720 20072
rect 20760 19960 20786 21080
rect 20800 20000 20872 21120
rect 21048 21120 29432 21192
rect 21048 21040 21120 21120
rect 21134 21080 29346 21106
rect 19754 19934 20786 19960
rect 21134 19960 21160 21080
rect 21200 21014 29280 21040
rect 21200 20072 21272 21014
rect 29254 20160 29280 21014
rect 29320 20160 29346 21080
rect 29360 20160 29432 21120
rect 33528 21120 40320 21192
rect 33528 21040 33600 21120
rect 33614 21080 40320 21106
rect 33614 20160 33640 21080
rect 33680 21014 40320 21040
rect 33680 20160 33752 21014
rect 21200 20000 22166 20072
rect 21134 19934 22166 19960
rect 19754 19680 20872 19752
rect 19754 19640 20786 19666
rect 19754 19574 20720 19600
rect 20694 18632 20720 19574
rect 19754 18560 20720 18632
rect 20760 18520 20786 19640
rect 20800 18560 20872 19680
rect 21048 19680 22166 19752
rect 21048 19600 21120 19680
rect 21134 19640 22166 19666
rect 19754 18494 20786 18520
rect 21134 18520 21160 19640
rect 21200 19574 22166 19600
rect 21200 18632 21272 19574
rect 21200 18560 22166 18632
rect 21134 18494 22166 18520
rect 19754 15840 20872 15912
rect 19754 15800 20786 15826
rect 19754 15734 20720 15760
rect 20694 14792 20720 15734
rect 19754 14720 20720 14792
rect 20760 14680 20786 15800
rect 20800 14720 20872 15840
rect 21048 15840 22166 15912
rect 21048 15760 21120 15840
rect 21134 15800 22166 15826
rect 19754 14654 20786 14680
rect 21134 14680 21160 15800
rect 21200 15734 22166 15760
rect 21200 14792 21272 15734
rect 21200 14720 22166 14792
rect 21134 14654 22166 14680
rect 19754 14400 20872 14472
rect 19754 14360 20786 14386
rect 19754 14294 20720 14320
rect 20694 13352 20720 14294
rect 19754 13280 20720 13352
rect 20760 13240 20786 14360
rect 20800 13280 20872 14400
rect 21048 14400 22166 14472
rect 21048 14320 21120 14400
rect 21134 14360 22166 14386
rect 19754 13214 20786 13240
rect 21134 13240 21160 14360
rect 21200 14294 22166 14320
rect 21200 13352 21272 14294
rect 21200 13280 22166 13352
rect 21134 13214 22166 13240
rect 19754 12960 20872 13032
rect 19754 12920 20786 12946
rect 19754 12854 20720 12880
rect 20694 11912 20720 12854
rect 19754 11840 20720 11912
rect 20760 11800 20786 12920
rect 20800 11840 20872 12960
rect 21048 12960 22166 13032
rect 21048 12880 21120 12960
rect 21134 12920 22166 12946
rect 19754 11774 20786 11800
rect 21134 11800 21160 12920
rect 21200 12854 22166 12880
rect 21200 11912 21272 12854
rect 21200 11840 22166 11912
rect 21134 11774 22166 11800
rect 19754 11520 20872 11592
rect 19754 11480 20786 11506
rect 19754 11414 20720 11440
rect 20694 10472 20720 11414
rect 19754 10400 20720 10472
rect 20760 10360 20786 11480
rect 20800 10400 20872 11520
rect 21048 11520 22166 11592
rect 21048 11440 21120 11520
rect 21134 11480 22166 11506
rect 19754 10334 20786 10360
rect 21134 10360 21160 11480
rect 21200 11414 22166 11440
rect 21200 10472 21272 11414
rect 21200 10400 22166 10472
rect 21134 10334 22166 10360
rect 19754 8880 20872 8952
rect 19754 8840 20786 8866
rect 19754 8774 20720 8800
rect 20694 7832 20720 8774
rect 19754 7760 20720 7832
rect 20760 7720 20786 8840
rect 20800 7760 20872 8880
rect 21048 8880 22166 8952
rect 21048 8800 21120 8880
rect 21134 8840 22166 8866
rect 19754 7694 20786 7720
rect 21134 7720 21160 8840
rect 21200 8774 22166 8800
rect 21200 7832 21272 8774
rect 21200 7760 22166 7832
rect 21134 7694 22166 7720
rect 19754 4240 20872 4312
rect 19754 4200 20786 4226
rect 19754 4134 20720 4160
rect 20694 3192 20720 4134
rect 19754 3120 20720 3192
rect 20760 3080 20786 4200
rect 20800 3120 20872 4240
rect 21048 4240 22166 4312
rect 21048 4160 21120 4240
rect 21134 4200 22166 4226
rect 19754 3054 20786 3080
rect 21134 3080 21160 4200
rect 21200 4134 22166 4160
rect 21200 3192 21272 4134
rect 21200 3120 22166 3192
rect 21134 3054 22166 3080
rect 19754 2800 20872 2872
rect 19754 2760 20786 2786
rect 19754 2694 20720 2720
rect 20694 1752 20720 2694
rect 19754 1680 20720 1752
rect 20760 1640 20786 2760
rect 20800 1680 20872 2800
rect 21048 2800 22166 2872
rect 21048 2720 21120 2800
rect 21134 2760 22166 2786
rect 19754 1614 20786 1640
rect 21134 1640 21160 2760
rect 21200 2694 22166 2720
rect 21200 1752 21272 2694
rect 21200 1680 22166 1752
rect 21134 1614 22166 1640
rect 19754 1360 20872 1432
rect 19754 1320 20786 1346
rect 19754 1254 20720 1280
rect 20694 312 20720 1254
rect 19754 240 20720 312
rect 20760 200 20786 1320
rect 20800 240 20872 1360
rect 21048 1360 22166 1432
rect 21048 1280 21120 1360
rect 21134 1320 22166 1346
rect 19754 174 20786 200
rect 21134 200 21160 1320
rect 21200 1254 22166 1280
rect 21200 312 21272 1254
rect 21200 240 22166 312
rect 21134 174 22166 200
<< locali >>
rect 0 37337 80 37360
rect 0 37303 23 37337
rect 57 37303 80 37337
rect 0 37017 80 37303
rect 0 36983 23 37017
rect 57 36983 80 37017
rect 0 36960 80 36983
rect 160 37337 240 37360
rect 160 37303 183 37337
rect 217 37303 240 37337
rect 160 37017 240 37303
rect 160 36983 183 37017
rect 217 36983 240 37017
rect 160 36960 240 36983
rect 320 37337 400 37360
rect 320 37303 343 37337
rect 377 37303 400 37337
rect 320 37017 400 37303
rect 320 36983 343 37017
rect 377 36983 400 37017
rect 320 36960 400 36983
rect 480 37337 560 37360
rect 480 37303 503 37337
rect 537 37303 560 37337
rect 480 37017 560 37303
rect 480 36983 503 37017
rect 537 36983 560 37017
rect 480 36960 560 36983
rect 640 37337 720 37360
rect 640 37303 663 37337
rect 697 37303 720 37337
rect 640 37017 720 37303
rect 640 36983 663 37017
rect 697 36983 720 37017
rect 640 36960 720 36983
rect 800 37337 880 37360
rect 800 37303 823 37337
rect 857 37303 880 37337
rect 800 37017 880 37303
rect 800 36983 823 37017
rect 857 36983 880 37017
rect 800 36960 880 36983
rect 960 37337 1040 37360
rect 960 37303 983 37337
rect 1017 37303 1040 37337
rect 960 37017 1040 37303
rect 960 36983 983 37017
rect 1017 36983 1040 37017
rect 960 36960 1040 36983
rect 1120 37337 1200 37360
rect 1120 37303 1143 37337
rect 1177 37303 1200 37337
rect 1120 37017 1200 37303
rect 1120 36983 1143 37017
rect 1177 36983 1200 37017
rect 1120 36960 1200 36983
rect 1280 37337 1360 37360
rect 1280 37303 1303 37337
rect 1337 37303 1360 37337
rect 1280 37017 1360 37303
rect 1280 36983 1303 37017
rect 1337 36983 1360 37017
rect 1280 36960 1360 36983
rect 1440 37337 1520 37360
rect 1440 37303 1463 37337
rect 1497 37303 1520 37337
rect 1440 37017 1520 37303
rect 1440 36983 1463 37017
rect 1497 36983 1520 37017
rect 1440 36960 1520 36983
rect 1600 37337 1680 37360
rect 1600 37303 1623 37337
rect 1657 37303 1680 37337
rect 1600 37017 1680 37303
rect 1600 36983 1623 37017
rect 1657 36983 1680 37017
rect 1600 36960 1680 36983
rect 1760 37337 1840 37360
rect 1760 37303 1783 37337
rect 1817 37303 1840 37337
rect 1760 37017 1840 37303
rect 1760 36983 1783 37017
rect 1817 36983 1840 37017
rect 1760 36960 1840 36983
rect 1920 37337 2000 37360
rect 1920 37303 1943 37337
rect 1977 37303 2000 37337
rect 1920 37017 2000 37303
rect 1920 36983 1943 37017
rect 1977 36983 2000 37017
rect 1920 36960 2000 36983
rect 2080 37337 2160 37360
rect 2080 37303 2103 37337
rect 2137 37303 2160 37337
rect 2080 37017 2160 37303
rect 2080 36983 2103 37017
rect 2137 36983 2160 37017
rect 2080 36960 2160 36983
rect 2240 37337 2320 37360
rect 2240 37303 2263 37337
rect 2297 37303 2320 37337
rect 2240 37017 2320 37303
rect 2240 36983 2263 37017
rect 2297 36983 2320 37017
rect 2240 36960 2320 36983
rect 2400 37337 2480 37360
rect 2400 37303 2423 37337
rect 2457 37303 2480 37337
rect 2400 37017 2480 37303
rect 2400 36983 2423 37017
rect 2457 36983 2480 37017
rect 2400 36960 2480 36983
rect 2560 37337 2640 37360
rect 2560 37303 2583 37337
rect 2617 37303 2640 37337
rect 2560 37017 2640 37303
rect 2560 36983 2583 37017
rect 2617 36983 2640 37017
rect 2560 36960 2640 36983
rect 2720 37337 2800 37360
rect 2720 37303 2743 37337
rect 2777 37303 2800 37337
rect 2720 37017 2800 37303
rect 2720 36983 2743 37017
rect 2777 36983 2800 37017
rect 2720 36960 2800 36983
rect 2880 37337 2960 37360
rect 2880 37303 2903 37337
rect 2937 37303 2960 37337
rect 2880 37017 2960 37303
rect 2880 36983 2903 37017
rect 2937 36983 2960 37017
rect 2880 36960 2960 36983
rect 3040 37337 3120 37360
rect 3040 37303 3063 37337
rect 3097 37303 3120 37337
rect 3040 37017 3120 37303
rect 3040 36983 3063 37017
rect 3097 36983 3120 37017
rect 3040 36960 3120 36983
rect 3200 37337 3280 37360
rect 3200 37303 3223 37337
rect 3257 37303 3280 37337
rect 3200 37017 3280 37303
rect 3200 36983 3223 37017
rect 3257 36983 3280 37017
rect 3200 36960 3280 36983
rect 3360 37337 3440 37360
rect 3360 37303 3383 37337
rect 3417 37303 3440 37337
rect 3360 37017 3440 37303
rect 3360 36983 3383 37017
rect 3417 36983 3440 37017
rect 3360 36960 3440 36983
rect 3520 37337 3600 37360
rect 3520 37303 3543 37337
rect 3577 37303 3600 37337
rect 3520 37017 3600 37303
rect 3520 36983 3543 37017
rect 3577 36983 3600 37017
rect 3520 36960 3600 36983
rect 3680 37337 3760 37360
rect 3680 37303 3703 37337
rect 3737 37303 3760 37337
rect 3680 37017 3760 37303
rect 3680 36983 3703 37017
rect 3737 36983 3760 37017
rect 3680 36960 3760 36983
rect 3840 37337 3920 37360
rect 3840 37303 3863 37337
rect 3897 37303 3920 37337
rect 3840 37017 3920 37303
rect 3840 36983 3863 37017
rect 3897 36983 3920 37017
rect 3840 36960 3920 36983
rect 4000 37337 4080 37360
rect 4000 37303 4023 37337
rect 4057 37303 4080 37337
rect 4000 37017 4080 37303
rect 4000 36983 4023 37017
rect 4057 36983 4080 37017
rect 4000 36960 4080 36983
rect 4160 37337 4240 37360
rect 4160 37303 4183 37337
rect 4217 37303 4240 37337
rect 4160 37017 4240 37303
rect 4160 36983 4183 37017
rect 4217 36983 4240 37017
rect 4160 36960 4240 36983
rect 4320 37337 4400 37360
rect 4320 37303 4343 37337
rect 4377 37303 4400 37337
rect 4320 37017 4400 37303
rect 4320 36983 4343 37017
rect 4377 36983 4400 37017
rect 4320 36960 4400 36983
rect 4480 37337 4560 37360
rect 4480 37303 4503 37337
rect 4537 37303 4560 37337
rect 4480 37017 4560 37303
rect 4480 36983 4503 37017
rect 4537 36983 4560 37017
rect 4480 36960 4560 36983
rect 4640 37337 4720 37360
rect 4640 37303 4663 37337
rect 4697 37303 4720 37337
rect 4640 37017 4720 37303
rect 4640 36983 4663 37017
rect 4697 36983 4720 37017
rect 4640 36960 4720 36983
rect 4800 37337 4880 37360
rect 4800 37303 4823 37337
rect 4857 37303 4880 37337
rect 4800 37017 4880 37303
rect 4800 36983 4823 37017
rect 4857 36983 4880 37017
rect 4800 36960 4880 36983
rect 4960 37337 5040 37360
rect 4960 37303 4983 37337
rect 5017 37303 5040 37337
rect 4960 37017 5040 37303
rect 4960 36983 4983 37017
rect 5017 36983 5040 37017
rect 4960 36960 5040 36983
rect 5120 37337 5200 37360
rect 5120 37303 5143 37337
rect 5177 37303 5200 37337
rect 5120 37017 5200 37303
rect 5120 36983 5143 37017
rect 5177 36983 5200 37017
rect 5120 36960 5200 36983
rect 5280 37337 5360 37360
rect 5280 37303 5303 37337
rect 5337 37303 5360 37337
rect 5280 37017 5360 37303
rect 5280 36983 5303 37017
rect 5337 36983 5360 37017
rect 5280 36960 5360 36983
rect 5440 37337 5520 37360
rect 5440 37303 5463 37337
rect 5497 37303 5520 37337
rect 5440 37017 5520 37303
rect 5440 36983 5463 37017
rect 5497 36983 5520 37017
rect 5440 36960 5520 36983
rect 5600 37337 5680 37360
rect 5600 37303 5623 37337
rect 5657 37303 5680 37337
rect 5600 37017 5680 37303
rect 5600 36983 5623 37017
rect 5657 36983 5680 37017
rect 5600 36960 5680 36983
rect 5760 37337 5840 37360
rect 5760 37303 5783 37337
rect 5817 37303 5840 37337
rect 5760 37017 5840 37303
rect 5760 36983 5783 37017
rect 5817 36983 5840 37017
rect 5760 36960 5840 36983
rect 5920 37337 6000 37360
rect 5920 37303 5943 37337
rect 5977 37303 6000 37337
rect 5920 37017 6000 37303
rect 5920 36983 5943 37017
rect 5977 36983 6000 37017
rect 5920 36960 6000 36983
rect 6080 37337 6160 37360
rect 6080 37303 6103 37337
rect 6137 37303 6160 37337
rect 6080 37017 6160 37303
rect 6080 36983 6103 37017
rect 6137 36983 6160 37017
rect 6080 36960 6160 36983
rect 6240 37337 6320 37360
rect 6240 37303 6263 37337
rect 6297 37303 6320 37337
rect 6240 37017 6320 37303
rect 6240 36983 6263 37017
rect 6297 36983 6320 37017
rect 6240 36960 6320 36983
rect 6400 37337 6480 37360
rect 6400 37303 6423 37337
rect 6457 37303 6480 37337
rect 6400 37017 6480 37303
rect 6400 36983 6423 37017
rect 6457 36983 6480 37017
rect 6400 36960 6480 36983
rect 6560 37337 6640 37360
rect 6560 37303 6583 37337
rect 6617 37303 6640 37337
rect 6560 37017 6640 37303
rect 6560 36983 6583 37017
rect 6617 36983 6640 37017
rect 6560 36960 6640 36983
rect 6720 37337 6800 37360
rect 6720 37303 6743 37337
rect 6777 37303 6800 37337
rect 6720 37017 6800 37303
rect 6720 36983 6743 37017
rect 6777 36983 6800 37017
rect 6720 36960 6800 36983
rect 6880 37337 6960 37360
rect 6880 37303 6903 37337
rect 6937 37303 6960 37337
rect 6880 37017 6960 37303
rect 6880 36983 6903 37017
rect 6937 36983 6960 37017
rect 6880 36960 6960 36983
rect 7040 37337 7120 37360
rect 7040 37303 7063 37337
rect 7097 37303 7120 37337
rect 7040 37017 7120 37303
rect 7040 36983 7063 37017
rect 7097 36983 7120 37017
rect 7040 36960 7120 36983
rect 7200 37337 7280 37360
rect 7200 37303 7223 37337
rect 7257 37303 7280 37337
rect 7200 37017 7280 37303
rect 7200 36983 7223 37017
rect 7257 36983 7280 37017
rect 7200 36960 7280 36983
rect 7360 37337 7440 37360
rect 7360 37303 7383 37337
rect 7417 37303 7440 37337
rect 7360 37017 7440 37303
rect 7360 36983 7383 37017
rect 7417 36983 7440 37017
rect 7360 36960 7440 36983
rect 7520 37337 7600 37360
rect 7520 37303 7543 37337
rect 7577 37303 7600 37337
rect 7520 37017 7600 37303
rect 7520 36983 7543 37017
rect 7577 36983 7600 37017
rect 7520 36960 7600 36983
rect 7680 37337 7760 37360
rect 7680 37303 7703 37337
rect 7737 37303 7760 37337
rect 7680 37017 7760 37303
rect 7680 36983 7703 37017
rect 7737 36983 7760 37017
rect 7680 36960 7760 36983
rect 7840 37337 7920 37360
rect 7840 37303 7863 37337
rect 7897 37303 7920 37337
rect 7840 37017 7920 37303
rect 7840 36983 7863 37017
rect 7897 36983 7920 37017
rect 7840 36960 7920 36983
rect 8000 37337 8080 37360
rect 8000 37303 8023 37337
rect 8057 37303 8080 37337
rect 8000 37017 8080 37303
rect 8000 36983 8023 37017
rect 8057 36983 8080 37017
rect 8000 36960 8080 36983
rect 8160 37337 8240 37360
rect 8160 37303 8183 37337
rect 8217 37303 8240 37337
rect 8160 37017 8240 37303
rect 8160 36983 8183 37017
rect 8217 36983 8240 37017
rect 8160 36960 8240 36983
rect 8320 37337 8400 37360
rect 8320 37303 8343 37337
rect 8377 37303 8400 37337
rect 8320 37017 8400 37303
rect 8320 36983 8343 37017
rect 8377 36983 8400 37017
rect 8320 36960 8400 36983
rect 8480 36960 8560 37360
rect 8640 36960 8720 37360
rect 8800 36960 8880 37360
rect 8960 36960 9040 37360
rect 9120 36960 9200 37360
rect 9280 36960 9360 37360
rect 9440 36960 9520 37360
rect 9600 36960 9680 37360
rect 9760 36960 9840 37360
rect 9920 36960 10000 37360
rect 10080 36960 10160 37360
rect 10240 36960 10320 37360
rect 10400 36960 10480 37360
rect 10560 36960 10640 37360
rect 10720 36960 10800 37360
rect 10880 36960 10960 37360
rect 11040 36960 11120 37360
rect 11200 36960 11280 37360
rect 11360 36960 11440 37360
rect 11520 36960 11600 37360
rect 11680 36960 11760 37360
rect 11840 36960 11920 37360
rect 12000 36960 12080 37360
rect 12160 36960 12240 37360
rect 12320 36960 12400 37360
rect 12480 37337 12560 37360
rect 12480 37303 12503 37337
rect 12537 37303 12560 37337
rect 12480 37017 12560 37303
rect 12480 36983 12503 37017
rect 12537 36983 12560 37017
rect 12480 36960 12560 36983
rect 12640 37337 12720 37360
rect 12640 37303 12663 37337
rect 12697 37303 12720 37337
rect 12640 37017 12720 37303
rect 12640 36983 12663 37017
rect 12697 36983 12720 37017
rect 12640 36960 12720 36983
rect 12800 37337 12880 37360
rect 12800 37303 12823 37337
rect 12857 37303 12880 37337
rect 12800 37017 12880 37303
rect 12800 36983 12823 37017
rect 12857 36983 12880 37017
rect 12800 36960 12880 36983
rect 12960 37337 13040 37360
rect 12960 37303 12983 37337
rect 13017 37303 13040 37337
rect 12960 37017 13040 37303
rect 12960 36983 12983 37017
rect 13017 36983 13040 37017
rect 12960 36960 13040 36983
rect 13120 37337 13200 37360
rect 13120 37303 13143 37337
rect 13177 37303 13200 37337
rect 13120 37017 13200 37303
rect 13120 36983 13143 37017
rect 13177 36983 13200 37017
rect 13120 36960 13200 36983
rect 13280 37337 13360 37360
rect 13280 37303 13303 37337
rect 13337 37303 13360 37337
rect 13280 37017 13360 37303
rect 13280 36983 13303 37017
rect 13337 36983 13360 37017
rect 13280 36960 13360 36983
rect 13440 37337 13520 37360
rect 13440 37303 13463 37337
rect 13497 37303 13520 37337
rect 13440 37017 13520 37303
rect 13440 36983 13463 37017
rect 13497 36983 13520 37017
rect 13440 36960 13520 36983
rect 13600 37337 13680 37360
rect 13600 37303 13623 37337
rect 13657 37303 13680 37337
rect 13600 37017 13680 37303
rect 13600 36983 13623 37017
rect 13657 36983 13680 37017
rect 13600 36960 13680 36983
rect 13760 37337 13840 37360
rect 13760 37303 13783 37337
rect 13817 37303 13840 37337
rect 13760 37017 13840 37303
rect 13760 36983 13783 37017
rect 13817 36983 13840 37017
rect 13760 36960 13840 36983
rect 13920 37337 14000 37360
rect 13920 37303 13943 37337
rect 13977 37303 14000 37337
rect 13920 37017 14000 37303
rect 13920 36983 13943 37017
rect 13977 36983 14000 37017
rect 13920 36960 14000 36983
rect 14080 37337 14160 37360
rect 14080 37303 14103 37337
rect 14137 37303 14160 37337
rect 14080 37017 14160 37303
rect 14080 36983 14103 37017
rect 14137 36983 14160 37017
rect 14080 36960 14160 36983
rect 14240 37337 14320 37360
rect 14240 37303 14263 37337
rect 14297 37303 14320 37337
rect 14240 37017 14320 37303
rect 14240 36983 14263 37017
rect 14297 36983 14320 37017
rect 14240 36960 14320 36983
rect 14400 37337 14480 37360
rect 14400 37303 14423 37337
rect 14457 37303 14480 37337
rect 14400 37017 14480 37303
rect 14400 36983 14423 37017
rect 14457 36983 14480 37017
rect 14400 36960 14480 36983
rect 14560 37337 14640 37360
rect 14560 37303 14583 37337
rect 14617 37303 14640 37337
rect 14560 37017 14640 37303
rect 14560 36983 14583 37017
rect 14617 36983 14640 37017
rect 14560 36960 14640 36983
rect 14720 37337 14800 37360
rect 14720 37303 14743 37337
rect 14777 37303 14800 37337
rect 14720 37017 14800 37303
rect 14720 36983 14743 37017
rect 14777 36983 14800 37017
rect 14720 36960 14800 36983
rect 14880 37337 14960 37360
rect 14880 37303 14903 37337
rect 14937 37303 14960 37337
rect 14880 37017 14960 37303
rect 14880 36983 14903 37017
rect 14937 36983 14960 37017
rect 14880 36960 14960 36983
rect 15040 37337 15120 37360
rect 15040 37303 15063 37337
rect 15097 37303 15120 37337
rect 15040 37017 15120 37303
rect 15040 36983 15063 37017
rect 15097 36983 15120 37017
rect 15040 36960 15120 36983
rect 15200 37337 15280 37360
rect 15200 37303 15223 37337
rect 15257 37303 15280 37337
rect 15200 37017 15280 37303
rect 15200 36983 15223 37017
rect 15257 36983 15280 37017
rect 15200 36960 15280 36983
rect 15360 37337 15440 37360
rect 15360 37303 15383 37337
rect 15417 37303 15440 37337
rect 15360 37017 15440 37303
rect 15360 36983 15383 37017
rect 15417 36983 15440 37017
rect 15360 36960 15440 36983
rect 15520 37337 15600 37360
rect 15520 37303 15543 37337
rect 15577 37303 15600 37337
rect 15520 37017 15600 37303
rect 15520 36983 15543 37017
rect 15577 36983 15600 37017
rect 15520 36960 15600 36983
rect 15680 37337 15760 37360
rect 15680 37303 15703 37337
rect 15737 37303 15760 37337
rect 15680 37017 15760 37303
rect 15680 36983 15703 37017
rect 15737 36983 15760 37017
rect 15680 36960 15760 36983
rect 15840 37337 15920 37360
rect 15840 37303 15863 37337
rect 15897 37303 15920 37337
rect 15840 37017 15920 37303
rect 15840 36983 15863 37017
rect 15897 36983 15920 37017
rect 15840 36960 15920 36983
rect 16000 37337 16080 37360
rect 16000 37303 16023 37337
rect 16057 37303 16080 37337
rect 16000 37017 16080 37303
rect 16000 36983 16023 37017
rect 16057 36983 16080 37017
rect 16000 36960 16080 36983
rect 16160 37337 16240 37360
rect 16160 37303 16183 37337
rect 16217 37303 16240 37337
rect 16160 37017 16240 37303
rect 16160 36983 16183 37017
rect 16217 36983 16240 37017
rect 16160 36960 16240 36983
rect 16320 37337 16400 37360
rect 16320 37303 16343 37337
rect 16377 37303 16400 37337
rect 16320 37017 16400 37303
rect 16320 36983 16343 37017
rect 16377 36983 16400 37017
rect 16320 36960 16400 36983
rect 16480 37337 16560 37360
rect 16480 37303 16503 37337
rect 16537 37303 16560 37337
rect 16480 37017 16560 37303
rect 16480 36983 16503 37017
rect 16537 36983 16560 37017
rect 16480 36960 16560 36983
rect 16640 37337 16720 37360
rect 16640 37303 16663 37337
rect 16697 37303 16720 37337
rect 16640 37017 16720 37303
rect 16640 36983 16663 37017
rect 16697 36983 16720 37017
rect 16640 36960 16720 36983
rect 16800 37337 16880 37360
rect 16800 37303 16823 37337
rect 16857 37303 16880 37337
rect 16800 37017 16880 37303
rect 16800 36983 16823 37017
rect 16857 36983 16880 37017
rect 16800 36960 16880 36983
rect 16960 37337 17040 37360
rect 16960 37303 16983 37337
rect 17017 37303 17040 37337
rect 16960 37017 17040 37303
rect 16960 36983 16983 37017
rect 17017 36983 17040 37017
rect 16960 36960 17040 36983
rect 17120 37337 17200 37360
rect 17120 37303 17143 37337
rect 17177 37303 17200 37337
rect 17120 37017 17200 37303
rect 17120 36983 17143 37017
rect 17177 36983 17200 37017
rect 17120 36960 17200 36983
rect 17280 37337 17360 37360
rect 17280 37303 17303 37337
rect 17337 37303 17360 37337
rect 17280 37017 17360 37303
rect 17280 36983 17303 37017
rect 17337 36983 17360 37017
rect 17280 36960 17360 36983
rect 17440 37337 17520 37360
rect 17440 37303 17463 37337
rect 17497 37303 17520 37337
rect 17440 37017 17520 37303
rect 17440 36983 17463 37017
rect 17497 36983 17520 37017
rect 17440 36960 17520 36983
rect 17600 37337 17680 37360
rect 17600 37303 17623 37337
rect 17657 37303 17680 37337
rect 17600 37017 17680 37303
rect 17600 36983 17623 37017
rect 17657 36983 17680 37017
rect 17600 36960 17680 36983
rect 17760 37337 17840 37360
rect 17760 37303 17783 37337
rect 17817 37303 17840 37337
rect 17760 37017 17840 37303
rect 17760 36983 17783 37017
rect 17817 36983 17840 37017
rect 17760 36960 17840 36983
rect 17920 37337 18000 37360
rect 17920 37303 17943 37337
rect 17977 37303 18000 37337
rect 17920 37017 18000 37303
rect 17920 36983 17943 37017
rect 17977 36983 18000 37017
rect 17920 36960 18000 36983
rect 18080 37337 18160 37360
rect 18080 37303 18103 37337
rect 18137 37303 18160 37337
rect 18080 37017 18160 37303
rect 18080 36983 18103 37017
rect 18137 36983 18160 37017
rect 18080 36960 18160 36983
rect 18240 37337 18320 37360
rect 18240 37303 18263 37337
rect 18297 37303 18320 37337
rect 18240 37017 18320 37303
rect 18240 36983 18263 37017
rect 18297 36983 18320 37017
rect 18240 36960 18320 36983
rect 18400 37337 18480 37360
rect 18400 37303 18423 37337
rect 18457 37303 18480 37337
rect 18400 37017 18480 37303
rect 18400 36983 18423 37017
rect 18457 36983 18480 37017
rect 18400 36960 18480 36983
rect 18560 37337 18640 37360
rect 18560 37303 18583 37337
rect 18617 37303 18640 37337
rect 18560 37017 18640 37303
rect 18560 36983 18583 37017
rect 18617 36983 18640 37017
rect 18560 36960 18640 36983
rect 18720 37337 18800 37360
rect 18720 37303 18743 37337
rect 18777 37303 18800 37337
rect 18720 37017 18800 37303
rect 18720 36983 18743 37017
rect 18777 36983 18800 37017
rect 18720 36960 18800 36983
rect 18880 37337 18960 37360
rect 18880 37303 18903 37337
rect 18937 37303 18960 37337
rect 18880 37017 18960 37303
rect 18880 36983 18903 37017
rect 18937 36983 18960 37017
rect 18880 36960 18960 36983
rect 19040 36960 19120 37360
rect 19200 36960 19280 37360
rect 19360 36960 19440 37360
rect 19520 36960 19600 37360
rect 19680 36960 19760 37360
rect 19840 36960 19920 37360
rect 20000 36960 20080 37360
rect 20160 36960 20240 37360
rect 20320 36960 20400 37360
rect 20480 36960 20560 37360
rect 20640 36960 20720 37360
rect 20800 36960 20880 37360
rect 20960 36960 21040 37360
rect 21120 36960 21200 37360
rect 21280 36960 21360 37360
rect 21440 36960 21520 37360
rect 21600 36960 21680 37360
rect 21760 36960 21840 37360
rect 21920 36960 22000 37360
rect 22080 36960 22160 37360
rect 22240 36960 22320 37360
rect 22400 36960 22480 37360
rect 22560 36960 22640 37360
rect 22720 36960 22800 37360
rect 22880 36960 22960 37360
rect 23120 37337 23200 37360
rect 23120 37303 23143 37337
rect 23177 37303 23200 37337
rect 23120 37017 23200 37303
rect 23120 36983 23143 37017
rect 23177 36983 23200 37017
rect 23120 36960 23200 36983
rect 23280 37337 23360 37360
rect 23280 37303 23303 37337
rect 23337 37303 23360 37337
rect 23280 37017 23360 37303
rect 23280 36983 23303 37017
rect 23337 36983 23360 37017
rect 23280 36960 23360 36983
rect 23440 37337 23520 37360
rect 23440 37303 23463 37337
rect 23497 37303 23520 37337
rect 23440 37017 23520 37303
rect 23440 36983 23463 37017
rect 23497 36983 23520 37017
rect 23440 36960 23520 36983
rect 23600 37337 23680 37360
rect 23600 37303 23623 37337
rect 23657 37303 23680 37337
rect 23600 37017 23680 37303
rect 23600 36983 23623 37017
rect 23657 36983 23680 37017
rect 23600 36960 23680 36983
rect 23760 37337 23840 37360
rect 23760 37303 23783 37337
rect 23817 37303 23840 37337
rect 23760 37017 23840 37303
rect 23760 36983 23783 37017
rect 23817 36983 23840 37017
rect 23760 36960 23840 36983
rect 23920 37337 24000 37360
rect 23920 37303 23943 37337
rect 23977 37303 24000 37337
rect 23920 37017 24000 37303
rect 23920 36983 23943 37017
rect 23977 36983 24000 37017
rect 23920 36960 24000 36983
rect 24080 37337 24160 37360
rect 24080 37303 24103 37337
rect 24137 37303 24160 37337
rect 24080 37017 24160 37303
rect 24080 36983 24103 37017
rect 24137 36983 24160 37017
rect 24080 36960 24160 36983
rect 24240 37337 24320 37360
rect 24240 37303 24263 37337
rect 24297 37303 24320 37337
rect 24240 37017 24320 37303
rect 24240 36983 24263 37017
rect 24297 36983 24320 37017
rect 24240 36960 24320 36983
rect 24400 37337 24480 37360
rect 24400 37303 24423 37337
rect 24457 37303 24480 37337
rect 24400 37017 24480 37303
rect 24400 36983 24423 37017
rect 24457 36983 24480 37017
rect 24400 36960 24480 36983
rect 24560 37337 24640 37360
rect 24560 37303 24583 37337
rect 24617 37303 24640 37337
rect 24560 37017 24640 37303
rect 24560 36983 24583 37017
rect 24617 36983 24640 37017
rect 24560 36960 24640 36983
rect 24720 37337 24800 37360
rect 24720 37303 24743 37337
rect 24777 37303 24800 37337
rect 24720 37017 24800 37303
rect 24720 36983 24743 37017
rect 24777 36983 24800 37017
rect 24720 36960 24800 36983
rect 24880 37337 24960 37360
rect 24880 37303 24903 37337
rect 24937 37303 24960 37337
rect 24880 37017 24960 37303
rect 24880 36983 24903 37017
rect 24937 36983 24960 37017
rect 24880 36960 24960 36983
rect 25040 37337 25120 37360
rect 25040 37303 25063 37337
rect 25097 37303 25120 37337
rect 25040 37017 25120 37303
rect 25040 36983 25063 37017
rect 25097 36983 25120 37017
rect 25040 36960 25120 36983
rect 25200 37337 25280 37360
rect 25200 37303 25223 37337
rect 25257 37303 25280 37337
rect 25200 37017 25280 37303
rect 25200 36983 25223 37017
rect 25257 36983 25280 37017
rect 25200 36960 25280 36983
rect 25360 37337 25440 37360
rect 25360 37303 25383 37337
rect 25417 37303 25440 37337
rect 25360 37017 25440 37303
rect 25360 36983 25383 37017
rect 25417 36983 25440 37017
rect 25360 36960 25440 36983
rect 25520 37337 25600 37360
rect 25520 37303 25543 37337
rect 25577 37303 25600 37337
rect 25520 37017 25600 37303
rect 25520 36983 25543 37017
rect 25577 36983 25600 37017
rect 25520 36960 25600 36983
rect 25680 37337 25760 37360
rect 25680 37303 25703 37337
rect 25737 37303 25760 37337
rect 25680 37017 25760 37303
rect 25680 36983 25703 37017
rect 25737 36983 25760 37017
rect 25680 36960 25760 36983
rect 25840 37337 25920 37360
rect 25840 37303 25863 37337
rect 25897 37303 25920 37337
rect 25840 37017 25920 37303
rect 25840 36983 25863 37017
rect 25897 36983 25920 37017
rect 25840 36960 25920 36983
rect 26000 37337 26080 37360
rect 26000 37303 26023 37337
rect 26057 37303 26080 37337
rect 26000 37017 26080 37303
rect 26000 36983 26023 37017
rect 26057 36983 26080 37017
rect 26000 36960 26080 36983
rect 26160 37337 26240 37360
rect 26160 37303 26183 37337
rect 26217 37303 26240 37337
rect 26160 37017 26240 37303
rect 26160 36983 26183 37017
rect 26217 36983 26240 37017
rect 26160 36960 26240 36983
rect 26320 37337 26400 37360
rect 26320 37303 26343 37337
rect 26377 37303 26400 37337
rect 26320 37017 26400 37303
rect 26320 36983 26343 37017
rect 26377 36983 26400 37017
rect 26320 36960 26400 36983
rect 26480 37337 26560 37360
rect 26480 37303 26503 37337
rect 26537 37303 26560 37337
rect 26480 37017 26560 37303
rect 26480 36983 26503 37017
rect 26537 36983 26560 37017
rect 26480 36960 26560 36983
rect 26640 37337 26720 37360
rect 26640 37303 26663 37337
rect 26697 37303 26720 37337
rect 26640 37017 26720 37303
rect 26640 36983 26663 37017
rect 26697 36983 26720 37017
rect 26640 36960 26720 36983
rect 26800 37337 26880 37360
rect 26800 37303 26823 37337
rect 26857 37303 26880 37337
rect 26800 37017 26880 37303
rect 26800 36983 26823 37017
rect 26857 36983 26880 37017
rect 26800 36960 26880 36983
rect 26960 37337 27040 37360
rect 26960 37303 26983 37337
rect 27017 37303 27040 37337
rect 26960 37017 27040 37303
rect 26960 36983 26983 37017
rect 27017 36983 27040 37017
rect 26960 36960 27040 36983
rect 27120 37337 27200 37360
rect 27120 37303 27143 37337
rect 27177 37303 27200 37337
rect 27120 37017 27200 37303
rect 27120 36983 27143 37017
rect 27177 36983 27200 37017
rect 27120 36960 27200 36983
rect 27280 37337 27360 37360
rect 27280 37303 27303 37337
rect 27337 37303 27360 37337
rect 27280 37017 27360 37303
rect 27280 36983 27303 37017
rect 27337 36983 27360 37017
rect 27280 36960 27360 36983
rect 27440 37337 27520 37360
rect 27440 37303 27463 37337
rect 27497 37303 27520 37337
rect 27440 37017 27520 37303
rect 27440 36983 27463 37017
rect 27497 36983 27520 37017
rect 27440 36960 27520 36983
rect 27600 37337 27680 37360
rect 27600 37303 27623 37337
rect 27657 37303 27680 37337
rect 27600 37017 27680 37303
rect 27600 36983 27623 37017
rect 27657 36983 27680 37017
rect 27600 36960 27680 36983
rect 27760 37337 27840 37360
rect 27760 37303 27783 37337
rect 27817 37303 27840 37337
rect 27760 37017 27840 37303
rect 27760 36983 27783 37017
rect 27817 36983 27840 37017
rect 27760 36960 27840 36983
rect 27920 37337 28000 37360
rect 27920 37303 27943 37337
rect 27977 37303 28000 37337
rect 27920 37017 28000 37303
rect 27920 36983 27943 37017
rect 27977 36983 28000 37017
rect 27920 36960 28000 36983
rect 28080 37337 28160 37360
rect 28080 37303 28103 37337
rect 28137 37303 28160 37337
rect 28080 37017 28160 37303
rect 28080 36983 28103 37017
rect 28137 36983 28160 37017
rect 28080 36960 28160 36983
rect 28240 37337 28320 37360
rect 28240 37303 28263 37337
rect 28297 37303 28320 37337
rect 28240 37017 28320 37303
rect 28240 36983 28263 37017
rect 28297 36983 28320 37017
rect 28240 36960 28320 36983
rect 28400 37337 28480 37360
rect 28400 37303 28423 37337
rect 28457 37303 28480 37337
rect 28400 37017 28480 37303
rect 28400 36983 28423 37017
rect 28457 36983 28480 37017
rect 28400 36960 28480 36983
rect 28560 37337 28640 37360
rect 28560 37303 28583 37337
rect 28617 37303 28640 37337
rect 28560 37017 28640 37303
rect 28560 36983 28583 37017
rect 28617 36983 28640 37017
rect 28560 36960 28640 36983
rect 28720 37337 28800 37360
rect 28720 37303 28743 37337
rect 28777 37303 28800 37337
rect 28720 37017 28800 37303
rect 28720 36983 28743 37017
rect 28777 36983 28800 37017
rect 28720 36960 28800 36983
rect 28880 37337 28960 37360
rect 28880 37303 28903 37337
rect 28937 37303 28960 37337
rect 28880 37017 28960 37303
rect 28880 36983 28903 37017
rect 28937 36983 28960 37017
rect 28880 36960 28960 36983
rect 29040 37337 29120 37360
rect 29040 37303 29063 37337
rect 29097 37303 29120 37337
rect 29040 37017 29120 37303
rect 29040 36983 29063 37017
rect 29097 36983 29120 37017
rect 29040 36960 29120 36983
rect 29200 37337 29280 37360
rect 29200 37303 29223 37337
rect 29257 37303 29280 37337
rect 29200 37017 29280 37303
rect 29200 36983 29223 37017
rect 29257 36983 29280 37017
rect 29200 36960 29280 36983
rect 29360 37337 29440 37360
rect 29360 37303 29383 37337
rect 29417 37303 29440 37337
rect 29360 37017 29440 37303
rect 29360 36983 29383 37017
rect 29417 36983 29440 37017
rect 29360 36960 29440 36983
rect 29520 36960 29600 37360
rect 29680 36960 29760 37360
rect 29840 36960 29920 37360
rect 30000 36960 30080 37360
rect 30160 36960 30240 37360
rect 30320 36960 30400 37360
rect 30480 36960 30560 37360
rect 30640 36960 30720 37360
rect 30800 36960 30880 37360
rect 30960 36960 31040 37360
rect 31120 36960 31200 37360
rect 31280 36960 31360 37360
rect 31440 36960 31520 37360
rect 31600 36960 31680 37360
rect 31760 36960 31840 37360
rect 31920 36960 32000 37360
rect 32080 36960 32160 37360
rect 32240 36960 32320 37360
rect 32400 36960 32480 37360
rect 32560 36960 32640 37360
rect 32720 36960 32800 37360
rect 32880 36960 32960 37360
rect 33040 36960 33120 37360
rect 33200 36960 33280 37360
rect 33360 36960 33440 37360
rect 33520 37337 33600 37360
rect 33520 37303 33543 37337
rect 33577 37303 33600 37337
rect 33520 37017 33600 37303
rect 33520 36983 33543 37017
rect 33577 36983 33600 37017
rect 33520 36960 33600 36983
rect 33680 37337 33760 37360
rect 33680 37303 33703 37337
rect 33737 37303 33760 37337
rect 33680 37017 33760 37303
rect 33680 36983 33703 37017
rect 33737 36983 33760 37017
rect 33680 36960 33760 36983
rect 33840 37337 33920 37360
rect 33840 37303 33863 37337
rect 33897 37303 33920 37337
rect 33840 37017 33920 37303
rect 33840 36983 33863 37017
rect 33897 36983 33920 37017
rect 33840 36960 33920 36983
rect 34000 37337 34080 37360
rect 34000 37303 34023 37337
rect 34057 37303 34080 37337
rect 34000 37017 34080 37303
rect 34000 36983 34023 37017
rect 34057 36983 34080 37017
rect 34000 36960 34080 36983
rect 34160 37337 34240 37360
rect 34160 37303 34183 37337
rect 34217 37303 34240 37337
rect 34160 37017 34240 37303
rect 34160 36983 34183 37017
rect 34217 36983 34240 37017
rect 34160 36960 34240 36983
rect 34320 37337 34400 37360
rect 34320 37303 34343 37337
rect 34377 37303 34400 37337
rect 34320 37017 34400 37303
rect 34320 36983 34343 37017
rect 34377 36983 34400 37017
rect 34320 36960 34400 36983
rect 34480 37337 34560 37360
rect 34480 37303 34503 37337
rect 34537 37303 34560 37337
rect 34480 37017 34560 37303
rect 34480 36983 34503 37017
rect 34537 36983 34560 37017
rect 34480 36960 34560 36983
rect 34640 37337 34720 37360
rect 34640 37303 34663 37337
rect 34697 37303 34720 37337
rect 34640 37017 34720 37303
rect 34640 36983 34663 37017
rect 34697 36983 34720 37017
rect 34640 36960 34720 36983
rect 34800 37337 34880 37360
rect 34800 37303 34823 37337
rect 34857 37303 34880 37337
rect 34800 37017 34880 37303
rect 34800 36983 34823 37017
rect 34857 36983 34880 37017
rect 34800 36960 34880 36983
rect 34960 37337 35040 37360
rect 34960 37303 34983 37337
rect 35017 37303 35040 37337
rect 34960 37017 35040 37303
rect 34960 36983 34983 37017
rect 35017 36983 35040 37017
rect 34960 36960 35040 36983
rect 35120 37337 35200 37360
rect 35120 37303 35143 37337
rect 35177 37303 35200 37337
rect 35120 37017 35200 37303
rect 35120 36983 35143 37017
rect 35177 36983 35200 37017
rect 35120 36960 35200 36983
rect 35280 37337 35360 37360
rect 35280 37303 35303 37337
rect 35337 37303 35360 37337
rect 35280 37017 35360 37303
rect 35280 36983 35303 37017
rect 35337 36983 35360 37017
rect 35280 36960 35360 36983
rect 35440 37337 35520 37360
rect 35440 37303 35463 37337
rect 35497 37303 35520 37337
rect 35440 37017 35520 37303
rect 35440 36983 35463 37017
rect 35497 36983 35520 37017
rect 35440 36960 35520 36983
rect 35600 37337 35680 37360
rect 35600 37303 35623 37337
rect 35657 37303 35680 37337
rect 35600 37017 35680 37303
rect 35600 36983 35623 37017
rect 35657 36983 35680 37017
rect 35600 36960 35680 36983
rect 35760 37337 35840 37360
rect 35760 37303 35783 37337
rect 35817 37303 35840 37337
rect 35760 37017 35840 37303
rect 35760 36983 35783 37017
rect 35817 36983 35840 37017
rect 35760 36960 35840 36983
rect 35920 37337 36000 37360
rect 35920 37303 35943 37337
rect 35977 37303 36000 37337
rect 35920 37017 36000 37303
rect 35920 36983 35943 37017
rect 35977 36983 36000 37017
rect 35920 36960 36000 36983
rect 36080 37337 36160 37360
rect 36080 37303 36103 37337
rect 36137 37303 36160 37337
rect 36080 37017 36160 37303
rect 36080 36983 36103 37017
rect 36137 36983 36160 37017
rect 36080 36960 36160 36983
rect 36240 37337 36320 37360
rect 36240 37303 36263 37337
rect 36297 37303 36320 37337
rect 36240 37017 36320 37303
rect 36240 36983 36263 37017
rect 36297 36983 36320 37017
rect 36240 36960 36320 36983
rect 36400 37337 36480 37360
rect 36400 37303 36423 37337
rect 36457 37303 36480 37337
rect 36400 37017 36480 37303
rect 36400 36983 36423 37017
rect 36457 36983 36480 37017
rect 36400 36960 36480 36983
rect 36560 37337 36640 37360
rect 36560 37303 36583 37337
rect 36617 37303 36640 37337
rect 36560 37017 36640 37303
rect 36560 36983 36583 37017
rect 36617 36983 36640 37017
rect 36560 36960 36640 36983
rect 36720 37337 36800 37360
rect 36720 37303 36743 37337
rect 36777 37303 36800 37337
rect 36720 37017 36800 37303
rect 36720 36983 36743 37017
rect 36777 36983 36800 37017
rect 36720 36960 36800 36983
rect 36880 37337 36960 37360
rect 36880 37303 36903 37337
rect 36937 37303 36960 37337
rect 36880 37017 36960 37303
rect 36880 36983 36903 37017
rect 36937 36983 36960 37017
rect 36880 36960 36960 36983
rect 37040 37337 37120 37360
rect 37040 37303 37063 37337
rect 37097 37303 37120 37337
rect 37040 37017 37120 37303
rect 37040 36983 37063 37017
rect 37097 36983 37120 37017
rect 37040 36960 37120 36983
rect 37200 37337 37280 37360
rect 37200 37303 37223 37337
rect 37257 37303 37280 37337
rect 37200 37017 37280 37303
rect 37200 36983 37223 37017
rect 37257 36983 37280 37017
rect 37200 36960 37280 36983
rect 37360 37337 37440 37360
rect 37360 37303 37383 37337
rect 37417 37303 37440 37337
rect 37360 37017 37440 37303
rect 37360 36983 37383 37017
rect 37417 36983 37440 37017
rect 37360 36960 37440 36983
rect 37520 37337 37600 37360
rect 37520 37303 37543 37337
rect 37577 37303 37600 37337
rect 37520 37017 37600 37303
rect 37520 36983 37543 37017
rect 37577 36983 37600 37017
rect 37520 36960 37600 36983
rect 37680 37337 37760 37360
rect 37680 37303 37703 37337
rect 37737 37303 37760 37337
rect 37680 37017 37760 37303
rect 37680 36983 37703 37017
rect 37737 36983 37760 37017
rect 37680 36960 37760 36983
rect 37840 37337 37920 37360
rect 37840 37303 37863 37337
rect 37897 37303 37920 37337
rect 37840 37017 37920 37303
rect 37840 36983 37863 37017
rect 37897 36983 37920 37017
rect 37840 36960 37920 36983
rect 38000 37337 38080 37360
rect 38000 37303 38023 37337
rect 38057 37303 38080 37337
rect 38000 37017 38080 37303
rect 38000 36983 38023 37017
rect 38057 36983 38080 37017
rect 38000 36960 38080 36983
rect 38160 37337 38240 37360
rect 38160 37303 38183 37337
rect 38217 37303 38240 37337
rect 38160 37017 38240 37303
rect 38160 36983 38183 37017
rect 38217 36983 38240 37017
rect 38160 36960 38240 36983
rect 38320 37337 38400 37360
rect 38320 37303 38343 37337
rect 38377 37303 38400 37337
rect 38320 37017 38400 37303
rect 38320 36983 38343 37017
rect 38377 36983 38400 37017
rect 38320 36960 38400 36983
rect 38480 37337 38560 37360
rect 38480 37303 38503 37337
rect 38537 37303 38560 37337
rect 38480 37017 38560 37303
rect 38480 36983 38503 37017
rect 38537 36983 38560 37017
rect 38480 36960 38560 36983
rect 38640 37337 38720 37360
rect 38640 37303 38663 37337
rect 38697 37303 38720 37337
rect 38640 37017 38720 37303
rect 38640 36983 38663 37017
rect 38697 36983 38720 37017
rect 38640 36960 38720 36983
rect 38800 37337 38880 37360
rect 38800 37303 38823 37337
rect 38857 37303 38880 37337
rect 38800 37017 38880 37303
rect 38800 36983 38823 37017
rect 38857 36983 38880 37017
rect 38800 36960 38880 36983
rect 38960 37337 39040 37360
rect 38960 37303 38983 37337
rect 39017 37303 39040 37337
rect 38960 37017 39040 37303
rect 38960 36983 38983 37017
rect 39017 36983 39040 37017
rect 38960 36960 39040 36983
rect 39120 37337 39200 37360
rect 39120 37303 39143 37337
rect 39177 37303 39200 37337
rect 39120 37017 39200 37303
rect 39120 36983 39143 37017
rect 39177 36983 39200 37017
rect 39120 36960 39200 36983
rect 39280 37337 39360 37360
rect 39280 37303 39303 37337
rect 39337 37303 39360 37337
rect 39280 37017 39360 37303
rect 39280 36983 39303 37017
rect 39337 36983 39360 37017
rect 39280 36960 39360 36983
rect 39440 37337 39520 37360
rect 39440 37303 39463 37337
rect 39497 37303 39520 37337
rect 39440 37017 39520 37303
rect 39440 36983 39463 37017
rect 39497 36983 39520 37017
rect 39440 36960 39520 36983
rect 39600 37337 39680 37360
rect 39600 37303 39623 37337
rect 39657 37303 39680 37337
rect 39600 37017 39680 37303
rect 39600 36983 39623 37017
rect 39657 36983 39680 37017
rect 39600 36960 39680 36983
rect 39760 37337 39840 37360
rect 39760 37303 39783 37337
rect 39817 37303 39840 37337
rect 39760 37017 39840 37303
rect 39760 36983 39783 37017
rect 39817 36983 39840 37017
rect 39760 36960 39840 36983
rect 39920 37337 40000 37360
rect 39920 37303 39943 37337
rect 39977 37303 40000 37337
rect 39920 37017 40000 37303
rect 39920 36983 39943 37017
rect 39977 36983 40000 37017
rect 39920 36960 40000 36983
rect 40080 37337 40160 37360
rect 40080 37303 40103 37337
rect 40137 37303 40160 37337
rect 40080 37017 40160 37303
rect 40080 36983 40103 37017
rect 40137 36983 40160 37017
rect 40080 36960 40160 36983
rect 40240 37337 40320 37360
rect 40240 37303 40263 37337
rect 40297 37303 40320 37337
rect 40240 37017 40320 37303
rect 40240 36983 40263 37017
rect 40297 36983 40320 37017
rect 40240 36960 40320 36983
rect 40400 37337 40480 37360
rect 40400 37303 40423 37337
rect 40457 37303 40480 37337
rect 40400 37017 40480 37303
rect 40400 36983 40423 37017
rect 40457 36983 40480 37017
rect 40400 36960 40480 36983
rect 40560 37337 40640 37360
rect 40560 37303 40583 37337
rect 40617 37303 40640 37337
rect 40560 37017 40640 37303
rect 40560 36983 40583 37017
rect 40617 36983 40640 37017
rect 40560 36960 40640 36983
rect 40720 37337 40800 37360
rect 40720 37303 40743 37337
rect 40777 37303 40800 37337
rect 40720 37017 40800 37303
rect 40720 36983 40743 37017
rect 40777 36983 40800 37017
rect 40720 36960 40800 36983
rect 40880 37337 40960 37360
rect 40880 37303 40903 37337
rect 40937 37303 40960 37337
rect 40880 37017 40960 37303
rect 40880 36983 40903 37017
rect 40937 36983 40960 37017
rect 40880 36960 40960 36983
rect 41040 37337 41120 37360
rect 41040 37303 41063 37337
rect 41097 37303 41120 37337
rect 41040 37017 41120 37303
rect 41040 36983 41063 37017
rect 41097 36983 41120 37017
rect 41040 36960 41120 36983
rect 41200 37337 41280 37360
rect 41200 37303 41223 37337
rect 41257 37303 41280 37337
rect 41200 37017 41280 37303
rect 41200 36983 41223 37017
rect 41257 36983 41280 37017
rect 41200 36960 41280 36983
rect 41360 37337 41440 37360
rect 41360 37303 41383 37337
rect 41417 37303 41440 37337
rect 41360 37017 41440 37303
rect 41360 36983 41383 37017
rect 41417 36983 41440 37017
rect 41360 36960 41440 36983
rect 41520 37337 41600 37360
rect 41520 37303 41543 37337
rect 41577 37303 41600 37337
rect 41520 37017 41600 37303
rect 41520 36983 41543 37017
rect 41577 36983 41600 37017
rect 41520 36960 41600 36983
rect 41680 37337 41760 37360
rect 41680 37303 41703 37337
rect 41737 37303 41760 37337
rect 41680 37017 41760 37303
rect 41680 36983 41703 37017
rect 41737 36983 41760 37017
rect 41680 36960 41760 36983
rect 41840 37337 41920 37360
rect 41840 37303 41863 37337
rect 41897 37303 41920 37337
rect 41840 37017 41920 37303
rect 41840 36983 41863 37017
rect 41897 36983 41920 37017
rect 41840 36960 41920 36983
rect 0 36857 80 36880
rect 0 36823 23 36857
rect 57 36823 80 36857
rect 0 36537 80 36823
rect 0 36503 23 36537
rect 57 36503 80 36537
rect 0 36480 80 36503
rect 160 36857 240 36880
rect 160 36823 183 36857
rect 217 36823 240 36857
rect 160 36537 240 36823
rect 160 36503 183 36537
rect 217 36503 240 36537
rect 160 36480 240 36503
rect 320 36857 400 36880
rect 320 36823 343 36857
rect 377 36823 400 36857
rect 320 36537 400 36823
rect 320 36503 343 36537
rect 377 36503 400 36537
rect 320 36480 400 36503
rect 480 36857 560 36880
rect 480 36823 503 36857
rect 537 36823 560 36857
rect 480 36537 560 36823
rect 480 36503 503 36537
rect 537 36503 560 36537
rect 480 36480 560 36503
rect 640 36857 720 36880
rect 640 36823 663 36857
rect 697 36823 720 36857
rect 640 36537 720 36823
rect 640 36503 663 36537
rect 697 36503 720 36537
rect 640 36480 720 36503
rect 800 36857 880 36880
rect 800 36823 823 36857
rect 857 36823 880 36857
rect 800 36537 880 36823
rect 800 36503 823 36537
rect 857 36503 880 36537
rect 800 36480 880 36503
rect 960 36857 1040 36880
rect 960 36823 983 36857
rect 1017 36823 1040 36857
rect 960 36537 1040 36823
rect 960 36503 983 36537
rect 1017 36503 1040 36537
rect 960 36480 1040 36503
rect 1120 36857 1200 36880
rect 1120 36823 1143 36857
rect 1177 36823 1200 36857
rect 1120 36537 1200 36823
rect 1120 36503 1143 36537
rect 1177 36503 1200 36537
rect 1120 36480 1200 36503
rect 1280 36857 1360 36880
rect 1280 36823 1303 36857
rect 1337 36823 1360 36857
rect 1280 36537 1360 36823
rect 1280 36503 1303 36537
rect 1337 36503 1360 36537
rect 1280 36480 1360 36503
rect 1440 36857 1520 36880
rect 1440 36823 1463 36857
rect 1497 36823 1520 36857
rect 1440 36537 1520 36823
rect 1440 36503 1463 36537
rect 1497 36503 1520 36537
rect 1440 36480 1520 36503
rect 1600 36857 1680 36880
rect 1600 36823 1623 36857
rect 1657 36823 1680 36857
rect 1600 36537 1680 36823
rect 1600 36503 1623 36537
rect 1657 36503 1680 36537
rect 1600 36480 1680 36503
rect 1760 36857 1840 36880
rect 1760 36823 1783 36857
rect 1817 36823 1840 36857
rect 1760 36537 1840 36823
rect 1760 36503 1783 36537
rect 1817 36503 1840 36537
rect 1760 36480 1840 36503
rect 1920 36857 2000 36880
rect 1920 36823 1943 36857
rect 1977 36823 2000 36857
rect 1920 36537 2000 36823
rect 1920 36503 1943 36537
rect 1977 36503 2000 36537
rect 1920 36480 2000 36503
rect 2080 36857 2160 36880
rect 2080 36823 2103 36857
rect 2137 36823 2160 36857
rect 2080 36537 2160 36823
rect 2080 36503 2103 36537
rect 2137 36503 2160 36537
rect 2080 36480 2160 36503
rect 2240 36857 2320 36880
rect 2240 36823 2263 36857
rect 2297 36823 2320 36857
rect 2240 36537 2320 36823
rect 2240 36503 2263 36537
rect 2297 36503 2320 36537
rect 2240 36480 2320 36503
rect 2400 36857 2480 36880
rect 2400 36823 2423 36857
rect 2457 36823 2480 36857
rect 2400 36537 2480 36823
rect 2400 36503 2423 36537
rect 2457 36503 2480 36537
rect 2400 36480 2480 36503
rect 2560 36857 2640 36880
rect 2560 36823 2583 36857
rect 2617 36823 2640 36857
rect 2560 36537 2640 36823
rect 2560 36503 2583 36537
rect 2617 36503 2640 36537
rect 2560 36480 2640 36503
rect 2720 36857 2800 36880
rect 2720 36823 2743 36857
rect 2777 36823 2800 36857
rect 2720 36537 2800 36823
rect 2720 36503 2743 36537
rect 2777 36503 2800 36537
rect 2720 36480 2800 36503
rect 2880 36857 2960 36880
rect 2880 36823 2903 36857
rect 2937 36823 2960 36857
rect 2880 36537 2960 36823
rect 2880 36503 2903 36537
rect 2937 36503 2960 36537
rect 2880 36480 2960 36503
rect 3040 36857 3120 36880
rect 3040 36823 3063 36857
rect 3097 36823 3120 36857
rect 3040 36537 3120 36823
rect 3040 36503 3063 36537
rect 3097 36503 3120 36537
rect 3040 36480 3120 36503
rect 3200 36857 3280 36880
rect 3200 36823 3223 36857
rect 3257 36823 3280 36857
rect 3200 36537 3280 36823
rect 3200 36503 3223 36537
rect 3257 36503 3280 36537
rect 3200 36480 3280 36503
rect 3360 36857 3440 36880
rect 3360 36823 3383 36857
rect 3417 36823 3440 36857
rect 3360 36537 3440 36823
rect 3360 36503 3383 36537
rect 3417 36503 3440 36537
rect 3360 36480 3440 36503
rect 3520 36857 3600 36880
rect 3520 36823 3543 36857
rect 3577 36823 3600 36857
rect 3520 36537 3600 36823
rect 3520 36503 3543 36537
rect 3577 36503 3600 36537
rect 3520 36480 3600 36503
rect 3680 36857 3760 36880
rect 3680 36823 3703 36857
rect 3737 36823 3760 36857
rect 3680 36537 3760 36823
rect 3680 36503 3703 36537
rect 3737 36503 3760 36537
rect 3680 36480 3760 36503
rect 3840 36857 3920 36880
rect 3840 36823 3863 36857
rect 3897 36823 3920 36857
rect 3840 36537 3920 36823
rect 3840 36503 3863 36537
rect 3897 36503 3920 36537
rect 3840 36480 3920 36503
rect 4000 36857 4080 36880
rect 4000 36823 4023 36857
rect 4057 36823 4080 36857
rect 4000 36537 4080 36823
rect 4000 36503 4023 36537
rect 4057 36503 4080 36537
rect 4000 36480 4080 36503
rect 4160 36857 4240 36880
rect 4160 36823 4183 36857
rect 4217 36823 4240 36857
rect 4160 36537 4240 36823
rect 4160 36503 4183 36537
rect 4217 36503 4240 36537
rect 4160 36480 4240 36503
rect 4320 36857 4400 36880
rect 4320 36823 4343 36857
rect 4377 36823 4400 36857
rect 4320 36537 4400 36823
rect 4320 36503 4343 36537
rect 4377 36503 4400 36537
rect 4320 36480 4400 36503
rect 4480 36857 4560 36880
rect 4480 36823 4503 36857
rect 4537 36823 4560 36857
rect 4480 36537 4560 36823
rect 4480 36503 4503 36537
rect 4537 36503 4560 36537
rect 4480 36480 4560 36503
rect 4640 36857 4720 36880
rect 4640 36823 4663 36857
rect 4697 36823 4720 36857
rect 4640 36537 4720 36823
rect 4640 36503 4663 36537
rect 4697 36503 4720 36537
rect 4640 36480 4720 36503
rect 4800 36857 4880 36880
rect 4800 36823 4823 36857
rect 4857 36823 4880 36857
rect 4800 36537 4880 36823
rect 4800 36503 4823 36537
rect 4857 36503 4880 36537
rect 4800 36480 4880 36503
rect 4960 36857 5040 36880
rect 4960 36823 4983 36857
rect 5017 36823 5040 36857
rect 4960 36537 5040 36823
rect 4960 36503 4983 36537
rect 5017 36503 5040 36537
rect 4960 36480 5040 36503
rect 5120 36857 5200 36880
rect 5120 36823 5143 36857
rect 5177 36823 5200 36857
rect 5120 36537 5200 36823
rect 5120 36503 5143 36537
rect 5177 36503 5200 36537
rect 5120 36480 5200 36503
rect 5280 36857 5360 36880
rect 5280 36823 5303 36857
rect 5337 36823 5360 36857
rect 5280 36537 5360 36823
rect 5280 36503 5303 36537
rect 5337 36503 5360 36537
rect 5280 36480 5360 36503
rect 5440 36857 5520 36880
rect 5440 36823 5463 36857
rect 5497 36823 5520 36857
rect 5440 36537 5520 36823
rect 5440 36503 5463 36537
rect 5497 36503 5520 36537
rect 5440 36480 5520 36503
rect 5600 36857 5680 36880
rect 5600 36823 5623 36857
rect 5657 36823 5680 36857
rect 5600 36537 5680 36823
rect 5600 36503 5623 36537
rect 5657 36503 5680 36537
rect 5600 36480 5680 36503
rect 5760 36857 5840 36880
rect 5760 36823 5783 36857
rect 5817 36823 5840 36857
rect 5760 36537 5840 36823
rect 5760 36503 5783 36537
rect 5817 36503 5840 36537
rect 5760 36480 5840 36503
rect 5920 36857 6000 36880
rect 5920 36823 5943 36857
rect 5977 36823 6000 36857
rect 5920 36537 6000 36823
rect 5920 36503 5943 36537
rect 5977 36503 6000 36537
rect 5920 36480 6000 36503
rect 6080 36857 6160 36880
rect 6080 36823 6103 36857
rect 6137 36823 6160 36857
rect 6080 36537 6160 36823
rect 6080 36503 6103 36537
rect 6137 36503 6160 36537
rect 6080 36480 6160 36503
rect 6240 36857 6320 36880
rect 6240 36823 6263 36857
rect 6297 36823 6320 36857
rect 6240 36537 6320 36823
rect 6240 36503 6263 36537
rect 6297 36503 6320 36537
rect 6240 36480 6320 36503
rect 6400 36857 6480 36880
rect 6400 36823 6423 36857
rect 6457 36823 6480 36857
rect 6400 36537 6480 36823
rect 6400 36503 6423 36537
rect 6457 36503 6480 36537
rect 6400 36480 6480 36503
rect 6560 36857 6640 36880
rect 6560 36823 6583 36857
rect 6617 36823 6640 36857
rect 6560 36537 6640 36823
rect 6560 36503 6583 36537
rect 6617 36503 6640 36537
rect 6560 36480 6640 36503
rect 6720 36857 6800 36880
rect 6720 36823 6743 36857
rect 6777 36823 6800 36857
rect 6720 36537 6800 36823
rect 6720 36503 6743 36537
rect 6777 36503 6800 36537
rect 6720 36480 6800 36503
rect 6880 36857 6960 36880
rect 6880 36823 6903 36857
rect 6937 36823 6960 36857
rect 6880 36537 6960 36823
rect 6880 36503 6903 36537
rect 6937 36503 6960 36537
rect 6880 36480 6960 36503
rect 7040 36857 7120 36880
rect 7040 36823 7063 36857
rect 7097 36823 7120 36857
rect 7040 36537 7120 36823
rect 7040 36503 7063 36537
rect 7097 36503 7120 36537
rect 7040 36480 7120 36503
rect 7200 36857 7280 36880
rect 7200 36823 7223 36857
rect 7257 36823 7280 36857
rect 7200 36537 7280 36823
rect 7200 36503 7223 36537
rect 7257 36503 7280 36537
rect 7200 36480 7280 36503
rect 7360 36857 7440 36880
rect 7360 36823 7383 36857
rect 7417 36823 7440 36857
rect 7360 36537 7440 36823
rect 7360 36503 7383 36537
rect 7417 36503 7440 36537
rect 7360 36480 7440 36503
rect 7520 36857 7600 36880
rect 7520 36823 7543 36857
rect 7577 36823 7600 36857
rect 7520 36537 7600 36823
rect 7520 36503 7543 36537
rect 7577 36503 7600 36537
rect 7520 36480 7600 36503
rect 7680 36857 7760 36880
rect 7680 36823 7703 36857
rect 7737 36823 7760 36857
rect 7680 36537 7760 36823
rect 7680 36503 7703 36537
rect 7737 36503 7760 36537
rect 7680 36480 7760 36503
rect 7840 36857 7920 36880
rect 7840 36823 7863 36857
rect 7897 36823 7920 36857
rect 7840 36537 7920 36823
rect 7840 36503 7863 36537
rect 7897 36503 7920 36537
rect 7840 36480 7920 36503
rect 8000 36857 8080 36880
rect 8000 36823 8023 36857
rect 8057 36823 8080 36857
rect 8000 36537 8080 36823
rect 8000 36503 8023 36537
rect 8057 36503 8080 36537
rect 8000 36480 8080 36503
rect 8160 36857 8240 36880
rect 8160 36823 8183 36857
rect 8217 36823 8240 36857
rect 8160 36537 8240 36823
rect 8160 36503 8183 36537
rect 8217 36503 8240 36537
rect 8160 36480 8240 36503
rect 8320 36857 8400 36880
rect 8320 36823 8343 36857
rect 8377 36823 8400 36857
rect 8320 36537 8400 36823
rect 8320 36503 8343 36537
rect 8377 36503 8400 36537
rect 8320 36480 8400 36503
rect 8480 36480 8560 36880
rect 8640 36480 8720 36880
rect 8800 36480 8880 36880
rect 8960 36480 9040 36880
rect 9120 36480 9200 36880
rect 9280 36480 9360 36880
rect 9440 36480 9520 36880
rect 9600 36480 9680 36880
rect 9760 36480 9840 36880
rect 9920 36480 10000 36880
rect 10080 36480 10160 36880
rect 10240 36480 10320 36880
rect 10400 36480 10480 36880
rect 10560 36480 10640 36880
rect 10720 36480 10800 36880
rect 10880 36480 10960 36880
rect 11040 36480 11120 36880
rect 11200 36480 11280 36880
rect 11360 36480 11440 36880
rect 11520 36480 11600 36880
rect 11680 36480 11760 36880
rect 11840 36480 11920 36880
rect 12000 36480 12080 36880
rect 12160 36480 12240 36880
rect 12320 36480 12400 36880
rect 12480 36857 12560 36880
rect 12480 36823 12503 36857
rect 12537 36823 12560 36857
rect 12480 36537 12560 36823
rect 12480 36503 12503 36537
rect 12537 36503 12560 36537
rect 12480 36480 12560 36503
rect 12640 36857 12720 36880
rect 12640 36823 12663 36857
rect 12697 36823 12720 36857
rect 12640 36537 12720 36823
rect 12640 36503 12663 36537
rect 12697 36503 12720 36537
rect 12640 36480 12720 36503
rect 12800 36857 12880 36880
rect 12800 36823 12823 36857
rect 12857 36823 12880 36857
rect 12800 36537 12880 36823
rect 12800 36503 12823 36537
rect 12857 36503 12880 36537
rect 12800 36480 12880 36503
rect 12960 36857 13040 36880
rect 12960 36823 12983 36857
rect 13017 36823 13040 36857
rect 12960 36537 13040 36823
rect 12960 36503 12983 36537
rect 13017 36503 13040 36537
rect 12960 36480 13040 36503
rect 13120 36857 13200 36880
rect 13120 36823 13143 36857
rect 13177 36823 13200 36857
rect 13120 36537 13200 36823
rect 13120 36503 13143 36537
rect 13177 36503 13200 36537
rect 13120 36480 13200 36503
rect 13280 36857 13360 36880
rect 13280 36823 13303 36857
rect 13337 36823 13360 36857
rect 13280 36537 13360 36823
rect 13280 36503 13303 36537
rect 13337 36503 13360 36537
rect 13280 36480 13360 36503
rect 13440 36857 13520 36880
rect 13440 36823 13463 36857
rect 13497 36823 13520 36857
rect 13440 36537 13520 36823
rect 13440 36503 13463 36537
rect 13497 36503 13520 36537
rect 13440 36480 13520 36503
rect 13600 36857 13680 36880
rect 13600 36823 13623 36857
rect 13657 36823 13680 36857
rect 13600 36537 13680 36823
rect 13600 36503 13623 36537
rect 13657 36503 13680 36537
rect 13600 36480 13680 36503
rect 13760 36857 13840 36880
rect 13760 36823 13783 36857
rect 13817 36823 13840 36857
rect 13760 36537 13840 36823
rect 13760 36503 13783 36537
rect 13817 36503 13840 36537
rect 13760 36480 13840 36503
rect 13920 36857 14000 36880
rect 13920 36823 13943 36857
rect 13977 36823 14000 36857
rect 13920 36537 14000 36823
rect 13920 36503 13943 36537
rect 13977 36503 14000 36537
rect 13920 36480 14000 36503
rect 14080 36857 14160 36880
rect 14080 36823 14103 36857
rect 14137 36823 14160 36857
rect 14080 36537 14160 36823
rect 14080 36503 14103 36537
rect 14137 36503 14160 36537
rect 14080 36480 14160 36503
rect 14240 36857 14320 36880
rect 14240 36823 14263 36857
rect 14297 36823 14320 36857
rect 14240 36537 14320 36823
rect 14240 36503 14263 36537
rect 14297 36503 14320 36537
rect 14240 36480 14320 36503
rect 14400 36857 14480 36880
rect 14400 36823 14423 36857
rect 14457 36823 14480 36857
rect 14400 36537 14480 36823
rect 14400 36503 14423 36537
rect 14457 36503 14480 36537
rect 14400 36480 14480 36503
rect 14560 36857 14640 36880
rect 14560 36823 14583 36857
rect 14617 36823 14640 36857
rect 14560 36537 14640 36823
rect 14560 36503 14583 36537
rect 14617 36503 14640 36537
rect 14560 36480 14640 36503
rect 14720 36857 14800 36880
rect 14720 36823 14743 36857
rect 14777 36823 14800 36857
rect 14720 36537 14800 36823
rect 14720 36503 14743 36537
rect 14777 36503 14800 36537
rect 14720 36480 14800 36503
rect 14880 36857 14960 36880
rect 14880 36823 14903 36857
rect 14937 36823 14960 36857
rect 14880 36537 14960 36823
rect 14880 36503 14903 36537
rect 14937 36503 14960 36537
rect 14880 36480 14960 36503
rect 15040 36857 15120 36880
rect 15040 36823 15063 36857
rect 15097 36823 15120 36857
rect 15040 36537 15120 36823
rect 15040 36503 15063 36537
rect 15097 36503 15120 36537
rect 15040 36480 15120 36503
rect 15200 36857 15280 36880
rect 15200 36823 15223 36857
rect 15257 36823 15280 36857
rect 15200 36537 15280 36823
rect 15200 36503 15223 36537
rect 15257 36503 15280 36537
rect 15200 36480 15280 36503
rect 15360 36857 15440 36880
rect 15360 36823 15383 36857
rect 15417 36823 15440 36857
rect 15360 36537 15440 36823
rect 15360 36503 15383 36537
rect 15417 36503 15440 36537
rect 15360 36480 15440 36503
rect 15520 36857 15600 36880
rect 15520 36823 15543 36857
rect 15577 36823 15600 36857
rect 15520 36537 15600 36823
rect 15520 36503 15543 36537
rect 15577 36503 15600 36537
rect 15520 36480 15600 36503
rect 15680 36857 15760 36880
rect 15680 36823 15703 36857
rect 15737 36823 15760 36857
rect 15680 36537 15760 36823
rect 15680 36503 15703 36537
rect 15737 36503 15760 36537
rect 15680 36480 15760 36503
rect 15840 36857 15920 36880
rect 15840 36823 15863 36857
rect 15897 36823 15920 36857
rect 15840 36537 15920 36823
rect 15840 36503 15863 36537
rect 15897 36503 15920 36537
rect 15840 36480 15920 36503
rect 16000 36857 16080 36880
rect 16000 36823 16023 36857
rect 16057 36823 16080 36857
rect 16000 36537 16080 36823
rect 16000 36503 16023 36537
rect 16057 36503 16080 36537
rect 16000 36480 16080 36503
rect 16160 36857 16240 36880
rect 16160 36823 16183 36857
rect 16217 36823 16240 36857
rect 16160 36537 16240 36823
rect 16160 36503 16183 36537
rect 16217 36503 16240 36537
rect 16160 36480 16240 36503
rect 16320 36857 16400 36880
rect 16320 36823 16343 36857
rect 16377 36823 16400 36857
rect 16320 36537 16400 36823
rect 16320 36503 16343 36537
rect 16377 36503 16400 36537
rect 16320 36480 16400 36503
rect 16480 36857 16560 36880
rect 16480 36823 16503 36857
rect 16537 36823 16560 36857
rect 16480 36537 16560 36823
rect 16480 36503 16503 36537
rect 16537 36503 16560 36537
rect 16480 36480 16560 36503
rect 16640 36857 16720 36880
rect 16640 36823 16663 36857
rect 16697 36823 16720 36857
rect 16640 36537 16720 36823
rect 16640 36503 16663 36537
rect 16697 36503 16720 36537
rect 16640 36480 16720 36503
rect 16800 36857 16880 36880
rect 16800 36823 16823 36857
rect 16857 36823 16880 36857
rect 16800 36537 16880 36823
rect 16800 36503 16823 36537
rect 16857 36503 16880 36537
rect 16800 36480 16880 36503
rect 16960 36857 17040 36880
rect 16960 36823 16983 36857
rect 17017 36823 17040 36857
rect 16960 36537 17040 36823
rect 16960 36503 16983 36537
rect 17017 36503 17040 36537
rect 16960 36480 17040 36503
rect 17120 36857 17200 36880
rect 17120 36823 17143 36857
rect 17177 36823 17200 36857
rect 17120 36537 17200 36823
rect 17120 36503 17143 36537
rect 17177 36503 17200 36537
rect 17120 36480 17200 36503
rect 17280 36857 17360 36880
rect 17280 36823 17303 36857
rect 17337 36823 17360 36857
rect 17280 36537 17360 36823
rect 17280 36503 17303 36537
rect 17337 36503 17360 36537
rect 17280 36480 17360 36503
rect 17440 36857 17520 36880
rect 17440 36823 17463 36857
rect 17497 36823 17520 36857
rect 17440 36537 17520 36823
rect 17440 36503 17463 36537
rect 17497 36503 17520 36537
rect 17440 36480 17520 36503
rect 17600 36857 17680 36880
rect 17600 36823 17623 36857
rect 17657 36823 17680 36857
rect 17600 36537 17680 36823
rect 17600 36503 17623 36537
rect 17657 36503 17680 36537
rect 17600 36480 17680 36503
rect 17760 36857 17840 36880
rect 17760 36823 17783 36857
rect 17817 36823 17840 36857
rect 17760 36537 17840 36823
rect 17760 36503 17783 36537
rect 17817 36503 17840 36537
rect 17760 36480 17840 36503
rect 17920 36857 18000 36880
rect 17920 36823 17943 36857
rect 17977 36823 18000 36857
rect 17920 36537 18000 36823
rect 17920 36503 17943 36537
rect 17977 36503 18000 36537
rect 17920 36480 18000 36503
rect 18080 36857 18160 36880
rect 18080 36823 18103 36857
rect 18137 36823 18160 36857
rect 18080 36537 18160 36823
rect 18080 36503 18103 36537
rect 18137 36503 18160 36537
rect 18080 36480 18160 36503
rect 18240 36857 18320 36880
rect 18240 36823 18263 36857
rect 18297 36823 18320 36857
rect 18240 36537 18320 36823
rect 18240 36503 18263 36537
rect 18297 36503 18320 36537
rect 18240 36480 18320 36503
rect 18400 36857 18480 36880
rect 18400 36823 18423 36857
rect 18457 36823 18480 36857
rect 18400 36537 18480 36823
rect 18400 36503 18423 36537
rect 18457 36503 18480 36537
rect 18400 36480 18480 36503
rect 18560 36857 18640 36880
rect 18560 36823 18583 36857
rect 18617 36823 18640 36857
rect 18560 36537 18640 36823
rect 18560 36503 18583 36537
rect 18617 36503 18640 36537
rect 18560 36480 18640 36503
rect 18720 36857 18800 36880
rect 18720 36823 18743 36857
rect 18777 36823 18800 36857
rect 18720 36537 18800 36823
rect 18720 36503 18743 36537
rect 18777 36503 18800 36537
rect 18720 36480 18800 36503
rect 18880 36857 18960 36880
rect 18880 36823 18903 36857
rect 18937 36823 18960 36857
rect 18880 36537 18960 36823
rect 18880 36503 18903 36537
rect 18937 36503 18960 36537
rect 18880 36480 18960 36503
rect 19040 36480 19120 36880
rect 19200 36480 19280 36880
rect 19360 36480 19440 36880
rect 19520 36480 19600 36880
rect 19680 36480 19760 36880
rect 19840 36480 19920 36880
rect 20000 36480 20080 36880
rect 20160 36480 20240 36880
rect 20320 36480 20400 36880
rect 20480 36480 20560 36880
rect 20640 36480 20720 36880
rect 20800 36480 20880 36880
rect 20960 36480 21040 36880
rect 21120 36480 21200 36880
rect 21280 36480 21360 36880
rect 21440 36480 21520 36880
rect 21600 36480 21680 36880
rect 21760 36480 21840 36880
rect 21920 36480 22000 36880
rect 22080 36480 22160 36880
rect 22240 36480 22320 36880
rect 22400 36480 22480 36880
rect 22560 36480 22640 36880
rect 22720 36480 22800 36880
rect 22880 36480 22960 36880
rect 23120 36857 23200 36880
rect 23120 36823 23143 36857
rect 23177 36823 23200 36857
rect 23120 36537 23200 36823
rect 23120 36503 23143 36537
rect 23177 36503 23200 36537
rect 23120 36480 23200 36503
rect 23280 36857 23360 36880
rect 23280 36823 23303 36857
rect 23337 36823 23360 36857
rect 23280 36537 23360 36823
rect 23280 36503 23303 36537
rect 23337 36503 23360 36537
rect 23280 36480 23360 36503
rect 23440 36857 23520 36880
rect 23440 36823 23463 36857
rect 23497 36823 23520 36857
rect 23440 36537 23520 36823
rect 23440 36503 23463 36537
rect 23497 36503 23520 36537
rect 23440 36480 23520 36503
rect 23600 36857 23680 36880
rect 23600 36823 23623 36857
rect 23657 36823 23680 36857
rect 23600 36537 23680 36823
rect 23600 36503 23623 36537
rect 23657 36503 23680 36537
rect 23600 36480 23680 36503
rect 23760 36857 23840 36880
rect 23760 36823 23783 36857
rect 23817 36823 23840 36857
rect 23760 36537 23840 36823
rect 23760 36503 23783 36537
rect 23817 36503 23840 36537
rect 23760 36480 23840 36503
rect 23920 36857 24000 36880
rect 23920 36823 23943 36857
rect 23977 36823 24000 36857
rect 23920 36537 24000 36823
rect 23920 36503 23943 36537
rect 23977 36503 24000 36537
rect 23920 36480 24000 36503
rect 24080 36857 24160 36880
rect 24080 36823 24103 36857
rect 24137 36823 24160 36857
rect 24080 36537 24160 36823
rect 24080 36503 24103 36537
rect 24137 36503 24160 36537
rect 24080 36480 24160 36503
rect 24240 36857 24320 36880
rect 24240 36823 24263 36857
rect 24297 36823 24320 36857
rect 24240 36537 24320 36823
rect 24240 36503 24263 36537
rect 24297 36503 24320 36537
rect 24240 36480 24320 36503
rect 24400 36857 24480 36880
rect 24400 36823 24423 36857
rect 24457 36823 24480 36857
rect 24400 36537 24480 36823
rect 24400 36503 24423 36537
rect 24457 36503 24480 36537
rect 24400 36480 24480 36503
rect 24560 36857 24640 36880
rect 24560 36823 24583 36857
rect 24617 36823 24640 36857
rect 24560 36537 24640 36823
rect 24560 36503 24583 36537
rect 24617 36503 24640 36537
rect 24560 36480 24640 36503
rect 24720 36857 24800 36880
rect 24720 36823 24743 36857
rect 24777 36823 24800 36857
rect 24720 36537 24800 36823
rect 24720 36503 24743 36537
rect 24777 36503 24800 36537
rect 24720 36480 24800 36503
rect 24880 36857 24960 36880
rect 24880 36823 24903 36857
rect 24937 36823 24960 36857
rect 24880 36537 24960 36823
rect 24880 36503 24903 36537
rect 24937 36503 24960 36537
rect 24880 36480 24960 36503
rect 25040 36857 25120 36880
rect 25040 36823 25063 36857
rect 25097 36823 25120 36857
rect 25040 36537 25120 36823
rect 25040 36503 25063 36537
rect 25097 36503 25120 36537
rect 25040 36480 25120 36503
rect 25200 36857 25280 36880
rect 25200 36823 25223 36857
rect 25257 36823 25280 36857
rect 25200 36537 25280 36823
rect 25200 36503 25223 36537
rect 25257 36503 25280 36537
rect 25200 36480 25280 36503
rect 25360 36857 25440 36880
rect 25360 36823 25383 36857
rect 25417 36823 25440 36857
rect 25360 36537 25440 36823
rect 25360 36503 25383 36537
rect 25417 36503 25440 36537
rect 25360 36480 25440 36503
rect 25520 36857 25600 36880
rect 25520 36823 25543 36857
rect 25577 36823 25600 36857
rect 25520 36537 25600 36823
rect 25520 36503 25543 36537
rect 25577 36503 25600 36537
rect 25520 36480 25600 36503
rect 25680 36857 25760 36880
rect 25680 36823 25703 36857
rect 25737 36823 25760 36857
rect 25680 36537 25760 36823
rect 25680 36503 25703 36537
rect 25737 36503 25760 36537
rect 25680 36480 25760 36503
rect 25840 36857 25920 36880
rect 25840 36823 25863 36857
rect 25897 36823 25920 36857
rect 25840 36537 25920 36823
rect 25840 36503 25863 36537
rect 25897 36503 25920 36537
rect 25840 36480 25920 36503
rect 26000 36857 26080 36880
rect 26000 36823 26023 36857
rect 26057 36823 26080 36857
rect 26000 36537 26080 36823
rect 26000 36503 26023 36537
rect 26057 36503 26080 36537
rect 26000 36480 26080 36503
rect 26160 36857 26240 36880
rect 26160 36823 26183 36857
rect 26217 36823 26240 36857
rect 26160 36537 26240 36823
rect 26160 36503 26183 36537
rect 26217 36503 26240 36537
rect 26160 36480 26240 36503
rect 26320 36857 26400 36880
rect 26320 36823 26343 36857
rect 26377 36823 26400 36857
rect 26320 36537 26400 36823
rect 26320 36503 26343 36537
rect 26377 36503 26400 36537
rect 26320 36480 26400 36503
rect 26480 36857 26560 36880
rect 26480 36823 26503 36857
rect 26537 36823 26560 36857
rect 26480 36537 26560 36823
rect 26480 36503 26503 36537
rect 26537 36503 26560 36537
rect 26480 36480 26560 36503
rect 26640 36857 26720 36880
rect 26640 36823 26663 36857
rect 26697 36823 26720 36857
rect 26640 36537 26720 36823
rect 26640 36503 26663 36537
rect 26697 36503 26720 36537
rect 26640 36480 26720 36503
rect 26800 36857 26880 36880
rect 26800 36823 26823 36857
rect 26857 36823 26880 36857
rect 26800 36537 26880 36823
rect 26800 36503 26823 36537
rect 26857 36503 26880 36537
rect 26800 36480 26880 36503
rect 26960 36857 27040 36880
rect 26960 36823 26983 36857
rect 27017 36823 27040 36857
rect 26960 36537 27040 36823
rect 26960 36503 26983 36537
rect 27017 36503 27040 36537
rect 26960 36480 27040 36503
rect 27120 36857 27200 36880
rect 27120 36823 27143 36857
rect 27177 36823 27200 36857
rect 27120 36537 27200 36823
rect 27120 36503 27143 36537
rect 27177 36503 27200 36537
rect 27120 36480 27200 36503
rect 27280 36857 27360 36880
rect 27280 36823 27303 36857
rect 27337 36823 27360 36857
rect 27280 36537 27360 36823
rect 27280 36503 27303 36537
rect 27337 36503 27360 36537
rect 27280 36480 27360 36503
rect 27440 36857 27520 36880
rect 27440 36823 27463 36857
rect 27497 36823 27520 36857
rect 27440 36537 27520 36823
rect 27440 36503 27463 36537
rect 27497 36503 27520 36537
rect 27440 36480 27520 36503
rect 27600 36857 27680 36880
rect 27600 36823 27623 36857
rect 27657 36823 27680 36857
rect 27600 36537 27680 36823
rect 27600 36503 27623 36537
rect 27657 36503 27680 36537
rect 27600 36480 27680 36503
rect 27760 36857 27840 36880
rect 27760 36823 27783 36857
rect 27817 36823 27840 36857
rect 27760 36537 27840 36823
rect 27760 36503 27783 36537
rect 27817 36503 27840 36537
rect 27760 36480 27840 36503
rect 27920 36857 28000 36880
rect 27920 36823 27943 36857
rect 27977 36823 28000 36857
rect 27920 36537 28000 36823
rect 27920 36503 27943 36537
rect 27977 36503 28000 36537
rect 27920 36480 28000 36503
rect 28080 36857 28160 36880
rect 28080 36823 28103 36857
rect 28137 36823 28160 36857
rect 28080 36537 28160 36823
rect 28080 36503 28103 36537
rect 28137 36503 28160 36537
rect 28080 36480 28160 36503
rect 28240 36857 28320 36880
rect 28240 36823 28263 36857
rect 28297 36823 28320 36857
rect 28240 36537 28320 36823
rect 28240 36503 28263 36537
rect 28297 36503 28320 36537
rect 28240 36480 28320 36503
rect 28400 36857 28480 36880
rect 28400 36823 28423 36857
rect 28457 36823 28480 36857
rect 28400 36537 28480 36823
rect 28400 36503 28423 36537
rect 28457 36503 28480 36537
rect 28400 36480 28480 36503
rect 28560 36857 28640 36880
rect 28560 36823 28583 36857
rect 28617 36823 28640 36857
rect 28560 36537 28640 36823
rect 28560 36503 28583 36537
rect 28617 36503 28640 36537
rect 28560 36480 28640 36503
rect 28720 36857 28800 36880
rect 28720 36823 28743 36857
rect 28777 36823 28800 36857
rect 28720 36537 28800 36823
rect 28720 36503 28743 36537
rect 28777 36503 28800 36537
rect 28720 36480 28800 36503
rect 28880 36857 28960 36880
rect 28880 36823 28903 36857
rect 28937 36823 28960 36857
rect 28880 36537 28960 36823
rect 28880 36503 28903 36537
rect 28937 36503 28960 36537
rect 28880 36480 28960 36503
rect 29040 36857 29120 36880
rect 29040 36823 29063 36857
rect 29097 36823 29120 36857
rect 29040 36537 29120 36823
rect 29040 36503 29063 36537
rect 29097 36503 29120 36537
rect 29040 36480 29120 36503
rect 29200 36857 29280 36880
rect 29200 36823 29223 36857
rect 29257 36823 29280 36857
rect 29200 36537 29280 36823
rect 29200 36503 29223 36537
rect 29257 36503 29280 36537
rect 29200 36480 29280 36503
rect 29360 36857 29440 36880
rect 29360 36823 29383 36857
rect 29417 36823 29440 36857
rect 29360 36537 29440 36823
rect 29360 36503 29383 36537
rect 29417 36503 29440 36537
rect 29360 36480 29440 36503
rect 29520 36480 29600 36880
rect 29680 36480 29760 36880
rect 29840 36480 29920 36880
rect 30000 36480 30080 36880
rect 30160 36480 30240 36880
rect 30320 36480 30400 36880
rect 30480 36480 30560 36880
rect 30640 36480 30720 36880
rect 30800 36480 30880 36880
rect 30960 36480 31040 36880
rect 31120 36480 31200 36880
rect 31280 36480 31360 36880
rect 31440 36480 31520 36880
rect 31600 36480 31680 36880
rect 31760 36480 31840 36880
rect 31920 36480 32000 36880
rect 32080 36480 32160 36880
rect 32240 36480 32320 36880
rect 32400 36480 32480 36880
rect 32560 36480 32640 36880
rect 32720 36480 32800 36880
rect 32880 36480 32960 36880
rect 33040 36480 33120 36880
rect 33200 36480 33280 36880
rect 33360 36480 33440 36880
rect 33520 36857 33600 36880
rect 33520 36823 33543 36857
rect 33577 36823 33600 36857
rect 33520 36537 33600 36823
rect 33520 36503 33543 36537
rect 33577 36503 33600 36537
rect 33520 36480 33600 36503
rect 33680 36857 33760 36880
rect 33680 36823 33703 36857
rect 33737 36823 33760 36857
rect 33680 36537 33760 36823
rect 33680 36503 33703 36537
rect 33737 36503 33760 36537
rect 33680 36480 33760 36503
rect 33840 36857 33920 36880
rect 33840 36823 33863 36857
rect 33897 36823 33920 36857
rect 33840 36537 33920 36823
rect 33840 36503 33863 36537
rect 33897 36503 33920 36537
rect 33840 36480 33920 36503
rect 34000 36857 34080 36880
rect 34000 36823 34023 36857
rect 34057 36823 34080 36857
rect 34000 36537 34080 36823
rect 34000 36503 34023 36537
rect 34057 36503 34080 36537
rect 34000 36480 34080 36503
rect 34160 36857 34240 36880
rect 34160 36823 34183 36857
rect 34217 36823 34240 36857
rect 34160 36537 34240 36823
rect 34160 36503 34183 36537
rect 34217 36503 34240 36537
rect 34160 36480 34240 36503
rect 34320 36857 34400 36880
rect 34320 36823 34343 36857
rect 34377 36823 34400 36857
rect 34320 36537 34400 36823
rect 34320 36503 34343 36537
rect 34377 36503 34400 36537
rect 34320 36480 34400 36503
rect 34480 36857 34560 36880
rect 34480 36823 34503 36857
rect 34537 36823 34560 36857
rect 34480 36537 34560 36823
rect 34480 36503 34503 36537
rect 34537 36503 34560 36537
rect 34480 36480 34560 36503
rect 34640 36857 34720 36880
rect 34640 36823 34663 36857
rect 34697 36823 34720 36857
rect 34640 36537 34720 36823
rect 34640 36503 34663 36537
rect 34697 36503 34720 36537
rect 34640 36480 34720 36503
rect 34800 36857 34880 36880
rect 34800 36823 34823 36857
rect 34857 36823 34880 36857
rect 34800 36537 34880 36823
rect 34800 36503 34823 36537
rect 34857 36503 34880 36537
rect 34800 36480 34880 36503
rect 34960 36857 35040 36880
rect 34960 36823 34983 36857
rect 35017 36823 35040 36857
rect 34960 36537 35040 36823
rect 34960 36503 34983 36537
rect 35017 36503 35040 36537
rect 34960 36480 35040 36503
rect 35120 36857 35200 36880
rect 35120 36823 35143 36857
rect 35177 36823 35200 36857
rect 35120 36537 35200 36823
rect 35120 36503 35143 36537
rect 35177 36503 35200 36537
rect 35120 36480 35200 36503
rect 35280 36857 35360 36880
rect 35280 36823 35303 36857
rect 35337 36823 35360 36857
rect 35280 36537 35360 36823
rect 35280 36503 35303 36537
rect 35337 36503 35360 36537
rect 35280 36480 35360 36503
rect 35440 36857 35520 36880
rect 35440 36823 35463 36857
rect 35497 36823 35520 36857
rect 35440 36537 35520 36823
rect 35440 36503 35463 36537
rect 35497 36503 35520 36537
rect 35440 36480 35520 36503
rect 35600 36857 35680 36880
rect 35600 36823 35623 36857
rect 35657 36823 35680 36857
rect 35600 36537 35680 36823
rect 35600 36503 35623 36537
rect 35657 36503 35680 36537
rect 35600 36480 35680 36503
rect 35760 36857 35840 36880
rect 35760 36823 35783 36857
rect 35817 36823 35840 36857
rect 35760 36537 35840 36823
rect 35760 36503 35783 36537
rect 35817 36503 35840 36537
rect 35760 36480 35840 36503
rect 35920 36857 36000 36880
rect 35920 36823 35943 36857
rect 35977 36823 36000 36857
rect 35920 36537 36000 36823
rect 35920 36503 35943 36537
rect 35977 36503 36000 36537
rect 35920 36480 36000 36503
rect 36080 36857 36160 36880
rect 36080 36823 36103 36857
rect 36137 36823 36160 36857
rect 36080 36537 36160 36823
rect 36080 36503 36103 36537
rect 36137 36503 36160 36537
rect 36080 36480 36160 36503
rect 36240 36857 36320 36880
rect 36240 36823 36263 36857
rect 36297 36823 36320 36857
rect 36240 36537 36320 36823
rect 36240 36503 36263 36537
rect 36297 36503 36320 36537
rect 36240 36480 36320 36503
rect 36400 36857 36480 36880
rect 36400 36823 36423 36857
rect 36457 36823 36480 36857
rect 36400 36537 36480 36823
rect 36400 36503 36423 36537
rect 36457 36503 36480 36537
rect 36400 36480 36480 36503
rect 36560 36857 36640 36880
rect 36560 36823 36583 36857
rect 36617 36823 36640 36857
rect 36560 36537 36640 36823
rect 36560 36503 36583 36537
rect 36617 36503 36640 36537
rect 36560 36480 36640 36503
rect 36720 36857 36800 36880
rect 36720 36823 36743 36857
rect 36777 36823 36800 36857
rect 36720 36537 36800 36823
rect 36720 36503 36743 36537
rect 36777 36503 36800 36537
rect 36720 36480 36800 36503
rect 36880 36857 36960 36880
rect 36880 36823 36903 36857
rect 36937 36823 36960 36857
rect 36880 36537 36960 36823
rect 36880 36503 36903 36537
rect 36937 36503 36960 36537
rect 36880 36480 36960 36503
rect 37040 36857 37120 36880
rect 37040 36823 37063 36857
rect 37097 36823 37120 36857
rect 37040 36537 37120 36823
rect 37040 36503 37063 36537
rect 37097 36503 37120 36537
rect 37040 36480 37120 36503
rect 37200 36857 37280 36880
rect 37200 36823 37223 36857
rect 37257 36823 37280 36857
rect 37200 36537 37280 36823
rect 37200 36503 37223 36537
rect 37257 36503 37280 36537
rect 37200 36480 37280 36503
rect 37360 36857 37440 36880
rect 37360 36823 37383 36857
rect 37417 36823 37440 36857
rect 37360 36537 37440 36823
rect 37360 36503 37383 36537
rect 37417 36503 37440 36537
rect 37360 36480 37440 36503
rect 37520 36857 37600 36880
rect 37520 36823 37543 36857
rect 37577 36823 37600 36857
rect 37520 36537 37600 36823
rect 37520 36503 37543 36537
rect 37577 36503 37600 36537
rect 37520 36480 37600 36503
rect 37680 36857 37760 36880
rect 37680 36823 37703 36857
rect 37737 36823 37760 36857
rect 37680 36537 37760 36823
rect 37680 36503 37703 36537
rect 37737 36503 37760 36537
rect 37680 36480 37760 36503
rect 37840 36857 37920 36880
rect 37840 36823 37863 36857
rect 37897 36823 37920 36857
rect 37840 36537 37920 36823
rect 37840 36503 37863 36537
rect 37897 36503 37920 36537
rect 37840 36480 37920 36503
rect 38000 36857 38080 36880
rect 38000 36823 38023 36857
rect 38057 36823 38080 36857
rect 38000 36537 38080 36823
rect 38000 36503 38023 36537
rect 38057 36503 38080 36537
rect 38000 36480 38080 36503
rect 38160 36857 38240 36880
rect 38160 36823 38183 36857
rect 38217 36823 38240 36857
rect 38160 36537 38240 36823
rect 38160 36503 38183 36537
rect 38217 36503 38240 36537
rect 38160 36480 38240 36503
rect 38320 36857 38400 36880
rect 38320 36823 38343 36857
rect 38377 36823 38400 36857
rect 38320 36537 38400 36823
rect 38320 36503 38343 36537
rect 38377 36503 38400 36537
rect 38320 36480 38400 36503
rect 38480 36857 38560 36880
rect 38480 36823 38503 36857
rect 38537 36823 38560 36857
rect 38480 36537 38560 36823
rect 38480 36503 38503 36537
rect 38537 36503 38560 36537
rect 38480 36480 38560 36503
rect 38640 36857 38720 36880
rect 38640 36823 38663 36857
rect 38697 36823 38720 36857
rect 38640 36537 38720 36823
rect 38640 36503 38663 36537
rect 38697 36503 38720 36537
rect 38640 36480 38720 36503
rect 38800 36857 38880 36880
rect 38800 36823 38823 36857
rect 38857 36823 38880 36857
rect 38800 36537 38880 36823
rect 38800 36503 38823 36537
rect 38857 36503 38880 36537
rect 38800 36480 38880 36503
rect 38960 36857 39040 36880
rect 38960 36823 38983 36857
rect 39017 36823 39040 36857
rect 38960 36537 39040 36823
rect 38960 36503 38983 36537
rect 39017 36503 39040 36537
rect 38960 36480 39040 36503
rect 39120 36857 39200 36880
rect 39120 36823 39143 36857
rect 39177 36823 39200 36857
rect 39120 36537 39200 36823
rect 39120 36503 39143 36537
rect 39177 36503 39200 36537
rect 39120 36480 39200 36503
rect 39280 36857 39360 36880
rect 39280 36823 39303 36857
rect 39337 36823 39360 36857
rect 39280 36537 39360 36823
rect 39280 36503 39303 36537
rect 39337 36503 39360 36537
rect 39280 36480 39360 36503
rect 39440 36857 39520 36880
rect 39440 36823 39463 36857
rect 39497 36823 39520 36857
rect 39440 36537 39520 36823
rect 39440 36503 39463 36537
rect 39497 36503 39520 36537
rect 39440 36480 39520 36503
rect 39600 36857 39680 36880
rect 39600 36823 39623 36857
rect 39657 36823 39680 36857
rect 39600 36537 39680 36823
rect 39600 36503 39623 36537
rect 39657 36503 39680 36537
rect 39600 36480 39680 36503
rect 39760 36857 39840 36880
rect 39760 36823 39783 36857
rect 39817 36823 39840 36857
rect 39760 36537 39840 36823
rect 39760 36503 39783 36537
rect 39817 36503 39840 36537
rect 39760 36480 39840 36503
rect 39920 36857 40000 36880
rect 39920 36823 39943 36857
rect 39977 36823 40000 36857
rect 39920 36537 40000 36823
rect 39920 36503 39943 36537
rect 39977 36503 40000 36537
rect 39920 36480 40000 36503
rect 40080 36857 40160 36880
rect 40080 36823 40103 36857
rect 40137 36823 40160 36857
rect 40080 36537 40160 36823
rect 40080 36503 40103 36537
rect 40137 36503 40160 36537
rect 40080 36480 40160 36503
rect 40240 36857 40320 36880
rect 40240 36823 40263 36857
rect 40297 36823 40320 36857
rect 40240 36537 40320 36823
rect 40240 36503 40263 36537
rect 40297 36503 40320 36537
rect 40240 36480 40320 36503
rect 40400 36857 40480 36880
rect 40400 36823 40423 36857
rect 40457 36823 40480 36857
rect 40400 36537 40480 36823
rect 40400 36503 40423 36537
rect 40457 36503 40480 36537
rect 40400 36480 40480 36503
rect 40560 36857 40640 36880
rect 40560 36823 40583 36857
rect 40617 36823 40640 36857
rect 40560 36537 40640 36823
rect 40560 36503 40583 36537
rect 40617 36503 40640 36537
rect 40560 36480 40640 36503
rect 40720 36857 40800 36880
rect 40720 36823 40743 36857
rect 40777 36823 40800 36857
rect 40720 36537 40800 36823
rect 40720 36503 40743 36537
rect 40777 36503 40800 36537
rect 40720 36480 40800 36503
rect 40880 36857 40960 36880
rect 40880 36823 40903 36857
rect 40937 36823 40960 36857
rect 40880 36537 40960 36823
rect 40880 36503 40903 36537
rect 40937 36503 40960 36537
rect 40880 36480 40960 36503
rect 41040 36857 41120 36880
rect 41040 36823 41063 36857
rect 41097 36823 41120 36857
rect 41040 36537 41120 36823
rect 41040 36503 41063 36537
rect 41097 36503 41120 36537
rect 41040 36480 41120 36503
rect 41200 36857 41280 36880
rect 41200 36823 41223 36857
rect 41257 36823 41280 36857
rect 41200 36537 41280 36823
rect 41200 36503 41223 36537
rect 41257 36503 41280 36537
rect 41200 36480 41280 36503
rect 41360 36857 41440 36880
rect 41360 36823 41383 36857
rect 41417 36823 41440 36857
rect 41360 36537 41440 36823
rect 41360 36503 41383 36537
rect 41417 36503 41440 36537
rect 41360 36480 41440 36503
rect 41520 36857 41600 36880
rect 41520 36823 41543 36857
rect 41577 36823 41600 36857
rect 41520 36537 41600 36823
rect 41520 36503 41543 36537
rect 41577 36503 41600 36537
rect 41520 36480 41600 36503
rect 41680 36857 41760 36880
rect 41680 36823 41703 36857
rect 41737 36823 41760 36857
rect 41680 36537 41760 36823
rect 41680 36503 41703 36537
rect 41737 36503 41760 36537
rect 41680 36480 41760 36503
rect 41840 36857 41920 36880
rect 41840 36823 41863 36857
rect 41897 36823 41920 36857
rect 41840 36537 41920 36823
rect 41840 36503 41863 36537
rect 41897 36503 41920 36537
rect 41840 36480 41920 36503
rect 0 36377 80 36400
rect 0 36343 23 36377
rect 57 36343 80 36377
rect 0 36057 80 36343
rect 0 36023 23 36057
rect 57 36023 80 36057
rect 0 35737 80 36023
rect 0 35703 23 35737
rect 57 35703 80 35737
rect 0 35417 80 35703
rect 0 35383 23 35417
rect 57 35383 80 35417
rect 0 35097 80 35383
rect 0 35063 23 35097
rect 57 35063 80 35097
rect 0 34777 80 35063
rect 0 34743 23 34777
rect 57 34743 80 34777
rect 0 34457 80 34743
rect 0 34423 23 34457
rect 57 34423 80 34457
rect 0 34400 80 34423
rect 160 36377 240 36400
rect 160 36343 183 36377
rect 217 36343 240 36377
rect 160 36057 240 36343
rect 160 36023 183 36057
rect 217 36023 240 36057
rect 160 35737 240 36023
rect 160 35703 183 35737
rect 217 35703 240 35737
rect 160 35417 240 35703
rect 160 35383 183 35417
rect 217 35383 240 35417
rect 160 35097 240 35383
rect 160 35063 183 35097
rect 217 35063 240 35097
rect 160 34777 240 35063
rect 160 34743 183 34777
rect 217 34743 240 34777
rect 160 34457 240 34743
rect 160 34423 183 34457
rect 217 34423 240 34457
rect 160 34400 240 34423
rect 320 36377 400 36400
rect 320 36343 343 36377
rect 377 36343 400 36377
rect 320 36057 400 36343
rect 320 36023 343 36057
rect 377 36023 400 36057
rect 320 35737 400 36023
rect 320 35703 343 35737
rect 377 35703 400 35737
rect 320 35417 400 35703
rect 320 35383 343 35417
rect 377 35383 400 35417
rect 320 35097 400 35383
rect 320 35063 343 35097
rect 377 35063 400 35097
rect 320 34777 400 35063
rect 320 34743 343 34777
rect 377 34743 400 34777
rect 320 34457 400 34743
rect 320 34423 343 34457
rect 377 34423 400 34457
rect 320 34400 400 34423
rect 480 36377 560 36400
rect 480 36343 503 36377
rect 537 36343 560 36377
rect 480 36057 560 36343
rect 480 36023 503 36057
rect 537 36023 560 36057
rect 480 35737 560 36023
rect 480 35703 503 35737
rect 537 35703 560 35737
rect 480 35417 560 35703
rect 480 35383 503 35417
rect 537 35383 560 35417
rect 480 35097 560 35383
rect 480 35063 503 35097
rect 537 35063 560 35097
rect 480 34777 560 35063
rect 480 34743 503 34777
rect 537 34743 560 34777
rect 480 34457 560 34743
rect 480 34423 503 34457
rect 537 34423 560 34457
rect 480 34400 560 34423
rect 640 36377 720 36400
rect 640 36343 663 36377
rect 697 36343 720 36377
rect 640 36057 720 36343
rect 640 36023 663 36057
rect 697 36023 720 36057
rect 640 35737 720 36023
rect 640 35703 663 35737
rect 697 35703 720 35737
rect 640 35417 720 35703
rect 640 35383 663 35417
rect 697 35383 720 35417
rect 640 35097 720 35383
rect 640 35063 663 35097
rect 697 35063 720 35097
rect 640 34777 720 35063
rect 640 34743 663 34777
rect 697 34743 720 34777
rect 640 34457 720 34743
rect 640 34423 663 34457
rect 697 34423 720 34457
rect 640 34400 720 34423
rect 800 36377 880 36400
rect 800 36343 823 36377
rect 857 36343 880 36377
rect 800 36057 880 36343
rect 800 36023 823 36057
rect 857 36023 880 36057
rect 800 35737 880 36023
rect 800 35703 823 35737
rect 857 35703 880 35737
rect 800 35417 880 35703
rect 800 35383 823 35417
rect 857 35383 880 35417
rect 800 35097 880 35383
rect 800 35063 823 35097
rect 857 35063 880 35097
rect 800 34777 880 35063
rect 800 34743 823 34777
rect 857 34743 880 34777
rect 800 34457 880 34743
rect 800 34423 823 34457
rect 857 34423 880 34457
rect 800 34400 880 34423
rect 960 36377 1040 36400
rect 960 36343 983 36377
rect 1017 36343 1040 36377
rect 960 36057 1040 36343
rect 960 36023 983 36057
rect 1017 36023 1040 36057
rect 960 35737 1040 36023
rect 960 35703 983 35737
rect 1017 35703 1040 35737
rect 960 35417 1040 35703
rect 960 35383 983 35417
rect 1017 35383 1040 35417
rect 960 35097 1040 35383
rect 960 35063 983 35097
rect 1017 35063 1040 35097
rect 960 34777 1040 35063
rect 960 34743 983 34777
rect 1017 34743 1040 34777
rect 960 34457 1040 34743
rect 960 34423 983 34457
rect 1017 34423 1040 34457
rect 960 34400 1040 34423
rect 1120 36377 1200 36400
rect 1120 36343 1143 36377
rect 1177 36343 1200 36377
rect 1120 36057 1200 36343
rect 1120 36023 1143 36057
rect 1177 36023 1200 36057
rect 1120 35737 1200 36023
rect 1120 35703 1143 35737
rect 1177 35703 1200 35737
rect 1120 35417 1200 35703
rect 1120 35383 1143 35417
rect 1177 35383 1200 35417
rect 1120 35097 1200 35383
rect 1120 35063 1143 35097
rect 1177 35063 1200 35097
rect 1120 34777 1200 35063
rect 1120 34743 1143 34777
rect 1177 34743 1200 34777
rect 1120 34457 1200 34743
rect 1120 34423 1143 34457
rect 1177 34423 1200 34457
rect 1120 34400 1200 34423
rect 1280 36377 1360 36400
rect 1280 36343 1303 36377
rect 1337 36343 1360 36377
rect 1280 36057 1360 36343
rect 1280 36023 1303 36057
rect 1337 36023 1360 36057
rect 1280 35737 1360 36023
rect 1280 35703 1303 35737
rect 1337 35703 1360 35737
rect 1280 35417 1360 35703
rect 1280 35383 1303 35417
rect 1337 35383 1360 35417
rect 1280 35097 1360 35383
rect 1280 35063 1303 35097
rect 1337 35063 1360 35097
rect 1280 34777 1360 35063
rect 1280 34743 1303 34777
rect 1337 34743 1360 34777
rect 1280 34457 1360 34743
rect 1280 34423 1303 34457
rect 1337 34423 1360 34457
rect 1280 34400 1360 34423
rect 1440 36377 1520 36400
rect 1440 36343 1463 36377
rect 1497 36343 1520 36377
rect 1440 36057 1520 36343
rect 1440 36023 1463 36057
rect 1497 36023 1520 36057
rect 1440 35737 1520 36023
rect 1440 35703 1463 35737
rect 1497 35703 1520 35737
rect 1440 35417 1520 35703
rect 1440 35383 1463 35417
rect 1497 35383 1520 35417
rect 1440 35097 1520 35383
rect 1440 35063 1463 35097
rect 1497 35063 1520 35097
rect 1440 34777 1520 35063
rect 1440 34743 1463 34777
rect 1497 34743 1520 34777
rect 1440 34457 1520 34743
rect 1440 34423 1463 34457
rect 1497 34423 1520 34457
rect 1440 34400 1520 34423
rect 1600 36377 1680 36400
rect 1600 36343 1623 36377
rect 1657 36343 1680 36377
rect 1600 36057 1680 36343
rect 1600 36023 1623 36057
rect 1657 36023 1680 36057
rect 1600 35737 1680 36023
rect 1600 35703 1623 35737
rect 1657 35703 1680 35737
rect 1600 35417 1680 35703
rect 1600 35383 1623 35417
rect 1657 35383 1680 35417
rect 1600 35097 1680 35383
rect 1600 35063 1623 35097
rect 1657 35063 1680 35097
rect 1600 34777 1680 35063
rect 1600 34743 1623 34777
rect 1657 34743 1680 34777
rect 1600 34457 1680 34743
rect 1600 34423 1623 34457
rect 1657 34423 1680 34457
rect 1600 34400 1680 34423
rect 1760 36377 1840 36400
rect 1760 36343 1783 36377
rect 1817 36343 1840 36377
rect 1760 36057 1840 36343
rect 1760 36023 1783 36057
rect 1817 36023 1840 36057
rect 1760 35737 1840 36023
rect 1760 35703 1783 35737
rect 1817 35703 1840 35737
rect 1760 35417 1840 35703
rect 1760 35383 1783 35417
rect 1817 35383 1840 35417
rect 1760 35097 1840 35383
rect 1760 35063 1783 35097
rect 1817 35063 1840 35097
rect 1760 34777 1840 35063
rect 1760 34743 1783 34777
rect 1817 34743 1840 34777
rect 1760 34457 1840 34743
rect 1760 34423 1783 34457
rect 1817 34423 1840 34457
rect 1760 34400 1840 34423
rect 1920 36377 2000 36400
rect 1920 36343 1943 36377
rect 1977 36343 2000 36377
rect 1920 36057 2000 36343
rect 1920 36023 1943 36057
rect 1977 36023 2000 36057
rect 1920 35737 2000 36023
rect 1920 35703 1943 35737
rect 1977 35703 2000 35737
rect 1920 35417 2000 35703
rect 1920 35383 1943 35417
rect 1977 35383 2000 35417
rect 1920 35097 2000 35383
rect 1920 35063 1943 35097
rect 1977 35063 2000 35097
rect 1920 34777 2000 35063
rect 1920 34743 1943 34777
rect 1977 34743 2000 34777
rect 1920 34457 2000 34743
rect 1920 34423 1943 34457
rect 1977 34423 2000 34457
rect 1920 34400 2000 34423
rect 2080 36377 2160 36400
rect 2080 36343 2103 36377
rect 2137 36343 2160 36377
rect 2080 36057 2160 36343
rect 2080 36023 2103 36057
rect 2137 36023 2160 36057
rect 2080 35737 2160 36023
rect 2080 35703 2103 35737
rect 2137 35703 2160 35737
rect 2080 35417 2160 35703
rect 2080 35383 2103 35417
rect 2137 35383 2160 35417
rect 2080 35097 2160 35383
rect 2080 35063 2103 35097
rect 2137 35063 2160 35097
rect 2080 34777 2160 35063
rect 2080 34743 2103 34777
rect 2137 34743 2160 34777
rect 2080 34457 2160 34743
rect 2080 34423 2103 34457
rect 2137 34423 2160 34457
rect 2080 34400 2160 34423
rect 2240 36377 2320 36400
rect 2240 36343 2263 36377
rect 2297 36343 2320 36377
rect 2240 36057 2320 36343
rect 2240 36023 2263 36057
rect 2297 36023 2320 36057
rect 2240 35737 2320 36023
rect 2240 35703 2263 35737
rect 2297 35703 2320 35737
rect 2240 35417 2320 35703
rect 2240 35383 2263 35417
rect 2297 35383 2320 35417
rect 2240 35097 2320 35383
rect 2240 35063 2263 35097
rect 2297 35063 2320 35097
rect 2240 34777 2320 35063
rect 2240 34743 2263 34777
rect 2297 34743 2320 34777
rect 2240 34457 2320 34743
rect 2240 34423 2263 34457
rect 2297 34423 2320 34457
rect 2240 34400 2320 34423
rect 2400 36377 2480 36400
rect 2400 36343 2423 36377
rect 2457 36343 2480 36377
rect 2400 36057 2480 36343
rect 2400 36023 2423 36057
rect 2457 36023 2480 36057
rect 2400 35737 2480 36023
rect 2400 35703 2423 35737
rect 2457 35703 2480 35737
rect 2400 35417 2480 35703
rect 2400 35383 2423 35417
rect 2457 35383 2480 35417
rect 2400 35097 2480 35383
rect 2400 35063 2423 35097
rect 2457 35063 2480 35097
rect 2400 34777 2480 35063
rect 2400 34743 2423 34777
rect 2457 34743 2480 34777
rect 2400 34457 2480 34743
rect 2400 34423 2423 34457
rect 2457 34423 2480 34457
rect 2400 34400 2480 34423
rect 2560 36377 2640 36400
rect 2560 36343 2583 36377
rect 2617 36343 2640 36377
rect 2560 36057 2640 36343
rect 2560 36023 2583 36057
rect 2617 36023 2640 36057
rect 2560 35737 2640 36023
rect 2560 35703 2583 35737
rect 2617 35703 2640 35737
rect 2560 35417 2640 35703
rect 2560 35383 2583 35417
rect 2617 35383 2640 35417
rect 2560 35097 2640 35383
rect 2560 35063 2583 35097
rect 2617 35063 2640 35097
rect 2560 34777 2640 35063
rect 2560 34743 2583 34777
rect 2617 34743 2640 34777
rect 2560 34457 2640 34743
rect 2560 34423 2583 34457
rect 2617 34423 2640 34457
rect 2560 34400 2640 34423
rect 2720 36377 2800 36400
rect 2720 36343 2743 36377
rect 2777 36343 2800 36377
rect 2720 36057 2800 36343
rect 2720 36023 2743 36057
rect 2777 36023 2800 36057
rect 2720 35737 2800 36023
rect 2720 35703 2743 35737
rect 2777 35703 2800 35737
rect 2720 35417 2800 35703
rect 2720 35383 2743 35417
rect 2777 35383 2800 35417
rect 2720 35097 2800 35383
rect 2720 35063 2743 35097
rect 2777 35063 2800 35097
rect 2720 34777 2800 35063
rect 2720 34743 2743 34777
rect 2777 34743 2800 34777
rect 2720 34457 2800 34743
rect 2720 34423 2743 34457
rect 2777 34423 2800 34457
rect 2720 34400 2800 34423
rect 2880 36377 2960 36400
rect 2880 36343 2903 36377
rect 2937 36343 2960 36377
rect 2880 36057 2960 36343
rect 2880 36023 2903 36057
rect 2937 36023 2960 36057
rect 2880 35737 2960 36023
rect 2880 35703 2903 35737
rect 2937 35703 2960 35737
rect 2880 35417 2960 35703
rect 2880 35383 2903 35417
rect 2937 35383 2960 35417
rect 2880 35097 2960 35383
rect 2880 35063 2903 35097
rect 2937 35063 2960 35097
rect 2880 34777 2960 35063
rect 2880 34743 2903 34777
rect 2937 34743 2960 34777
rect 2880 34457 2960 34743
rect 2880 34423 2903 34457
rect 2937 34423 2960 34457
rect 2880 34400 2960 34423
rect 3040 36377 3120 36400
rect 3040 36343 3063 36377
rect 3097 36343 3120 36377
rect 3040 36057 3120 36343
rect 3040 36023 3063 36057
rect 3097 36023 3120 36057
rect 3040 35737 3120 36023
rect 3040 35703 3063 35737
rect 3097 35703 3120 35737
rect 3040 35417 3120 35703
rect 3040 35383 3063 35417
rect 3097 35383 3120 35417
rect 3040 35097 3120 35383
rect 3040 35063 3063 35097
rect 3097 35063 3120 35097
rect 3040 34777 3120 35063
rect 3040 34743 3063 34777
rect 3097 34743 3120 34777
rect 3040 34457 3120 34743
rect 3040 34423 3063 34457
rect 3097 34423 3120 34457
rect 3040 34400 3120 34423
rect 3200 36377 3280 36400
rect 3200 36343 3223 36377
rect 3257 36343 3280 36377
rect 3200 36057 3280 36343
rect 3200 36023 3223 36057
rect 3257 36023 3280 36057
rect 3200 35737 3280 36023
rect 3200 35703 3223 35737
rect 3257 35703 3280 35737
rect 3200 35417 3280 35703
rect 3200 35383 3223 35417
rect 3257 35383 3280 35417
rect 3200 35097 3280 35383
rect 3200 35063 3223 35097
rect 3257 35063 3280 35097
rect 3200 34777 3280 35063
rect 3200 34743 3223 34777
rect 3257 34743 3280 34777
rect 3200 34457 3280 34743
rect 3200 34423 3223 34457
rect 3257 34423 3280 34457
rect 3200 34400 3280 34423
rect 3360 36377 3440 36400
rect 3360 36343 3383 36377
rect 3417 36343 3440 36377
rect 3360 36057 3440 36343
rect 3360 36023 3383 36057
rect 3417 36023 3440 36057
rect 3360 35737 3440 36023
rect 3360 35703 3383 35737
rect 3417 35703 3440 35737
rect 3360 35417 3440 35703
rect 3360 35383 3383 35417
rect 3417 35383 3440 35417
rect 3360 35097 3440 35383
rect 3360 35063 3383 35097
rect 3417 35063 3440 35097
rect 3360 34777 3440 35063
rect 3360 34743 3383 34777
rect 3417 34743 3440 34777
rect 3360 34457 3440 34743
rect 3360 34423 3383 34457
rect 3417 34423 3440 34457
rect 3360 34400 3440 34423
rect 3520 36377 3600 36400
rect 3520 36343 3543 36377
rect 3577 36343 3600 36377
rect 3520 36057 3600 36343
rect 3520 36023 3543 36057
rect 3577 36023 3600 36057
rect 3520 35737 3600 36023
rect 3520 35703 3543 35737
rect 3577 35703 3600 35737
rect 3520 35417 3600 35703
rect 3520 35383 3543 35417
rect 3577 35383 3600 35417
rect 3520 35097 3600 35383
rect 3520 35063 3543 35097
rect 3577 35063 3600 35097
rect 3520 34777 3600 35063
rect 3520 34743 3543 34777
rect 3577 34743 3600 34777
rect 3520 34457 3600 34743
rect 3520 34423 3543 34457
rect 3577 34423 3600 34457
rect 3520 34400 3600 34423
rect 3680 36377 3760 36400
rect 3680 36343 3703 36377
rect 3737 36343 3760 36377
rect 3680 36057 3760 36343
rect 3680 36023 3703 36057
rect 3737 36023 3760 36057
rect 3680 35737 3760 36023
rect 3680 35703 3703 35737
rect 3737 35703 3760 35737
rect 3680 35417 3760 35703
rect 3680 35383 3703 35417
rect 3737 35383 3760 35417
rect 3680 35097 3760 35383
rect 3680 35063 3703 35097
rect 3737 35063 3760 35097
rect 3680 34777 3760 35063
rect 3680 34743 3703 34777
rect 3737 34743 3760 34777
rect 3680 34457 3760 34743
rect 3680 34423 3703 34457
rect 3737 34423 3760 34457
rect 3680 34400 3760 34423
rect 3840 36377 3920 36400
rect 3840 36343 3863 36377
rect 3897 36343 3920 36377
rect 3840 36057 3920 36343
rect 3840 36023 3863 36057
rect 3897 36023 3920 36057
rect 3840 35737 3920 36023
rect 3840 35703 3863 35737
rect 3897 35703 3920 35737
rect 3840 35417 3920 35703
rect 3840 35383 3863 35417
rect 3897 35383 3920 35417
rect 3840 35097 3920 35383
rect 3840 35063 3863 35097
rect 3897 35063 3920 35097
rect 3840 34777 3920 35063
rect 3840 34743 3863 34777
rect 3897 34743 3920 34777
rect 3840 34457 3920 34743
rect 3840 34423 3863 34457
rect 3897 34423 3920 34457
rect 3840 34400 3920 34423
rect 4000 36377 4080 36400
rect 4000 36343 4023 36377
rect 4057 36343 4080 36377
rect 4000 36057 4080 36343
rect 4000 36023 4023 36057
rect 4057 36023 4080 36057
rect 4000 35737 4080 36023
rect 4000 35703 4023 35737
rect 4057 35703 4080 35737
rect 4000 35417 4080 35703
rect 4000 35383 4023 35417
rect 4057 35383 4080 35417
rect 4000 35097 4080 35383
rect 4000 35063 4023 35097
rect 4057 35063 4080 35097
rect 4000 34777 4080 35063
rect 4000 34743 4023 34777
rect 4057 34743 4080 34777
rect 4000 34457 4080 34743
rect 4000 34423 4023 34457
rect 4057 34423 4080 34457
rect 4000 34400 4080 34423
rect 4160 36377 4240 36400
rect 4160 36343 4183 36377
rect 4217 36343 4240 36377
rect 4160 36057 4240 36343
rect 4160 36023 4183 36057
rect 4217 36023 4240 36057
rect 4160 35737 4240 36023
rect 4160 35703 4183 35737
rect 4217 35703 4240 35737
rect 4160 35417 4240 35703
rect 4160 35383 4183 35417
rect 4217 35383 4240 35417
rect 4160 35097 4240 35383
rect 4160 35063 4183 35097
rect 4217 35063 4240 35097
rect 4160 34777 4240 35063
rect 4160 34743 4183 34777
rect 4217 34743 4240 34777
rect 4160 34457 4240 34743
rect 4160 34423 4183 34457
rect 4217 34423 4240 34457
rect 4160 34400 4240 34423
rect 4320 36377 4400 36400
rect 4320 36343 4343 36377
rect 4377 36343 4400 36377
rect 4320 36057 4400 36343
rect 4320 36023 4343 36057
rect 4377 36023 4400 36057
rect 4320 35737 4400 36023
rect 4320 35703 4343 35737
rect 4377 35703 4400 35737
rect 4320 35417 4400 35703
rect 4320 35383 4343 35417
rect 4377 35383 4400 35417
rect 4320 35097 4400 35383
rect 4320 35063 4343 35097
rect 4377 35063 4400 35097
rect 4320 34777 4400 35063
rect 4320 34743 4343 34777
rect 4377 34743 4400 34777
rect 4320 34457 4400 34743
rect 4320 34423 4343 34457
rect 4377 34423 4400 34457
rect 4320 34400 4400 34423
rect 4480 36377 4560 36400
rect 4480 36343 4503 36377
rect 4537 36343 4560 36377
rect 4480 36057 4560 36343
rect 4480 36023 4503 36057
rect 4537 36023 4560 36057
rect 4480 35737 4560 36023
rect 4480 35703 4503 35737
rect 4537 35703 4560 35737
rect 4480 35417 4560 35703
rect 4480 35383 4503 35417
rect 4537 35383 4560 35417
rect 4480 35097 4560 35383
rect 4480 35063 4503 35097
rect 4537 35063 4560 35097
rect 4480 34777 4560 35063
rect 4480 34743 4503 34777
rect 4537 34743 4560 34777
rect 4480 34457 4560 34743
rect 4480 34423 4503 34457
rect 4537 34423 4560 34457
rect 4480 34400 4560 34423
rect 4640 36377 4720 36400
rect 4640 36343 4663 36377
rect 4697 36343 4720 36377
rect 4640 36057 4720 36343
rect 4640 36023 4663 36057
rect 4697 36023 4720 36057
rect 4640 35737 4720 36023
rect 4640 35703 4663 35737
rect 4697 35703 4720 35737
rect 4640 35417 4720 35703
rect 4640 35383 4663 35417
rect 4697 35383 4720 35417
rect 4640 35097 4720 35383
rect 4640 35063 4663 35097
rect 4697 35063 4720 35097
rect 4640 34777 4720 35063
rect 4640 34743 4663 34777
rect 4697 34743 4720 34777
rect 4640 34457 4720 34743
rect 4640 34423 4663 34457
rect 4697 34423 4720 34457
rect 4640 34400 4720 34423
rect 4800 36377 4880 36400
rect 4800 36343 4823 36377
rect 4857 36343 4880 36377
rect 4800 36057 4880 36343
rect 4800 36023 4823 36057
rect 4857 36023 4880 36057
rect 4800 35737 4880 36023
rect 4800 35703 4823 35737
rect 4857 35703 4880 35737
rect 4800 35417 4880 35703
rect 4800 35383 4823 35417
rect 4857 35383 4880 35417
rect 4800 35097 4880 35383
rect 4800 35063 4823 35097
rect 4857 35063 4880 35097
rect 4800 34777 4880 35063
rect 4800 34743 4823 34777
rect 4857 34743 4880 34777
rect 4800 34457 4880 34743
rect 4800 34423 4823 34457
rect 4857 34423 4880 34457
rect 4800 34400 4880 34423
rect 4960 36377 5040 36400
rect 4960 36343 4983 36377
rect 5017 36343 5040 36377
rect 4960 36057 5040 36343
rect 4960 36023 4983 36057
rect 5017 36023 5040 36057
rect 4960 35737 5040 36023
rect 4960 35703 4983 35737
rect 5017 35703 5040 35737
rect 4960 35417 5040 35703
rect 4960 35383 4983 35417
rect 5017 35383 5040 35417
rect 4960 35097 5040 35383
rect 4960 35063 4983 35097
rect 5017 35063 5040 35097
rect 4960 34777 5040 35063
rect 4960 34743 4983 34777
rect 5017 34743 5040 34777
rect 4960 34457 5040 34743
rect 4960 34423 4983 34457
rect 5017 34423 5040 34457
rect 4960 34400 5040 34423
rect 5120 36377 5200 36400
rect 5120 36343 5143 36377
rect 5177 36343 5200 36377
rect 5120 36057 5200 36343
rect 5120 36023 5143 36057
rect 5177 36023 5200 36057
rect 5120 35737 5200 36023
rect 5120 35703 5143 35737
rect 5177 35703 5200 35737
rect 5120 35417 5200 35703
rect 5120 35383 5143 35417
rect 5177 35383 5200 35417
rect 5120 35097 5200 35383
rect 5120 35063 5143 35097
rect 5177 35063 5200 35097
rect 5120 34777 5200 35063
rect 5120 34743 5143 34777
rect 5177 34743 5200 34777
rect 5120 34457 5200 34743
rect 5120 34423 5143 34457
rect 5177 34423 5200 34457
rect 5120 34400 5200 34423
rect 5280 36377 5360 36400
rect 5280 36343 5303 36377
rect 5337 36343 5360 36377
rect 5280 36057 5360 36343
rect 5280 36023 5303 36057
rect 5337 36023 5360 36057
rect 5280 35737 5360 36023
rect 5280 35703 5303 35737
rect 5337 35703 5360 35737
rect 5280 35417 5360 35703
rect 5280 35383 5303 35417
rect 5337 35383 5360 35417
rect 5280 35097 5360 35383
rect 5280 35063 5303 35097
rect 5337 35063 5360 35097
rect 5280 34777 5360 35063
rect 5280 34743 5303 34777
rect 5337 34743 5360 34777
rect 5280 34457 5360 34743
rect 5280 34423 5303 34457
rect 5337 34423 5360 34457
rect 5280 34400 5360 34423
rect 5440 36377 5520 36400
rect 5440 36343 5463 36377
rect 5497 36343 5520 36377
rect 5440 36057 5520 36343
rect 5440 36023 5463 36057
rect 5497 36023 5520 36057
rect 5440 35737 5520 36023
rect 5440 35703 5463 35737
rect 5497 35703 5520 35737
rect 5440 35417 5520 35703
rect 5440 35383 5463 35417
rect 5497 35383 5520 35417
rect 5440 35097 5520 35383
rect 5440 35063 5463 35097
rect 5497 35063 5520 35097
rect 5440 34777 5520 35063
rect 5440 34743 5463 34777
rect 5497 34743 5520 34777
rect 5440 34457 5520 34743
rect 5440 34423 5463 34457
rect 5497 34423 5520 34457
rect 5440 34400 5520 34423
rect 5600 36377 5680 36400
rect 5600 36343 5623 36377
rect 5657 36343 5680 36377
rect 5600 36057 5680 36343
rect 5600 36023 5623 36057
rect 5657 36023 5680 36057
rect 5600 35737 5680 36023
rect 5600 35703 5623 35737
rect 5657 35703 5680 35737
rect 5600 35417 5680 35703
rect 5600 35383 5623 35417
rect 5657 35383 5680 35417
rect 5600 35097 5680 35383
rect 5600 35063 5623 35097
rect 5657 35063 5680 35097
rect 5600 34777 5680 35063
rect 5600 34743 5623 34777
rect 5657 34743 5680 34777
rect 5600 34457 5680 34743
rect 5600 34423 5623 34457
rect 5657 34423 5680 34457
rect 5600 34400 5680 34423
rect 5760 36377 5840 36400
rect 5760 36343 5783 36377
rect 5817 36343 5840 36377
rect 5760 36057 5840 36343
rect 5760 36023 5783 36057
rect 5817 36023 5840 36057
rect 5760 35737 5840 36023
rect 5760 35703 5783 35737
rect 5817 35703 5840 35737
rect 5760 35417 5840 35703
rect 5760 35383 5783 35417
rect 5817 35383 5840 35417
rect 5760 35097 5840 35383
rect 5760 35063 5783 35097
rect 5817 35063 5840 35097
rect 5760 34777 5840 35063
rect 5760 34743 5783 34777
rect 5817 34743 5840 34777
rect 5760 34457 5840 34743
rect 5760 34423 5783 34457
rect 5817 34423 5840 34457
rect 5760 34400 5840 34423
rect 5920 36377 6000 36400
rect 5920 36343 5943 36377
rect 5977 36343 6000 36377
rect 5920 36057 6000 36343
rect 5920 36023 5943 36057
rect 5977 36023 6000 36057
rect 5920 35737 6000 36023
rect 5920 35703 5943 35737
rect 5977 35703 6000 35737
rect 5920 35417 6000 35703
rect 5920 35383 5943 35417
rect 5977 35383 6000 35417
rect 5920 35097 6000 35383
rect 5920 35063 5943 35097
rect 5977 35063 6000 35097
rect 5920 34777 6000 35063
rect 5920 34743 5943 34777
rect 5977 34743 6000 34777
rect 5920 34457 6000 34743
rect 5920 34423 5943 34457
rect 5977 34423 6000 34457
rect 5920 34400 6000 34423
rect 6080 36377 6160 36400
rect 6080 36343 6103 36377
rect 6137 36343 6160 36377
rect 6080 36057 6160 36343
rect 6080 36023 6103 36057
rect 6137 36023 6160 36057
rect 6080 35737 6160 36023
rect 6080 35703 6103 35737
rect 6137 35703 6160 35737
rect 6080 35417 6160 35703
rect 6080 35383 6103 35417
rect 6137 35383 6160 35417
rect 6080 35097 6160 35383
rect 6080 35063 6103 35097
rect 6137 35063 6160 35097
rect 6080 34777 6160 35063
rect 6080 34743 6103 34777
rect 6137 34743 6160 34777
rect 6080 34457 6160 34743
rect 6080 34423 6103 34457
rect 6137 34423 6160 34457
rect 6080 34400 6160 34423
rect 6240 36377 6320 36400
rect 6240 36343 6263 36377
rect 6297 36343 6320 36377
rect 6240 36057 6320 36343
rect 6240 36023 6263 36057
rect 6297 36023 6320 36057
rect 6240 35737 6320 36023
rect 6240 35703 6263 35737
rect 6297 35703 6320 35737
rect 6240 35417 6320 35703
rect 6240 35383 6263 35417
rect 6297 35383 6320 35417
rect 6240 35097 6320 35383
rect 6240 35063 6263 35097
rect 6297 35063 6320 35097
rect 6240 34777 6320 35063
rect 6240 34743 6263 34777
rect 6297 34743 6320 34777
rect 6240 34457 6320 34743
rect 6240 34423 6263 34457
rect 6297 34423 6320 34457
rect 6240 34400 6320 34423
rect 6400 36377 6480 36400
rect 6400 36343 6423 36377
rect 6457 36343 6480 36377
rect 6400 36057 6480 36343
rect 6400 36023 6423 36057
rect 6457 36023 6480 36057
rect 6400 35737 6480 36023
rect 6400 35703 6423 35737
rect 6457 35703 6480 35737
rect 6400 35417 6480 35703
rect 6400 35383 6423 35417
rect 6457 35383 6480 35417
rect 6400 35097 6480 35383
rect 6400 35063 6423 35097
rect 6457 35063 6480 35097
rect 6400 34777 6480 35063
rect 6400 34743 6423 34777
rect 6457 34743 6480 34777
rect 6400 34457 6480 34743
rect 6400 34423 6423 34457
rect 6457 34423 6480 34457
rect 6400 34400 6480 34423
rect 6560 36377 6640 36400
rect 6560 36343 6583 36377
rect 6617 36343 6640 36377
rect 6560 36057 6640 36343
rect 6560 36023 6583 36057
rect 6617 36023 6640 36057
rect 6560 35737 6640 36023
rect 6560 35703 6583 35737
rect 6617 35703 6640 35737
rect 6560 35417 6640 35703
rect 6560 35383 6583 35417
rect 6617 35383 6640 35417
rect 6560 35097 6640 35383
rect 6560 35063 6583 35097
rect 6617 35063 6640 35097
rect 6560 34777 6640 35063
rect 6560 34743 6583 34777
rect 6617 34743 6640 34777
rect 6560 34457 6640 34743
rect 6560 34423 6583 34457
rect 6617 34423 6640 34457
rect 6560 34400 6640 34423
rect 6720 36377 6800 36400
rect 6720 36343 6743 36377
rect 6777 36343 6800 36377
rect 6720 36057 6800 36343
rect 6720 36023 6743 36057
rect 6777 36023 6800 36057
rect 6720 35737 6800 36023
rect 6720 35703 6743 35737
rect 6777 35703 6800 35737
rect 6720 35417 6800 35703
rect 6720 35383 6743 35417
rect 6777 35383 6800 35417
rect 6720 35097 6800 35383
rect 6720 35063 6743 35097
rect 6777 35063 6800 35097
rect 6720 34777 6800 35063
rect 6720 34743 6743 34777
rect 6777 34743 6800 34777
rect 6720 34457 6800 34743
rect 6720 34423 6743 34457
rect 6777 34423 6800 34457
rect 6720 34400 6800 34423
rect 6880 36377 6960 36400
rect 6880 36343 6903 36377
rect 6937 36343 6960 36377
rect 6880 36057 6960 36343
rect 6880 36023 6903 36057
rect 6937 36023 6960 36057
rect 6880 35737 6960 36023
rect 6880 35703 6903 35737
rect 6937 35703 6960 35737
rect 6880 35417 6960 35703
rect 6880 35383 6903 35417
rect 6937 35383 6960 35417
rect 6880 35097 6960 35383
rect 6880 35063 6903 35097
rect 6937 35063 6960 35097
rect 6880 34777 6960 35063
rect 6880 34743 6903 34777
rect 6937 34743 6960 34777
rect 6880 34457 6960 34743
rect 6880 34423 6903 34457
rect 6937 34423 6960 34457
rect 6880 34400 6960 34423
rect 7040 36377 7120 36400
rect 7040 36343 7063 36377
rect 7097 36343 7120 36377
rect 7040 36057 7120 36343
rect 7040 36023 7063 36057
rect 7097 36023 7120 36057
rect 7040 35737 7120 36023
rect 7040 35703 7063 35737
rect 7097 35703 7120 35737
rect 7040 35417 7120 35703
rect 7040 35383 7063 35417
rect 7097 35383 7120 35417
rect 7040 35097 7120 35383
rect 7040 35063 7063 35097
rect 7097 35063 7120 35097
rect 7040 34777 7120 35063
rect 7040 34743 7063 34777
rect 7097 34743 7120 34777
rect 7040 34457 7120 34743
rect 7040 34423 7063 34457
rect 7097 34423 7120 34457
rect 7040 34400 7120 34423
rect 7200 36377 7280 36400
rect 7200 36343 7223 36377
rect 7257 36343 7280 36377
rect 7200 36057 7280 36343
rect 7200 36023 7223 36057
rect 7257 36023 7280 36057
rect 7200 35737 7280 36023
rect 7200 35703 7223 35737
rect 7257 35703 7280 35737
rect 7200 35417 7280 35703
rect 7200 35383 7223 35417
rect 7257 35383 7280 35417
rect 7200 35097 7280 35383
rect 7200 35063 7223 35097
rect 7257 35063 7280 35097
rect 7200 34777 7280 35063
rect 7200 34743 7223 34777
rect 7257 34743 7280 34777
rect 7200 34457 7280 34743
rect 7200 34423 7223 34457
rect 7257 34423 7280 34457
rect 7200 34400 7280 34423
rect 7360 36377 7440 36400
rect 7360 36343 7383 36377
rect 7417 36343 7440 36377
rect 7360 36057 7440 36343
rect 7360 36023 7383 36057
rect 7417 36023 7440 36057
rect 7360 35737 7440 36023
rect 7360 35703 7383 35737
rect 7417 35703 7440 35737
rect 7360 35417 7440 35703
rect 7360 35383 7383 35417
rect 7417 35383 7440 35417
rect 7360 35097 7440 35383
rect 7360 35063 7383 35097
rect 7417 35063 7440 35097
rect 7360 34777 7440 35063
rect 7360 34743 7383 34777
rect 7417 34743 7440 34777
rect 7360 34457 7440 34743
rect 7360 34423 7383 34457
rect 7417 34423 7440 34457
rect 7360 34400 7440 34423
rect 7520 36377 7600 36400
rect 7520 36343 7543 36377
rect 7577 36343 7600 36377
rect 7520 36057 7600 36343
rect 7520 36023 7543 36057
rect 7577 36023 7600 36057
rect 7520 35737 7600 36023
rect 7520 35703 7543 35737
rect 7577 35703 7600 35737
rect 7520 35417 7600 35703
rect 7520 35383 7543 35417
rect 7577 35383 7600 35417
rect 7520 35097 7600 35383
rect 7520 35063 7543 35097
rect 7577 35063 7600 35097
rect 7520 34777 7600 35063
rect 7520 34743 7543 34777
rect 7577 34743 7600 34777
rect 7520 34457 7600 34743
rect 7520 34423 7543 34457
rect 7577 34423 7600 34457
rect 7520 34400 7600 34423
rect 7680 36377 7760 36400
rect 7680 36343 7703 36377
rect 7737 36343 7760 36377
rect 7680 36057 7760 36343
rect 7680 36023 7703 36057
rect 7737 36023 7760 36057
rect 7680 35737 7760 36023
rect 7680 35703 7703 35737
rect 7737 35703 7760 35737
rect 7680 35417 7760 35703
rect 7680 35383 7703 35417
rect 7737 35383 7760 35417
rect 7680 35097 7760 35383
rect 7680 35063 7703 35097
rect 7737 35063 7760 35097
rect 7680 34777 7760 35063
rect 7680 34743 7703 34777
rect 7737 34743 7760 34777
rect 7680 34457 7760 34743
rect 7680 34423 7703 34457
rect 7737 34423 7760 34457
rect 7680 34400 7760 34423
rect 7840 36377 7920 36400
rect 7840 36343 7863 36377
rect 7897 36343 7920 36377
rect 7840 36057 7920 36343
rect 7840 36023 7863 36057
rect 7897 36023 7920 36057
rect 7840 35737 7920 36023
rect 7840 35703 7863 35737
rect 7897 35703 7920 35737
rect 7840 35417 7920 35703
rect 7840 35383 7863 35417
rect 7897 35383 7920 35417
rect 7840 35097 7920 35383
rect 7840 35063 7863 35097
rect 7897 35063 7920 35097
rect 7840 34777 7920 35063
rect 7840 34743 7863 34777
rect 7897 34743 7920 34777
rect 7840 34457 7920 34743
rect 7840 34423 7863 34457
rect 7897 34423 7920 34457
rect 7840 34400 7920 34423
rect 8000 36377 8080 36400
rect 8000 36343 8023 36377
rect 8057 36343 8080 36377
rect 8000 36057 8080 36343
rect 8000 36023 8023 36057
rect 8057 36023 8080 36057
rect 8000 35737 8080 36023
rect 8000 35703 8023 35737
rect 8057 35703 8080 35737
rect 8000 35417 8080 35703
rect 8000 35383 8023 35417
rect 8057 35383 8080 35417
rect 8000 35097 8080 35383
rect 8000 35063 8023 35097
rect 8057 35063 8080 35097
rect 8000 34777 8080 35063
rect 8000 34743 8023 34777
rect 8057 34743 8080 34777
rect 8000 34457 8080 34743
rect 8000 34423 8023 34457
rect 8057 34423 8080 34457
rect 8000 34400 8080 34423
rect 8160 36377 8240 36400
rect 8160 36343 8183 36377
rect 8217 36343 8240 36377
rect 8160 36057 8240 36343
rect 8160 36023 8183 36057
rect 8217 36023 8240 36057
rect 8160 35737 8240 36023
rect 8160 35703 8183 35737
rect 8217 35703 8240 35737
rect 8160 35417 8240 35703
rect 8160 35383 8183 35417
rect 8217 35383 8240 35417
rect 8160 35097 8240 35383
rect 8160 35063 8183 35097
rect 8217 35063 8240 35097
rect 8160 34777 8240 35063
rect 8160 34743 8183 34777
rect 8217 34743 8240 34777
rect 8160 34457 8240 34743
rect 8160 34423 8183 34457
rect 8217 34423 8240 34457
rect 8160 34400 8240 34423
rect 8320 36377 8400 36400
rect 8320 36343 8343 36377
rect 8377 36343 8400 36377
rect 8320 36057 8400 36343
rect 8320 36023 8343 36057
rect 8377 36023 8400 36057
rect 8320 35737 8400 36023
rect 8320 35703 8343 35737
rect 8377 35703 8400 35737
rect 8320 35417 8400 35703
rect 8320 35383 8343 35417
rect 8377 35383 8400 35417
rect 8320 35097 8400 35383
rect 8320 35063 8343 35097
rect 8377 35063 8400 35097
rect 8320 34777 8400 35063
rect 8320 34743 8343 34777
rect 8377 34743 8400 34777
rect 8320 34457 8400 34743
rect 8320 34423 8343 34457
rect 8377 34423 8400 34457
rect 8320 34400 8400 34423
rect 8480 34400 8560 36400
rect 8640 34400 8720 36400
rect 8800 34400 8880 36400
rect 8960 34400 9040 36400
rect 9120 34400 9200 36400
rect 9280 34400 9360 36400
rect 9440 34400 9520 36400
rect 9600 34400 9680 36400
rect 9760 34400 9840 36400
rect 9920 34400 10000 36400
rect 10080 34400 10160 36400
rect 10240 34400 10320 36400
rect 10400 34400 10480 36400
rect 10560 34400 10640 36400
rect 10720 34400 10800 36400
rect 10880 34400 10960 36400
rect 11040 34400 11120 36400
rect 11200 34400 11280 36400
rect 11360 34400 11440 36400
rect 11520 34400 11600 36400
rect 11680 34400 11760 36400
rect 11840 34400 11920 36400
rect 12000 34400 12080 36400
rect 12160 34400 12240 36400
rect 12320 34400 12400 36400
rect 12480 36377 12560 36400
rect 12480 36343 12503 36377
rect 12537 36343 12560 36377
rect 12480 36057 12560 36343
rect 12480 36023 12503 36057
rect 12537 36023 12560 36057
rect 12480 35737 12560 36023
rect 12480 35703 12503 35737
rect 12537 35703 12560 35737
rect 12480 35417 12560 35703
rect 12480 35383 12503 35417
rect 12537 35383 12560 35417
rect 12480 35097 12560 35383
rect 12480 35063 12503 35097
rect 12537 35063 12560 35097
rect 12480 34777 12560 35063
rect 12480 34743 12503 34777
rect 12537 34743 12560 34777
rect 12480 34457 12560 34743
rect 12480 34423 12503 34457
rect 12537 34423 12560 34457
rect 12480 34400 12560 34423
rect 12640 36377 12720 36400
rect 12640 36343 12663 36377
rect 12697 36343 12720 36377
rect 12640 36057 12720 36343
rect 12640 36023 12663 36057
rect 12697 36023 12720 36057
rect 12640 35737 12720 36023
rect 12640 35703 12663 35737
rect 12697 35703 12720 35737
rect 12640 35417 12720 35703
rect 12640 35383 12663 35417
rect 12697 35383 12720 35417
rect 12640 35097 12720 35383
rect 12640 35063 12663 35097
rect 12697 35063 12720 35097
rect 12640 34777 12720 35063
rect 12640 34743 12663 34777
rect 12697 34743 12720 34777
rect 12640 34457 12720 34743
rect 12640 34423 12663 34457
rect 12697 34423 12720 34457
rect 12640 34400 12720 34423
rect 12800 36377 12880 36400
rect 12800 36343 12823 36377
rect 12857 36343 12880 36377
rect 12800 36057 12880 36343
rect 12800 36023 12823 36057
rect 12857 36023 12880 36057
rect 12800 35737 12880 36023
rect 12800 35703 12823 35737
rect 12857 35703 12880 35737
rect 12800 35417 12880 35703
rect 12800 35383 12823 35417
rect 12857 35383 12880 35417
rect 12800 35097 12880 35383
rect 12800 35063 12823 35097
rect 12857 35063 12880 35097
rect 12800 34777 12880 35063
rect 12800 34743 12823 34777
rect 12857 34743 12880 34777
rect 12800 34457 12880 34743
rect 12800 34423 12823 34457
rect 12857 34423 12880 34457
rect 12800 34400 12880 34423
rect 12960 36377 13040 36400
rect 12960 36343 12983 36377
rect 13017 36343 13040 36377
rect 12960 36057 13040 36343
rect 12960 36023 12983 36057
rect 13017 36023 13040 36057
rect 12960 35737 13040 36023
rect 12960 35703 12983 35737
rect 13017 35703 13040 35737
rect 12960 35417 13040 35703
rect 12960 35383 12983 35417
rect 13017 35383 13040 35417
rect 12960 35097 13040 35383
rect 12960 35063 12983 35097
rect 13017 35063 13040 35097
rect 12960 34777 13040 35063
rect 12960 34743 12983 34777
rect 13017 34743 13040 34777
rect 12960 34457 13040 34743
rect 12960 34423 12983 34457
rect 13017 34423 13040 34457
rect 12960 34400 13040 34423
rect 13120 36377 13200 36400
rect 13120 36343 13143 36377
rect 13177 36343 13200 36377
rect 13120 36057 13200 36343
rect 13120 36023 13143 36057
rect 13177 36023 13200 36057
rect 13120 35737 13200 36023
rect 13120 35703 13143 35737
rect 13177 35703 13200 35737
rect 13120 35417 13200 35703
rect 13120 35383 13143 35417
rect 13177 35383 13200 35417
rect 13120 35097 13200 35383
rect 13120 35063 13143 35097
rect 13177 35063 13200 35097
rect 13120 34777 13200 35063
rect 13120 34743 13143 34777
rect 13177 34743 13200 34777
rect 13120 34457 13200 34743
rect 13120 34423 13143 34457
rect 13177 34423 13200 34457
rect 13120 34400 13200 34423
rect 13280 36377 13360 36400
rect 13280 36343 13303 36377
rect 13337 36343 13360 36377
rect 13280 36057 13360 36343
rect 13280 36023 13303 36057
rect 13337 36023 13360 36057
rect 13280 35737 13360 36023
rect 13280 35703 13303 35737
rect 13337 35703 13360 35737
rect 13280 35417 13360 35703
rect 13280 35383 13303 35417
rect 13337 35383 13360 35417
rect 13280 35097 13360 35383
rect 13280 35063 13303 35097
rect 13337 35063 13360 35097
rect 13280 34777 13360 35063
rect 13280 34743 13303 34777
rect 13337 34743 13360 34777
rect 13280 34457 13360 34743
rect 13280 34423 13303 34457
rect 13337 34423 13360 34457
rect 13280 34400 13360 34423
rect 13440 36377 13520 36400
rect 13440 36343 13463 36377
rect 13497 36343 13520 36377
rect 13440 36057 13520 36343
rect 13440 36023 13463 36057
rect 13497 36023 13520 36057
rect 13440 35737 13520 36023
rect 13440 35703 13463 35737
rect 13497 35703 13520 35737
rect 13440 35417 13520 35703
rect 13440 35383 13463 35417
rect 13497 35383 13520 35417
rect 13440 35097 13520 35383
rect 13440 35063 13463 35097
rect 13497 35063 13520 35097
rect 13440 34777 13520 35063
rect 13440 34743 13463 34777
rect 13497 34743 13520 34777
rect 13440 34457 13520 34743
rect 13440 34423 13463 34457
rect 13497 34423 13520 34457
rect 13440 34400 13520 34423
rect 13600 36377 13680 36400
rect 13600 36343 13623 36377
rect 13657 36343 13680 36377
rect 13600 36057 13680 36343
rect 13600 36023 13623 36057
rect 13657 36023 13680 36057
rect 13600 35737 13680 36023
rect 13600 35703 13623 35737
rect 13657 35703 13680 35737
rect 13600 35417 13680 35703
rect 13600 35383 13623 35417
rect 13657 35383 13680 35417
rect 13600 35097 13680 35383
rect 13600 35063 13623 35097
rect 13657 35063 13680 35097
rect 13600 34777 13680 35063
rect 13600 34743 13623 34777
rect 13657 34743 13680 34777
rect 13600 34457 13680 34743
rect 13600 34423 13623 34457
rect 13657 34423 13680 34457
rect 13600 34400 13680 34423
rect 13760 36377 13840 36400
rect 13760 36343 13783 36377
rect 13817 36343 13840 36377
rect 13760 36057 13840 36343
rect 13760 36023 13783 36057
rect 13817 36023 13840 36057
rect 13760 35737 13840 36023
rect 13760 35703 13783 35737
rect 13817 35703 13840 35737
rect 13760 35417 13840 35703
rect 13760 35383 13783 35417
rect 13817 35383 13840 35417
rect 13760 35097 13840 35383
rect 13760 35063 13783 35097
rect 13817 35063 13840 35097
rect 13760 34777 13840 35063
rect 13760 34743 13783 34777
rect 13817 34743 13840 34777
rect 13760 34457 13840 34743
rect 13760 34423 13783 34457
rect 13817 34423 13840 34457
rect 13760 34400 13840 34423
rect 13920 36377 14000 36400
rect 13920 36343 13943 36377
rect 13977 36343 14000 36377
rect 13920 36057 14000 36343
rect 13920 36023 13943 36057
rect 13977 36023 14000 36057
rect 13920 35737 14000 36023
rect 13920 35703 13943 35737
rect 13977 35703 14000 35737
rect 13920 35417 14000 35703
rect 13920 35383 13943 35417
rect 13977 35383 14000 35417
rect 13920 35097 14000 35383
rect 13920 35063 13943 35097
rect 13977 35063 14000 35097
rect 13920 34777 14000 35063
rect 13920 34743 13943 34777
rect 13977 34743 14000 34777
rect 13920 34457 14000 34743
rect 13920 34423 13943 34457
rect 13977 34423 14000 34457
rect 13920 34400 14000 34423
rect 14080 36377 14160 36400
rect 14080 36343 14103 36377
rect 14137 36343 14160 36377
rect 14080 36057 14160 36343
rect 14080 36023 14103 36057
rect 14137 36023 14160 36057
rect 14080 35737 14160 36023
rect 14080 35703 14103 35737
rect 14137 35703 14160 35737
rect 14080 35417 14160 35703
rect 14080 35383 14103 35417
rect 14137 35383 14160 35417
rect 14080 35097 14160 35383
rect 14080 35063 14103 35097
rect 14137 35063 14160 35097
rect 14080 34777 14160 35063
rect 14080 34743 14103 34777
rect 14137 34743 14160 34777
rect 14080 34457 14160 34743
rect 14080 34423 14103 34457
rect 14137 34423 14160 34457
rect 14080 34400 14160 34423
rect 14240 36377 14320 36400
rect 14240 36343 14263 36377
rect 14297 36343 14320 36377
rect 14240 36057 14320 36343
rect 14240 36023 14263 36057
rect 14297 36023 14320 36057
rect 14240 35737 14320 36023
rect 14240 35703 14263 35737
rect 14297 35703 14320 35737
rect 14240 35417 14320 35703
rect 14240 35383 14263 35417
rect 14297 35383 14320 35417
rect 14240 35097 14320 35383
rect 14240 35063 14263 35097
rect 14297 35063 14320 35097
rect 14240 34777 14320 35063
rect 14240 34743 14263 34777
rect 14297 34743 14320 34777
rect 14240 34457 14320 34743
rect 14240 34423 14263 34457
rect 14297 34423 14320 34457
rect 14240 34400 14320 34423
rect 14400 36377 14480 36400
rect 14400 36343 14423 36377
rect 14457 36343 14480 36377
rect 14400 36057 14480 36343
rect 14400 36023 14423 36057
rect 14457 36023 14480 36057
rect 14400 35737 14480 36023
rect 14400 35703 14423 35737
rect 14457 35703 14480 35737
rect 14400 35417 14480 35703
rect 14400 35383 14423 35417
rect 14457 35383 14480 35417
rect 14400 35097 14480 35383
rect 14400 35063 14423 35097
rect 14457 35063 14480 35097
rect 14400 34777 14480 35063
rect 14400 34743 14423 34777
rect 14457 34743 14480 34777
rect 14400 34457 14480 34743
rect 14400 34423 14423 34457
rect 14457 34423 14480 34457
rect 14400 34400 14480 34423
rect 14560 36377 14640 36400
rect 14560 36343 14583 36377
rect 14617 36343 14640 36377
rect 14560 36057 14640 36343
rect 14560 36023 14583 36057
rect 14617 36023 14640 36057
rect 14560 35737 14640 36023
rect 14560 35703 14583 35737
rect 14617 35703 14640 35737
rect 14560 35417 14640 35703
rect 14560 35383 14583 35417
rect 14617 35383 14640 35417
rect 14560 35097 14640 35383
rect 14560 35063 14583 35097
rect 14617 35063 14640 35097
rect 14560 34777 14640 35063
rect 14560 34743 14583 34777
rect 14617 34743 14640 34777
rect 14560 34457 14640 34743
rect 14560 34423 14583 34457
rect 14617 34423 14640 34457
rect 14560 34400 14640 34423
rect 14720 36377 14800 36400
rect 14720 36343 14743 36377
rect 14777 36343 14800 36377
rect 14720 36057 14800 36343
rect 14720 36023 14743 36057
rect 14777 36023 14800 36057
rect 14720 35737 14800 36023
rect 14720 35703 14743 35737
rect 14777 35703 14800 35737
rect 14720 35417 14800 35703
rect 14720 35383 14743 35417
rect 14777 35383 14800 35417
rect 14720 35097 14800 35383
rect 14720 35063 14743 35097
rect 14777 35063 14800 35097
rect 14720 34777 14800 35063
rect 14720 34743 14743 34777
rect 14777 34743 14800 34777
rect 14720 34457 14800 34743
rect 14720 34423 14743 34457
rect 14777 34423 14800 34457
rect 14720 34400 14800 34423
rect 14880 36377 14960 36400
rect 14880 36343 14903 36377
rect 14937 36343 14960 36377
rect 14880 36057 14960 36343
rect 14880 36023 14903 36057
rect 14937 36023 14960 36057
rect 14880 35737 14960 36023
rect 14880 35703 14903 35737
rect 14937 35703 14960 35737
rect 14880 35417 14960 35703
rect 14880 35383 14903 35417
rect 14937 35383 14960 35417
rect 14880 35097 14960 35383
rect 14880 35063 14903 35097
rect 14937 35063 14960 35097
rect 14880 34777 14960 35063
rect 14880 34743 14903 34777
rect 14937 34743 14960 34777
rect 14880 34457 14960 34743
rect 14880 34423 14903 34457
rect 14937 34423 14960 34457
rect 14880 34400 14960 34423
rect 15040 36377 15120 36400
rect 15040 36343 15063 36377
rect 15097 36343 15120 36377
rect 15040 36057 15120 36343
rect 15040 36023 15063 36057
rect 15097 36023 15120 36057
rect 15040 35737 15120 36023
rect 15040 35703 15063 35737
rect 15097 35703 15120 35737
rect 15040 35417 15120 35703
rect 15040 35383 15063 35417
rect 15097 35383 15120 35417
rect 15040 35097 15120 35383
rect 15040 35063 15063 35097
rect 15097 35063 15120 35097
rect 15040 34777 15120 35063
rect 15040 34743 15063 34777
rect 15097 34743 15120 34777
rect 15040 34457 15120 34743
rect 15040 34423 15063 34457
rect 15097 34423 15120 34457
rect 15040 34400 15120 34423
rect 15200 36377 15280 36400
rect 15200 36343 15223 36377
rect 15257 36343 15280 36377
rect 15200 36057 15280 36343
rect 15200 36023 15223 36057
rect 15257 36023 15280 36057
rect 15200 35737 15280 36023
rect 15200 35703 15223 35737
rect 15257 35703 15280 35737
rect 15200 35417 15280 35703
rect 15200 35383 15223 35417
rect 15257 35383 15280 35417
rect 15200 35097 15280 35383
rect 15200 35063 15223 35097
rect 15257 35063 15280 35097
rect 15200 34777 15280 35063
rect 15200 34743 15223 34777
rect 15257 34743 15280 34777
rect 15200 34457 15280 34743
rect 15200 34423 15223 34457
rect 15257 34423 15280 34457
rect 15200 34400 15280 34423
rect 15360 36377 15440 36400
rect 15360 36343 15383 36377
rect 15417 36343 15440 36377
rect 15360 36057 15440 36343
rect 15360 36023 15383 36057
rect 15417 36023 15440 36057
rect 15360 35737 15440 36023
rect 15360 35703 15383 35737
rect 15417 35703 15440 35737
rect 15360 35417 15440 35703
rect 15360 35383 15383 35417
rect 15417 35383 15440 35417
rect 15360 35097 15440 35383
rect 15360 35063 15383 35097
rect 15417 35063 15440 35097
rect 15360 34777 15440 35063
rect 15360 34743 15383 34777
rect 15417 34743 15440 34777
rect 15360 34457 15440 34743
rect 15360 34423 15383 34457
rect 15417 34423 15440 34457
rect 15360 34400 15440 34423
rect 15520 36377 15600 36400
rect 15520 36343 15543 36377
rect 15577 36343 15600 36377
rect 15520 36057 15600 36343
rect 15520 36023 15543 36057
rect 15577 36023 15600 36057
rect 15520 35737 15600 36023
rect 15520 35703 15543 35737
rect 15577 35703 15600 35737
rect 15520 35417 15600 35703
rect 15520 35383 15543 35417
rect 15577 35383 15600 35417
rect 15520 35097 15600 35383
rect 15520 35063 15543 35097
rect 15577 35063 15600 35097
rect 15520 34777 15600 35063
rect 15520 34743 15543 34777
rect 15577 34743 15600 34777
rect 15520 34457 15600 34743
rect 15520 34423 15543 34457
rect 15577 34423 15600 34457
rect 15520 34400 15600 34423
rect 15680 36377 15760 36400
rect 15680 36343 15703 36377
rect 15737 36343 15760 36377
rect 15680 36057 15760 36343
rect 15680 36023 15703 36057
rect 15737 36023 15760 36057
rect 15680 35737 15760 36023
rect 15680 35703 15703 35737
rect 15737 35703 15760 35737
rect 15680 35417 15760 35703
rect 15680 35383 15703 35417
rect 15737 35383 15760 35417
rect 15680 35097 15760 35383
rect 15680 35063 15703 35097
rect 15737 35063 15760 35097
rect 15680 34777 15760 35063
rect 15680 34743 15703 34777
rect 15737 34743 15760 34777
rect 15680 34457 15760 34743
rect 15680 34423 15703 34457
rect 15737 34423 15760 34457
rect 15680 34400 15760 34423
rect 15840 36377 15920 36400
rect 15840 36343 15863 36377
rect 15897 36343 15920 36377
rect 15840 36057 15920 36343
rect 15840 36023 15863 36057
rect 15897 36023 15920 36057
rect 15840 35737 15920 36023
rect 15840 35703 15863 35737
rect 15897 35703 15920 35737
rect 15840 35417 15920 35703
rect 15840 35383 15863 35417
rect 15897 35383 15920 35417
rect 15840 35097 15920 35383
rect 15840 35063 15863 35097
rect 15897 35063 15920 35097
rect 15840 34777 15920 35063
rect 15840 34743 15863 34777
rect 15897 34743 15920 34777
rect 15840 34457 15920 34743
rect 15840 34423 15863 34457
rect 15897 34423 15920 34457
rect 15840 34400 15920 34423
rect 16000 36377 16080 36400
rect 16000 36343 16023 36377
rect 16057 36343 16080 36377
rect 16000 36057 16080 36343
rect 16000 36023 16023 36057
rect 16057 36023 16080 36057
rect 16000 35737 16080 36023
rect 16000 35703 16023 35737
rect 16057 35703 16080 35737
rect 16000 35417 16080 35703
rect 16000 35383 16023 35417
rect 16057 35383 16080 35417
rect 16000 35097 16080 35383
rect 16000 35063 16023 35097
rect 16057 35063 16080 35097
rect 16000 34777 16080 35063
rect 16000 34743 16023 34777
rect 16057 34743 16080 34777
rect 16000 34457 16080 34743
rect 16000 34423 16023 34457
rect 16057 34423 16080 34457
rect 16000 34400 16080 34423
rect 16160 36377 16240 36400
rect 16160 36343 16183 36377
rect 16217 36343 16240 36377
rect 16160 36057 16240 36343
rect 16160 36023 16183 36057
rect 16217 36023 16240 36057
rect 16160 35737 16240 36023
rect 16160 35703 16183 35737
rect 16217 35703 16240 35737
rect 16160 35417 16240 35703
rect 16160 35383 16183 35417
rect 16217 35383 16240 35417
rect 16160 35097 16240 35383
rect 16160 35063 16183 35097
rect 16217 35063 16240 35097
rect 16160 34777 16240 35063
rect 16160 34743 16183 34777
rect 16217 34743 16240 34777
rect 16160 34457 16240 34743
rect 16160 34423 16183 34457
rect 16217 34423 16240 34457
rect 16160 34400 16240 34423
rect 16320 36377 16400 36400
rect 16320 36343 16343 36377
rect 16377 36343 16400 36377
rect 16320 36057 16400 36343
rect 16320 36023 16343 36057
rect 16377 36023 16400 36057
rect 16320 35737 16400 36023
rect 16320 35703 16343 35737
rect 16377 35703 16400 35737
rect 16320 35417 16400 35703
rect 16320 35383 16343 35417
rect 16377 35383 16400 35417
rect 16320 35097 16400 35383
rect 16320 35063 16343 35097
rect 16377 35063 16400 35097
rect 16320 34777 16400 35063
rect 16320 34743 16343 34777
rect 16377 34743 16400 34777
rect 16320 34457 16400 34743
rect 16320 34423 16343 34457
rect 16377 34423 16400 34457
rect 16320 34400 16400 34423
rect 16480 36377 16560 36400
rect 16480 36343 16503 36377
rect 16537 36343 16560 36377
rect 16480 36057 16560 36343
rect 16480 36023 16503 36057
rect 16537 36023 16560 36057
rect 16480 35737 16560 36023
rect 16480 35703 16503 35737
rect 16537 35703 16560 35737
rect 16480 35417 16560 35703
rect 16480 35383 16503 35417
rect 16537 35383 16560 35417
rect 16480 35097 16560 35383
rect 16480 35063 16503 35097
rect 16537 35063 16560 35097
rect 16480 34777 16560 35063
rect 16480 34743 16503 34777
rect 16537 34743 16560 34777
rect 16480 34457 16560 34743
rect 16480 34423 16503 34457
rect 16537 34423 16560 34457
rect 16480 34400 16560 34423
rect 16640 36377 16720 36400
rect 16640 36343 16663 36377
rect 16697 36343 16720 36377
rect 16640 36057 16720 36343
rect 16640 36023 16663 36057
rect 16697 36023 16720 36057
rect 16640 35737 16720 36023
rect 16640 35703 16663 35737
rect 16697 35703 16720 35737
rect 16640 35417 16720 35703
rect 16640 35383 16663 35417
rect 16697 35383 16720 35417
rect 16640 35097 16720 35383
rect 16640 35063 16663 35097
rect 16697 35063 16720 35097
rect 16640 34777 16720 35063
rect 16640 34743 16663 34777
rect 16697 34743 16720 34777
rect 16640 34457 16720 34743
rect 16640 34423 16663 34457
rect 16697 34423 16720 34457
rect 16640 34400 16720 34423
rect 16800 36377 16880 36400
rect 16800 36343 16823 36377
rect 16857 36343 16880 36377
rect 16800 36057 16880 36343
rect 16800 36023 16823 36057
rect 16857 36023 16880 36057
rect 16800 35737 16880 36023
rect 16800 35703 16823 35737
rect 16857 35703 16880 35737
rect 16800 35417 16880 35703
rect 16800 35383 16823 35417
rect 16857 35383 16880 35417
rect 16800 35097 16880 35383
rect 16800 35063 16823 35097
rect 16857 35063 16880 35097
rect 16800 34777 16880 35063
rect 16800 34743 16823 34777
rect 16857 34743 16880 34777
rect 16800 34457 16880 34743
rect 16800 34423 16823 34457
rect 16857 34423 16880 34457
rect 16800 34400 16880 34423
rect 16960 36377 17040 36400
rect 16960 36343 16983 36377
rect 17017 36343 17040 36377
rect 16960 36057 17040 36343
rect 16960 36023 16983 36057
rect 17017 36023 17040 36057
rect 16960 35737 17040 36023
rect 16960 35703 16983 35737
rect 17017 35703 17040 35737
rect 16960 35417 17040 35703
rect 16960 35383 16983 35417
rect 17017 35383 17040 35417
rect 16960 35097 17040 35383
rect 16960 35063 16983 35097
rect 17017 35063 17040 35097
rect 16960 34777 17040 35063
rect 16960 34743 16983 34777
rect 17017 34743 17040 34777
rect 16960 34457 17040 34743
rect 16960 34423 16983 34457
rect 17017 34423 17040 34457
rect 16960 34400 17040 34423
rect 17120 36377 17200 36400
rect 17120 36343 17143 36377
rect 17177 36343 17200 36377
rect 17120 36057 17200 36343
rect 17120 36023 17143 36057
rect 17177 36023 17200 36057
rect 17120 35737 17200 36023
rect 17120 35703 17143 35737
rect 17177 35703 17200 35737
rect 17120 35417 17200 35703
rect 17120 35383 17143 35417
rect 17177 35383 17200 35417
rect 17120 35097 17200 35383
rect 17120 35063 17143 35097
rect 17177 35063 17200 35097
rect 17120 34777 17200 35063
rect 17120 34743 17143 34777
rect 17177 34743 17200 34777
rect 17120 34457 17200 34743
rect 17120 34423 17143 34457
rect 17177 34423 17200 34457
rect 17120 34400 17200 34423
rect 17280 36377 17360 36400
rect 17280 36343 17303 36377
rect 17337 36343 17360 36377
rect 17280 36057 17360 36343
rect 17280 36023 17303 36057
rect 17337 36023 17360 36057
rect 17280 35737 17360 36023
rect 17280 35703 17303 35737
rect 17337 35703 17360 35737
rect 17280 35417 17360 35703
rect 17280 35383 17303 35417
rect 17337 35383 17360 35417
rect 17280 35097 17360 35383
rect 17280 35063 17303 35097
rect 17337 35063 17360 35097
rect 17280 34777 17360 35063
rect 17280 34743 17303 34777
rect 17337 34743 17360 34777
rect 17280 34457 17360 34743
rect 17280 34423 17303 34457
rect 17337 34423 17360 34457
rect 17280 34400 17360 34423
rect 17440 36377 17520 36400
rect 17440 36343 17463 36377
rect 17497 36343 17520 36377
rect 17440 36057 17520 36343
rect 17440 36023 17463 36057
rect 17497 36023 17520 36057
rect 17440 35737 17520 36023
rect 17440 35703 17463 35737
rect 17497 35703 17520 35737
rect 17440 35417 17520 35703
rect 17440 35383 17463 35417
rect 17497 35383 17520 35417
rect 17440 35097 17520 35383
rect 17440 35063 17463 35097
rect 17497 35063 17520 35097
rect 17440 34777 17520 35063
rect 17440 34743 17463 34777
rect 17497 34743 17520 34777
rect 17440 34457 17520 34743
rect 17440 34423 17463 34457
rect 17497 34423 17520 34457
rect 17440 34400 17520 34423
rect 17600 36377 17680 36400
rect 17600 36343 17623 36377
rect 17657 36343 17680 36377
rect 17600 36057 17680 36343
rect 17600 36023 17623 36057
rect 17657 36023 17680 36057
rect 17600 35737 17680 36023
rect 17600 35703 17623 35737
rect 17657 35703 17680 35737
rect 17600 35417 17680 35703
rect 17600 35383 17623 35417
rect 17657 35383 17680 35417
rect 17600 35097 17680 35383
rect 17600 35063 17623 35097
rect 17657 35063 17680 35097
rect 17600 34777 17680 35063
rect 17600 34743 17623 34777
rect 17657 34743 17680 34777
rect 17600 34457 17680 34743
rect 17600 34423 17623 34457
rect 17657 34423 17680 34457
rect 17600 34400 17680 34423
rect 17760 36377 17840 36400
rect 17760 36343 17783 36377
rect 17817 36343 17840 36377
rect 17760 36057 17840 36343
rect 17760 36023 17783 36057
rect 17817 36023 17840 36057
rect 17760 35737 17840 36023
rect 17760 35703 17783 35737
rect 17817 35703 17840 35737
rect 17760 35417 17840 35703
rect 17760 35383 17783 35417
rect 17817 35383 17840 35417
rect 17760 35097 17840 35383
rect 17760 35063 17783 35097
rect 17817 35063 17840 35097
rect 17760 34777 17840 35063
rect 17760 34743 17783 34777
rect 17817 34743 17840 34777
rect 17760 34457 17840 34743
rect 17760 34423 17783 34457
rect 17817 34423 17840 34457
rect 17760 34400 17840 34423
rect 17920 36377 18000 36400
rect 17920 36343 17943 36377
rect 17977 36343 18000 36377
rect 17920 36057 18000 36343
rect 17920 36023 17943 36057
rect 17977 36023 18000 36057
rect 17920 35737 18000 36023
rect 17920 35703 17943 35737
rect 17977 35703 18000 35737
rect 17920 35417 18000 35703
rect 17920 35383 17943 35417
rect 17977 35383 18000 35417
rect 17920 35097 18000 35383
rect 17920 35063 17943 35097
rect 17977 35063 18000 35097
rect 17920 34777 18000 35063
rect 17920 34743 17943 34777
rect 17977 34743 18000 34777
rect 17920 34457 18000 34743
rect 17920 34423 17943 34457
rect 17977 34423 18000 34457
rect 17920 34400 18000 34423
rect 18080 36377 18160 36400
rect 18080 36343 18103 36377
rect 18137 36343 18160 36377
rect 18080 36057 18160 36343
rect 18080 36023 18103 36057
rect 18137 36023 18160 36057
rect 18080 35737 18160 36023
rect 18080 35703 18103 35737
rect 18137 35703 18160 35737
rect 18080 35417 18160 35703
rect 18080 35383 18103 35417
rect 18137 35383 18160 35417
rect 18080 35097 18160 35383
rect 18080 35063 18103 35097
rect 18137 35063 18160 35097
rect 18080 34777 18160 35063
rect 18080 34743 18103 34777
rect 18137 34743 18160 34777
rect 18080 34457 18160 34743
rect 18080 34423 18103 34457
rect 18137 34423 18160 34457
rect 18080 34400 18160 34423
rect 18240 36377 18320 36400
rect 18240 36343 18263 36377
rect 18297 36343 18320 36377
rect 18240 36057 18320 36343
rect 18240 36023 18263 36057
rect 18297 36023 18320 36057
rect 18240 35737 18320 36023
rect 18240 35703 18263 35737
rect 18297 35703 18320 35737
rect 18240 35417 18320 35703
rect 18240 35383 18263 35417
rect 18297 35383 18320 35417
rect 18240 35097 18320 35383
rect 18240 35063 18263 35097
rect 18297 35063 18320 35097
rect 18240 34777 18320 35063
rect 18240 34743 18263 34777
rect 18297 34743 18320 34777
rect 18240 34457 18320 34743
rect 18240 34423 18263 34457
rect 18297 34423 18320 34457
rect 18240 34400 18320 34423
rect 18400 36377 18480 36400
rect 18400 36343 18423 36377
rect 18457 36343 18480 36377
rect 18400 36057 18480 36343
rect 18400 36023 18423 36057
rect 18457 36023 18480 36057
rect 18400 35737 18480 36023
rect 18400 35703 18423 35737
rect 18457 35703 18480 35737
rect 18400 35417 18480 35703
rect 18400 35383 18423 35417
rect 18457 35383 18480 35417
rect 18400 35097 18480 35383
rect 18400 35063 18423 35097
rect 18457 35063 18480 35097
rect 18400 34777 18480 35063
rect 18400 34743 18423 34777
rect 18457 34743 18480 34777
rect 18400 34457 18480 34743
rect 18400 34423 18423 34457
rect 18457 34423 18480 34457
rect 18400 34400 18480 34423
rect 18560 36377 18640 36400
rect 18560 36343 18583 36377
rect 18617 36343 18640 36377
rect 18560 36057 18640 36343
rect 18560 36023 18583 36057
rect 18617 36023 18640 36057
rect 18560 35737 18640 36023
rect 18560 35703 18583 35737
rect 18617 35703 18640 35737
rect 18560 35417 18640 35703
rect 18560 35383 18583 35417
rect 18617 35383 18640 35417
rect 18560 35097 18640 35383
rect 18560 35063 18583 35097
rect 18617 35063 18640 35097
rect 18560 34777 18640 35063
rect 18560 34743 18583 34777
rect 18617 34743 18640 34777
rect 18560 34457 18640 34743
rect 18560 34423 18583 34457
rect 18617 34423 18640 34457
rect 18560 34400 18640 34423
rect 18720 36377 18800 36400
rect 18720 36343 18743 36377
rect 18777 36343 18800 36377
rect 18720 36057 18800 36343
rect 18720 36023 18743 36057
rect 18777 36023 18800 36057
rect 18720 35737 18800 36023
rect 18720 35703 18743 35737
rect 18777 35703 18800 35737
rect 18720 35417 18800 35703
rect 18720 35383 18743 35417
rect 18777 35383 18800 35417
rect 18720 35097 18800 35383
rect 18720 35063 18743 35097
rect 18777 35063 18800 35097
rect 18720 34777 18800 35063
rect 18720 34743 18743 34777
rect 18777 34743 18800 34777
rect 18720 34457 18800 34743
rect 18720 34423 18743 34457
rect 18777 34423 18800 34457
rect 18720 34400 18800 34423
rect 18880 36377 18960 36400
rect 18880 36343 18903 36377
rect 18937 36343 18960 36377
rect 18880 36057 18960 36343
rect 18880 36023 18903 36057
rect 18937 36023 18960 36057
rect 18880 35737 18960 36023
rect 18880 35703 18903 35737
rect 18937 35703 18960 35737
rect 18880 35417 18960 35703
rect 18880 35383 18903 35417
rect 18937 35383 18960 35417
rect 18880 35097 18960 35383
rect 18880 35063 18903 35097
rect 18937 35063 18960 35097
rect 18880 34777 18960 35063
rect 18880 34743 18903 34777
rect 18937 34743 18960 34777
rect 18880 34457 18960 34743
rect 18880 34423 18903 34457
rect 18937 34423 18960 34457
rect 18880 34400 18960 34423
rect 19040 34400 19120 36400
rect 19200 34400 19280 36400
rect 19360 34400 19440 36400
rect 19520 34400 19600 36400
rect 19680 34400 19760 36400
rect 19840 34400 19920 36400
rect 20000 34400 20080 36400
rect 20160 34400 20240 36400
rect 20320 34400 20400 36400
rect 20480 34400 20560 36400
rect 20640 34400 20720 36400
rect 20800 34400 20880 36400
rect 20960 34400 21040 36400
rect 21120 34400 21200 36400
rect 21280 34400 21360 36400
rect 21440 34400 21520 36400
rect 21600 34400 21680 36400
rect 21760 34400 21840 36400
rect 21920 34400 22000 36400
rect 22080 34400 22160 36400
rect 22240 34400 22320 36400
rect 22400 34400 22480 36400
rect 22560 34400 22640 36400
rect 22720 34400 22800 36400
rect 22880 34400 22960 36400
rect 23120 36377 23200 36400
rect 23120 36343 23143 36377
rect 23177 36343 23200 36377
rect 23120 36057 23200 36343
rect 23120 36023 23143 36057
rect 23177 36023 23200 36057
rect 23120 35737 23200 36023
rect 23120 35703 23143 35737
rect 23177 35703 23200 35737
rect 23120 35417 23200 35703
rect 23120 35383 23143 35417
rect 23177 35383 23200 35417
rect 23120 35097 23200 35383
rect 23120 35063 23143 35097
rect 23177 35063 23200 35097
rect 23120 34777 23200 35063
rect 23120 34743 23143 34777
rect 23177 34743 23200 34777
rect 23120 34457 23200 34743
rect 23120 34423 23143 34457
rect 23177 34423 23200 34457
rect 23120 34400 23200 34423
rect 23280 36377 23360 36400
rect 23280 36343 23303 36377
rect 23337 36343 23360 36377
rect 23280 36057 23360 36343
rect 23280 36023 23303 36057
rect 23337 36023 23360 36057
rect 23280 35737 23360 36023
rect 23280 35703 23303 35737
rect 23337 35703 23360 35737
rect 23280 35417 23360 35703
rect 23280 35383 23303 35417
rect 23337 35383 23360 35417
rect 23280 35097 23360 35383
rect 23280 35063 23303 35097
rect 23337 35063 23360 35097
rect 23280 34777 23360 35063
rect 23280 34743 23303 34777
rect 23337 34743 23360 34777
rect 23280 34457 23360 34743
rect 23280 34423 23303 34457
rect 23337 34423 23360 34457
rect 23280 34400 23360 34423
rect 23440 36377 23520 36400
rect 23440 36343 23463 36377
rect 23497 36343 23520 36377
rect 23440 36057 23520 36343
rect 23440 36023 23463 36057
rect 23497 36023 23520 36057
rect 23440 35737 23520 36023
rect 23440 35703 23463 35737
rect 23497 35703 23520 35737
rect 23440 35417 23520 35703
rect 23440 35383 23463 35417
rect 23497 35383 23520 35417
rect 23440 35097 23520 35383
rect 23440 35063 23463 35097
rect 23497 35063 23520 35097
rect 23440 34777 23520 35063
rect 23440 34743 23463 34777
rect 23497 34743 23520 34777
rect 23440 34457 23520 34743
rect 23440 34423 23463 34457
rect 23497 34423 23520 34457
rect 23440 34400 23520 34423
rect 23600 36377 23680 36400
rect 23600 36343 23623 36377
rect 23657 36343 23680 36377
rect 23600 36057 23680 36343
rect 23600 36023 23623 36057
rect 23657 36023 23680 36057
rect 23600 35737 23680 36023
rect 23600 35703 23623 35737
rect 23657 35703 23680 35737
rect 23600 35417 23680 35703
rect 23600 35383 23623 35417
rect 23657 35383 23680 35417
rect 23600 35097 23680 35383
rect 23600 35063 23623 35097
rect 23657 35063 23680 35097
rect 23600 34777 23680 35063
rect 23600 34743 23623 34777
rect 23657 34743 23680 34777
rect 23600 34457 23680 34743
rect 23600 34423 23623 34457
rect 23657 34423 23680 34457
rect 23600 34400 23680 34423
rect 23760 36377 23840 36400
rect 23760 36343 23783 36377
rect 23817 36343 23840 36377
rect 23760 36057 23840 36343
rect 23760 36023 23783 36057
rect 23817 36023 23840 36057
rect 23760 35737 23840 36023
rect 23760 35703 23783 35737
rect 23817 35703 23840 35737
rect 23760 35417 23840 35703
rect 23760 35383 23783 35417
rect 23817 35383 23840 35417
rect 23760 35097 23840 35383
rect 23760 35063 23783 35097
rect 23817 35063 23840 35097
rect 23760 34777 23840 35063
rect 23760 34743 23783 34777
rect 23817 34743 23840 34777
rect 23760 34457 23840 34743
rect 23760 34423 23783 34457
rect 23817 34423 23840 34457
rect 23760 34400 23840 34423
rect 23920 36377 24000 36400
rect 23920 36343 23943 36377
rect 23977 36343 24000 36377
rect 23920 36057 24000 36343
rect 23920 36023 23943 36057
rect 23977 36023 24000 36057
rect 23920 35737 24000 36023
rect 23920 35703 23943 35737
rect 23977 35703 24000 35737
rect 23920 35417 24000 35703
rect 23920 35383 23943 35417
rect 23977 35383 24000 35417
rect 23920 35097 24000 35383
rect 23920 35063 23943 35097
rect 23977 35063 24000 35097
rect 23920 34777 24000 35063
rect 23920 34743 23943 34777
rect 23977 34743 24000 34777
rect 23920 34457 24000 34743
rect 23920 34423 23943 34457
rect 23977 34423 24000 34457
rect 23920 34400 24000 34423
rect 24080 36377 24160 36400
rect 24080 36343 24103 36377
rect 24137 36343 24160 36377
rect 24080 36057 24160 36343
rect 24080 36023 24103 36057
rect 24137 36023 24160 36057
rect 24080 35737 24160 36023
rect 24080 35703 24103 35737
rect 24137 35703 24160 35737
rect 24080 35417 24160 35703
rect 24080 35383 24103 35417
rect 24137 35383 24160 35417
rect 24080 35097 24160 35383
rect 24080 35063 24103 35097
rect 24137 35063 24160 35097
rect 24080 34777 24160 35063
rect 24080 34743 24103 34777
rect 24137 34743 24160 34777
rect 24080 34457 24160 34743
rect 24080 34423 24103 34457
rect 24137 34423 24160 34457
rect 24080 34400 24160 34423
rect 24240 36377 24320 36400
rect 24240 36343 24263 36377
rect 24297 36343 24320 36377
rect 24240 36057 24320 36343
rect 24240 36023 24263 36057
rect 24297 36023 24320 36057
rect 24240 35737 24320 36023
rect 24240 35703 24263 35737
rect 24297 35703 24320 35737
rect 24240 35417 24320 35703
rect 24240 35383 24263 35417
rect 24297 35383 24320 35417
rect 24240 35097 24320 35383
rect 24240 35063 24263 35097
rect 24297 35063 24320 35097
rect 24240 34777 24320 35063
rect 24240 34743 24263 34777
rect 24297 34743 24320 34777
rect 24240 34457 24320 34743
rect 24240 34423 24263 34457
rect 24297 34423 24320 34457
rect 24240 34400 24320 34423
rect 24400 36377 24480 36400
rect 24400 36343 24423 36377
rect 24457 36343 24480 36377
rect 24400 36057 24480 36343
rect 24400 36023 24423 36057
rect 24457 36023 24480 36057
rect 24400 35737 24480 36023
rect 24400 35703 24423 35737
rect 24457 35703 24480 35737
rect 24400 35417 24480 35703
rect 24400 35383 24423 35417
rect 24457 35383 24480 35417
rect 24400 35097 24480 35383
rect 24400 35063 24423 35097
rect 24457 35063 24480 35097
rect 24400 34777 24480 35063
rect 24400 34743 24423 34777
rect 24457 34743 24480 34777
rect 24400 34457 24480 34743
rect 24400 34423 24423 34457
rect 24457 34423 24480 34457
rect 24400 34400 24480 34423
rect 24560 36377 24640 36400
rect 24560 36343 24583 36377
rect 24617 36343 24640 36377
rect 24560 36057 24640 36343
rect 24560 36023 24583 36057
rect 24617 36023 24640 36057
rect 24560 35737 24640 36023
rect 24560 35703 24583 35737
rect 24617 35703 24640 35737
rect 24560 35417 24640 35703
rect 24560 35383 24583 35417
rect 24617 35383 24640 35417
rect 24560 35097 24640 35383
rect 24560 35063 24583 35097
rect 24617 35063 24640 35097
rect 24560 34777 24640 35063
rect 24560 34743 24583 34777
rect 24617 34743 24640 34777
rect 24560 34457 24640 34743
rect 24560 34423 24583 34457
rect 24617 34423 24640 34457
rect 24560 34400 24640 34423
rect 24720 36377 24800 36400
rect 24720 36343 24743 36377
rect 24777 36343 24800 36377
rect 24720 36057 24800 36343
rect 24720 36023 24743 36057
rect 24777 36023 24800 36057
rect 24720 35737 24800 36023
rect 24720 35703 24743 35737
rect 24777 35703 24800 35737
rect 24720 35417 24800 35703
rect 24720 35383 24743 35417
rect 24777 35383 24800 35417
rect 24720 35097 24800 35383
rect 24720 35063 24743 35097
rect 24777 35063 24800 35097
rect 24720 34777 24800 35063
rect 24720 34743 24743 34777
rect 24777 34743 24800 34777
rect 24720 34457 24800 34743
rect 24720 34423 24743 34457
rect 24777 34423 24800 34457
rect 24720 34400 24800 34423
rect 24880 36377 24960 36400
rect 24880 36343 24903 36377
rect 24937 36343 24960 36377
rect 24880 36057 24960 36343
rect 24880 36023 24903 36057
rect 24937 36023 24960 36057
rect 24880 35737 24960 36023
rect 24880 35703 24903 35737
rect 24937 35703 24960 35737
rect 24880 35417 24960 35703
rect 24880 35383 24903 35417
rect 24937 35383 24960 35417
rect 24880 35097 24960 35383
rect 24880 35063 24903 35097
rect 24937 35063 24960 35097
rect 24880 34777 24960 35063
rect 24880 34743 24903 34777
rect 24937 34743 24960 34777
rect 24880 34457 24960 34743
rect 24880 34423 24903 34457
rect 24937 34423 24960 34457
rect 24880 34400 24960 34423
rect 25040 36377 25120 36400
rect 25040 36343 25063 36377
rect 25097 36343 25120 36377
rect 25040 36057 25120 36343
rect 25040 36023 25063 36057
rect 25097 36023 25120 36057
rect 25040 35737 25120 36023
rect 25040 35703 25063 35737
rect 25097 35703 25120 35737
rect 25040 35417 25120 35703
rect 25040 35383 25063 35417
rect 25097 35383 25120 35417
rect 25040 35097 25120 35383
rect 25040 35063 25063 35097
rect 25097 35063 25120 35097
rect 25040 34777 25120 35063
rect 25040 34743 25063 34777
rect 25097 34743 25120 34777
rect 25040 34457 25120 34743
rect 25040 34423 25063 34457
rect 25097 34423 25120 34457
rect 25040 34400 25120 34423
rect 25200 36377 25280 36400
rect 25200 36343 25223 36377
rect 25257 36343 25280 36377
rect 25200 36057 25280 36343
rect 25200 36023 25223 36057
rect 25257 36023 25280 36057
rect 25200 35737 25280 36023
rect 25200 35703 25223 35737
rect 25257 35703 25280 35737
rect 25200 35417 25280 35703
rect 25200 35383 25223 35417
rect 25257 35383 25280 35417
rect 25200 35097 25280 35383
rect 25200 35063 25223 35097
rect 25257 35063 25280 35097
rect 25200 34777 25280 35063
rect 25200 34743 25223 34777
rect 25257 34743 25280 34777
rect 25200 34457 25280 34743
rect 25200 34423 25223 34457
rect 25257 34423 25280 34457
rect 25200 34400 25280 34423
rect 25360 36377 25440 36400
rect 25360 36343 25383 36377
rect 25417 36343 25440 36377
rect 25360 36057 25440 36343
rect 25360 36023 25383 36057
rect 25417 36023 25440 36057
rect 25360 35737 25440 36023
rect 25360 35703 25383 35737
rect 25417 35703 25440 35737
rect 25360 35417 25440 35703
rect 25360 35383 25383 35417
rect 25417 35383 25440 35417
rect 25360 35097 25440 35383
rect 25360 35063 25383 35097
rect 25417 35063 25440 35097
rect 25360 34777 25440 35063
rect 25360 34743 25383 34777
rect 25417 34743 25440 34777
rect 25360 34457 25440 34743
rect 25360 34423 25383 34457
rect 25417 34423 25440 34457
rect 25360 34400 25440 34423
rect 25520 36377 25600 36400
rect 25520 36343 25543 36377
rect 25577 36343 25600 36377
rect 25520 36057 25600 36343
rect 25520 36023 25543 36057
rect 25577 36023 25600 36057
rect 25520 35737 25600 36023
rect 25520 35703 25543 35737
rect 25577 35703 25600 35737
rect 25520 35417 25600 35703
rect 25520 35383 25543 35417
rect 25577 35383 25600 35417
rect 25520 35097 25600 35383
rect 25520 35063 25543 35097
rect 25577 35063 25600 35097
rect 25520 34777 25600 35063
rect 25520 34743 25543 34777
rect 25577 34743 25600 34777
rect 25520 34457 25600 34743
rect 25520 34423 25543 34457
rect 25577 34423 25600 34457
rect 25520 34400 25600 34423
rect 25680 36377 25760 36400
rect 25680 36343 25703 36377
rect 25737 36343 25760 36377
rect 25680 36057 25760 36343
rect 25680 36023 25703 36057
rect 25737 36023 25760 36057
rect 25680 35737 25760 36023
rect 25680 35703 25703 35737
rect 25737 35703 25760 35737
rect 25680 35417 25760 35703
rect 25680 35383 25703 35417
rect 25737 35383 25760 35417
rect 25680 35097 25760 35383
rect 25680 35063 25703 35097
rect 25737 35063 25760 35097
rect 25680 34777 25760 35063
rect 25680 34743 25703 34777
rect 25737 34743 25760 34777
rect 25680 34457 25760 34743
rect 25680 34423 25703 34457
rect 25737 34423 25760 34457
rect 25680 34400 25760 34423
rect 25840 36377 25920 36400
rect 25840 36343 25863 36377
rect 25897 36343 25920 36377
rect 25840 36057 25920 36343
rect 25840 36023 25863 36057
rect 25897 36023 25920 36057
rect 25840 35737 25920 36023
rect 25840 35703 25863 35737
rect 25897 35703 25920 35737
rect 25840 35417 25920 35703
rect 25840 35383 25863 35417
rect 25897 35383 25920 35417
rect 25840 35097 25920 35383
rect 25840 35063 25863 35097
rect 25897 35063 25920 35097
rect 25840 34777 25920 35063
rect 25840 34743 25863 34777
rect 25897 34743 25920 34777
rect 25840 34457 25920 34743
rect 25840 34423 25863 34457
rect 25897 34423 25920 34457
rect 25840 34400 25920 34423
rect 26000 36377 26080 36400
rect 26000 36343 26023 36377
rect 26057 36343 26080 36377
rect 26000 36057 26080 36343
rect 26000 36023 26023 36057
rect 26057 36023 26080 36057
rect 26000 35737 26080 36023
rect 26000 35703 26023 35737
rect 26057 35703 26080 35737
rect 26000 35417 26080 35703
rect 26000 35383 26023 35417
rect 26057 35383 26080 35417
rect 26000 35097 26080 35383
rect 26000 35063 26023 35097
rect 26057 35063 26080 35097
rect 26000 34777 26080 35063
rect 26000 34743 26023 34777
rect 26057 34743 26080 34777
rect 26000 34457 26080 34743
rect 26000 34423 26023 34457
rect 26057 34423 26080 34457
rect 26000 34400 26080 34423
rect 26160 36377 26240 36400
rect 26160 36343 26183 36377
rect 26217 36343 26240 36377
rect 26160 36057 26240 36343
rect 26160 36023 26183 36057
rect 26217 36023 26240 36057
rect 26160 35737 26240 36023
rect 26160 35703 26183 35737
rect 26217 35703 26240 35737
rect 26160 35417 26240 35703
rect 26160 35383 26183 35417
rect 26217 35383 26240 35417
rect 26160 35097 26240 35383
rect 26160 35063 26183 35097
rect 26217 35063 26240 35097
rect 26160 34777 26240 35063
rect 26160 34743 26183 34777
rect 26217 34743 26240 34777
rect 26160 34457 26240 34743
rect 26160 34423 26183 34457
rect 26217 34423 26240 34457
rect 26160 34400 26240 34423
rect 26320 36377 26400 36400
rect 26320 36343 26343 36377
rect 26377 36343 26400 36377
rect 26320 36057 26400 36343
rect 26320 36023 26343 36057
rect 26377 36023 26400 36057
rect 26320 35737 26400 36023
rect 26320 35703 26343 35737
rect 26377 35703 26400 35737
rect 26320 35417 26400 35703
rect 26320 35383 26343 35417
rect 26377 35383 26400 35417
rect 26320 35097 26400 35383
rect 26320 35063 26343 35097
rect 26377 35063 26400 35097
rect 26320 34777 26400 35063
rect 26320 34743 26343 34777
rect 26377 34743 26400 34777
rect 26320 34457 26400 34743
rect 26320 34423 26343 34457
rect 26377 34423 26400 34457
rect 26320 34400 26400 34423
rect 26480 36377 26560 36400
rect 26480 36343 26503 36377
rect 26537 36343 26560 36377
rect 26480 36057 26560 36343
rect 26480 36023 26503 36057
rect 26537 36023 26560 36057
rect 26480 35737 26560 36023
rect 26480 35703 26503 35737
rect 26537 35703 26560 35737
rect 26480 35417 26560 35703
rect 26480 35383 26503 35417
rect 26537 35383 26560 35417
rect 26480 35097 26560 35383
rect 26480 35063 26503 35097
rect 26537 35063 26560 35097
rect 26480 34777 26560 35063
rect 26480 34743 26503 34777
rect 26537 34743 26560 34777
rect 26480 34457 26560 34743
rect 26480 34423 26503 34457
rect 26537 34423 26560 34457
rect 26480 34400 26560 34423
rect 26640 36377 26720 36400
rect 26640 36343 26663 36377
rect 26697 36343 26720 36377
rect 26640 36057 26720 36343
rect 26640 36023 26663 36057
rect 26697 36023 26720 36057
rect 26640 35737 26720 36023
rect 26640 35703 26663 35737
rect 26697 35703 26720 35737
rect 26640 35417 26720 35703
rect 26640 35383 26663 35417
rect 26697 35383 26720 35417
rect 26640 35097 26720 35383
rect 26640 35063 26663 35097
rect 26697 35063 26720 35097
rect 26640 34777 26720 35063
rect 26640 34743 26663 34777
rect 26697 34743 26720 34777
rect 26640 34457 26720 34743
rect 26640 34423 26663 34457
rect 26697 34423 26720 34457
rect 26640 34400 26720 34423
rect 26800 36377 26880 36400
rect 26800 36343 26823 36377
rect 26857 36343 26880 36377
rect 26800 36057 26880 36343
rect 26800 36023 26823 36057
rect 26857 36023 26880 36057
rect 26800 35737 26880 36023
rect 26800 35703 26823 35737
rect 26857 35703 26880 35737
rect 26800 35417 26880 35703
rect 26800 35383 26823 35417
rect 26857 35383 26880 35417
rect 26800 35097 26880 35383
rect 26800 35063 26823 35097
rect 26857 35063 26880 35097
rect 26800 34777 26880 35063
rect 26800 34743 26823 34777
rect 26857 34743 26880 34777
rect 26800 34457 26880 34743
rect 26800 34423 26823 34457
rect 26857 34423 26880 34457
rect 26800 34400 26880 34423
rect 26960 36377 27040 36400
rect 26960 36343 26983 36377
rect 27017 36343 27040 36377
rect 26960 36057 27040 36343
rect 26960 36023 26983 36057
rect 27017 36023 27040 36057
rect 26960 35737 27040 36023
rect 26960 35703 26983 35737
rect 27017 35703 27040 35737
rect 26960 35417 27040 35703
rect 26960 35383 26983 35417
rect 27017 35383 27040 35417
rect 26960 35097 27040 35383
rect 26960 35063 26983 35097
rect 27017 35063 27040 35097
rect 26960 34777 27040 35063
rect 26960 34743 26983 34777
rect 27017 34743 27040 34777
rect 26960 34457 27040 34743
rect 26960 34423 26983 34457
rect 27017 34423 27040 34457
rect 26960 34400 27040 34423
rect 27120 36377 27200 36400
rect 27120 36343 27143 36377
rect 27177 36343 27200 36377
rect 27120 36057 27200 36343
rect 27120 36023 27143 36057
rect 27177 36023 27200 36057
rect 27120 35737 27200 36023
rect 27120 35703 27143 35737
rect 27177 35703 27200 35737
rect 27120 35417 27200 35703
rect 27120 35383 27143 35417
rect 27177 35383 27200 35417
rect 27120 35097 27200 35383
rect 27120 35063 27143 35097
rect 27177 35063 27200 35097
rect 27120 34777 27200 35063
rect 27120 34743 27143 34777
rect 27177 34743 27200 34777
rect 27120 34457 27200 34743
rect 27120 34423 27143 34457
rect 27177 34423 27200 34457
rect 27120 34400 27200 34423
rect 27280 36377 27360 36400
rect 27280 36343 27303 36377
rect 27337 36343 27360 36377
rect 27280 36057 27360 36343
rect 27280 36023 27303 36057
rect 27337 36023 27360 36057
rect 27280 35737 27360 36023
rect 27280 35703 27303 35737
rect 27337 35703 27360 35737
rect 27280 35417 27360 35703
rect 27280 35383 27303 35417
rect 27337 35383 27360 35417
rect 27280 35097 27360 35383
rect 27280 35063 27303 35097
rect 27337 35063 27360 35097
rect 27280 34777 27360 35063
rect 27280 34743 27303 34777
rect 27337 34743 27360 34777
rect 27280 34457 27360 34743
rect 27280 34423 27303 34457
rect 27337 34423 27360 34457
rect 27280 34400 27360 34423
rect 27440 36377 27520 36400
rect 27440 36343 27463 36377
rect 27497 36343 27520 36377
rect 27440 36057 27520 36343
rect 27440 36023 27463 36057
rect 27497 36023 27520 36057
rect 27440 35737 27520 36023
rect 27440 35703 27463 35737
rect 27497 35703 27520 35737
rect 27440 35417 27520 35703
rect 27440 35383 27463 35417
rect 27497 35383 27520 35417
rect 27440 35097 27520 35383
rect 27440 35063 27463 35097
rect 27497 35063 27520 35097
rect 27440 34777 27520 35063
rect 27440 34743 27463 34777
rect 27497 34743 27520 34777
rect 27440 34457 27520 34743
rect 27440 34423 27463 34457
rect 27497 34423 27520 34457
rect 27440 34400 27520 34423
rect 27600 36377 27680 36400
rect 27600 36343 27623 36377
rect 27657 36343 27680 36377
rect 27600 36057 27680 36343
rect 27600 36023 27623 36057
rect 27657 36023 27680 36057
rect 27600 35737 27680 36023
rect 27600 35703 27623 35737
rect 27657 35703 27680 35737
rect 27600 35417 27680 35703
rect 27600 35383 27623 35417
rect 27657 35383 27680 35417
rect 27600 35097 27680 35383
rect 27600 35063 27623 35097
rect 27657 35063 27680 35097
rect 27600 34777 27680 35063
rect 27600 34743 27623 34777
rect 27657 34743 27680 34777
rect 27600 34457 27680 34743
rect 27600 34423 27623 34457
rect 27657 34423 27680 34457
rect 27600 34400 27680 34423
rect 27760 36377 27840 36400
rect 27760 36343 27783 36377
rect 27817 36343 27840 36377
rect 27760 36057 27840 36343
rect 27760 36023 27783 36057
rect 27817 36023 27840 36057
rect 27760 35737 27840 36023
rect 27760 35703 27783 35737
rect 27817 35703 27840 35737
rect 27760 35417 27840 35703
rect 27760 35383 27783 35417
rect 27817 35383 27840 35417
rect 27760 35097 27840 35383
rect 27760 35063 27783 35097
rect 27817 35063 27840 35097
rect 27760 34777 27840 35063
rect 27760 34743 27783 34777
rect 27817 34743 27840 34777
rect 27760 34457 27840 34743
rect 27760 34423 27783 34457
rect 27817 34423 27840 34457
rect 27760 34400 27840 34423
rect 27920 36377 28000 36400
rect 27920 36343 27943 36377
rect 27977 36343 28000 36377
rect 27920 36057 28000 36343
rect 27920 36023 27943 36057
rect 27977 36023 28000 36057
rect 27920 35737 28000 36023
rect 27920 35703 27943 35737
rect 27977 35703 28000 35737
rect 27920 35417 28000 35703
rect 27920 35383 27943 35417
rect 27977 35383 28000 35417
rect 27920 35097 28000 35383
rect 27920 35063 27943 35097
rect 27977 35063 28000 35097
rect 27920 34777 28000 35063
rect 27920 34743 27943 34777
rect 27977 34743 28000 34777
rect 27920 34457 28000 34743
rect 27920 34423 27943 34457
rect 27977 34423 28000 34457
rect 27920 34400 28000 34423
rect 28080 36377 28160 36400
rect 28080 36343 28103 36377
rect 28137 36343 28160 36377
rect 28080 36057 28160 36343
rect 28080 36023 28103 36057
rect 28137 36023 28160 36057
rect 28080 35737 28160 36023
rect 28080 35703 28103 35737
rect 28137 35703 28160 35737
rect 28080 35417 28160 35703
rect 28080 35383 28103 35417
rect 28137 35383 28160 35417
rect 28080 35097 28160 35383
rect 28080 35063 28103 35097
rect 28137 35063 28160 35097
rect 28080 34777 28160 35063
rect 28080 34743 28103 34777
rect 28137 34743 28160 34777
rect 28080 34457 28160 34743
rect 28080 34423 28103 34457
rect 28137 34423 28160 34457
rect 28080 34400 28160 34423
rect 28240 36377 28320 36400
rect 28240 36343 28263 36377
rect 28297 36343 28320 36377
rect 28240 36057 28320 36343
rect 28240 36023 28263 36057
rect 28297 36023 28320 36057
rect 28240 35737 28320 36023
rect 28240 35703 28263 35737
rect 28297 35703 28320 35737
rect 28240 35417 28320 35703
rect 28240 35383 28263 35417
rect 28297 35383 28320 35417
rect 28240 35097 28320 35383
rect 28240 35063 28263 35097
rect 28297 35063 28320 35097
rect 28240 34777 28320 35063
rect 28240 34743 28263 34777
rect 28297 34743 28320 34777
rect 28240 34457 28320 34743
rect 28240 34423 28263 34457
rect 28297 34423 28320 34457
rect 28240 34400 28320 34423
rect 28400 36377 28480 36400
rect 28400 36343 28423 36377
rect 28457 36343 28480 36377
rect 28400 36057 28480 36343
rect 28400 36023 28423 36057
rect 28457 36023 28480 36057
rect 28400 35737 28480 36023
rect 28400 35703 28423 35737
rect 28457 35703 28480 35737
rect 28400 35417 28480 35703
rect 28400 35383 28423 35417
rect 28457 35383 28480 35417
rect 28400 35097 28480 35383
rect 28400 35063 28423 35097
rect 28457 35063 28480 35097
rect 28400 34777 28480 35063
rect 28400 34743 28423 34777
rect 28457 34743 28480 34777
rect 28400 34457 28480 34743
rect 28400 34423 28423 34457
rect 28457 34423 28480 34457
rect 28400 34400 28480 34423
rect 28560 36377 28640 36400
rect 28560 36343 28583 36377
rect 28617 36343 28640 36377
rect 28560 36057 28640 36343
rect 28560 36023 28583 36057
rect 28617 36023 28640 36057
rect 28560 35737 28640 36023
rect 28560 35703 28583 35737
rect 28617 35703 28640 35737
rect 28560 35417 28640 35703
rect 28560 35383 28583 35417
rect 28617 35383 28640 35417
rect 28560 35097 28640 35383
rect 28560 35063 28583 35097
rect 28617 35063 28640 35097
rect 28560 34777 28640 35063
rect 28560 34743 28583 34777
rect 28617 34743 28640 34777
rect 28560 34457 28640 34743
rect 28560 34423 28583 34457
rect 28617 34423 28640 34457
rect 28560 34400 28640 34423
rect 28720 36377 28800 36400
rect 28720 36343 28743 36377
rect 28777 36343 28800 36377
rect 28720 36057 28800 36343
rect 28720 36023 28743 36057
rect 28777 36023 28800 36057
rect 28720 35737 28800 36023
rect 28720 35703 28743 35737
rect 28777 35703 28800 35737
rect 28720 35417 28800 35703
rect 28720 35383 28743 35417
rect 28777 35383 28800 35417
rect 28720 35097 28800 35383
rect 28720 35063 28743 35097
rect 28777 35063 28800 35097
rect 28720 34777 28800 35063
rect 28720 34743 28743 34777
rect 28777 34743 28800 34777
rect 28720 34457 28800 34743
rect 28720 34423 28743 34457
rect 28777 34423 28800 34457
rect 28720 34400 28800 34423
rect 28880 36377 28960 36400
rect 28880 36343 28903 36377
rect 28937 36343 28960 36377
rect 28880 36057 28960 36343
rect 28880 36023 28903 36057
rect 28937 36023 28960 36057
rect 28880 35737 28960 36023
rect 28880 35703 28903 35737
rect 28937 35703 28960 35737
rect 28880 35417 28960 35703
rect 28880 35383 28903 35417
rect 28937 35383 28960 35417
rect 28880 35097 28960 35383
rect 28880 35063 28903 35097
rect 28937 35063 28960 35097
rect 28880 34777 28960 35063
rect 28880 34743 28903 34777
rect 28937 34743 28960 34777
rect 28880 34457 28960 34743
rect 28880 34423 28903 34457
rect 28937 34423 28960 34457
rect 28880 34400 28960 34423
rect 29040 36377 29120 36400
rect 29040 36343 29063 36377
rect 29097 36343 29120 36377
rect 29040 36057 29120 36343
rect 29040 36023 29063 36057
rect 29097 36023 29120 36057
rect 29040 35737 29120 36023
rect 29040 35703 29063 35737
rect 29097 35703 29120 35737
rect 29040 35417 29120 35703
rect 29040 35383 29063 35417
rect 29097 35383 29120 35417
rect 29040 35097 29120 35383
rect 29040 35063 29063 35097
rect 29097 35063 29120 35097
rect 29040 34777 29120 35063
rect 29040 34743 29063 34777
rect 29097 34743 29120 34777
rect 29040 34457 29120 34743
rect 29040 34423 29063 34457
rect 29097 34423 29120 34457
rect 29040 34400 29120 34423
rect 29200 36377 29280 36400
rect 29200 36343 29223 36377
rect 29257 36343 29280 36377
rect 29200 36057 29280 36343
rect 29200 36023 29223 36057
rect 29257 36023 29280 36057
rect 29200 35737 29280 36023
rect 29200 35703 29223 35737
rect 29257 35703 29280 35737
rect 29200 35417 29280 35703
rect 29200 35383 29223 35417
rect 29257 35383 29280 35417
rect 29200 35097 29280 35383
rect 29200 35063 29223 35097
rect 29257 35063 29280 35097
rect 29200 34777 29280 35063
rect 29200 34743 29223 34777
rect 29257 34743 29280 34777
rect 29200 34457 29280 34743
rect 29200 34423 29223 34457
rect 29257 34423 29280 34457
rect 29200 34400 29280 34423
rect 29360 36377 29440 36400
rect 29360 36343 29383 36377
rect 29417 36343 29440 36377
rect 29360 36057 29440 36343
rect 29360 36023 29383 36057
rect 29417 36023 29440 36057
rect 29360 35737 29440 36023
rect 29360 35703 29383 35737
rect 29417 35703 29440 35737
rect 29360 35417 29440 35703
rect 29360 35383 29383 35417
rect 29417 35383 29440 35417
rect 29360 35097 29440 35383
rect 29360 35063 29383 35097
rect 29417 35063 29440 35097
rect 29360 34777 29440 35063
rect 29360 34743 29383 34777
rect 29417 34743 29440 34777
rect 29360 34457 29440 34743
rect 29360 34423 29383 34457
rect 29417 34423 29440 34457
rect 29360 34400 29440 34423
rect 29520 34400 29600 36400
rect 29680 34400 29760 36400
rect 29840 34400 29920 36400
rect 30000 34400 30080 36400
rect 30160 34400 30240 36400
rect 30320 34400 30400 36400
rect 30480 34400 30560 36400
rect 30640 34400 30720 36400
rect 30800 34400 30880 36400
rect 30960 34400 31040 36400
rect 31120 34400 31200 36400
rect 31280 34400 31360 36400
rect 31440 34400 31520 36400
rect 31600 34400 31680 36400
rect 31760 34400 31840 36400
rect 31920 34400 32000 36400
rect 32080 34400 32160 36400
rect 32240 34400 32320 36400
rect 32400 34400 32480 36400
rect 32560 34400 32640 36400
rect 32720 34400 32800 36400
rect 32880 34400 32960 36400
rect 33040 34400 33120 36400
rect 33200 34400 33280 36400
rect 33360 34400 33440 36400
rect 33520 36377 33600 36400
rect 33520 36343 33543 36377
rect 33577 36343 33600 36377
rect 33520 36057 33600 36343
rect 33520 36023 33543 36057
rect 33577 36023 33600 36057
rect 33520 35737 33600 36023
rect 33520 35703 33543 35737
rect 33577 35703 33600 35737
rect 33520 35417 33600 35703
rect 33520 35383 33543 35417
rect 33577 35383 33600 35417
rect 33520 35097 33600 35383
rect 33520 35063 33543 35097
rect 33577 35063 33600 35097
rect 33520 34777 33600 35063
rect 33520 34743 33543 34777
rect 33577 34743 33600 34777
rect 33520 34457 33600 34743
rect 33520 34423 33543 34457
rect 33577 34423 33600 34457
rect 33520 34400 33600 34423
rect 33680 36377 33760 36400
rect 33680 36343 33703 36377
rect 33737 36343 33760 36377
rect 33680 36057 33760 36343
rect 33680 36023 33703 36057
rect 33737 36023 33760 36057
rect 33680 35737 33760 36023
rect 33680 35703 33703 35737
rect 33737 35703 33760 35737
rect 33680 35417 33760 35703
rect 33680 35383 33703 35417
rect 33737 35383 33760 35417
rect 33680 35097 33760 35383
rect 33680 35063 33703 35097
rect 33737 35063 33760 35097
rect 33680 34777 33760 35063
rect 33680 34743 33703 34777
rect 33737 34743 33760 34777
rect 33680 34457 33760 34743
rect 33680 34423 33703 34457
rect 33737 34423 33760 34457
rect 33680 34400 33760 34423
rect 33840 36377 33920 36400
rect 33840 36343 33863 36377
rect 33897 36343 33920 36377
rect 33840 36057 33920 36343
rect 33840 36023 33863 36057
rect 33897 36023 33920 36057
rect 33840 35737 33920 36023
rect 33840 35703 33863 35737
rect 33897 35703 33920 35737
rect 33840 35417 33920 35703
rect 33840 35383 33863 35417
rect 33897 35383 33920 35417
rect 33840 35097 33920 35383
rect 33840 35063 33863 35097
rect 33897 35063 33920 35097
rect 33840 34777 33920 35063
rect 33840 34743 33863 34777
rect 33897 34743 33920 34777
rect 33840 34457 33920 34743
rect 33840 34423 33863 34457
rect 33897 34423 33920 34457
rect 33840 34400 33920 34423
rect 34000 36377 34080 36400
rect 34000 36343 34023 36377
rect 34057 36343 34080 36377
rect 34000 36057 34080 36343
rect 34000 36023 34023 36057
rect 34057 36023 34080 36057
rect 34000 35737 34080 36023
rect 34000 35703 34023 35737
rect 34057 35703 34080 35737
rect 34000 35417 34080 35703
rect 34000 35383 34023 35417
rect 34057 35383 34080 35417
rect 34000 35097 34080 35383
rect 34000 35063 34023 35097
rect 34057 35063 34080 35097
rect 34000 34777 34080 35063
rect 34000 34743 34023 34777
rect 34057 34743 34080 34777
rect 34000 34457 34080 34743
rect 34000 34423 34023 34457
rect 34057 34423 34080 34457
rect 34000 34400 34080 34423
rect 34160 36377 34240 36400
rect 34160 36343 34183 36377
rect 34217 36343 34240 36377
rect 34160 36057 34240 36343
rect 34160 36023 34183 36057
rect 34217 36023 34240 36057
rect 34160 35737 34240 36023
rect 34160 35703 34183 35737
rect 34217 35703 34240 35737
rect 34160 35417 34240 35703
rect 34160 35383 34183 35417
rect 34217 35383 34240 35417
rect 34160 35097 34240 35383
rect 34160 35063 34183 35097
rect 34217 35063 34240 35097
rect 34160 34777 34240 35063
rect 34160 34743 34183 34777
rect 34217 34743 34240 34777
rect 34160 34457 34240 34743
rect 34160 34423 34183 34457
rect 34217 34423 34240 34457
rect 34160 34400 34240 34423
rect 34320 36377 34400 36400
rect 34320 36343 34343 36377
rect 34377 36343 34400 36377
rect 34320 36057 34400 36343
rect 34320 36023 34343 36057
rect 34377 36023 34400 36057
rect 34320 35737 34400 36023
rect 34320 35703 34343 35737
rect 34377 35703 34400 35737
rect 34320 35417 34400 35703
rect 34320 35383 34343 35417
rect 34377 35383 34400 35417
rect 34320 35097 34400 35383
rect 34320 35063 34343 35097
rect 34377 35063 34400 35097
rect 34320 34777 34400 35063
rect 34320 34743 34343 34777
rect 34377 34743 34400 34777
rect 34320 34457 34400 34743
rect 34320 34423 34343 34457
rect 34377 34423 34400 34457
rect 34320 34400 34400 34423
rect 34480 36377 34560 36400
rect 34480 36343 34503 36377
rect 34537 36343 34560 36377
rect 34480 36057 34560 36343
rect 34480 36023 34503 36057
rect 34537 36023 34560 36057
rect 34480 35737 34560 36023
rect 34480 35703 34503 35737
rect 34537 35703 34560 35737
rect 34480 35417 34560 35703
rect 34480 35383 34503 35417
rect 34537 35383 34560 35417
rect 34480 35097 34560 35383
rect 34480 35063 34503 35097
rect 34537 35063 34560 35097
rect 34480 34777 34560 35063
rect 34480 34743 34503 34777
rect 34537 34743 34560 34777
rect 34480 34457 34560 34743
rect 34480 34423 34503 34457
rect 34537 34423 34560 34457
rect 34480 34400 34560 34423
rect 34640 36377 34720 36400
rect 34640 36343 34663 36377
rect 34697 36343 34720 36377
rect 34640 36057 34720 36343
rect 34640 36023 34663 36057
rect 34697 36023 34720 36057
rect 34640 35737 34720 36023
rect 34640 35703 34663 35737
rect 34697 35703 34720 35737
rect 34640 35417 34720 35703
rect 34640 35383 34663 35417
rect 34697 35383 34720 35417
rect 34640 35097 34720 35383
rect 34640 35063 34663 35097
rect 34697 35063 34720 35097
rect 34640 34777 34720 35063
rect 34640 34743 34663 34777
rect 34697 34743 34720 34777
rect 34640 34457 34720 34743
rect 34640 34423 34663 34457
rect 34697 34423 34720 34457
rect 34640 34400 34720 34423
rect 34800 36377 34880 36400
rect 34800 36343 34823 36377
rect 34857 36343 34880 36377
rect 34800 36057 34880 36343
rect 34800 36023 34823 36057
rect 34857 36023 34880 36057
rect 34800 35737 34880 36023
rect 34800 35703 34823 35737
rect 34857 35703 34880 35737
rect 34800 35417 34880 35703
rect 34800 35383 34823 35417
rect 34857 35383 34880 35417
rect 34800 35097 34880 35383
rect 34800 35063 34823 35097
rect 34857 35063 34880 35097
rect 34800 34777 34880 35063
rect 34800 34743 34823 34777
rect 34857 34743 34880 34777
rect 34800 34457 34880 34743
rect 34800 34423 34823 34457
rect 34857 34423 34880 34457
rect 34800 34400 34880 34423
rect 34960 36377 35040 36400
rect 34960 36343 34983 36377
rect 35017 36343 35040 36377
rect 34960 36057 35040 36343
rect 34960 36023 34983 36057
rect 35017 36023 35040 36057
rect 34960 35737 35040 36023
rect 34960 35703 34983 35737
rect 35017 35703 35040 35737
rect 34960 35417 35040 35703
rect 34960 35383 34983 35417
rect 35017 35383 35040 35417
rect 34960 35097 35040 35383
rect 34960 35063 34983 35097
rect 35017 35063 35040 35097
rect 34960 34777 35040 35063
rect 34960 34743 34983 34777
rect 35017 34743 35040 34777
rect 34960 34457 35040 34743
rect 34960 34423 34983 34457
rect 35017 34423 35040 34457
rect 34960 34400 35040 34423
rect 35120 36377 35200 36400
rect 35120 36343 35143 36377
rect 35177 36343 35200 36377
rect 35120 36057 35200 36343
rect 35120 36023 35143 36057
rect 35177 36023 35200 36057
rect 35120 35737 35200 36023
rect 35120 35703 35143 35737
rect 35177 35703 35200 35737
rect 35120 35417 35200 35703
rect 35120 35383 35143 35417
rect 35177 35383 35200 35417
rect 35120 35097 35200 35383
rect 35120 35063 35143 35097
rect 35177 35063 35200 35097
rect 35120 34777 35200 35063
rect 35120 34743 35143 34777
rect 35177 34743 35200 34777
rect 35120 34457 35200 34743
rect 35120 34423 35143 34457
rect 35177 34423 35200 34457
rect 35120 34400 35200 34423
rect 35280 36377 35360 36400
rect 35280 36343 35303 36377
rect 35337 36343 35360 36377
rect 35280 36057 35360 36343
rect 35280 36023 35303 36057
rect 35337 36023 35360 36057
rect 35280 35737 35360 36023
rect 35280 35703 35303 35737
rect 35337 35703 35360 35737
rect 35280 35417 35360 35703
rect 35280 35383 35303 35417
rect 35337 35383 35360 35417
rect 35280 35097 35360 35383
rect 35280 35063 35303 35097
rect 35337 35063 35360 35097
rect 35280 34777 35360 35063
rect 35280 34743 35303 34777
rect 35337 34743 35360 34777
rect 35280 34457 35360 34743
rect 35280 34423 35303 34457
rect 35337 34423 35360 34457
rect 35280 34400 35360 34423
rect 35440 36377 35520 36400
rect 35440 36343 35463 36377
rect 35497 36343 35520 36377
rect 35440 36057 35520 36343
rect 35440 36023 35463 36057
rect 35497 36023 35520 36057
rect 35440 35737 35520 36023
rect 35440 35703 35463 35737
rect 35497 35703 35520 35737
rect 35440 35417 35520 35703
rect 35440 35383 35463 35417
rect 35497 35383 35520 35417
rect 35440 35097 35520 35383
rect 35440 35063 35463 35097
rect 35497 35063 35520 35097
rect 35440 34777 35520 35063
rect 35440 34743 35463 34777
rect 35497 34743 35520 34777
rect 35440 34457 35520 34743
rect 35440 34423 35463 34457
rect 35497 34423 35520 34457
rect 35440 34400 35520 34423
rect 35600 36377 35680 36400
rect 35600 36343 35623 36377
rect 35657 36343 35680 36377
rect 35600 36057 35680 36343
rect 35600 36023 35623 36057
rect 35657 36023 35680 36057
rect 35600 35737 35680 36023
rect 35600 35703 35623 35737
rect 35657 35703 35680 35737
rect 35600 35417 35680 35703
rect 35600 35383 35623 35417
rect 35657 35383 35680 35417
rect 35600 35097 35680 35383
rect 35600 35063 35623 35097
rect 35657 35063 35680 35097
rect 35600 34777 35680 35063
rect 35600 34743 35623 34777
rect 35657 34743 35680 34777
rect 35600 34457 35680 34743
rect 35600 34423 35623 34457
rect 35657 34423 35680 34457
rect 35600 34400 35680 34423
rect 35760 36377 35840 36400
rect 35760 36343 35783 36377
rect 35817 36343 35840 36377
rect 35760 36057 35840 36343
rect 35760 36023 35783 36057
rect 35817 36023 35840 36057
rect 35760 35737 35840 36023
rect 35760 35703 35783 35737
rect 35817 35703 35840 35737
rect 35760 35417 35840 35703
rect 35760 35383 35783 35417
rect 35817 35383 35840 35417
rect 35760 35097 35840 35383
rect 35760 35063 35783 35097
rect 35817 35063 35840 35097
rect 35760 34777 35840 35063
rect 35760 34743 35783 34777
rect 35817 34743 35840 34777
rect 35760 34457 35840 34743
rect 35760 34423 35783 34457
rect 35817 34423 35840 34457
rect 35760 34400 35840 34423
rect 35920 36377 36000 36400
rect 35920 36343 35943 36377
rect 35977 36343 36000 36377
rect 35920 36057 36000 36343
rect 35920 36023 35943 36057
rect 35977 36023 36000 36057
rect 35920 35737 36000 36023
rect 35920 35703 35943 35737
rect 35977 35703 36000 35737
rect 35920 35417 36000 35703
rect 35920 35383 35943 35417
rect 35977 35383 36000 35417
rect 35920 35097 36000 35383
rect 35920 35063 35943 35097
rect 35977 35063 36000 35097
rect 35920 34777 36000 35063
rect 35920 34743 35943 34777
rect 35977 34743 36000 34777
rect 35920 34457 36000 34743
rect 35920 34423 35943 34457
rect 35977 34423 36000 34457
rect 35920 34400 36000 34423
rect 36080 36377 36160 36400
rect 36080 36343 36103 36377
rect 36137 36343 36160 36377
rect 36080 36057 36160 36343
rect 36080 36023 36103 36057
rect 36137 36023 36160 36057
rect 36080 35737 36160 36023
rect 36080 35703 36103 35737
rect 36137 35703 36160 35737
rect 36080 35417 36160 35703
rect 36080 35383 36103 35417
rect 36137 35383 36160 35417
rect 36080 35097 36160 35383
rect 36080 35063 36103 35097
rect 36137 35063 36160 35097
rect 36080 34777 36160 35063
rect 36080 34743 36103 34777
rect 36137 34743 36160 34777
rect 36080 34457 36160 34743
rect 36080 34423 36103 34457
rect 36137 34423 36160 34457
rect 36080 34400 36160 34423
rect 36240 36377 36320 36400
rect 36240 36343 36263 36377
rect 36297 36343 36320 36377
rect 36240 36057 36320 36343
rect 36240 36023 36263 36057
rect 36297 36023 36320 36057
rect 36240 35737 36320 36023
rect 36240 35703 36263 35737
rect 36297 35703 36320 35737
rect 36240 35417 36320 35703
rect 36240 35383 36263 35417
rect 36297 35383 36320 35417
rect 36240 35097 36320 35383
rect 36240 35063 36263 35097
rect 36297 35063 36320 35097
rect 36240 34777 36320 35063
rect 36240 34743 36263 34777
rect 36297 34743 36320 34777
rect 36240 34457 36320 34743
rect 36240 34423 36263 34457
rect 36297 34423 36320 34457
rect 36240 34400 36320 34423
rect 36400 36377 36480 36400
rect 36400 36343 36423 36377
rect 36457 36343 36480 36377
rect 36400 36057 36480 36343
rect 36400 36023 36423 36057
rect 36457 36023 36480 36057
rect 36400 35737 36480 36023
rect 36400 35703 36423 35737
rect 36457 35703 36480 35737
rect 36400 35417 36480 35703
rect 36400 35383 36423 35417
rect 36457 35383 36480 35417
rect 36400 35097 36480 35383
rect 36400 35063 36423 35097
rect 36457 35063 36480 35097
rect 36400 34777 36480 35063
rect 36400 34743 36423 34777
rect 36457 34743 36480 34777
rect 36400 34457 36480 34743
rect 36400 34423 36423 34457
rect 36457 34423 36480 34457
rect 36400 34400 36480 34423
rect 36560 36377 36640 36400
rect 36560 36343 36583 36377
rect 36617 36343 36640 36377
rect 36560 36057 36640 36343
rect 36560 36023 36583 36057
rect 36617 36023 36640 36057
rect 36560 35737 36640 36023
rect 36560 35703 36583 35737
rect 36617 35703 36640 35737
rect 36560 35417 36640 35703
rect 36560 35383 36583 35417
rect 36617 35383 36640 35417
rect 36560 35097 36640 35383
rect 36560 35063 36583 35097
rect 36617 35063 36640 35097
rect 36560 34777 36640 35063
rect 36560 34743 36583 34777
rect 36617 34743 36640 34777
rect 36560 34457 36640 34743
rect 36560 34423 36583 34457
rect 36617 34423 36640 34457
rect 36560 34400 36640 34423
rect 36720 36377 36800 36400
rect 36720 36343 36743 36377
rect 36777 36343 36800 36377
rect 36720 36057 36800 36343
rect 36720 36023 36743 36057
rect 36777 36023 36800 36057
rect 36720 35737 36800 36023
rect 36720 35703 36743 35737
rect 36777 35703 36800 35737
rect 36720 35417 36800 35703
rect 36720 35383 36743 35417
rect 36777 35383 36800 35417
rect 36720 35097 36800 35383
rect 36720 35063 36743 35097
rect 36777 35063 36800 35097
rect 36720 34777 36800 35063
rect 36720 34743 36743 34777
rect 36777 34743 36800 34777
rect 36720 34457 36800 34743
rect 36720 34423 36743 34457
rect 36777 34423 36800 34457
rect 36720 34400 36800 34423
rect 36880 36377 36960 36400
rect 36880 36343 36903 36377
rect 36937 36343 36960 36377
rect 36880 36057 36960 36343
rect 36880 36023 36903 36057
rect 36937 36023 36960 36057
rect 36880 35737 36960 36023
rect 36880 35703 36903 35737
rect 36937 35703 36960 35737
rect 36880 35417 36960 35703
rect 36880 35383 36903 35417
rect 36937 35383 36960 35417
rect 36880 35097 36960 35383
rect 36880 35063 36903 35097
rect 36937 35063 36960 35097
rect 36880 34777 36960 35063
rect 36880 34743 36903 34777
rect 36937 34743 36960 34777
rect 36880 34457 36960 34743
rect 36880 34423 36903 34457
rect 36937 34423 36960 34457
rect 36880 34400 36960 34423
rect 37040 36377 37120 36400
rect 37040 36343 37063 36377
rect 37097 36343 37120 36377
rect 37040 36057 37120 36343
rect 37040 36023 37063 36057
rect 37097 36023 37120 36057
rect 37040 35737 37120 36023
rect 37040 35703 37063 35737
rect 37097 35703 37120 35737
rect 37040 35417 37120 35703
rect 37040 35383 37063 35417
rect 37097 35383 37120 35417
rect 37040 35097 37120 35383
rect 37040 35063 37063 35097
rect 37097 35063 37120 35097
rect 37040 34777 37120 35063
rect 37040 34743 37063 34777
rect 37097 34743 37120 34777
rect 37040 34457 37120 34743
rect 37040 34423 37063 34457
rect 37097 34423 37120 34457
rect 37040 34400 37120 34423
rect 37200 36377 37280 36400
rect 37200 36343 37223 36377
rect 37257 36343 37280 36377
rect 37200 36057 37280 36343
rect 37200 36023 37223 36057
rect 37257 36023 37280 36057
rect 37200 35737 37280 36023
rect 37200 35703 37223 35737
rect 37257 35703 37280 35737
rect 37200 35417 37280 35703
rect 37200 35383 37223 35417
rect 37257 35383 37280 35417
rect 37200 35097 37280 35383
rect 37200 35063 37223 35097
rect 37257 35063 37280 35097
rect 37200 34777 37280 35063
rect 37200 34743 37223 34777
rect 37257 34743 37280 34777
rect 37200 34457 37280 34743
rect 37200 34423 37223 34457
rect 37257 34423 37280 34457
rect 37200 34400 37280 34423
rect 37360 36377 37440 36400
rect 37360 36343 37383 36377
rect 37417 36343 37440 36377
rect 37360 36057 37440 36343
rect 37360 36023 37383 36057
rect 37417 36023 37440 36057
rect 37360 35737 37440 36023
rect 37360 35703 37383 35737
rect 37417 35703 37440 35737
rect 37360 35417 37440 35703
rect 37360 35383 37383 35417
rect 37417 35383 37440 35417
rect 37360 35097 37440 35383
rect 37360 35063 37383 35097
rect 37417 35063 37440 35097
rect 37360 34777 37440 35063
rect 37360 34743 37383 34777
rect 37417 34743 37440 34777
rect 37360 34457 37440 34743
rect 37360 34423 37383 34457
rect 37417 34423 37440 34457
rect 37360 34400 37440 34423
rect 37520 36377 37600 36400
rect 37520 36343 37543 36377
rect 37577 36343 37600 36377
rect 37520 36057 37600 36343
rect 37520 36023 37543 36057
rect 37577 36023 37600 36057
rect 37520 35737 37600 36023
rect 37520 35703 37543 35737
rect 37577 35703 37600 35737
rect 37520 35417 37600 35703
rect 37520 35383 37543 35417
rect 37577 35383 37600 35417
rect 37520 35097 37600 35383
rect 37520 35063 37543 35097
rect 37577 35063 37600 35097
rect 37520 34777 37600 35063
rect 37520 34743 37543 34777
rect 37577 34743 37600 34777
rect 37520 34457 37600 34743
rect 37520 34423 37543 34457
rect 37577 34423 37600 34457
rect 37520 34400 37600 34423
rect 37680 36377 37760 36400
rect 37680 36343 37703 36377
rect 37737 36343 37760 36377
rect 37680 36057 37760 36343
rect 37680 36023 37703 36057
rect 37737 36023 37760 36057
rect 37680 35737 37760 36023
rect 37680 35703 37703 35737
rect 37737 35703 37760 35737
rect 37680 35417 37760 35703
rect 37680 35383 37703 35417
rect 37737 35383 37760 35417
rect 37680 35097 37760 35383
rect 37680 35063 37703 35097
rect 37737 35063 37760 35097
rect 37680 34777 37760 35063
rect 37680 34743 37703 34777
rect 37737 34743 37760 34777
rect 37680 34457 37760 34743
rect 37680 34423 37703 34457
rect 37737 34423 37760 34457
rect 37680 34400 37760 34423
rect 37840 36377 37920 36400
rect 37840 36343 37863 36377
rect 37897 36343 37920 36377
rect 37840 36057 37920 36343
rect 37840 36023 37863 36057
rect 37897 36023 37920 36057
rect 37840 35737 37920 36023
rect 37840 35703 37863 35737
rect 37897 35703 37920 35737
rect 37840 35417 37920 35703
rect 37840 35383 37863 35417
rect 37897 35383 37920 35417
rect 37840 35097 37920 35383
rect 37840 35063 37863 35097
rect 37897 35063 37920 35097
rect 37840 34777 37920 35063
rect 37840 34743 37863 34777
rect 37897 34743 37920 34777
rect 37840 34457 37920 34743
rect 37840 34423 37863 34457
rect 37897 34423 37920 34457
rect 37840 34400 37920 34423
rect 38000 36377 38080 36400
rect 38000 36343 38023 36377
rect 38057 36343 38080 36377
rect 38000 36057 38080 36343
rect 38000 36023 38023 36057
rect 38057 36023 38080 36057
rect 38000 35737 38080 36023
rect 38000 35703 38023 35737
rect 38057 35703 38080 35737
rect 38000 35417 38080 35703
rect 38000 35383 38023 35417
rect 38057 35383 38080 35417
rect 38000 35097 38080 35383
rect 38000 35063 38023 35097
rect 38057 35063 38080 35097
rect 38000 34777 38080 35063
rect 38000 34743 38023 34777
rect 38057 34743 38080 34777
rect 38000 34457 38080 34743
rect 38000 34423 38023 34457
rect 38057 34423 38080 34457
rect 38000 34400 38080 34423
rect 38160 36377 38240 36400
rect 38160 36343 38183 36377
rect 38217 36343 38240 36377
rect 38160 36057 38240 36343
rect 38160 36023 38183 36057
rect 38217 36023 38240 36057
rect 38160 35737 38240 36023
rect 38160 35703 38183 35737
rect 38217 35703 38240 35737
rect 38160 35417 38240 35703
rect 38160 35383 38183 35417
rect 38217 35383 38240 35417
rect 38160 35097 38240 35383
rect 38160 35063 38183 35097
rect 38217 35063 38240 35097
rect 38160 34777 38240 35063
rect 38160 34743 38183 34777
rect 38217 34743 38240 34777
rect 38160 34457 38240 34743
rect 38160 34423 38183 34457
rect 38217 34423 38240 34457
rect 38160 34400 38240 34423
rect 38320 36377 38400 36400
rect 38320 36343 38343 36377
rect 38377 36343 38400 36377
rect 38320 36057 38400 36343
rect 38320 36023 38343 36057
rect 38377 36023 38400 36057
rect 38320 35737 38400 36023
rect 38320 35703 38343 35737
rect 38377 35703 38400 35737
rect 38320 35417 38400 35703
rect 38320 35383 38343 35417
rect 38377 35383 38400 35417
rect 38320 35097 38400 35383
rect 38320 35063 38343 35097
rect 38377 35063 38400 35097
rect 38320 34777 38400 35063
rect 38320 34743 38343 34777
rect 38377 34743 38400 34777
rect 38320 34457 38400 34743
rect 38320 34423 38343 34457
rect 38377 34423 38400 34457
rect 38320 34400 38400 34423
rect 38480 36377 38560 36400
rect 38480 36343 38503 36377
rect 38537 36343 38560 36377
rect 38480 36057 38560 36343
rect 38480 36023 38503 36057
rect 38537 36023 38560 36057
rect 38480 35737 38560 36023
rect 38480 35703 38503 35737
rect 38537 35703 38560 35737
rect 38480 35417 38560 35703
rect 38480 35383 38503 35417
rect 38537 35383 38560 35417
rect 38480 35097 38560 35383
rect 38480 35063 38503 35097
rect 38537 35063 38560 35097
rect 38480 34777 38560 35063
rect 38480 34743 38503 34777
rect 38537 34743 38560 34777
rect 38480 34457 38560 34743
rect 38480 34423 38503 34457
rect 38537 34423 38560 34457
rect 38480 34400 38560 34423
rect 38640 36377 38720 36400
rect 38640 36343 38663 36377
rect 38697 36343 38720 36377
rect 38640 36057 38720 36343
rect 38640 36023 38663 36057
rect 38697 36023 38720 36057
rect 38640 35737 38720 36023
rect 38640 35703 38663 35737
rect 38697 35703 38720 35737
rect 38640 35417 38720 35703
rect 38640 35383 38663 35417
rect 38697 35383 38720 35417
rect 38640 35097 38720 35383
rect 38640 35063 38663 35097
rect 38697 35063 38720 35097
rect 38640 34777 38720 35063
rect 38640 34743 38663 34777
rect 38697 34743 38720 34777
rect 38640 34457 38720 34743
rect 38640 34423 38663 34457
rect 38697 34423 38720 34457
rect 38640 34400 38720 34423
rect 38800 36377 38880 36400
rect 38800 36343 38823 36377
rect 38857 36343 38880 36377
rect 38800 36057 38880 36343
rect 38800 36023 38823 36057
rect 38857 36023 38880 36057
rect 38800 35737 38880 36023
rect 38800 35703 38823 35737
rect 38857 35703 38880 35737
rect 38800 35417 38880 35703
rect 38800 35383 38823 35417
rect 38857 35383 38880 35417
rect 38800 35097 38880 35383
rect 38800 35063 38823 35097
rect 38857 35063 38880 35097
rect 38800 34777 38880 35063
rect 38800 34743 38823 34777
rect 38857 34743 38880 34777
rect 38800 34457 38880 34743
rect 38800 34423 38823 34457
rect 38857 34423 38880 34457
rect 38800 34400 38880 34423
rect 38960 36377 39040 36400
rect 38960 36343 38983 36377
rect 39017 36343 39040 36377
rect 38960 36057 39040 36343
rect 38960 36023 38983 36057
rect 39017 36023 39040 36057
rect 38960 35737 39040 36023
rect 38960 35703 38983 35737
rect 39017 35703 39040 35737
rect 38960 35417 39040 35703
rect 38960 35383 38983 35417
rect 39017 35383 39040 35417
rect 38960 35097 39040 35383
rect 38960 35063 38983 35097
rect 39017 35063 39040 35097
rect 38960 34777 39040 35063
rect 38960 34743 38983 34777
rect 39017 34743 39040 34777
rect 38960 34457 39040 34743
rect 38960 34423 38983 34457
rect 39017 34423 39040 34457
rect 38960 34400 39040 34423
rect 39120 36377 39200 36400
rect 39120 36343 39143 36377
rect 39177 36343 39200 36377
rect 39120 36057 39200 36343
rect 39120 36023 39143 36057
rect 39177 36023 39200 36057
rect 39120 35737 39200 36023
rect 39120 35703 39143 35737
rect 39177 35703 39200 35737
rect 39120 35417 39200 35703
rect 39120 35383 39143 35417
rect 39177 35383 39200 35417
rect 39120 35097 39200 35383
rect 39120 35063 39143 35097
rect 39177 35063 39200 35097
rect 39120 34777 39200 35063
rect 39120 34743 39143 34777
rect 39177 34743 39200 34777
rect 39120 34457 39200 34743
rect 39120 34423 39143 34457
rect 39177 34423 39200 34457
rect 39120 34400 39200 34423
rect 39280 36377 39360 36400
rect 39280 36343 39303 36377
rect 39337 36343 39360 36377
rect 39280 36057 39360 36343
rect 39280 36023 39303 36057
rect 39337 36023 39360 36057
rect 39280 35737 39360 36023
rect 39280 35703 39303 35737
rect 39337 35703 39360 35737
rect 39280 35417 39360 35703
rect 39280 35383 39303 35417
rect 39337 35383 39360 35417
rect 39280 35097 39360 35383
rect 39280 35063 39303 35097
rect 39337 35063 39360 35097
rect 39280 34777 39360 35063
rect 39280 34743 39303 34777
rect 39337 34743 39360 34777
rect 39280 34457 39360 34743
rect 39280 34423 39303 34457
rect 39337 34423 39360 34457
rect 39280 34400 39360 34423
rect 39440 36377 39520 36400
rect 39440 36343 39463 36377
rect 39497 36343 39520 36377
rect 39440 36057 39520 36343
rect 39440 36023 39463 36057
rect 39497 36023 39520 36057
rect 39440 35737 39520 36023
rect 39440 35703 39463 35737
rect 39497 35703 39520 35737
rect 39440 35417 39520 35703
rect 39440 35383 39463 35417
rect 39497 35383 39520 35417
rect 39440 35097 39520 35383
rect 39440 35063 39463 35097
rect 39497 35063 39520 35097
rect 39440 34777 39520 35063
rect 39440 34743 39463 34777
rect 39497 34743 39520 34777
rect 39440 34457 39520 34743
rect 39440 34423 39463 34457
rect 39497 34423 39520 34457
rect 39440 34400 39520 34423
rect 39600 36377 39680 36400
rect 39600 36343 39623 36377
rect 39657 36343 39680 36377
rect 39600 36057 39680 36343
rect 39600 36023 39623 36057
rect 39657 36023 39680 36057
rect 39600 35737 39680 36023
rect 39600 35703 39623 35737
rect 39657 35703 39680 35737
rect 39600 35417 39680 35703
rect 39600 35383 39623 35417
rect 39657 35383 39680 35417
rect 39600 35097 39680 35383
rect 39600 35063 39623 35097
rect 39657 35063 39680 35097
rect 39600 34777 39680 35063
rect 39600 34743 39623 34777
rect 39657 34743 39680 34777
rect 39600 34457 39680 34743
rect 39600 34423 39623 34457
rect 39657 34423 39680 34457
rect 39600 34400 39680 34423
rect 39760 36377 39840 36400
rect 39760 36343 39783 36377
rect 39817 36343 39840 36377
rect 39760 36057 39840 36343
rect 39760 36023 39783 36057
rect 39817 36023 39840 36057
rect 39760 35737 39840 36023
rect 39760 35703 39783 35737
rect 39817 35703 39840 35737
rect 39760 35417 39840 35703
rect 39760 35383 39783 35417
rect 39817 35383 39840 35417
rect 39760 35097 39840 35383
rect 39760 35063 39783 35097
rect 39817 35063 39840 35097
rect 39760 34777 39840 35063
rect 39760 34743 39783 34777
rect 39817 34743 39840 34777
rect 39760 34457 39840 34743
rect 39760 34423 39783 34457
rect 39817 34423 39840 34457
rect 39760 34400 39840 34423
rect 39920 36377 40000 36400
rect 39920 36343 39943 36377
rect 39977 36343 40000 36377
rect 39920 36057 40000 36343
rect 39920 36023 39943 36057
rect 39977 36023 40000 36057
rect 39920 35737 40000 36023
rect 39920 35703 39943 35737
rect 39977 35703 40000 35737
rect 39920 35417 40000 35703
rect 39920 35383 39943 35417
rect 39977 35383 40000 35417
rect 39920 35097 40000 35383
rect 39920 35063 39943 35097
rect 39977 35063 40000 35097
rect 39920 34777 40000 35063
rect 39920 34743 39943 34777
rect 39977 34743 40000 34777
rect 39920 34457 40000 34743
rect 39920 34423 39943 34457
rect 39977 34423 40000 34457
rect 39920 34400 40000 34423
rect 40080 36377 40160 36400
rect 40080 36343 40103 36377
rect 40137 36343 40160 36377
rect 40080 36057 40160 36343
rect 40080 36023 40103 36057
rect 40137 36023 40160 36057
rect 40080 35737 40160 36023
rect 40080 35703 40103 35737
rect 40137 35703 40160 35737
rect 40080 35417 40160 35703
rect 40080 35383 40103 35417
rect 40137 35383 40160 35417
rect 40080 35097 40160 35383
rect 40080 35063 40103 35097
rect 40137 35063 40160 35097
rect 40080 34777 40160 35063
rect 40080 34743 40103 34777
rect 40137 34743 40160 34777
rect 40080 34457 40160 34743
rect 40080 34423 40103 34457
rect 40137 34423 40160 34457
rect 40080 34400 40160 34423
rect 40240 36377 40320 36400
rect 40240 36343 40263 36377
rect 40297 36343 40320 36377
rect 40240 36057 40320 36343
rect 40240 36023 40263 36057
rect 40297 36023 40320 36057
rect 40240 35737 40320 36023
rect 40240 35703 40263 35737
rect 40297 35703 40320 35737
rect 40240 35417 40320 35703
rect 40240 35383 40263 35417
rect 40297 35383 40320 35417
rect 40240 35097 40320 35383
rect 40240 35063 40263 35097
rect 40297 35063 40320 35097
rect 40240 34777 40320 35063
rect 40240 34743 40263 34777
rect 40297 34743 40320 34777
rect 40240 34457 40320 34743
rect 40240 34423 40263 34457
rect 40297 34423 40320 34457
rect 40240 34400 40320 34423
rect 40400 36377 40480 36400
rect 40400 36343 40423 36377
rect 40457 36343 40480 36377
rect 40400 36057 40480 36343
rect 40400 36023 40423 36057
rect 40457 36023 40480 36057
rect 40400 35737 40480 36023
rect 40400 35703 40423 35737
rect 40457 35703 40480 35737
rect 40400 35417 40480 35703
rect 40400 35383 40423 35417
rect 40457 35383 40480 35417
rect 40400 35097 40480 35383
rect 40400 35063 40423 35097
rect 40457 35063 40480 35097
rect 40400 34777 40480 35063
rect 40400 34743 40423 34777
rect 40457 34743 40480 34777
rect 40400 34457 40480 34743
rect 40400 34423 40423 34457
rect 40457 34423 40480 34457
rect 40400 34400 40480 34423
rect 40560 36377 40640 36400
rect 40560 36343 40583 36377
rect 40617 36343 40640 36377
rect 40560 36057 40640 36343
rect 40560 36023 40583 36057
rect 40617 36023 40640 36057
rect 40560 35737 40640 36023
rect 40560 35703 40583 35737
rect 40617 35703 40640 35737
rect 40560 35417 40640 35703
rect 40560 35383 40583 35417
rect 40617 35383 40640 35417
rect 40560 35097 40640 35383
rect 40560 35063 40583 35097
rect 40617 35063 40640 35097
rect 40560 34777 40640 35063
rect 40560 34743 40583 34777
rect 40617 34743 40640 34777
rect 40560 34457 40640 34743
rect 40560 34423 40583 34457
rect 40617 34423 40640 34457
rect 40560 34400 40640 34423
rect 40720 36377 40800 36400
rect 40720 36343 40743 36377
rect 40777 36343 40800 36377
rect 40720 36057 40800 36343
rect 40720 36023 40743 36057
rect 40777 36023 40800 36057
rect 40720 35737 40800 36023
rect 40720 35703 40743 35737
rect 40777 35703 40800 35737
rect 40720 35417 40800 35703
rect 40720 35383 40743 35417
rect 40777 35383 40800 35417
rect 40720 35097 40800 35383
rect 40720 35063 40743 35097
rect 40777 35063 40800 35097
rect 40720 34777 40800 35063
rect 40720 34743 40743 34777
rect 40777 34743 40800 34777
rect 40720 34457 40800 34743
rect 40720 34423 40743 34457
rect 40777 34423 40800 34457
rect 40720 34400 40800 34423
rect 40880 36377 40960 36400
rect 40880 36343 40903 36377
rect 40937 36343 40960 36377
rect 40880 36057 40960 36343
rect 40880 36023 40903 36057
rect 40937 36023 40960 36057
rect 40880 35737 40960 36023
rect 40880 35703 40903 35737
rect 40937 35703 40960 35737
rect 40880 35417 40960 35703
rect 40880 35383 40903 35417
rect 40937 35383 40960 35417
rect 40880 35097 40960 35383
rect 40880 35063 40903 35097
rect 40937 35063 40960 35097
rect 40880 34777 40960 35063
rect 40880 34743 40903 34777
rect 40937 34743 40960 34777
rect 40880 34457 40960 34743
rect 40880 34423 40903 34457
rect 40937 34423 40960 34457
rect 40880 34400 40960 34423
rect 41040 36377 41120 36400
rect 41040 36343 41063 36377
rect 41097 36343 41120 36377
rect 41040 36057 41120 36343
rect 41040 36023 41063 36057
rect 41097 36023 41120 36057
rect 41040 35737 41120 36023
rect 41040 35703 41063 35737
rect 41097 35703 41120 35737
rect 41040 35417 41120 35703
rect 41040 35383 41063 35417
rect 41097 35383 41120 35417
rect 41040 35097 41120 35383
rect 41040 35063 41063 35097
rect 41097 35063 41120 35097
rect 41040 34777 41120 35063
rect 41040 34743 41063 34777
rect 41097 34743 41120 34777
rect 41040 34457 41120 34743
rect 41040 34423 41063 34457
rect 41097 34423 41120 34457
rect 41040 34400 41120 34423
rect 41200 36377 41280 36400
rect 41200 36343 41223 36377
rect 41257 36343 41280 36377
rect 41200 36057 41280 36343
rect 41200 36023 41223 36057
rect 41257 36023 41280 36057
rect 41200 35737 41280 36023
rect 41200 35703 41223 35737
rect 41257 35703 41280 35737
rect 41200 35417 41280 35703
rect 41200 35383 41223 35417
rect 41257 35383 41280 35417
rect 41200 35097 41280 35383
rect 41200 35063 41223 35097
rect 41257 35063 41280 35097
rect 41200 34777 41280 35063
rect 41200 34743 41223 34777
rect 41257 34743 41280 34777
rect 41200 34457 41280 34743
rect 41200 34423 41223 34457
rect 41257 34423 41280 34457
rect 41200 34400 41280 34423
rect 41360 36377 41440 36400
rect 41360 36343 41383 36377
rect 41417 36343 41440 36377
rect 41360 36057 41440 36343
rect 41360 36023 41383 36057
rect 41417 36023 41440 36057
rect 41360 35737 41440 36023
rect 41360 35703 41383 35737
rect 41417 35703 41440 35737
rect 41360 35417 41440 35703
rect 41360 35383 41383 35417
rect 41417 35383 41440 35417
rect 41360 35097 41440 35383
rect 41360 35063 41383 35097
rect 41417 35063 41440 35097
rect 41360 34777 41440 35063
rect 41360 34743 41383 34777
rect 41417 34743 41440 34777
rect 41360 34457 41440 34743
rect 41360 34423 41383 34457
rect 41417 34423 41440 34457
rect 41360 34400 41440 34423
rect 41520 36377 41600 36400
rect 41520 36343 41543 36377
rect 41577 36343 41600 36377
rect 41520 36057 41600 36343
rect 41520 36023 41543 36057
rect 41577 36023 41600 36057
rect 41520 35737 41600 36023
rect 41520 35703 41543 35737
rect 41577 35703 41600 35737
rect 41520 35417 41600 35703
rect 41520 35383 41543 35417
rect 41577 35383 41600 35417
rect 41520 35097 41600 35383
rect 41520 35063 41543 35097
rect 41577 35063 41600 35097
rect 41520 34777 41600 35063
rect 41520 34743 41543 34777
rect 41577 34743 41600 34777
rect 41520 34457 41600 34743
rect 41520 34423 41543 34457
rect 41577 34423 41600 34457
rect 41520 34400 41600 34423
rect 41680 36377 41760 36400
rect 41680 36343 41703 36377
rect 41737 36343 41760 36377
rect 41680 36057 41760 36343
rect 41680 36023 41703 36057
rect 41737 36023 41760 36057
rect 41680 35737 41760 36023
rect 41680 35703 41703 35737
rect 41737 35703 41760 35737
rect 41680 35417 41760 35703
rect 41680 35383 41703 35417
rect 41737 35383 41760 35417
rect 41680 35097 41760 35383
rect 41680 35063 41703 35097
rect 41737 35063 41760 35097
rect 41680 34777 41760 35063
rect 41680 34743 41703 34777
rect 41737 34743 41760 34777
rect 41680 34457 41760 34743
rect 41680 34423 41703 34457
rect 41737 34423 41760 34457
rect 41680 34400 41760 34423
rect 41840 36377 41920 36400
rect 41840 36343 41863 36377
rect 41897 36343 41920 36377
rect 41840 36057 41920 36343
rect 41840 36023 41863 36057
rect 41897 36023 41920 36057
rect 41840 35737 41920 36023
rect 41840 35703 41863 35737
rect 41897 35703 41920 35737
rect 41840 35417 41920 35703
rect 41840 35383 41863 35417
rect 41897 35383 41920 35417
rect 41840 35097 41920 35383
rect 41840 35063 41863 35097
rect 41897 35063 41920 35097
rect 41840 34777 41920 35063
rect 41840 34743 41863 34777
rect 41897 34743 41920 34777
rect 41840 34457 41920 34743
rect 41840 34423 41863 34457
rect 41897 34423 41920 34457
rect 41840 34400 41920 34423
rect 0 34297 80 34320
rect 0 34263 23 34297
rect 57 34263 80 34297
rect 0 33977 80 34263
rect 0 33943 23 33977
rect 57 33943 80 33977
rect 0 33920 80 33943
rect 160 34297 240 34320
rect 160 34263 183 34297
rect 217 34263 240 34297
rect 160 33977 240 34263
rect 160 33943 183 33977
rect 217 33943 240 33977
rect 160 33920 240 33943
rect 320 34297 400 34320
rect 320 34263 343 34297
rect 377 34263 400 34297
rect 320 33977 400 34263
rect 320 33943 343 33977
rect 377 33943 400 33977
rect 320 33920 400 33943
rect 480 34297 560 34320
rect 480 34263 503 34297
rect 537 34263 560 34297
rect 480 33977 560 34263
rect 480 33943 503 33977
rect 537 33943 560 33977
rect 480 33920 560 33943
rect 640 34297 720 34320
rect 640 34263 663 34297
rect 697 34263 720 34297
rect 640 33977 720 34263
rect 640 33943 663 33977
rect 697 33943 720 33977
rect 640 33920 720 33943
rect 800 34297 880 34320
rect 800 34263 823 34297
rect 857 34263 880 34297
rect 800 33977 880 34263
rect 800 33943 823 33977
rect 857 33943 880 33977
rect 800 33920 880 33943
rect 960 34297 1040 34320
rect 960 34263 983 34297
rect 1017 34263 1040 34297
rect 960 33977 1040 34263
rect 960 33943 983 33977
rect 1017 33943 1040 33977
rect 960 33920 1040 33943
rect 1120 34297 1200 34320
rect 1120 34263 1143 34297
rect 1177 34263 1200 34297
rect 1120 33977 1200 34263
rect 1120 33943 1143 33977
rect 1177 33943 1200 33977
rect 1120 33920 1200 33943
rect 1280 34297 1360 34320
rect 1280 34263 1303 34297
rect 1337 34263 1360 34297
rect 1280 33977 1360 34263
rect 1280 33943 1303 33977
rect 1337 33943 1360 33977
rect 1280 33920 1360 33943
rect 1440 34297 1520 34320
rect 1440 34263 1463 34297
rect 1497 34263 1520 34297
rect 1440 33977 1520 34263
rect 1440 33943 1463 33977
rect 1497 33943 1520 33977
rect 1440 33920 1520 33943
rect 1600 34297 1680 34320
rect 1600 34263 1623 34297
rect 1657 34263 1680 34297
rect 1600 33977 1680 34263
rect 1600 33943 1623 33977
rect 1657 33943 1680 33977
rect 1600 33920 1680 33943
rect 1760 34297 1840 34320
rect 1760 34263 1783 34297
rect 1817 34263 1840 34297
rect 1760 33977 1840 34263
rect 1760 33943 1783 33977
rect 1817 33943 1840 33977
rect 1760 33920 1840 33943
rect 1920 34297 2000 34320
rect 1920 34263 1943 34297
rect 1977 34263 2000 34297
rect 1920 33977 2000 34263
rect 1920 33943 1943 33977
rect 1977 33943 2000 33977
rect 1920 33920 2000 33943
rect 2080 34297 2160 34320
rect 2080 34263 2103 34297
rect 2137 34263 2160 34297
rect 2080 33977 2160 34263
rect 2080 33943 2103 33977
rect 2137 33943 2160 33977
rect 2080 33920 2160 33943
rect 2240 34297 2320 34320
rect 2240 34263 2263 34297
rect 2297 34263 2320 34297
rect 2240 33977 2320 34263
rect 2240 33943 2263 33977
rect 2297 33943 2320 33977
rect 2240 33920 2320 33943
rect 2400 34297 2480 34320
rect 2400 34263 2423 34297
rect 2457 34263 2480 34297
rect 2400 33977 2480 34263
rect 2400 33943 2423 33977
rect 2457 33943 2480 33977
rect 2400 33920 2480 33943
rect 2560 34297 2640 34320
rect 2560 34263 2583 34297
rect 2617 34263 2640 34297
rect 2560 33977 2640 34263
rect 2560 33943 2583 33977
rect 2617 33943 2640 33977
rect 2560 33920 2640 33943
rect 2720 34297 2800 34320
rect 2720 34263 2743 34297
rect 2777 34263 2800 34297
rect 2720 33977 2800 34263
rect 2720 33943 2743 33977
rect 2777 33943 2800 33977
rect 2720 33920 2800 33943
rect 2880 34297 2960 34320
rect 2880 34263 2903 34297
rect 2937 34263 2960 34297
rect 2880 33977 2960 34263
rect 2880 33943 2903 33977
rect 2937 33943 2960 33977
rect 2880 33920 2960 33943
rect 3040 34297 3120 34320
rect 3040 34263 3063 34297
rect 3097 34263 3120 34297
rect 3040 33977 3120 34263
rect 3040 33943 3063 33977
rect 3097 33943 3120 33977
rect 3040 33920 3120 33943
rect 3200 34297 3280 34320
rect 3200 34263 3223 34297
rect 3257 34263 3280 34297
rect 3200 33977 3280 34263
rect 3200 33943 3223 33977
rect 3257 33943 3280 33977
rect 3200 33920 3280 33943
rect 3360 34297 3440 34320
rect 3360 34263 3383 34297
rect 3417 34263 3440 34297
rect 3360 33977 3440 34263
rect 3360 33943 3383 33977
rect 3417 33943 3440 33977
rect 3360 33920 3440 33943
rect 3520 34297 3600 34320
rect 3520 34263 3543 34297
rect 3577 34263 3600 34297
rect 3520 33977 3600 34263
rect 3520 33943 3543 33977
rect 3577 33943 3600 33977
rect 3520 33920 3600 33943
rect 3680 34297 3760 34320
rect 3680 34263 3703 34297
rect 3737 34263 3760 34297
rect 3680 33977 3760 34263
rect 3680 33943 3703 33977
rect 3737 33943 3760 33977
rect 3680 33920 3760 33943
rect 3840 34297 3920 34320
rect 3840 34263 3863 34297
rect 3897 34263 3920 34297
rect 3840 33977 3920 34263
rect 3840 33943 3863 33977
rect 3897 33943 3920 33977
rect 3840 33920 3920 33943
rect 4000 34297 4080 34320
rect 4000 34263 4023 34297
rect 4057 34263 4080 34297
rect 4000 33977 4080 34263
rect 4000 33943 4023 33977
rect 4057 33943 4080 33977
rect 4000 33920 4080 33943
rect 4160 34297 4240 34320
rect 4160 34263 4183 34297
rect 4217 34263 4240 34297
rect 4160 33977 4240 34263
rect 4160 33943 4183 33977
rect 4217 33943 4240 33977
rect 4160 33920 4240 33943
rect 4320 34297 4400 34320
rect 4320 34263 4343 34297
rect 4377 34263 4400 34297
rect 4320 33977 4400 34263
rect 4320 33943 4343 33977
rect 4377 33943 4400 33977
rect 4320 33920 4400 33943
rect 4480 34297 4560 34320
rect 4480 34263 4503 34297
rect 4537 34263 4560 34297
rect 4480 33977 4560 34263
rect 4480 33943 4503 33977
rect 4537 33943 4560 33977
rect 4480 33920 4560 33943
rect 4640 34297 4720 34320
rect 4640 34263 4663 34297
rect 4697 34263 4720 34297
rect 4640 33977 4720 34263
rect 4640 33943 4663 33977
rect 4697 33943 4720 33977
rect 4640 33920 4720 33943
rect 4800 34297 4880 34320
rect 4800 34263 4823 34297
rect 4857 34263 4880 34297
rect 4800 33977 4880 34263
rect 4800 33943 4823 33977
rect 4857 33943 4880 33977
rect 4800 33920 4880 33943
rect 4960 34297 5040 34320
rect 4960 34263 4983 34297
rect 5017 34263 5040 34297
rect 4960 33977 5040 34263
rect 4960 33943 4983 33977
rect 5017 33943 5040 33977
rect 4960 33920 5040 33943
rect 5120 34297 5200 34320
rect 5120 34263 5143 34297
rect 5177 34263 5200 34297
rect 5120 33977 5200 34263
rect 5120 33943 5143 33977
rect 5177 33943 5200 33977
rect 5120 33920 5200 33943
rect 5280 34297 5360 34320
rect 5280 34263 5303 34297
rect 5337 34263 5360 34297
rect 5280 33977 5360 34263
rect 5280 33943 5303 33977
rect 5337 33943 5360 33977
rect 5280 33920 5360 33943
rect 5440 34297 5520 34320
rect 5440 34263 5463 34297
rect 5497 34263 5520 34297
rect 5440 33977 5520 34263
rect 5440 33943 5463 33977
rect 5497 33943 5520 33977
rect 5440 33920 5520 33943
rect 5600 34297 5680 34320
rect 5600 34263 5623 34297
rect 5657 34263 5680 34297
rect 5600 33977 5680 34263
rect 5600 33943 5623 33977
rect 5657 33943 5680 33977
rect 5600 33920 5680 33943
rect 5760 34297 5840 34320
rect 5760 34263 5783 34297
rect 5817 34263 5840 34297
rect 5760 33977 5840 34263
rect 5760 33943 5783 33977
rect 5817 33943 5840 33977
rect 5760 33920 5840 33943
rect 5920 34297 6000 34320
rect 5920 34263 5943 34297
rect 5977 34263 6000 34297
rect 5920 33977 6000 34263
rect 5920 33943 5943 33977
rect 5977 33943 6000 33977
rect 5920 33920 6000 33943
rect 6080 34297 6160 34320
rect 6080 34263 6103 34297
rect 6137 34263 6160 34297
rect 6080 33977 6160 34263
rect 6080 33943 6103 33977
rect 6137 33943 6160 33977
rect 6080 33920 6160 33943
rect 6240 34297 6320 34320
rect 6240 34263 6263 34297
rect 6297 34263 6320 34297
rect 6240 33977 6320 34263
rect 6240 33943 6263 33977
rect 6297 33943 6320 33977
rect 6240 33920 6320 33943
rect 6400 34297 6480 34320
rect 6400 34263 6423 34297
rect 6457 34263 6480 34297
rect 6400 33977 6480 34263
rect 6400 33943 6423 33977
rect 6457 33943 6480 33977
rect 6400 33920 6480 33943
rect 6560 34297 6640 34320
rect 6560 34263 6583 34297
rect 6617 34263 6640 34297
rect 6560 33977 6640 34263
rect 6560 33943 6583 33977
rect 6617 33943 6640 33977
rect 6560 33920 6640 33943
rect 6720 34297 6800 34320
rect 6720 34263 6743 34297
rect 6777 34263 6800 34297
rect 6720 33977 6800 34263
rect 6720 33943 6743 33977
rect 6777 33943 6800 33977
rect 6720 33920 6800 33943
rect 6880 34297 6960 34320
rect 6880 34263 6903 34297
rect 6937 34263 6960 34297
rect 6880 33977 6960 34263
rect 6880 33943 6903 33977
rect 6937 33943 6960 33977
rect 6880 33920 6960 33943
rect 7040 34297 7120 34320
rect 7040 34263 7063 34297
rect 7097 34263 7120 34297
rect 7040 33977 7120 34263
rect 7040 33943 7063 33977
rect 7097 33943 7120 33977
rect 7040 33920 7120 33943
rect 7200 34297 7280 34320
rect 7200 34263 7223 34297
rect 7257 34263 7280 34297
rect 7200 33977 7280 34263
rect 7200 33943 7223 33977
rect 7257 33943 7280 33977
rect 7200 33920 7280 33943
rect 7360 34297 7440 34320
rect 7360 34263 7383 34297
rect 7417 34263 7440 34297
rect 7360 33977 7440 34263
rect 7360 33943 7383 33977
rect 7417 33943 7440 33977
rect 7360 33920 7440 33943
rect 7520 34297 7600 34320
rect 7520 34263 7543 34297
rect 7577 34263 7600 34297
rect 7520 33977 7600 34263
rect 7520 33943 7543 33977
rect 7577 33943 7600 33977
rect 7520 33920 7600 33943
rect 7680 34297 7760 34320
rect 7680 34263 7703 34297
rect 7737 34263 7760 34297
rect 7680 33977 7760 34263
rect 7680 33943 7703 33977
rect 7737 33943 7760 33977
rect 7680 33920 7760 33943
rect 7840 34297 7920 34320
rect 7840 34263 7863 34297
rect 7897 34263 7920 34297
rect 7840 33977 7920 34263
rect 7840 33943 7863 33977
rect 7897 33943 7920 33977
rect 7840 33920 7920 33943
rect 8000 34297 8080 34320
rect 8000 34263 8023 34297
rect 8057 34263 8080 34297
rect 8000 33977 8080 34263
rect 8000 33943 8023 33977
rect 8057 33943 8080 33977
rect 8000 33920 8080 33943
rect 8160 34297 8240 34320
rect 8160 34263 8183 34297
rect 8217 34263 8240 34297
rect 8160 33977 8240 34263
rect 8160 33943 8183 33977
rect 8217 33943 8240 33977
rect 8160 33920 8240 33943
rect 8320 34297 8400 34320
rect 8320 34263 8343 34297
rect 8377 34263 8400 34297
rect 8320 33977 8400 34263
rect 8320 33943 8343 33977
rect 8377 33943 8400 33977
rect 8320 33920 8400 33943
rect 8480 33920 8560 34320
rect 8640 33920 8720 34320
rect 8800 33920 8880 34320
rect 8960 33920 9040 34320
rect 9120 33920 9200 34320
rect 9280 33920 9360 34320
rect 9440 33920 9520 34320
rect 9600 33920 9680 34320
rect 9760 33920 9840 34320
rect 9920 33920 10000 34320
rect 10080 33920 10160 34320
rect 10240 33920 10320 34320
rect 10400 33920 10480 34320
rect 10560 33920 10640 34320
rect 10720 33920 10800 34320
rect 10880 33920 10960 34320
rect 11040 33920 11120 34320
rect 11200 33920 11280 34320
rect 11360 33920 11440 34320
rect 11520 33920 11600 34320
rect 11680 33920 11760 34320
rect 11840 33920 11920 34320
rect 12000 33920 12080 34320
rect 12160 33920 12240 34320
rect 12320 33920 12400 34320
rect 12480 34297 12560 34320
rect 12480 34263 12503 34297
rect 12537 34263 12560 34297
rect 12480 33977 12560 34263
rect 12480 33943 12503 33977
rect 12537 33943 12560 33977
rect 12480 33920 12560 33943
rect 12640 34297 12720 34320
rect 12640 34263 12663 34297
rect 12697 34263 12720 34297
rect 12640 33977 12720 34263
rect 12640 33943 12663 33977
rect 12697 33943 12720 33977
rect 12640 33920 12720 33943
rect 12800 34297 12880 34320
rect 12800 34263 12823 34297
rect 12857 34263 12880 34297
rect 12800 33977 12880 34263
rect 12800 33943 12823 33977
rect 12857 33943 12880 33977
rect 12800 33920 12880 33943
rect 12960 34297 13040 34320
rect 12960 34263 12983 34297
rect 13017 34263 13040 34297
rect 12960 33977 13040 34263
rect 12960 33943 12983 33977
rect 13017 33943 13040 33977
rect 12960 33920 13040 33943
rect 13120 34297 13200 34320
rect 13120 34263 13143 34297
rect 13177 34263 13200 34297
rect 13120 33977 13200 34263
rect 13120 33943 13143 33977
rect 13177 33943 13200 33977
rect 13120 33920 13200 33943
rect 13280 34297 13360 34320
rect 13280 34263 13303 34297
rect 13337 34263 13360 34297
rect 13280 33977 13360 34263
rect 13280 33943 13303 33977
rect 13337 33943 13360 33977
rect 13280 33920 13360 33943
rect 13440 34297 13520 34320
rect 13440 34263 13463 34297
rect 13497 34263 13520 34297
rect 13440 33977 13520 34263
rect 13440 33943 13463 33977
rect 13497 33943 13520 33977
rect 13440 33920 13520 33943
rect 13600 34297 13680 34320
rect 13600 34263 13623 34297
rect 13657 34263 13680 34297
rect 13600 33977 13680 34263
rect 13600 33943 13623 33977
rect 13657 33943 13680 33977
rect 13600 33920 13680 33943
rect 13760 34297 13840 34320
rect 13760 34263 13783 34297
rect 13817 34263 13840 34297
rect 13760 33977 13840 34263
rect 13760 33943 13783 33977
rect 13817 33943 13840 33977
rect 13760 33920 13840 33943
rect 13920 34297 14000 34320
rect 13920 34263 13943 34297
rect 13977 34263 14000 34297
rect 13920 33977 14000 34263
rect 13920 33943 13943 33977
rect 13977 33943 14000 33977
rect 13920 33920 14000 33943
rect 14080 34297 14160 34320
rect 14080 34263 14103 34297
rect 14137 34263 14160 34297
rect 14080 33977 14160 34263
rect 14080 33943 14103 33977
rect 14137 33943 14160 33977
rect 14080 33920 14160 33943
rect 14240 34297 14320 34320
rect 14240 34263 14263 34297
rect 14297 34263 14320 34297
rect 14240 33977 14320 34263
rect 14240 33943 14263 33977
rect 14297 33943 14320 33977
rect 14240 33920 14320 33943
rect 14400 34297 14480 34320
rect 14400 34263 14423 34297
rect 14457 34263 14480 34297
rect 14400 33977 14480 34263
rect 14400 33943 14423 33977
rect 14457 33943 14480 33977
rect 14400 33920 14480 33943
rect 14560 34297 14640 34320
rect 14560 34263 14583 34297
rect 14617 34263 14640 34297
rect 14560 33977 14640 34263
rect 14560 33943 14583 33977
rect 14617 33943 14640 33977
rect 14560 33920 14640 33943
rect 14720 34297 14800 34320
rect 14720 34263 14743 34297
rect 14777 34263 14800 34297
rect 14720 33977 14800 34263
rect 14720 33943 14743 33977
rect 14777 33943 14800 33977
rect 14720 33920 14800 33943
rect 14880 34297 14960 34320
rect 14880 34263 14903 34297
rect 14937 34263 14960 34297
rect 14880 33977 14960 34263
rect 14880 33943 14903 33977
rect 14937 33943 14960 33977
rect 14880 33920 14960 33943
rect 15040 34297 15120 34320
rect 15040 34263 15063 34297
rect 15097 34263 15120 34297
rect 15040 33977 15120 34263
rect 15040 33943 15063 33977
rect 15097 33943 15120 33977
rect 15040 33920 15120 33943
rect 15200 34297 15280 34320
rect 15200 34263 15223 34297
rect 15257 34263 15280 34297
rect 15200 33977 15280 34263
rect 15200 33943 15223 33977
rect 15257 33943 15280 33977
rect 15200 33920 15280 33943
rect 15360 34297 15440 34320
rect 15360 34263 15383 34297
rect 15417 34263 15440 34297
rect 15360 33977 15440 34263
rect 15360 33943 15383 33977
rect 15417 33943 15440 33977
rect 15360 33920 15440 33943
rect 15520 34297 15600 34320
rect 15520 34263 15543 34297
rect 15577 34263 15600 34297
rect 15520 33977 15600 34263
rect 15520 33943 15543 33977
rect 15577 33943 15600 33977
rect 15520 33920 15600 33943
rect 15680 34297 15760 34320
rect 15680 34263 15703 34297
rect 15737 34263 15760 34297
rect 15680 33977 15760 34263
rect 15680 33943 15703 33977
rect 15737 33943 15760 33977
rect 15680 33920 15760 33943
rect 15840 34297 15920 34320
rect 15840 34263 15863 34297
rect 15897 34263 15920 34297
rect 15840 33977 15920 34263
rect 15840 33943 15863 33977
rect 15897 33943 15920 33977
rect 15840 33920 15920 33943
rect 16000 34297 16080 34320
rect 16000 34263 16023 34297
rect 16057 34263 16080 34297
rect 16000 33977 16080 34263
rect 16000 33943 16023 33977
rect 16057 33943 16080 33977
rect 16000 33920 16080 33943
rect 16160 34297 16240 34320
rect 16160 34263 16183 34297
rect 16217 34263 16240 34297
rect 16160 33977 16240 34263
rect 16160 33943 16183 33977
rect 16217 33943 16240 33977
rect 16160 33920 16240 33943
rect 16320 34297 16400 34320
rect 16320 34263 16343 34297
rect 16377 34263 16400 34297
rect 16320 33977 16400 34263
rect 16320 33943 16343 33977
rect 16377 33943 16400 33977
rect 16320 33920 16400 33943
rect 16480 34297 16560 34320
rect 16480 34263 16503 34297
rect 16537 34263 16560 34297
rect 16480 33977 16560 34263
rect 16480 33943 16503 33977
rect 16537 33943 16560 33977
rect 16480 33920 16560 33943
rect 16640 34297 16720 34320
rect 16640 34263 16663 34297
rect 16697 34263 16720 34297
rect 16640 33977 16720 34263
rect 16640 33943 16663 33977
rect 16697 33943 16720 33977
rect 16640 33920 16720 33943
rect 16800 34297 16880 34320
rect 16800 34263 16823 34297
rect 16857 34263 16880 34297
rect 16800 33977 16880 34263
rect 16800 33943 16823 33977
rect 16857 33943 16880 33977
rect 16800 33920 16880 33943
rect 16960 34297 17040 34320
rect 16960 34263 16983 34297
rect 17017 34263 17040 34297
rect 16960 33977 17040 34263
rect 16960 33943 16983 33977
rect 17017 33943 17040 33977
rect 16960 33920 17040 33943
rect 17120 34297 17200 34320
rect 17120 34263 17143 34297
rect 17177 34263 17200 34297
rect 17120 33977 17200 34263
rect 17120 33943 17143 33977
rect 17177 33943 17200 33977
rect 17120 33920 17200 33943
rect 17280 34297 17360 34320
rect 17280 34263 17303 34297
rect 17337 34263 17360 34297
rect 17280 33977 17360 34263
rect 17280 33943 17303 33977
rect 17337 33943 17360 33977
rect 17280 33920 17360 33943
rect 17440 34297 17520 34320
rect 17440 34263 17463 34297
rect 17497 34263 17520 34297
rect 17440 33977 17520 34263
rect 17440 33943 17463 33977
rect 17497 33943 17520 33977
rect 17440 33920 17520 33943
rect 17600 34297 17680 34320
rect 17600 34263 17623 34297
rect 17657 34263 17680 34297
rect 17600 33977 17680 34263
rect 17600 33943 17623 33977
rect 17657 33943 17680 33977
rect 17600 33920 17680 33943
rect 17760 34297 17840 34320
rect 17760 34263 17783 34297
rect 17817 34263 17840 34297
rect 17760 33977 17840 34263
rect 17760 33943 17783 33977
rect 17817 33943 17840 33977
rect 17760 33920 17840 33943
rect 17920 34297 18000 34320
rect 17920 34263 17943 34297
rect 17977 34263 18000 34297
rect 17920 33977 18000 34263
rect 17920 33943 17943 33977
rect 17977 33943 18000 33977
rect 17920 33920 18000 33943
rect 18080 34297 18160 34320
rect 18080 34263 18103 34297
rect 18137 34263 18160 34297
rect 18080 33977 18160 34263
rect 18080 33943 18103 33977
rect 18137 33943 18160 33977
rect 18080 33920 18160 33943
rect 18240 34297 18320 34320
rect 18240 34263 18263 34297
rect 18297 34263 18320 34297
rect 18240 33977 18320 34263
rect 18240 33943 18263 33977
rect 18297 33943 18320 33977
rect 18240 33920 18320 33943
rect 18400 34297 18480 34320
rect 18400 34263 18423 34297
rect 18457 34263 18480 34297
rect 18400 33977 18480 34263
rect 18400 33943 18423 33977
rect 18457 33943 18480 33977
rect 18400 33920 18480 33943
rect 18560 34297 18640 34320
rect 18560 34263 18583 34297
rect 18617 34263 18640 34297
rect 18560 33977 18640 34263
rect 18560 33943 18583 33977
rect 18617 33943 18640 33977
rect 18560 33920 18640 33943
rect 18720 34297 18800 34320
rect 18720 34263 18743 34297
rect 18777 34263 18800 34297
rect 18720 33977 18800 34263
rect 18720 33943 18743 33977
rect 18777 33943 18800 33977
rect 18720 33920 18800 33943
rect 18880 34297 18960 34320
rect 18880 34263 18903 34297
rect 18937 34263 18960 34297
rect 18880 33977 18960 34263
rect 18880 33943 18903 33977
rect 18937 33943 18960 33977
rect 18880 33920 18960 33943
rect 19040 33920 19120 34320
rect 19200 33920 19280 34320
rect 19360 33920 19440 34320
rect 19520 33920 19600 34320
rect 19680 33920 19760 34320
rect 19840 33920 19920 34320
rect 20000 33920 20080 34320
rect 20160 33920 20240 34320
rect 20320 33920 20400 34320
rect 20480 33920 20560 34320
rect 20640 33920 20720 34320
rect 20800 33920 20880 34320
rect 20960 33920 21040 34320
rect 21120 33920 21200 34320
rect 21280 33920 21360 34320
rect 21440 33920 21520 34320
rect 21600 33920 21680 34320
rect 21760 33920 21840 34320
rect 21920 33920 22000 34320
rect 22080 33920 22160 34320
rect 22240 33920 22320 34320
rect 22400 33920 22480 34320
rect 22560 33920 22640 34320
rect 22720 33920 22800 34320
rect 22880 33920 22960 34320
rect 23120 34297 23200 34320
rect 23120 34263 23143 34297
rect 23177 34263 23200 34297
rect 23120 33977 23200 34263
rect 23120 33943 23143 33977
rect 23177 33943 23200 33977
rect 23120 33920 23200 33943
rect 23280 34297 23360 34320
rect 23280 34263 23303 34297
rect 23337 34263 23360 34297
rect 23280 33977 23360 34263
rect 23280 33943 23303 33977
rect 23337 33943 23360 33977
rect 23280 33920 23360 33943
rect 23440 34297 23520 34320
rect 23440 34263 23463 34297
rect 23497 34263 23520 34297
rect 23440 33977 23520 34263
rect 23440 33943 23463 33977
rect 23497 33943 23520 33977
rect 23440 33920 23520 33943
rect 23600 34297 23680 34320
rect 23600 34263 23623 34297
rect 23657 34263 23680 34297
rect 23600 33977 23680 34263
rect 23600 33943 23623 33977
rect 23657 33943 23680 33977
rect 23600 33920 23680 33943
rect 23760 34297 23840 34320
rect 23760 34263 23783 34297
rect 23817 34263 23840 34297
rect 23760 33977 23840 34263
rect 23760 33943 23783 33977
rect 23817 33943 23840 33977
rect 23760 33920 23840 33943
rect 23920 34297 24000 34320
rect 23920 34263 23943 34297
rect 23977 34263 24000 34297
rect 23920 33977 24000 34263
rect 23920 33943 23943 33977
rect 23977 33943 24000 33977
rect 23920 33920 24000 33943
rect 24080 34297 24160 34320
rect 24080 34263 24103 34297
rect 24137 34263 24160 34297
rect 24080 33977 24160 34263
rect 24080 33943 24103 33977
rect 24137 33943 24160 33977
rect 24080 33920 24160 33943
rect 24240 34297 24320 34320
rect 24240 34263 24263 34297
rect 24297 34263 24320 34297
rect 24240 33977 24320 34263
rect 24240 33943 24263 33977
rect 24297 33943 24320 33977
rect 24240 33920 24320 33943
rect 24400 34297 24480 34320
rect 24400 34263 24423 34297
rect 24457 34263 24480 34297
rect 24400 33977 24480 34263
rect 24400 33943 24423 33977
rect 24457 33943 24480 33977
rect 24400 33920 24480 33943
rect 24560 34297 24640 34320
rect 24560 34263 24583 34297
rect 24617 34263 24640 34297
rect 24560 33977 24640 34263
rect 24560 33943 24583 33977
rect 24617 33943 24640 33977
rect 24560 33920 24640 33943
rect 24720 34297 24800 34320
rect 24720 34263 24743 34297
rect 24777 34263 24800 34297
rect 24720 33977 24800 34263
rect 24720 33943 24743 33977
rect 24777 33943 24800 33977
rect 24720 33920 24800 33943
rect 24880 34297 24960 34320
rect 24880 34263 24903 34297
rect 24937 34263 24960 34297
rect 24880 33977 24960 34263
rect 24880 33943 24903 33977
rect 24937 33943 24960 33977
rect 24880 33920 24960 33943
rect 25040 34297 25120 34320
rect 25040 34263 25063 34297
rect 25097 34263 25120 34297
rect 25040 33977 25120 34263
rect 25040 33943 25063 33977
rect 25097 33943 25120 33977
rect 25040 33920 25120 33943
rect 25200 34297 25280 34320
rect 25200 34263 25223 34297
rect 25257 34263 25280 34297
rect 25200 33977 25280 34263
rect 25200 33943 25223 33977
rect 25257 33943 25280 33977
rect 25200 33920 25280 33943
rect 25360 34297 25440 34320
rect 25360 34263 25383 34297
rect 25417 34263 25440 34297
rect 25360 33977 25440 34263
rect 25360 33943 25383 33977
rect 25417 33943 25440 33977
rect 25360 33920 25440 33943
rect 25520 34297 25600 34320
rect 25520 34263 25543 34297
rect 25577 34263 25600 34297
rect 25520 33977 25600 34263
rect 25520 33943 25543 33977
rect 25577 33943 25600 33977
rect 25520 33920 25600 33943
rect 25680 34297 25760 34320
rect 25680 34263 25703 34297
rect 25737 34263 25760 34297
rect 25680 33977 25760 34263
rect 25680 33943 25703 33977
rect 25737 33943 25760 33977
rect 25680 33920 25760 33943
rect 25840 34297 25920 34320
rect 25840 34263 25863 34297
rect 25897 34263 25920 34297
rect 25840 33977 25920 34263
rect 25840 33943 25863 33977
rect 25897 33943 25920 33977
rect 25840 33920 25920 33943
rect 26000 34297 26080 34320
rect 26000 34263 26023 34297
rect 26057 34263 26080 34297
rect 26000 33977 26080 34263
rect 26000 33943 26023 33977
rect 26057 33943 26080 33977
rect 26000 33920 26080 33943
rect 26160 34297 26240 34320
rect 26160 34263 26183 34297
rect 26217 34263 26240 34297
rect 26160 33977 26240 34263
rect 26160 33943 26183 33977
rect 26217 33943 26240 33977
rect 26160 33920 26240 33943
rect 26320 34297 26400 34320
rect 26320 34263 26343 34297
rect 26377 34263 26400 34297
rect 26320 33977 26400 34263
rect 26320 33943 26343 33977
rect 26377 33943 26400 33977
rect 26320 33920 26400 33943
rect 26480 34297 26560 34320
rect 26480 34263 26503 34297
rect 26537 34263 26560 34297
rect 26480 33977 26560 34263
rect 26480 33943 26503 33977
rect 26537 33943 26560 33977
rect 26480 33920 26560 33943
rect 26640 34297 26720 34320
rect 26640 34263 26663 34297
rect 26697 34263 26720 34297
rect 26640 33977 26720 34263
rect 26640 33943 26663 33977
rect 26697 33943 26720 33977
rect 26640 33920 26720 33943
rect 26800 34297 26880 34320
rect 26800 34263 26823 34297
rect 26857 34263 26880 34297
rect 26800 33977 26880 34263
rect 26800 33943 26823 33977
rect 26857 33943 26880 33977
rect 26800 33920 26880 33943
rect 26960 34297 27040 34320
rect 26960 34263 26983 34297
rect 27017 34263 27040 34297
rect 26960 33977 27040 34263
rect 26960 33943 26983 33977
rect 27017 33943 27040 33977
rect 26960 33920 27040 33943
rect 27120 34297 27200 34320
rect 27120 34263 27143 34297
rect 27177 34263 27200 34297
rect 27120 33977 27200 34263
rect 27120 33943 27143 33977
rect 27177 33943 27200 33977
rect 27120 33920 27200 33943
rect 27280 34297 27360 34320
rect 27280 34263 27303 34297
rect 27337 34263 27360 34297
rect 27280 33977 27360 34263
rect 27280 33943 27303 33977
rect 27337 33943 27360 33977
rect 27280 33920 27360 33943
rect 27440 34297 27520 34320
rect 27440 34263 27463 34297
rect 27497 34263 27520 34297
rect 27440 33977 27520 34263
rect 27440 33943 27463 33977
rect 27497 33943 27520 33977
rect 27440 33920 27520 33943
rect 27600 34297 27680 34320
rect 27600 34263 27623 34297
rect 27657 34263 27680 34297
rect 27600 33977 27680 34263
rect 27600 33943 27623 33977
rect 27657 33943 27680 33977
rect 27600 33920 27680 33943
rect 27760 34297 27840 34320
rect 27760 34263 27783 34297
rect 27817 34263 27840 34297
rect 27760 33977 27840 34263
rect 27760 33943 27783 33977
rect 27817 33943 27840 33977
rect 27760 33920 27840 33943
rect 27920 34297 28000 34320
rect 27920 34263 27943 34297
rect 27977 34263 28000 34297
rect 27920 33977 28000 34263
rect 27920 33943 27943 33977
rect 27977 33943 28000 33977
rect 27920 33920 28000 33943
rect 28080 34297 28160 34320
rect 28080 34263 28103 34297
rect 28137 34263 28160 34297
rect 28080 33977 28160 34263
rect 28080 33943 28103 33977
rect 28137 33943 28160 33977
rect 28080 33920 28160 33943
rect 28240 34297 28320 34320
rect 28240 34263 28263 34297
rect 28297 34263 28320 34297
rect 28240 33977 28320 34263
rect 28240 33943 28263 33977
rect 28297 33943 28320 33977
rect 28240 33920 28320 33943
rect 28400 34297 28480 34320
rect 28400 34263 28423 34297
rect 28457 34263 28480 34297
rect 28400 33977 28480 34263
rect 28400 33943 28423 33977
rect 28457 33943 28480 33977
rect 28400 33920 28480 33943
rect 28560 34297 28640 34320
rect 28560 34263 28583 34297
rect 28617 34263 28640 34297
rect 28560 33977 28640 34263
rect 28560 33943 28583 33977
rect 28617 33943 28640 33977
rect 28560 33920 28640 33943
rect 28720 34297 28800 34320
rect 28720 34263 28743 34297
rect 28777 34263 28800 34297
rect 28720 33977 28800 34263
rect 28720 33943 28743 33977
rect 28777 33943 28800 33977
rect 28720 33920 28800 33943
rect 28880 34297 28960 34320
rect 28880 34263 28903 34297
rect 28937 34263 28960 34297
rect 28880 33977 28960 34263
rect 28880 33943 28903 33977
rect 28937 33943 28960 33977
rect 28880 33920 28960 33943
rect 29040 34297 29120 34320
rect 29040 34263 29063 34297
rect 29097 34263 29120 34297
rect 29040 33977 29120 34263
rect 29040 33943 29063 33977
rect 29097 33943 29120 33977
rect 29040 33920 29120 33943
rect 29200 34297 29280 34320
rect 29200 34263 29223 34297
rect 29257 34263 29280 34297
rect 29200 33977 29280 34263
rect 29200 33943 29223 33977
rect 29257 33943 29280 33977
rect 29200 33920 29280 33943
rect 29360 34297 29440 34320
rect 29360 34263 29383 34297
rect 29417 34263 29440 34297
rect 29360 33977 29440 34263
rect 29360 33943 29383 33977
rect 29417 33943 29440 33977
rect 29360 33920 29440 33943
rect 29520 33920 29600 34320
rect 29680 33920 29760 34320
rect 29840 33920 29920 34320
rect 30000 33920 30080 34320
rect 30160 33920 30240 34320
rect 30320 33920 30400 34320
rect 30480 33920 30560 34320
rect 30640 33920 30720 34320
rect 30800 33920 30880 34320
rect 30960 33920 31040 34320
rect 31120 33920 31200 34320
rect 31280 33920 31360 34320
rect 31440 33920 31520 34320
rect 31600 33920 31680 34320
rect 31760 33920 31840 34320
rect 31920 33920 32000 34320
rect 32080 33920 32160 34320
rect 32240 33920 32320 34320
rect 32400 33920 32480 34320
rect 32560 33920 32640 34320
rect 32720 33920 32800 34320
rect 32880 33920 32960 34320
rect 33040 33920 33120 34320
rect 33200 33920 33280 34320
rect 33360 33920 33440 34320
rect 33520 34297 33600 34320
rect 33520 34263 33543 34297
rect 33577 34263 33600 34297
rect 33520 33977 33600 34263
rect 33520 33943 33543 33977
rect 33577 33943 33600 33977
rect 33520 33920 33600 33943
rect 33680 34297 33760 34320
rect 33680 34263 33703 34297
rect 33737 34263 33760 34297
rect 33680 33977 33760 34263
rect 33680 33943 33703 33977
rect 33737 33943 33760 33977
rect 33680 33920 33760 33943
rect 33840 34297 33920 34320
rect 33840 34263 33863 34297
rect 33897 34263 33920 34297
rect 33840 33977 33920 34263
rect 33840 33943 33863 33977
rect 33897 33943 33920 33977
rect 33840 33920 33920 33943
rect 34000 34297 34080 34320
rect 34000 34263 34023 34297
rect 34057 34263 34080 34297
rect 34000 33977 34080 34263
rect 34000 33943 34023 33977
rect 34057 33943 34080 33977
rect 34000 33920 34080 33943
rect 34160 34297 34240 34320
rect 34160 34263 34183 34297
rect 34217 34263 34240 34297
rect 34160 33977 34240 34263
rect 34160 33943 34183 33977
rect 34217 33943 34240 33977
rect 34160 33920 34240 33943
rect 34320 34297 34400 34320
rect 34320 34263 34343 34297
rect 34377 34263 34400 34297
rect 34320 33977 34400 34263
rect 34320 33943 34343 33977
rect 34377 33943 34400 33977
rect 34320 33920 34400 33943
rect 34480 34297 34560 34320
rect 34480 34263 34503 34297
rect 34537 34263 34560 34297
rect 34480 33977 34560 34263
rect 34480 33943 34503 33977
rect 34537 33943 34560 33977
rect 34480 33920 34560 33943
rect 34640 34297 34720 34320
rect 34640 34263 34663 34297
rect 34697 34263 34720 34297
rect 34640 33977 34720 34263
rect 34640 33943 34663 33977
rect 34697 33943 34720 33977
rect 34640 33920 34720 33943
rect 34800 34297 34880 34320
rect 34800 34263 34823 34297
rect 34857 34263 34880 34297
rect 34800 33977 34880 34263
rect 34800 33943 34823 33977
rect 34857 33943 34880 33977
rect 34800 33920 34880 33943
rect 34960 34297 35040 34320
rect 34960 34263 34983 34297
rect 35017 34263 35040 34297
rect 34960 33977 35040 34263
rect 34960 33943 34983 33977
rect 35017 33943 35040 33977
rect 34960 33920 35040 33943
rect 35120 34297 35200 34320
rect 35120 34263 35143 34297
rect 35177 34263 35200 34297
rect 35120 33977 35200 34263
rect 35120 33943 35143 33977
rect 35177 33943 35200 33977
rect 35120 33920 35200 33943
rect 35280 34297 35360 34320
rect 35280 34263 35303 34297
rect 35337 34263 35360 34297
rect 35280 33977 35360 34263
rect 35280 33943 35303 33977
rect 35337 33943 35360 33977
rect 35280 33920 35360 33943
rect 35440 34297 35520 34320
rect 35440 34263 35463 34297
rect 35497 34263 35520 34297
rect 35440 33977 35520 34263
rect 35440 33943 35463 33977
rect 35497 33943 35520 33977
rect 35440 33920 35520 33943
rect 35600 34297 35680 34320
rect 35600 34263 35623 34297
rect 35657 34263 35680 34297
rect 35600 33977 35680 34263
rect 35600 33943 35623 33977
rect 35657 33943 35680 33977
rect 35600 33920 35680 33943
rect 35760 34297 35840 34320
rect 35760 34263 35783 34297
rect 35817 34263 35840 34297
rect 35760 33977 35840 34263
rect 35760 33943 35783 33977
rect 35817 33943 35840 33977
rect 35760 33920 35840 33943
rect 35920 34297 36000 34320
rect 35920 34263 35943 34297
rect 35977 34263 36000 34297
rect 35920 33977 36000 34263
rect 35920 33943 35943 33977
rect 35977 33943 36000 33977
rect 35920 33920 36000 33943
rect 36080 34297 36160 34320
rect 36080 34263 36103 34297
rect 36137 34263 36160 34297
rect 36080 33977 36160 34263
rect 36080 33943 36103 33977
rect 36137 33943 36160 33977
rect 36080 33920 36160 33943
rect 36240 34297 36320 34320
rect 36240 34263 36263 34297
rect 36297 34263 36320 34297
rect 36240 33977 36320 34263
rect 36240 33943 36263 33977
rect 36297 33943 36320 33977
rect 36240 33920 36320 33943
rect 36400 34297 36480 34320
rect 36400 34263 36423 34297
rect 36457 34263 36480 34297
rect 36400 33977 36480 34263
rect 36400 33943 36423 33977
rect 36457 33943 36480 33977
rect 36400 33920 36480 33943
rect 36560 34297 36640 34320
rect 36560 34263 36583 34297
rect 36617 34263 36640 34297
rect 36560 33977 36640 34263
rect 36560 33943 36583 33977
rect 36617 33943 36640 33977
rect 36560 33920 36640 33943
rect 36720 34297 36800 34320
rect 36720 34263 36743 34297
rect 36777 34263 36800 34297
rect 36720 33977 36800 34263
rect 36720 33943 36743 33977
rect 36777 33943 36800 33977
rect 36720 33920 36800 33943
rect 36880 34297 36960 34320
rect 36880 34263 36903 34297
rect 36937 34263 36960 34297
rect 36880 33977 36960 34263
rect 36880 33943 36903 33977
rect 36937 33943 36960 33977
rect 36880 33920 36960 33943
rect 37040 34297 37120 34320
rect 37040 34263 37063 34297
rect 37097 34263 37120 34297
rect 37040 33977 37120 34263
rect 37040 33943 37063 33977
rect 37097 33943 37120 33977
rect 37040 33920 37120 33943
rect 37200 34297 37280 34320
rect 37200 34263 37223 34297
rect 37257 34263 37280 34297
rect 37200 33977 37280 34263
rect 37200 33943 37223 33977
rect 37257 33943 37280 33977
rect 37200 33920 37280 33943
rect 37360 34297 37440 34320
rect 37360 34263 37383 34297
rect 37417 34263 37440 34297
rect 37360 33977 37440 34263
rect 37360 33943 37383 33977
rect 37417 33943 37440 33977
rect 37360 33920 37440 33943
rect 37520 34297 37600 34320
rect 37520 34263 37543 34297
rect 37577 34263 37600 34297
rect 37520 33977 37600 34263
rect 37520 33943 37543 33977
rect 37577 33943 37600 33977
rect 37520 33920 37600 33943
rect 37680 34297 37760 34320
rect 37680 34263 37703 34297
rect 37737 34263 37760 34297
rect 37680 33977 37760 34263
rect 37680 33943 37703 33977
rect 37737 33943 37760 33977
rect 37680 33920 37760 33943
rect 37840 34297 37920 34320
rect 37840 34263 37863 34297
rect 37897 34263 37920 34297
rect 37840 33977 37920 34263
rect 37840 33943 37863 33977
rect 37897 33943 37920 33977
rect 37840 33920 37920 33943
rect 38000 34297 38080 34320
rect 38000 34263 38023 34297
rect 38057 34263 38080 34297
rect 38000 33977 38080 34263
rect 38000 33943 38023 33977
rect 38057 33943 38080 33977
rect 38000 33920 38080 33943
rect 38160 34297 38240 34320
rect 38160 34263 38183 34297
rect 38217 34263 38240 34297
rect 38160 33977 38240 34263
rect 38160 33943 38183 33977
rect 38217 33943 38240 33977
rect 38160 33920 38240 33943
rect 38320 34297 38400 34320
rect 38320 34263 38343 34297
rect 38377 34263 38400 34297
rect 38320 33977 38400 34263
rect 38320 33943 38343 33977
rect 38377 33943 38400 33977
rect 38320 33920 38400 33943
rect 38480 34297 38560 34320
rect 38480 34263 38503 34297
rect 38537 34263 38560 34297
rect 38480 33977 38560 34263
rect 38480 33943 38503 33977
rect 38537 33943 38560 33977
rect 38480 33920 38560 33943
rect 38640 34297 38720 34320
rect 38640 34263 38663 34297
rect 38697 34263 38720 34297
rect 38640 33977 38720 34263
rect 38640 33943 38663 33977
rect 38697 33943 38720 33977
rect 38640 33920 38720 33943
rect 38800 34297 38880 34320
rect 38800 34263 38823 34297
rect 38857 34263 38880 34297
rect 38800 33977 38880 34263
rect 38800 33943 38823 33977
rect 38857 33943 38880 33977
rect 38800 33920 38880 33943
rect 38960 34297 39040 34320
rect 38960 34263 38983 34297
rect 39017 34263 39040 34297
rect 38960 33977 39040 34263
rect 38960 33943 38983 33977
rect 39017 33943 39040 33977
rect 38960 33920 39040 33943
rect 39120 34297 39200 34320
rect 39120 34263 39143 34297
rect 39177 34263 39200 34297
rect 39120 33977 39200 34263
rect 39120 33943 39143 33977
rect 39177 33943 39200 33977
rect 39120 33920 39200 33943
rect 39280 34297 39360 34320
rect 39280 34263 39303 34297
rect 39337 34263 39360 34297
rect 39280 33977 39360 34263
rect 39280 33943 39303 33977
rect 39337 33943 39360 33977
rect 39280 33920 39360 33943
rect 39440 34297 39520 34320
rect 39440 34263 39463 34297
rect 39497 34263 39520 34297
rect 39440 33977 39520 34263
rect 39440 33943 39463 33977
rect 39497 33943 39520 33977
rect 39440 33920 39520 33943
rect 39600 34297 39680 34320
rect 39600 34263 39623 34297
rect 39657 34263 39680 34297
rect 39600 33977 39680 34263
rect 39600 33943 39623 33977
rect 39657 33943 39680 33977
rect 39600 33920 39680 33943
rect 39760 34297 39840 34320
rect 39760 34263 39783 34297
rect 39817 34263 39840 34297
rect 39760 33977 39840 34263
rect 39760 33943 39783 33977
rect 39817 33943 39840 33977
rect 39760 33920 39840 33943
rect 39920 34297 40000 34320
rect 39920 34263 39943 34297
rect 39977 34263 40000 34297
rect 39920 33977 40000 34263
rect 39920 33943 39943 33977
rect 39977 33943 40000 33977
rect 39920 33920 40000 33943
rect 40080 34297 40160 34320
rect 40080 34263 40103 34297
rect 40137 34263 40160 34297
rect 40080 33977 40160 34263
rect 40080 33943 40103 33977
rect 40137 33943 40160 33977
rect 40080 33920 40160 33943
rect 40240 34297 40320 34320
rect 40240 34263 40263 34297
rect 40297 34263 40320 34297
rect 40240 33977 40320 34263
rect 40240 33943 40263 33977
rect 40297 33943 40320 33977
rect 40240 33920 40320 33943
rect 40400 34297 40480 34320
rect 40400 34263 40423 34297
rect 40457 34263 40480 34297
rect 40400 33977 40480 34263
rect 40400 33943 40423 33977
rect 40457 33943 40480 33977
rect 40400 33920 40480 33943
rect 40560 34297 40640 34320
rect 40560 34263 40583 34297
rect 40617 34263 40640 34297
rect 40560 33977 40640 34263
rect 40560 33943 40583 33977
rect 40617 33943 40640 33977
rect 40560 33920 40640 33943
rect 40720 34297 40800 34320
rect 40720 34263 40743 34297
rect 40777 34263 40800 34297
rect 40720 33977 40800 34263
rect 40720 33943 40743 33977
rect 40777 33943 40800 33977
rect 40720 33920 40800 33943
rect 40880 34297 40960 34320
rect 40880 34263 40903 34297
rect 40937 34263 40960 34297
rect 40880 33977 40960 34263
rect 40880 33943 40903 33977
rect 40937 33943 40960 33977
rect 40880 33920 40960 33943
rect 41040 34297 41120 34320
rect 41040 34263 41063 34297
rect 41097 34263 41120 34297
rect 41040 33977 41120 34263
rect 41040 33943 41063 33977
rect 41097 33943 41120 33977
rect 41040 33920 41120 33943
rect 41200 34297 41280 34320
rect 41200 34263 41223 34297
rect 41257 34263 41280 34297
rect 41200 33977 41280 34263
rect 41200 33943 41223 33977
rect 41257 33943 41280 33977
rect 41200 33920 41280 33943
rect 41360 34297 41440 34320
rect 41360 34263 41383 34297
rect 41417 34263 41440 34297
rect 41360 33977 41440 34263
rect 41360 33943 41383 33977
rect 41417 33943 41440 33977
rect 41360 33920 41440 33943
rect 41520 34297 41600 34320
rect 41520 34263 41543 34297
rect 41577 34263 41600 34297
rect 41520 33977 41600 34263
rect 41520 33943 41543 33977
rect 41577 33943 41600 33977
rect 41520 33920 41600 33943
rect 41680 34297 41760 34320
rect 41680 34263 41703 34297
rect 41737 34263 41760 34297
rect 41680 33977 41760 34263
rect 41680 33943 41703 33977
rect 41737 33943 41760 33977
rect 41680 33920 41760 33943
rect 41840 34297 41920 34320
rect 41840 34263 41863 34297
rect 41897 34263 41920 34297
rect 41840 33977 41920 34263
rect 41840 33943 41863 33977
rect 41897 33943 41920 33977
rect 41840 33920 41920 33943
rect 0 33817 80 33840
rect 0 33783 23 33817
rect 57 33783 80 33817
rect 0 33497 80 33783
rect 0 33463 23 33497
rect 57 33463 80 33497
rect 0 33440 80 33463
rect 160 33817 240 33840
rect 160 33783 183 33817
rect 217 33783 240 33817
rect 160 33497 240 33783
rect 160 33463 183 33497
rect 217 33463 240 33497
rect 160 33440 240 33463
rect 320 33817 400 33840
rect 320 33783 343 33817
rect 377 33783 400 33817
rect 320 33497 400 33783
rect 320 33463 343 33497
rect 377 33463 400 33497
rect 320 33440 400 33463
rect 480 33817 560 33840
rect 480 33783 503 33817
rect 537 33783 560 33817
rect 480 33497 560 33783
rect 480 33463 503 33497
rect 537 33463 560 33497
rect 480 33440 560 33463
rect 640 33817 720 33840
rect 640 33783 663 33817
rect 697 33783 720 33817
rect 640 33497 720 33783
rect 640 33463 663 33497
rect 697 33463 720 33497
rect 640 33440 720 33463
rect 800 33817 880 33840
rect 800 33783 823 33817
rect 857 33783 880 33817
rect 800 33497 880 33783
rect 800 33463 823 33497
rect 857 33463 880 33497
rect 800 33440 880 33463
rect 960 33817 1040 33840
rect 960 33783 983 33817
rect 1017 33783 1040 33817
rect 960 33497 1040 33783
rect 960 33463 983 33497
rect 1017 33463 1040 33497
rect 960 33440 1040 33463
rect 1120 33817 1200 33840
rect 1120 33783 1143 33817
rect 1177 33783 1200 33817
rect 1120 33497 1200 33783
rect 1120 33463 1143 33497
rect 1177 33463 1200 33497
rect 1120 33440 1200 33463
rect 1280 33817 1360 33840
rect 1280 33783 1303 33817
rect 1337 33783 1360 33817
rect 1280 33497 1360 33783
rect 1280 33463 1303 33497
rect 1337 33463 1360 33497
rect 1280 33440 1360 33463
rect 1440 33817 1520 33840
rect 1440 33783 1463 33817
rect 1497 33783 1520 33817
rect 1440 33497 1520 33783
rect 1440 33463 1463 33497
rect 1497 33463 1520 33497
rect 1440 33440 1520 33463
rect 1600 33817 1680 33840
rect 1600 33783 1623 33817
rect 1657 33783 1680 33817
rect 1600 33497 1680 33783
rect 1600 33463 1623 33497
rect 1657 33463 1680 33497
rect 1600 33440 1680 33463
rect 1760 33817 1840 33840
rect 1760 33783 1783 33817
rect 1817 33783 1840 33817
rect 1760 33497 1840 33783
rect 1760 33463 1783 33497
rect 1817 33463 1840 33497
rect 1760 33440 1840 33463
rect 1920 33817 2000 33840
rect 1920 33783 1943 33817
rect 1977 33783 2000 33817
rect 1920 33497 2000 33783
rect 1920 33463 1943 33497
rect 1977 33463 2000 33497
rect 1920 33440 2000 33463
rect 2080 33817 2160 33840
rect 2080 33783 2103 33817
rect 2137 33783 2160 33817
rect 2080 33497 2160 33783
rect 2080 33463 2103 33497
rect 2137 33463 2160 33497
rect 2080 33440 2160 33463
rect 2240 33817 2320 33840
rect 2240 33783 2263 33817
rect 2297 33783 2320 33817
rect 2240 33497 2320 33783
rect 2240 33463 2263 33497
rect 2297 33463 2320 33497
rect 2240 33440 2320 33463
rect 2400 33817 2480 33840
rect 2400 33783 2423 33817
rect 2457 33783 2480 33817
rect 2400 33497 2480 33783
rect 2400 33463 2423 33497
rect 2457 33463 2480 33497
rect 2400 33440 2480 33463
rect 2560 33817 2640 33840
rect 2560 33783 2583 33817
rect 2617 33783 2640 33817
rect 2560 33497 2640 33783
rect 2560 33463 2583 33497
rect 2617 33463 2640 33497
rect 2560 33440 2640 33463
rect 2720 33817 2800 33840
rect 2720 33783 2743 33817
rect 2777 33783 2800 33817
rect 2720 33497 2800 33783
rect 2720 33463 2743 33497
rect 2777 33463 2800 33497
rect 2720 33440 2800 33463
rect 2880 33817 2960 33840
rect 2880 33783 2903 33817
rect 2937 33783 2960 33817
rect 2880 33497 2960 33783
rect 2880 33463 2903 33497
rect 2937 33463 2960 33497
rect 2880 33440 2960 33463
rect 3040 33817 3120 33840
rect 3040 33783 3063 33817
rect 3097 33783 3120 33817
rect 3040 33497 3120 33783
rect 3040 33463 3063 33497
rect 3097 33463 3120 33497
rect 3040 33440 3120 33463
rect 3200 33817 3280 33840
rect 3200 33783 3223 33817
rect 3257 33783 3280 33817
rect 3200 33497 3280 33783
rect 3200 33463 3223 33497
rect 3257 33463 3280 33497
rect 3200 33440 3280 33463
rect 3360 33817 3440 33840
rect 3360 33783 3383 33817
rect 3417 33783 3440 33817
rect 3360 33497 3440 33783
rect 3360 33463 3383 33497
rect 3417 33463 3440 33497
rect 3360 33440 3440 33463
rect 3520 33817 3600 33840
rect 3520 33783 3543 33817
rect 3577 33783 3600 33817
rect 3520 33497 3600 33783
rect 3520 33463 3543 33497
rect 3577 33463 3600 33497
rect 3520 33440 3600 33463
rect 3680 33817 3760 33840
rect 3680 33783 3703 33817
rect 3737 33783 3760 33817
rect 3680 33497 3760 33783
rect 3680 33463 3703 33497
rect 3737 33463 3760 33497
rect 3680 33440 3760 33463
rect 3840 33817 3920 33840
rect 3840 33783 3863 33817
rect 3897 33783 3920 33817
rect 3840 33497 3920 33783
rect 3840 33463 3863 33497
rect 3897 33463 3920 33497
rect 3840 33440 3920 33463
rect 4000 33817 4080 33840
rect 4000 33783 4023 33817
rect 4057 33783 4080 33817
rect 4000 33497 4080 33783
rect 4000 33463 4023 33497
rect 4057 33463 4080 33497
rect 4000 33440 4080 33463
rect 4160 33817 4240 33840
rect 4160 33783 4183 33817
rect 4217 33783 4240 33817
rect 4160 33497 4240 33783
rect 4160 33463 4183 33497
rect 4217 33463 4240 33497
rect 4160 33440 4240 33463
rect 4320 33817 4400 33840
rect 4320 33783 4343 33817
rect 4377 33783 4400 33817
rect 4320 33497 4400 33783
rect 4320 33463 4343 33497
rect 4377 33463 4400 33497
rect 4320 33440 4400 33463
rect 4480 33817 4560 33840
rect 4480 33783 4503 33817
rect 4537 33783 4560 33817
rect 4480 33497 4560 33783
rect 4480 33463 4503 33497
rect 4537 33463 4560 33497
rect 4480 33440 4560 33463
rect 4640 33817 4720 33840
rect 4640 33783 4663 33817
rect 4697 33783 4720 33817
rect 4640 33497 4720 33783
rect 4640 33463 4663 33497
rect 4697 33463 4720 33497
rect 4640 33440 4720 33463
rect 4800 33817 4880 33840
rect 4800 33783 4823 33817
rect 4857 33783 4880 33817
rect 4800 33497 4880 33783
rect 4800 33463 4823 33497
rect 4857 33463 4880 33497
rect 4800 33440 4880 33463
rect 4960 33817 5040 33840
rect 4960 33783 4983 33817
rect 5017 33783 5040 33817
rect 4960 33497 5040 33783
rect 4960 33463 4983 33497
rect 5017 33463 5040 33497
rect 4960 33440 5040 33463
rect 5120 33817 5200 33840
rect 5120 33783 5143 33817
rect 5177 33783 5200 33817
rect 5120 33497 5200 33783
rect 5120 33463 5143 33497
rect 5177 33463 5200 33497
rect 5120 33440 5200 33463
rect 5280 33817 5360 33840
rect 5280 33783 5303 33817
rect 5337 33783 5360 33817
rect 5280 33497 5360 33783
rect 5280 33463 5303 33497
rect 5337 33463 5360 33497
rect 5280 33440 5360 33463
rect 5440 33817 5520 33840
rect 5440 33783 5463 33817
rect 5497 33783 5520 33817
rect 5440 33497 5520 33783
rect 5440 33463 5463 33497
rect 5497 33463 5520 33497
rect 5440 33440 5520 33463
rect 5600 33817 5680 33840
rect 5600 33783 5623 33817
rect 5657 33783 5680 33817
rect 5600 33497 5680 33783
rect 5600 33463 5623 33497
rect 5657 33463 5680 33497
rect 5600 33440 5680 33463
rect 5760 33817 5840 33840
rect 5760 33783 5783 33817
rect 5817 33783 5840 33817
rect 5760 33497 5840 33783
rect 5760 33463 5783 33497
rect 5817 33463 5840 33497
rect 5760 33440 5840 33463
rect 5920 33817 6000 33840
rect 5920 33783 5943 33817
rect 5977 33783 6000 33817
rect 5920 33497 6000 33783
rect 5920 33463 5943 33497
rect 5977 33463 6000 33497
rect 5920 33440 6000 33463
rect 6080 33817 6160 33840
rect 6080 33783 6103 33817
rect 6137 33783 6160 33817
rect 6080 33497 6160 33783
rect 6080 33463 6103 33497
rect 6137 33463 6160 33497
rect 6080 33440 6160 33463
rect 6240 33817 6320 33840
rect 6240 33783 6263 33817
rect 6297 33783 6320 33817
rect 6240 33497 6320 33783
rect 6240 33463 6263 33497
rect 6297 33463 6320 33497
rect 6240 33440 6320 33463
rect 6400 33817 6480 33840
rect 6400 33783 6423 33817
rect 6457 33783 6480 33817
rect 6400 33497 6480 33783
rect 6400 33463 6423 33497
rect 6457 33463 6480 33497
rect 6400 33440 6480 33463
rect 6560 33817 6640 33840
rect 6560 33783 6583 33817
rect 6617 33783 6640 33817
rect 6560 33497 6640 33783
rect 6560 33463 6583 33497
rect 6617 33463 6640 33497
rect 6560 33440 6640 33463
rect 6720 33817 6800 33840
rect 6720 33783 6743 33817
rect 6777 33783 6800 33817
rect 6720 33497 6800 33783
rect 6720 33463 6743 33497
rect 6777 33463 6800 33497
rect 6720 33440 6800 33463
rect 6880 33817 6960 33840
rect 6880 33783 6903 33817
rect 6937 33783 6960 33817
rect 6880 33497 6960 33783
rect 6880 33463 6903 33497
rect 6937 33463 6960 33497
rect 6880 33440 6960 33463
rect 7040 33817 7120 33840
rect 7040 33783 7063 33817
rect 7097 33783 7120 33817
rect 7040 33497 7120 33783
rect 7040 33463 7063 33497
rect 7097 33463 7120 33497
rect 7040 33440 7120 33463
rect 7200 33817 7280 33840
rect 7200 33783 7223 33817
rect 7257 33783 7280 33817
rect 7200 33497 7280 33783
rect 7200 33463 7223 33497
rect 7257 33463 7280 33497
rect 7200 33440 7280 33463
rect 7360 33817 7440 33840
rect 7360 33783 7383 33817
rect 7417 33783 7440 33817
rect 7360 33497 7440 33783
rect 7360 33463 7383 33497
rect 7417 33463 7440 33497
rect 7360 33440 7440 33463
rect 7520 33817 7600 33840
rect 7520 33783 7543 33817
rect 7577 33783 7600 33817
rect 7520 33497 7600 33783
rect 7520 33463 7543 33497
rect 7577 33463 7600 33497
rect 7520 33440 7600 33463
rect 7680 33817 7760 33840
rect 7680 33783 7703 33817
rect 7737 33783 7760 33817
rect 7680 33497 7760 33783
rect 7680 33463 7703 33497
rect 7737 33463 7760 33497
rect 7680 33440 7760 33463
rect 7840 33817 7920 33840
rect 7840 33783 7863 33817
rect 7897 33783 7920 33817
rect 7840 33497 7920 33783
rect 7840 33463 7863 33497
rect 7897 33463 7920 33497
rect 7840 33440 7920 33463
rect 8000 33817 8080 33840
rect 8000 33783 8023 33817
rect 8057 33783 8080 33817
rect 8000 33497 8080 33783
rect 8000 33463 8023 33497
rect 8057 33463 8080 33497
rect 8000 33440 8080 33463
rect 8160 33817 8240 33840
rect 8160 33783 8183 33817
rect 8217 33783 8240 33817
rect 8160 33497 8240 33783
rect 8160 33463 8183 33497
rect 8217 33463 8240 33497
rect 8160 33440 8240 33463
rect 8320 33817 8400 33840
rect 8320 33783 8343 33817
rect 8377 33783 8400 33817
rect 8320 33497 8400 33783
rect 8320 33463 8343 33497
rect 8377 33463 8400 33497
rect 8320 33440 8400 33463
rect 8480 33440 8560 33840
rect 8640 33440 8720 33840
rect 8800 33440 8880 33840
rect 8960 33440 9040 33840
rect 9120 33440 9200 33840
rect 9280 33440 9360 33840
rect 9440 33440 9520 33840
rect 9600 33440 9680 33840
rect 9760 33440 9840 33840
rect 9920 33440 10000 33840
rect 10080 33440 10160 33840
rect 10240 33440 10320 33840
rect 10400 33440 10480 33840
rect 10560 33440 10640 33840
rect 10720 33440 10800 33840
rect 10880 33440 10960 33840
rect 11040 33440 11120 33840
rect 11200 33440 11280 33840
rect 11360 33440 11440 33840
rect 11520 33440 11600 33840
rect 11680 33440 11760 33840
rect 11840 33440 11920 33840
rect 12000 33440 12080 33840
rect 12160 33440 12240 33840
rect 12320 33440 12400 33840
rect 12480 33817 12560 33840
rect 12480 33783 12503 33817
rect 12537 33783 12560 33817
rect 12480 33497 12560 33783
rect 12480 33463 12503 33497
rect 12537 33463 12560 33497
rect 12480 33440 12560 33463
rect 12640 33817 12720 33840
rect 12640 33783 12663 33817
rect 12697 33783 12720 33817
rect 12640 33497 12720 33783
rect 12640 33463 12663 33497
rect 12697 33463 12720 33497
rect 12640 33440 12720 33463
rect 12800 33817 12880 33840
rect 12800 33783 12823 33817
rect 12857 33783 12880 33817
rect 12800 33497 12880 33783
rect 12800 33463 12823 33497
rect 12857 33463 12880 33497
rect 12800 33440 12880 33463
rect 12960 33817 13040 33840
rect 12960 33783 12983 33817
rect 13017 33783 13040 33817
rect 12960 33497 13040 33783
rect 12960 33463 12983 33497
rect 13017 33463 13040 33497
rect 12960 33440 13040 33463
rect 13120 33817 13200 33840
rect 13120 33783 13143 33817
rect 13177 33783 13200 33817
rect 13120 33497 13200 33783
rect 13120 33463 13143 33497
rect 13177 33463 13200 33497
rect 13120 33440 13200 33463
rect 13280 33817 13360 33840
rect 13280 33783 13303 33817
rect 13337 33783 13360 33817
rect 13280 33497 13360 33783
rect 13280 33463 13303 33497
rect 13337 33463 13360 33497
rect 13280 33440 13360 33463
rect 13440 33817 13520 33840
rect 13440 33783 13463 33817
rect 13497 33783 13520 33817
rect 13440 33497 13520 33783
rect 13440 33463 13463 33497
rect 13497 33463 13520 33497
rect 13440 33440 13520 33463
rect 13600 33817 13680 33840
rect 13600 33783 13623 33817
rect 13657 33783 13680 33817
rect 13600 33497 13680 33783
rect 13600 33463 13623 33497
rect 13657 33463 13680 33497
rect 13600 33440 13680 33463
rect 13760 33817 13840 33840
rect 13760 33783 13783 33817
rect 13817 33783 13840 33817
rect 13760 33497 13840 33783
rect 13760 33463 13783 33497
rect 13817 33463 13840 33497
rect 13760 33440 13840 33463
rect 13920 33817 14000 33840
rect 13920 33783 13943 33817
rect 13977 33783 14000 33817
rect 13920 33497 14000 33783
rect 13920 33463 13943 33497
rect 13977 33463 14000 33497
rect 13920 33440 14000 33463
rect 14080 33817 14160 33840
rect 14080 33783 14103 33817
rect 14137 33783 14160 33817
rect 14080 33497 14160 33783
rect 14080 33463 14103 33497
rect 14137 33463 14160 33497
rect 14080 33440 14160 33463
rect 14240 33817 14320 33840
rect 14240 33783 14263 33817
rect 14297 33783 14320 33817
rect 14240 33497 14320 33783
rect 14240 33463 14263 33497
rect 14297 33463 14320 33497
rect 14240 33440 14320 33463
rect 14400 33817 14480 33840
rect 14400 33783 14423 33817
rect 14457 33783 14480 33817
rect 14400 33497 14480 33783
rect 14400 33463 14423 33497
rect 14457 33463 14480 33497
rect 14400 33440 14480 33463
rect 14560 33817 14640 33840
rect 14560 33783 14583 33817
rect 14617 33783 14640 33817
rect 14560 33497 14640 33783
rect 14560 33463 14583 33497
rect 14617 33463 14640 33497
rect 14560 33440 14640 33463
rect 14720 33817 14800 33840
rect 14720 33783 14743 33817
rect 14777 33783 14800 33817
rect 14720 33497 14800 33783
rect 14720 33463 14743 33497
rect 14777 33463 14800 33497
rect 14720 33440 14800 33463
rect 14880 33817 14960 33840
rect 14880 33783 14903 33817
rect 14937 33783 14960 33817
rect 14880 33497 14960 33783
rect 14880 33463 14903 33497
rect 14937 33463 14960 33497
rect 14880 33440 14960 33463
rect 15040 33817 15120 33840
rect 15040 33783 15063 33817
rect 15097 33783 15120 33817
rect 15040 33497 15120 33783
rect 15040 33463 15063 33497
rect 15097 33463 15120 33497
rect 15040 33440 15120 33463
rect 15200 33817 15280 33840
rect 15200 33783 15223 33817
rect 15257 33783 15280 33817
rect 15200 33497 15280 33783
rect 15200 33463 15223 33497
rect 15257 33463 15280 33497
rect 15200 33440 15280 33463
rect 15360 33817 15440 33840
rect 15360 33783 15383 33817
rect 15417 33783 15440 33817
rect 15360 33497 15440 33783
rect 15360 33463 15383 33497
rect 15417 33463 15440 33497
rect 15360 33440 15440 33463
rect 15520 33817 15600 33840
rect 15520 33783 15543 33817
rect 15577 33783 15600 33817
rect 15520 33497 15600 33783
rect 15520 33463 15543 33497
rect 15577 33463 15600 33497
rect 15520 33440 15600 33463
rect 15680 33817 15760 33840
rect 15680 33783 15703 33817
rect 15737 33783 15760 33817
rect 15680 33497 15760 33783
rect 15680 33463 15703 33497
rect 15737 33463 15760 33497
rect 15680 33440 15760 33463
rect 15840 33817 15920 33840
rect 15840 33783 15863 33817
rect 15897 33783 15920 33817
rect 15840 33497 15920 33783
rect 15840 33463 15863 33497
rect 15897 33463 15920 33497
rect 15840 33440 15920 33463
rect 16000 33817 16080 33840
rect 16000 33783 16023 33817
rect 16057 33783 16080 33817
rect 16000 33497 16080 33783
rect 16000 33463 16023 33497
rect 16057 33463 16080 33497
rect 16000 33440 16080 33463
rect 16160 33817 16240 33840
rect 16160 33783 16183 33817
rect 16217 33783 16240 33817
rect 16160 33497 16240 33783
rect 16160 33463 16183 33497
rect 16217 33463 16240 33497
rect 16160 33440 16240 33463
rect 16320 33817 16400 33840
rect 16320 33783 16343 33817
rect 16377 33783 16400 33817
rect 16320 33497 16400 33783
rect 16320 33463 16343 33497
rect 16377 33463 16400 33497
rect 16320 33440 16400 33463
rect 16480 33817 16560 33840
rect 16480 33783 16503 33817
rect 16537 33783 16560 33817
rect 16480 33497 16560 33783
rect 16480 33463 16503 33497
rect 16537 33463 16560 33497
rect 16480 33440 16560 33463
rect 16640 33817 16720 33840
rect 16640 33783 16663 33817
rect 16697 33783 16720 33817
rect 16640 33497 16720 33783
rect 16640 33463 16663 33497
rect 16697 33463 16720 33497
rect 16640 33440 16720 33463
rect 16800 33817 16880 33840
rect 16800 33783 16823 33817
rect 16857 33783 16880 33817
rect 16800 33497 16880 33783
rect 16800 33463 16823 33497
rect 16857 33463 16880 33497
rect 16800 33440 16880 33463
rect 16960 33817 17040 33840
rect 16960 33783 16983 33817
rect 17017 33783 17040 33817
rect 16960 33497 17040 33783
rect 16960 33463 16983 33497
rect 17017 33463 17040 33497
rect 16960 33440 17040 33463
rect 17120 33817 17200 33840
rect 17120 33783 17143 33817
rect 17177 33783 17200 33817
rect 17120 33497 17200 33783
rect 17120 33463 17143 33497
rect 17177 33463 17200 33497
rect 17120 33440 17200 33463
rect 17280 33817 17360 33840
rect 17280 33783 17303 33817
rect 17337 33783 17360 33817
rect 17280 33497 17360 33783
rect 17280 33463 17303 33497
rect 17337 33463 17360 33497
rect 17280 33440 17360 33463
rect 17440 33817 17520 33840
rect 17440 33783 17463 33817
rect 17497 33783 17520 33817
rect 17440 33497 17520 33783
rect 17440 33463 17463 33497
rect 17497 33463 17520 33497
rect 17440 33440 17520 33463
rect 17600 33817 17680 33840
rect 17600 33783 17623 33817
rect 17657 33783 17680 33817
rect 17600 33497 17680 33783
rect 17600 33463 17623 33497
rect 17657 33463 17680 33497
rect 17600 33440 17680 33463
rect 17760 33817 17840 33840
rect 17760 33783 17783 33817
rect 17817 33783 17840 33817
rect 17760 33497 17840 33783
rect 17760 33463 17783 33497
rect 17817 33463 17840 33497
rect 17760 33440 17840 33463
rect 17920 33817 18000 33840
rect 17920 33783 17943 33817
rect 17977 33783 18000 33817
rect 17920 33497 18000 33783
rect 17920 33463 17943 33497
rect 17977 33463 18000 33497
rect 17920 33440 18000 33463
rect 18080 33817 18160 33840
rect 18080 33783 18103 33817
rect 18137 33783 18160 33817
rect 18080 33497 18160 33783
rect 18080 33463 18103 33497
rect 18137 33463 18160 33497
rect 18080 33440 18160 33463
rect 18240 33817 18320 33840
rect 18240 33783 18263 33817
rect 18297 33783 18320 33817
rect 18240 33497 18320 33783
rect 18240 33463 18263 33497
rect 18297 33463 18320 33497
rect 18240 33440 18320 33463
rect 18400 33817 18480 33840
rect 18400 33783 18423 33817
rect 18457 33783 18480 33817
rect 18400 33497 18480 33783
rect 18400 33463 18423 33497
rect 18457 33463 18480 33497
rect 18400 33440 18480 33463
rect 18560 33817 18640 33840
rect 18560 33783 18583 33817
rect 18617 33783 18640 33817
rect 18560 33497 18640 33783
rect 18560 33463 18583 33497
rect 18617 33463 18640 33497
rect 18560 33440 18640 33463
rect 18720 33817 18800 33840
rect 18720 33783 18743 33817
rect 18777 33783 18800 33817
rect 18720 33497 18800 33783
rect 18720 33463 18743 33497
rect 18777 33463 18800 33497
rect 18720 33440 18800 33463
rect 18880 33817 18960 33840
rect 18880 33783 18903 33817
rect 18937 33783 18960 33817
rect 18880 33497 18960 33783
rect 18880 33463 18903 33497
rect 18937 33463 18960 33497
rect 18880 33440 18960 33463
rect 19040 33440 19120 33840
rect 19200 33440 19280 33840
rect 19360 33440 19440 33840
rect 19520 33440 19600 33840
rect 19680 33440 19760 33840
rect 19840 33440 19920 33840
rect 20000 33440 20080 33840
rect 20160 33440 20240 33840
rect 20320 33440 20400 33840
rect 20480 33440 20560 33840
rect 20640 33440 20720 33840
rect 20800 33440 20880 33840
rect 20960 33440 21040 33840
rect 21120 33440 21200 33840
rect 21280 33440 21360 33840
rect 21440 33440 21520 33840
rect 21600 33440 21680 33840
rect 21760 33440 21840 33840
rect 21920 33440 22000 33840
rect 22080 33440 22160 33840
rect 22240 33440 22320 33840
rect 22400 33440 22480 33840
rect 22560 33440 22640 33840
rect 22720 33440 22800 33840
rect 22880 33440 22960 33840
rect 23120 33817 23200 33840
rect 23120 33783 23143 33817
rect 23177 33783 23200 33817
rect 23120 33497 23200 33783
rect 23120 33463 23143 33497
rect 23177 33463 23200 33497
rect 23120 33440 23200 33463
rect 23280 33817 23360 33840
rect 23280 33783 23303 33817
rect 23337 33783 23360 33817
rect 23280 33497 23360 33783
rect 23280 33463 23303 33497
rect 23337 33463 23360 33497
rect 23280 33440 23360 33463
rect 23440 33817 23520 33840
rect 23440 33783 23463 33817
rect 23497 33783 23520 33817
rect 23440 33497 23520 33783
rect 23440 33463 23463 33497
rect 23497 33463 23520 33497
rect 23440 33440 23520 33463
rect 23600 33817 23680 33840
rect 23600 33783 23623 33817
rect 23657 33783 23680 33817
rect 23600 33497 23680 33783
rect 23600 33463 23623 33497
rect 23657 33463 23680 33497
rect 23600 33440 23680 33463
rect 23760 33817 23840 33840
rect 23760 33783 23783 33817
rect 23817 33783 23840 33817
rect 23760 33497 23840 33783
rect 23760 33463 23783 33497
rect 23817 33463 23840 33497
rect 23760 33440 23840 33463
rect 23920 33817 24000 33840
rect 23920 33783 23943 33817
rect 23977 33783 24000 33817
rect 23920 33497 24000 33783
rect 23920 33463 23943 33497
rect 23977 33463 24000 33497
rect 23920 33440 24000 33463
rect 24080 33817 24160 33840
rect 24080 33783 24103 33817
rect 24137 33783 24160 33817
rect 24080 33497 24160 33783
rect 24080 33463 24103 33497
rect 24137 33463 24160 33497
rect 24080 33440 24160 33463
rect 24240 33817 24320 33840
rect 24240 33783 24263 33817
rect 24297 33783 24320 33817
rect 24240 33497 24320 33783
rect 24240 33463 24263 33497
rect 24297 33463 24320 33497
rect 24240 33440 24320 33463
rect 24400 33817 24480 33840
rect 24400 33783 24423 33817
rect 24457 33783 24480 33817
rect 24400 33497 24480 33783
rect 24400 33463 24423 33497
rect 24457 33463 24480 33497
rect 24400 33440 24480 33463
rect 24560 33817 24640 33840
rect 24560 33783 24583 33817
rect 24617 33783 24640 33817
rect 24560 33497 24640 33783
rect 24560 33463 24583 33497
rect 24617 33463 24640 33497
rect 24560 33440 24640 33463
rect 24720 33817 24800 33840
rect 24720 33783 24743 33817
rect 24777 33783 24800 33817
rect 24720 33497 24800 33783
rect 24720 33463 24743 33497
rect 24777 33463 24800 33497
rect 24720 33440 24800 33463
rect 24880 33817 24960 33840
rect 24880 33783 24903 33817
rect 24937 33783 24960 33817
rect 24880 33497 24960 33783
rect 24880 33463 24903 33497
rect 24937 33463 24960 33497
rect 24880 33440 24960 33463
rect 25040 33817 25120 33840
rect 25040 33783 25063 33817
rect 25097 33783 25120 33817
rect 25040 33497 25120 33783
rect 25040 33463 25063 33497
rect 25097 33463 25120 33497
rect 25040 33440 25120 33463
rect 25200 33817 25280 33840
rect 25200 33783 25223 33817
rect 25257 33783 25280 33817
rect 25200 33497 25280 33783
rect 25200 33463 25223 33497
rect 25257 33463 25280 33497
rect 25200 33440 25280 33463
rect 25360 33817 25440 33840
rect 25360 33783 25383 33817
rect 25417 33783 25440 33817
rect 25360 33497 25440 33783
rect 25360 33463 25383 33497
rect 25417 33463 25440 33497
rect 25360 33440 25440 33463
rect 25520 33817 25600 33840
rect 25520 33783 25543 33817
rect 25577 33783 25600 33817
rect 25520 33497 25600 33783
rect 25520 33463 25543 33497
rect 25577 33463 25600 33497
rect 25520 33440 25600 33463
rect 25680 33817 25760 33840
rect 25680 33783 25703 33817
rect 25737 33783 25760 33817
rect 25680 33497 25760 33783
rect 25680 33463 25703 33497
rect 25737 33463 25760 33497
rect 25680 33440 25760 33463
rect 25840 33817 25920 33840
rect 25840 33783 25863 33817
rect 25897 33783 25920 33817
rect 25840 33497 25920 33783
rect 25840 33463 25863 33497
rect 25897 33463 25920 33497
rect 25840 33440 25920 33463
rect 26000 33817 26080 33840
rect 26000 33783 26023 33817
rect 26057 33783 26080 33817
rect 26000 33497 26080 33783
rect 26000 33463 26023 33497
rect 26057 33463 26080 33497
rect 26000 33440 26080 33463
rect 26160 33817 26240 33840
rect 26160 33783 26183 33817
rect 26217 33783 26240 33817
rect 26160 33497 26240 33783
rect 26160 33463 26183 33497
rect 26217 33463 26240 33497
rect 26160 33440 26240 33463
rect 26320 33817 26400 33840
rect 26320 33783 26343 33817
rect 26377 33783 26400 33817
rect 26320 33497 26400 33783
rect 26320 33463 26343 33497
rect 26377 33463 26400 33497
rect 26320 33440 26400 33463
rect 26480 33817 26560 33840
rect 26480 33783 26503 33817
rect 26537 33783 26560 33817
rect 26480 33497 26560 33783
rect 26480 33463 26503 33497
rect 26537 33463 26560 33497
rect 26480 33440 26560 33463
rect 26640 33817 26720 33840
rect 26640 33783 26663 33817
rect 26697 33783 26720 33817
rect 26640 33497 26720 33783
rect 26640 33463 26663 33497
rect 26697 33463 26720 33497
rect 26640 33440 26720 33463
rect 26800 33817 26880 33840
rect 26800 33783 26823 33817
rect 26857 33783 26880 33817
rect 26800 33497 26880 33783
rect 26800 33463 26823 33497
rect 26857 33463 26880 33497
rect 26800 33440 26880 33463
rect 26960 33817 27040 33840
rect 26960 33783 26983 33817
rect 27017 33783 27040 33817
rect 26960 33497 27040 33783
rect 26960 33463 26983 33497
rect 27017 33463 27040 33497
rect 26960 33440 27040 33463
rect 27120 33817 27200 33840
rect 27120 33783 27143 33817
rect 27177 33783 27200 33817
rect 27120 33497 27200 33783
rect 27120 33463 27143 33497
rect 27177 33463 27200 33497
rect 27120 33440 27200 33463
rect 27280 33817 27360 33840
rect 27280 33783 27303 33817
rect 27337 33783 27360 33817
rect 27280 33497 27360 33783
rect 27280 33463 27303 33497
rect 27337 33463 27360 33497
rect 27280 33440 27360 33463
rect 27440 33817 27520 33840
rect 27440 33783 27463 33817
rect 27497 33783 27520 33817
rect 27440 33497 27520 33783
rect 27440 33463 27463 33497
rect 27497 33463 27520 33497
rect 27440 33440 27520 33463
rect 27600 33817 27680 33840
rect 27600 33783 27623 33817
rect 27657 33783 27680 33817
rect 27600 33497 27680 33783
rect 27600 33463 27623 33497
rect 27657 33463 27680 33497
rect 27600 33440 27680 33463
rect 27760 33817 27840 33840
rect 27760 33783 27783 33817
rect 27817 33783 27840 33817
rect 27760 33497 27840 33783
rect 27760 33463 27783 33497
rect 27817 33463 27840 33497
rect 27760 33440 27840 33463
rect 27920 33817 28000 33840
rect 27920 33783 27943 33817
rect 27977 33783 28000 33817
rect 27920 33497 28000 33783
rect 27920 33463 27943 33497
rect 27977 33463 28000 33497
rect 27920 33440 28000 33463
rect 28080 33817 28160 33840
rect 28080 33783 28103 33817
rect 28137 33783 28160 33817
rect 28080 33497 28160 33783
rect 28080 33463 28103 33497
rect 28137 33463 28160 33497
rect 28080 33440 28160 33463
rect 28240 33817 28320 33840
rect 28240 33783 28263 33817
rect 28297 33783 28320 33817
rect 28240 33497 28320 33783
rect 28240 33463 28263 33497
rect 28297 33463 28320 33497
rect 28240 33440 28320 33463
rect 28400 33817 28480 33840
rect 28400 33783 28423 33817
rect 28457 33783 28480 33817
rect 28400 33497 28480 33783
rect 28400 33463 28423 33497
rect 28457 33463 28480 33497
rect 28400 33440 28480 33463
rect 28560 33817 28640 33840
rect 28560 33783 28583 33817
rect 28617 33783 28640 33817
rect 28560 33497 28640 33783
rect 28560 33463 28583 33497
rect 28617 33463 28640 33497
rect 28560 33440 28640 33463
rect 28720 33817 28800 33840
rect 28720 33783 28743 33817
rect 28777 33783 28800 33817
rect 28720 33497 28800 33783
rect 28720 33463 28743 33497
rect 28777 33463 28800 33497
rect 28720 33440 28800 33463
rect 28880 33817 28960 33840
rect 28880 33783 28903 33817
rect 28937 33783 28960 33817
rect 28880 33497 28960 33783
rect 28880 33463 28903 33497
rect 28937 33463 28960 33497
rect 28880 33440 28960 33463
rect 29040 33817 29120 33840
rect 29040 33783 29063 33817
rect 29097 33783 29120 33817
rect 29040 33497 29120 33783
rect 29040 33463 29063 33497
rect 29097 33463 29120 33497
rect 29040 33440 29120 33463
rect 29200 33817 29280 33840
rect 29200 33783 29223 33817
rect 29257 33783 29280 33817
rect 29200 33497 29280 33783
rect 29200 33463 29223 33497
rect 29257 33463 29280 33497
rect 29200 33440 29280 33463
rect 29360 33817 29440 33840
rect 29360 33783 29383 33817
rect 29417 33783 29440 33817
rect 29360 33497 29440 33783
rect 29360 33463 29383 33497
rect 29417 33463 29440 33497
rect 29360 33440 29440 33463
rect 29520 33440 29600 33840
rect 29680 33440 29760 33840
rect 29840 33440 29920 33840
rect 30000 33440 30080 33840
rect 30160 33440 30240 33840
rect 30320 33440 30400 33840
rect 30480 33440 30560 33840
rect 30640 33440 30720 33840
rect 30800 33440 30880 33840
rect 30960 33440 31040 33840
rect 31120 33440 31200 33840
rect 31280 33440 31360 33840
rect 31440 33440 31520 33840
rect 31600 33440 31680 33840
rect 31760 33440 31840 33840
rect 31920 33440 32000 33840
rect 32080 33440 32160 33840
rect 32240 33440 32320 33840
rect 32400 33440 32480 33840
rect 32560 33440 32640 33840
rect 32720 33440 32800 33840
rect 32880 33440 32960 33840
rect 33040 33440 33120 33840
rect 33200 33440 33280 33840
rect 33360 33440 33440 33840
rect 33520 33817 33600 33840
rect 33520 33783 33543 33817
rect 33577 33783 33600 33817
rect 33520 33497 33600 33783
rect 33520 33463 33543 33497
rect 33577 33463 33600 33497
rect 33520 33440 33600 33463
rect 33680 33817 33760 33840
rect 33680 33783 33703 33817
rect 33737 33783 33760 33817
rect 33680 33497 33760 33783
rect 33680 33463 33703 33497
rect 33737 33463 33760 33497
rect 33680 33440 33760 33463
rect 33840 33817 33920 33840
rect 33840 33783 33863 33817
rect 33897 33783 33920 33817
rect 33840 33497 33920 33783
rect 33840 33463 33863 33497
rect 33897 33463 33920 33497
rect 33840 33440 33920 33463
rect 34000 33817 34080 33840
rect 34000 33783 34023 33817
rect 34057 33783 34080 33817
rect 34000 33497 34080 33783
rect 34000 33463 34023 33497
rect 34057 33463 34080 33497
rect 34000 33440 34080 33463
rect 34160 33817 34240 33840
rect 34160 33783 34183 33817
rect 34217 33783 34240 33817
rect 34160 33497 34240 33783
rect 34160 33463 34183 33497
rect 34217 33463 34240 33497
rect 34160 33440 34240 33463
rect 34320 33817 34400 33840
rect 34320 33783 34343 33817
rect 34377 33783 34400 33817
rect 34320 33497 34400 33783
rect 34320 33463 34343 33497
rect 34377 33463 34400 33497
rect 34320 33440 34400 33463
rect 34480 33817 34560 33840
rect 34480 33783 34503 33817
rect 34537 33783 34560 33817
rect 34480 33497 34560 33783
rect 34480 33463 34503 33497
rect 34537 33463 34560 33497
rect 34480 33440 34560 33463
rect 34640 33817 34720 33840
rect 34640 33783 34663 33817
rect 34697 33783 34720 33817
rect 34640 33497 34720 33783
rect 34640 33463 34663 33497
rect 34697 33463 34720 33497
rect 34640 33440 34720 33463
rect 34800 33817 34880 33840
rect 34800 33783 34823 33817
rect 34857 33783 34880 33817
rect 34800 33497 34880 33783
rect 34800 33463 34823 33497
rect 34857 33463 34880 33497
rect 34800 33440 34880 33463
rect 34960 33817 35040 33840
rect 34960 33783 34983 33817
rect 35017 33783 35040 33817
rect 34960 33497 35040 33783
rect 34960 33463 34983 33497
rect 35017 33463 35040 33497
rect 34960 33440 35040 33463
rect 35120 33817 35200 33840
rect 35120 33783 35143 33817
rect 35177 33783 35200 33817
rect 35120 33497 35200 33783
rect 35120 33463 35143 33497
rect 35177 33463 35200 33497
rect 35120 33440 35200 33463
rect 35280 33817 35360 33840
rect 35280 33783 35303 33817
rect 35337 33783 35360 33817
rect 35280 33497 35360 33783
rect 35280 33463 35303 33497
rect 35337 33463 35360 33497
rect 35280 33440 35360 33463
rect 35440 33817 35520 33840
rect 35440 33783 35463 33817
rect 35497 33783 35520 33817
rect 35440 33497 35520 33783
rect 35440 33463 35463 33497
rect 35497 33463 35520 33497
rect 35440 33440 35520 33463
rect 35600 33817 35680 33840
rect 35600 33783 35623 33817
rect 35657 33783 35680 33817
rect 35600 33497 35680 33783
rect 35600 33463 35623 33497
rect 35657 33463 35680 33497
rect 35600 33440 35680 33463
rect 35760 33817 35840 33840
rect 35760 33783 35783 33817
rect 35817 33783 35840 33817
rect 35760 33497 35840 33783
rect 35760 33463 35783 33497
rect 35817 33463 35840 33497
rect 35760 33440 35840 33463
rect 35920 33817 36000 33840
rect 35920 33783 35943 33817
rect 35977 33783 36000 33817
rect 35920 33497 36000 33783
rect 35920 33463 35943 33497
rect 35977 33463 36000 33497
rect 35920 33440 36000 33463
rect 36080 33817 36160 33840
rect 36080 33783 36103 33817
rect 36137 33783 36160 33817
rect 36080 33497 36160 33783
rect 36080 33463 36103 33497
rect 36137 33463 36160 33497
rect 36080 33440 36160 33463
rect 36240 33817 36320 33840
rect 36240 33783 36263 33817
rect 36297 33783 36320 33817
rect 36240 33497 36320 33783
rect 36240 33463 36263 33497
rect 36297 33463 36320 33497
rect 36240 33440 36320 33463
rect 36400 33817 36480 33840
rect 36400 33783 36423 33817
rect 36457 33783 36480 33817
rect 36400 33497 36480 33783
rect 36400 33463 36423 33497
rect 36457 33463 36480 33497
rect 36400 33440 36480 33463
rect 36560 33817 36640 33840
rect 36560 33783 36583 33817
rect 36617 33783 36640 33817
rect 36560 33497 36640 33783
rect 36560 33463 36583 33497
rect 36617 33463 36640 33497
rect 36560 33440 36640 33463
rect 36720 33817 36800 33840
rect 36720 33783 36743 33817
rect 36777 33783 36800 33817
rect 36720 33497 36800 33783
rect 36720 33463 36743 33497
rect 36777 33463 36800 33497
rect 36720 33440 36800 33463
rect 36880 33817 36960 33840
rect 36880 33783 36903 33817
rect 36937 33783 36960 33817
rect 36880 33497 36960 33783
rect 36880 33463 36903 33497
rect 36937 33463 36960 33497
rect 36880 33440 36960 33463
rect 37040 33817 37120 33840
rect 37040 33783 37063 33817
rect 37097 33783 37120 33817
rect 37040 33497 37120 33783
rect 37040 33463 37063 33497
rect 37097 33463 37120 33497
rect 37040 33440 37120 33463
rect 37200 33817 37280 33840
rect 37200 33783 37223 33817
rect 37257 33783 37280 33817
rect 37200 33497 37280 33783
rect 37200 33463 37223 33497
rect 37257 33463 37280 33497
rect 37200 33440 37280 33463
rect 37360 33817 37440 33840
rect 37360 33783 37383 33817
rect 37417 33783 37440 33817
rect 37360 33497 37440 33783
rect 37360 33463 37383 33497
rect 37417 33463 37440 33497
rect 37360 33440 37440 33463
rect 37520 33817 37600 33840
rect 37520 33783 37543 33817
rect 37577 33783 37600 33817
rect 37520 33497 37600 33783
rect 37520 33463 37543 33497
rect 37577 33463 37600 33497
rect 37520 33440 37600 33463
rect 37680 33817 37760 33840
rect 37680 33783 37703 33817
rect 37737 33783 37760 33817
rect 37680 33497 37760 33783
rect 37680 33463 37703 33497
rect 37737 33463 37760 33497
rect 37680 33440 37760 33463
rect 37840 33817 37920 33840
rect 37840 33783 37863 33817
rect 37897 33783 37920 33817
rect 37840 33497 37920 33783
rect 37840 33463 37863 33497
rect 37897 33463 37920 33497
rect 37840 33440 37920 33463
rect 38000 33817 38080 33840
rect 38000 33783 38023 33817
rect 38057 33783 38080 33817
rect 38000 33497 38080 33783
rect 38000 33463 38023 33497
rect 38057 33463 38080 33497
rect 38000 33440 38080 33463
rect 38160 33817 38240 33840
rect 38160 33783 38183 33817
rect 38217 33783 38240 33817
rect 38160 33497 38240 33783
rect 38160 33463 38183 33497
rect 38217 33463 38240 33497
rect 38160 33440 38240 33463
rect 38320 33817 38400 33840
rect 38320 33783 38343 33817
rect 38377 33783 38400 33817
rect 38320 33497 38400 33783
rect 38320 33463 38343 33497
rect 38377 33463 38400 33497
rect 38320 33440 38400 33463
rect 38480 33817 38560 33840
rect 38480 33783 38503 33817
rect 38537 33783 38560 33817
rect 38480 33497 38560 33783
rect 38480 33463 38503 33497
rect 38537 33463 38560 33497
rect 38480 33440 38560 33463
rect 38640 33817 38720 33840
rect 38640 33783 38663 33817
rect 38697 33783 38720 33817
rect 38640 33497 38720 33783
rect 38640 33463 38663 33497
rect 38697 33463 38720 33497
rect 38640 33440 38720 33463
rect 38800 33817 38880 33840
rect 38800 33783 38823 33817
rect 38857 33783 38880 33817
rect 38800 33497 38880 33783
rect 38800 33463 38823 33497
rect 38857 33463 38880 33497
rect 38800 33440 38880 33463
rect 38960 33817 39040 33840
rect 38960 33783 38983 33817
rect 39017 33783 39040 33817
rect 38960 33497 39040 33783
rect 38960 33463 38983 33497
rect 39017 33463 39040 33497
rect 38960 33440 39040 33463
rect 39120 33817 39200 33840
rect 39120 33783 39143 33817
rect 39177 33783 39200 33817
rect 39120 33497 39200 33783
rect 39120 33463 39143 33497
rect 39177 33463 39200 33497
rect 39120 33440 39200 33463
rect 39280 33817 39360 33840
rect 39280 33783 39303 33817
rect 39337 33783 39360 33817
rect 39280 33497 39360 33783
rect 39280 33463 39303 33497
rect 39337 33463 39360 33497
rect 39280 33440 39360 33463
rect 39440 33817 39520 33840
rect 39440 33783 39463 33817
rect 39497 33783 39520 33817
rect 39440 33497 39520 33783
rect 39440 33463 39463 33497
rect 39497 33463 39520 33497
rect 39440 33440 39520 33463
rect 39600 33817 39680 33840
rect 39600 33783 39623 33817
rect 39657 33783 39680 33817
rect 39600 33497 39680 33783
rect 39600 33463 39623 33497
rect 39657 33463 39680 33497
rect 39600 33440 39680 33463
rect 39760 33817 39840 33840
rect 39760 33783 39783 33817
rect 39817 33783 39840 33817
rect 39760 33497 39840 33783
rect 39760 33463 39783 33497
rect 39817 33463 39840 33497
rect 39760 33440 39840 33463
rect 39920 33817 40000 33840
rect 39920 33783 39943 33817
rect 39977 33783 40000 33817
rect 39920 33497 40000 33783
rect 39920 33463 39943 33497
rect 39977 33463 40000 33497
rect 39920 33440 40000 33463
rect 40080 33817 40160 33840
rect 40080 33783 40103 33817
rect 40137 33783 40160 33817
rect 40080 33497 40160 33783
rect 40080 33463 40103 33497
rect 40137 33463 40160 33497
rect 40080 33440 40160 33463
rect 40240 33817 40320 33840
rect 40240 33783 40263 33817
rect 40297 33783 40320 33817
rect 40240 33497 40320 33783
rect 40240 33463 40263 33497
rect 40297 33463 40320 33497
rect 40240 33440 40320 33463
rect 40400 33817 40480 33840
rect 40400 33783 40423 33817
rect 40457 33783 40480 33817
rect 40400 33497 40480 33783
rect 40400 33463 40423 33497
rect 40457 33463 40480 33497
rect 40400 33440 40480 33463
rect 40560 33817 40640 33840
rect 40560 33783 40583 33817
rect 40617 33783 40640 33817
rect 40560 33497 40640 33783
rect 40560 33463 40583 33497
rect 40617 33463 40640 33497
rect 40560 33440 40640 33463
rect 40720 33817 40800 33840
rect 40720 33783 40743 33817
rect 40777 33783 40800 33817
rect 40720 33497 40800 33783
rect 40720 33463 40743 33497
rect 40777 33463 40800 33497
rect 40720 33440 40800 33463
rect 40880 33817 40960 33840
rect 40880 33783 40903 33817
rect 40937 33783 40960 33817
rect 40880 33497 40960 33783
rect 40880 33463 40903 33497
rect 40937 33463 40960 33497
rect 40880 33440 40960 33463
rect 41040 33817 41120 33840
rect 41040 33783 41063 33817
rect 41097 33783 41120 33817
rect 41040 33497 41120 33783
rect 41040 33463 41063 33497
rect 41097 33463 41120 33497
rect 41040 33440 41120 33463
rect 41200 33817 41280 33840
rect 41200 33783 41223 33817
rect 41257 33783 41280 33817
rect 41200 33497 41280 33783
rect 41200 33463 41223 33497
rect 41257 33463 41280 33497
rect 41200 33440 41280 33463
rect 41360 33817 41440 33840
rect 41360 33783 41383 33817
rect 41417 33783 41440 33817
rect 41360 33497 41440 33783
rect 41360 33463 41383 33497
rect 41417 33463 41440 33497
rect 41360 33440 41440 33463
rect 41520 33817 41600 33840
rect 41520 33783 41543 33817
rect 41577 33783 41600 33817
rect 41520 33497 41600 33783
rect 41520 33463 41543 33497
rect 41577 33463 41600 33497
rect 41520 33440 41600 33463
rect 41680 33817 41760 33840
rect 41680 33783 41703 33817
rect 41737 33783 41760 33817
rect 41680 33497 41760 33783
rect 41680 33463 41703 33497
rect 41737 33463 41760 33497
rect 41680 33440 41760 33463
rect 41840 33817 41920 33840
rect 41840 33783 41863 33817
rect 41897 33783 41920 33817
rect 41840 33497 41920 33783
rect 41840 33463 41863 33497
rect 41897 33463 41920 33497
rect 41840 33440 41920 33463
rect 0 33337 80 33360
rect 0 33303 23 33337
rect 57 33303 80 33337
rect 0 33017 80 33303
rect 0 32983 23 33017
rect 57 32983 80 33017
rect 0 32960 80 32983
rect 160 33337 240 33360
rect 160 33303 183 33337
rect 217 33303 240 33337
rect 160 33017 240 33303
rect 160 32983 183 33017
rect 217 32983 240 33017
rect 160 32960 240 32983
rect 320 33337 400 33360
rect 320 33303 343 33337
rect 377 33303 400 33337
rect 320 33017 400 33303
rect 320 32983 343 33017
rect 377 32983 400 33017
rect 320 32960 400 32983
rect 480 33337 560 33360
rect 480 33303 503 33337
rect 537 33303 560 33337
rect 480 33017 560 33303
rect 480 32983 503 33017
rect 537 32983 560 33017
rect 480 32960 560 32983
rect 640 33337 720 33360
rect 640 33303 663 33337
rect 697 33303 720 33337
rect 640 33017 720 33303
rect 640 32983 663 33017
rect 697 32983 720 33017
rect 640 32960 720 32983
rect 800 33337 880 33360
rect 800 33303 823 33337
rect 857 33303 880 33337
rect 800 33017 880 33303
rect 800 32983 823 33017
rect 857 32983 880 33017
rect 800 32960 880 32983
rect 960 33337 1040 33360
rect 960 33303 983 33337
rect 1017 33303 1040 33337
rect 960 33017 1040 33303
rect 960 32983 983 33017
rect 1017 32983 1040 33017
rect 960 32960 1040 32983
rect 1120 33337 1200 33360
rect 1120 33303 1143 33337
rect 1177 33303 1200 33337
rect 1120 33017 1200 33303
rect 1120 32983 1143 33017
rect 1177 32983 1200 33017
rect 1120 32960 1200 32983
rect 1280 33337 1360 33360
rect 1280 33303 1303 33337
rect 1337 33303 1360 33337
rect 1280 33017 1360 33303
rect 1280 32983 1303 33017
rect 1337 32983 1360 33017
rect 1280 32960 1360 32983
rect 1440 33337 1520 33360
rect 1440 33303 1463 33337
rect 1497 33303 1520 33337
rect 1440 33017 1520 33303
rect 1440 32983 1463 33017
rect 1497 32983 1520 33017
rect 1440 32960 1520 32983
rect 1600 33337 1680 33360
rect 1600 33303 1623 33337
rect 1657 33303 1680 33337
rect 1600 33017 1680 33303
rect 1600 32983 1623 33017
rect 1657 32983 1680 33017
rect 1600 32960 1680 32983
rect 1760 33337 1840 33360
rect 1760 33303 1783 33337
rect 1817 33303 1840 33337
rect 1760 33017 1840 33303
rect 1760 32983 1783 33017
rect 1817 32983 1840 33017
rect 1760 32960 1840 32983
rect 1920 33337 2000 33360
rect 1920 33303 1943 33337
rect 1977 33303 2000 33337
rect 1920 33017 2000 33303
rect 1920 32983 1943 33017
rect 1977 32983 2000 33017
rect 1920 32960 2000 32983
rect 2080 33337 2160 33360
rect 2080 33303 2103 33337
rect 2137 33303 2160 33337
rect 2080 33017 2160 33303
rect 2080 32983 2103 33017
rect 2137 32983 2160 33017
rect 2080 32960 2160 32983
rect 2240 33337 2320 33360
rect 2240 33303 2263 33337
rect 2297 33303 2320 33337
rect 2240 33017 2320 33303
rect 2240 32983 2263 33017
rect 2297 32983 2320 33017
rect 2240 32960 2320 32983
rect 2400 33337 2480 33360
rect 2400 33303 2423 33337
rect 2457 33303 2480 33337
rect 2400 33017 2480 33303
rect 2400 32983 2423 33017
rect 2457 32983 2480 33017
rect 2400 32960 2480 32983
rect 2560 33337 2640 33360
rect 2560 33303 2583 33337
rect 2617 33303 2640 33337
rect 2560 33017 2640 33303
rect 2560 32983 2583 33017
rect 2617 32983 2640 33017
rect 2560 32960 2640 32983
rect 2720 33337 2800 33360
rect 2720 33303 2743 33337
rect 2777 33303 2800 33337
rect 2720 33017 2800 33303
rect 2720 32983 2743 33017
rect 2777 32983 2800 33017
rect 2720 32960 2800 32983
rect 2880 33337 2960 33360
rect 2880 33303 2903 33337
rect 2937 33303 2960 33337
rect 2880 33017 2960 33303
rect 2880 32983 2903 33017
rect 2937 32983 2960 33017
rect 2880 32960 2960 32983
rect 3040 33337 3120 33360
rect 3040 33303 3063 33337
rect 3097 33303 3120 33337
rect 3040 33017 3120 33303
rect 3040 32983 3063 33017
rect 3097 32983 3120 33017
rect 3040 32960 3120 32983
rect 3200 33337 3280 33360
rect 3200 33303 3223 33337
rect 3257 33303 3280 33337
rect 3200 33017 3280 33303
rect 3200 32983 3223 33017
rect 3257 32983 3280 33017
rect 3200 32960 3280 32983
rect 3360 33337 3440 33360
rect 3360 33303 3383 33337
rect 3417 33303 3440 33337
rect 3360 33017 3440 33303
rect 3360 32983 3383 33017
rect 3417 32983 3440 33017
rect 3360 32960 3440 32983
rect 3520 33337 3600 33360
rect 3520 33303 3543 33337
rect 3577 33303 3600 33337
rect 3520 33017 3600 33303
rect 3520 32983 3543 33017
rect 3577 32983 3600 33017
rect 3520 32960 3600 32983
rect 3680 33337 3760 33360
rect 3680 33303 3703 33337
rect 3737 33303 3760 33337
rect 3680 33017 3760 33303
rect 3680 32983 3703 33017
rect 3737 32983 3760 33017
rect 3680 32960 3760 32983
rect 3840 33337 3920 33360
rect 3840 33303 3863 33337
rect 3897 33303 3920 33337
rect 3840 33017 3920 33303
rect 3840 32983 3863 33017
rect 3897 32983 3920 33017
rect 3840 32960 3920 32983
rect 4000 33337 4080 33360
rect 4000 33303 4023 33337
rect 4057 33303 4080 33337
rect 4000 33017 4080 33303
rect 4000 32983 4023 33017
rect 4057 32983 4080 33017
rect 4000 32960 4080 32983
rect 4160 33337 4240 33360
rect 4160 33303 4183 33337
rect 4217 33303 4240 33337
rect 4160 33017 4240 33303
rect 4160 32983 4183 33017
rect 4217 32983 4240 33017
rect 4160 32960 4240 32983
rect 4320 33337 4400 33360
rect 4320 33303 4343 33337
rect 4377 33303 4400 33337
rect 4320 33017 4400 33303
rect 4320 32983 4343 33017
rect 4377 32983 4400 33017
rect 4320 32960 4400 32983
rect 4480 33337 4560 33360
rect 4480 33303 4503 33337
rect 4537 33303 4560 33337
rect 4480 33017 4560 33303
rect 4480 32983 4503 33017
rect 4537 32983 4560 33017
rect 4480 32960 4560 32983
rect 4640 33337 4720 33360
rect 4640 33303 4663 33337
rect 4697 33303 4720 33337
rect 4640 33017 4720 33303
rect 4640 32983 4663 33017
rect 4697 32983 4720 33017
rect 4640 32960 4720 32983
rect 4800 33337 4880 33360
rect 4800 33303 4823 33337
rect 4857 33303 4880 33337
rect 4800 33017 4880 33303
rect 4800 32983 4823 33017
rect 4857 32983 4880 33017
rect 4800 32960 4880 32983
rect 4960 33337 5040 33360
rect 4960 33303 4983 33337
rect 5017 33303 5040 33337
rect 4960 33017 5040 33303
rect 4960 32983 4983 33017
rect 5017 32983 5040 33017
rect 4960 32960 5040 32983
rect 5120 33337 5200 33360
rect 5120 33303 5143 33337
rect 5177 33303 5200 33337
rect 5120 33017 5200 33303
rect 5120 32983 5143 33017
rect 5177 32983 5200 33017
rect 5120 32960 5200 32983
rect 5280 33337 5360 33360
rect 5280 33303 5303 33337
rect 5337 33303 5360 33337
rect 5280 33017 5360 33303
rect 5280 32983 5303 33017
rect 5337 32983 5360 33017
rect 5280 32960 5360 32983
rect 5440 33337 5520 33360
rect 5440 33303 5463 33337
rect 5497 33303 5520 33337
rect 5440 33017 5520 33303
rect 5440 32983 5463 33017
rect 5497 32983 5520 33017
rect 5440 32960 5520 32983
rect 5600 33337 5680 33360
rect 5600 33303 5623 33337
rect 5657 33303 5680 33337
rect 5600 33017 5680 33303
rect 5600 32983 5623 33017
rect 5657 32983 5680 33017
rect 5600 32960 5680 32983
rect 5760 33337 5840 33360
rect 5760 33303 5783 33337
rect 5817 33303 5840 33337
rect 5760 33017 5840 33303
rect 5760 32983 5783 33017
rect 5817 32983 5840 33017
rect 5760 32960 5840 32983
rect 5920 33337 6000 33360
rect 5920 33303 5943 33337
rect 5977 33303 6000 33337
rect 5920 33017 6000 33303
rect 5920 32983 5943 33017
rect 5977 32983 6000 33017
rect 5920 32960 6000 32983
rect 6080 33337 6160 33360
rect 6080 33303 6103 33337
rect 6137 33303 6160 33337
rect 6080 33017 6160 33303
rect 6080 32983 6103 33017
rect 6137 32983 6160 33017
rect 6080 32960 6160 32983
rect 6240 33337 6320 33360
rect 6240 33303 6263 33337
rect 6297 33303 6320 33337
rect 6240 33017 6320 33303
rect 6240 32983 6263 33017
rect 6297 32983 6320 33017
rect 6240 32960 6320 32983
rect 6400 33337 6480 33360
rect 6400 33303 6423 33337
rect 6457 33303 6480 33337
rect 6400 33017 6480 33303
rect 6400 32983 6423 33017
rect 6457 32983 6480 33017
rect 6400 32960 6480 32983
rect 6560 33337 6640 33360
rect 6560 33303 6583 33337
rect 6617 33303 6640 33337
rect 6560 33017 6640 33303
rect 6560 32983 6583 33017
rect 6617 32983 6640 33017
rect 6560 32960 6640 32983
rect 6720 33337 6800 33360
rect 6720 33303 6743 33337
rect 6777 33303 6800 33337
rect 6720 33017 6800 33303
rect 6720 32983 6743 33017
rect 6777 32983 6800 33017
rect 6720 32960 6800 32983
rect 6880 33337 6960 33360
rect 6880 33303 6903 33337
rect 6937 33303 6960 33337
rect 6880 33017 6960 33303
rect 6880 32983 6903 33017
rect 6937 32983 6960 33017
rect 6880 32960 6960 32983
rect 7040 33337 7120 33360
rect 7040 33303 7063 33337
rect 7097 33303 7120 33337
rect 7040 33017 7120 33303
rect 7040 32983 7063 33017
rect 7097 32983 7120 33017
rect 7040 32960 7120 32983
rect 7200 33337 7280 33360
rect 7200 33303 7223 33337
rect 7257 33303 7280 33337
rect 7200 33017 7280 33303
rect 7200 32983 7223 33017
rect 7257 32983 7280 33017
rect 7200 32960 7280 32983
rect 7360 33337 7440 33360
rect 7360 33303 7383 33337
rect 7417 33303 7440 33337
rect 7360 33017 7440 33303
rect 7360 32983 7383 33017
rect 7417 32983 7440 33017
rect 7360 32960 7440 32983
rect 7520 33337 7600 33360
rect 7520 33303 7543 33337
rect 7577 33303 7600 33337
rect 7520 33017 7600 33303
rect 7520 32983 7543 33017
rect 7577 32983 7600 33017
rect 7520 32960 7600 32983
rect 7680 33337 7760 33360
rect 7680 33303 7703 33337
rect 7737 33303 7760 33337
rect 7680 33017 7760 33303
rect 7680 32983 7703 33017
rect 7737 32983 7760 33017
rect 7680 32960 7760 32983
rect 7840 33337 7920 33360
rect 7840 33303 7863 33337
rect 7897 33303 7920 33337
rect 7840 33017 7920 33303
rect 7840 32983 7863 33017
rect 7897 32983 7920 33017
rect 7840 32960 7920 32983
rect 8000 33337 8080 33360
rect 8000 33303 8023 33337
rect 8057 33303 8080 33337
rect 8000 33017 8080 33303
rect 8000 32983 8023 33017
rect 8057 32983 8080 33017
rect 8000 32960 8080 32983
rect 8160 33337 8240 33360
rect 8160 33303 8183 33337
rect 8217 33303 8240 33337
rect 8160 33017 8240 33303
rect 8160 32983 8183 33017
rect 8217 32983 8240 33017
rect 8160 32960 8240 32983
rect 8320 33337 8400 33360
rect 8320 33303 8343 33337
rect 8377 33303 8400 33337
rect 8320 33017 8400 33303
rect 8320 32983 8343 33017
rect 8377 32983 8400 33017
rect 8320 32960 8400 32983
rect 8480 32960 8560 33360
rect 8640 32960 8720 33360
rect 8800 32960 8880 33360
rect 8960 32960 9040 33360
rect 9120 32960 9200 33360
rect 9280 32960 9360 33360
rect 9440 32960 9520 33360
rect 9600 32960 9680 33360
rect 9760 32960 9840 33360
rect 9920 32960 10000 33360
rect 10080 32960 10160 33360
rect 10240 32960 10320 33360
rect 10400 32960 10480 33360
rect 10560 32960 10640 33360
rect 10720 32960 10800 33360
rect 10880 32960 10960 33360
rect 11040 32960 11120 33360
rect 11200 32960 11280 33360
rect 11360 32960 11440 33360
rect 11520 32960 11600 33360
rect 11680 32960 11760 33360
rect 11840 32960 11920 33360
rect 12000 32960 12080 33360
rect 12160 32960 12240 33360
rect 12320 32960 12400 33360
rect 12480 33337 12560 33360
rect 12480 33303 12503 33337
rect 12537 33303 12560 33337
rect 12480 33017 12560 33303
rect 12480 32983 12503 33017
rect 12537 32983 12560 33017
rect 12480 32960 12560 32983
rect 12640 33337 12720 33360
rect 12640 33303 12663 33337
rect 12697 33303 12720 33337
rect 12640 33017 12720 33303
rect 12640 32983 12663 33017
rect 12697 32983 12720 33017
rect 12640 32960 12720 32983
rect 12800 33337 12880 33360
rect 12800 33303 12823 33337
rect 12857 33303 12880 33337
rect 12800 33017 12880 33303
rect 12800 32983 12823 33017
rect 12857 32983 12880 33017
rect 12800 32960 12880 32983
rect 12960 33337 13040 33360
rect 12960 33303 12983 33337
rect 13017 33303 13040 33337
rect 12960 33017 13040 33303
rect 12960 32983 12983 33017
rect 13017 32983 13040 33017
rect 12960 32960 13040 32983
rect 13120 33337 13200 33360
rect 13120 33303 13143 33337
rect 13177 33303 13200 33337
rect 13120 33017 13200 33303
rect 13120 32983 13143 33017
rect 13177 32983 13200 33017
rect 13120 32960 13200 32983
rect 13280 33337 13360 33360
rect 13280 33303 13303 33337
rect 13337 33303 13360 33337
rect 13280 33017 13360 33303
rect 13280 32983 13303 33017
rect 13337 32983 13360 33017
rect 13280 32960 13360 32983
rect 13440 33337 13520 33360
rect 13440 33303 13463 33337
rect 13497 33303 13520 33337
rect 13440 33017 13520 33303
rect 13440 32983 13463 33017
rect 13497 32983 13520 33017
rect 13440 32960 13520 32983
rect 13600 33337 13680 33360
rect 13600 33303 13623 33337
rect 13657 33303 13680 33337
rect 13600 33017 13680 33303
rect 13600 32983 13623 33017
rect 13657 32983 13680 33017
rect 13600 32960 13680 32983
rect 13760 33337 13840 33360
rect 13760 33303 13783 33337
rect 13817 33303 13840 33337
rect 13760 33017 13840 33303
rect 13760 32983 13783 33017
rect 13817 32983 13840 33017
rect 13760 32960 13840 32983
rect 13920 33337 14000 33360
rect 13920 33303 13943 33337
rect 13977 33303 14000 33337
rect 13920 33017 14000 33303
rect 13920 32983 13943 33017
rect 13977 32983 14000 33017
rect 13920 32960 14000 32983
rect 14080 33337 14160 33360
rect 14080 33303 14103 33337
rect 14137 33303 14160 33337
rect 14080 33017 14160 33303
rect 14080 32983 14103 33017
rect 14137 32983 14160 33017
rect 14080 32960 14160 32983
rect 14240 33337 14320 33360
rect 14240 33303 14263 33337
rect 14297 33303 14320 33337
rect 14240 33017 14320 33303
rect 14240 32983 14263 33017
rect 14297 32983 14320 33017
rect 14240 32960 14320 32983
rect 14400 33337 14480 33360
rect 14400 33303 14423 33337
rect 14457 33303 14480 33337
rect 14400 33017 14480 33303
rect 14400 32983 14423 33017
rect 14457 32983 14480 33017
rect 14400 32960 14480 32983
rect 14560 33337 14640 33360
rect 14560 33303 14583 33337
rect 14617 33303 14640 33337
rect 14560 33017 14640 33303
rect 14560 32983 14583 33017
rect 14617 32983 14640 33017
rect 14560 32960 14640 32983
rect 14720 33337 14800 33360
rect 14720 33303 14743 33337
rect 14777 33303 14800 33337
rect 14720 33017 14800 33303
rect 14720 32983 14743 33017
rect 14777 32983 14800 33017
rect 14720 32960 14800 32983
rect 14880 33337 14960 33360
rect 14880 33303 14903 33337
rect 14937 33303 14960 33337
rect 14880 33017 14960 33303
rect 14880 32983 14903 33017
rect 14937 32983 14960 33017
rect 14880 32960 14960 32983
rect 15040 33337 15120 33360
rect 15040 33303 15063 33337
rect 15097 33303 15120 33337
rect 15040 33017 15120 33303
rect 15040 32983 15063 33017
rect 15097 32983 15120 33017
rect 15040 32960 15120 32983
rect 15200 33337 15280 33360
rect 15200 33303 15223 33337
rect 15257 33303 15280 33337
rect 15200 33017 15280 33303
rect 15200 32983 15223 33017
rect 15257 32983 15280 33017
rect 15200 32960 15280 32983
rect 15360 33337 15440 33360
rect 15360 33303 15383 33337
rect 15417 33303 15440 33337
rect 15360 33017 15440 33303
rect 15360 32983 15383 33017
rect 15417 32983 15440 33017
rect 15360 32960 15440 32983
rect 15520 33337 15600 33360
rect 15520 33303 15543 33337
rect 15577 33303 15600 33337
rect 15520 33017 15600 33303
rect 15520 32983 15543 33017
rect 15577 32983 15600 33017
rect 15520 32960 15600 32983
rect 15680 33337 15760 33360
rect 15680 33303 15703 33337
rect 15737 33303 15760 33337
rect 15680 33017 15760 33303
rect 15680 32983 15703 33017
rect 15737 32983 15760 33017
rect 15680 32960 15760 32983
rect 15840 33337 15920 33360
rect 15840 33303 15863 33337
rect 15897 33303 15920 33337
rect 15840 33017 15920 33303
rect 15840 32983 15863 33017
rect 15897 32983 15920 33017
rect 15840 32960 15920 32983
rect 16000 33337 16080 33360
rect 16000 33303 16023 33337
rect 16057 33303 16080 33337
rect 16000 33017 16080 33303
rect 16000 32983 16023 33017
rect 16057 32983 16080 33017
rect 16000 32960 16080 32983
rect 16160 33337 16240 33360
rect 16160 33303 16183 33337
rect 16217 33303 16240 33337
rect 16160 33017 16240 33303
rect 16160 32983 16183 33017
rect 16217 32983 16240 33017
rect 16160 32960 16240 32983
rect 16320 33337 16400 33360
rect 16320 33303 16343 33337
rect 16377 33303 16400 33337
rect 16320 33017 16400 33303
rect 16320 32983 16343 33017
rect 16377 32983 16400 33017
rect 16320 32960 16400 32983
rect 16480 33337 16560 33360
rect 16480 33303 16503 33337
rect 16537 33303 16560 33337
rect 16480 33017 16560 33303
rect 16480 32983 16503 33017
rect 16537 32983 16560 33017
rect 16480 32960 16560 32983
rect 16640 33337 16720 33360
rect 16640 33303 16663 33337
rect 16697 33303 16720 33337
rect 16640 33017 16720 33303
rect 16640 32983 16663 33017
rect 16697 32983 16720 33017
rect 16640 32960 16720 32983
rect 16800 33337 16880 33360
rect 16800 33303 16823 33337
rect 16857 33303 16880 33337
rect 16800 33017 16880 33303
rect 16800 32983 16823 33017
rect 16857 32983 16880 33017
rect 16800 32960 16880 32983
rect 16960 33337 17040 33360
rect 16960 33303 16983 33337
rect 17017 33303 17040 33337
rect 16960 33017 17040 33303
rect 16960 32983 16983 33017
rect 17017 32983 17040 33017
rect 16960 32960 17040 32983
rect 17120 33337 17200 33360
rect 17120 33303 17143 33337
rect 17177 33303 17200 33337
rect 17120 33017 17200 33303
rect 17120 32983 17143 33017
rect 17177 32983 17200 33017
rect 17120 32960 17200 32983
rect 17280 33337 17360 33360
rect 17280 33303 17303 33337
rect 17337 33303 17360 33337
rect 17280 33017 17360 33303
rect 17280 32983 17303 33017
rect 17337 32983 17360 33017
rect 17280 32960 17360 32983
rect 17440 33337 17520 33360
rect 17440 33303 17463 33337
rect 17497 33303 17520 33337
rect 17440 33017 17520 33303
rect 17440 32983 17463 33017
rect 17497 32983 17520 33017
rect 17440 32960 17520 32983
rect 17600 33337 17680 33360
rect 17600 33303 17623 33337
rect 17657 33303 17680 33337
rect 17600 33017 17680 33303
rect 17600 32983 17623 33017
rect 17657 32983 17680 33017
rect 17600 32960 17680 32983
rect 17760 33337 17840 33360
rect 17760 33303 17783 33337
rect 17817 33303 17840 33337
rect 17760 33017 17840 33303
rect 17760 32983 17783 33017
rect 17817 32983 17840 33017
rect 17760 32960 17840 32983
rect 17920 33337 18000 33360
rect 17920 33303 17943 33337
rect 17977 33303 18000 33337
rect 17920 33017 18000 33303
rect 17920 32983 17943 33017
rect 17977 32983 18000 33017
rect 17920 32960 18000 32983
rect 18080 33337 18160 33360
rect 18080 33303 18103 33337
rect 18137 33303 18160 33337
rect 18080 33017 18160 33303
rect 18080 32983 18103 33017
rect 18137 32983 18160 33017
rect 18080 32960 18160 32983
rect 18240 33337 18320 33360
rect 18240 33303 18263 33337
rect 18297 33303 18320 33337
rect 18240 33017 18320 33303
rect 18240 32983 18263 33017
rect 18297 32983 18320 33017
rect 18240 32960 18320 32983
rect 18400 33337 18480 33360
rect 18400 33303 18423 33337
rect 18457 33303 18480 33337
rect 18400 33017 18480 33303
rect 18400 32983 18423 33017
rect 18457 32983 18480 33017
rect 18400 32960 18480 32983
rect 18560 33337 18640 33360
rect 18560 33303 18583 33337
rect 18617 33303 18640 33337
rect 18560 33017 18640 33303
rect 18560 32983 18583 33017
rect 18617 32983 18640 33017
rect 18560 32960 18640 32983
rect 18720 33337 18800 33360
rect 18720 33303 18743 33337
rect 18777 33303 18800 33337
rect 18720 33017 18800 33303
rect 18720 32983 18743 33017
rect 18777 32983 18800 33017
rect 18720 32960 18800 32983
rect 18880 33337 18960 33360
rect 18880 33303 18903 33337
rect 18937 33303 18960 33337
rect 18880 33017 18960 33303
rect 18880 32983 18903 33017
rect 18937 32983 18960 33017
rect 18880 32960 18960 32983
rect 19040 32960 19120 33360
rect 19200 32960 19280 33360
rect 19360 32960 19440 33360
rect 19520 32960 19600 33360
rect 19680 32960 19760 33360
rect 19840 32960 19920 33360
rect 20000 32960 20080 33360
rect 20160 32960 20240 33360
rect 20320 32960 20400 33360
rect 20480 32960 20560 33360
rect 20640 32960 20720 33360
rect 20800 32960 20880 33360
rect 20960 32960 21040 33360
rect 21120 32960 21200 33360
rect 21280 32960 21360 33360
rect 21440 32960 21520 33360
rect 21600 32960 21680 33360
rect 21760 32960 21840 33360
rect 21920 32960 22000 33360
rect 22080 32960 22160 33360
rect 22240 32960 22320 33360
rect 22400 32960 22480 33360
rect 22560 32960 22640 33360
rect 22720 32960 22800 33360
rect 22880 32960 22960 33360
rect 23120 33337 23200 33360
rect 23120 33303 23143 33337
rect 23177 33303 23200 33337
rect 23120 33017 23200 33303
rect 23120 32983 23143 33017
rect 23177 32983 23200 33017
rect 23120 32960 23200 32983
rect 23280 33337 23360 33360
rect 23280 33303 23303 33337
rect 23337 33303 23360 33337
rect 23280 33017 23360 33303
rect 23280 32983 23303 33017
rect 23337 32983 23360 33017
rect 23280 32960 23360 32983
rect 23440 33337 23520 33360
rect 23440 33303 23463 33337
rect 23497 33303 23520 33337
rect 23440 33017 23520 33303
rect 23440 32983 23463 33017
rect 23497 32983 23520 33017
rect 23440 32960 23520 32983
rect 23600 33337 23680 33360
rect 23600 33303 23623 33337
rect 23657 33303 23680 33337
rect 23600 33017 23680 33303
rect 23600 32983 23623 33017
rect 23657 32983 23680 33017
rect 23600 32960 23680 32983
rect 23760 33337 23840 33360
rect 23760 33303 23783 33337
rect 23817 33303 23840 33337
rect 23760 33017 23840 33303
rect 23760 32983 23783 33017
rect 23817 32983 23840 33017
rect 23760 32960 23840 32983
rect 23920 33337 24000 33360
rect 23920 33303 23943 33337
rect 23977 33303 24000 33337
rect 23920 33017 24000 33303
rect 23920 32983 23943 33017
rect 23977 32983 24000 33017
rect 23920 32960 24000 32983
rect 24080 33337 24160 33360
rect 24080 33303 24103 33337
rect 24137 33303 24160 33337
rect 24080 33017 24160 33303
rect 24080 32983 24103 33017
rect 24137 32983 24160 33017
rect 24080 32960 24160 32983
rect 24240 33337 24320 33360
rect 24240 33303 24263 33337
rect 24297 33303 24320 33337
rect 24240 33017 24320 33303
rect 24240 32983 24263 33017
rect 24297 32983 24320 33017
rect 24240 32960 24320 32983
rect 24400 33337 24480 33360
rect 24400 33303 24423 33337
rect 24457 33303 24480 33337
rect 24400 33017 24480 33303
rect 24400 32983 24423 33017
rect 24457 32983 24480 33017
rect 24400 32960 24480 32983
rect 24560 33337 24640 33360
rect 24560 33303 24583 33337
rect 24617 33303 24640 33337
rect 24560 33017 24640 33303
rect 24560 32983 24583 33017
rect 24617 32983 24640 33017
rect 24560 32960 24640 32983
rect 24720 33337 24800 33360
rect 24720 33303 24743 33337
rect 24777 33303 24800 33337
rect 24720 33017 24800 33303
rect 24720 32983 24743 33017
rect 24777 32983 24800 33017
rect 24720 32960 24800 32983
rect 24880 33337 24960 33360
rect 24880 33303 24903 33337
rect 24937 33303 24960 33337
rect 24880 33017 24960 33303
rect 24880 32983 24903 33017
rect 24937 32983 24960 33017
rect 24880 32960 24960 32983
rect 25040 33337 25120 33360
rect 25040 33303 25063 33337
rect 25097 33303 25120 33337
rect 25040 33017 25120 33303
rect 25040 32983 25063 33017
rect 25097 32983 25120 33017
rect 25040 32960 25120 32983
rect 25200 33337 25280 33360
rect 25200 33303 25223 33337
rect 25257 33303 25280 33337
rect 25200 33017 25280 33303
rect 25200 32983 25223 33017
rect 25257 32983 25280 33017
rect 25200 32960 25280 32983
rect 25360 33337 25440 33360
rect 25360 33303 25383 33337
rect 25417 33303 25440 33337
rect 25360 33017 25440 33303
rect 25360 32983 25383 33017
rect 25417 32983 25440 33017
rect 25360 32960 25440 32983
rect 25520 33337 25600 33360
rect 25520 33303 25543 33337
rect 25577 33303 25600 33337
rect 25520 33017 25600 33303
rect 25520 32983 25543 33017
rect 25577 32983 25600 33017
rect 25520 32960 25600 32983
rect 25680 33337 25760 33360
rect 25680 33303 25703 33337
rect 25737 33303 25760 33337
rect 25680 33017 25760 33303
rect 25680 32983 25703 33017
rect 25737 32983 25760 33017
rect 25680 32960 25760 32983
rect 25840 33337 25920 33360
rect 25840 33303 25863 33337
rect 25897 33303 25920 33337
rect 25840 33017 25920 33303
rect 25840 32983 25863 33017
rect 25897 32983 25920 33017
rect 25840 32960 25920 32983
rect 26000 33337 26080 33360
rect 26000 33303 26023 33337
rect 26057 33303 26080 33337
rect 26000 33017 26080 33303
rect 26000 32983 26023 33017
rect 26057 32983 26080 33017
rect 26000 32960 26080 32983
rect 26160 33337 26240 33360
rect 26160 33303 26183 33337
rect 26217 33303 26240 33337
rect 26160 33017 26240 33303
rect 26160 32983 26183 33017
rect 26217 32983 26240 33017
rect 26160 32960 26240 32983
rect 26320 33337 26400 33360
rect 26320 33303 26343 33337
rect 26377 33303 26400 33337
rect 26320 33017 26400 33303
rect 26320 32983 26343 33017
rect 26377 32983 26400 33017
rect 26320 32960 26400 32983
rect 26480 33337 26560 33360
rect 26480 33303 26503 33337
rect 26537 33303 26560 33337
rect 26480 33017 26560 33303
rect 26480 32983 26503 33017
rect 26537 32983 26560 33017
rect 26480 32960 26560 32983
rect 26640 33337 26720 33360
rect 26640 33303 26663 33337
rect 26697 33303 26720 33337
rect 26640 33017 26720 33303
rect 26640 32983 26663 33017
rect 26697 32983 26720 33017
rect 26640 32960 26720 32983
rect 26800 33337 26880 33360
rect 26800 33303 26823 33337
rect 26857 33303 26880 33337
rect 26800 33017 26880 33303
rect 26800 32983 26823 33017
rect 26857 32983 26880 33017
rect 26800 32960 26880 32983
rect 26960 33337 27040 33360
rect 26960 33303 26983 33337
rect 27017 33303 27040 33337
rect 26960 33017 27040 33303
rect 26960 32983 26983 33017
rect 27017 32983 27040 33017
rect 26960 32960 27040 32983
rect 27120 33337 27200 33360
rect 27120 33303 27143 33337
rect 27177 33303 27200 33337
rect 27120 33017 27200 33303
rect 27120 32983 27143 33017
rect 27177 32983 27200 33017
rect 27120 32960 27200 32983
rect 27280 33337 27360 33360
rect 27280 33303 27303 33337
rect 27337 33303 27360 33337
rect 27280 33017 27360 33303
rect 27280 32983 27303 33017
rect 27337 32983 27360 33017
rect 27280 32960 27360 32983
rect 27440 33337 27520 33360
rect 27440 33303 27463 33337
rect 27497 33303 27520 33337
rect 27440 33017 27520 33303
rect 27440 32983 27463 33017
rect 27497 32983 27520 33017
rect 27440 32960 27520 32983
rect 27600 33337 27680 33360
rect 27600 33303 27623 33337
rect 27657 33303 27680 33337
rect 27600 33017 27680 33303
rect 27600 32983 27623 33017
rect 27657 32983 27680 33017
rect 27600 32960 27680 32983
rect 27760 33337 27840 33360
rect 27760 33303 27783 33337
rect 27817 33303 27840 33337
rect 27760 33017 27840 33303
rect 27760 32983 27783 33017
rect 27817 32983 27840 33017
rect 27760 32960 27840 32983
rect 27920 33337 28000 33360
rect 27920 33303 27943 33337
rect 27977 33303 28000 33337
rect 27920 33017 28000 33303
rect 27920 32983 27943 33017
rect 27977 32983 28000 33017
rect 27920 32960 28000 32983
rect 28080 33337 28160 33360
rect 28080 33303 28103 33337
rect 28137 33303 28160 33337
rect 28080 33017 28160 33303
rect 28080 32983 28103 33017
rect 28137 32983 28160 33017
rect 28080 32960 28160 32983
rect 28240 33337 28320 33360
rect 28240 33303 28263 33337
rect 28297 33303 28320 33337
rect 28240 33017 28320 33303
rect 28240 32983 28263 33017
rect 28297 32983 28320 33017
rect 28240 32960 28320 32983
rect 28400 33337 28480 33360
rect 28400 33303 28423 33337
rect 28457 33303 28480 33337
rect 28400 33017 28480 33303
rect 28400 32983 28423 33017
rect 28457 32983 28480 33017
rect 28400 32960 28480 32983
rect 28560 33337 28640 33360
rect 28560 33303 28583 33337
rect 28617 33303 28640 33337
rect 28560 33017 28640 33303
rect 28560 32983 28583 33017
rect 28617 32983 28640 33017
rect 28560 32960 28640 32983
rect 28720 33337 28800 33360
rect 28720 33303 28743 33337
rect 28777 33303 28800 33337
rect 28720 33017 28800 33303
rect 28720 32983 28743 33017
rect 28777 32983 28800 33017
rect 28720 32960 28800 32983
rect 28880 33337 28960 33360
rect 28880 33303 28903 33337
rect 28937 33303 28960 33337
rect 28880 33017 28960 33303
rect 28880 32983 28903 33017
rect 28937 32983 28960 33017
rect 28880 32960 28960 32983
rect 29040 33337 29120 33360
rect 29040 33303 29063 33337
rect 29097 33303 29120 33337
rect 29040 33017 29120 33303
rect 29040 32983 29063 33017
rect 29097 32983 29120 33017
rect 29040 32960 29120 32983
rect 29200 33337 29280 33360
rect 29200 33303 29223 33337
rect 29257 33303 29280 33337
rect 29200 33017 29280 33303
rect 29200 32983 29223 33017
rect 29257 32983 29280 33017
rect 29200 32960 29280 32983
rect 29360 33337 29440 33360
rect 29360 33303 29383 33337
rect 29417 33303 29440 33337
rect 29360 33017 29440 33303
rect 29360 32983 29383 33017
rect 29417 32983 29440 33017
rect 29360 32960 29440 32983
rect 29520 32960 29600 33360
rect 29680 32960 29760 33360
rect 29840 32960 29920 33360
rect 30000 32960 30080 33360
rect 30160 32960 30240 33360
rect 30320 32960 30400 33360
rect 30480 32960 30560 33360
rect 30640 32960 30720 33360
rect 30800 32960 30880 33360
rect 30960 32960 31040 33360
rect 31120 32960 31200 33360
rect 31280 32960 31360 33360
rect 31440 32960 31520 33360
rect 31600 32960 31680 33360
rect 31760 32960 31840 33360
rect 31920 32960 32000 33360
rect 32080 32960 32160 33360
rect 32240 32960 32320 33360
rect 32400 32960 32480 33360
rect 32560 32960 32640 33360
rect 32720 32960 32800 33360
rect 32880 32960 32960 33360
rect 33040 32960 33120 33360
rect 33200 32960 33280 33360
rect 33360 32960 33440 33360
rect 33520 33337 33600 33360
rect 33520 33303 33543 33337
rect 33577 33303 33600 33337
rect 33520 33017 33600 33303
rect 33520 32983 33543 33017
rect 33577 32983 33600 33017
rect 33520 32960 33600 32983
rect 33680 33337 33760 33360
rect 33680 33303 33703 33337
rect 33737 33303 33760 33337
rect 33680 33017 33760 33303
rect 33680 32983 33703 33017
rect 33737 32983 33760 33017
rect 33680 32960 33760 32983
rect 33840 33337 33920 33360
rect 33840 33303 33863 33337
rect 33897 33303 33920 33337
rect 33840 33017 33920 33303
rect 33840 32983 33863 33017
rect 33897 32983 33920 33017
rect 33840 32960 33920 32983
rect 34000 33337 34080 33360
rect 34000 33303 34023 33337
rect 34057 33303 34080 33337
rect 34000 33017 34080 33303
rect 34000 32983 34023 33017
rect 34057 32983 34080 33017
rect 34000 32960 34080 32983
rect 34160 33337 34240 33360
rect 34160 33303 34183 33337
rect 34217 33303 34240 33337
rect 34160 33017 34240 33303
rect 34160 32983 34183 33017
rect 34217 32983 34240 33017
rect 34160 32960 34240 32983
rect 34320 33337 34400 33360
rect 34320 33303 34343 33337
rect 34377 33303 34400 33337
rect 34320 33017 34400 33303
rect 34320 32983 34343 33017
rect 34377 32983 34400 33017
rect 34320 32960 34400 32983
rect 34480 33337 34560 33360
rect 34480 33303 34503 33337
rect 34537 33303 34560 33337
rect 34480 33017 34560 33303
rect 34480 32983 34503 33017
rect 34537 32983 34560 33017
rect 34480 32960 34560 32983
rect 34640 33337 34720 33360
rect 34640 33303 34663 33337
rect 34697 33303 34720 33337
rect 34640 33017 34720 33303
rect 34640 32983 34663 33017
rect 34697 32983 34720 33017
rect 34640 32960 34720 32983
rect 34800 33337 34880 33360
rect 34800 33303 34823 33337
rect 34857 33303 34880 33337
rect 34800 33017 34880 33303
rect 34800 32983 34823 33017
rect 34857 32983 34880 33017
rect 34800 32960 34880 32983
rect 34960 33337 35040 33360
rect 34960 33303 34983 33337
rect 35017 33303 35040 33337
rect 34960 33017 35040 33303
rect 34960 32983 34983 33017
rect 35017 32983 35040 33017
rect 34960 32960 35040 32983
rect 35120 33337 35200 33360
rect 35120 33303 35143 33337
rect 35177 33303 35200 33337
rect 35120 33017 35200 33303
rect 35120 32983 35143 33017
rect 35177 32983 35200 33017
rect 35120 32960 35200 32983
rect 35280 33337 35360 33360
rect 35280 33303 35303 33337
rect 35337 33303 35360 33337
rect 35280 33017 35360 33303
rect 35280 32983 35303 33017
rect 35337 32983 35360 33017
rect 35280 32960 35360 32983
rect 35440 33337 35520 33360
rect 35440 33303 35463 33337
rect 35497 33303 35520 33337
rect 35440 33017 35520 33303
rect 35440 32983 35463 33017
rect 35497 32983 35520 33017
rect 35440 32960 35520 32983
rect 35600 33337 35680 33360
rect 35600 33303 35623 33337
rect 35657 33303 35680 33337
rect 35600 33017 35680 33303
rect 35600 32983 35623 33017
rect 35657 32983 35680 33017
rect 35600 32960 35680 32983
rect 35760 33337 35840 33360
rect 35760 33303 35783 33337
rect 35817 33303 35840 33337
rect 35760 33017 35840 33303
rect 35760 32983 35783 33017
rect 35817 32983 35840 33017
rect 35760 32960 35840 32983
rect 35920 33337 36000 33360
rect 35920 33303 35943 33337
rect 35977 33303 36000 33337
rect 35920 33017 36000 33303
rect 35920 32983 35943 33017
rect 35977 32983 36000 33017
rect 35920 32960 36000 32983
rect 36080 33337 36160 33360
rect 36080 33303 36103 33337
rect 36137 33303 36160 33337
rect 36080 33017 36160 33303
rect 36080 32983 36103 33017
rect 36137 32983 36160 33017
rect 36080 32960 36160 32983
rect 36240 33337 36320 33360
rect 36240 33303 36263 33337
rect 36297 33303 36320 33337
rect 36240 33017 36320 33303
rect 36240 32983 36263 33017
rect 36297 32983 36320 33017
rect 36240 32960 36320 32983
rect 36400 33337 36480 33360
rect 36400 33303 36423 33337
rect 36457 33303 36480 33337
rect 36400 33017 36480 33303
rect 36400 32983 36423 33017
rect 36457 32983 36480 33017
rect 36400 32960 36480 32983
rect 36560 33337 36640 33360
rect 36560 33303 36583 33337
rect 36617 33303 36640 33337
rect 36560 33017 36640 33303
rect 36560 32983 36583 33017
rect 36617 32983 36640 33017
rect 36560 32960 36640 32983
rect 36720 33337 36800 33360
rect 36720 33303 36743 33337
rect 36777 33303 36800 33337
rect 36720 33017 36800 33303
rect 36720 32983 36743 33017
rect 36777 32983 36800 33017
rect 36720 32960 36800 32983
rect 36880 33337 36960 33360
rect 36880 33303 36903 33337
rect 36937 33303 36960 33337
rect 36880 33017 36960 33303
rect 36880 32983 36903 33017
rect 36937 32983 36960 33017
rect 36880 32960 36960 32983
rect 37040 33337 37120 33360
rect 37040 33303 37063 33337
rect 37097 33303 37120 33337
rect 37040 33017 37120 33303
rect 37040 32983 37063 33017
rect 37097 32983 37120 33017
rect 37040 32960 37120 32983
rect 37200 33337 37280 33360
rect 37200 33303 37223 33337
rect 37257 33303 37280 33337
rect 37200 33017 37280 33303
rect 37200 32983 37223 33017
rect 37257 32983 37280 33017
rect 37200 32960 37280 32983
rect 37360 33337 37440 33360
rect 37360 33303 37383 33337
rect 37417 33303 37440 33337
rect 37360 33017 37440 33303
rect 37360 32983 37383 33017
rect 37417 32983 37440 33017
rect 37360 32960 37440 32983
rect 37520 33337 37600 33360
rect 37520 33303 37543 33337
rect 37577 33303 37600 33337
rect 37520 33017 37600 33303
rect 37520 32983 37543 33017
rect 37577 32983 37600 33017
rect 37520 32960 37600 32983
rect 37680 33337 37760 33360
rect 37680 33303 37703 33337
rect 37737 33303 37760 33337
rect 37680 33017 37760 33303
rect 37680 32983 37703 33017
rect 37737 32983 37760 33017
rect 37680 32960 37760 32983
rect 37840 33337 37920 33360
rect 37840 33303 37863 33337
rect 37897 33303 37920 33337
rect 37840 33017 37920 33303
rect 37840 32983 37863 33017
rect 37897 32983 37920 33017
rect 37840 32960 37920 32983
rect 38000 33337 38080 33360
rect 38000 33303 38023 33337
rect 38057 33303 38080 33337
rect 38000 33017 38080 33303
rect 38000 32983 38023 33017
rect 38057 32983 38080 33017
rect 38000 32960 38080 32983
rect 38160 33337 38240 33360
rect 38160 33303 38183 33337
rect 38217 33303 38240 33337
rect 38160 33017 38240 33303
rect 38160 32983 38183 33017
rect 38217 32983 38240 33017
rect 38160 32960 38240 32983
rect 38320 33337 38400 33360
rect 38320 33303 38343 33337
rect 38377 33303 38400 33337
rect 38320 33017 38400 33303
rect 38320 32983 38343 33017
rect 38377 32983 38400 33017
rect 38320 32960 38400 32983
rect 38480 33337 38560 33360
rect 38480 33303 38503 33337
rect 38537 33303 38560 33337
rect 38480 33017 38560 33303
rect 38480 32983 38503 33017
rect 38537 32983 38560 33017
rect 38480 32960 38560 32983
rect 38640 33337 38720 33360
rect 38640 33303 38663 33337
rect 38697 33303 38720 33337
rect 38640 33017 38720 33303
rect 38640 32983 38663 33017
rect 38697 32983 38720 33017
rect 38640 32960 38720 32983
rect 38800 33337 38880 33360
rect 38800 33303 38823 33337
rect 38857 33303 38880 33337
rect 38800 33017 38880 33303
rect 38800 32983 38823 33017
rect 38857 32983 38880 33017
rect 38800 32960 38880 32983
rect 38960 33337 39040 33360
rect 38960 33303 38983 33337
rect 39017 33303 39040 33337
rect 38960 33017 39040 33303
rect 38960 32983 38983 33017
rect 39017 32983 39040 33017
rect 38960 32960 39040 32983
rect 39120 33337 39200 33360
rect 39120 33303 39143 33337
rect 39177 33303 39200 33337
rect 39120 33017 39200 33303
rect 39120 32983 39143 33017
rect 39177 32983 39200 33017
rect 39120 32960 39200 32983
rect 39280 33337 39360 33360
rect 39280 33303 39303 33337
rect 39337 33303 39360 33337
rect 39280 33017 39360 33303
rect 39280 32983 39303 33017
rect 39337 32983 39360 33017
rect 39280 32960 39360 32983
rect 39440 33337 39520 33360
rect 39440 33303 39463 33337
rect 39497 33303 39520 33337
rect 39440 33017 39520 33303
rect 39440 32983 39463 33017
rect 39497 32983 39520 33017
rect 39440 32960 39520 32983
rect 39600 33337 39680 33360
rect 39600 33303 39623 33337
rect 39657 33303 39680 33337
rect 39600 33017 39680 33303
rect 39600 32983 39623 33017
rect 39657 32983 39680 33017
rect 39600 32960 39680 32983
rect 39760 33337 39840 33360
rect 39760 33303 39783 33337
rect 39817 33303 39840 33337
rect 39760 33017 39840 33303
rect 39760 32983 39783 33017
rect 39817 32983 39840 33017
rect 39760 32960 39840 32983
rect 39920 33337 40000 33360
rect 39920 33303 39943 33337
rect 39977 33303 40000 33337
rect 39920 33017 40000 33303
rect 39920 32983 39943 33017
rect 39977 32983 40000 33017
rect 39920 32960 40000 32983
rect 40080 33337 40160 33360
rect 40080 33303 40103 33337
rect 40137 33303 40160 33337
rect 40080 33017 40160 33303
rect 40080 32983 40103 33017
rect 40137 32983 40160 33017
rect 40080 32960 40160 32983
rect 40240 33337 40320 33360
rect 40240 33303 40263 33337
rect 40297 33303 40320 33337
rect 40240 33017 40320 33303
rect 40240 32983 40263 33017
rect 40297 32983 40320 33017
rect 40240 32960 40320 32983
rect 40400 33337 40480 33360
rect 40400 33303 40423 33337
rect 40457 33303 40480 33337
rect 40400 33017 40480 33303
rect 40400 32983 40423 33017
rect 40457 32983 40480 33017
rect 40400 32960 40480 32983
rect 40560 33337 40640 33360
rect 40560 33303 40583 33337
rect 40617 33303 40640 33337
rect 40560 33017 40640 33303
rect 40560 32983 40583 33017
rect 40617 32983 40640 33017
rect 40560 32960 40640 32983
rect 40720 33337 40800 33360
rect 40720 33303 40743 33337
rect 40777 33303 40800 33337
rect 40720 33017 40800 33303
rect 40720 32983 40743 33017
rect 40777 32983 40800 33017
rect 40720 32960 40800 32983
rect 40880 33337 40960 33360
rect 40880 33303 40903 33337
rect 40937 33303 40960 33337
rect 40880 33017 40960 33303
rect 40880 32983 40903 33017
rect 40937 32983 40960 33017
rect 40880 32960 40960 32983
rect 41040 33337 41120 33360
rect 41040 33303 41063 33337
rect 41097 33303 41120 33337
rect 41040 33017 41120 33303
rect 41040 32983 41063 33017
rect 41097 32983 41120 33017
rect 41040 32960 41120 32983
rect 41200 33337 41280 33360
rect 41200 33303 41223 33337
rect 41257 33303 41280 33337
rect 41200 33017 41280 33303
rect 41200 32983 41223 33017
rect 41257 32983 41280 33017
rect 41200 32960 41280 32983
rect 41360 33337 41440 33360
rect 41360 33303 41383 33337
rect 41417 33303 41440 33337
rect 41360 33017 41440 33303
rect 41360 32983 41383 33017
rect 41417 32983 41440 33017
rect 41360 32960 41440 32983
rect 41520 33337 41600 33360
rect 41520 33303 41543 33337
rect 41577 33303 41600 33337
rect 41520 33017 41600 33303
rect 41520 32983 41543 33017
rect 41577 32983 41600 33017
rect 41520 32960 41600 32983
rect 41680 33337 41760 33360
rect 41680 33303 41703 33337
rect 41737 33303 41760 33337
rect 41680 33017 41760 33303
rect 41680 32983 41703 33017
rect 41737 32983 41760 33017
rect 41680 32960 41760 32983
rect 41840 33337 41920 33360
rect 41840 33303 41863 33337
rect 41897 33303 41920 33337
rect 41840 33017 41920 33303
rect 41840 32983 41863 33017
rect 41897 32983 41920 33017
rect 41840 32960 41920 32983
rect 0 32857 80 32880
rect 0 32823 23 32857
rect 57 32823 80 32857
rect 0 32537 80 32823
rect 0 32503 23 32537
rect 57 32503 80 32537
rect 0 32480 80 32503
rect 160 32857 240 32880
rect 160 32823 183 32857
rect 217 32823 240 32857
rect 160 32537 240 32823
rect 160 32503 183 32537
rect 217 32503 240 32537
rect 160 32480 240 32503
rect 320 32857 400 32880
rect 320 32823 343 32857
rect 377 32823 400 32857
rect 320 32537 400 32823
rect 320 32503 343 32537
rect 377 32503 400 32537
rect 320 32480 400 32503
rect 480 32857 560 32880
rect 480 32823 503 32857
rect 537 32823 560 32857
rect 480 32537 560 32823
rect 480 32503 503 32537
rect 537 32503 560 32537
rect 480 32480 560 32503
rect 640 32857 720 32880
rect 640 32823 663 32857
rect 697 32823 720 32857
rect 640 32537 720 32823
rect 640 32503 663 32537
rect 697 32503 720 32537
rect 640 32480 720 32503
rect 800 32857 880 32880
rect 800 32823 823 32857
rect 857 32823 880 32857
rect 800 32537 880 32823
rect 800 32503 823 32537
rect 857 32503 880 32537
rect 800 32480 880 32503
rect 960 32857 1040 32880
rect 960 32823 983 32857
rect 1017 32823 1040 32857
rect 960 32537 1040 32823
rect 960 32503 983 32537
rect 1017 32503 1040 32537
rect 960 32480 1040 32503
rect 1120 32857 1200 32880
rect 1120 32823 1143 32857
rect 1177 32823 1200 32857
rect 1120 32537 1200 32823
rect 1120 32503 1143 32537
rect 1177 32503 1200 32537
rect 1120 32480 1200 32503
rect 1280 32857 1360 32880
rect 1280 32823 1303 32857
rect 1337 32823 1360 32857
rect 1280 32537 1360 32823
rect 1280 32503 1303 32537
rect 1337 32503 1360 32537
rect 1280 32480 1360 32503
rect 1440 32857 1520 32880
rect 1440 32823 1463 32857
rect 1497 32823 1520 32857
rect 1440 32537 1520 32823
rect 1440 32503 1463 32537
rect 1497 32503 1520 32537
rect 1440 32480 1520 32503
rect 1600 32857 1680 32880
rect 1600 32823 1623 32857
rect 1657 32823 1680 32857
rect 1600 32537 1680 32823
rect 1600 32503 1623 32537
rect 1657 32503 1680 32537
rect 1600 32480 1680 32503
rect 1760 32857 1840 32880
rect 1760 32823 1783 32857
rect 1817 32823 1840 32857
rect 1760 32537 1840 32823
rect 1760 32503 1783 32537
rect 1817 32503 1840 32537
rect 1760 32480 1840 32503
rect 1920 32857 2000 32880
rect 1920 32823 1943 32857
rect 1977 32823 2000 32857
rect 1920 32537 2000 32823
rect 1920 32503 1943 32537
rect 1977 32503 2000 32537
rect 1920 32480 2000 32503
rect 2080 32857 2160 32880
rect 2080 32823 2103 32857
rect 2137 32823 2160 32857
rect 2080 32537 2160 32823
rect 2080 32503 2103 32537
rect 2137 32503 2160 32537
rect 2080 32480 2160 32503
rect 2240 32857 2320 32880
rect 2240 32823 2263 32857
rect 2297 32823 2320 32857
rect 2240 32537 2320 32823
rect 2240 32503 2263 32537
rect 2297 32503 2320 32537
rect 2240 32480 2320 32503
rect 2400 32857 2480 32880
rect 2400 32823 2423 32857
rect 2457 32823 2480 32857
rect 2400 32537 2480 32823
rect 2400 32503 2423 32537
rect 2457 32503 2480 32537
rect 2400 32480 2480 32503
rect 2560 32857 2640 32880
rect 2560 32823 2583 32857
rect 2617 32823 2640 32857
rect 2560 32537 2640 32823
rect 2560 32503 2583 32537
rect 2617 32503 2640 32537
rect 2560 32480 2640 32503
rect 2720 32857 2800 32880
rect 2720 32823 2743 32857
rect 2777 32823 2800 32857
rect 2720 32537 2800 32823
rect 2720 32503 2743 32537
rect 2777 32503 2800 32537
rect 2720 32480 2800 32503
rect 2880 32857 2960 32880
rect 2880 32823 2903 32857
rect 2937 32823 2960 32857
rect 2880 32537 2960 32823
rect 2880 32503 2903 32537
rect 2937 32503 2960 32537
rect 2880 32480 2960 32503
rect 3040 32857 3120 32880
rect 3040 32823 3063 32857
rect 3097 32823 3120 32857
rect 3040 32537 3120 32823
rect 3040 32503 3063 32537
rect 3097 32503 3120 32537
rect 3040 32480 3120 32503
rect 3200 32857 3280 32880
rect 3200 32823 3223 32857
rect 3257 32823 3280 32857
rect 3200 32537 3280 32823
rect 3200 32503 3223 32537
rect 3257 32503 3280 32537
rect 3200 32480 3280 32503
rect 3360 32857 3440 32880
rect 3360 32823 3383 32857
rect 3417 32823 3440 32857
rect 3360 32537 3440 32823
rect 3360 32503 3383 32537
rect 3417 32503 3440 32537
rect 3360 32480 3440 32503
rect 3520 32857 3600 32880
rect 3520 32823 3543 32857
rect 3577 32823 3600 32857
rect 3520 32537 3600 32823
rect 3520 32503 3543 32537
rect 3577 32503 3600 32537
rect 3520 32480 3600 32503
rect 3680 32857 3760 32880
rect 3680 32823 3703 32857
rect 3737 32823 3760 32857
rect 3680 32537 3760 32823
rect 3680 32503 3703 32537
rect 3737 32503 3760 32537
rect 3680 32480 3760 32503
rect 3840 32857 3920 32880
rect 3840 32823 3863 32857
rect 3897 32823 3920 32857
rect 3840 32537 3920 32823
rect 3840 32503 3863 32537
rect 3897 32503 3920 32537
rect 3840 32480 3920 32503
rect 4000 32857 4080 32880
rect 4000 32823 4023 32857
rect 4057 32823 4080 32857
rect 4000 32537 4080 32823
rect 4000 32503 4023 32537
rect 4057 32503 4080 32537
rect 4000 32480 4080 32503
rect 4160 32857 4240 32880
rect 4160 32823 4183 32857
rect 4217 32823 4240 32857
rect 4160 32537 4240 32823
rect 4160 32503 4183 32537
rect 4217 32503 4240 32537
rect 4160 32480 4240 32503
rect 4320 32857 4400 32880
rect 4320 32823 4343 32857
rect 4377 32823 4400 32857
rect 4320 32537 4400 32823
rect 4320 32503 4343 32537
rect 4377 32503 4400 32537
rect 4320 32480 4400 32503
rect 4480 32857 4560 32880
rect 4480 32823 4503 32857
rect 4537 32823 4560 32857
rect 4480 32537 4560 32823
rect 4480 32503 4503 32537
rect 4537 32503 4560 32537
rect 4480 32480 4560 32503
rect 4640 32857 4720 32880
rect 4640 32823 4663 32857
rect 4697 32823 4720 32857
rect 4640 32537 4720 32823
rect 4640 32503 4663 32537
rect 4697 32503 4720 32537
rect 4640 32480 4720 32503
rect 4800 32857 4880 32880
rect 4800 32823 4823 32857
rect 4857 32823 4880 32857
rect 4800 32537 4880 32823
rect 4800 32503 4823 32537
rect 4857 32503 4880 32537
rect 4800 32480 4880 32503
rect 4960 32857 5040 32880
rect 4960 32823 4983 32857
rect 5017 32823 5040 32857
rect 4960 32537 5040 32823
rect 4960 32503 4983 32537
rect 5017 32503 5040 32537
rect 4960 32480 5040 32503
rect 5120 32857 5200 32880
rect 5120 32823 5143 32857
rect 5177 32823 5200 32857
rect 5120 32537 5200 32823
rect 5120 32503 5143 32537
rect 5177 32503 5200 32537
rect 5120 32480 5200 32503
rect 5280 32857 5360 32880
rect 5280 32823 5303 32857
rect 5337 32823 5360 32857
rect 5280 32537 5360 32823
rect 5280 32503 5303 32537
rect 5337 32503 5360 32537
rect 5280 32480 5360 32503
rect 5440 32857 5520 32880
rect 5440 32823 5463 32857
rect 5497 32823 5520 32857
rect 5440 32537 5520 32823
rect 5440 32503 5463 32537
rect 5497 32503 5520 32537
rect 5440 32480 5520 32503
rect 5600 32857 5680 32880
rect 5600 32823 5623 32857
rect 5657 32823 5680 32857
rect 5600 32537 5680 32823
rect 5600 32503 5623 32537
rect 5657 32503 5680 32537
rect 5600 32480 5680 32503
rect 5760 32857 5840 32880
rect 5760 32823 5783 32857
rect 5817 32823 5840 32857
rect 5760 32537 5840 32823
rect 5760 32503 5783 32537
rect 5817 32503 5840 32537
rect 5760 32480 5840 32503
rect 5920 32857 6000 32880
rect 5920 32823 5943 32857
rect 5977 32823 6000 32857
rect 5920 32537 6000 32823
rect 5920 32503 5943 32537
rect 5977 32503 6000 32537
rect 5920 32480 6000 32503
rect 6080 32857 6160 32880
rect 6080 32823 6103 32857
rect 6137 32823 6160 32857
rect 6080 32537 6160 32823
rect 6080 32503 6103 32537
rect 6137 32503 6160 32537
rect 6080 32480 6160 32503
rect 6240 32857 6320 32880
rect 6240 32823 6263 32857
rect 6297 32823 6320 32857
rect 6240 32537 6320 32823
rect 6240 32503 6263 32537
rect 6297 32503 6320 32537
rect 6240 32480 6320 32503
rect 6400 32857 6480 32880
rect 6400 32823 6423 32857
rect 6457 32823 6480 32857
rect 6400 32537 6480 32823
rect 6400 32503 6423 32537
rect 6457 32503 6480 32537
rect 6400 32480 6480 32503
rect 6560 32857 6640 32880
rect 6560 32823 6583 32857
rect 6617 32823 6640 32857
rect 6560 32537 6640 32823
rect 6560 32503 6583 32537
rect 6617 32503 6640 32537
rect 6560 32480 6640 32503
rect 6720 32857 6800 32880
rect 6720 32823 6743 32857
rect 6777 32823 6800 32857
rect 6720 32537 6800 32823
rect 6720 32503 6743 32537
rect 6777 32503 6800 32537
rect 6720 32480 6800 32503
rect 6880 32857 6960 32880
rect 6880 32823 6903 32857
rect 6937 32823 6960 32857
rect 6880 32537 6960 32823
rect 6880 32503 6903 32537
rect 6937 32503 6960 32537
rect 6880 32480 6960 32503
rect 7040 32857 7120 32880
rect 7040 32823 7063 32857
rect 7097 32823 7120 32857
rect 7040 32537 7120 32823
rect 7040 32503 7063 32537
rect 7097 32503 7120 32537
rect 7040 32480 7120 32503
rect 7200 32857 7280 32880
rect 7200 32823 7223 32857
rect 7257 32823 7280 32857
rect 7200 32537 7280 32823
rect 7200 32503 7223 32537
rect 7257 32503 7280 32537
rect 7200 32480 7280 32503
rect 7360 32857 7440 32880
rect 7360 32823 7383 32857
rect 7417 32823 7440 32857
rect 7360 32537 7440 32823
rect 7360 32503 7383 32537
rect 7417 32503 7440 32537
rect 7360 32480 7440 32503
rect 7520 32857 7600 32880
rect 7520 32823 7543 32857
rect 7577 32823 7600 32857
rect 7520 32537 7600 32823
rect 7520 32503 7543 32537
rect 7577 32503 7600 32537
rect 7520 32480 7600 32503
rect 7680 32857 7760 32880
rect 7680 32823 7703 32857
rect 7737 32823 7760 32857
rect 7680 32537 7760 32823
rect 7680 32503 7703 32537
rect 7737 32503 7760 32537
rect 7680 32480 7760 32503
rect 7840 32857 7920 32880
rect 7840 32823 7863 32857
rect 7897 32823 7920 32857
rect 7840 32537 7920 32823
rect 7840 32503 7863 32537
rect 7897 32503 7920 32537
rect 7840 32480 7920 32503
rect 8000 32857 8080 32880
rect 8000 32823 8023 32857
rect 8057 32823 8080 32857
rect 8000 32537 8080 32823
rect 8000 32503 8023 32537
rect 8057 32503 8080 32537
rect 8000 32480 8080 32503
rect 8160 32857 8240 32880
rect 8160 32823 8183 32857
rect 8217 32823 8240 32857
rect 8160 32537 8240 32823
rect 8160 32503 8183 32537
rect 8217 32503 8240 32537
rect 8160 32480 8240 32503
rect 8320 32857 8400 32880
rect 8320 32823 8343 32857
rect 8377 32823 8400 32857
rect 8320 32537 8400 32823
rect 8320 32503 8343 32537
rect 8377 32503 8400 32537
rect 8320 32480 8400 32503
rect 8480 32480 8560 32880
rect 8640 32480 8720 32880
rect 8800 32480 8880 32880
rect 8960 32480 9040 32880
rect 9120 32480 9200 32880
rect 9280 32480 9360 32880
rect 9440 32480 9520 32880
rect 9600 32480 9680 32880
rect 9760 32480 9840 32880
rect 9920 32480 10000 32880
rect 10080 32480 10160 32880
rect 10240 32480 10320 32880
rect 10400 32480 10480 32880
rect 10560 32480 10640 32880
rect 10720 32480 10800 32880
rect 10880 32480 10960 32880
rect 11040 32480 11120 32880
rect 11200 32480 11280 32880
rect 11360 32480 11440 32880
rect 11520 32480 11600 32880
rect 11680 32480 11760 32880
rect 11840 32480 11920 32880
rect 12000 32480 12080 32880
rect 12160 32480 12240 32880
rect 12320 32480 12400 32880
rect 12480 32857 12560 32880
rect 12480 32823 12503 32857
rect 12537 32823 12560 32857
rect 12480 32537 12560 32823
rect 12480 32503 12503 32537
rect 12537 32503 12560 32537
rect 12480 32480 12560 32503
rect 12640 32857 12720 32880
rect 12640 32823 12663 32857
rect 12697 32823 12720 32857
rect 12640 32537 12720 32823
rect 12640 32503 12663 32537
rect 12697 32503 12720 32537
rect 12640 32480 12720 32503
rect 12800 32857 12880 32880
rect 12800 32823 12823 32857
rect 12857 32823 12880 32857
rect 12800 32537 12880 32823
rect 12800 32503 12823 32537
rect 12857 32503 12880 32537
rect 12800 32480 12880 32503
rect 12960 32857 13040 32880
rect 12960 32823 12983 32857
rect 13017 32823 13040 32857
rect 12960 32537 13040 32823
rect 12960 32503 12983 32537
rect 13017 32503 13040 32537
rect 12960 32480 13040 32503
rect 13120 32857 13200 32880
rect 13120 32823 13143 32857
rect 13177 32823 13200 32857
rect 13120 32537 13200 32823
rect 13120 32503 13143 32537
rect 13177 32503 13200 32537
rect 13120 32480 13200 32503
rect 13280 32857 13360 32880
rect 13280 32823 13303 32857
rect 13337 32823 13360 32857
rect 13280 32537 13360 32823
rect 13280 32503 13303 32537
rect 13337 32503 13360 32537
rect 13280 32480 13360 32503
rect 13440 32857 13520 32880
rect 13440 32823 13463 32857
rect 13497 32823 13520 32857
rect 13440 32537 13520 32823
rect 13440 32503 13463 32537
rect 13497 32503 13520 32537
rect 13440 32480 13520 32503
rect 13600 32857 13680 32880
rect 13600 32823 13623 32857
rect 13657 32823 13680 32857
rect 13600 32537 13680 32823
rect 13600 32503 13623 32537
rect 13657 32503 13680 32537
rect 13600 32480 13680 32503
rect 13760 32857 13840 32880
rect 13760 32823 13783 32857
rect 13817 32823 13840 32857
rect 13760 32537 13840 32823
rect 13760 32503 13783 32537
rect 13817 32503 13840 32537
rect 13760 32480 13840 32503
rect 13920 32857 14000 32880
rect 13920 32823 13943 32857
rect 13977 32823 14000 32857
rect 13920 32537 14000 32823
rect 13920 32503 13943 32537
rect 13977 32503 14000 32537
rect 13920 32480 14000 32503
rect 14080 32857 14160 32880
rect 14080 32823 14103 32857
rect 14137 32823 14160 32857
rect 14080 32537 14160 32823
rect 14080 32503 14103 32537
rect 14137 32503 14160 32537
rect 14080 32480 14160 32503
rect 14240 32857 14320 32880
rect 14240 32823 14263 32857
rect 14297 32823 14320 32857
rect 14240 32537 14320 32823
rect 14240 32503 14263 32537
rect 14297 32503 14320 32537
rect 14240 32480 14320 32503
rect 14400 32857 14480 32880
rect 14400 32823 14423 32857
rect 14457 32823 14480 32857
rect 14400 32537 14480 32823
rect 14400 32503 14423 32537
rect 14457 32503 14480 32537
rect 14400 32480 14480 32503
rect 14560 32857 14640 32880
rect 14560 32823 14583 32857
rect 14617 32823 14640 32857
rect 14560 32537 14640 32823
rect 14560 32503 14583 32537
rect 14617 32503 14640 32537
rect 14560 32480 14640 32503
rect 14720 32857 14800 32880
rect 14720 32823 14743 32857
rect 14777 32823 14800 32857
rect 14720 32537 14800 32823
rect 14720 32503 14743 32537
rect 14777 32503 14800 32537
rect 14720 32480 14800 32503
rect 14880 32857 14960 32880
rect 14880 32823 14903 32857
rect 14937 32823 14960 32857
rect 14880 32537 14960 32823
rect 14880 32503 14903 32537
rect 14937 32503 14960 32537
rect 14880 32480 14960 32503
rect 15040 32857 15120 32880
rect 15040 32823 15063 32857
rect 15097 32823 15120 32857
rect 15040 32537 15120 32823
rect 15040 32503 15063 32537
rect 15097 32503 15120 32537
rect 15040 32480 15120 32503
rect 15200 32857 15280 32880
rect 15200 32823 15223 32857
rect 15257 32823 15280 32857
rect 15200 32537 15280 32823
rect 15200 32503 15223 32537
rect 15257 32503 15280 32537
rect 15200 32480 15280 32503
rect 15360 32857 15440 32880
rect 15360 32823 15383 32857
rect 15417 32823 15440 32857
rect 15360 32537 15440 32823
rect 15360 32503 15383 32537
rect 15417 32503 15440 32537
rect 15360 32480 15440 32503
rect 15520 32857 15600 32880
rect 15520 32823 15543 32857
rect 15577 32823 15600 32857
rect 15520 32537 15600 32823
rect 15520 32503 15543 32537
rect 15577 32503 15600 32537
rect 15520 32480 15600 32503
rect 15680 32857 15760 32880
rect 15680 32823 15703 32857
rect 15737 32823 15760 32857
rect 15680 32537 15760 32823
rect 15680 32503 15703 32537
rect 15737 32503 15760 32537
rect 15680 32480 15760 32503
rect 15840 32857 15920 32880
rect 15840 32823 15863 32857
rect 15897 32823 15920 32857
rect 15840 32537 15920 32823
rect 15840 32503 15863 32537
rect 15897 32503 15920 32537
rect 15840 32480 15920 32503
rect 16000 32857 16080 32880
rect 16000 32823 16023 32857
rect 16057 32823 16080 32857
rect 16000 32537 16080 32823
rect 16000 32503 16023 32537
rect 16057 32503 16080 32537
rect 16000 32480 16080 32503
rect 16160 32857 16240 32880
rect 16160 32823 16183 32857
rect 16217 32823 16240 32857
rect 16160 32537 16240 32823
rect 16160 32503 16183 32537
rect 16217 32503 16240 32537
rect 16160 32480 16240 32503
rect 16320 32857 16400 32880
rect 16320 32823 16343 32857
rect 16377 32823 16400 32857
rect 16320 32537 16400 32823
rect 16320 32503 16343 32537
rect 16377 32503 16400 32537
rect 16320 32480 16400 32503
rect 16480 32857 16560 32880
rect 16480 32823 16503 32857
rect 16537 32823 16560 32857
rect 16480 32537 16560 32823
rect 16480 32503 16503 32537
rect 16537 32503 16560 32537
rect 16480 32480 16560 32503
rect 16640 32857 16720 32880
rect 16640 32823 16663 32857
rect 16697 32823 16720 32857
rect 16640 32537 16720 32823
rect 16640 32503 16663 32537
rect 16697 32503 16720 32537
rect 16640 32480 16720 32503
rect 16800 32857 16880 32880
rect 16800 32823 16823 32857
rect 16857 32823 16880 32857
rect 16800 32537 16880 32823
rect 16800 32503 16823 32537
rect 16857 32503 16880 32537
rect 16800 32480 16880 32503
rect 16960 32857 17040 32880
rect 16960 32823 16983 32857
rect 17017 32823 17040 32857
rect 16960 32537 17040 32823
rect 16960 32503 16983 32537
rect 17017 32503 17040 32537
rect 16960 32480 17040 32503
rect 17120 32857 17200 32880
rect 17120 32823 17143 32857
rect 17177 32823 17200 32857
rect 17120 32537 17200 32823
rect 17120 32503 17143 32537
rect 17177 32503 17200 32537
rect 17120 32480 17200 32503
rect 17280 32857 17360 32880
rect 17280 32823 17303 32857
rect 17337 32823 17360 32857
rect 17280 32537 17360 32823
rect 17280 32503 17303 32537
rect 17337 32503 17360 32537
rect 17280 32480 17360 32503
rect 17440 32857 17520 32880
rect 17440 32823 17463 32857
rect 17497 32823 17520 32857
rect 17440 32537 17520 32823
rect 17440 32503 17463 32537
rect 17497 32503 17520 32537
rect 17440 32480 17520 32503
rect 17600 32857 17680 32880
rect 17600 32823 17623 32857
rect 17657 32823 17680 32857
rect 17600 32537 17680 32823
rect 17600 32503 17623 32537
rect 17657 32503 17680 32537
rect 17600 32480 17680 32503
rect 17760 32857 17840 32880
rect 17760 32823 17783 32857
rect 17817 32823 17840 32857
rect 17760 32537 17840 32823
rect 17760 32503 17783 32537
rect 17817 32503 17840 32537
rect 17760 32480 17840 32503
rect 17920 32857 18000 32880
rect 17920 32823 17943 32857
rect 17977 32823 18000 32857
rect 17920 32537 18000 32823
rect 17920 32503 17943 32537
rect 17977 32503 18000 32537
rect 17920 32480 18000 32503
rect 18080 32857 18160 32880
rect 18080 32823 18103 32857
rect 18137 32823 18160 32857
rect 18080 32537 18160 32823
rect 18080 32503 18103 32537
rect 18137 32503 18160 32537
rect 18080 32480 18160 32503
rect 18240 32857 18320 32880
rect 18240 32823 18263 32857
rect 18297 32823 18320 32857
rect 18240 32537 18320 32823
rect 18240 32503 18263 32537
rect 18297 32503 18320 32537
rect 18240 32480 18320 32503
rect 18400 32857 18480 32880
rect 18400 32823 18423 32857
rect 18457 32823 18480 32857
rect 18400 32537 18480 32823
rect 18400 32503 18423 32537
rect 18457 32503 18480 32537
rect 18400 32480 18480 32503
rect 18560 32857 18640 32880
rect 18560 32823 18583 32857
rect 18617 32823 18640 32857
rect 18560 32537 18640 32823
rect 18560 32503 18583 32537
rect 18617 32503 18640 32537
rect 18560 32480 18640 32503
rect 18720 32857 18800 32880
rect 18720 32823 18743 32857
rect 18777 32823 18800 32857
rect 18720 32537 18800 32823
rect 18720 32503 18743 32537
rect 18777 32503 18800 32537
rect 18720 32480 18800 32503
rect 18880 32857 18960 32880
rect 18880 32823 18903 32857
rect 18937 32823 18960 32857
rect 18880 32537 18960 32823
rect 18880 32503 18903 32537
rect 18937 32503 18960 32537
rect 18880 32480 18960 32503
rect 19040 32480 19120 32880
rect 19200 32480 19280 32880
rect 19360 32480 19440 32880
rect 19520 32480 19600 32880
rect 19680 32480 19760 32880
rect 19840 32480 19920 32880
rect 20000 32480 20080 32880
rect 20160 32480 20240 32880
rect 20320 32480 20400 32880
rect 20480 32480 20560 32880
rect 20640 32480 20720 32880
rect 20800 32480 20880 32880
rect 20960 32480 21040 32880
rect 21120 32480 21200 32880
rect 21280 32480 21360 32880
rect 21440 32480 21520 32880
rect 21600 32480 21680 32880
rect 21760 32480 21840 32880
rect 21920 32480 22000 32880
rect 22080 32480 22160 32880
rect 22240 32480 22320 32880
rect 22400 32480 22480 32880
rect 22560 32480 22640 32880
rect 22720 32480 22800 32880
rect 22880 32480 22960 32880
rect 23120 32857 23200 32880
rect 23120 32823 23143 32857
rect 23177 32823 23200 32857
rect 23120 32537 23200 32823
rect 23120 32503 23143 32537
rect 23177 32503 23200 32537
rect 23120 32480 23200 32503
rect 23280 32857 23360 32880
rect 23280 32823 23303 32857
rect 23337 32823 23360 32857
rect 23280 32537 23360 32823
rect 23280 32503 23303 32537
rect 23337 32503 23360 32537
rect 23280 32480 23360 32503
rect 23440 32857 23520 32880
rect 23440 32823 23463 32857
rect 23497 32823 23520 32857
rect 23440 32537 23520 32823
rect 23440 32503 23463 32537
rect 23497 32503 23520 32537
rect 23440 32480 23520 32503
rect 23600 32857 23680 32880
rect 23600 32823 23623 32857
rect 23657 32823 23680 32857
rect 23600 32537 23680 32823
rect 23600 32503 23623 32537
rect 23657 32503 23680 32537
rect 23600 32480 23680 32503
rect 23760 32857 23840 32880
rect 23760 32823 23783 32857
rect 23817 32823 23840 32857
rect 23760 32537 23840 32823
rect 23760 32503 23783 32537
rect 23817 32503 23840 32537
rect 23760 32480 23840 32503
rect 23920 32857 24000 32880
rect 23920 32823 23943 32857
rect 23977 32823 24000 32857
rect 23920 32537 24000 32823
rect 23920 32503 23943 32537
rect 23977 32503 24000 32537
rect 23920 32480 24000 32503
rect 24080 32857 24160 32880
rect 24080 32823 24103 32857
rect 24137 32823 24160 32857
rect 24080 32537 24160 32823
rect 24080 32503 24103 32537
rect 24137 32503 24160 32537
rect 24080 32480 24160 32503
rect 24240 32857 24320 32880
rect 24240 32823 24263 32857
rect 24297 32823 24320 32857
rect 24240 32537 24320 32823
rect 24240 32503 24263 32537
rect 24297 32503 24320 32537
rect 24240 32480 24320 32503
rect 24400 32857 24480 32880
rect 24400 32823 24423 32857
rect 24457 32823 24480 32857
rect 24400 32537 24480 32823
rect 24400 32503 24423 32537
rect 24457 32503 24480 32537
rect 24400 32480 24480 32503
rect 24560 32857 24640 32880
rect 24560 32823 24583 32857
rect 24617 32823 24640 32857
rect 24560 32537 24640 32823
rect 24560 32503 24583 32537
rect 24617 32503 24640 32537
rect 24560 32480 24640 32503
rect 24720 32857 24800 32880
rect 24720 32823 24743 32857
rect 24777 32823 24800 32857
rect 24720 32537 24800 32823
rect 24720 32503 24743 32537
rect 24777 32503 24800 32537
rect 24720 32480 24800 32503
rect 24880 32857 24960 32880
rect 24880 32823 24903 32857
rect 24937 32823 24960 32857
rect 24880 32537 24960 32823
rect 24880 32503 24903 32537
rect 24937 32503 24960 32537
rect 24880 32480 24960 32503
rect 25040 32857 25120 32880
rect 25040 32823 25063 32857
rect 25097 32823 25120 32857
rect 25040 32537 25120 32823
rect 25040 32503 25063 32537
rect 25097 32503 25120 32537
rect 25040 32480 25120 32503
rect 25200 32857 25280 32880
rect 25200 32823 25223 32857
rect 25257 32823 25280 32857
rect 25200 32537 25280 32823
rect 25200 32503 25223 32537
rect 25257 32503 25280 32537
rect 25200 32480 25280 32503
rect 25360 32857 25440 32880
rect 25360 32823 25383 32857
rect 25417 32823 25440 32857
rect 25360 32537 25440 32823
rect 25360 32503 25383 32537
rect 25417 32503 25440 32537
rect 25360 32480 25440 32503
rect 25520 32857 25600 32880
rect 25520 32823 25543 32857
rect 25577 32823 25600 32857
rect 25520 32537 25600 32823
rect 25520 32503 25543 32537
rect 25577 32503 25600 32537
rect 25520 32480 25600 32503
rect 25680 32857 25760 32880
rect 25680 32823 25703 32857
rect 25737 32823 25760 32857
rect 25680 32537 25760 32823
rect 25680 32503 25703 32537
rect 25737 32503 25760 32537
rect 25680 32480 25760 32503
rect 25840 32857 25920 32880
rect 25840 32823 25863 32857
rect 25897 32823 25920 32857
rect 25840 32537 25920 32823
rect 25840 32503 25863 32537
rect 25897 32503 25920 32537
rect 25840 32480 25920 32503
rect 26000 32857 26080 32880
rect 26000 32823 26023 32857
rect 26057 32823 26080 32857
rect 26000 32537 26080 32823
rect 26000 32503 26023 32537
rect 26057 32503 26080 32537
rect 26000 32480 26080 32503
rect 26160 32857 26240 32880
rect 26160 32823 26183 32857
rect 26217 32823 26240 32857
rect 26160 32537 26240 32823
rect 26160 32503 26183 32537
rect 26217 32503 26240 32537
rect 26160 32480 26240 32503
rect 26320 32857 26400 32880
rect 26320 32823 26343 32857
rect 26377 32823 26400 32857
rect 26320 32537 26400 32823
rect 26320 32503 26343 32537
rect 26377 32503 26400 32537
rect 26320 32480 26400 32503
rect 26480 32857 26560 32880
rect 26480 32823 26503 32857
rect 26537 32823 26560 32857
rect 26480 32537 26560 32823
rect 26480 32503 26503 32537
rect 26537 32503 26560 32537
rect 26480 32480 26560 32503
rect 26640 32857 26720 32880
rect 26640 32823 26663 32857
rect 26697 32823 26720 32857
rect 26640 32537 26720 32823
rect 26640 32503 26663 32537
rect 26697 32503 26720 32537
rect 26640 32480 26720 32503
rect 26800 32857 26880 32880
rect 26800 32823 26823 32857
rect 26857 32823 26880 32857
rect 26800 32537 26880 32823
rect 26800 32503 26823 32537
rect 26857 32503 26880 32537
rect 26800 32480 26880 32503
rect 26960 32857 27040 32880
rect 26960 32823 26983 32857
rect 27017 32823 27040 32857
rect 26960 32537 27040 32823
rect 26960 32503 26983 32537
rect 27017 32503 27040 32537
rect 26960 32480 27040 32503
rect 27120 32857 27200 32880
rect 27120 32823 27143 32857
rect 27177 32823 27200 32857
rect 27120 32537 27200 32823
rect 27120 32503 27143 32537
rect 27177 32503 27200 32537
rect 27120 32480 27200 32503
rect 27280 32857 27360 32880
rect 27280 32823 27303 32857
rect 27337 32823 27360 32857
rect 27280 32537 27360 32823
rect 27280 32503 27303 32537
rect 27337 32503 27360 32537
rect 27280 32480 27360 32503
rect 27440 32857 27520 32880
rect 27440 32823 27463 32857
rect 27497 32823 27520 32857
rect 27440 32537 27520 32823
rect 27440 32503 27463 32537
rect 27497 32503 27520 32537
rect 27440 32480 27520 32503
rect 27600 32857 27680 32880
rect 27600 32823 27623 32857
rect 27657 32823 27680 32857
rect 27600 32537 27680 32823
rect 27600 32503 27623 32537
rect 27657 32503 27680 32537
rect 27600 32480 27680 32503
rect 27760 32857 27840 32880
rect 27760 32823 27783 32857
rect 27817 32823 27840 32857
rect 27760 32537 27840 32823
rect 27760 32503 27783 32537
rect 27817 32503 27840 32537
rect 27760 32480 27840 32503
rect 27920 32857 28000 32880
rect 27920 32823 27943 32857
rect 27977 32823 28000 32857
rect 27920 32537 28000 32823
rect 27920 32503 27943 32537
rect 27977 32503 28000 32537
rect 27920 32480 28000 32503
rect 28080 32857 28160 32880
rect 28080 32823 28103 32857
rect 28137 32823 28160 32857
rect 28080 32537 28160 32823
rect 28080 32503 28103 32537
rect 28137 32503 28160 32537
rect 28080 32480 28160 32503
rect 28240 32857 28320 32880
rect 28240 32823 28263 32857
rect 28297 32823 28320 32857
rect 28240 32537 28320 32823
rect 28240 32503 28263 32537
rect 28297 32503 28320 32537
rect 28240 32480 28320 32503
rect 28400 32857 28480 32880
rect 28400 32823 28423 32857
rect 28457 32823 28480 32857
rect 28400 32537 28480 32823
rect 28400 32503 28423 32537
rect 28457 32503 28480 32537
rect 28400 32480 28480 32503
rect 28560 32857 28640 32880
rect 28560 32823 28583 32857
rect 28617 32823 28640 32857
rect 28560 32537 28640 32823
rect 28560 32503 28583 32537
rect 28617 32503 28640 32537
rect 28560 32480 28640 32503
rect 28720 32857 28800 32880
rect 28720 32823 28743 32857
rect 28777 32823 28800 32857
rect 28720 32537 28800 32823
rect 28720 32503 28743 32537
rect 28777 32503 28800 32537
rect 28720 32480 28800 32503
rect 28880 32857 28960 32880
rect 28880 32823 28903 32857
rect 28937 32823 28960 32857
rect 28880 32537 28960 32823
rect 28880 32503 28903 32537
rect 28937 32503 28960 32537
rect 28880 32480 28960 32503
rect 29040 32857 29120 32880
rect 29040 32823 29063 32857
rect 29097 32823 29120 32857
rect 29040 32537 29120 32823
rect 29040 32503 29063 32537
rect 29097 32503 29120 32537
rect 29040 32480 29120 32503
rect 29200 32857 29280 32880
rect 29200 32823 29223 32857
rect 29257 32823 29280 32857
rect 29200 32537 29280 32823
rect 29200 32503 29223 32537
rect 29257 32503 29280 32537
rect 29200 32480 29280 32503
rect 29360 32857 29440 32880
rect 29360 32823 29383 32857
rect 29417 32823 29440 32857
rect 29360 32537 29440 32823
rect 29360 32503 29383 32537
rect 29417 32503 29440 32537
rect 29360 32480 29440 32503
rect 29520 32480 29600 32880
rect 29680 32480 29760 32880
rect 29840 32480 29920 32880
rect 30000 32480 30080 32880
rect 30160 32480 30240 32880
rect 30320 32480 30400 32880
rect 30480 32480 30560 32880
rect 30640 32480 30720 32880
rect 30800 32480 30880 32880
rect 30960 32480 31040 32880
rect 31120 32480 31200 32880
rect 31280 32480 31360 32880
rect 31440 32480 31520 32880
rect 31600 32480 31680 32880
rect 31760 32480 31840 32880
rect 31920 32480 32000 32880
rect 32080 32480 32160 32880
rect 32240 32480 32320 32880
rect 32400 32480 32480 32880
rect 32560 32480 32640 32880
rect 32720 32480 32800 32880
rect 32880 32480 32960 32880
rect 33040 32480 33120 32880
rect 33200 32480 33280 32880
rect 33360 32480 33440 32880
rect 33520 32857 33600 32880
rect 33520 32823 33543 32857
rect 33577 32823 33600 32857
rect 33520 32537 33600 32823
rect 33520 32503 33543 32537
rect 33577 32503 33600 32537
rect 33520 32480 33600 32503
rect 33680 32857 33760 32880
rect 33680 32823 33703 32857
rect 33737 32823 33760 32857
rect 33680 32537 33760 32823
rect 33680 32503 33703 32537
rect 33737 32503 33760 32537
rect 33680 32480 33760 32503
rect 33840 32857 33920 32880
rect 33840 32823 33863 32857
rect 33897 32823 33920 32857
rect 33840 32537 33920 32823
rect 33840 32503 33863 32537
rect 33897 32503 33920 32537
rect 33840 32480 33920 32503
rect 34000 32857 34080 32880
rect 34000 32823 34023 32857
rect 34057 32823 34080 32857
rect 34000 32537 34080 32823
rect 34000 32503 34023 32537
rect 34057 32503 34080 32537
rect 34000 32480 34080 32503
rect 34160 32857 34240 32880
rect 34160 32823 34183 32857
rect 34217 32823 34240 32857
rect 34160 32537 34240 32823
rect 34160 32503 34183 32537
rect 34217 32503 34240 32537
rect 34160 32480 34240 32503
rect 34320 32857 34400 32880
rect 34320 32823 34343 32857
rect 34377 32823 34400 32857
rect 34320 32537 34400 32823
rect 34320 32503 34343 32537
rect 34377 32503 34400 32537
rect 34320 32480 34400 32503
rect 34480 32857 34560 32880
rect 34480 32823 34503 32857
rect 34537 32823 34560 32857
rect 34480 32537 34560 32823
rect 34480 32503 34503 32537
rect 34537 32503 34560 32537
rect 34480 32480 34560 32503
rect 34640 32857 34720 32880
rect 34640 32823 34663 32857
rect 34697 32823 34720 32857
rect 34640 32537 34720 32823
rect 34640 32503 34663 32537
rect 34697 32503 34720 32537
rect 34640 32480 34720 32503
rect 34800 32857 34880 32880
rect 34800 32823 34823 32857
rect 34857 32823 34880 32857
rect 34800 32537 34880 32823
rect 34800 32503 34823 32537
rect 34857 32503 34880 32537
rect 34800 32480 34880 32503
rect 34960 32857 35040 32880
rect 34960 32823 34983 32857
rect 35017 32823 35040 32857
rect 34960 32537 35040 32823
rect 34960 32503 34983 32537
rect 35017 32503 35040 32537
rect 34960 32480 35040 32503
rect 35120 32857 35200 32880
rect 35120 32823 35143 32857
rect 35177 32823 35200 32857
rect 35120 32537 35200 32823
rect 35120 32503 35143 32537
rect 35177 32503 35200 32537
rect 35120 32480 35200 32503
rect 35280 32857 35360 32880
rect 35280 32823 35303 32857
rect 35337 32823 35360 32857
rect 35280 32537 35360 32823
rect 35280 32503 35303 32537
rect 35337 32503 35360 32537
rect 35280 32480 35360 32503
rect 35440 32857 35520 32880
rect 35440 32823 35463 32857
rect 35497 32823 35520 32857
rect 35440 32537 35520 32823
rect 35440 32503 35463 32537
rect 35497 32503 35520 32537
rect 35440 32480 35520 32503
rect 35600 32857 35680 32880
rect 35600 32823 35623 32857
rect 35657 32823 35680 32857
rect 35600 32537 35680 32823
rect 35600 32503 35623 32537
rect 35657 32503 35680 32537
rect 35600 32480 35680 32503
rect 35760 32857 35840 32880
rect 35760 32823 35783 32857
rect 35817 32823 35840 32857
rect 35760 32537 35840 32823
rect 35760 32503 35783 32537
rect 35817 32503 35840 32537
rect 35760 32480 35840 32503
rect 35920 32857 36000 32880
rect 35920 32823 35943 32857
rect 35977 32823 36000 32857
rect 35920 32537 36000 32823
rect 35920 32503 35943 32537
rect 35977 32503 36000 32537
rect 35920 32480 36000 32503
rect 36080 32857 36160 32880
rect 36080 32823 36103 32857
rect 36137 32823 36160 32857
rect 36080 32537 36160 32823
rect 36080 32503 36103 32537
rect 36137 32503 36160 32537
rect 36080 32480 36160 32503
rect 36240 32857 36320 32880
rect 36240 32823 36263 32857
rect 36297 32823 36320 32857
rect 36240 32537 36320 32823
rect 36240 32503 36263 32537
rect 36297 32503 36320 32537
rect 36240 32480 36320 32503
rect 36400 32857 36480 32880
rect 36400 32823 36423 32857
rect 36457 32823 36480 32857
rect 36400 32537 36480 32823
rect 36400 32503 36423 32537
rect 36457 32503 36480 32537
rect 36400 32480 36480 32503
rect 36560 32857 36640 32880
rect 36560 32823 36583 32857
rect 36617 32823 36640 32857
rect 36560 32537 36640 32823
rect 36560 32503 36583 32537
rect 36617 32503 36640 32537
rect 36560 32480 36640 32503
rect 36720 32857 36800 32880
rect 36720 32823 36743 32857
rect 36777 32823 36800 32857
rect 36720 32537 36800 32823
rect 36720 32503 36743 32537
rect 36777 32503 36800 32537
rect 36720 32480 36800 32503
rect 36880 32857 36960 32880
rect 36880 32823 36903 32857
rect 36937 32823 36960 32857
rect 36880 32537 36960 32823
rect 36880 32503 36903 32537
rect 36937 32503 36960 32537
rect 36880 32480 36960 32503
rect 37040 32857 37120 32880
rect 37040 32823 37063 32857
rect 37097 32823 37120 32857
rect 37040 32537 37120 32823
rect 37040 32503 37063 32537
rect 37097 32503 37120 32537
rect 37040 32480 37120 32503
rect 37200 32857 37280 32880
rect 37200 32823 37223 32857
rect 37257 32823 37280 32857
rect 37200 32537 37280 32823
rect 37200 32503 37223 32537
rect 37257 32503 37280 32537
rect 37200 32480 37280 32503
rect 37360 32857 37440 32880
rect 37360 32823 37383 32857
rect 37417 32823 37440 32857
rect 37360 32537 37440 32823
rect 37360 32503 37383 32537
rect 37417 32503 37440 32537
rect 37360 32480 37440 32503
rect 37520 32857 37600 32880
rect 37520 32823 37543 32857
rect 37577 32823 37600 32857
rect 37520 32537 37600 32823
rect 37520 32503 37543 32537
rect 37577 32503 37600 32537
rect 37520 32480 37600 32503
rect 37680 32857 37760 32880
rect 37680 32823 37703 32857
rect 37737 32823 37760 32857
rect 37680 32537 37760 32823
rect 37680 32503 37703 32537
rect 37737 32503 37760 32537
rect 37680 32480 37760 32503
rect 37840 32857 37920 32880
rect 37840 32823 37863 32857
rect 37897 32823 37920 32857
rect 37840 32537 37920 32823
rect 37840 32503 37863 32537
rect 37897 32503 37920 32537
rect 37840 32480 37920 32503
rect 38000 32857 38080 32880
rect 38000 32823 38023 32857
rect 38057 32823 38080 32857
rect 38000 32537 38080 32823
rect 38000 32503 38023 32537
rect 38057 32503 38080 32537
rect 38000 32480 38080 32503
rect 38160 32857 38240 32880
rect 38160 32823 38183 32857
rect 38217 32823 38240 32857
rect 38160 32537 38240 32823
rect 38160 32503 38183 32537
rect 38217 32503 38240 32537
rect 38160 32480 38240 32503
rect 38320 32857 38400 32880
rect 38320 32823 38343 32857
rect 38377 32823 38400 32857
rect 38320 32537 38400 32823
rect 38320 32503 38343 32537
rect 38377 32503 38400 32537
rect 38320 32480 38400 32503
rect 38480 32857 38560 32880
rect 38480 32823 38503 32857
rect 38537 32823 38560 32857
rect 38480 32537 38560 32823
rect 38480 32503 38503 32537
rect 38537 32503 38560 32537
rect 38480 32480 38560 32503
rect 38640 32857 38720 32880
rect 38640 32823 38663 32857
rect 38697 32823 38720 32857
rect 38640 32537 38720 32823
rect 38640 32503 38663 32537
rect 38697 32503 38720 32537
rect 38640 32480 38720 32503
rect 38800 32857 38880 32880
rect 38800 32823 38823 32857
rect 38857 32823 38880 32857
rect 38800 32537 38880 32823
rect 38800 32503 38823 32537
rect 38857 32503 38880 32537
rect 38800 32480 38880 32503
rect 38960 32857 39040 32880
rect 38960 32823 38983 32857
rect 39017 32823 39040 32857
rect 38960 32537 39040 32823
rect 38960 32503 38983 32537
rect 39017 32503 39040 32537
rect 38960 32480 39040 32503
rect 39120 32857 39200 32880
rect 39120 32823 39143 32857
rect 39177 32823 39200 32857
rect 39120 32537 39200 32823
rect 39120 32503 39143 32537
rect 39177 32503 39200 32537
rect 39120 32480 39200 32503
rect 39280 32857 39360 32880
rect 39280 32823 39303 32857
rect 39337 32823 39360 32857
rect 39280 32537 39360 32823
rect 39280 32503 39303 32537
rect 39337 32503 39360 32537
rect 39280 32480 39360 32503
rect 39440 32857 39520 32880
rect 39440 32823 39463 32857
rect 39497 32823 39520 32857
rect 39440 32537 39520 32823
rect 39440 32503 39463 32537
rect 39497 32503 39520 32537
rect 39440 32480 39520 32503
rect 39600 32857 39680 32880
rect 39600 32823 39623 32857
rect 39657 32823 39680 32857
rect 39600 32537 39680 32823
rect 39600 32503 39623 32537
rect 39657 32503 39680 32537
rect 39600 32480 39680 32503
rect 39760 32857 39840 32880
rect 39760 32823 39783 32857
rect 39817 32823 39840 32857
rect 39760 32537 39840 32823
rect 39760 32503 39783 32537
rect 39817 32503 39840 32537
rect 39760 32480 39840 32503
rect 39920 32857 40000 32880
rect 39920 32823 39943 32857
rect 39977 32823 40000 32857
rect 39920 32537 40000 32823
rect 39920 32503 39943 32537
rect 39977 32503 40000 32537
rect 39920 32480 40000 32503
rect 40080 32857 40160 32880
rect 40080 32823 40103 32857
rect 40137 32823 40160 32857
rect 40080 32537 40160 32823
rect 40080 32503 40103 32537
rect 40137 32503 40160 32537
rect 40080 32480 40160 32503
rect 40240 32857 40320 32880
rect 40240 32823 40263 32857
rect 40297 32823 40320 32857
rect 40240 32537 40320 32823
rect 40240 32503 40263 32537
rect 40297 32503 40320 32537
rect 40240 32480 40320 32503
rect 40400 32857 40480 32880
rect 40400 32823 40423 32857
rect 40457 32823 40480 32857
rect 40400 32537 40480 32823
rect 40400 32503 40423 32537
rect 40457 32503 40480 32537
rect 40400 32480 40480 32503
rect 40560 32857 40640 32880
rect 40560 32823 40583 32857
rect 40617 32823 40640 32857
rect 40560 32537 40640 32823
rect 40560 32503 40583 32537
rect 40617 32503 40640 32537
rect 40560 32480 40640 32503
rect 40720 32857 40800 32880
rect 40720 32823 40743 32857
rect 40777 32823 40800 32857
rect 40720 32537 40800 32823
rect 40720 32503 40743 32537
rect 40777 32503 40800 32537
rect 40720 32480 40800 32503
rect 40880 32857 40960 32880
rect 40880 32823 40903 32857
rect 40937 32823 40960 32857
rect 40880 32537 40960 32823
rect 40880 32503 40903 32537
rect 40937 32503 40960 32537
rect 40880 32480 40960 32503
rect 41040 32857 41120 32880
rect 41040 32823 41063 32857
rect 41097 32823 41120 32857
rect 41040 32537 41120 32823
rect 41040 32503 41063 32537
rect 41097 32503 41120 32537
rect 41040 32480 41120 32503
rect 41200 32857 41280 32880
rect 41200 32823 41223 32857
rect 41257 32823 41280 32857
rect 41200 32537 41280 32823
rect 41200 32503 41223 32537
rect 41257 32503 41280 32537
rect 41200 32480 41280 32503
rect 41360 32857 41440 32880
rect 41360 32823 41383 32857
rect 41417 32823 41440 32857
rect 41360 32537 41440 32823
rect 41360 32503 41383 32537
rect 41417 32503 41440 32537
rect 41360 32480 41440 32503
rect 41520 32857 41600 32880
rect 41520 32823 41543 32857
rect 41577 32823 41600 32857
rect 41520 32537 41600 32823
rect 41520 32503 41543 32537
rect 41577 32503 41600 32537
rect 41520 32480 41600 32503
rect 41680 32857 41760 32880
rect 41680 32823 41703 32857
rect 41737 32823 41760 32857
rect 41680 32537 41760 32823
rect 41680 32503 41703 32537
rect 41737 32503 41760 32537
rect 41680 32480 41760 32503
rect 41840 32857 41920 32880
rect 41840 32823 41863 32857
rect 41897 32823 41920 32857
rect 41840 32537 41920 32823
rect 41840 32503 41863 32537
rect 41897 32503 41920 32537
rect 41840 32480 41920 32503
rect 0 32377 80 32400
rect 0 32343 23 32377
rect 57 32343 80 32377
rect 0 32057 80 32343
rect 0 32023 23 32057
rect 57 32023 80 32057
rect 0 31737 80 32023
rect 0 31703 23 31737
rect 57 31703 80 31737
rect 0 31417 80 31703
rect 0 31383 23 31417
rect 57 31383 80 31417
rect 0 31097 80 31383
rect 0 31063 23 31097
rect 57 31063 80 31097
rect 0 30777 80 31063
rect 0 30743 23 30777
rect 57 30743 80 30777
rect 0 30457 80 30743
rect 0 30423 23 30457
rect 57 30423 80 30457
rect 0 30400 80 30423
rect 160 32377 240 32400
rect 160 32343 183 32377
rect 217 32343 240 32377
rect 160 32057 240 32343
rect 160 32023 183 32057
rect 217 32023 240 32057
rect 160 31737 240 32023
rect 160 31703 183 31737
rect 217 31703 240 31737
rect 160 31417 240 31703
rect 160 31383 183 31417
rect 217 31383 240 31417
rect 160 31097 240 31383
rect 160 31063 183 31097
rect 217 31063 240 31097
rect 160 30777 240 31063
rect 160 30743 183 30777
rect 217 30743 240 30777
rect 160 30457 240 30743
rect 160 30423 183 30457
rect 217 30423 240 30457
rect 160 30400 240 30423
rect 320 32377 400 32400
rect 320 32343 343 32377
rect 377 32343 400 32377
rect 320 32057 400 32343
rect 320 32023 343 32057
rect 377 32023 400 32057
rect 320 31737 400 32023
rect 320 31703 343 31737
rect 377 31703 400 31737
rect 320 31417 400 31703
rect 320 31383 343 31417
rect 377 31383 400 31417
rect 320 31097 400 31383
rect 320 31063 343 31097
rect 377 31063 400 31097
rect 320 30777 400 31063
rect 320 30743 343 30777
rect 377 30743 400 30777
rect 320 30457 400 30743
rect 320 30423 343 30457
rect 377 30423 400 30457
rect 320 30400 400 30423
rect 480 32377 560 32400
rect 480 32343 503 32377
rect 537 32343 560 32377
rect 480 32057 560 32343
rect 480 32023 503 32057
rect 537 32023 560 32057
rect 480 31737 560 32023
rect 480 31703 503 31737
rect 537 31703 560 31737
rect 480 31417 560 31703
rect 480 31383 503 31417
rect 537 31383 560 31417
rect 480 31097 560 31383
rect 480 31063 503 31097
rect 537 31063 560 31097
rect 480 30777 560 31063
rect 480 30743 503 30777
rect 537 30743 560 30777
rect 480 30457 560 30743
rect 480 30423 503 30457
rect 537 30423 560 30457
rect 480 30400 560 30423
rect 640 32377 720 32400
rect 640 32343 663 32377
rect 697 32343 720 32377
rect 640 32057 720 32343
rect 640 32023 663 32057
rect 697 32023 720 32057
rect 640 31737 720 32023
rect 640 31703 663 31737
rect 697 31703 720 31737
rect 640 31417 720 31703
rect 640 31383 663 31417
rect 697 31383 720 31417
rect 640 31097 720 31383
rect 640 31063 663 31097
rect 697 31063 720 31097
rect 640 30777 720 31063
rect 640 30743 663 30777
rect 697 30743 720 30777
rect 640 30457 720 30743
rect 640 30423 663 30457
rect 697 30423 720 30457
rect 640 30400 720 30423
rect 800 32377 880 32400
rect 800 32343 823 32377
rect 857 32343 880 32377
rect 800 32057 880 32343
rect 800 32023 823 32057
rect 857 32023 880 32057
rect 800 31737 880 32023
rect 800 31703 823 31737
rect 857 31703 880 31737
rect 800 31417 880 31703
rect 800 31383 823 31417
rect 857 31383 880 31417
rect 800 31097 880 31383
rect 800 31063 823 31097
rect 857 31063 880 31097
rect 800 30777 880 31063
rect 800 30743 823 30777
rect 857 30743 880 30777
rect 800 30457 880 30743
rect 800 30423 823 30457
rect 857 30423 880 30457
rect 800 30400 880 30423
rect 960 32377 1040 32400
rect 960 32343 983 32377
rect 1017 32343 1040 32377
rect 960 32057 1040 32343
rect 960 32023 983 32057
rect 1017 32023 1040 32057
rect 960 31737 1040 32023
rect 960 31703 983 31737
rect 1017 31703 1040 31737
rect 960 31417 1040 31703
rect 960 31383 983 31417
rect 1017 31383 1040 31417
rect 960 31097 1040 31383
rect 960 31063 983 31097
rect 1017 31063 1040 31097
rect 960 30777 1040 31063
rect 960 30743 983 30777
rect 1017 30743 1040 30777
rect 960 30457 1040 30743
rect 960 30423 983 30457
rect 1017 30423 1040 30457
rect 960 30400 1040 30423
rect 1120 32377 1200 32400
rect 1120 32343 1143 32377
rect 1177 32343 1200 32377
rect 1120 32057 1200 32343
rect 1120 32023 1143 32057
rect 1177 32023 1200 32057
rect 1120 31737 1200 32023
rect 1120 31703 1143 31737
rect 1177 31703 1200 31737
rect 1120 31417 1200 31703
rect 1120 31383 1143 31417
rect 1177 31383 1200 31417
rect 1120 31097 1200 31383
rect 1120 31063 1143 31097
rect 1177 31063 1200 31097
rect 1120 30777 1200 31063
rect 1120 30743 1143 30777
rect 1177 30743 1200 30777
rect 1120 30457 1200 30743
rect 1120 30423 1143 30457
rect 1177 30423 1200 30457
rect 1120 30400 1200 30423
rect 1280 32377 1360 32400
rect 1280 32343 1303 32377
rect 1337 32343 1360 32377
rect 1280 32057 1360 32343
rect 1280 32023 1303 32057
rect 1337 32023 1360 32057
rect 1280 31737 1360 32023
rect 1280 31703 1303 31737
rect 1337 31703 1360 31737
rect 1280 31417 1360 31703
rect 1280 31383 1303 31417
rect 1337 31383 1360 31417
rect 1280 31097 1360 31383
rect 1280 31063 1303 31097
rect 1337 31063 1360 31097
rect 1280 30777 1360 31063
rect 1280 30743 1303 30777
rect 1337 30743 1360 30777
rect 1280 30457 1360 30743
rect 1280 30423 1303 30457
rect 1337 30423 1360 30457
rect 1280 30400 1360 30423
rect 1440 32377 1520 32400
rect 1440 32343 1463 32377
rect 1497 32343 1520 32377
rect 1440 32057 1520 32343
rect 1440 32023 1463 32057
rect 1497 32023 1520 32057
rect 1440 31737 1520 32023
rect 1440 31703 1463 31737
rect 1497 31703 1520 31737
rect 1440 31417 1520 31703
rect 1440 31383 1463 31417
rect 1497 31383 1520 31417
rect 1440 31097 1520 31383
rect 1440 31063 1463 31097
rect 1497 31063 1520 31097
rect 1440 30777 1520 31063
rect 1440 30743 1463 30777
rect 1497 30743 1520 30777
rect 1440 30457 1520 30743
rect 1440 30423 1463 30457
rect 1497 30423 1520 30457
rect 1440 30400 1520 30423
rect 1600 32377 1680 32400
rect 1600 32343 1623 32377
rect 1657 32343 1680 32377
rect 1600 32057 1680 32343
rect 1600 32023 1623 32057
rect 1657 32023 1680 32057
rect 1600 31737 1680 32023
rect 1600 31703 1623 31737
rect 1657 31703 1680 31737
rect 1600 31417 1680 31703
rect 1600 31383 1623 31417
rect 1657 31383 1680 31417
rect 1600 31097 1680 31383
rect 1600 31063 1623 31097
rect 1657 31063 1680 31097
rect 1600 30777 1680 31063
rect 1600 30743 1623 30777
rect 1657 30743 1680 30777
rect 1600 30457 1680 30743
rect 1600 30423 1623 30457
rect 1657 30423 1680 30457
rect 1600 30400 1680 30423
rect 1760 32377 1840 32400
rect 1760 32343 1783 32377
rect 1817 32343 1840 32377
rect 1760 32057 1840 32343
rect 1760 32023 1783 32057
rect 1817 32023 1840 32057
rect 1760 31737 1840 32023
rect 1760 31703 1783 31737
rect 1817 31703 1840 31737
rect 1760 31417 1840 31703
rect 1760 31383 1783 31417
rect 1817 31383 1840 31417
rect 1760 31097 1840 31383
rect 1760 31063 1783 31097
rect 1817 31063 1840 31097
rect 1760 30777 1840 31063
rect 1760 30743 1783 30777
rect 1817 30743 1840 30777
rect 1760 30457 1840 30743
rect 1760 30423 1783 30457
rect 1817 30423 1840 30457
rect 1760 30400 1840 30423
rect 1920 32377 2000 32400
rect 1920 32343 1943 32377
rect 1977 32343 2000 32377
rect 1920 32057 2000 32343
rect 1920 32023 1943 32057
rect 1977 32023 2000 32057
rect 1920 31737 2000 32023
rect 1920 31703 1943 31737
rect 1977 31703 2000 31737
rect 1920 31417 2000 31703
rect 1920 31383 1943 31417
rect 1977 31383 2000 31417
rect 1920 31097 2000 31383
rect 1920 31063 1943 31097
rect 1977 31063 2000 31097
rect 1920 30777 2000 31063
rect 1920 30743 1943 30777
rect 1977 30743 2000 30777
rect 1920 30457 2000 30743
rect 1920 30423 1943 30457
rect 1977 30423 2000 30457
rect 1920 30400 2000 30423
rect 2080 32377 2160 32400
rect 2080 32343 2103 32377
rect 2137 32343 2160 32377
rect 2080 32057 2160 32343
rect 2080 32023 2103 32057
rect 2137 32023 2160 32057
rect 2080 31737 2160 32023
rect 2080 31703 2103 31737
rect 2137 31703 2160 31737
rect 2080 31417 2160 31703
rect 2080 31383 2103 31417
rect 2137 31383 2160 31417
rect 2080 31097 2160 31383
rect 2080 31063 2103 31097
rect 2137 31063 2160 31097
rect 2080 30777 2160 31063
rect 2080 30743 2103 30777
rect 2137 30743 2160 30777
rect 2080 30457 2160 30743
rect 2080 30423 2103 30457
rect 2137 30423 2160 30457
rect 2080 30400 2160 30423
rect 2240 32377 2320 32400
rect 2240 32343 2263 32377
rect 2297 32343 2320 32377
rect 2240 32057 2320 32343
rect 2240 32023 2263 32057
rect 2297 32023 2320 32057
rect 2240 31737 2320 32023
rect 2240 31703 2263 31737
rect 2297 31703 2320 31737
rect 2240 31417 2320 31703
rect 2240 31383 2263 31417
rect 2297 31383 2320 31417
rect 2240 31097 2320 31383
rect 2240 31063 2263 31097
rect 2297 31063 2320 31097
rect 2240 30777 2320 31063
rect 2240 30743 2263 30777
rect 2297 30743 2320 30777
rect 2240 30457 2320 30743
rect 2240 30423 2263 30457
rect 2297 30423 2320 30457
rect 2240 30400 2320 30423
rect 2400 32377 2480 32400
rect 2400 32343 2423 32377
rect 2457 32343 2480 32377
rect 2400 32057 2480 32343
rect 2400 32023 2423 32057
rect 2457 32023 2480 32057
rect 2400 31737 2480 32023
rect 2400 31703 2423 31737
rect 2457 31703 2480 31737
rect 2400 31417 2480 31703
rect 2400 31383 2423 31417
rect 2457 31383 2480 31417
rect 2400 31097 2480 31383
rect 2400 31063 2423 31097
rect 2457 31063 2480 31097
rect 2400 30777 2480 31063
rect 2400 30743 2423 30777
rect 2457 30743 2480 30777
rect 2400 30457 2480 30743
rect 2400 30423 2423 30457
rect 2457 30423 2480 30457
rect 2400 30400 2480 30423
rect 2560 32377 2640 32400
rect 2560 32343 2583 32377
rect 2617 32343 2640 32377
rect 2560 32057 2640 32343
rect 2560 32023 2583 32057
rect 2617 32023 2640 32057
rect 2560 31737 2640 32023
rect 2560 31703 2583 31737
rect 2617 31703 2640 31737
rect 2560 31417 2640 31703
rect 2560 31383 2583 31417
rect 2617 31383 2640 31417
rect 2560 31097 2640 31383
rect 2560 31063 2583 31097
rect 2617 31063 2640 31097
rect 2560 30777 2640 31063
rect 2560 30743 2583 30777
rect 2617 30743 2640 30777
rect 2560 30457 2640 30743
rect 2560 30423 2583 30457
rect 2617 30423 2640 30457
rect 2560 30400 2640 30423
rect 2720 32377 2800 32400
rect 2720 32343 2743 32377
rect 2777 32343 2800 32377
rect 2720 32057 2800 32343
rect 2720 32023 2743 32057
rect 2777 32023 2800 32057
rect 2720 31737 2800 32023
rect 2720 31703 2743 31737
rect 2777 31703 2800 31737
rect 2720 31417 2800 31703
rect 2720 31383 2743 31417
rect 2777 31383 2800 31417
rect 2720 31097 2800 31383
rect 2720 31063 2743 31097
rect 2777 31063 2800 31097
rect 2720 30777 2800 31063
rect 2720 30743 2743 30777
rect 2777 30743 2800 30777
rect 2720 30457 2800 30743
rect 2720 30423 2743 30457
rect 2777 30423 2800 30457
rect 2720 30400 2800 30423
rect 2880 32377 2960 32400
rect 2880 32343 2903 32377
rect 2937 32343 2960 32377
rect 2880 32057 2960 32343
rect 2880 32023 2903 32057
rect 2937 32023 2960 32057
rect 2880 31737 2960 32023
rect 2880 31703 2903 31737
rect 2937 31703 2960 31737
rect 2880 31417 2960 31703
rect 2880 31383 2903 31417
rect 2937 31383 2960 31417
rect 2880 31097 2960 31383
rect 2880 31063 2903 31097
rect 2937 31063 2960 31097
rect 2880 30777 2960 31063
rect 2880 30743 2903 30777
rect 2937 30743 2960 30777
rect 2880 30457 2960 30743
rect 2880 30423 2903 30457
rect 2937 30423 2960 30457
rect 2880 30400 2960 30423
rect 3040 32377 3120 32400
rect 3040 32343 3063 32377
rect 3097 32343 3120 32377
rect 3040 32057 3120 32343
rect 3040 32023 3063 32057
rect 3097 32023 3120 32057
rect 3040 31737 3120 32023
rect 3040 31703 3063 31737
rect 3097 31703 3120 31737
rect 3040 31417 3120 31703
rect 3040 31383 3063 31417
rect 3097 31383 3120 31417
rect 3040 31097 3120 31383
rect 3040 31063 3063 31097
rect 3097 31063 3120 31097
rect 3040 30777 3120 31063
rect 3040 30743 3063 30777
rect 3097 30743 3120 30777
rect 3040 30457 3120 30743
rect 3040 30423 3063 30457
rect 3097 30423 3120 30457
rect 3040 30400 3120 30423
rect 3200 32377 3280 32400
rect 3200 32343 3223 32377
rect 3257 32343 3280 32377
rect 3200 32057 3280 32343
rect 3200 32023 3223 32057
rect 3257 32023 3280 32057
rect 3200 31737 3280 32023
rect 3200 31703 3223 31737
rect 3257 31703 3280 31737
rect 3200 31417 3280 31703
rect 3200 31383 3223 31417
rect 3257 31383 3280 31417
rect 3200 31097 3280 31383
rect 3200 31063 3223 31097
rect 3257 31063 3280 31097
rect 3200 30777 3280 31063
rect 3200 30743 3223 30777
rect 3257 30743 3280 30777
rect 3200 30457 3280 30743
rect 3200 30423 3223 30457
rect 3257 30423 3280 30457
rect 3200 30400 3280 30423
rect 3360 32377 3440 32400
rect 3360 32343 3383 32377
rect 3417 32343 3440 32377
rect 3360 32057 3440 32343
rect 3360 32023 3383 32057
rect 3417 32023 3440 32057
rect 3360 31737 3440 32023
rect 3360 31703 3383 31737
rect 3417 31703 3440 31737
rect 3360 31417 3440 31703
rect 3360 31383 3383 31417
rect 3417 31383 3440 31417
rect 3360 31097 3440 31383
rect 3360 31063 3383 31097
rect 3417 31063 3440 31097
rect 3360 30777 3440 31063
rect 3360 30743 3383 30777
rect 3417 30743 3440 30777
rect 3360 30457 3440 30743
rect 3360 30423 3383 30457
rect 3417 30423 3440 30457
rect 3360 30400 3440 30423
rect 3520 32377 3600 32400
rect 3520 32343 3543 32377
rect 3577 32343 3600 32377
rect 3520 32057 3600 32343
rect 3520 32023 3543 32057
rect 3577 32023 3600 32057
rect 3520 31737 3600 32023
rect 3520 31703 3543 31737
rect 3577 31703 3600 31737
rect 3520 31417 3600 31703
rect 3520 31383 3543 31417
rect 3577 31383 3600 31417
rect 3520 31097 3600 31383
rect 3520 31063 3543 31097
rect 3577 31063 3600 31097
rect 3520 30777 3600 31063
rect 3520 30743 3543 30777
rect 3577 30743 3600 30777
rect 3520 30457 3600 30743
rect 3520 30423 3543 30457
rect 3577 30423 3600 30457
rect 3520 30400 3600 30423
rect 3680 32377 3760 32400
rect 3680 32343 3703 32377
rect 3737 32343 3760 32377
rect 3680 32057 3760 32343
rect 3680 32023 3703 32057
rect 3737 32023 3760 32057
rect 3680 31737 3760 32023
rect 3680 31703 3703 31737
rect 3737 31703 3760 31737
rect 3680 31417 3760 31703
rect 3680 31383 3703 31417
rect 3737 31383 3760 31417
rect 3680 31097 3760 31383
rect 3680 31063 3703 31097
rect 3737 31063 3760 31097
rect 3680 30777 3760 31063
rect 3680 30743 3703 30777
rect 3737 30743 3760 30777
rect 3680 30457 3760 30743
rect 3680 30423 3703 30457
rect 3737 30423 3760 30457
rect 3680 30400 3760 30423
rect 3840 32377 3920 32400
rect 3840 32343 3863 32377
rect 3897 32343 3920 32377
rect 3840 32057 3920 32343
rect 3840 32023 3863 32057
rect 3897 32023 3920 32057
rect 3840 31737 3920 32023
rect 3840 31703 3863 31737
rect 3897 31703 3920 31737
rect 3840 31417 3920 31703
rect 3840 31383 3863 31417
rect 3897 31383 3920 31417
rect 3840 31097 3920 31383
rect 3840 31063 3863 31097
rect 3897 31063 3920 31097
rect 3840 30777 3920 31063
rect 3840 30743 3863 30777
rect 3897 30743 3920 30777
rect 3840 30457 3920 30743
rect 3840 30423 3863 30457
rect 3897 30423 3920 30457
rect 3840 30400 3920 30423
rect 4000 32377 4080 32400
rect 4000 32343 4023 32377
rect 4057 32343 4080 32377
rect 4000 32057 4080 32343
rect 4000 32023 4023 32057
rect 4057 32023 4080 32057
rect 4000 31737 4080 32023
rect 4000 31703 4023 31737
rect 4057 31703 4080 31737
rect 4000 31417 4080 31703
rect 4000 31383 4023 31417
rect 4057 31383 4080 31417
rect 4000 31097 4080 31383
rect 4000 31063 4023 31097
rect 4057 31063 4080 31097
rect 4000 30777 4080 31063
rect 4000 30743 4023 30777
rect 4057 30743 4080 30777
rect 4000 30457 4080 30743
rect 4000 30423 4023 30457
rect 4057 30423 4080 30457
rect 4000 30400 4080 30423
rect 4160 32377 4240 32400
rect 4160 32343 4183 32377
rect 4217 32343 4240 32377
rect 4160 32057 4240 32343
rect 4160 32023 4183 32057
rect 4217 32023 4240 32057
rect 4160 31737 4240 32023
rect 4160 31703 4183 31737
rect 4217 31703 4240 31737
rect 4160 31417 4240 31703
rect 4160 31383 4183 31417
rect 4217 31383 4240 31417
rect 4160 31097 4240 31383
rect 4160 31063 4183 31097
rect 4217 31063 4240 31097
rect 4160 30777 4240 31063
rect 4160 30743 4183 30777
rect 4217 30743 4240 30777
rect 4160 30457 4240 30743
rect 4160 30423 4183 30457
rect 4217 30423 4240 30457
rect 4160 30400 4240 30423
rect 4320 32377 4400 32400
rect 4320 32343 4343 32377
rect 4377 32343 4400 32377
rect 4320 32057 4400 32343
rect 4320 32023 4343 32057
rect 4377 32023 4400 32057
rect 4320 31737 4400 32023
rect 4320 31703 4343 31737
rect 4377 31703 4400 31737
rect 4320 31417 4400 31703
rect 4320 31383 4343 31417
rect 4377 31383 4400 31417
rect 4320 31097 4400 31383
rect 4320 31063 4343 31097
rect 4377 31063 4400 31097
rect 4320 30777 4400 31063
rect 4320 30743 4343 30777
rect 4377 30743 4400 30777
rect 4320 30457 4400 30743
rect 4320 30423 4343 30457
rect 4377 30423 4400 30457
rect 4320 30400 4400 30423
rect 4480 32377 4560 32400
rect 4480 32343 4503 32377
rect 4537 32343 4560 32377
rect 4480 32057 4560 32343
rect 4480 32023 4503 32057
rect 4537 32023 4560 32057
rect 4480 31737 4560 32023
rect 4480 31703 4503 31737
rect 4537 31703 4560 31737
rect 4480 31417 4560 31703
rect 4480 31383 4503 31417
rect 4537 31383 4560 31417
rect 4480 31097 4560 31383
rect 4480 31063 4503 31097
rect 4537 31063 4560 31097
rect 4480 30777 4560 31063
rect 4480 30743 4503 30777
rect 4537 30743 4560 30777
rect 4480 30457 4560 30743
rect 4480 30423 4503 30457
rect 4537 30423 4560 30457
rect 4480 30400 4560 30423
rect 4640 32377 4720 32400
rect 4640 32343 4663 32377
rect 4697 32343 4720 32377
rect 4640 32057 4720 32343
rect 4640 32023 4663 32057
rect 4697 32023 4720 32057
rect 4640 31737 4720 32023
rect 4640 31703 4663 31737
rect 4697 31703 4720 31737
rect 4640 31417 4720 31703
rect 4640 31383 4663 31417
rect 4697 31383 4720 31417
rect 4640 31097 4720 31383
rect 4640 31063 4663 31097
rect 4697 31063 4720 31097
rect 4640 30777 4720 31063
rect 4640 30743 4663 30777
rect 4697 30743 4720 30777
rect 4640 30457 4720 30743
rect 4640 30423 4663 30457
rect 4697 30423 4720 30457
rect 4640 30400 4720 30423
rect 4800 32377 4880 32400
rect 4800 32343 4823 32377
rect 4857 32343 4880 32377
rect 4800 32057 4880 32343
rect 4800 32023 4823 32057
rect 4857 32023 4880 32057
rect 4800 31737 4880 32023
rect 4800 31703 4823 31737
rect 4857 31703 4880 31737
rect 4800 31417 4880 31703
rect 4800 31383 4823 31417
rect 4857 31383 4880 31417
rect 4800 31097 4880 31383
rect 4800 31063 4823 31097
rect 4857 31063 4880 31097
rect 4800 30777 4880 31063
rect 4800 30743 4823 30777
rect 4857 30743 4880 30777
rect 4800 30457 4880 30743
rect 4800 30423 4823 30457
rect 4857 30423 4880 30457
rect 4800 30400 4880 30423
rect 4960 32377 5040 32400
rect 4960 32343 4983 32377
rect 5017 32343 5040 32377
rect 4960 32057 5040 32343
rect 4960 32023 4983 32057
rect 5017 32023 5040 32057
rect 4960 31737 5040 32023
rect 4960 31703 4983 31737
rect 5017 31703 5040 31737
rect 4960 31417 5040 31703
rect 4960 31383 4983 31417
rect 5017 31383 5040 31417
rect 4960 31097 5040 31383
rect 4960 31063 4983 31097
rect 5017 31063 5040 31097
rect 4960 30777 5040 31063
rect 4960 30743 4983 30777
rect 5017 30743 5040 30777
rect 4960 30457 5040 30743
rect 4960 30423 4983 30457
rect 5017 30423 5040 30457
rect 4960 30400 5040 30423
rect 5120 32377 5200 32400
rect 5120 32343 5143 32377
rect 5177 32343 5200 32377
rect 5120 32057 5200 32343
rect 5120 32023 5143 32057
rect 5177 32023 5200 32057
rect 5120 31737 5200 32023
rect 5120 31703 5143 31737
rect 5177 31703 5200 31737
rect 5120 31417 5200 31703
rect 5120 31383 5143 31417
rect 5177 31383 5200 31417
rect 5120 31097 5200 31383
rect 5120 31063 5143 31097
rect 5177 31063 5200 31097
rect 5120 30777 5200 31063
rect 5120 30743 5143 30777
rect 5177 30743 5200 30777
rect 5120 30457 5200 30743
rect 5120 30423 5143 30457
rect 5177 30423 5200 30457
rect 5120 30400 5200 30423
rect 5280 32377 5360 32400
rect 5280 32343 5303 32377
rect 5337 32343 5360 32377
rect 5280 32057 5360 32343
rect 5280 32023 5303 32057
rect 5337 32023 5360 32057
rect 5280 31737 5360 32023
rect 5280 31703 5303 31737
rect 5337 31703 5360 31737
rect 5280 31417 5360 31703
rect 5280 31383 5303 31417
rect 5337 31383 5360 31417
rect 5280 31097 5360 31383
rect 5280 31063 5303 31097
rect 5337 31063 5360 31097
rect 5280 30777 5360 31063
rect 5280 30743 5303 30777
rect 5337 30743 5360 30777
rect 5280 30457 5360 30743
rect 5280 30423 5303 30457
rect 5337 30423 5360 30457
rect 5280 30400 5360 30423
rect 5440 32377 5520 32400
rect 5440 32343 5463 32377
rect 5497 32343 5520 32377
rect 5440 32057 5520 32343
rect 5440 32023 5463 32057
rect 5497 32023 5520 32057
rect 5440 31737 5520 32023
rect 5440 31703 5463 31737
rect 5497 31703 5520 31737
rect 5440 31417 5520 31703
rect 5440 31383 5463 31417
rect 5497 31383 5520 31417
rect 5440 31097 5520 31383
rect 5440 31063 5463 31097
rect 5497 31063 5520 31097
rect 5440 30777 5520 31063
rect 5440 30743 5463 30777
rect 5497 30743 5520 30777
rect 5440 30457 5520 30743
rect 5440 30423 5463 30457
rect 5497 30423 5520 30457
rect 5440 30400 5520 30423
rect 5600 32377 5680 32400
rect 5600 32343 5623 32377
rect 5657 32343 5680 32377
rect 5600 32057 5680 32343
rect 5600 32023 5623 32057
rect 5657 32023 5680 32057
rect 5600 31737 5680 32023
rect 5600 31703 5623 31737
rect 5657 31703 5680 31737
rect 5600 31417 5680 31703
rect 5600 31383 5623 31417
rect 5657 31383 5680 31417
rect 5600 31097 5680 31383
rect 5600 31063 5623 31097
rect 5657 31063 5680 31097
rect 5600 30777 5680 31063
rect 5600 30743 5623 30777
rect 5657 30743 5680 30777
rect 5600 30457 5680 30743
rect 5600 30423 5623 30457
rect 5657 30423 5680 30457
rect 5600 30400 5680 30423
rect 5760 32377 5840 32400
rect 5760 32343 5783 32377
rect 5817 32343 5840 32377
rect 5760 32057 5840 32343
rect 5760 32023 5783 32057
rect 5817 32023 5840 32057
rect 5760 31737 5840 32023
rect 5760 31703 5783 31737
rect 5817 31703 5840 31737
rect 5760 31417 5840 31703
rect 5760 31383 5783 31417
rect 5817 31383 5840 31417
rect 5760 31097 5840 31383
rect 5760 31063 5783 31097
rect 5817 31063 5840 31097
rect 5760 30777 5840 31063
rect 5760 30743 5783 30777
rect 5817 30743 5840 30777
rect 5760 30457 5840 30743
rect 5760 30423 5783 30457
rect 5817 30423 5840 30457
rect 5760 30400 5840 30423
rect 5920 32377 6000 32400
rect 5920 32343 5943 32377
rect 5977 32343 6000 32377
rect 5920 32057 6000 32343
rect 5920 32023 5943 32057
rect 5977 32023 6000 32057
rect 5920 31737 6000 32023
rect 5920 31703 5943 31737
rect 5977 31703 6000 31737
rect 5920 31417 6000 31703
rect 5920 31383 5943 31417
rect 5977 31383 6000 31417
rect 5920 31097 6000 31383
rect 5920 31063 5943 31097
rect 5977 31063 6000 31097
rect 5920 30777 6000 31063
rect 5920 30743 5943 30777
rect 5977 30743 6000 30777
rect 5920 30457 6000 30743
rect 5920 30423 5943 30457
rect 5977 30423 6000 30457
rect 5920 30400 6000 30423
rect 6080 32377 6160 32400
rect 6080 32343 6103 32377
rect 6137 32343 6160 32377
rect 6080 32057 6160 32343
rect 6080 32023 6103 32057
rect 6137 32023 6160 32057
rect 6080 31737 6160 32023
rect 6080 31703 6103 31737
rect 6137 31703 6160 31737
rect 6080 31417 6160 31703
rect 6080 31383 6103 31417
rect 6137 31383 6160 31417
rect 6080 31097 6160 31383
rect 6080 31063 6103 31097
rect 6137 31063 6160 31097
rect 6080 30777 6160 31063
rect 6080 30743 6103 30777
rect 6137 30743 6160 30777
rect 6080 30457 6160 30743
rect 6080 30423 6103 30457
rect 6137 30423 6160 30457
rect 6080 30400 6160 30423
rect 6240 32377 6320 32400
rect 6240 32343 6263 32377
rect 6297 32343 6320 32377
rect 6240 32057 6320 32343
rect 6240 32023 6263 32057
rect 6297 32023 6320 32057
rect 6240 31737 6320 32023
rect 6240 31703 6263 31737
rect 6297 31703 6320 31737
rect 6240 31417 6320 31703
rect 6240 31383 6263 31417
rect 6297 31383 6320 31417
rect 6240 31097 6320 31383
rect 6240 31063 6263 31097
rect 6297 31063 6320 31097
rect 6240 30777 6320 31063
rect 6240 30743 6263 30777
rect 6297 30743 6320 30777
rect 6240 30457 6320 30743
rect 6240 30423 6263 30457
rect 6297 30423 6320 30457
rect 6240 30400 6320 30423
rect 6400 32377 6480 32400
rect 6400 32343 6423 32377
rect 6457 32343 6480 32377
rect 6400 32057 6480 32343
rect 6400 32023 6423 32057
rect 6457 32023 6480 32057
rect 6400 31737 6480 32023
rect 6400 31703 6423 31737
rect 6457 31703 6480 31737
rect 6400 31417 6480 31703
rect 6400 31383 6423 31417
rect 6457 31383 6480 31417
rect 6400 31097 6480 31383
rect 6400 31063 6423 31097
rect 6457 31063 6480 31097
rect 6400 30777 6480 31063
rect 6400 30743 6423 30777
rect 6457 30743 6480 30777
rect 6400 30457 6480 30743
rect 6400 30423 6423 30457
rect 6457 30423 6480 30457
rect 6400 30400 6480 30423
rect 6560 32377 6640 32400
rect 6560 32343 6583 32377
rect 6617 32343 6640 32377
rect 6560 32057 6640 32343
rect 6560 32023 6583 32057
rect 6617 32023 6640 32057
rect 6560 31737 6640 32023
rect 6560 31703 6583 31737
rect 6617 31703 6640 31737
rect 6560 31417 6640 31703
rect 6560 31383 6583 31417
rect 6617 31383 6640 31417
rect 6560 31097 6640 31383
rect 6560 31063 6583 31097
rect 6617 31063 6640 31097
rect 6560 30777 6640 31063
rect 6560 30743 6583 30777
rect 6617 30743 6640 30777
rect 6560 30457 6640 30743
rect 6560 30423 6583 30457
rect 6617 30423 6640 30457
rect 6560 30400 6640 30423
rect 6720 32377 6800 32400
rect 6720 32343 6743 32377
rect 6777 32343 6800 32377
rect 6720 32057 6800 32343
rect 6720 32023 6743 32057
rect 6777 32023 6800 32057
rect 6720 31737 6800 32023
rect 6720 31703 6743 31737
rect 6777 31703 6800 31737
rect 6720 31417 6800 31703
rect 6720 31383 6743 31417
rect 6777 31383 6800 31417
rect 6720 31097 6800 31383
rect 6720 31063 6743 31097
rect 6777 31063 6800 31097
rect 6720 30777 6800 31063
rect 6720 30743 6743 30777
rect 6777 30743 6800 30777
rect 6720 30457 6800 30743
rect 6720 30423 6743 30457
rect 6777 30423 6800 30457
rect 6720 30400 6800 30423
rect 6880 32377 6960 32400
rect 6880 32343 6903 32377
rect 6937 32343 6960 32377
rect 6880 32057 6960 32343
rect 6880 32023 6903 32057
rect 6937 32023 6960 32057
rect 6880 31737 6960 32023
rect 6880 31703 6903 31737
rect 6937 31703 6960 31737
rect 6880 31417 6960 31703
rect 6880 31383 6903 31417
rect 6937 31383 6960 31417
rect 6880 31097 6960 31383
rect 6880 31063 6903 31097
rect 6937 31063 6960 31097
rect 6880 30777 6960 31063
rect 6880 30743 6903 30777
rect 6937 30743 6960 30777
rect 6880 30457 6960 30743
rect 6880 30423 6903 30457
rect 6937 30423 6960 30457
rect 6880 30400 6960 30423
rect 7040 32377 7120 32400
rect 7040 32343 7063 32377
rect 7097 32343 7120 32377
rect 7040 32057 7120 32343
rect 7040 32023 7063 32057
rect 7097 32023 7120 32057
rect 7040 31737 7120 32023
rect 7040 31703 7063 31737
rect 7097 31703 7120 31737
rect 7040 31417 7120 31703
rect 7040 31383 7063 31417
rect 7097 31383 7120 31417
rect 7040 31097 7120 31383
rect 7040 31063 7063 31097
rect 7097 31063 7120 31097
rect 7040 30777 7120 31063
rect 7040 30743 7063 30777
rect 7097 30743 7120 30777
rect 7040 30457 7120 30743
rect 7040 30423 7063 30457
rect 7097 30423 7120 30457
rect 7040 30400 7120 30423
rect 7200 32377 7280 32400
rect 7200 32343 7223 32377
rect 7257 32343 7280 32377
rect 7200 32057 7280 32343
rect 7200 32023 7223 32057
rect 7257 32023 7280 32057
rect 7200 31737 7280 32023
rect 7200 31703 7223 31737
rect 7257 31703 7280 31737
rect 7200 31417 7280 31703
rect 7200 31383 7223 31417
rect 7257 31383 7280 31417
rect 7200 31097 7280 31383
rect 7200 31063 7223 31097
rect 7257 31063 7280 31097
rect 7200 30777 7280 31063
rect 7200 30743 7223 30777
rect 7257 30743 7280 30777
rect 7200 30457 7280 30743
rect 7200 30423 7223 30457
rect 7257 30423 7280 30457
rect 7200 30400 7280 30423
rect 7360 32377 7440 32400
rect 7360 32343 7383 32377
rect 7417 32343 7440 32377
rect 7360 32057 7440 32343
rect 7360 32023 7383 32057
rect 7417 32023 7440 32057
rect 7360 31737 7440 32023
rect 7360 31703 7383 31737
rect 7417 31703 7440 31737
rect 7360 31417 7440 31703
rect 7360 31383 7383 31417
rect 7417 31383 7440 31417
rect 7360 31097 7440 31383
rect 7360 31063 7383 31097
rect 7417 31063 7440 31097
rect 7360 30777 7440 31063
rect 7360 30743 7383 30777
rect 7417 30743 7440 30777
rect 7360 30457 7440 30743
rect 7360 30423 7383 30457
rect 7417 30423 7440 30457
rect 7360 30400 7440 30423
rect 7520 32377 7600 32400
rect 7520 32343 7543 32377
rect 7577 32343 7600 32377
rect 7520 32057 7600 32343
rect 7520 32023 7543 32057
rect 7577 32023 7600 32057
rect 7520 31737 7600 32023
rect 7520 31703 7543 31737
rect 7577 31703 7600 31737
rect 7520 31417 7600 31703
rect 7520 31383 7543 31417
rect 7577 31383 7600 31417
rect 7520 31097 7600 31383
rect 7520 31063 7543 31097
rect 7577 31063 7600 31097
rect 7520 30777 7600 31063
rect 7520 30743 7543 30777
rect 7577 30743 7600 30777
rect 7520 30457 7600 30743
rect 7520 30423 7543 30457
rect 7577 30423 7600 30457
rect 7520 30400 7600 30423
rect 7680 32377 7760 32400
rect 7680 32343 7703 32377
rect 7737 32343 7760 32377
rect 7680 32057 7760 32343
rect 7680 32023 7703 32057
rect 7737 32023 7760 32057
rect 7680 31737 7760 32023
rect 7680 31703 7703 31737
rect 7737 31703 7760 31737
rect 7680 31417 7760 31703
rect 7680 31383 7703 31417
rect 7737 31383 7760 31417
rect 7680 31097 7760 31383
rect 7680 31063 7703 31097
rect 7737 31063 7760 31097
rect 7680 30777 7760 31063
rect 7680 30743 7703 30777
rect 7737 30743 7760 30777
rect 7680 30457 7760 30743
rect 7680 30423 7703 30457
rect 7737 30423 7760 30457
rect 7680 30400 7760 30423
rect 7840 32377 7920 32400
rect 7840 32343 7863 32377
rect 7897 32343 7920 32377
rect 7840 32057 7920 32343
rect 7840 32023 7863 32057
rect 7897 32023 7920 32057
rect 7840 31737 7920 32023
rect 7840 31703 7863 31737
rect 7897 31703 7920 31737
rect 7840 31417 7920 31703
rect 7840 31383 7863 31417
rect 7897 31383 7920 31417
rect 7840 31097 7920 31383
rect 7840 31063 7863 31097
rect 7897 31063 7920 31097
rect 7840 30777 7920 31063
rect 7840 30743 7863 30777
rect 7897 30743 7920 30777
rect 7840 30457 7920 30743
rect 7840 30423 7863 30457
rect 7897 30423 7920 30457
rect 7840 30400 7920 30423
rect 8000 32377 8080 32400
rect 8000 32343 8023 32377
rect 8057 32343 8080 32377
rect 8000 32057 8080 32343
rect 8000 32023 8023 32057
rect 8057 32023 8080 32057
rect 8000 31737 8080 32023
rect 8000 31703 8023 31737
rect 8057 31703 8080 31737
rect 8000 31417 8080 31703
rect 8000 31383 8023 31417
rect 8057 31383 8080 31417
rect 8000 31097 8080 31383
rect 8000 31063 8023 31097
rect 8057 31063 8080 31097
rect 8000 30777 8080 31063
rect 8000 30743 8023 30777
rect 8057 30743 8080 30777
rect 8000 30457 8080 30743
rect 8000 30423 8023 30457
rect 8057 30423 8080 30457
rect 8000 30400 8080 30423
rect 8160 32377 8240 32400
rect 8160 32343 8183 32377
rect 8217 32343 8240 32377
rect 8160 32057 8240 32343
rect 8160 32023 8183 32057
rect 8217 32023 8240 32057
rect 8160 31737 8240 32023
rect 8160 31703 8183 31737
rect 8217 31703 8240 31737
rect 8160 31417 8240 31703
rect 8160 31383 8183 31417
rect 8217 31383 8240 31417
rect 8160 31097 8240 31383
rect 8160 31063 8183 31097
rect 8217 31063 8240 31097
rect 8160 30777 8240 31063
rect 8160 30743 8183 30777
rect 8217 30743 8240 30777
rect 8160 30457 8240 30743
rect 8160 30423 8183 30457
rect 8217 30423 8240 30457
rect 8160 30400 8240 30423
rect 8320 32377 8400 32400
rect 8320 32343 8343 32377
rect 8377 32343 8400 32377
rect 8320 32057 8400 32343
rect 8320 32023 8343 32057
rect 8377 32023 8400 32057
rect 8320 31737 8400 32023
rect 8320 31703 8343 31737
rect 8377 31703 8400 31737
rect 8320 31417 8400 31703
rect 8320 31383 8343 31417
rect 8377 31383 8400 31417
rect 8320 31097 8400 31383
rect 8320 31063 8343 31097
rect 8377 31063 8400 31097
rect 8320 30777 8400 31063
rect 8320 30743 8343 30777
rect 8377 30743 8400 30777
rect 8320 30457 8400 30743
rect 8320 30423 8343 30457
rect 8377 30423 8400 30457
rect 8320 30400 8400 30423
rect 8480 30400 8560 32400
rect 8640 30400 8720 32400
rect 8800 30400 8880 32400
rect 8960 30400 9040 32400
rect 9120 30400 9200 32400
rect 9280 30400 9360 32400
rect 9440 30400 9520 32400
rect 9600 30400 9680 32400
rect 9760 30400 9840 32400
rect 9920 30400 10000 32400
rect 10080 30400 10160 32400
rect 10240 30400 10320 32400
rect 10400 30400 10480 32400
rect 10560 30400 10640 32400
rect 10720 30400 10800 32400
rect 10880 30400 10960 32400
rect 11040 30400 11120 32400
rect 11200 30400 11280 32400
rect 11360 30400 11440 32400
rect 11520 30400 11600 32400
rect 11680 30400 11760 32400
rect 11840 30400 11920 32400
rect 12000 30400 12080 32400
rect 12160 30400 12240 32400
rect 12320 30400 12400 32400
rect 12480 32377 12560 32400
rect 12480 32343 12503 32377
rect 12537 32343 12560 32377
rect 12480 32057 12560 32343
rect 12480 32023 12503 32057
rect 12537 32023 12560 32057
rect 12480 31737 12560 32023
rect 12480 31703 12503 31737
rect 12537 31703 12560 31737
rect 12480 31417 12560 31703
rect 12480 31383 12503 31417
rect 12537 31383 12560 31417
rect 12480 31097 12560 31383
rect 12480 31063 12503 31097
rect 12537 31063 12560 31097
rect 12480 30777 12560 31063
rect 12480 30743 12503 30777
rect 12537 30743 12560 30777
rect 12480 30457 12560 30743
rect 12480 30423 12503 30457
rect 12537 30423 12560 30457
rect 12480 30400 12560 30423
rect 12640 32377 12720 32400
rect 12640 32343 12663 32377
rect 12697 32343 12720 32377
rect 12640 32057 12720 32343
rect 12640 32023 12663 32057
rect 12697 32023 12720 32057
rect 12640 31737 12720 32023
rect 12640 31703 12663 31737
rect 12697 31703 12720 31737
rect 12640 31417 12720 31703
rect 12640 31383 12663 31417
rect 12697 31383 12720 31417
rect 12640 31097 12720 31383
rect 12640 31063 12663 31097
rect 12697 31063 12720 31097
rect 12640 30777 12720 31063
rect 12640 30743 12663 30777
rect 12697 30743 12720 30777
rect 12640 30457 12720 30743
rect 12640 30423 12663 30457
rect 12697 30423 12720 30457
rect 12640 30400 12720 30423
rect 12800 32377 12880 32400
rect 12800 32343 12823 32377
rect 12857 32343 12880 32377
rect 12800 32057 12880 32343
rect 12800 32023 12823 32057
rect 12857 32023 12880 32057
rect 12800 31737 12880 32023
rect 12800 31703 12823 31737
rect 12857 31703 12880 31737
rect 12800 31417 12880 31703
rect 12800 31383 12823 31417
rect 12857 31383 12880 31417
rect 12800 31097 12880 31383
rect 12800 31063 12823 31097
rect 12857 31063 12880 31097
rect 12800 30777 12880 31063
rect 12800 30743 12823 30777
rect 12857 30743 12880 30777
rect 12800 30457 12880 30743
rect 12800 30423 12823 30457
rect 12857 30423 12880 30457
rect 12800 30400 12880 30423
rect 12960 32377 13040 32400
rect 12960 32343 12983 32377
rect 13017 32343 13040 32377
rect 12960 32057 13040 32343
rect 12960 32023 12983 32057
rect 13017 32023 13040 32057
rect 12960 31737 13040 32023
rect 12960 31703 12983 31737
rect 13017 31703 13040 31737
rect 12960 31417 13040 31703
rect 12960 31383 12983 31417
rect 13017 31383 13040 31417
rect 12960 31097 13040 31383
rect 12960 31063 12983 31097
rect 13017 31063 13040 31097
rect 12960 30777 13040 31063
rect 12960 30743 12983 30777
rect 13017 30743 13040 30777
rect 12960 30457 13040 30743
rect 12960 30423 12983 30457
rect 13017 30423 13040 30457
rect 12960 30400 13040 30423
rect 13120 32377 13200 32400
rect 13120 32343 13143 32377
rect 13177 32343 13200 32377
rect 13120 32057 13200 32343
rect 13120 32023 13143 32057
rect 13177 32023 13200 32057
rect 13120 31737 13200 32023
rect 13120 31703 13143 31737
rect 13177 31703 13200 31737
rect 13120 31417 13200 31703
rect 13120 31383 13143 31417
rect 13177 31383 13200 31417
rect 13120 31097 13200 31383
rect 13120 31063 13143 31097
rect 13177 31063 13200 31097
rect 13120 30777 13200 31063
rect 13120 30743 13143 30777
rect 13177 30743 13200 30777
rect 13120 30457 13200 30743
rect 13120 30423 13143 30457
rect 13177 30423 13200 30457
rect 13120 30400 13200 30423
rect 13280 32377 13360 32400
rect 13280 32343 13303 32377
rect 13337 32343 13360 32377
rect 13280 32057 13360 32343
rect 13280 32023 13303 32057
rect 13337 32023 13360 32057
rect 13280 31737 13360 32023
rect 13280 31703 13303 31737
rect 13337 31703 13360 31737
rect 13280 31417 13360 31703
rect 13280 31383 13303 31417
rect 13337 31383 13360 31417
rect 13280 31097 13360 31383
rect 13280 31063 13303 31097
rect 13337 31063 13360 31097
rect 13280 30777 13360 31063
rect 13280 30743 13303 30777
rect 13337 30743 13360 30777
rect 13280 30457 13360 30743
rect 13280 30423 13303 30457
rect 13337 30423 13360 30457
rect 13280 30400 13360 30423
rect 13440 32377 13520 32400
rect 13440 32343 13463 32377
rect 13497 32343 13520 32377
rect 13440 32057 13520 32343
rect 13440 32023 13463 32057
rect 13497 32023 13520 32057
rect 13440 31737 13520 32023
rect 13440 31703 13463 31737
rect 13497 31703 13520 31737
rect 13440 31417 13520 31703
rect 13440 31383 13463 31417
rect 13497 31383 13520 31417
rect 13440 31097 13520 31383
rect 13440 31063 13463 31097
rect 13497 31063 13520 31097
rect 13440 30777 13520 31063
rect 13440 30743 13463 30777
rect 13497 30743 13520 30777
rect 13440 30457 13520 30743
rect 13440 30423 13463 30457
rect 13497 30423 13520 30457
rect 13440 30400 13520 30423
rect 13600 32377 13680 32400
rect 13600 32343 13623 32377
rect 13657 32343 13680 32377
rect 13600 32057 13680 32343
rect 13600 32023 13623 32057
rect 13657 32023 13680 32057
rect 13600 31737 13680 32023
rect 13600 31703 13623 31737
rect 13657 31703 13680 31737
rect 13600 31417 13680 31703
rect 13600 31383 13623 31417
rect 13657 31383 13680 31417
rect 13600 31097 13680 31383
rect 13600 31063 13623 31097
rect 13657 31063 13680 31097
rect 13600 30777 13680 31063
rect 13600 30743 13623 30777
rect 13657 30743 13680 30777
rect 13600 30457 13680 30743
rect 13600 30423 13623 30457
rect 13657 30423 13680 30457
rect 13600 30400 13680 30423
rect 13760 32377 13840 32400
rect 13760 32343 13783 32377
rect 13817 32343 13840 32377
rect 13760 32057 13840 32343
rect 13760 32023 13783 32057
rect 13817 32023 13840 32057
rect 13760 31737 13840 32023
rect 13760 31703 13783 31737
rect 13817 31703 13840 31737
rect 13760 31417 13840 31703
rect 13760 31383 13783 31417
rect 13817 31383 13840 31417
rect 13760 31097 13840 31383
rect 13760 31063 13783 31097
rect 13817 31063 13840 31097
rect 13760 30777 13840 31063
rect 13760 30743 13783 30777
rect 13817 30743 13840 30777
rect 13760 30457 13840 30743
rect 13760 30423 13783 30457
rect 13817 30423 13840 30457
rect 13760 30400 13840 30423
rect 13920 32377 14000 32400
rect 13920 32343 13943 32377
rect 13977 32343 14000 32377
rect 13920 32057 14000 32343
rect 13920 32023 13943 32057
rect 13977 32023 14000 32057
rect 13920 31737 14000 32023
rect 13920 31703 13943 31737
rect 13977 31703 14000 31737
rect 13920 31417 14000 31703
rect 13920 31383 13943 31417
rect 13977 31383 14000 31417
rect 13920 31097 14000 31383
rect 13920 31063 13943 31097
rect 13977 31063 14000 31097
rect 13920 30777 14000 31063
rect 13920 30743 13943 30777
rect 13977 30743 14000 30777
rect 13920 30457 14000 30743
rect 13920 30423 13943 30457
rect 13977 30423 14000 30457
rect 13920 30400 14000 30423
rect 14080 32377 14160 32400
rect 14080 32343 14103 32377
rect 14137 32343 14160 32377
rect 14080 32057 14160 32343
rect 14080 32023 14103 32057
rect 14137 32023 14160 32057
rect 14080 31737 14160 32023
rect 14080 31703 14103 31737
rect 14137 31703 14160 31737
rect 14080 31417 14160 31703
rect 14080 31383 14103 31417
rect 14137 31383 14160 31417
rect 14080 31097 14160 31383
rect 14080 31063 14103 31097
rect 14137 31063 14160 31097
rect 14080 30777 14160 31063
rect 14080 30743 14103 30777
rect 14137 30743 14160 30777
rect 14080 30457 14160 30743
rect 14080 30423 14103 30457
rect 14137 30423 14160 30457
rect 14080 30400 14160 30423
rect 14240 32377 14320 32400
rect 14240 32343 14263 32377
rect 14297 32343 14320 32377
rect 14240 32057 14320 32343
rect 14240 32023 14263 32057
rect 14297 32023 14320 32057
rect 14240 31737 14320 32023
rect 14240 31703 14263 31737
rect 14297 31703 14320 31737
rect 14240 31417 14320 31703
rect 14240 31383 14263 31417
rect 14297 31383 14320 31417
rect 14240 31097 14320 31383
rect 14240 31063 14263 31097
rect 14297 31063 14320 31097
rect 14240 30777 14320 31063
rect 14240 30743 14263 30777
rect 14297 30743 14320 30777
rect 14240 30457 14320 30743
rect 14240 30423 14263 30457
rect 14297 30423 14320 30457
rect 14240 30400 14320 30423
rect 14400 32377 14480 32400
rect 14400 32343 14423 32377
rect 14457 32343 14480 32377
rect 14400 32057 14480 32343
rect 14400 32023 14423 32057
rect 14457 32023 14480 32057
rect 14400 31737 14480 32023
rect 14400 31703 14423 31737
rect 14457 31703 14480 31737
rect 14400 31417 14480 31703
rect 14400 31383 14423 31417
rect 14457 31383 14480 31417
rect 14400 31097 14480 31383
rect 14400 31063 14423 31097
rect 14457 31063 14480 31097
rect 14400 30777 14480 31063
rect 14400 30743 14423 30777
rect 14457 30743 14480 30777
rect 14400 30457 14480 30743
rect 14400 30423 14423 30457
rect 14457 30423 14480 30457
rect 14400 30400 14480 30423
rect 14560 32377 14640 32400
rect 14560 32343 14583 32377
rect 14617 32343 14640 32377
rect 14560 32057 14640 32343
rect 14560 32023 14583 32057
rect 14617 32023 14640 32057
rect 14560 31737 14640 32023
rect 14560 31703 14583 31737
rect 14617 31703 14640 31737
rect 14560 31417 14640 31703
rect 14560 31383 14583 31417
rect 14617 31383 14640 31417
rect 14560 31097 14640 31383
rect 14560 31063 14583 31097
rect 14617 31063 14640 31097
rect 14560 30777 14640 31063
rect 14560 30743 14583 30777
rect 14617 30743 14640 30777
rect 14560 30457 14640 30743
rect 14560 30423 14583 30457
rect 14617 30423 14640 30457
rect 14560 30400 14640 30423
rect 14720 32377 14800 32400
rect 14720 32343 14743 32377
rect 14777 32343 14800 32377
rect 14720 32057 14800 32343
rect 14720 32023 14743 32057
rect 14777 32023 14800 32057
rect 14720 31737 14800 32023
rect 14720 31703 14743 31737
rect 14777 31703 14800 31737
rect 14720 31417 14800 31703
rect 14720 31383 14743 31417
rect 14777 31383 14800 31417
rect 14720 31097 14800 31383
rect 14720 31063 14743 31097
rect 14777 31063 14800 31097
rect 14720 30777 14800 31063
rect 14720 30743 14743 30777
rect 14777 30743 14800 30777
rect 14720 30457 14800 30743
rect 14720 30423 14743 30457
rect 14777 30423 14800 30457
rect 14720 30400 14800 30423
rect 14880 32377 14960 32400
rect 14880 32343 14903 32377
rect 14937 32343 14960 32377
rect 14880 32057 14960 32343
rect 14880 32023 14903 32057
rect 14937 32023 14960 32057
rect 14880 31737 14960 32023
rect 14880 31703 14903 31737
rect 14937 31703 14960 31737
rect 14880 31417 14960 31703
rect 14880 31383 14903 31417
rect 14937 31383 14960 31417
rect 14880 31097 14960 31383
rect 14880 31063 14903 31097
rect 14937 31063 14960 31097
rect 14880 30777 14960 31063
rect 14880 30743 14903 30777
rect 14937 30743 14960 30777
rect 14880 30457 14960 30743
rect 14880 30423 14903 30457
rect 14937 30423 14960 30457
rect 14880 30400 14960 30423
rect 15040 32377 15120 32400
rect 15040 32343 15063 32377
rect 15097 32343 15120 32377
rect 15040 32057 15120 32343
rect 15040 32023 15063 32057
rect 15097 32023 15120 32057
rect 15040 31737 15120 32023
rect 15040 31703 15063 31737
rect 15097 31703 15120 31737
rect 15040 31417 15120 31703
rect 15040 31383 15063 31417
rect 15097 31383 15120 31417
rect 15040 31097 15120 31383
rect 15040 31063 15063 31097
rect 15097 31063 15120 31097
rect 15040 30777 15120 31063
rect 15040 30743 15063 30777
rect 15097 30743 15120 30777
rect 15040 30457 15120 30743
rect 15040 30423 15063 30457
rect 15097 30423 15120 30457
rect 15040 30400 15120 30423
rect 15200 32377 15280 32400
rect 15200 32343 15223 32377
rect 15257 32343 15280 32377
rect 15200 32057 15280 32343
rect 15200 32023 15223 32057
rect 15257 32023 15280 32057
rect 15200 31737 15280 32023
rect 15200 31703 15223 31737
rect 15257 31703 15280 31737
rect 15200 31417 15280 31703
rect 15200 31383 15223 31417
rect 15257 31383 15280 31417
rect 15200 31097 15280 31383
rect 15200 31063 15223 31097
rect 15257 31063 15280 31097
rect 15200 30777 15280 31063
rect 15200 30743 15223 30777
rect 15257 30743 15280 30777
rect 15200 30457 15280 30743
rect 15200 30423 15223 30457
rect 15257 30423 15280 30457
rect 15200 30400 15280 30423
rect 15360 32377 15440 32400
rect 15360 32343 15383 32377
rect 15417 32343 15440 32377
rect 15360 32057 15440 32343
rect 15360 32023 15383 32057
rect 15417 32023 15440 32057
rect 15360 31737 15440 32023
rect 15360 31703 15383 31737
rect 15417 31703 15440 31737
rect 15360 31417 15440 31703
rect 15360 31383 15383 31417
rect 15417 31383 15440 31417
rect 15360 31097 15440 31383
rect 15360 31063 15383 31097
rect 15417 31063 15440 31097
rect 15360 30777 15440 31063
rect 15360 30743 15383 30777
rect 15417 30743 15440 30777
rect 15360 30457 15440 30743
rect 15360 30423 15383 30457
rect 15417 30423 15440 30457
rect 15360 30400 15440 30423
rect 15520 32377 15600 32400
rect 15520 32343 15543 32377
rect 15577 32343 15600 32377
rect 15520 32057 15600 32343
rect 15520 32023 15543 32057
rect 15577 32023 15600 32057
rect 15520 31737 15600 32023
rect 15520 31703 15543 31737
rect 15577 31703 15600 31737
rect 15520 31417 15600 31703
rect 15520 31383 15543 31417
rect 15577 31383 15600 31417
rect 15520 31097 15600 31383
rect 15520 31063 15543 31097
rect 15577 31063 15600 31097
rect 15520 30777 15600 31063
rect 15520 30743 15543 30777
rect 15577 30743 15600 30777
rect 15520 30457 15600 30743
rect 15520 30423 15543 30457
rect 15577 30423 15600 30457
rect 15520 30400 15600 30423
rect 15680 32377 15760 32400
rect 15680 32343 15703 32377
rect 15737 32343 15760 32377
rect 15680 32057 15760 32343
rect 15680 32023 15703 32057
rect 15737 32023 15760 32057
rect 15680 31737 15760 32023
rect 15680 31703 15703 31737
rect 15737 31703 15760 31737
rect 15680 31417 15760 31703
rect 15680 31383 15703 31417
rect 15737 31383 15760 31417
rect 15680 31097 15760 31383
rect 15680 31063 15703 31097
rect 15737 31063 15760 31097
rect 15680 30777 15760 31063
rect 15680 30743 15703 30777
rect 15737 30743 15760 30777
rect 15680 30457 15760 30743
rect 15680 30423 15703 30457
rect 15737 30423 15760 30457
rect 15680 30400 15760 30423
rect 15840 32377 15920 32400
rect 15840 32343 15863 32377
rect 15897 32343 15920 32377
rect 15840 32057 15920 32343
rect 15840 32023 15863 32057
rect 15897 32023 15920 32057
rect 15840 31737 15920 32023
rect 15840 31703 15863 31737
rect 15897 31703 15920 31737
rect 15840 31417 15920 31703
rect 15840 31383 15863 31417
rect 15897 31383 15920 31417
rect 15840 31097 15920 31383
rect 15840 31063 15863 31097
rect 15897 31063 15920 31097
rect 15840 30777 15920 31063
rect 15840 30743 15863 30777
rect 15897 30743 15920 30777
rect 15840 30457 15920 30743
rect 15840 30423 15863 30457
rect 15897 30423 15920 30457
rect 15840 30400 15920 30423
rect 16000 32377 16080 32400
rect 16000 32343 16023 32377
rect 16057 32343 16080 32377
rect 16000 32057 16080 32343
rect 16000 32023 16023 32057
rect 16057 32023 16080 32057
rect 16000 31737 16080 32023
rect 16000 31703 16023 31737
rect 16057 31703 16080 31737
rect 16000 31417 16080 31703
rect 16000 31383 16023 31417
rect 16057 31383 16080 31417
rect 16000 31097 16080 31383
rect 16000 31063 16023 31097
rect 16057 31063 16080 31097
rect 16000 30777 16080 31063
rect 16000 30743 16023 30777
rect 16057 30743 16080 30777
rect 16000 30457 16080 30743
rect 16000 30423 16023 30457
rect 16057 30423 16080 30457
rect 16000 30400 16080 30423
rect 16160 32377 16240 32400
rect 16160 32343 16183 32377
rect 16217 32343 16240 32377
rect 16160 32057 16240 32343
rect 16160 32023 16183 32057
rect 16217 32023 16240 32057
rect 16160 31737 16240 32023
rect 16160 31703 16183 31737
rect 16217 31703 16240 31737
rect 16160 31417 16240 31703
rect 16160 31383 16183 31417
rect 16217 31383 16240 31417
rect 16160 31097 16240 31383
rect 16160 31063 16183 31097
rect 16217 31063 16240 31097
rect 16160 30777 16240 31063
rect 16160 30743 16183 30777
rect 16217 30743 16240 30777
rect 16160 30457 16240 30743
rect 16160 30423 16183 30457
rect 16217 30423 16240 30457
rect 16160 30400 16240 30423
rect 16320 32377 16400 32400
rect 16320 32343 16343 32377
rect 16377 32343 16400 32377
rect 16320 32057 16400 32343
rect 16320 32023 16343 32057
rect 16377 32023 16400 32057
rect 16320 31737 16400 32023
rect 16320 31703 16343 31737
rect 16377 31703 16400 31737
rect 16320 31417 16400 31703
rect 16320 31383 16343 31417
rect 16377 31383 16400 31417
rect 16320 31097 16400 31383
rect 16320 31063 16343 31097
rect 16377 31063 16400 31097
rect 16320 30777 16400 31063
rect 16320 30743 16343 30777
rect 16377 30743 16400 30777
rect 16320 30457 16400 30743
rect 16320 30423 16343 30457
rect 16377 30423 16400 30457
rect 16320 30400 16400 30423
rect 16480 32377 16560 32400
rect 16480 32343 16503 32377
rect 16537 32343 16560 32377
rect 16480 32057 16560 32343
rect 16480 32023 16503 32057
rect 16537 32023 16560 32057
rect 16480 31737 16560 32023
rect 16480 31703 16503 31737
rect 16537 31703 16560 31737
rect 16480 31417 16560 31703
rect 16480 31383 16503 31417
rect 16537 31383 16560 31417
rect 16480 31097 16560 31383
rect 16480 31063 16503 31097
rect 16537 31063 16560 31097
rect 16480 30777 16560 31063
rect 16480 30743 16503 30777
rect 16537 30743 16560 30777
rect 16480 30457 16560 30743
rect 16480 30423 16503 30457
rect 16537 30423 16560 30457
rect 16480 30400 16560 30423
rect 16640 32377 16720 32400
rect 16640 32343 16663 32377
rect 16697 32343 16720 32377
rect 16640 32057 16720 32343
rect 16640 32023 16663 32057
rect 16697 32023 16720 32057
rect 16640 31737 16720 32023
rect 16640 31703 16663 31737
rect 16697 31703 16720 31737
rect 16640 31417 16720 31703
rect 16640 31383 16663 31417
rect 16697 31383 16720 31417
rect 16640 31097 16720 31383
rect 16640 31063 16663 31097
rect 16697 31063 16720 31097
rect 16640 30777 16720 31063
rect 16640 30743 16663 30777
rect 16697 30743 16720 30777
rect 16640 30457 16720 30743
rect 16640 30423 16663 30457
rect 16697 30423 16720 30457
rect 16640 30400 16720 30423
rect 16800 32377 16880 32400
rect 16800 32343 16823 32377
rect 16857 32343 16880 32377
rect 16800 32057 16880 32343
rect 16800 32023 16823 32057
rect 16857 32023 16880 32057
rect 16800 31737 16880 32023
rect 16800 31703 16823 31737
rect 16857 31703 16880 31737
rect 16800 31417 16880 31703
rect 16800 31383 16823 31417
rect 16857 31383 16880 31417
rect 16800 31097 16880 31383
rect 16800 31063 16823 31097
rect 16857 31063 16880 31097
rect 16800 30777 16880 31063
rect 16800 30743 16823 30777
rect 16857 30743 16880 30777
rect 16800 30457 16880 30743
rect 16800 30423 16823 30457
rect 16857 30423 16880 30457
rect 16800 30400 16880 30423
rect 16960 32377 17040 32400
rect 16960 32343 16983 32377
rect 17017 32343 17040 32377
rect 16960 32057 17040 32343
rect 16960 32023 16983 32057
rect 17017 32023 17040 32057
rect 16960 31737 17040 32023
rect 16960 31703 16983 31737
rect 17017 31703 17040 31737
rect 16960 31417 17040 31703
rect 16960 31383 16983 31417
rect 17017 31383 17040 31417
rect 16960 31097 17040 31383
rect 16960 31063 16983 31097
rect 17017 31063 17040 31097
rect 16960 30777 17040 31063
rect 16960 30743 16983 30777
rect 17017 30743 17040 30777
rect 16960 30457 17040 30743
rect 16960 30423 16983 30457
rect 17017 30423 17040 30457
rect 16960 30400 17040 30423
rect 17120 32377 17200 32400
rect 17120 32343 17143 32377
rect 17177 32343 17200 32377
rect 17120 32057 17200 32343
rect 17120 32023 17143 32057
rect 17177 32023 17200 32057
rect 17120 31737 17200 32023
rect 17120 31703 17143 31737
rect 17177 31703 17200 31737
rect 17120 31417 17200 31703
rect 17120 31383 17143 31417
rect 17177 31383 17200 31417
rect 17120 31097 17200 31383
rect 17120 31063 17143 31097
rect 17177 31063 17200 31097
rect 17120 30777 17200 31063
rect 17120 30743 17143 30777
rect 17177 30743 17200 30777
rect 17120 30457 17200 30743
rect 17120 30423 17143 30457
rect 17177 30423 17200 30457
rect 17120 30400 17200 30423
rect 17280 32377 17360 32400
rect 17280 32343 17303 32377
rect 17337 32343 17360 32377
rect 17280 32057 17360 32343
rect 17280 32023 17303 32057
rect 17337 32023 17360 32057
rect 17280 31737 17360 32023
rect 17280 31703 17303 31737
rect 17337 31703 17360 31737
rect 17280 31417 17360 31703
rect 17280 31383 17303 31417
rect 17337 31383 17360 31417
rect 17280 31097 17360 31383
rect 17280 31063 17303 31097
rect 17337 31063 17360 31097
rect 17280 30777 17360 31063
rect 17280 30743 17303 30777
rect 17337 30743 17360 30777
rect 17280 30457 17360 30743
rect 17280 30423 17303 30457
rect 17337 30423 17360 30457
rect 17280 30400 17360 30423
rect 17440 32377 17520 32400
rect 17440 32343 17463 32377
rect 17497 32343 17520 32377
rect 17440 32057 17520 32343
rect 17440 32023 17463 32057
rect 17497 32023 17520 32057
rect 17440 31737 17520 32023
rect 17440 31703 17463 31737
rect 17497 31703 17520 31737
rect 17440 31417 17520 31703
rect 17440 31383 17463 31417
rect 17497 31383 17520 31417
rect 17440 31097 17520 31383
rect 17440 31063 17463 31097
rect 17497 31063 17520 31097
rect 17440 30777 17520 31063
rect 17440 30743 17463 30777
rect 17497 30743 17520 30777
rect 17440 30457 17520 30743
rect 17440 30423 17463 30457
rect 17497 30423 17520 30457
rect 17440 30400 17520 30423
rect 17600 32377 17680 32400
rect 17600 32343 17623 32377
rect 17657 32343 17680 32377
rect 17600 32057 17680 32343
rect 17600 32023 17623 32057
rect 17657 32023 17680 32057
rect 17600 31737 17680 32023
rect 17600 31703 17623 31737
rect 17657 31703 17680 31737
rect 17600 31417 17680 31703
rect 17600 31383 17623 31417
rect 17657 31383 17680 31417
rect 17600 31097 17680 31383
rect 17600 31063 17623 31097
rect 17657 31063 17680 31097
rect 17600 30777 17680 31063
rect 17600 30743 17623 30777
rect 17657 30743 17680 30777
rect 17600 30457 17680 30743
rect 17600 30423 17623 30457
rect 17657 30423 17680 30457
rect 17600 30400 17680 30423
rect 17760 32377 17840 32400
rect 17760 32343 17783 32377
rect 17817 32343 17840 32377
rect 17760 32057 17840 32343
rect 17760 32023 17783 32057
rect 17817 32023 17840 32057
rect 17760 31737 17840 32023
rect 17760 31703 17783 31737
rect 17817 31703 17840 31737
rect 17760 31417 17840 31703
rect 17760 31383 17783 31417
rect 17817 31383 17840 31417
rect 17760 31097 17840 31383
rect 17760 31063 17783 31097
rect 17817 31063 17840 31097
rect 17760 30777 17840 31063
rect 17760 30743 17783 30777
rect 17817 30743 17840 30777
rect 17760 30457 17840 30743
rect 17760 30423 17783 30457
rect 17817 30423 17840 30457
rect 17760 30400 17840 30423
rect 17920 32377 18000 32400
rect 17920 32343 17943 32377
rect 17977 32343 18000 32377
rect 17920 32057 18000 32343
rect 17920 32023 17943 32057
rect 17977 32023 18000 32057
rect 17920 31737 18000 32023
rect 17920 31703 17943 31737
rect 17977 31703 18000 31737
rect 17920 31417 18000 31703
rect 17920 31383 17943 31417
rect 17977 31383 18000 31417
rect 17920 31097 18000 31383
rect 17920 31063 17943 31097
rect 17977 31063 18000 31097
rect 17920 30777 18000 31063
rect 17920 30743 17943 30777
rect 17977 30743 18000 30777
rect 17920 30457 18000 30743
rect 17920 30423 17943 30457
rect 17977 30423 18000 30457
rect 17920 30400 18000 30423
rect 18080 32377 18160 32400
rect 18080 32343 18103 32377
rect 18137 32343 18160 32377
rect 18080 32057 18160 32343
rect 18080 32023 18103 32057
rect 18137 32023 18160 32057
rect 18080 31737 18160 32023
rect 18080 31703 18103 31737
rect 18137 31703 18160 31737
rect 18080 31417 18160 31703
rect 18080 31383 18103 31417
rect 18137 31383 18160 31417
rect 18080 31097 18160 31383
rect 18080 31063 18103 31097
rect 18137 31063 18160 31097
rect 18080 30777 18160 31063
rect 18080 30743 18103 30777
rect 18137 30743 18160 30777
rect 18080 30457 18160 30743
rect 18080 30423 18103 30457
rect 18137 30423 18160 30457
rect 18080 30400 18160 30423
rect 18240 32377 18320 32400
rect 18240 32343 18263 32377
rect 18297 32343 18320 32377
rect 18240 32057 18320 32343
rect 18240 32023 18263 32057
rect 18297 32023 18320 32057
rect 18240 31737 18320 32023
rect 18240 31703 18263 31737
rect 18297 31703 18320 31737
rect 18240 31417 18320 31703
rect 18240 31383 18263 31417
rect 18297 31383 18320 31417
rect 18240 31097 18320 31383
rect 18240 31063 18263 31097
rect 18297 31063 18320 31097
rect 18240 30777 18320 31063
rect 18240 30743 18263 30777
rect 18297 30743 18320 30777
rect 18240 30457 18320 30743
rect 18240 30423 18263 30457
rect 18297 30423 18320 30457
rect 18240 30400 18320 30423
rect 18400 32377 18480 32400
rect 18400 32343 18423 32377
rect 18457 32343 18480 32377
rect 18400 32057 18480 32343
rect 18400 32023 18423 32057
rect 18457 32023 18480 32057
rect 18400 31737 18480 32023
rect 18400 31703 18423 31737
rect 18457 31703 18480 31737
rect 18400 31417 18480 31703
rect 18400 31383 18423 31417
rect 18457 31383 18480 31417
rect 18400 31097 18480 31383
rect 18400 31063 18423 31097
rect 18457 31063 18480 31097
rect 18400 30777 18480 31063
rect 18400 30743 18423 30777
rect 18457 30743 18480 30777
rect 18400 30457 18480 30743
rect 18400 30423 18423 30457
rect 18457 30423 18480 30457
rect 18400 30400 18480 30423
rect 18560 32377 18640 32400
rect 18560 32343 18583 32377
rect 18617 32343 18640 32377
rect 18560 32057 18640 32343
rect 18560 32023 18583 32057
rect 18617 32023 18640 32057
rect 18560 31737 18640 32023
rect 18560 31703 18583 31737
rect 18617 31703 18640 31737
rect 18560 31417 18640 31703
rect 18560 31383 18583 31417
rect 18617 31383 18640 31417
rect 18560 31097 18640 31383
rect 18560 31063 18583 31097
rect 18617 31063 18640 31097
rect 18560 30777 18640 31063
rect 18560 30743 18583 30777
rect 18617 30743 18640 30777
rect 18560 30457 18640 30743
rect 18560 30423 18583 30457
rect 18617 30423 18640 30457
rect 18560 30400 18640 30423
rect 18720 32377 18800 32400
rect 18720 32343 18743 32377
rect 18777 32343 18800 32377
rect 18720 32057 18800 32343
rect 18720 32023 18743 32057
rect 18777 32023 18800 32057
rect 18720 31737 18800 32023
rect 18720 31703 18743 31737
rect 18777 31703 18800 31737
rect 18720 31417 18800 31703
rect 18720 31383 18743 31417
rect 18777 31383 18800 31417
rect 18720 31097 18800 31383
rect 18720 31063 18743 31097
rect 18777 31063 18800 31097
rect 18720 30777 18800 31063
rect 18720 30743 18743 30777
rect 18777 30743 18800 30777
rect 18720 30457 18800 30743
rect 18720 30423 18743 30457
rect 18777 30423 18800 30457
rect 18720 30400 18800 30423
rect 18880 32377 18960 32400
rect 18880 32343 18903 32377
rect 18937 32343 18960 32377
rect 18880 32057 18960 32343
rect 18880 32023 18903 32057
rect 18937 32023 18960 32057
rect 18880 31737 18960 32023
rect 18880 31703 18903 31737
rect 18937 31703 18960 31737
rect 18880 31417 18960 31703
rect 18880 31383 18903 31417
rect 18937 31383 18960 31417
rect 18880 31097 18960 31383
rect 18880 31063 18903 31097
rect 18937 31063 18960 31097
rect 18880 30777 18960 31063
rect 18880 30743 18903 30777
rect 18937 30743 18960 30777
rect 18880 30457 18960 30743
rect 18880 30423 18903 30457
rect 18937 30423 18960 30457
rect 18880 30400 18960 30423
rect 19040 30400 19120 32400
rect 19200 30400 19280 32400
rect 19360 30400 19440 32400
rect 19520 30400 19600 32400
rect 19680 30400 19760 32400
rect 19840 30400 19920 32400
rect 20000 30400 20080 32400
rect 20160 30400 20240 32400
rect 20320 30400 20400 32400
rect 20480 30400 20560 32400
rect 20640 30400 20720 32400
rect 20800 30400 20880 32400
rect 20960 30400 21040 32400
rect 21120 30400 21200 32400
rect 21280 30400 21360 32400
rect 21440 30400 21520 32400
rect 21600 30400 21680 32400
rect 21760 30400 21840 32400
rect 21920 30400 22000 32400
rect 22080 30400 22160 32400
rect 22240 30400 22320 32400
rect 22400 30400 22480 32400
rect 22560 30400 22640 32400
rect 22720 30400 22800 32400
rect 22880 30400 22960 32400
rect 23120 32377 23200 32400
rect 23120 32343 23143 32377
rect 23177 32343 23200 32377
rect 23120 32057 23200 32343
rect 23120 32023 23143 32057
rect 23177 32023 23200 32057
rect 23120 31737 23200 32023
rect 23120 31703 23143 31737
rect 23177 31703 23200 31737
rect 23120 31417 23200 31703
rect 23120 31383 23143 31417
rect 23177 31383 23200 31417
rect 23120 31097 23200 31383
rect 23120 31063 23143 31097
rect 23177 31063 23200 31097
rect 23120 30777 23200 31063
rect 23120 30743 23143 30777
rect 23177 30743 23200 30777
rect 23120 30457 23200 30743
rect 23120 30423 23143 30457
rect 23177 30423 23200 30457
rect 23120 30400 23200 30423
rect 23280 32377 23360 32400
rect 23280 32343 23303 32377
rect 23337 32343 23360 32377
rect 23280 32057 23360 32343
rect 23280 32023 23303 32057
rect 23337 32023 23360 32057
rect 23280 31737 23360 32023
rect 23280 31703 23303 31737
rect 23337 31703 23360 31737
rect 23280 31417 23360 31703
rect 23280 31383 23303 31417
rect 23337 31383 23360 31417
rect 23280 31097 23360 31383
rect 23280 31063 23303 31097
rect 23337 31063 23360 31097
rect 23280 30777 23360 31063
rect 23280 30743 23303 30777
rect 23337 30743 23360 30777
rect 23280 30457 23360 30743
rect 23280 30423 23303 30457
rect 23337 30423 23360 30457
rect 23280 30400 23360 30423
rect 23440 32377 23520 32400
rect 23440 32343 23463 32377
rect 23497 32343 23520 32377
rect 23440 32057 23520 32343
rect 23440 32023 23463 32057
rect 23497 32023 23520 32057
rect 23440 31737 23520 32023
rect 23440 31703 23463 31737
rect 23497 31703 23520 31737
rect 23440 31417 23520 31703
rect 23440 31383 23463 31417
rect 23497 31383 23520 31417
rect 23440 31097 23520 31383
rect 23440 31063 23463 31097
rect 23497 31063 23520 31097
rect 23440 30777 23520 31063
rect 23440 30743 23463 30777
rect 23497 30743 23520 30777
rect 23440 30457 23520 30743
rect 23440 30423 23463 30457
rect 23497 30423 23520 30457
rect 23440 30400 23520 30423
rect 23600 32377 23680 32400
rect 23600 32343 23623 32377
rect 23657 32343 23680 32377
rect 23600 32057 23680 32343
rect 23600 32023 23623 32057
rect 23657 32023 23680 32057
rect 23600 31737 23680 32023
rect 23600 31703 23623 31737
rect 23657 31703 23680 31737
rect 23600 31417 23680 31703
rect 23600 31383 23623 31417
rect 23657 31383 23680 31417
rect 23600 31097 23680 31383
rect 23600 31063 23623 31097
rect 23657 31063 23680 31097
rect 23600 30777 23680 31063
rect 23600 30743 23623 30777
rect 23657 30743 23680 30777
rect 23600 30457 23680 30743
rect 23600 30423 23623 30457
rect 23657 30423 23680 30457
rect 23600 30400 23680 30423
rect 23760 32377 23840 32400
rect 23760 32343 23783 32377
rect 23817 32343 23840 32377
rect 23760 32057 23840 32343
rect 23760 32023 23783 32057
rect 23817 32023 23840 32057
rect 23760 31737 23840 32023
rect 23760 31703 23783 31737
rect 23817 31703 23840 31737
rect 23760 31417 23840 31703
rect 23760 31383 23783 31417
rect 23817 31383 23840 31417
rect 23760 31097 23840 31383
rect 23760 31063 23783 31097
rect 23817 31063 23840 31097
rect 23760 30777 23840 31063
rect 23760 30743 23783 30777
rect 23817 30743 23840 30777
rect 23760 30457 23840 30743
rect 23760 30423 23783 30457
rect 23817 30423 23840 30457
rect 23760 30400 23840 30423
rect 23920 32377 24000 32400
rect 23920 32343 23943 32377
rect 23977 32343 24000 32377
rect 23920 32057 24000 32343
rect 23920 32023 23943 32057
rect 23977 32023 24000 32057
rect 23920 31737 24000 32023
rect 23920 31703 23943 31737
rect 23977 31703 24000 31737
rect 23920 31417 24000 31703
rect 23920 31383 23943 31417
rect 23977 31383 24000 31417
rect 23920 31097 24000 31383
rect 23920 31063 23943 31097
rect 23977 31063 24000 31097
rect 23920 30777 24000 31063
rect 23920 30743 23943 30777
rect 23977 30743 24000 30777
rect 23920 30457 24000 30743
rect 23920 30423 23943 30457
rect 23977 30423 24000 30457
rect 23920 30400 24000 30423
rect 24080 32377 24160 32400
rect 24080 32343 24103 32377
rect 24137 32343 24160 32377
rect 24080 32057 24160 32343
rect 24080 32023 24103 32057
rect 24137 32023 24160 32057
rect 24080 31737 24160 32023
rect 24080 31703 24103 31737
rect 24137 31703 24160 31737
rect 24080 31417 24160 31703
rect 24080 31383 24103 31417
rect 24137 31383 24160 31417
rect 24080 31097 24160 31383
rect 24080 31063 24103 31097
rect 24137 31063 24160 31097
rect 24080 30777 24160 31063
rect 24080 30743 24103 30777
rect 24137 30743 24160 30777
rect 24080 30457 24160 30743
rect 24080 30423 24103 30457
rect 24137 30423 24160 30457
rect 24080 30400 24160 30423
rect 24240 32377 24320 32400
rect 24240 32343 24263 32377
rect 24297 32343 24320 32377
rect 24240 32057 24320 32343
rect 24240 32023 24263 32057
rect 24297 32023 24320 32057
rect 24240 31737 24320 32023
rect 24240 31703 24263 31737
rect 24297 31703 24320 31737
rect 24240 31417 24320 31703
rect 24240 31383 24263 31417
rect 24297 31383 24320 31417
rect 24240 31097 24320 31383
rect 24240 31063 24263 31097
rect 24297 31063 24320 31097
rect 24240 30777 24320 31063
rect 24240 30743 24263 30777
rect 24297 30743 24320 30777
rect 24240 30457 24320 30743
rect 24240 30423 24263 30457
rect 24297 30423 24320 30457
rect 24240 30400 24320 30423
rect 24400 32377 24480 32400
rect 24400 32343 24423 32377
rect 24457 32343 24480 32377
rect 24400 32057 24480 32343
rect 24400 32023 24423 32057
rect 24457 32023 24480 32057
rect 24400 31737 24480 32023
rect 24400 31703 24423 31737
rect 24457 31703 24480 31737
rect 24400 31417 24480 31703
rect 24400 31383 24423 31417
rect 24457 31383 24480 31417
rect 24400 31097 24480 31383
rect 24400 31063 24423 31097
rect 24457 31063 24480 31097
rect 24400 30777 24480 31063
rect 24400 30743 24423 30777
rect 24457 30743 24480 30777
rect 24400 30457 24480 30743
rect 24400 30423 24423 30457
rect 24457 30423 24480 30457
rect 24400 30400 24480 30423
rect 24560 32377 24640 32400
rect 24560 32343 24583 32377
rect 24617 32343 24640 32377
rect 24560 32057 24640 32343
rect 24560 32023 24583 32057
rect 24617 32023 24640 32057
rect 24560 31737 24640 32023
rect 24560 31703 24583 31737
rect 24617 31703 24640 31737
rect 24560 31417 24640 31703
rect 24560 31383 24583 31417
rect 24617 31383 24640 31417
rect 24560 31097 24640 31383
rect 24560 31063 24583 31097
rect 24617 31063 24640 31097
rect 24560 30777 24640 31063
rect 24560 30743 24583 30777
rect 24617 30743 24640 30777
rect 24560 30457 24640 30743
rect 24560 30423 24583 30457
rect 24617 30423 24640 30457
rect 24560 30400 24640 30423
rect 24720 32377 24800 32400
rect 24720 32343 24743 32377
rect 24777 32343 24800 32377
rect 24720 32057 24800 32343
rect 24720 32023 24743 32057
rect 24777 32023 24800 32057
rect 24720 31737 24800 32023
rect 24720 31703 24743 31737
rect 24777 31703 24800 31737
rect 24720 31417 24800 31703
rect 24720 31383 24743 31417
rect 24777 31383 24800 31417
rect 24720 31097 24800 31383
rect 24720 31063 24743 31097
rect 24777 31063 24800 31097
rect 24720 30777 24800 31063
rect 24720 30743 24743 30777
rect 24777 30743 24800 30777
rect 24720 30457 24800 30743
rect 24720 30423 24743 30457
rect 24777 30423 24800 30457
rect 24720 30400 24800 30423
rect 24880 32377 24960 32400
rect 24880 32343 24903 32377
rect 24937 32343 24960 32377
rect 24880 32057 24960 32343
rect 24880 32023 24903 32057
rect 24937 32023 24960 32057
rect 24880 31737 24960 32023
rect 24880 31703 24903 31737
rect 24937 31703 24960 31737
rect 24880 31417 24960 31703
rect 24880 31383 24903 31417
rect 24937 31383 24960 31417
rect 24880 31097 24960 31383
rect 24880 31063 24903 31097
rect 24937 31063 24960 31097
rect 24880 30777 24960 31063
rect 24880 30743 24903 30777
rect 24937 30743 24960 30777
rect 24880 30457 24960 30743
rect 24880 30423 24903 30457
rect 24937 30423 24960 30457
rect 24880 30400 24960 30423
rect 25040 32377 25120 32400
rect 25040 32343 25063 32377
rect 25097 32343 25120 32377
rect 25040 32057 25120 32343
rect 25040 32023 25063 32057
rect 25097 32023 25120 32057
rect 25040 31737 25120 32023
rect 25040 31703 25063 31737
rect 25097 31703 25120 31737
rect 25040 31417 25120 31703
rect 25040 31383 25063 31417
rect 25097 31383 25120 31417
rect 25040 31097 25120 31383
rect 25040 31063 25063 31097
rect 25097 31063 25120 31097
rect 25040 30777 25120 31063
rect 25040 30743 25063 30777
rect 25097 30743 25120 30777
rect 25040 30457 25120 30743
rect 25040 30423 25063 30457
rect 25097 30423 25120 30457
rect 25040 30400 25120 30423
rect 25200 32377 25280 32400
rect 25200 32343 25223 32377
rect 25257 32343 25280 32377
rect 25200 32057 25280 32343
rect 25200 32023 25223 32057
rect 25257 32023 25280 32057
rect 25200 31737 25280 32023
rect 25200 31703 25223 31737
rect 25257 31703 25280 31737
rect 25200 31417 25280 31703
rect 25200 31383 25223 31417
rect 25257 31383 25280 31417
rect 25200 31097 25280 31383
rect 25200 31063 25223 31097
rect 25257 31063 25280 31097
rect 25200 30777 25280 31063
rect 25200 30743 25223 30777
rect 25257 30743 25280 30777
rect 25200 30457 25280 30743
rect 25200 30423 25223 30457
rect 25257 30423 25280 30457
rect 25200 30400 25280 30423
rect 25360 32377 25440 32400
rect 25360 32343 25383 32377
rect 25417 32343 25440 32377
rect 25360 32057 25440 32343
rect 25360 32023 25383 32057
rect 25417 32023 25440 32057
rect 25360 31737 25440 32023
rect 25360 31703 25383 31737
rect 25417 31703 25440 31737
rect 25360 31417 25440 31703
rect 25360 31383 25383 31417
rect 25417 31383 25440 31417
rect 25360 31097 25440 31383
rect 25360 31063 25383 31097
rect 25417 31063 25440 31097
rect 25360 30777 25440 31063
rect 25360 30743 25383 30777
rect 25417 30743 25440 30777
rect 25360 30457 25440 30743
rect 25360 30423 25383 30457
rect 25417 30423 25440 30457
rect 25360 30400 25440 30423
rect 25520 32377 25600 32400
rect 25520 32343 25543 32377
rect 25577 32343 25600 32377
rect 25520 32057 25600 32343
rect 25520 32023 25543 32057
rect 25577 32023 25600 32057
rect 25520 31737 25600 32023
rect 25520 31703 25543 31737
rect 25577 31703 25600 31737
rect 25520 31417 25600 31703
rect 25520 31383 25543 31417
rect 25577 31383 25600 31417
rect 25520 31097 25600 31383
rect 25520 31063 25543 31097
rect 25577 31063 25600 31097
rect 25520 30777 25600 31063
rect 25520 30743 25543 30777
rect 25577 30743 25600 30777
rect 25520 30457 25600 30743
rect 25520 30423 25543 30457
rect 25577 30423 25600 30457
rect 25520 30400 25600 30423
rect 25680 32377 25760 32400
rect 25680 32343 25703 32377
rect 25737 32343 25760 32377
rect 25680 32057 25760 32343
rect 25680 32023 25703 32057
rect 25737 32023 25760 32057
rect 25680 31737 25760 32023
rect 25680 31703 25703 31737
rect 25737 31703 25760 31737
rect 25680 31417 25760 31703
rect 25680 31383 25703 31417
rect 25737 31383 25760 31417
rect 25680 31097 25760 31383
rect 25680 31063 25703 31097
rect 25737 31063 25760 31097
rect 25680 30777 25760 31063
rect 25680 30743 25703 30777
rect 25737 30743 25760 30777
rect 25680 30457 25760 30743
rect 25680 30423 25703 30457
rect 25737 30423 25760 30457
rect 25680 30400 25760 30423
rect 25840 32377 25920 32400
rect 25840 32343 25863 32377
rect 25897 32343 25920 32377
rect 25840 32057 25920 32343
rect 25840 32023 25863 32057
rect 25897 32023 25920 32057
rect 25840 31737 25920 32023
rect 25840 31703 25863 31737
rect 25897 31703 25920 31737
rect 25840 31417 25920 31703
rect 25840 31383 25863 31417
rect 25897 31383 25920 31417
rect 25840 31097 25920 31383
rect 25840 31063 25863 31097
rect 25897 31063 25920 31097
rect 25840 30777 25920 31063
rect 25840 30743 25863 30777
rect 25897 30743 25920 30777
rect 25840 30457 25920 30743
rect 25840 30423 25863 30457
rect 25897 30423 25920 30457
rect 25840 30400 25920 30423
rect 26000 32377 26080 32400
rect 26000 32343 26023 32377
rect 26057 32343 26080 32377
rect 26000 32057 26080 32343
rect 26000 32023 26023 32057
rect 26057 32023 26080 32057
rect 26000 31737 26080 32023
rect 26000 31703 26023 31737
rect 26057 31703 26080 31737
rect 26000 31417 26080 31703
rect 26000 31383 26023 31417
rect 26057 31383 26080 31417
rect 26000 31097 26080 31383
rect 26000 31063 26023 31097
rect 26057 31063 26080 31097
rect 26000 30777 26080 31063
rect 26000 30743 26023 30777
rect 26057 30743 26080 30777
rect 26000 30457 26080 30743
rect 26000 30423 26023 30457
rect 26057 30423 26080 30457
rect 26000 30400 26080 30423
rect 26160 32377 26240 32400
rect 26160 32343 26183 32377
rect 26217 32343 26240 32377
rect 26160 32057 26240 32343
rect 26160 32023 26183 32057
rect 26217 32023 26240 32057
rect 26160 31737 26240 32023
rect 26160 31703 26183 31737
rect 26217 31703 26240 31737
rect 26160 31417 26240 31703
rect 26160 31383 26183 31417
rect 26217 31383 26240 31417
rect 26160 31097 26240 31383
rect 26160 31063 26183 31097
rect 26217 31063 26240 31097
rect 26160 30777 26240 31063
rect 26160 30743 26183 30777
rect 26217 30743 26240 30777
rect 26160 30457 26240 30743
rect 26160 30423 26183 30457
rect 26217 30423 26240 30457
rect 26160 30400 26240 30423
rect 26320 32377 26400 32400
rect 26320 32343 26343 32377
rect 26377 32343 26400 32377
rect 26320 32057 26400 32343
rect 26320 32023 26343 32057
rect 26377 32023 26400 32057
rect 26320 31737 26400 32023
rect 26320 31703 26343 31737
rect 26377 31703 26400 31737
rect 26320 31417 26400 31703
rect 26320 31383 26343 31417
rect 26377 31383 26400 31417
rect 26320 31097 26400 31383
rect 26320 31063 26343 31097
rect 26377 31063 26400 31097
rect 26320 30777 26400 31063
rect 26320 30743 26343 30777
rect 26377 30743 26400 30777
rect 26320 30457 26400 30743
rect 26320 30423 26343 30457
rect 26377 30423 26400 30457
rect 26320 30400 26400 30423
rect 26480 32377 26560 32400
rect 26480 32343 26503 32377
rect 26537 32343 26560 32377
rect 26480 32057 26560 32343
rect 26480 32023 26503 32057
rect 26537 32023 26560 32057
rect 26480 31737 26560 32023
rect 26480 31703 26503 31737
rect 26537 31703 26560 31737
rect 26480 31417 26560 31703
rect 26480 31383 26503 31417
rect 26537 31383 26560 31417
rect 26480 31097 26560 31383
rect 26480 31063 26503 31097
rect 26537 31063 26560 31097
rect 26480 30777 26560 31063
rect 26480 30743 26503 30777
rect 26537 30743 26560 30777
rect 26480 30457 26560 30743
rect 26480 30423 26503 30457
rect 26537 30423 26560 30457
rect 26480 30400 26560 30423
rect 26640 32377 26720 32400
rect 26640 32343 26663 32377
rect 26697 32343 26720 32377
rect 26640 32057 26720 32343
rect 26640 32023 26663 32057
rect 26697 32023 26720 32057
rect 26640 31737 26720 32023
rect 26640 31703 26663 31737
rect 26697 31703 26720 31737
rect 26640 31417 26720 31703
rect 26640 31383 26663 31417
rect 26697 31383 26720 31417
rect 26640 31097 26720 31383
rect 26640 31063 26663 31097
rect 26697 31063 26720 31097
rect 26640 30777 26720 31063
rect 26640 30743 26663 30777
rect 26697 30743 26720 30777
rect 26640 30457 26720 30743
rect 26640 30423 26663 30457
rect 26697 30423 26720 30457
rect 26640 30400 26720 30423
rect 26800 32377 26880 32400
rect 26800 32343 26823 32377
rect 26857 32343 26880 32377
rect 26800 32057 26880 32343
rect 26800 32023 26823 32057
rect 26857 32023 26880 32057
rect 26800 31737 26880 32023
rect 26800 31703 26823 31737
rect 26857 31703 26880 31737
rect 26800 31417 26880 31703
rect 26800 31383 26823 31417
rect 26857 31383 26880 31417
rect 26800 31097 26880 31383
rect 26800 31063 26823 31097
rect 26857 31063 26880 31097
rect 26800 30777 26880 31063
rect 26800 30743 26823 30777
rect 26857 30743 26880 30777
rect 26800 30457 26880 30743
rect 26800 30423 26823 30457
rect 26857 30423 26880 30457
rect 26800 30400 26880 30423
rect 26960 32377 27040 32400
rect 26960 32343 26983 32377
rect 27017 32343 27040 32377
rect 26960 32057 27040 32343
rect 26960 32023 26983 32057
rect 27017 32023 27040 32057
rect 26960 31737 27040 32023
rect 26960 31703 26983 31737
rect 27017 31703 27040 31737
rect 26960 31417 27040 31703
rect 26960 31383 26983 31417
rect 27017 31383 27040 31417
rect 26960 31097 27040 31383
rect 26960 31063 26983 31097
rect 27017 31063 27040 31097
rect 26960 30777 27040 31063
rect 26960 30743 26983 30777
rect 27017 30743 27040 30777
rect 26960 30457 27040 30743
rect 26960 30423 26983 30457
rect 27017 30423 27040 30457
rect 26960 30400 27040 30423
rect 27120 32377 27200 32400
rect 27120 32343 27143 32377
rect 27177 32343 27200 32377
rect 27120 32057 27200 32343
rect 27120 32023 27143 32057
rect 27177 32023 27200 32057
rect 27120 31737 27200 32023
rect 27120 31703 27143 31737
rect 27177 31703 27200 31737
rect 27120 31417 27200 31703
rect 27120 31383 27143 31417
rect 27177 31383 27200 31417
rect 27120 31097 27200 31383
rect 27120 31063 27143 31097
rect 27177 31063 27200 31097
rect 27120 30777 27200 31063
rect 27120 30743 27143 30777
rect 27177 30743 27200 30777
rect 27120 30457 27200 30743
rect 27120 30423 27143 30457
rect 27177 30423 27200 30457
rect 27120 30400 27200 30423
rect 27280 32377 27360 32400
rect 27280 32343 27303 32377
rect 27337 32343 27360 32377
rect 27280 32057 27360 32343
rect 27280 32023 27303 32057
rect 27337 32023 27360 32057
rect 27280 31737 27360 32023
rect 27280 31703 27303 31737
rect 27337 31703 27360 31737
rect 27280 31417 27360 31703
rect 27280 31383 27303 31417
rect 27337 31383 27360 31417
rect 27280 31097 27360 31383
rect 27280 31063 27303 31097
rect 27337 31063 27360 31097
rect 27280 30777 27360 31063
rect 27280 30743 27303 30777
rect 27337 30743 27360 30777
rect 27280 30457 27360 30743
rect 27280 30423 27303 30457
rect 27337 30423 27360 30457
rect 27280 30400 27360 30423
rect 27440 32377 27520 32400
rect 27440 32343 27463 32377
rect 27497 32343 27520 32377
rect 27440 32057 27520 32343
rect 27440 32023 27463 32057
rect 27497 32023 27520 32057
rect 27440 31737 27520 32023
rect 27440 31703 27463 31737
rect 27497 31703 27520 31737
rect 27440 31417 27520 31703
rect 27440 31383 27463 31417
rect 27497 31383 27520 31417
rect 27440 31097 27520 31383
rect 27440 31063 27463 31097
rect 27497 31063 27520 31097
rect 27440 30777 27520 31063
rect 27440 30743 27463 30777
rect 27497 30743 27520 30777
rect 27440 30457 27520 30743
rect 27440 30423 27463 30457
rect 27497 30423 27520 30457
rect 27440 30400 27520 30423
rect 27600 32377 27680 32400
rect 27600 32343 27623 32377
rect 27657 32343 27680 32377
rect 27600 32057 27680 32343
rect 27600 32023 27623 32057
rect 27657 32023 27680 32057
rect 27600 31737 27680 32023
rect 27600 31703 27623 31737
rect 27657 31703 27680 31737
rect 27600 31417 27680 31703
rect 27600 31383 27623 31417
rect 27657 31383 27680 31417
rect 27600 31097 27680 31383
rect 27600 31063 27623 31097
rect 27657 31063 27680 31097
rect 27600 30777 27680 31063
rect 27600 30743 27623 30777
rect 27657 30743 27680 30777
rect 27600 30457 27680 30743
rect 27600 30423 27623 30457
rect 27657 30423 27680 30457
rect 27600 30400 27680 30423
rect 27760 32377 27840 32400
rect 27760 32343 27783 32377
rect 27817 32343 27840 32377
rect 27760 32057 27840 32343
rect 27760 32023 27783 32057
rect 27817 32023 27840 32057
rect 27760 31737 27840 32023
rect 27760 31703 27783 31737
rect 27817 31703 27840 31737
rect 27760 31417 27840 31703
rect 27760 31383 27783 31417
rect 27817 31383 27840 31417
rect 27760 31097 27840 31383
rect 27760 31063 27783 31097
rect 27817 31063 27840 31097
rect 27760 30777 27840 31063
rect 27760 30743 27783 30777
rect 27817 30743 27840 30777
rect 27760 30457 27840 30743
rect 27760 30423 27783 30457
rect 27817 30423 27840 30457
rect 27760 30400 27840 30423
rect 27920 32377 28000 32400
rect 27920 32343 27943 32377
rect 27977 32343 28000 32377
rect 27920 32057 28000 32343
rect 27920 32023 27943 32057
rect 27977 32023 28000 32057
rect 27920 31737 28000 32023
rect 27920 31703 27943 31737
rect 27977 31703 28000 31737
rect 27920 31417 28000 31703
rect 27920 31383 27943 31417
rect 27977 31383 28000 31417
rect 27920 31097 28000 31383
rect 27920 31063 27943 31097
rect 27977 31063 28000 31097
rect 27920 30777 28000 31063
rect 27920 30743 27943 30777
rect 27977 30743 28000 30777
rect 27920 30457 28000 30743
rect 27920 30423 27943 30457
rect 27977 30423 28000 30457
rect 27920 30400 28000 30423
rect 28080 32377 28160 32400
rect 28080 32343 28103 32377
rect 28137 32343 28160 32377
rect 28080 32057 28160 32343
rect 28080 32023 28103 32057
rect 28137 32023 28160 32057
rect 28080 31737 28160 32023
rect 28080 31703 28103 31737
rect 28137 31703 28160 31737
rect 28080 31417 28160 31703
rect 28080 31383 28103 31417
rect 28137 31383 28160 31417
rect 28080 31097 28160 31383
rect 28080 31063 28103 31097
rect 28137 31063 28160 31097
rect 28080 30777 28160 31063
rect 28080 30743 28103 30777
rect 28137 30743 28160 30777
rect 28080 30457 28160 30743
rect 28080 30423 28103 30457
rect 28137 30423 28160 30457
rect 28080 30400 28160 30423
rect 28240 32377 28320 32400
rect 28240 32343 28263 32377
rect 28297 32343 28320 32377
rect 28240 32057 28320 32343
rect 28240 32023 28263 32057
rect 28297 32023 28320 32057
rect 28240 31737 28320 32023
rect 28240 31703 28263 31737
rect 28297 31703 28320 31737
rect 28240 31417 28320 31703
rect 28240 31383 28263 31417
rect 28297 31383 28320 31417
rect 28240 31097 28320 31383
rect 28240 31063 28263 31097
rect 28297 31063 28320 31097
rect 28240 30777 28320 31063
rect 28240 30743 28263 30777
rect 28297 30743 28320 30777
rect 28240 30457 28320 30743
rect 28240 30423 28263 30457
rect 28297 30423 28320 30457
rect 28240 30400 28320 30423
rect 28400 32377 28480 32400
rect 28400 32343 28423 32377
rect 28457 32343 28480 32377
rect 28400 32057 28480 32343
rect 28400 32023 28423 32057
rect 28457 32023 28480 32057
rect 28400 31737 28480 32023
rect 28400 31703 28423 31737
rect 28457 31703 28480 31737
rect 28400 31417 28480 31703
rect 28400 31383 28423 31417
rect 28457 31383 28480 31417
rect 28400 31097 28480 31383
rect 28400 31063 28423 31097
rect 28457 31063 28480 31097
rect 28400 30777 28480 31063
rect 28400 30743 28423 30777
rect 28457 30743 28480 30777
rect 28400 30457 28480 30743
rect 28400 30423 28423 30457
rect 28457 30423 28480 30457
rect 28400 30400 28480 30423
rect 28560 32377 28640 32400
rect 28560 32343 28583 32377
rect 28617 32343 28640 32377
rect 28560 32057 28640 32343
rect 28560 32023 28583 32057
rect 28617 32023 28640 32057
rect 28560 31737 28640 32023
rect 28560 31703 28583 31737
rect 28617 31703 28640 31737
rect 28560 31417 28640 31703
rect 28560 31383 28583 31417
rect 28617 31383 28640 31417
rect 28560 31097 28640 31383
rect 28560 31063 28583 31097
rect 28617 31063 28640 31097
rect 28560 30777 28640 31063
rect 28560 30743 28583 30777
rect 28617 30743 28640 30777
rect 28560 30457 28640 30743
rect 28560 30423 28583 30457
rect 28617 30423 28640 30457
rect 28560 30400 28640 30423
rect 28720 32377 28800 32400
rect 28720 32343 28743 32377
rect 28777 32343 28800 32377
rect 28720 32057 28800 32343
rect 28720 32023 28743 32057
rect 28777 32023 28800 32057
rect 28720 31737 28800 32023
rect 28720 31703 28743 31737
rect 28777 31703 28800 31737
rect 28720 31417 28800 31703
rect 28720 31383 28743 31417
rect 28777 31383 28800 31417
rect 28720 31097 28800 31383
rect 28720 31063 28743 31097
rect 28777 31063 28800 31097
rect 28720 30777 28800 31063
rect 28720 30743 28743 30777
rect 28777 30743 28800 30777
rect 28720 30457 28800 30743
rect 28720 30423 28743 30457
rect 28777 30423 28800 30457
rect 28720 30400 28800 30423
rect 28880 32377 28960 32400
rect 28880 32343 28903 32377
rect 28937 32343 28960 32377
rect 28880 32057 28960 32343
rect 28880 32023 28903 32057
rect 28937 32023 28960 32057
rect 28880 31737 28960 32023
rect 28880 31703 28903 31737
rect 28937 31703 28960 31737
rect 28880 31417 28960 31703
rect 28880 31383 28903 31417
rect 28937 31383 28960 31417
rect 28880 31097 28960 31383
rect 28880 31063 28903 31097
rect 28937 31063 28960 31097
rect 28880 30777 28960 31063
rect 28880 30743 28903 30777
rect 28937 30743 28960 30777
rect 28880 30457 28960 30743
rect 28880 30423 28903 30457
rect 28937 30423 28960 30457
rect 28880 30400 28960 30423
rect 29040 32377 29120 32400
rect 29040 32343 29063 32377
rect 29097 32343 29120 32377
rect 29040 32057 29120 32343
rect 29040 32023 29063 32057
rect 29097 32023 29120 32057
rect 29040 31737 29120 32023
rect 29040 31703 29063 31737
rect 29097 31703 29120 31737
rect 29040 31417 29120 31703
rect 29040 31383 29063 31417
rect 29097 31383 29120 31417
rect 29040 31097 29120 31383
rect 29040 31063 29063 31097
rect 29097 31063 29120 31097
rect 29040 30777 29120 31063
rect 29040 30743 29063 30777
rect 29097 30743 29120 30777
rect 29040 30457 29120 30743
rect 29040 30423 29063 30457
rect 29097 30423 29120 30457
rect 29040 30400 29120 30423
rect 29200 32377 29280 32400
rect 29200 32343 29223 32377
rect 29257 32343 29280 32377
rect 29200 32057 29280 32343
rect 29200 32023 29223 32057
rect 29257 32023 29280 32057
rect 29200 31737 29280 32023
rect 29200 31703 29223 31737
rect 29257 31703 29280 31737
rect 29200 31417 29280 31703
rect 29200 31383 29223 31417
rect 29257 31383 29280 31417
rect 29200 31097 29280 31383
rect 29200 31063 29223 31097
rect 29257 31063 29280 31097
rect 29200 30777 29280 31063
rect 29200 30743 29223 30777
rect 29257 30743 29280 30777
rect 29200 30457 29280 30743
rect 29200 30423 29223 30457
rect 29257 30423 29280 30457
rect 29200 30400 29280 30423
rect 29360 32377 29440 32400
rect 29360 32343 29383 32377
rect 29417 32343 29440 32377
rect 29360 32057 29440 32343
rect 29360 32023 29383 32057
rect 29417 32023 29440 32057
rect 29360 31737 29440 32023
rect 29360 31703 29383 31737
rect 29417 31703 29440 31737
rect 29360 31417 29440 31703
rect 29360 31383 29383 31417
rect 29417 31383 29440 31417
rect 29360 31097 29440 31383
rect 29360 31063 29383 31097
rect 29417 31063 29440 31097
rect 29360 30777 29440 31063
rect 29360 30743 29383 30777
rect 29417 30743 29440 30777
rect 29360 30457 29440 30743
rect 29360 30423 29383 30457
rect 29417 30423 29440 30457
rect 29360 30400 29440 30423
rect 29520 30400 29600 32400
rect 29680 30400 29760 32400
rect 29840 30400 29920 32400
rect 30000 30400 30080 32400
rect 30160 30400 30240 32400
rect 30320 30400 30400 32400
rect 30480 30400 30560 32400
rect 30640 30400 30720 32400
rect 30800 30400 30880 32400
rect 30960 30400 31040 32400
rect 31120 30400 31200 32400
rect 31280 30400 31360 32400
rect 31440 30400 31520 32400
rect 31600 30400 31680 32400
rect 31760 30400 31840 32400
rect 31920 30400 32000 32400
rect 32080 30400 32160 32400
rect 32240 30400 32320 32400
rect 32400 30400 32480 32400
rect 32560 30400 32640 32400
rect 32720 30400 32800 32400
rect 32880 30400 32960 32400
rect 33040 30400 33120 32400
rect 33200 30400 33280 32400
rect 33360 30400 33440 32400
rect 33520 32377 33600 32400
rect 33520 32343 33543 32377
rect 33577 32343 33600 32377
rect 33520 32057 33600 32343
rect 33520 32023 33543 32057
rect 33577 32023 33600 32057
rect 33520 31737 33600 32023
rect 33520 31703 33543 31737
rect 33577 31703 33600 31737
rect 33520 31417 33600 31703
rect 33520 31383 33543 31417
rect 33577 31383 33600 31417
rect 33520 31097 33600 31383
rect 33520 31063 33543 31097
rect 33577 31063 33600 31097
rect 33520 30777 33600 31063
rect 33520 30743 33543 30777
rect 33577 30743 33600 30777
rect 33520 30457 33600 30743
rect 33520 30423 33543 30457
rect 33577 30423 33600 30457
rect 33520 30400 33600 30423
rect 33680 32377 33760 32400
rect 33680 32343 33703 32377
rect 33737 32343 33760 32377
rect 33680 32057 33760 32343
rect 33680 32023 33703 32057
rect 33737 32023 33760 32057
rect 33680 31737 33760 32023
rect 33680 31703 33703 31737
rect 33737 31703 33760 31737
rect 33680 31417 33760 31703
rect 33680 31383 33703 31417
rect 33737 31383 33760 31417
rect 33680 31097 33760 31383
rect 33680 31063 33703 31097
rect 33737 31063 33760 31097
rect 33680 30777 33760 31063
rect 33680 30743 33703 30777
rect 33737 30743 33760 30777
rect 33680 30457 33760 30743
rect 33680 30423 33703 30457
rect 33737 30423 33760 30457
rect 33680 30400 33760 30423
rect 33840 32377 33920 32400
rect 33840 32343 33863 32377
rect 33897 32343 33920 32377
rect 33840 32057 33920 32343
rect 33840 32023 33863 32057
rect 33897 32023 33920 32057
rect 33840 31737 33920 32023
rect 33840 31703 33863 31737
rect 33897 31703 33920 31737
rect 33840 31417 33920 31703
rect 33840 31383 33863 31417
rect 33897 31383 33920 31417
rect 33840 31097 33920 31383
rect 33840 31063 33863 31097
rect 33897 31063 33920 31097
rect 33840 30777 33920 31063
rect 33840 30743 33863 30777
rect 33897 30743 33920 30777
rect 33840 30457 33920 30743
rect 33840 30423 33863 30457
rect 33897 30423 33920 30457
rect 33840 30400 33920 30423
rect 34000 32377 34080 32400
rect 34000 32343 34023 32377
rect 34057 32343 34080 32377
rect 34000 32057 34080 32343
rect 34000 32023 34023 32057
rect 34057 32023 34080 32057
rect 34000 31737 34080 32023
rect 34000 31703 34023 31737
rect 34057 31703 34080 31737
rect 34000 31417 34080 31703
rect 34000 31383 34023 31417
rect 34057 31383 34080 31417
rect 34000 31097 34080 31383
rect 34000 31063 34023 31097
rect 34057 31063 34080 31097
rect 34000 30777 34080 31063
rect 34000 30743 34023 30777
rect 34057 30743 34080 30777
rect 34000 30457 34080 30743
rect 34000 30423 34023 30457
rect 34057 30423 34080 30457
rect 34000 30400 34080 30423
rect 34160 32377 34240 32400
rect 34160 32343 34183 32377
rect 34217 32343 34240 32377
rect 34160 32057 34240 32343
rect 34160 32023 34183 32057
rect 34217 32023 34240 32057
rect 34160 31737 34240 32023
rect 34160 31703 34183 31737
rect 34217 31703 34240 31737
rect 34160 31417 34240 31703
rect 34160 31383 34183 31417
rect 34217 31383 34240 31417
rect 34160 31097 34240 31383
rect 34160 31063 34183 31097
rect 34217 31063 34240 31097
rect 34160 30777 34240 31063
rect 34160 30743 34183 30777
rect 34217 30743 34240 30777
rect 34160 30457 34240 30743
rect 34160 30423 34183 30457
rect 34217 30423 34240 30457
rect 34160 30400 34240 30423
rect 34320 32377 34400 32400
rect 34320 32343 34343 32377
rect 34377 32343 34400 32377
rect 34320 32057 34400 32343
rect 34320 32023 34343 32057
rect 34377 32023 34400 32057
rect 34320 31737 34400 32023
rect 34320 31703 34343 31737
rect 34377 31703 34400 31737
rect 34320 31417 34400 31703
rect 34320 31383 34343 31417
rect 34377 31383 34400 31417
rect 34320 31097 34400 31383
rect 34320 31063 34343 31097
rect 34377 31063 34400 31097
rect 34320 30777 34400 31063
rect 34320 30743 34343 30777
rect 34377 30743 34400 30777
rect 34320 30457 34400 30743
rect 34320 30423 34343 30457
rect 34377 30423 34400 30457
rect 34320 30400 34400 30423
rect 34480 32377 34560 32400
rect 34480 32343 34503 32377
rect 34537 32343 34560 32377
rect 34480 32057 34560 32343
rect 34480 32023 34503 32057
rect 34537 32023 34560 32057
rect 34480 31737 34560 32023
rect 34480 31703 34503 31737
rect 34537 31703 34560 31737
rect 34480 31417 34560 31703
rect 34480 31383 34503 31417
rect 34537 31383 34560 31417
rect 34480 31097 34560 31383
rect 34480 31063 34503 31097
rect 34537 31063 34560 31097
rect 34480 30777 34560 31063
rect 34480 30743 34503 30777
rect 34537 30743 34560 30777
rect 34480 30457 34560 30743
rect 34480 30423 34503 30457
rect 34537 30423 34560 30457
rect 34480 30400 34560 30423
rect 34640 32377 34720 32400
rect 34640 32343 34663 32377
rect 34697 32343 34720 32377
rect 34640 32057 34720 32343
rect 34640 32023 34663 32057
rect 34697 32023 34720 32057
rect 34640 31737 34720 32023
rect 34640 31703 34663 31737
rect 34697 31703 34720 31737
rect 34640 31417 34720 31703
rect 34640 31383 34663 31417
rect 34697 31383 34720 31417
rect 34640 31097 34720 31383
rect 34640 31063 34663 31097
rect 34697 31063 34720 31097
rect 34640 30777 34720 31063
rect 34640 30743 34663 30777
rect 34697 30743 34720 30777
rect 34640 30457 34720 30743
rect 34640 30423 34663 30457
rect 34697 30423 34720 30457
rect 34640 30400 34720 30423
rect 34800 32377 34880 32400
rect 34800 32343 34823 32377
rect 34857 32343 34880 32377
rect 34800 32057 34880 32343
rect 34800 32023 34823 32057
rect 34857 32023 34880 32057
rect 34800 31737 34880 32023
rect 34800 31703 34823 31737
rect 34857 31703 34880 31737
rect 34800 31417 34880 31703
rect 34800 31383 34823 31417
rect 34857 31383 34880 31417
rect 34800 31097 34880 31383
rect 34800 31063 34823 31097
rect 34857 31063 34880 31097
rect 34800 30777 34880 31063
rect 34800 30743 34823 30777
rect 34857 30743 34880 30777
rect 34800 30457 34880 30743
rect 34800 30423 34823 30457
rect 34857 30423 34880 30457
rect 34800 30400 34880 30423
rect 34960 32377 35040 32400
rect 34960 32343 34983 32377
rect 35017 32343 35040 32377
rect 34960 32057 35040 32343
rect 34960 32023 34983 32057
rect 35017 32023 35040 32057
rect 34960 31737 35040 32023
rect 34960 31703 34983 31737
rect 35017 31703 35040 31737
rect 34960 31417 35040 31703
rect 34960 31383 34983 31417
rect 35017 31383 35040 31417
rect 34960 31097 35040 31383
rect 34960 31063 34983 31097
rect 35017 31063 35040 31097
rect 34960 30777 35040 31063
rect 34960 30743 34983 30777
rect 35017 30743 35040 30777
rect 34960 30457 35040 30743
rect 34960 30423 34983 30457
rect 35017 30423 35040 30457
rect 34960 30400 35040 30423
rect 35120 32377 35200 32400
rect 35120 32343 35143 32377
rect 35177 32343 35200 32377
rect 35120 32057 35200 32343
rect 35120 32023 35143 32057
rect 35177 32023 35200 32057
rect 35120 31737 35200 32023
rect 35120 31703 35143 31737
rect 35177 31703 35200 31737
rect 35120 31417 35200 31703
rect 35120 31383 35143 31417
rect 35177 31383 35200 31417
rect 35120 31097 35200 31383
rect 35120 31063 35143 31097
rect 35177 31063 35200 31097
rect 35120 30777 35200 31063
rect 35120 30743 35143 30777
rect 35177 30743 35200 30777
rect 35120 30457 35200 30743
rect 35120 30423 35143 30457
rect 35177 30423 35200 30457
rect 35120 30400 35200 30423
rect 35280 32377 35360 32400
rect 35280 32343 35303 32377
rect 35337 32343 35360 32377
rect 35280 32057 35360 32343
rect 35280 32023 35303 32057
rect 35337 32023 35360 32057
rect 35280 31737 35360 32023
rect 35280 31703 35303 31737
rect 35337 31703 35360 31737
rect 35280 31417 35360 31703
rect 35280 31383 35303 31417
rect 35337 31383 35360 31417
rect 35280 31097 35360 31383
rect 35280 31063 35303 31097
rect 35337 31063 35360 31097
rect 35280 30777 35360 31063
rect 35280 30743 35303 30777
rect 35337 30743 35360 30777
rect 35280 30457 35360 30743
rect 35280 30423 35303 30457
rect 35337 30423 35360 30457
rect 35280 30400 35360 30423
rect 35440 32377 35520 32400
rect 35440 32343 35463 32377
rect 35497 32343 35520 32377
rect 35440 32057 35520 32343
rect 35440 32023 35463 32057
rect 35497 32023 35520 32057
rect 35440 31737 35520 32023
rect 35440 31703 35463 31737
rect 35497 31703 35520 31737
rect 35440 31417 35520 31703
rect 35440 31383 35463 31417
rect 35497 31383 35520 31417
rect 35440 31097 35520 31383
rect 35440 31063 35463 31097
rect 35497 31063 35520 31097
rect 35440 30777 35520 31063
rect 35440 30743 35463 30777
rect 35497 30743 35520 30777
rect 35440 30457 35520 30743
rect 35440 30423 35463 30457
rect 35497 30423 35520 30457
rect 35440 30400 35520 30423
rect 35600 32377 35680 32400
rect 35600 32343 35623 32377
rect 35657 32343 35680 32377
rect 35600 32057 35680 32343
rect 35600 32023 35623 32057
rect 35657 32023 35680 32057
rect 35600 31737 35680 32023
rect 35600 31703 35623 31737
rect 35657 31703 35680 31737
rect 35600 31417 35680 31703
rect 35600 31383 35623 31417
rect 35657 31383 35680 31417
rect 35600 31097 35680 31383
rect 35600 31063 35623 31097
rect 35657 31063 35680 31097
rect 35600 30777 35680 31063
rect 35600 30743 35623 30777
rect 35657 30743 35680 30777
rect 35600 30457 35680 30743
rect 35600 30423 35623 30457
rect 35657 30423 35680 30457
rect 35600 30400 35680 30423
rect 35760 32377 35840 32400
rect 35760 32343 35783 32377
rect 35817 32343 35840 32377
rect 35760 32057 35840 32343
rect 35760 32023 35783 32057
rect 35817 32023 35840 32057
rect 35760 31737 35840 32023
rect 35760 31703 35783 31737
rect 35817 31703 35840 31737
rect 35760 31417 35840 31703
rect 35760 31383 35783 31417
rect 35817 31383 35840 31417
rect 35760 31097 35840 31383
rect 35760 31063 35783 31097
rect 35817 31063 35840 31097
rect 35760 30777 35840 31063
rect 35760 30743 35783 30777
rect 35817 30743 35840 30777
rect 35760 30457 35840 30743
rect 35760 30423 35783 30457
rect 35817 30423 35840 30457
rect 35760 30400 35840 30423
rect 35920 32377 36000 32400
rect 35920 32343 35943 32377
rect 35977 32343 36000 32377
rect 35920 32057 36000 32343
rect 35920 32023 35943 32057
rect 35977 32023 36000 32057
rect 35920 31737 36000 32023
rect 35920 31703 35943 31737
rect 35977 31703 36000 31737
rect 35920 31417 36000 31703
rect 35920 31383 35943 31417
rect 35977 31383 36000 31417
rect 35920 31097 36000 31383
rect 35920 31063 35943 31097
rect 35977 31063 36000 31097
rect 35920 30777 36000 31063
rect 35920 30743 35943 30777
rect 35977 30743 36000 30777
rect 35920 30457 36000 30743
rect 35920 30423 35943 30457
rect 35977 30423 36000 30457
rect 35920 30400 36000 30423
rect 36080 32377 36160 32400
rect 36080 32343 36103 32377
rect 36137 32343 36160 32377
rect 36080 32057 36160 32343
rect 36080 32023 36103 32057
rect 36137 32023 36160 32057
rect 36080 31737 36160 32023
rect 36080 31703 36103 31737
rect 36137 31703 36160 31737
rect 36080 31417 36160 31703
rect 36080 31383 36103 31417
rect 36137 31383 36160 31417
rect 36080 31097 36160 31383
rect 36080 31063 36103 31097
rect 36137 31063 36160 31097
rect 36080 30777 36160 31063
rect 36080 30743 36103 30777
rect 36137 30743 36160 30777
rect 36080 30457 36160 30743
rect 36080 30423 36103 30457
rect 36137 30423 36160 30457
rect 36080 30400 36160 30423
rect 36240 32377 36320 32400
rect 36240 32343 36263 32377
rect 36297 32343 36320 32377
rect 36240 32057 36320 32343
rect 36240 32023 36263 32057
rect 36297 32023 36320 32057
rect 36240 31737 36320 32023
rect 36240 31703 36263 31737
rect 36297 31703 36320 31737
rect 36240 31417 36320 31703
rect 36240 31383 36263 31417
rect 36297 31383 36320 31417
rect 36240 31097 36320 31383
rect 36240 31063 36263 31097
rect 36297 31063 36320 31097
rect 36240 30777 36320 31063
rect 36240 30743 36263 30777
rect 36297 30743 36320 30777
rect 36240 30457 36320 30743
rect 36240 30423 36263 30457
rect 36297 30423 36320 30457
rect 36240 30400 36320 30423
rect 36400 32377 36480 32400
rect 36400 32343 36423 32377
rect 36457 32343 36480 32377
rect 36400 32057 36480 32343
rect 36400 32023 36423 32057
rect 36457 32023 36480 32057
rect 36400 31737 36480 32023
rect 36400 31703 36423 31737
rect 36457 31703 36480 31737
rect 36400 31417 36480 31703
rect 36400 31383 36423 31417
rect 36457 31383 36480 31417
rect 36400 31097 36480 31383
rect 36400 31063 36423 31097
rect 36457 31063 36480 31097
rect 36400 30777 36480 31063
rect 36400 30743 36423 30777
rect 36457 30743 36480 30777
rect 36400 30457 36480 30743
rect 36400 30423 36423 30457
rect 36457 30423 36480 30457
rect 36400 30400 36480 30423
rect 36560 32377 36640 32400
rect 36560 32343 36583 32377
rect 36617 32343 36640 32377
rect 36560 32057 36640 32343
rect 36560 32023 36583 32057
rect 36617 32023 36640 32057
rect 36560 31737 36640 32023
rect 36560 31703 36583 31737
rect 36617 31703 36640 31737
rect 36560 31417 36640 31703
rect 36560 31383 36583 31417
rect 36617 31383 36640 31417
rect 36560 31097 36640 31383
rect 36560 31063 36583 31097
rect 36617 31063 36640 31097
rect 36560 30777 36640 31063
rect 36560 30743 36583 30777
rect 36617 30743 36640 30777
rect 36560 30457 36640 30743
rect 36560 30423 36583 30457
rect 36617 30423 36640 30457
rect 36560 30400 36640 30423
rect 36720 32377 36800 32400
rect 36720 32343 36743 32377
rect 36777 32343 36800 32377
rect 36720 32057 36800 32343
rect 36720 32023 36743 32057
rect 36777 32023 36800 32057
rect 36720 31737 36800 32023
rect 36720 31703 36743 31737
rect 36777 31703 36800 31737
rect 36720 31417 36800 31703
rect 36720 31383 36743 31417
rect 36777 31383 36800 31417
rect 36720 31097 36800 31383
rect 36720 31063 36743 31097
rect 36777 31063 36800 31097
rect 36720 30777 36800 31063
rect 36720 30743 36743 30777
rect 36777 30743 36800 30777
rect 36720 30457 36800 30743
rect 36720 30423 36743 30457
rect 36777 30423 36800 30457
rect 36720 30400 36800 30423
rect 36880 32377 36960 32400
rect 36880 32343 36903 32377
rect 36937 32343 36960 32377
rect 36880 32057 36960 32343
rect 36880 32023 36903 32057
rect 36937 32023 36960 32057
rect 36880 31737 36960 32023
rect 36880 31703 36903 31737
rect 36937 31703 36960 31737
rect 36880 31417 36960 31703
rect 36880 31383 36903 31417
rect 36937 31383 36960 31417
rect 36880 31097 36960 31383
rect 36880 31063 36903 31097
rect 36937 31063 36960 31097
rect 36880 30777 36960 31063
rect 36880 30743 36903 30777
rect 36937 30743 36960 30777
rect 36880 30457 36960 30743
rect 36880 30423 36903 30457
rect 36937 30423 36960 30457
rect 36880 30400 36960 30423
rect 37040 32377 37120 32400
rect 37040 32343 37063 32377
rect 37097 32343 37120 32377
rect 37040 32057 37120 32343
rect 37040 32023 37063 32057
rect 37097 32023 37120 32057
rect 37040 31737 37120 32023
rect 37040 31703 37063 31737
rect 37097 31703 37120 31737
rect 37040 31417 37120 31703
rect 37040 31383 37063 31417
rect 37097 31383 37120 31417
rect 37040 31097 37120 31383
rect 37040 31063 37063 31097
rect 37097 31063 37120 31097
rect 37040 30777 37120 31063
rect 37040 30743 37063 30777
rect 37097 30743 37120 30777
rect 37040 30457 37120 30743
rect 37040 30423 37063 30457
rect 37097 30423 37120 30457
rect 37040 30400 37120 30423
rect 37200 32377 37280 32400
rect 37200 32343 37223 32377
rect 37257 32343 37280 32377
rect 37200 32057 37280 32343
rect 37200 32023 37223 32057
rect 37257 32023 37280 32057
rect 37200 31737 37280 32023
rect 37200 31703 37223 31737
rect 37257 31703 37280 31737
rect 37200 31417 37280 31703
rect 37200 31383 37223 31417
rect 37257 31383 37280 31417
rect 37200 31097 37280 31383
rect 37200 31063 37223 31097
rect 37257 31063 37280 31097
rect 37200 30777 37280 31063
rect 37200 30743 37223 30777
rect 37257 30743 37280 30777
rect 37200 30457 37280 30743
rect 37200 30423 37223 30457
rect 37257 30423 37280 30457
rect 37200 30400 37280 30423
rect 37360 32377 37440 32400
rect 37360 32343 37383 32377
rect 37417 32343 37440 32377
rect 37360 32057 37440 32343
rect 37360 32023 37383 32057
rect 37417 32023 37440 32057
rect 37360 31737 37440 32023
rect 37360 31703 37383 31737
rect 37417 31703 37440 31737
rect 37360 31417 37440 31703
rect 37360 31383 37383 31417
rect 37417 31383 37440 31417
rect 37360 31097 37440 31383
rect 37360 31063 37383 31097
rect 37417 31063 37440 31097
rect 37360 30777 37440 31063
rect 37360 30743 37383 30777
rect 37417 30743 37440 30777
rect 37360 30457 37440 30743
rect 37360 30423 37383 30457
rect 37417 30423 37440 30457
rect 37360 30400 37440 30423
rect 37520 32377 37600 32400
rect 37520 32343 37543 32377
rect 37577 32343 37600 32377
rect 37520 32057 37600 32343
rect 37520 32023 37543 32057
rect 37577 32023 37600 32057
rect 37520 31737 37600 32023
rect 37520 31703 37543 31737
rect 37577 31703 37600 31737
rect 37520 31417 37600 31703
rect 37520 31383 37543 31417
rect 37577 31383 37600 31417
rect 37520 31097 37600 31383
rect 37520 31063 37543 31097
rect 37577 31063 37600 31097
rect 37520 30777 37600 31063
rect 37520 30743 37543 30777
rect 37577 30743 37600 30777
rect 37520 30457 37600 30743
rect 37520 30423 37543 30457
rect 37577 30423 37600 30457
rect 37520 30400 37600 30423
rect 37680 32377 37760 32400
rect 37680 32343 37703 32377
rect 37737 32343 37760 32377
rect 37680 32057 37760 32343
rect 37680 32023 37703 32057
rect 37737 32023 37760 32057
rect 37680 31737 37760 32023
rect 37680 31703 37703 31737
rect 37737 31703 37760 31737
rect 37680 31417 37760 31703
rect 37680 31383 37703 31417
rect 37737 31383 37760 31417
rect 37680 31097 37760 31383
rect 37680 31063 37703 31097
rect 37737 31063 37760 31097
rect 37680 30777 37760 31063
rect 37680 30743 37703 30777
rect 37737 30743 37760 30777
rect 37680 30457 37760 30743
rect 37680 30423 37703 30457
rect 37737 30423 37760 30457
rect 37680 30400 37760 30423
rect 37840 32377 37920 32400
rect 37840 32343 37863 32377
rect 37897 32343 37920 32377
rect 37840 32057 37920 32343
rect 37840 32023 37863 32057
rect 37897 32023 37920 32057
rect 37840 31737 37920 32023
rect 37840 31703 37863 31737
rect 37897 31703 37920 31737
rect 37840 31417 37920 31703
rect 37840 31383 37863 31417
rect 37897 31383 37920 31417
rect 37840 31097 37920 31383
rect 37840 31063 37863 31097
rect 37897 31063 37920 31097
rect 37840 30777 37920 31063
rect 37840 30743 37863 30777
rect 37897 30743 37920 30777
rect 37840 30457 37920 30743
rect 37840 30423 37863 30457
rect 37897 30423 37920 30457
rect 37840 30400 37920 30423
rect 38000 32377 38080 32400
rect 38000 32343 38023 32377
rect 38057 32343 38080 32377
rect 38000 32057 38080 32343
rect 38000 32023 38023 32057
rect 38057 32023 38080 32057
rect 38000 31737 38080 32023
rect 38000 31703 38023 31737
rect 38057 31703 38080 31737
rect 38000 31417 38080 31703
rect 38000 31383 38023 31417
rect 38057 31383 38080 31417
rect 38000 31097 38080 31383
rect 38000 31063 38023 31097
rect 38057 31063 38080 31097
rect 38000 30777 38080 31063
rect 38000 30743 38023 30777
rect 38057 30743 38080 30777
rect 38000 30457 38080 30743
rect 38000 30423 38023 30457
rect 38057 30423 38080 30457
rect 38000 30400 38080 30423
rect 38160 32377 38240 32400
rect 38160 32343 38183 32377
rect 38217 32343 38240 32377
rect 38160 32057 38240 32343
rect 38160 32023 38183 32057
rect 38217 32023 38240 32057
rect 38160 31737 38240 32023
rect 38160 31703 38183 31737
rect 38217 31703 38240 31737
rect 38160 31417 38240 31703
rect 38160 31383 38183 31417
rect 38217 31383 38240 31417
rect 38160 31097 38240 31383
rect 38160 31063 38183 31097
rect 38217 31063 38240 31097
rect 38160 30777 38240 31063
rect 38160 30743 38183 30777
rect 38217 30743 38240 30777
rect 38160 30457 38240 30743
rect 38160 30423 38183 30457
rect 38217 30423 38240 30457
rect 38160 30400 38240 30423
rect 38320 32377 38400 32400
rect 38320 32343 38343 32377
rect 38377 32343 38400 32377
rect 38320 32057 38400 32343
rect 38320 32023 38343 32057
rect 38377 32023 38400 32057
rect 38320 31737 38400 32023
rect 38320 31703 38343 31737
rect 38377 31703 38400 31737
rect 38320 31417 38400 31703
rect 38320 31383 38343 31417
rect 38377 31383 38400 31417
rect 38320 31097 38400 31383
rect 38320 31063 38343 31097
rect 38377 31063 38400 31097
rect 38320 30777 38400 31063
rect 38320 30743 38343 30777
rect 38377 30743 38400 30777
rect 38320 30457 38400 30743
rect 38320 30423 38343 30457
rect 38377 30423 38400 30457
rect 38320 30400 38400 30423
rect 38480 32377 38560 32400
rect 38480 32343 38503 32377
rect 38537 32343 38560 32377
rect 38480 32057 38560 32343
rect 38480 32023 38503 32057
rect 38537 32023 38560 32057
rect 38480 31737 38560 32023
rect 38480 31703 38503 31737
rect 38537 31703 38560 31737
rect 38480 31417 38560 31703
rect 38480 31383 38503 31417
rect 38537 31383 38560 31417
rect 38480 31097 38560 31383
rect 38480 31063 38503 31097
rect 38537 31063 38560 31097
rect 38480 30777 38560 31063
rect 38480 30743 38503 30777
rect 38537 30743 38560 30777
rect 38480 30457 38560 30743
rect 38480 30423 38503 30457
rect 38537 30423 38560 30457
rect 38480 30400 38560 30423
rect 38640 32377 38720 32400
rect 38640 32343 38663 32377
rect 38697 32343 38720 32377
rect 38640 32057 38720 32343
rect 38640 32023 38663 32057
rect 38697 32023 38720 32057
rect 38640 31737 38720 32023
rect 38640 31703 38663 31737
rect 38697 31703 38720 31737
rect 38640 31417 38720 31703
rect 38640 31383 38663 31417
rect 38697 31383 38720 31417
rect 38640 31097 38720 31383
rect 38640 31063 38663 31097
rect 38697 31063 38720 31097
rect 38640 30777 38720 31063
rect 38640 30743 38663 30777
rect 38697 30743 38720 30777
rect 38640 30457 38720 30743
rect 38640 30423 38663 30457
rect 38697 30423 38720 30457
rect 38640 30400 38720 30423
rect 38800 32377 38880 32400
rect 38800 32343 38823 32377
rect 38857 32343 38880 32377
rect 38800 32057 38880 32343
rect 38800 32023 38823 32057
rect 38857 32023 38880 32057
rect 38800 31737 38880 32023
rect 38800 31703 38823 31737
rect 38857 31703 38880 31737
rect 38800 31417 38880 31703
rect 38800 31383 38823 31417
rect 38857 31383 38880 31417
rect 38800 31097 38880 31383
rect 38800 31063 38823 31097
rect 38857 31063 38880 31097
rect 38800 30777 38880 31063
rect 38800 30743 38823 30777
rect 38857 30743 38880 30777
rect 38800 30457 38880 30743
rect 38800 30423 38823 30457
rect 38857 30423 38880 30457
rect 38800 30400 38880 30423
rect 38960 32377 39040 32400
rect 38960 32343 38983 32377
rect 39017 32343 39040 32377
rect 38960 32057 39040 32343
rect 38960 32023 38983 32057
rect 39017 32023 39040 32057
rect 38960 31737 39040 32023
rect 38960 31703 38983 31737
rect 39017 31703 39040 31737
rect 38960 31417 39040 31703
rect 38960 31383 38983 31417
rect 39017 31383 39040 31417
rect 38960 31097 39040 31383
rect 38960 31063 38983 31097
rect 39017 31063 39040 31097
rect 38960 30777 39040 31063
rect 38960 30743 38983 30777
rect 39017 30743 39040 30777
rect 38960 30457 39040 30743
rect 38960 30423 38983 30457
rect 39017 30423 39040 30457
rect 38960 30400 39040 30423
rect 39120 32377 39200 32400
rect 39120 32343 39143 32377
rect 39177 32343 39200 32377
rect 39120 32057 39200 32343
rect 39120 32023 39143 32057
rect 39177 32023 39200 32057
rect 39120 31737 39200 32023
rect 39120 31703 39143 31737
rect 39177 31703 39200 31737
rect 39120 31417 39200 31703
rect 39120 31383 39143 31417
rect 39177 31383 39200 31417
rect 39120 31097 39200 31383
rect 39120 31063 39143 31097
rect 39177 31063 39200 31097
rect 39120 30777 39200 31063
rect 39120 30743 39143 30777
rect 39177 30743 39200 30777
rect 39120 30457 39200 30743
rect 39120 30423 39143 30457
rect 39177 30423 39200 30457
rect 39120 30400 39200 30423
rect 39280 32377 39360 32400
rect 39280 32343 39303 32377
rect 39337 32343 39360 32377
rect 39280 32057 39360 32343
rect 39280 32023 39303 32057
rect 39337 32023 39360 32057
rect 39280 31737 39360 32023
rect 39280 31703 39303 31737
rect 39337 31703 39360 31737
rect 39280 31417 39360 31703
rect 39280 31383 39303 31417
rect 39337 31383 39360 31417
rect 39280 31097 39360 31383
rect 39280 31063 39303 31097
rect 39337 31063 39360 31097
rect 39280 30777 39360 31063
rect 39280 30743 39303 30777
rect 39337 30743 39360 30777
rect 39280 30457 39360 30743
rect 39280 30423 39303 30457
rect 39337 30423 39360 30457
rect 39280 30400 39360 30423
rect 39440 32377 39520 32400
rect 39440 32343 39463 32377
rect 39497 32343 39520 32377
rect 39440 32057 39520 32343
rect 39440 32023 39463 32057
rect 39497 32023 39520 32057
rect 39440 31737 39520 32023
rect 39440 31703 39463 31737
rect 39497 31703 39520 31737
rect 39440 31417 39520 31703
rect 39440 31383 39463 31417
rect 39497 31383 39520 31417
rect 39440 31097 39520 31383
rect 39440 31063 39463 31097
rect 39497 31063 39520 31097
rect 39440 30777 39520 31063
rect 39440 30743 39463 30777
rect 39497 30743 39520 30777
rect 39440 30457 39520 30743
rect 39440 30423 39463 30457
rect 39497 30423 39520 30457
rect 39440 30400 39520 30423
rect 39600 32377 39680 32400
rect 39600 32343 39623 32377
rect 39657 32343 39680 32377
rect 39600 32057 39680 32343
rect 39600 32023 39623 32057
rect 39657 32023 39680 32057
rect 39600 31737 39680 32023
rect 39600 31703 39623 31737
rect 39657 31703 39680 31737
rect 39600 31417 39680 31703
rect 39600 31383 39623 31417
rect 39657 31383 39680 31417
rect 39600 31097 39680 31383
rect 39600 31063 39623 31097
rect 39657 31063 39680 31097
rect 39600 30777 39680 31063
rect 39600 30743 39623 30777
rect 39657 30743 39680 30777
rect 39600 30457 39680 30743
rect 39600 30423 39623 30457
rect 39657 30423 39680 30457
rect 39600 30400 39680 30423
rect 39760 32377 39840 32400
rect 39760 32343 39783 32377
rect 39817 32343 39840 32377
rect 39760 32057 39840 32343
rect 39760 32023 39783 32057
rect 39817 32023 39840 32057
rect 39760 31737 39840 32023
rect 39760 31703 39783 31737
rect 39817 31703 39840 31737
rect 39760 31417 39840 31703
rect 39760 31383 39783 31417
rect 39817 31383 39840 31417
rect 39760 31097 39840 31383
rect 39760 31063 39783 31097
rect 39817 31063 39840 31097
rect 39760 30777 39840 31063
rect 39760 30743 39783 30777
rect 39817 30743 39840 30777
rect 39760 30457 39840 30743
rect 39760 30423 39783 30457
rect 39817 30423 39840 30457
rect 39760 30400 39840 30423
rect 39920 32377 40000 32400
rect 39920 32343 39943 32377
rect 39977 32343 40000 32377
rect 39920 32057 40000 32343
rect 39920 32023 39943 32057
rect 39977 32023 40000 32057
rect 39920 31737 40000 32023
rect 39920 31703 39943 31737
rect 39977 31703 40000 31737
rect 39920 31417 40000 31703
rect 39920 31383 39943 31417
rect 39977 31383 40000 31417
rect 39920 31097 40000 31383
rect 39920 31063 39943 31097
rect 39977 31063 40000 31097
rect 39920 30777 40000 31063
rect 39920 30743 39943 30777
rect 39977 30743 40000 30777
rect 39920 30457 40000 30743
rect 39920 30423 39943 30457
rect 39977 30423 40000 30457
rect 39920 30400 40000 30423
rect 40080 32377 40160 32400
rect 40080 32343 40103 32377
rect 40137 32343 40160 32377
rect 40080 32057 40160 32343
rect 40080 32023 40103 32057
rect 40137 32023 40160 32057
rect 40080 31737 40160 32023
rect 40080 31703 40103 31737
rect 40137 31703 40160 31737
rect 40080 31417 40160 31703
rect 40080 31383 40103 31417
rect 40137 31383 40160 31417
rect 40080 31097 40160 31383
rect 40080 31063 40103 31097
rect 40137 31063 40160 31097
rect 40080 30777 40160 31063
rect 40080 30743 40103 30777
rect 40137 30743 40160 30777
rect 40080 30457 40160 30743
rect 40080 30423 40103 30457
rect 40137 30423 40160 30457
rect 40080 30400 40160 30423
rect 40240 32377 40320 32400
rect 40240 32343 40263 32377
rect 40297 32343 40320 32377
rect 40240 32057 40320 32343
rect 40240 32023 40263 32057
rect 40297 32023 40320 32057
rect 40240 31737 40320 32023
rect 40240 31703 40263 31737
rect 40297 31703 40320 31737
rect 40240 31417 40320 31703
rect 40240 31383 40263 31417
rect 40297 31383 40320 31417
rect 40240 31097 40320 31383
rect 40240 31063 40263 31097
rect 40297 31063 40320 31097
rect 40240 30777 40320 31063
rect 40240 30743 40263 30777
rect 40297 30743 40320 30777
rect 40240 30457 40320 30743
rect 40240 30423 40263 30457
rect 40297 30423 40320 30457
rect 40240 30400 40320 30423
rect 40400 32377 40480 32400
rect 40400 32343 40423 32377
rect 40457 32343 40480 32377
rect 40400 32057 40480 32343
rect 40400 32023 40423 32057
rect 40457 32023 40480 32057
rect 40400 31737 40480 32023
rect 40400 31703 40423 31737
rect 40457 31703 40480 31737
rect 40400 31417 40480 31703
rect 40400 31383 40423 31417
rect 40457 31383 40480 31417
rect 40400 31097 40480 31383
rect 40400 31063 40423 31097
rect 40457 31063 40480 31097
rect 40400 30777 40480 31063
rect 40400 30743 40423 30777
rect 40457 30743 40480 30777
rect 40400 30457 40480 30743
rect 40400 30423 40423 30457
rect 40457 30423 40480 30457
rect 40400 30400 40480 30423
rect 40560 32377 40640 32400
rect 40560 32343 40583 32377
rect 40617 32343 40640 32377
rect 40560 32057 40640 32343
rect 40560 32023 40583 32057
rect 40617 32023 40640 32057
rect 40560 31737 40640 32023
rect 40560 31703 40583 31737
rect 40617 31703 40640 31737
rect 40560 31417 40640 31703
rect 40560 31383 40583 31417
rect 40617 31383 40640 31417
rect 40560 31097 40640 31383
rect 40560 31063 40583 31097
rect 40617 31063 40640 31097
rect 40560 30777 40640 31063
rect 40560 30743 40583 30777
rect 40617 30743 40640 30777
rect 40560 30457 40640 30743
rect 40560 30423 40583 30457
rect 40617 30423 40640 30457
rect 40560 30400 40640 30423
rect 40720 32377 40800 32400
rect 40720 32343 40743 32377
rect 40777 32343 40800 32377
rect 40720 32057 40800 32343
rect 40720 32023 40743 32057
rect 40777 32023 40800 32057
rect 40720 31737 40800 32023
rect 40720 31703 40743 31737
rect 40777 31703 40800 31737
rect 40720 31417 40800 31703
rect 40720 31383 40743 31417
rect 40777 31383 40800 31417
rect 40720 31097 40800 31383
rect 40720 31063 40743 31097
rect 40777 31063 40800 31097
rect 40720 30777 40800 31063
rect 40720 30743 40743 30777
rect 40777 30743 40800 30777
rect 40720 30457 40800 30743
rect 40720 30423 40743 30457
rect 40777 30423 40800 30457
rect 40720 30400 40800 30423
rect 40880 32377 40960 32400
rect 40880 32343 40903 32377
rect 40937 32343 40960 32377
rect 40880 32057 40960 32343
rect 40880 32023 40903 32057
rect 40937 32023 40960 32057
rect 40880 31737 40960 32023
rect 40880 31703 40903 31737
rect 40937 31703 40960 31737
rect 40880 31417 40960 31703
rect 40880 31383 40903 31417
rect 40937 31383 40960 31417
rect 40880 31097 40960 31383
rect 40880 31063 40903 31097
rect 40937 31063 40960 31097
rect 40880 30777 40960 31063
rect 40880 30743 40903 30777
rect 40937 30743 40960 30777
rect 40880 30457 40960 30743
rect 40880 30423 40903 30457
rect 40937 30423 40960 30457
rect 40880 30400 40960 30423
rect 41040 32377 41120 32400
rect 41040 32343 41063 32377
rect 41097 32343 41120 32377
rect 41040 32057 41120 32343
rect 41040 32023 41063 32057
rect 41097 32023 41120 32057
rect 41040 31737 41120 32023
rect 41040 31703 41063 31737
rect 41097 31703 41120 31737
rect 41040 31417 41120 31703
rect 41040 31383 41063 31417
rect 41097 31383 41120 31417
rect 41040 31097 41120 31383
rect 41040 31063 41063 31097
rect 41097 31063 41120 31097
rect 41040 30777 41120 31063
rect 41040 30743 41063 30777
rect 41097 30743 41120 30777
rect 41040 30457 41120 30743
rect 41040 30423 41063 30457
rect 41097 30423 41120 30457
rect 41040 30400 41120 30423
rect 41200 32377 41280 32400
rect 41200 32343 41223 32377
rect 41257 32343 41280 32377
rect 41200 32057 41280 32343
rect 41200 32023 41223 32057
rect 41257 32023 41280 32057
rect 41200 31737 41280 32023
rect 41200 31703 41223 31737
rect 41257 31703 41280 31737
rect 41200 31417 41280 31703
rect 41200 31383 41223 31417
rect 41257 31383 41280 31417
rect 41200 31097 41280 31383
rect 41200 31063 41223 31097
rect 41257 31063 41280 31097
rect 41200 30777 41280 31063
rect 41200 30743 41223 30777
rect 41257 30743 41280 30777
rect 41200 30457 41280 30743
rect 41200 30423 41223 30457
rect 41257 30423 41280 30457
rect 41200 30400 41280 30423
rect 41360 32377 41440 32400
rect 41360 32343 41383 32377
rect 41417 32343 41440 32377
rect 41360 32057 41440 32343
rect 41360 32023 41383 32057
rect 41417 32023 41440 32057
rect 41360 31737 41440 32023
rect 41360 31703 41383 31737
rect 41417 31703 41440 31737
rect 41360 31417 41440 31703
rect 41360 31383 41383 31417
rect 41417 31383 41440 31417
rect 41360 31097 41440 31383
rect 41360 31063 41383 31097
rect 41417 31063 41440 31097
rect 41360 30777 41440 31063
rect 41360 30743 41383 30777
rect 41417 30743 41440 30777
rect 41360 30457 41440 30743
rect 41360 30423 41383 30457
rect 41417 30423 41440 30457
rect 41360 30400 41440 30423
rect 41520 32377 41600 32400
rect 41520 32343 41543 32377
rect 41577 32343 41600 32377
rect 41520 32057 41600 32343
rect 41520 32023 41543 32057
rect 41577 32023 41600 32057
rect 41520 31737 41600 32023
rect 41520 31703 41543 31737
rect 41577 31703 41600 31737
rect 41520 31417 41600 31703
rect 41520 31383 41543 31417
rect 41577 31383 41600 31417
rect 41520 31097 41600 31383
rect 41520 31063 41543 31097
rect 41577 31063 41600 31097
rect 41520 30777 41600 31063
rect 41520 30743 41543 30777
rect 41577 30743 41600 30777
rect 41520 30457 41600 30743
rect 41520 30423 41543 30457
rect 41577 30423 41600 30457
rect 41520 30400 41600 30423
rect 41680 32377 41760 32400
rect 41680 32343 41703 32377
rect 41737 32343 41760 32377
rect 41680 32057 41760 32343
rect 41680 32023 41703 32057
rect 41737 32023 41760 32057
rect 41680 31737 41760 32023
rect 41680 31703 41703 31737
rect 41737 31703 41760 31737
rect 41680 31417 41760 31703
rect 41680 31383 41703 31417
rect 41737 31383 41760 31417
rect 41680 31097 41760 31383
rect 41680 31063 41703 31097
rect 41737 31063 41760 31097
rect 41680 30777 41760 31063
rect 41680 30743 41703 30777
rect 41737 30743 41760 30777
rect 41680 30457 41760 30743
rect 41680 30423 41703 30457
rect 41737 30423 41760 30457
rect 41680 30400 41760 30423
rect 41840 32377 41920 32400
rect 41840 32343 41863 32377
rect 41897 32343 41920 32377
rect 41840 32057 41920 32343
rect 41840 32023 41863 32057
rect 41897 32023 41920 32057
rect 41840 31737 41920 32023
rect 41840 31703 41863 31737
rect 41897 31703 41920 31737
rect 41840 31417 41920 31703
rect 41840 31383 41863 31417
rect 41897 31383 41920 31417
rect 41840 31097 41920 31383
rect 41840 31063 41863 31097
rect 41897 31063 41920 31097
rect 41840 30777 41920 31063
rect 41840 30743 41863 30777
rect 41897 30743 41920 30777
rect 41840 30457 41920 30743
rect 41840 30423 41863 30457
rect 41897 30423 41920 30457
rect 41840 30400 41920 30423
rect 0 30297 80 30320
rect 0 30263 23 30297
rect 57 30263 80 30297
rect 0 29977 80 30263
rect 0 29943 23 29977
rect 57 29943 80 29977
rect 0 29920 80 29943
rect 160 30297 240 30320
rect 160 30263 183 30297
rect 217 30263 240 30297
rect 160 29977 240 30263
rect 160 29943 183 29977
rect 217 29943 240 29977
rect 160 29920 240 29943
rect 320 30297 400 30320
rect 320 30263 343 30297
rect 377 30263 400 30297
rect 320 29977 400 30263
rect 320 29943 343 29977
rect 377 29943 400 29977
rect 320 29920 400 29943
rect 480 30297 560 30320
rect 480 30263 503 30297
rect 537 30263 560 30297
rect 480 29977 560 30263
rect 480 29943 503 29977
rect 537 29943 560 29977
rect 480 29920 560 29943
rect 640 30297 720 30320
rect 640 30263 663 30297
rect 697 30263 720 30297
rect 640 29977 720 30263
rect 640 29943 663 29977
rect 697 29943 720 29977
rect 640 29920 720 29943
rect 800 30297 880 30320
rect 800 30263 823 30297
rect 857 30263 880 30297
rect 800 29977 880 30263
rect 800 29943 823 29977
rect 857 29943 880 29977
rect 800 29920 880 29943
rect 960 30297 1040 30320
rect 960 30263 983 30297
rect 1017 30263 1040 30297
rect 960 29977 1040 30263
rect 960 29943 983 29977
rect 1017 29943 1040 29977
rect 960 29920 1040 29943
rect 1120 30297 1200 30320
rect 1120 30263 1143 30297
rect 1177 30263 1200 30297
rect 1120 29977 1200 30263
rect 1120 29943 1143 29977
rect 1177 29943 1200 29977
rect 1120 29920 1200 29943
rect 1280 30297 1360 30320
rect 1280 30263 1303 30297
rect 1337 30263 1360 30297
rect 1280 29977 1360 30263
rect 1280 29943 1303 29977
rect 1337 29943 1360 29977
rect 1280 29920 1360 29943
rect 1440 30297 1520 30320
rect 1440 30263 1463 30297
rect 1497 30263 1520 30297
rect 1440 29977 1520 30263
rect 1440 29943 1463 29977
rect 1497 29943 1520 29977
rect 1440 29920 1520 29943
rect 1600 30297 1680 30320
rect 1600 30263 1623 30297
rect 1657 30263 1680 30297
rect 1600 29977 1680 30263
rect 1600 29943 1623 29977
rect 1657 29943 1680 29977
rect 1600 29920 1680 29943
rect 1760 30297 1840 30320
rect 1760 30263 1783 30297
rect 1817 30263 1840 30297
rect 1760 29977 1840 30263
rect 1760 29943 1783 29977
rect 1817 29943 1840 29977
rect 1760 29920 1840 29943
rect 1920 30297 2000 30320
rect 1920 30263 1943 30297
rect 1977 30263 2000 30297
rect 1920 29977 2000 30263
rect 1920 29943 1943 29977
rect 1977 29943 2000 29977
rect 1920 29920 2000 29943
rect 2080 30297 2160 30320
rect 2080 30263 2103 30297
rect 2137 30263 2160 30297
rect 2080 29977 2160 30263
rect 2080 29943 2103 29977
rect 2137 29943 2160 29977
rect 2080 29920 2160 29943
rect 2240 30297 2320 30320
rect 2240 30263 2263 30297
rect 2297 30263 2320 30297
rect 2240 29977 2320 30263
rect 2240 29943 2263 29977
rect 2297 29943 2320 29977
rect 2240 29920 2320 29943
rect 2400 30297 2480 30320
rect 2400 30263 2423 30297
rect 2457 30263 2480 30297
rect 2400 29977 2480 30263
rect 2400 29943 2423 29977
rect 2457 29943 2480 29977
rect 2400 29920 2480 29943
rect 2560 30297 2640 30320
rect 2560 30263 2583 30297
rect 2617 30263 2640 30297
rect 2560 29977 2640 30263
rect 2560 29943 2583 29977
rect 2617 29943 2640 29977
rect 2560 29920 2640 29943
rect 2720 30297 2800 30320
rect 2720 30263 2743 30297
rect 2777 30263 2800 30297
rect 2720 29977 2800 30263
rect 2720 29943 2743 29977
rect 2777 29943 2800 29977
rect 2720 29920 2800 29943
rect 2880 30297 2960 30320
rect 2880 30263 2903 30297
rect 2937 30263 2960 30297
rect 2880 29977 2960 30263
rect 2880 29943 2903 29977
rect 2937 29943 2960 29977
rect 2880 29920 2960 29943
rect 3040 30297 3120 30320
rect 3040 30263 3063 30297
rect 3097 30263 3120 30297
rect 3040 29977 3120 30263
rect 3040 29943 3063 29977
rect 3097 29943 3120 29977
rect 3040 29920 3120 29943
rect 3200 30297 3280 30320
rect 3200 30263 3223 30297
rect 3257 30263 3280 30297
rect 3200 29977 3280 30263
rect 3200 29943 3223 29977
rect 3257 29943 3280 29977
rect 3200 29920 3280 29943
rect 3360 30297 3440 30320
rect 3360 30263 3383 30297
rect 3417 30263 3440 30297
rect 3360 29977 3440 30263
rect 3360 29943 3383 29977
rect 3417 29943 3440 29977
rect 3360 29920 3440 29943
rect 3520 30297 3600 30320
rect 3520 30263 3543 30297
rect 3577 30263 3600 30297
rect 3520 29977 3600 30263
rect 3520 29943 3543 29977
rect 3577 29943 3600 29977
rect 3520 29920 3600 29943
rect 3680 30297 3760 30320
rect 3680 30263 3703 30297
rect 3737 30263 3760 30297
rect 3680 29977 3760 30263
rect 3680 29943 3703 29977
rect 3737 29943 3760 29977
rect 3680 29920 3760 29943
rect 3840 30297 3920 30320
rect 3840 30263 3863 30297
rect 3897 30263 3920 30297
rect 3840 29977 3920 30263
rect 3840 29943 3863 29977
rect 3897 29943 3920 29977
rect 3840 29920 3920 29943
rect 4000 30297 4080 30320
rect 4000 30263 4023 30297
rect 4057 30263 4080 30297
rect 4000 29977 4080 30263
rect 4000 29943 4023 29977
rect 4057 29943 4080 29977
rect 4000 29920 4080 29943
rect 4160 30297 4240 30320
rect 4160 30263 4183 30297
rect 4217 30263 4240 30297
rect 4160 29977 4240 30263
rect 4160 29943 4183 29977
rect 4217 29943 4240 29977
rect 4160 29920 4240 29943
rect 4320 30297 4400 30320
rect 4320 30263 4343 30297
rect 4377 30263 4400 30297
rect 4320 29977 4400 30263
rect 4320 29943 4343 29977
rect 4377 29943 4400 29977
rect 4320 29920 4400 29943
rect 4480 30297 4560 30320
rect 4480 30263 4503 30297
rect 4537 30263 4560 30297
rect 4480 29977 4560 30263
rect 4480 29943 4503 29977
rect 4537 29943 4560 29977
rect 4480 29920 4560 29943
rect 4640 30297 4720 30320
rect 4640 30263 4663 30297
rect 4697 30263 4720 30297
rect 4640 29977 4720 30263
rect 4640 29943 4663 29977
rect 4697 29943 4720 29977
rect 4640 29920 4720 29943
rect 4800 30297 4880 30320
rect 4800 30263 4823 30297
rect 4857 30263 4880 30297
rect 4800 29977 4880 30263
rect 4800 29943 4823 29977
rect 4857 29943 4880 29977
rect 4800 29920 4880 29943
rect 4960 30297 5040 30320
rect 4960 30263 4983 30297
rect 5017 30263 5040 30297
rect 4960 29977 5040 30263
rect 4960 29943 4983 29977
rect 5017 29943 5040 29977
rect 4960 29920 5040 29943
rect 5120 30297 5200 30320
rect 5120 30263 5143 30297
rect 5177 30263 5200 30297
rect 5120 29977 5200 30263
rect 5120 29943 5143 29977
rect 5177 29943 5200 29977
rect 5120 29920 5200 29943
rect 5280 30297 5360 30320
rect 5280 30263 5303 30297
rect 5337 30263 5360 30297
rect 5280 29977 5360 30263
rect 5280 29943 5303 29977
rect 5337 29943 5360 29977
rect 5280 29920 5360 29943
rect 5440 30297 5520 30320
rect 5440 30263 5463 30297
rect 5497 30263 5520 30297
rect 5440 29977 5520 30263
rect 5440 29943 5463 29977
rect 5497 29943 5520 29977
rect 5440 29920 5520 29943
rect 5600 30297 5680 30320
rect 5600 30263 5623 30297
rect 5657 30263 5680 30297
rect 5600 29977 5680 30263
rect 5600 29943 5623 29977
rect 5657 29943 5680 29977
rect 5600 29920 5680 29943
rect 5760 30297 5840 30320
rect 5760 30263 5783 30297
rect 5817 30263 5840 30297
rect 5760 29977 5840 30263
rect 5760 29943 5783 29977
rect 5817 29943 5840 29977
rect 5760 29920 5840 29943
rect 5920 30297 6000 30320
rect 5920 30263 5943 30297
rect 5977 30263 6000 30297
rect 5920 29977 6000 30263
rect 5920 29943 5943 29977
rect 5977 29943 6000 29977
rect 5920 29920 6000 29943
rect 6080 30297 6160 30320
rect 6080 30263 6103 30297
rect 6137 30263 6160 30297
rect 6080 29977 6160 30263
rect 6080 29943 6103 29977
rect 6137 29943 6160 29977
rect 6080 29920 6160 29943
rect 6240 30297 6320 30320
rect 6240 30263 6263 30297
rect 6297 30263 6320 30297
rect 6240 29977 6320 30263
rect 6240 29943 6263 29977
rect 6297 29943 6320 29977
rect 6240 29920 6320 29943
rect 6400 30297 6480 30320
rect 6400 30263 6423 30297
rect 6457 30263 6480 30297
rect 6400 29977 6480 30263
rect 6400 29943 6423 29977
rect 6457 29943 6480 29977
rect 6400 29920 6480 29943
rect 6560 30297 6640 30320
rect 6560 30263 6583 30297
rect 6617 30263 6640 30297
rect 6560 29977 6640 30263
rect 6560 29943 6583 29977
rect 6617 29943 6640 29977
rect 6560 29920 6640 29943
rect 6720 30297 6800 30320
rect 6720 30263 6743 30297
rect 6777 30263 6800 30297
rect 6720 29977 6800 30263
rect 6720 29943 6743 29977
rect 6777 29943 6800 29977
rect 6720 29920 6800 29943
rect 6880 30297 6960 30320
rect 6880 30263 6903 30297
rect 6937 30263 6960 30297
rect 6880 29977 6960 30263
rect 6880 29943 6903 29977
rect 6937 29943 6960 29977
rect 6880 29920 6960 29943
rect 7040 30297 7120 30320
rect 7040 30263 7063 30297
rect 7097 30263 7120 30297
rect 7040 29977 7120 30263
rect 7040 29943 7063 29977
rect 7097 29943 7120 29977
rect 7040 29920 7120 29943
rect 7200 30297 7280 30320
rect 7200 30263 7223 30297
rect 7257 30263 7280 30297
rect 7200 29977 7280 30263
rect 7200 29943 7223 29977
rect 7257 29943 7280 29977
rect 7200 29920 7280 29943
rect 7360 30297 7440 30320
rect 7360 30263 7383 30297
rect 7417 30263 7440 30297
rect 7360 29977 7440 30263
rect 7360 29943 7383 29977
rect 7417 29943 7440 29977
rect 7360 29920 7440 29943
rect 7520 30297 7600 30320
rect 7520 30263 7543 30297
rect 7577 30263 7600 30297
rect 7520 29977 7600 30263
rect 7520 29943 7543 29977
rect 7577 29943 7600 29977
rect 7520 29920 7600 29943
rect 7680 30297 7760 30320
rect 7680 30263 7703 30297
rect 7737 30263 7760 30297
rect 7680 29977 7760 30263
rect 7680 29943 7703 29977
rect 7737 29943 7760 29977
rect 7680 29920 7760 29943
rect 7840 30297 7920 30320
rect 7840 30263 7863 30297
rect 7897 30263 7920 30297
rect 7840 29977 7920 30263
rect 7840 29943 7863 29977
rect 7897 29943 7920 29977
rect 7840 29920 7920 29943
rect 8000 30297 8080 30320
rect 8000 30263 8023 30297
rect 8057 30263 8080 30297
rect 8000 29977 8080 30263
rect 8000 29943 8023 29977
rect 8057 29943 8080 29977
rect 8000 29920 8080 29943
rect 8160 30297 8240 30320
rect 8160 30263 8183 30297
rect 8217 30263 8240 30297
rect 8160 29977 8240 30263
rect 8160 29943 8183 29977
rect 8217 29943 8240 29977
rect 8160 29920 8240 29943
rect 8320 30297 8400 30320
rect 8320 30263 8343 30297
rect 8377 30263 8400 30297
rect 8320 29977 8400 30263
rect 8320 29943 8343 29977
rect 8377 29943 8400 29977
rect 8320 29920 8400 29943
rect 8480 29920 8560 30320
rect 8640 29920 8720 30320
rect 8800 29920 8880 30320
rect 8960 29920 9040 30320
rect 9120 29920 9200 30320
rect 9280 29920 9360 30320
rect 9440 29920 9520 30320
rect 9600 29920 9680 30320
rect 9760 29920 9840 30320
rect 9920 29920 10000 30320
rect 10080 29920 10160 30320
rect 10240 29920 10320 30320
rect 10400 29920 10480 30320
rect 10560 29920 10640 30320
rect 10720 29920 10800 30320
rect 10880 29920 10960 30320
rect 11040 29920 11120 30320
rect 11200 29920 11280 30320
rect 11360 29920 11440 30320
rect 11520 29920 11600 30320
rect 11680 29920 11760 30320
rect 11840 29920 11920 30320
rect 12000 29920 12080 30320
rect 12160 29920 12240 30320
rect 12320 29920 12400 30320
rect 12480 30297 12560 30320
rect 12480 30263 12503 30297
rect 12537 30263 12560 30297
rect 12480 29977 12560 30263
rect 12480 29943 12503 29977
rect 12537 29943 12560 29977
rect 12480 29920 12560 29943
rect 12640 30297 12720 30320
rect 12640 30263 12663 30297
rect 12697 30263 12720 30297
rect 12640 29977 12720 30263
rect 12640 29943 12663 29977
rect 12697 29943 12720 29977
rect 12640 29920 12720 29943
rect 12800 30297 12880 30320
rect 12800 30263 12823 30297
rect 12857 30263 12880 30297
rect 12800 29977 12880 30263
rect 12800 29943 12823 29977
rect 12857 29943 12880 29977
rect 12800 29920 12880 29943
rect 12960 30297 13040 30320
rect 12960 30263 12983 30297
rect 13017 30263 13040 30297
rect 12960 29977 13040 30263
rect 12960 29943 12983 29977
rect 13017 29943 13040 29977
rect 12960 29920 13040 29943
rect 13120 30297 13200 30320
rect 13120 30263 13143 30297
rect 13177 30263 13200 30297
rect 13120 29977 13200 30263
rect 13120 29943 13143 29977
rect 13177 29943 13200 29977
rect 13120 29920 13200 29943
rect 13280 30297 13360 30320
rect 13280 30263 13303 30297
rect 13337 30263 13360 30297
rect 13280 29977 13360 30263
rect 13280 29943 13303 29977
rect 13337 29943 13360 29977
rect 13280 29920 13360 29943
rect 13440 30297 13520 30320
rect 13440 30263 13463 30297
rect 13497 30263 13520 30297
rect 13440 29977 13520 30263
rect 13440 29943 13463 29977
rect 13497 29943 13520 29977
rect 13440 29920 13520 29943
rect 13600 30297 13680 30320
rect 13600 30263 13623 30297
rect 13657 30263 13680 30297
rect 13600 29977 13680 30263
rect 13600 29943 13623 29977
rect 13657 29943 13680 29977
rect 13600 29920 13680 29943
rect 13760 30297 13840 30320
rect 13760 30263 13783 30297
rect 13817 30263 13840 30297
rect 13760 29977 13840 30263
rect 13760 29943 13783 29977
rect 13817 29943 13840 29977
rect 13760 29920 13840 29943
rect 13920 30297 14000 30320
rect 13920 30263 13943 30297
rect 13977 30263 14000 30297
rect 13920 29977 14000 30263
rect 13920 29943 13943 29977
rect 13977 29943 14000 29977
rect 13920 29920 14000 29943
rect 14080 30297 14160 30320
rect 14080 30263 14103 30297
rect 14137 30263 14160 30297
rect 14080 29977 14160 30263
rect 14080 29943 14103 29977
rect 14137 29943 14160 29977
rect 14080 29920 14160 29943
rect 14240 30297 14320 30320
rect 14240 30263 14263 30297
rect 14297 30263 14320 30297
rect 14240 29977 14320 30263
rect 14240 29943 14263 29977
rect 14297 29943 14320 29977
rect 14240 29920 14320 29943
rect 14400 30297 14480 30320
rect 14400 30263 14423 30297
rect 14457 30263 14480 30297
rect 14400 29977 14480 30263
rect 14400 29943 14423 29977
rect 14457 29943 14480 29977
rect 14400 29920 14480 29943
rect 14560 30297 14640 30320
rect 14560 30263 14583 30297
rect 14617 30263 14640 30297
rect 14560 29977 14640 30263
rect 14560 29943 14583 29977
rect 14617 29943 14640 29977
rect 14560 29920 14640 29943
rect 14720 30297 14800 30320
rect 14720 30263 14743 30297
rect 14777 30263 14800 30297
rect 14720 29977 14800 30263
rect 14720 29943 14743 29977
rect 14777 29943 14800 29977
rect 14720 29920 14800 29943
rect 14880 30297 14960 30320
rect 14880 30263 14903 30297
rect 14937 30263 14960 30297
rect 14880 29977 14960 30263
rect 14880 29943 14903 29977
rect 14937 29943 14960 29977
rect 14880 29920 14960 29943
rect 15040 30297 15120 30320
rect 15040 30263 15063 30297
rect 15097 30263 15120 30297
rect 15040 29977 15120 30263
rect 15040 29943 15063 29977
rect 15097 29943 15120 29977
rect 15040 29920 15120 29943
rect 15200 30297 15280 30320
rect 15200 30263 15223 30297
rect 15257 30263 15280 30297
rect 15200 29977 15280 30263
rect 15200 29943 15223 29977
rect 15257 29943 15280 29977
rect 15200 29920 15280 29943
rect 15360 30297 15440 30320
rect 15360 30263 15383 30297
rect 15417 30263 15440 30297
rect 15360 29977 15440 30263
rect 15360 29943 15383 29977
rect 15417 29943 15440 29977
rect 15360 29920 15440 29943
rect 15520 30297 15600 30320
rect 15520 30263 15543 30297
rect 15577 30263 15600 30297
rect 15520 29977 15600 30263
rect 15520 29943 15543 29977
rect 15577 29943 15600 29977
rect 15520 29920 15600 29943
rect 15680 30297 15760 30320
rect 15680 30263 15703 30297
rect 15737 30263 15760 30297
rect 15680 29977 15760 30263
rect 15680 29943 15703 29977
rect 15737 29943 15760 29977
rect 15680 29920 15760 29943
rect 15840 30297 15920 30320
rect 15840 30263 15863 30297
rect 15897 30263 15920 30297
rect 15840 29977 15920 30263
rect 15840 29943 15863 29977
rect 15897 29943 15920 29977
rect 15840 29920 15920 29943
rect 16000 30297 16080 30320
rect 16000 30263 16023 30297
rect 16057 30263 16080 30297
rect 16000 29977 16080 30263
rect 16000 29943 16023 29977
rect 16057 29943 16080 29977
rect 16000 29920 16080 29943
rect 16160 30297 16240 30320
rect 16160 30263 16183 30297
rect 16217 30263 16240 30297
rect 16160 29977 16240 30263
rect 16160 29943 16183 29977
rect 16217 29943 16240 29977
rect 16160 29920 16240 29943
rect 16320 30297 16400 30320
rect 16320 30263 16343 30297
rect 16377 30263 16400 30297
rect 16320 29977 16400 30263
rect 16320 29943 16343 29977
rect 16377 29943 16400 29977
rect 16320 29920 16400 29943
rect 16480 30297 16560 30320
rect 16480 30263 16503 30297
rect 16537 30263 16560 30297
rect 16480 29977 16560 30263
rect 16480 29943 16503 29977
rect 16537 29943 16560 29977
rect 16480 29920 16560 29943
rect 16640 30297 16720 30320
rect 16640 30263 16663 30297
rect 16697 30263 16720 30297
rect 16640 29977 16720 30263
rect 16640 29943 16663 29977
rect 16697 29943 16720 29977
rect 16640 29920 16720 29943
rect 16800 30297 16880 30320
rect 16800 30263 16823 30297
rect 16857 30263 16880 30297
rect 16800 29977 16880 30263
rect 16800 29943 16823 29977
rect 16857 29943 16880 29977
rect 16800 29920 16880 29943
rect 16960 30297 17040 30320
rect 16960 30263 16983 30297
rect 17017 30263 17040 30297
rect 16960 29977 17040 30263
rect 16960 29943 16983 29977
rect 17017 29943 17040 29977
rect 16960 29920 17040 29943
rect 17120 30297 17200 30320
rect 17120 30263 17143 30297
rect 17177 30263 17200 30297
rect 17120 29977 17200 30263
rect 17120 29943 17143 29977
rect 17177 29943 17200 29977
rect 17120 29920 17200 29943
rect 17280 30297 17360 30320
rect 17280 30263 17303 30297
rect 17337 30263 17360 30297
rect 17280 29977 17360 30263
rect 17280 29943 17303 29977
rect 17337 29943 17360 29977
rect 17280 29920 17360 29943
rect 17440 30297 17520 30320
rect 17440 30263 17463 30297
rect 17497 30263 17520 30297
rect 17440 29977 17520 30263
rect 17440 29943 17463 29977
rect 17497 29943 17520 29977
rect 17440 29920 17520 29943
rect 17600 30297 17680 30320
rect 17600 30263 17623 30297
rect 17657 30263 17680 30297
rect 17600 29977 17680 30263
rect 17600 29943 17623 29977
rect 17657 29943 17680 29977
rect 17600 29920 17680 29943
rect 17760 30297 17840 30320
rect 17760 30263 17783 30297
rect 17817 30263 17840 30297
rect 17760 29977 17840 30263
rect 17760 29943 17783 29977
rect 17817 29943 17840 29977
rect 17760 29920 17840 29943
rect 17920 30297 18000 30320
rect 17920 30263 17943 30297
rect 17977 30263 18000 30297
rect 17920 29977 18000 30263
rect 17920 29943 17943 29977
rect 17977 29943 18000 29977
rect 17920 29920 18000 29943
rect 18080 30297 18160 30320
rect 18080 30263 18103 30297
rect 18137 30263 18160 30297
rect 18080 29977 18160 30263
rect 18080 29943 18103 29977
rect 18137 29943 18160 29977
rect 18080 29920 18160 29943
rect 18240 30297 18320 30320
rect 18240 30263 18263 30297
rect 18297 30263 18320 30297
rect 18240 29977 18320 30263
rect 18240 29943 18263 29977
rect 18297 29943 18320 29977
rect 18240 29920 18320 29943
rect 18400 30297 18480 30320
rect 18400 30263 18423 30297
rect 18457 30263 18480 30297
rect 18400 29977 18480 30263
rect 18400 29943 18423 29977
rect 18457 29943 18480 29977
rect 18400 29920 18480 29943
rect 18560 30297 18640 30320
rect 18560 30263 18583 30297
rect 18617 30263 18640 30297
rect 18560 29977 18640 30263
rect 18560 29943 18583 29977
rect 18617 29943 18640 29977
rect 18560 29920 18640 29943
rect 18720 30297 18800 30320
rect 18720 30263 18743 30297
rect 18777 30263 18800 30297
rect 18720 29977 18800 30263
rect 18720 29943 18743 29977
rect 18777 29943 18800 29977
rect 18720 29920 18800 29943
rect 18880 30297 18960 30320
rect 18880 30263 18903 30297
rect 18937 30263 18960 30297
rect 18880 29977 18960 30263
rect 18880 29943 18903 29977
rect 18937 29943 18960 29977
rect 18880 29920 18960 29943
rect 19040 29920 19120 30320
rect 19200 29920 19280 30320
rect 19360 29920 19440 30320
rect 19520 29920 19600 30320
rect 19680 29920 19760 30320
rect 19840 29920 19920 30320
rect 20000 29920 20080 30320
rect 20160 29920 20240 30320
rect 20320 29920 20400 30320
rect 20480 29920 20560 30320
rect 20640 29920 20720 30320
rect 20800 29920 20880 30320
rect 20960 29920 21040 30320
rect 21120 29920 21200 30320
rect 21280 29920 21360 30320
rect 21440 29920 21520 30320
rect 21600 29920 21680 30320
rect 21760 29920 21840 30320
rect 21920 29920 22000 30320
rect 22080 29920 22160 30320
rect 22240 29920 22320 30320
rect 22400 29920 22480 30320
rect 22560 29920 22640 30320
rect 22720 29920 22800 30320
rect 22880 29920 22960 30320
rect 23120 30297 23200 30320
rect 23120 30263 23143 30297
rect 23177 30263 23200 30297
rect 23120 29977 23200 30263
rect 23120 29943 23143 29977
rect 23177 29943 23200 29977
rect 23120 29920 23200 29943
rect 23280 30297 23360 30320
rect 23280 30263 23303 30297
rect 23337 30263 23360 30297
rect 23280 29977 23360 30263
rect 23280 29943 23303 29977
rect 23337 29943 23360 29977
rect 23280 29920 23360 29943
rect 23440 30297 23520 30320
rect 23440 30263 23463 30297
rect 23497 30263 23520 30297
rect 23440 29977 23520 30263
rect 23440 29943 23463 29977
rect 23497 29943 23520 29977
rect 23440 29920 23520 29943
rect 23600 30297 23680 30320
rect 23600 30263 23623 30297
rect 23657 30263 23680 30297
rect 23600 29977 23680 30263
rect 23600 29943 23623 29977
rect 23657 29943 23680 29977
rect 23600 29920 23680 29943
rect 23760 30297 23840 30320
rect 23760 30263 23783 30297
rect 23817 30263 23840 30297
rect 23760 29977 23840 30263
rect 23760 29943 23783 29977
rect 23817 29943 23840 29977
rect 23760 29920 23840 29943
rect 23920 30297 24000 30320
rect 23920 30263 23943 30297
rect 23977 30263 24000 30297
rect 23920 29977 24000 30263
rect 23920 29943 23943 29977
rect 23977 29943 24000 29977
rect 23920 29920 24000 29943
rect 24080 30297 24160 30320
rect 24080 30263 24103 30297
rect 24137 30263 24160 30297
rect 24080 29977 24160 30263
rect 24080 29943 24103 29977
rect 24137 29943 24160 29977
rect 24080 29920 24160 29943
rect 24240 30297 24320 30320
rect 24240 30263 24263 30297
rect 24297 30263 24320 30297
rect 24240 29977 24320 30263
rect 24240 29943 24263 29977
rect 24297 29943 24320 29977
rect 24240 29920 24320 29943
rect 24400 30297 24480 30320
rect 24400 30263 24423 30297
rect 24457 30263 24480 30297
rect 24400 29977 24480 30263
rect 24400 29943 24423 29977
rect 24457 29943 24480 29977
rect 24400 29920 24480 29943
rect 24560 30297 24640 30320
rect 24560 30263 24583 30297
rect 24617 30263 24640 30297
rect 24560 29977 24640 30263
rect 24560 29943 24583 29977
rect 24617 29943 24640 29977
rect 24560 29920 24640 29943
rect 24720 30297 24800 30320
rect 24720 30263 24743 30297
rect 24777 30263 24800 30297
rect 24720 29977 24800 30263
rect 24720 29943 24743 29977
rect 24777 29943 24800 29977
rect 24720 29920 24800 29943
rect 24880 30297 24960 30320
rect 24880 30263 24903 30297
rect 24937 30263 24960 30297
rect 24880 29977 24960 30263
rect 24880 29943 24903 29977
rect 24937 29943 24960 29977
rect 24880 29920 24960 29943
rect 25040 30297 25120 30320
rect 25040 30263 25063 30297
rect 25097 30263 25120 30297
rect 25040 29977 25120 30263
rect 25040 29943 25063 29977
rect 25097 29943 25120 29977
rect 25040 29920 25120 29943
rect 25200 30297 25280 30320
rect 25200 30263 25223 30297
rect 25257 30263 25280 30297
rect 25200 29977 25280 30263
rect 25200 29943 25223 29977
rect 25257 29943 25280 29977
rect 25200 29920 25280 29943
rect 25360 30297 25440 30320
rect 25360 30263 25383 30297
rect 25417 30263 25440 30297
rect 25360 29977 25440 30263
rect 25360 29943 25383 29977
rect 25417 29943 25440 29977
rect 25360 29920 25440 29943
rect 25520 30297 25600 30320
rect 25520 30263 25543 30297
rect 25577 30263 25600 30297
rect 25520 29977 25600 30263
rect 25520 29943 25543 29977
rect 25577 29943 25600 29977
rect 25520 29920 25600 29943
rect 25680 30297 25760 30320
rect 25680 30263 25703 30297
rect 25737 30263 25760 30297
rect 25680 29977 25760 30263
rect 25680 29943 25703 29977
rect 25737 29943 25760 29977
rect 25680 29920 25760 29943
rect 25840 30297 25920 30320
rect 25840 30263 25863 30297
rect 25897 30263 25920 30297
rect 25840 29977 25920 30263
rect 25840 29943 25863 29977
rect 25897 29943 25920 29977
rect 25840 29920 25920 29943
rect 26000 30297 26080 30320
rect 26000 30263 26023 30297
rect 26057 30263 26080 30297
rect 26000 29977 26080 30263
rect 26000 29943 26023 29977
rect 26057 29943 26080 29977
rect 26000 29920 26080 29943
rect 26160 30297 26240 30320
rect 26160 30263 26183 30297
rect 26217 30263 26240 30297
rect 26160 29977 26240 30263
rect 26160 29943 26183 29977
rect 26217 29943 26240 29977
rect 26160 29920 26240 29943
rect 26320 30297 26400 30320
rect 26320 30263 26343 30297
rect 26377 30263 26400 30297
rect 26320 29977 26400 30263
rect 26320 29943 26343 29977
rect 26377 29943 26400 29977
rect 26320 29920 26400 29943
rect 26480 30297 26560 30320
rect 26480 30263 26503 30297
rect 26537 30263 26560 30297
rect 26480 29977 26560 30263
rect 26480 29943 26503 29977
rect 26537 29943 26560 29977
rect 26480 29920 26560 29943
rect 26640 30297 26720 30320
rect 26640 30263 26663 30297
rect 26697 30263 26720 30297
rect 26640 29977 26720 30263
rect 26640 29943 26663 29977
rect 26697 29943 26720 29977
rect 26640 29920 26720 29943
rect 26800 30297 26880 30320
rect 26800 30263 26823 30297
rect 26857 30263 26880 30297
rect 26800 29977 26880 30263
rect 26800 29943 26823 29977
rect 26857 29943 26880 29977
rect 26800 29920 26880 29943
rect 26960 30297 27040 30320
rect 26960 30263 26983 30297
rect 27017 30263 27040 30297
rect 26960 29977 27040 30263
rect 26960 29943 26983 29977
rect 27017 29943 27040 29977
rect 26960 29920 27040 29943
rect 27120 30297 27200 30320
rect 27120 30263 27143 30297
rect 27177 30263 27200 30297
rect 27120 29977 27200 30263
rect 27120 29943 27143 29977
rect 27177 29943 27200 29977
rect 27120 29920 27200 29943
rect 27280 30297 27360 30320
rect 27280 30263 27303 30297
rect 27337 30263 27360 30297
rect 27280 29977 27360 30263
rect 27280 29943 27303 29977
rect 27337 29943 27360 29977
rect 27280 29920 27360 29943
rect 27440 30297 27520 30320
rect 27440 30263 27463 30297
rect 27497 30263 27520 30297
rect 27440 29977 27520 30263
rect 27440 29943 27463 29977
rect 27497 29943 27520 29977
rect 27440 29920 27520 29943
rect 27600 30297 27680 30320
rect 27600 30263 27623 30297
rect 27657 30263 27680 30297
rect 27600 29977 27680 30263
rect 27600 29943 27623 29977
rect 27657 29943 27680 29977
rect 27600 29920 27680 29943
rect 27760 30297 27840 30320
rect 27760 30263 27783 30297
rect 27817 30263 27840 30297
rect 27760 29977 27840 30263
rect 27760 29943 27783 29977
rect 27817 29943 27840 29977
rect 27760 29920 27840 29943
rect 27920 30297 28000 30320
rect 27920 30263 27943 30297
rect 27977 30263 28000 30297
rect 27920 29977 28000 30263
rect 27920 29943 27943 29977
rect 27977 29943 28000 29977
rect 27920 29920 28000 29943
rect 28080 30297 28160 30320
rect 28080 30263 28103 30297
rect 28137 30263 28160 30297
rect 28080 29977 28160 30263
rect 28080 29943 28103 29977
rect 28137 29943 28160 29977
rect 28080 29920 28160 29943
rect 28240 30297 28320 30320
rect 28240 30263 28263 30297
rect 28297 30263 28320 30297
rect 28240 29977 28320 30263
rect 28240 29943 28263 29977
rect 28297 29943 28320 29977
rect 28240 29920 28320 29943
rect 28400 30297 28480 30320
rect 28400 30263 28423 30297
rect 28457 30263 28480 30297
rect 28400 29977 28480 30263
rect 28400 29943 28423 29977
rect 28457 29943 28480 29977
rect 28400 29920 28480 29943
rect 28560 30297 28640 30320
rect 28560 30263 28583 30297
rect 28617 30263 28640 30297
rect 28560 29977 28640 30263
rect 28560 29943 28583 29977
rect 28617 29943 28640 29977
rect 28560 29920 28640 29943
rect 28720 30297 28800 30320
rect 28720 30263 28743 30297
rect 28777 30263 28800 30297
rect 28720 29977 28800 30263
rect 28720 29943 28743 29977
rect 28777 29943 28800 29977
rect 28720 29920 28800 29943
rect 28880 30297 28960 30320
rect 28880 30263 28903 30297
rect 28937 30263 28960 30297
rect 28880 29977 28960 30263
rect 28880 29943 28903 29977
rect 28937 29943 28960 29977
rect 28880 29920 28960 29943
rect 29040 30297 29120 30320
rect 29040 30263 29063 30297
rect 29097 30263 29120 30297
rect 29040 29977 29120 30263
rect 29040 29943 29063 29977
rect 29097 29943 29120 29977
rect 29040 29920 29120 29943
rect 29200 30297 29280 30320
rect 29200 30263 29223 30297
rect 29257 30263 29280 30297
rect 29200 29977 29280 30263
rect 29200 29943 29223 29977
rect 29257 29943 29280 29977
rect 29200 29920 29280 29943
rect 29360 30297 29440 30320
rect 29360 30263 29383 30297
rect 29417 30263 29440 30297
rect 29360 29977 29440 30263
rect 29360 29943 29383 29977
rect 29417 29943 29440 29977
rect 29360 29920 29440 29943
rect 29520 29920 29600 30320
rect 29680 29920 29760 30320
rect 29840 29920 29920 30320
rect 30000 29920 30080 30320
rect 30160 29920 30240 30320
rect 30320 29920 30400 30320
rect 30480 29920 30560 30320
rect 30640 29920 30720 30320
rect 30800 29920 30880 30320
rect 30960 29920 31040 30320
rect 31120 29920 31200 30320
rect 31280 29920 31360 30320
rect 31440 29920 31520 30320
rect 31600 29920 31680 30320
rect 31760 29920 31840 30320
rect 31920 29920 32000 30320
rect 32080 29920 32160 30320
rect 32240 29920 32320 30320
rect 32400 29920 32480 30320
rect 32560 29920 32640 30320
rect 32720 29920 32800 30320
rect 32880 29920 32960 30320
rect 33040 29920 33120 30320
rect 33200 29920 33280 30320
rect 33360 29920 33440 30320
rect 33520 30297 33600 30320
rect 33520 30263 33543 30297
rect 33577 30263 33600 30297
rect 33520 29977 33600 30263
rect 33520 29943 33543 29977
rect 33577 29943 33600 29977
rect 33520 29920 33600 29943
rect 33680 30297 33760 30320
rect 33680 30263 33703 30297
rect 33737 30263 33760 30297
rect 33680 29977 33760 30263
rect 33680 29943 33703 29977
rect 33737 29943 33760 29977
rect 33680 29920 33760 29943
rect 33840 30297 33920 30320
rect 33840 30263 33863 30297
rect 33897 30263 33920 30297
rect 33840 29977 33920 30263
rect 33840 29943 33863 29977
rect 33897 29943 33920 29977
rect 33840 29920 33920 29943
rect 34000 30297 34080 30320
rect 34000 30263 34023 30297
rect 34057 30263 34080 30297
rect 34000 29977 34080 30263
rect 34000 29943 34023 29977
rect 34057 29943 34080 29977
rect 34000 29920 34080 29943
rect 34160 30297 34240 30320
rect 34160 30263 34183 30297
rect 34217 30263 34240 30297
rect 34160 29977 34240 30263
rect 34160 29943 34183 29977
rect 34217 29943 34240 29977
rect 34160 29920 34240 29943
rect 34320 30297 34400 30320
rect 34320 30263 34343 30297
rect 34377 30263 34400 30297
rect 34320 29977 34400 30263
rect 34320 29943 34343 29977
rect 34377 29943 34400 29977
rect 34320 29920 34400 29943
rect 34480 30297 34560 30320
rect 34480 30263 34503 30297
rect 34537 30263 34560 30297
rect 34480 29977 34560 30263
rect 34480 29943 34503 29977
rect 34537 29943 34560 29977
rect 34480 29920 34560 29943
rect 34640 30297 34720 30320
rect 34640 30263 34663 30297
rect 34697 30263 34720 30297
rect 34640 29977 34720 30263
rect 34640 29943 34663 29977
rect 34697 29943 34720 29977
rect 34640 29920 34720 29943
rect 34800 30297 34880 30320
rect 34800 30263 34823 30297
rect 34857 30263 34880 30297
rect 34800 29977 34880 30263
rect 34800 29943 34823 29977
rect 34857 29943 34880 29977
rect 34800 29920 34880 29943
rect 34960 30297 35040 30320
rect 34960 30263 34983 30297
rect 35017 30263 35040 30297
rect 34960 29977 35040 30263
rect 34960 29943 34983 29977
rect 35017 29943 35040 29977
rect 34960 29920 35040 29943
rect 35120 30297 35200 30320
rect 35120 30263 35143 30297
rect 35177 30263 35200 30297
rect 35120 29977 35200 30263
rect 35120 29943 35143 29977
rect 35177 29943 35200 29977
rect 35120 29920 35200 29943
rect 35280 30297 35360 30320
rect 35280 30263 35303 30297
rect 35337 30263 35360 30297
rect 35280 29977 35360 30263
rect 35280 29943 35303 29977
rect 35337 29943 35360 29977
rect 35280 29920 35360 29943
rect 35440 30297 35520 30320
rect 35440 30263 35463 30297
rect 35497 30263 35520 30297
rect 35440 29977 35520 30263
rect 35440 29943 35463 29977
rect 35497 29943 35520 29977
rect 35440 29920 35520 29943
rect 35600 30297 35680 30320
rect 35600 30263 35623 30297
rect 35657 30263 35680 30297
rect 35600 29977 35680 30263
rect 35600 29943 35623 29977
rect 35657 29943 35680 29977
rect 35600 29920 35680 29943
rect 35760 30297 35840 30320
rect 35760 30263 35783 30297
rect 35817 30263 35840 30297
rect 35760 29977 35840 30263
rect 35760 29943 35783 29977
rect 35817 29943 35840 29977
rect 35760 29920 35840 29943
rect 35920 30297 36000 30320
rect 35920 30263 35943 30297
rect 35977 30263 36000 30297
rect 35920 29977 36000 30263
rect 35920 29943 35943 29977
rect 35977 29943 36000 29977
rect 35920 29920 36000 29943
rect 36080 30297 36160 30320
rect 36080 30263 36103 30297
rect 36137 30263 36160 30297
rect 36080 29977 36160 30263
rect 36080 29943 36103 29977
rect 36137 29943 36160 29977
rect 36080 29920 36160 29943
rect 36240 30297 36320 30320
rect 36240 30263 36263 30297
rect 36297 30263 36320 30297
rect 36240 29977 36320 30263
rect 36240 29943 36263 29977
rect 36297 29943 36320 29977
rect 36240 29920 36320 29943
rect 36400 30297 36480 30320
rect 36400 30263 36423 30297
rect 36457 30263 36480 30297
rect 36400 29977 36480 30263
rect 36400 29943 36423 29977
rect 36457 29943 36480 29977
rect 36400 29920 36480 29943
rect 36560 30297 36640 30320
rect 36560 30263 36583 30297
rect 36617 30263 36640 30297
rect 36560 29977 36640 30263
rect 36560 29943 36583 29977
rect 36617 29943 36640 29977
rect 36560 29920 36640 29943
rect 36720 30297 36800 30320
rect 36720 30263 36743 30297
rect 36777 30263 36800 30297
rect 36720 29977 36800 30263
rect 36720 29943 36743 29977
rect 36777 29943 36800 29977
rect 36720 29920 36800 29943
rect 36880 30297 36960 30320
rect 36880 30263 36903 30297
rect 36937 30263 36960 30297
rect 36880 29977 36960 30263
rect 36880 29943 36903 29977
rect 36937 29943 36960 29977
rect 36880 29920 36960 29943
rect 37040 30297 37120 30320
rect 37040 30263 37063 30297
rect 37097 30263 37120 30297
rect 37040 29977 37120 30263
rect 37040 29943 37063 29977
rect 37097 29943 37120 29977
rect 37040 29920 37120 29943
rect 37200 30297 37280 30320
rect 37200 30263 37223 30297
rect 37257 30263 37280 30297
rect 37200 29977 37280 30263
rect 37200 29943 37223 29977
rect 37257 29943 37280 29977
rect 37200 29920 37280 29943
rect 37360 30297 37440 30320
rect 37360 30263 37383 30297
rect 37417 30263 37440 30297
rect 37360 29977 37440 30263
rect 37360 29943 37383 29977
rect 37417 29943 37440 29977
rect 37360 29920 37440 29943
rect 37520 30297 37600 30320
rect 37520 30263 37543 30297
rect 37577 30263 37600 30297
rect 37520 29977 37600 30263
rect 37520 29943 37543 29977
rect 37577 29943 37600 29977
rect 37520 29920 37600 29943
rect 37680 30297 37760 30320
rect 37680 30263 37703 30297
rect 37737 30263 37760 30297
rect 37680 29977 37760 30263
rect 37680 29943 37703 29977
rect 37737 29943 37760 29977
rect 37680 29920 37760 29943
rect 37840 30297 37920 30320
rect 37840 30263 37863 30297
rect 37897 30263 37920 30297
rect 37840 29977 37920 30263
rect 37840 29943 37863 29977
rect 37897 29943 37920 29977
rect 37840 29920 37920 29943
rect 38000 30297 38080 30320
rect 38000 30263 38023 30297
rect 38057 30263 38080 30297
rect 38000 29977 38080 30263
rect 38000 29943 38023 29977
rect 38057 29943 38080 29977
rect 38000 29920 38080 29943
rect 38160 30297 38240 30320
rect 38160 30263 38183 30297
rect 38217 30263 38240 30297
rect 38160 29977 38240 30263
rect 38160 29943 38183 29977
rect 38217 29943 38240 29977
rect 38160 29920 38240 29943
rect 38320 30297 38400 30320
rect 38320 30263 38343 30297
rect 38377 30263 38400 30297
rect 38320 29977 38400 30263
rect 38320 29943 38343 29977
rect 38377 29943 38400 29977
rect 38320 29920 38400 29943
rect 38480 30297 38560 30320
rect 38480 30263 38503 30297
rect 38537 30263 38560 30297
rect 38480 29977 38560 30263
rect 38480 29943 38503 29977
rect 38537 29943 38560 29977
rect 38480 29920 38560 29943
rect 38640 30297 38720 30320
rect 38640 30263 38663 30297
rect 38697 30263 38720 30297
rect 38640 29977 38720 30263
rect 38640 29943 38663 29977
rect 38697 29943 38720 29977
rect 38640 29920 38720 29943
rect 38800 30297 38880 30320
rect 38800 30263 38823 30297
rect 38857 30263 38880 30297
rect 38800 29977 38880 30263
rect 38800 29943 38823 29977
rect 38857 29943 38880 29977
rect 38800 29920 38880 29943
rect 38960 30297 39040 30320
rect 38960 30263 38983 30297
rect 39017 30263 39040 30297
rect 38960 29977 39040 30263
rect 38960 29943 38983 29977
rect 39017 29943 39040 29977
rect 38960 29920 39040 29943
rect 39120 30297 39200 30320
rect 39120 30263 39143 30297
rect 39177 30263 39200 30297
rect 39120 29977 39200 30263
rect 39120 29943 39143 29977
rect 39177 29943 39200 29977
rect 39120 29920 39200 29943
rect 39280 30297 39360 30320
rect 39280 30263 39303 30297
rect 39337 30263 39360 30297
rect 39280 29977 39360 30263
rect 39280 29943 39303 29977
rect 39337 29943 39360 29977
rect 39280 29920 39360 29943
rect 39440 30297 39520 30320
rect 39440 30263 39463 30297
rect 39497 30263 39520 30297
rect 39440 29977 39520 30263
rect 39440 29943 39463 29977
rect 39497 29943 39520 29977
rect 39440 29920 39520 29943
rect 39600 30297 39680 30320
rect 39600 30263 39623 30297
rect 39657 30263 39680 30297
rect 39600 29977 39680 30263
rect 39600 29943 39623 29977
rect 39657 29943 39680 29977
rect 39600 29920 39680 29943
rect 39760 30297 39840 30320
rect 39760 30263 39783 30297
rect 39817 30263 39840 30297
rect 39760 29977 39840 30263
rect 39760 29943 39783 29977
rect 39817 29943 39840 29977
rect 39760 29920 39840 29943
rect 39920 30297 40000 30320
rect 39920 30263 39943 30297
rect 39977 30263 40000 30297
rect 39920 29977 40000 30263
rect 39920 29943 39943 29977
rect 39977 29943 40000 29977
rect 39920 29920 40000 29943
rect 40080 30297 40160 30320
rect 40080 30263 40103 30297
rect 40137 30263 40160 30297
rect 40080 29977 40160 30263
rect 40080 29943 40103 29977
rect 40137 29943 40160 29977
rect 40080 29920 40160 29943
rect 40240 30297 40320 30320
rect 40240 30263 40263 30297
rect 40297 30263 40320 30297
rect 40240 29977 40320 30263
rect 40240 29943 40263 29977
rect 40297 29943 40320 29977
rect 40240 29920 40320 29943
rect 40400 30297 40480 30320
rect 40400 30263 40423 30297
rect 40457 30263 40480 30297
rect 40400 29977 40480 30263
rect 40400 29943 40423 29977
rect 40457 29943 40480 29977
rect 40400 29920 40480 29943
rect 40560 30297 40640 30320
rect 40560 30263 40583 30297
rect 40617 30263 40640 30297
rect 40560 29977 40640 30263
rect 40560 29943 40583 29977
rect 40617 29943 40640 29977
rect 40560 29920 40640 29943
rect 40720 30297 40800 30320
rect 40720 30263 40743 30297
rect 40777 30263 40800 30297
rect 40720 29977 40800 30263
rect 40720 29943 40743 29977
rect 40777 29943 40800 29977
rect 40720 29920 40800 29943
rect 40880 30297 40960 30320
rect 40880 30263 40903 30297
rect 40937 30263 40960 30297
rect 40880 29977 40960 30263
rect 40880 29943 40903 29977
rect 40937 29943 40960 29977
rect 40880 29920 40960 29943
rect 41040 30297 41120 30320
rect 41040 30263 41063 30297
rect 41097 30263 41120 30297
rect 41040 29977 41120 30263
rect 41040 29943 41063 29977
rect 41097 29943 41120 29977
rect 41040 29920 41120 29943
rect 41200 30297 41280 30320
rect 41200 30263 41223 30297
rect 41257 30263 41280 30297
rect 41200 29977 41280 30263
rect 41200 29943 41223 29977
rect 41257 29943 41280 29977
rect 41200 29920 41280 29943
rect 41360 30297 41440 30320
rect 41360 30263 41383 30297
rect 41417 30263 41440 30297
rect 41360 29977 41440 30263
rect 41360 29943 41383 29977
rect 41417 29943 41440 29977
rect 41360 29920 41440 29943
rect 41520 30297 41600 30320
rect 41520 30263 41543 30297
rect 41577 30263 41600 30297
rect 41520 29977 41600 30263
rect 41520 29943 41543 29977
rect 41577 29943 41600 29977
rect 41520 29920 41600 29943
rect 41680 30297 41760 30320
rect 41680 30263 41703 30297
rect 41737 30263 41760 30297
rect 41680 29977 41760 30263
rect 41680 29943 41703 29977
rect 41737 29943 41760 29977
rect 41680 29920 41760 29943
rect 41840 30297 41920 30320
rect 41840 30263 41863 30297
rect 41897 30263 41920 30297
rect 41840 29977 41920 30263
rect 41840 29943 41863 29977
rect 41897 29943 41920 29977
rect 41840 29920 41920 29943
rect 0 29817 80 29840
rect 0 29783 23 29817
rect 57 29783 80 29817
rect 0 29497 80 29783
rect 0 29463 23 29497
rect 57 29463 80 29497
rect 0 29440 80 29463
rect 160 29817 240 29840
rect 160 29783 183 29817
rect 217 29783 240 29817
rect 160 29497 240 29783
rect 160 29463 183 29497
rect 217 29463 240 29497
rect 160 29440 240 29463
rect 320 29817 400 29840
rect 320 29783 343 29817
rect 377 29783 400 29817
rect 320 29497 400 29783
rect 320 29463 343 29497
rect 377 29463 400 29497
rect 320 29440 400 29463
rect 480 29817 560 29840
rect 480 29783 503 29817
rect 537 29783 560 29817
rect 480 29497 560 29783
rect 480 29463 503 29497
rect 537 29463 560 29497
rect 480 29440 560 29463
rect 640 29817 720 29840
rect 640 29783 663 29817
rect 697 29783 720 29817
rect 640 29497 720 29783
rect 640 29463 663 29497
rect 697 29463 720 29497
rect 640 29440 720 29463
rect 800 29817 880 29840
rect 800 29783 823 29817
rect 857 29783 880 29817
rect 800 29497 880 29783
rect 800 29463 823 29497
rect 857 29463 880 29497
rect 800 29440 880 29463
rect 960 29817 1040 29840
rect 960 29783 983 29817
rect 1017 29783 1040 29817
rect 960 29497 1040 29783
rect 960 29463 983 29497
rect 1017 29463 1040 29497
rect 960 29440 1040 29463
rect 1120 29817 1200 29840
rect 1120 29783 1143 29817
rect 1177 29783 1200 29817
rect 1120 29497 1200 29783
rect 1120 29463 1143 29497
rect 1177 29463 1200 29497
rect 1120 29440 1200 29463
rect 1280 29817 1360 29840
rect 1280 29783 1303 29817
rect 1337 29783 1360 29817
rect 1280 29497 1360 29783
rect 1280 29463 1303 29497
rect 1337 29463 1360 29497
rect 1280 29440 1360 29463
rect 1440 29817 1520 29840
rect 1440 29783 1463 29817
rect 1497 29783 1520 29817
rect 1440 29497 1520 29783
rect 1440 29463 1463 29497
rect 1497 29463 1520 29497
rect 1440 29440 1520 29463
rect 1600 29817 1680 29840
rect 1600 29783 1623 29817
rect 1657 29783 1680 29817
rect 1600 29497 1680 29783
rect 1600 29463 1623 29497
rect 1657 29463 1680 29497
rect 1600 29440 1680 29463
rect 1760 29817 1840 29840
rect 1760 29783 1783 29817
rect 1817 29783 1840 29817
rect 1760 29497 1840 29783
rect 1760 29463 1783 29497
rect 1817 29463 1840 29497
rect 1760 29440 1840 29463
rect 1920 29817 2000 29840
rect 1920 29783 1943 29817
rect 1977 29783 2000 29817
rect 1920 29497 2000 29783
rect 1920 29463 1943 29497
rect 1977 29463 2000 29497
rect 1920 29440 2000 29463
rect 2080 29817 2160 29840
rect 2080 29783 2103 29817
rect 2137 29783 2160 29817
rect 2080 29497 2160 29783
rect 2080 29463 2103 29497
rect 2137 29463 2160 29497
rect 2080 29440 2160 29463
rect 2240 29817 2320 29840
rect 2240 29783 2263 29817
rect 2297 29783 2320 29817
rect 2240 29497 2320 29783
rect 2240 29463 2263 29497
rect 2297 29463 2320 29497
rect 2240 29440 2320 29463
rect 2400 29817 2480 29840
rect 2400 29783 2423 29817
rect 2457 29783 2480 29817
rect 2400 29497 2480 29783
rect 2400 29463 2423 29497
rect 2457 29463 2480 29497
rect 2400 29440 2480 29463
rect 2560 29817 2640 29840
rect 2560 29783 2583 29817
rect 2617 29783 2640 29817
rect 2560 29497 2640 29783
rect 2560 29463 2583 29497
rect 2617 29463 2640 29497
rect 2560 29440 2640 29463
rect 2720 29817 2800 29840
rect 2720 29783 2743 29817
rect 2777 29783 2800 29817
rect 2720 29497 2800 29783
rect 2720 29463 2743 29497
rect 2777 29463 2800 29497
rect 2720 29440 2800 29463
rect 2880 29817 2960 29840
rect 2880 29783 2903 29817
rect 2937 29783 2960 29817
rect 2880 29497 2960 29783
rect 2880 29463 2903 29497
rect 2937 29463 2960 29497
rect 2880 29440 2960 29463
rect 3040 29817 3120 29840
rect 3040 29783 3063 29817
rect 3097 29783 3120 29817
rect 3040 29497 3120 29783
rect 3040 29463 3063 29497
rect 3097 29463 3120 29497
rect 3040 29440 3120 29463
rect 3200 29817 3280 29840
rect 3200 29783 3223 29817
rect 3257 29783 3280 29817
rect 3200 29497 3280 29783
rect 3200 29463 3223 29497
rect 3257 29463 3280 29497
rect 3200 29440 3280 29463
rect 3360 29817 3440 29840
rect 3360 29783 3383 29817
rect 3417 29783 3440 29817
rect 3360 29497 3440 29783
rect 3360 29463 3383 29497
rect 3417 29463 3440 29497
rect 3360 29440 3440 29463
rect 3520 29817 3600 29840
rect 3520 29783 3543 29817
rect 3577 29783 3600 29817
rect 3520 29497 3600 29783
rect 3520 29463 3543 29497
rect 3577 29463 3600 29497
rect 3520 29440 3600 29463
rect 3680 29817 3760 29840
rect 3680 29783 3703 29817
rect 3737 29783 3760 29817
rect 3680 29497 3760 29783
rect 3680 29463 3703 29497
rect 3737 29463 3760 29497
rect 3680 29440 3760 29463
rect 3840 29817 3920 29840
rect 3840 29783 3863 29817
rect 3897 29783 3920 29817
rect 3840 29497 3920 29783
rect 3840 29463 3863 29497
rect 3897 29463 3920 29497
rect 3840 29440 3920 29463
rect 4000 29817 4080 29840
rect 4000 29783 4023 29817
rect 4057 29783 4080 29817
rect 4000 29497 4080 29783
rect 4000 29463 4023 29497
rect 4057 29463 4080 29497
rect 4000 29440 4080 29463
rect 4160 29817 4240 29840
rect 4160 29783 4183 29817
rect 4217 29783 4240 29817
rect 4160 29497 4240 29783
rect 4160 29463 4183 29497
rect 4217 29463 4240 29497
rect 4160 29440 4240 29463
rect 4320 29817 4400 29840
rect 4320 29783 4343 29817
rect 4377 29783 4400 29817
rect 4320 29497 4400 29783
rect 4320 29463 4343 29497
rect 4377 29463 4400 29497
rect 4320 29440 4400 29463
rect 4480 29817 4560 29840
rect 4480 29783 4503 29817
rect 4537 29783 4560 29817
rect 4480 29497 4560 29783
rect 4480 29463 4503 29497
rect 4537 29463 4560 29497
rect 4480 29440 4560 29463
rect 4640 29817 4720 29840
rect 4640 29783 4663 29817
rect 4697 29783 4720 29817
rect 4640 29497 4720 29783
rect 4640 29463 4663 29497
rect 4697 29463 4720 29497
rect 4640 29440 4720 29463
rect 4800 29817 4880 29840
rect 4800 29783 4823 29817
rect 4857 29783 4880 29817
rect 4800 29497 4880 29783
rect 4800 29463 4823 29497
rect 4857 29463 4880 29497
rect 4800 29440 4880 29463
rect 4960 29817 5040 29840
rect 4960 29783 4983 29817
rect 5017 29783 5040 29817
rect 4960 29497 5040 29783
rect 4960 29463 4983 29497
rect 5017 29463 5040 29497
rect 4960 29440 5040 29463
rect 5120 29817 5200 29840
rect 5120 29783 5143 29817
rect 5177 29783 5200 29817
rect 5120 29497 5200 29783
rect 5120 29463 5143 29497
rect 5177 29463 5200 29497
rect 5120 29440 5200 29463
rect 5280 29817 5360 29840
rect 5280 29783 5303 29817
rect 5337 29783 5360 29817
rect 5280 29497 5360 29783
rect 5280 29463 5303 29497
rect 5337 29463 5360 29497
rect 5280 29440 5360 29463
rect 5440 29817 5520 29840
rect 5440 29783 5463 29817
rect 5497 29783 5520 29817
rect 5440 29497 5520 29783
rect 5440 29463 5463 29497
rect 5497 29463 5520 29497
rect 5440 29440 5520 29463
rect 5600 29817 5680 29840
rect 5600 29783 5623 29817
rect 5657 29783 5680 29817
rect 5600 29497 5680 29783
rect 5600 29463 5623 29497
rect 5657 29463 5680 29497
rect 5600 29440 5680 29463
rect 5760 29817 5840 29840
rect 5760 29783 5783 29817
rect 5817 29783 5840 29817
rect 5760 29497 5840 29783
rect 5760 29463 5783 29497
rect 5817 29463 5840 29497
rect 5760 29440 5840 29463
rect 5920 29817 6000 29840
rect 5920 29783 5943 29817
rect 5977 29783 6000 29817
rect 5920 29497 6000 29783
rect 5920 29463 5943 29497
rect 5977 29463 6000 29497
rect 5920 29440 6000 29463
rect 6080 29817 6160 29840
rect 6080 29783 6103 29817
rect 6137 29783 6160 29817
rect 6080 29497 6160 29783
rect 6080 29463 6103 29497
rect 6137 29463 6160 29497
rect 6080 29440 6160 29463
rect 6240 29817 6320 29840
rect 6240 29783 6263 29817
rect 6297 29783 6320 29817
rect 6240 29497 6320 29783
rect 6240 29463 6263 29497
rect 6297 29463 6320 29497
rect 6240 29440 6320 29463
rect 6400 29817 6480 29840
rect 6400 29783 6423 29817
rect 6457 29783 6480 29817
rect 6400 29497 6480 29783
rect 6400 29463 6423 29497
rect 6457 29463 6480 29497
rect 6400 29440 6480 29463
rect 6560 29817 6640 29840
rect 6560 29783 6583 29817
rect 6617 29783 6640 29817
rect 6560 29497 6640 29783
rect 6560 29463 6583 29497
rect 6617 29463 6640 29497
rect 6560 29440 6640 29463
rect 6720 29817 6800 29840
rect 6720 29783 6743 29817
rect 6777 29783 6800 29817
rect 6720 29497 6800 29783
rect 6720 29463 6743 29497
rect 6777 29463 6800 29497
rect 6720 29440 6800 29463
rect 6880 29817 6960 29840
rect 6880 29783 6903 29817
rect 6937 29783 6960 29817
rect 6880 29497 6960 29783
rect 6880 29463 6903 29497
rect 6937 29463 6960 29497
rect 6880 29440 6960 29463
rect 7040 29817 7120 29840
rect 7040 29783 7063 29817
rect 7097 29783 7120 29817
rect 7040 29497 7120 29783
rect 7040 29463 7063 29497
rect 7097 29463 7120 29497
rect 7040 29440 7120 29463
rect 7200 29817 7280 29840
rect 7200 29783 7223 29817
rect 7257 29783 7280 29817
rect 7200 29497 7280 29783
rect 7200 29463 7223 29497
rect 7257 29463 7280 29497
rect 7200 29440 7280 29463
rect 7360 29817 7440 29840
rect 7360 29783 7383 29817
rect 7417 29783 7440 29817
rect 7360 29497 7440 29783
rect 7360 29463 7383 29497
rect 7417 29463 7440 29497
rect 7360 29440 7440 29463
rect 7520 29817 7600 29840
rect 7520 29783 7543 29817
rect 7577 29783 7600 29817
rect 7520 29497 7600 29783
rect 7520 29463 7543 29497
rect 7577 29463 7600 29497
rect 7520 29440 7600 29463
rect 7680 29817 7760 29840
rect 7680 29783 7703 29817
rect 7737 29783 7760 29817
rect 7680 29497 7760 29783
rect 7680 29463 7703 29497
rect 7737 29463 7760 29497
rect 7680 29440 7760 29463
rect 7840 29817 7920 29840
rect 7840 29783 7863 29817
rect 7897 29783 7920 29817
rect 7840 29497 7920 29783
rect 7840 29463 7863 29497
rect 7897 29463 7920 29497
rect 7840 29440 7920 29463
rect 8000 29817 8080 29840
rect 8000 29783 8023 29817
rect 8057 29783 8080 29817
rect 8000 29497 8080 29783
rect 8000 29463 8023 29497
rect 8057 29463 8080 29497
rect 8000 29440 8080 29463
rect 8160 29817 8240 29840
rect 8160 29783 8183 29817
rect 8217 29783 8240 29817
rect 8160 29497 8240 29783
rect 8160 29463 8183 29497
rect 8217 29463 8240 29497
rect 8160 29440 8240 29463
rect 8320 29817 8400 29840
rect 8320 29783 8343 29817
rect 8377 29783 8400 29817
rect 8320 29497 8400 29783
rect 8320 29463 8343 29497
rect 8377 29463 8400 29497
rect 8320 29440 8400 29463
rect 8480 29440 8560 29840
rect 8640 29440 8720 29840
rect 8800 29440 8880 29840
rect 8960 29440 9040 29840
rect 9120 29440 9200 29840
rect 9280 29440 9360 29840
rect 9440 29440 9520 29840
rect 9600 29440 9680 29840
rect 9760 29440 9840 29840
rect 9920 29440 10000 29840
rect 10080 29440 10160 29840
rect 10240 29440 10320 29840
rect 10400 29440 10480 29840
rect 10560 29440 10640 29840
rect 10720 29440 10800 29840
rect 10880 29440 10960 29840
rect 11040 29440 11120 29840
rect 11200 29440 11280 29840
rect 11360 29440 11440 29840
rect 11520 29440 11600 29840
rect 11680 29440 11760 29840
rect 11840 29440 11920 29840
rect 12000 29440 12080 29840
rect 12160 29440 12240 29840
rect 12320 29440 12400 29840
rect 12480 29817 12560 29840
rect 12480 29783 12503 29817
rect 12537 29783 12560 29817
rect 12480 29497 12560 29783
rect 12480 29463 12503 29497
rect 12537 29463 12560 29497
rect 12480 29440 12560 29463
rect 12640 29817 12720 29840
rect 12640 29783 12663 29817
rect 12697 29783 12720 29817
rect 12640 29497 12720 29783
rect 12640 29463 12663 29497
rect 12697 29463 12720 29497
rect 12640 29440 12720 29463
rect 12800 29817 12880 29840
rect 12800 29783 12823 29817
rect 12857 29783 12880 29817
rect 12800 29497 12880 29783
rect 12800 29463 12823 29497
rect 12857 29463 12880 29497
rect 12800 29440 12880 29463
rect 12960 29817 13040 29840
rect 12960 29783 12983 29817
rect 13017 29783 13040 29817
rect 12960 29497 13040 29783
rect 12960 29463 12983 29497
rect 13017 29463 13040 29497
rect 12960 29440 13040 29463
rect 13120 29817 13200 29840
rect 13120 29783 13143 29817
rect 13177 29783 13200 29817
rect 13120 29497 13200 29783
rect 13120 29463 13143 29497
rect 13177 29463 13200 29497
rect 13120 29440 13200 29463
rect 13280 29817 13360 29840
rect 13280 29783 13303 29817
rect 13337 29783 13360 29817
rect 13280 29497 13360 29783
rect 13280 29463 13303 29497
rect 13337 29463 13360 29497
rect 13280 29440 13360 29463
rect 13440 29817 13520 29840
rect 13440 29783 13463 29817
rect 13497 29783 13520 29817
rect 13440 29497 13520 29783
rect 13440 29463 13463 29497
rect 13497 29463 13520 29497
rect 13440 29440 13520 29463
rect 13600 29817 13680 29840
rect 13600 29783 13623 29817
rect 13657 29783 13680 29817
rect 13600 29497 13680 29783
rect 13600 29463 13623 29497
rect 13657 29463 13680 29497
rect 13600 29440 13680 29463
rect 13760 29817 13840 29840
rect 13760 29783 13783 29817
rect 13817 29783 13840 29817
rect 13760 29497 13840 29783
rect 13760 29463 13783 29497
rect 13817 29463 13840 29497
rect 13760 29440 13840 29463
rect 13920 29817 14000 29840
rect 13920 29783 13943 29817
rect 13977 29783 14000 29817
rect 13920 29497 14000 29783
rect 13920 29463 13943 29497
rect 13977 29463 14000 29497
rect 13920 29440 14000 29463
rect 14080 29817 14160 29840
rect 14080 29783 14103 29817
rect 14137 29783 14160 29817
rect 14080 29497 14160 29783
rect 14080 29463 14103 29497
rect 14137 29463 14160 29497
rect 14080 29440 14160 29463
rect 14240 29817 14320 29840
rect 14240 29783 14263 29817
rect 14297 29783 14320 29817
rect 14240 29497 14320 29783
rect 14240 29463 14263 29497
rect 14297 29463 14320 29497
rect 14240 29440 14320 29463
rect 14400 29817 14480 29840
rect 14400 29783 14423 29817
rect 14457 29783 14480 29817
rect 14400 29497 14480 29783
rect 14400 29463 14423 29497
rect 14457 29463 14480 29497
rect 14400 29440 14480 29463
rect 14560 29817 14640 29840
rect 14560 29783 14583 29817
rect 14617 29783 14640 29817
rect 14560 29497 14640 29783
rect 14560 29463 14583 29497
rect 14617 29463 14640 29497
rect 14560 29440 14640 29463
rect 14720 29817 14800 29840
rect 14720 29783 14743 29817
rect 14777 29783 14800 29817
rect 14720 29497 14800 29783
rect 14720 29463 14743 29497
rect 14777 29463 14800 29497
rect 14720 29440 14800 29463
rect 14880 29817 14960 29840
rect 14880 29783 14903 29817
rect 14937 29783 14960 29817
rect 14880 29497 14960 29783
rect 14880 29463 14903 29497
rect 14937 29463 14960 29497
rect 14880 29440 14960 29463
rect 15040 29817 15120 29840
rect 15040 29783 15063 29817
rect 15097 29783 15120 29817
rect 15040 29497 15120 29783
rect 15040 29463 15063 29497
rect 15097 29463 15120 29497
rect 15040 29440 15120 29463
rect 15200 29817 15280 29840
rect 15200 29783 15223 29817
rect 15257 29783 15280 29817
rect 15200 29497 15280 29783
rect 15200 29463 15223 29497
rect 15257 29463 15280 29497
rect 15200 29440 15280 29463
rect 15360 29817 15440 29840
rect 15360 29783 15383 29817
rect 15417 29783 15440 29817
rect 15360 29497 15440 29783
rect 15360 29463 15383 29497
rect 15417 29463 15440 29497
rect 15360 29440 15440 29463
rect 15520 29817 15600 29840
rect 15520 29783 15543 29817
rect 15577 29783 15600 29817
rect 15520 29497 15600 29783
rect 15520 29463 15543 29497
rect 15577 29463 15600 29497
rect 15520 29440 15600 29463
rect 15680 29817 15760 29840
rect 15680 29783 15703 29817
rect 15737 29783 15760 29817
rect 15680 29497 15760 29783
rect 15680 29463 15703 29497
rect 15737 29463 15760 29497
rect 15680 29440 15760 29463
rect 15840 29817 15920 29840
rect 15840 29783 15863 29817
rect 15897 29783 15920 29817
rect 15840 29497 15920 29783
rect 15840 29463 15863 29497
rect 15897 29463 15920 29497
rect 15840 29440 15920 29463
rect 16000 29817 16080 29840
rect 16000 29783 16023 29817
rect 16057 29783 16080 29817
rect 16000 29497 16080 29783
rect 16000 29463 16023 29497
rect 16057 29463 16080 29497
rect 16000 29440 16080 29463
rect 16160 29817 16240 29840
rect 16160 29783 16183 29817
rect 16217 29783 16240 29817
rect 16160 29497 16240 29783
rect 16160 29463 16183 29497
rect 16217 29463 16240 29497
rect 16160 29440 16240 29463
rect 16320 29817 16400 29840
rect 16320 29783 16343 29817
rect 16377 29783 16400 29817
rect 16320 29497 16400 29783
rect 16320 29463 16343 29497
rect 16377 29463 16400 29497
rect 16320 29440 16400 29463
rect 16480 29817 16560 29840
rect 16480 29783 16503 29817
rect 16537 29783 16560 29817
rect 16480 29497 16560 29783
rect 16480 29463 16503 29497
rect 16537 29463 16560 29497
rect 16480 29440 16560 29463
rect 16640 29817 16720 29840
rect 16640 29783 16663 29817
rect 16697 29783 16720 29817
rect 16640 29497 16720 29783
rect 16640 29463 16663 29497
rect 16697 29463 16720 29497
rect 16640 29440 16720 29463
rect 16800 29817 16880 29840
rect 16800 29783 16823 29817
rect 16857 29783 16880 29817
rect 16800 29497 16880 29783
rect 16800 29463 16823 29497
rect 16857 29463 16880 29497
rect 16800 29440 16880 29463
rect 16960 29817 17040 29840
rect 16960 29783 16983 29817
rect 17017 29783 17040 29817
rect 16960 29497 17040 29783
rect 16960 29463 16983 29497
rect 17017 29463 17040 29497
rect 16960 29440 17040 29463
rect 17120 29817 17200 29840
rect 17120 29783 17143 29817
rect 17177 29783 17200 29817
rect 17120 29497 17200 29783
rect 17120 29463 17143 29497
rect 17177 29463 17200 29497
rect 17120 29440 17200 29463
rect 17280 29817 17360 29840
rect 17280 29783 17303 29817
rect 17337 29783 17360 29817
rect 17280 29497 17360 29783
rect 17280 29463 17303 29497
rect 17337 29463 17360 29497
rect 17280 29440 17360 29463
rect 17440 29817 17520 29840
rect 17440 29783 17463 29817
rect 17497 29783 17520 29817
rect 17440 29497 17520 29783
rect 17440 29463 17463 29497
rect 17497 29463 17520 29497
rect 17440 29440 17520 29463
rect 17600 29817 17680 29840
rect 17600 29783 17623 29817
rect 17657 29783 17680 29817
rect 17600 29497 17680 29783
rect 17600 29463 17623 29497
rect 17657 29463 17680 29497
rect 17600 29440 17680 29463
rect 17760 29817 17840 29840
rect 17760 29783 17783 29817
rect 17817 29783 17840 29817
rect 17760 29497 17840 29783
rect 17760 29463 17783 29497
rect 17817 29463 17840 29497
rect 17760 29440 17840 29463
rect 17920 29817 18000 29840
rect 17920 29783 17943 29817
rect 17977 29783 18000 29817
rect 17920 29497 18000 29783
rect 17920 29463 17943 29497
rect 17977 29463 18000 29497
rect 17920 29440 18000 29463
rect 18080 29817 18160 29840
rect 18080 29783 18103 29817
rect 18137 29783 18160 29817
rect 18080 29497 18160 29783
rect 18080 29463 18103 29497
rect 18137 29463 18160 29497
rect 18080 29440 18160 29463
rect 18240 29817 18320 29840
rect 18240 29783 18263 29817
rect 18297 29783 18320 29817
rect 18240 29497 18320 29783
rect 18240 29463 18263 29497
rect 18297 29463 18320 29497
rect 18240 29440 18320 29463
rect 18400 29817 18480 29840
rect 18400 29783 18423 29817
rect 18457 29783 18480 29817
rect 18400 29497 18480 29783
rect 18400 29463 18423 29497
rect 18457 29463 18480 29497
rect 18400 29440 18480 29463
rect 18560 29817 18640 29840
rect 18560 29783 18583 29817
rect 18617 29783 18640 29817
rect 18560 29497 18640 29783
rect 18560 29463 18583 29497
rect 18617 29463 18640 29497
rect 18560 29440 18640 29463
rect 18720 29817 18800 29840
rect 18720 29783 18743 29817
rect 18777 29783 18800 29817
rect 18720 29497 18800 29783
rect 18720 29463 18743 29497
rect 18777 29463 18800 29497
rect 18720 29440 18800 29463
rect 18880 29817 18960 29840
rect 18880 29783 18903 29817
rect 18937 29783 18960 29817
rect 18880 29497 18960 29783
rect 18880 29463 18903 29497
rect 18937 29463 18960 29497
rect 18880 29440 18960 29463
rect 19040 29440 19120 29840
rect 19200 29440 19280 29840
rect 19360 29440 19440 29840
rect 19520 29440 19600 29840
rect 19680 29440 19760 29840
rect 19840 29440 19920 29840
rect 20000 29440 20080 29840
rect 20160 29440 20240 29840
rect 20320 29440 20400 29840
rect 20480 29440 20560 29840
rect 20640 29440 20720 29840
rect 20800 29440 20880 29840
rect 20960 29440 21040 29840
rect 21120 29440 21200 29840
rect 21280 29440 21360 29840
rect 21440 29440 21520 29840
rect 21600 29440 21680 29840
rect 21760 29440 21840 29840
rect 21920 29440 22000 29840
rect 22080 29440 22160 29840
rect 22240 29440 22320 29840
rect 22400 29440 22480 29840
rect 22560 29440 22640 29840
rect 22720 29440 22800 29840
rect 22880 29440 22960 29840
rect 23120 29817 23200 29840
rect 23120 29783 23143 29817
rect 23177 29783 23200 29817
rect 23120 29497 23200 29783
rect 23120 29463 23143 29497
rect 23177 29463 23200 29497
rect 23120 29440 23200 29463
rect 23280 29817 23360 29840
rect 23280 29783 23303 29817
rect 23337 29783 23360 29817
rect 23280 29497 23360 29783
rect 23280 29463 23303 29497
rect 23337 29463 23360 29497
rect 23280 29440 23360 29463
rect 23440 29817 23520 29840
rect 23440 29783 23463 29817
rect 23497 29783 23520 29817
rect 23440 29497 23520 29783
rect 23440 29463 23463 29497
rect 23497 29463 23520 29497
rect 23440 29440 23520 29463
rect 23600 29817 23680 29840
rect 23600 29783 23623 29817
rect 23657 29783 23680 29817
rect 23600 29497 23680 29783
rect 23600 29463 23623 29497
rect 23657 29463 23680 29497
rect 23600 29440 23680 29463
rect 23760 29817 23840 29840
rect 23760 29783 23783 29817
rect 23817 29783 23840 29817
rect 23760 29497 23840 29783
rect 23760 29463 23783 29497
rect 23817 29463 23840 29497
rect 23760 29440 23840 29463
rect 23920 29817 24000 29840
rect 23920 29783 23943 29817
rect 23977 29783 24000 29817
rect 23920 29497 24000 29783
rect 23920 29463 23943 29497
rect 23977 29463 24000 29497
rect 23920 29440 24000 29463
rect 24080 29817 24160 29840
rect 24080 29783 24103 29817
rect 24137 29783 24160 29817
rect 24080 29497 24160 29783
rect 24080 29463 24103 29497
rect 24137 29463 24160 29497
rect 24080 29440 24160 29463
rect 24240 29817 24320 29840
rect 24240 29783 24263 29817
rect 24297 29783 24320 29817
rect 24240 29497 24320 29783
rect 24240 29463 24263 29497
rect 24297 29463 24320 29497
rect 24240 29440 24320 29463
rect 24400 29817 24480 29840
rect 24400 29783 24423 29817
rect 24457 29783 24480 29817
rect 24400 29497 24480 29783
rect 24400 29463 24423 29497
rect 24457 29463 24480 29497
rect 24400 29440 24480 29463
rect 24560 29817 24640 29840
rect 24560 29783 24583 29817
rect 24617 29783 24640 29817
rect 24560 29497 24640 29783
rect 24560 29463 24583 29497
rect 24617 29463 24640 29497
rect 24560 29440 24640 29463
rect 24720 29817 24800 29840
rect 24720 29783 24743 29817
rect 24777 29783 24800 29817
rect 24720 29497 24800 29783
rect 24720 29463 24743 29497
rect 24777 29463 24800 29497
rect 24720 29440 24800 29463
rect 24880 29817 24960 29840
rect 24880 29783 24903 29817
rect 24937 29783 24960 29817
rect 24880 29497 24960 29783
rect 24880 29463 24903 29497
rect 24937 29463 24960 29497
rect 24880 29440 24960 29463
rect 25040 29817 25120 29840
rect 25040 29783 25063 29817
rect 25097 29783 25120 29817
rect 25040 29497 25120 29783
rect 25040 29463 25063 29497
rect 25097 29463 25120 29497
rect 25040 29440 25120 29463
rect 25200 29817 25280 29840
rect 25200 29783 25223 29817
rect 25257 29783 25280 29817
rect 25200 29497 25280 29783
rect 25200 29463 25223 29497
rect 25257 29463 25280 29497
rect 25200 29440 25280 29463
rect 25360 29817 25440 29840
rect 25360 29783 25383 29817
rect 25417 29783 25440 29817
rect 25360 29497 25440 29783
rect 25360 29463 25383 29497
rect 25417 29463 25440 29497
rect 25360 29440 25440 29463
rect 25520 29817 25600 29840
rect 25520 29783 25543 29817
rect 25577 29783 25600 29817
rect 25520 29497 25600 29783
rect 25520 29463 25543 29497
rect 25577 29463 25600 29497
rect 25520 29440 25600 29463
rect 25680 29817 25760 29840
rect 25680 29783 25703 29817
rect 25737 29783 25760 29817
rect 25680 29497 25760 29783
rect 25680 29463 25703 29497
rect 25737 29463 25760 29497
rect 25680 29440 25760 29463
rect 25840 29817 25920 29840
rect 25840 29783 25863 29817
rect 25897 29783 25920 29817
rect 25840 29497 25920 29783
rect 25840 29463 25863 29497
rect 25897 29463 25920 29497
rect 25840 29440 25920 29463
rect 26000 29817 26080 29840
rect 26000 29783 26023 29817
rect 26057 29783 26080 29817
rect 26000 29497 26080 29783
rect 26000 29463 26023 29497
rect 26057 29463 26080 29497
rect 26000 29440 26080 29463
rect 26160 29817 26240 29840
rect 26160 29783 26183 29817
rect 26217 29783 26240 29817
rect 26160 29497 26240 29783
rect 26160 29463 26183 29497
rect 26217 29463 26240 29497
rect 26160 29440 26240 29463
rect 26320 29817 26400 29840
rect 26320 29783 26343 29817
rect 26377 29783 26400 29817
rect 26320 29497 26400 29783
rect 26320 29463 26343 29497
rect 26377 29463 26400 29497
rect 26320 29440 26400 29463
rect 26480 29817 26560 29840
rect 26480 29783 26503 29817
rect 26537 29783 26560 29817
rect 26480 29497 26560 29783
rect 26480 29463 26503 29497
rect 26537 29463 26560 29497
rect 26480 29440 26560 29463
rect 26640 29817 26720 29840
rect 26640 29783 26663 29817
rect 26697 29783 26720 29817
rect 26640 29497 26720 29783
rect 26640 29463 26663 29497
rect 26697 29463 26720 29497
rect 26640 29440 26720 29463
rect 26800 29817 26880 29840
rect 26800 29783 26823 29817
rect 26857 29783 26880 29817
rect 26800 29497 26880 29783
rect 26800 29463 26823 29497
rect 26857 29463 26880 29497
rect 26800 29440 26880 29463
rect 26960 29817 27040 29840
rect 26960 29783 26983 29817
rect 27017 29783 27040 29817
rect 26960 29497 27040 29783
rect 26960 29463 26983 29497
rect 27017 29463 27040 29497
rect 26960 29440 27040 29463
rect 27120 29817 27200 29840
rect 27120 29783 27143 29817
rect 27177 29783 27200 29817
rect 27120 29497 27200 29783
rect 27120 29463 27143 29497
rect 27177 29463 27200 29497
rect 27120 29440 27200 29463
rect 27280 29817 27360 29840
rect 27280 29783 27303 29817
rect 27337 29783 27360 29817
rect 27280 29497 27360 29783
rect 27280 29463 27303 29497
rect 27337 29463 27360 29497
rect 27280 29440 27360 29463
rect 27440 29817 27520 29840
rect 27440 29783 27463 29817
rect 27497 29783 27520 29817
rect 27440 29497 27520 29783
rect 27440 29463 27463 29497
rect 27497 29463 27520 29497
rect 27440 29440 27520 29463
rect 27600 29817 27680 29840
rect 27600 29783 27623 29817
rect 27657 29783 27680 29817
rect 27600 29497 27680 29783
rect 27600 29463 27623 29497
rect 27657 29463 27680 29497
rect 27600 29440 27680 29463
rect 27760 29817 27840 29840
rect 27760 29783 27783 29817
rect 27817 29783 27840 29817
rect 27760 29497 27840 29783
rect 27760 29463 27783 29497
rect 27817 29463 27840 29497
rect 27760 29440 27840 29463
rect 27920 29817 28000 29840
rect 27920 29783 27943 29817
rect 27977 29783 28000 29817
rect 27920 29497 28000 29783
rect 27920 29463 27943 29497
rect 27977 29463 28000 29497
rect 27920 29440 28000 29463
rect 28080 29817 28160 29840
rect 28080 29783 28103 29817
rect 28137 29783 28160 29817
rect 28080 29497 28160 29783
rect 28080 29463 28103 29497
rect 28137 29463 28160 29497
rect 28080 29440 28160 29463
rect 28240 29817 28320 29840
rect 28240 29783 28263 29817
rect 28297 29783 28320 29817
rect 28240 29497 28320 29783
rect 28240 29463 28263 29497
rect 28297 29463 28320 29497
rect 28240 29440 28320 29463
rect 28400 29817 28480 29840
rect 28400 29783 28423 29817
rect 28457 29783 28480 29817
rect 28400 29497 28480 29783
rect 28400 29463 28423 29497
rect 28457 29463 28480 29497
rect 28400 29440 28480 29463
rect 28560 29817 28640 29840
rect 28560 29783 28583 29817
rect 28617 29783 28640 29817
rect 28560 29497 28640 29783
rect 28560 29463 28583 29497
rect 28617 29463 28640 29497
rect 28560 29440 28640 29463
rect 28720 29817 28800 29840
rect 28720 29783 28743 29817
rect 28777 29783 28800 29817
rect 28720 29497 28800 29783
rect 28720 29463 28743 29497
rect 28777 29463 28800 29497
rect 28720 29440 28800 29463
rect 28880 29817 28960 29840
rect 28880 29783 28903 29817
rect 28937 29783 28960 29817
rect 28880 29497 28960 29783
rect 28880 29463 28903 29497
rect 28937 29463 28960 29497
rect 28880 29440 28960 29463
rect 29040 29817 29120 29840
rect 29040 29783 29063 29817
rect 29097 29783 29120 29817
rect 29040 29497 29120 29783
rect 29040 29463 29063 29497
rect 29097 29463 29120 29497
rect 29040 29440 29120 29463
rect 29200 29817 29280 29840
rect 29200 29783 29223 29817
rect 29257 29783 29280 29817
rect 29200 29497 29280 29783
rect 29200 29463 29223 29497
rect 29257 29463 29280 29497
rect 29200 29440 29280 29463
rect 29360 29817 29440 29840
rect 29360 29783 29383 29817
rect 29417 29783 29440 29817
rect 29360 29497 29440 29783
rect 29360 29463 29383 29497
rect 29417 29463 29440 29497
rect 29360 29440 29440 29463
rect 29520 29440 29600 29840
rect 29680 29440 29760 29840
rect 29840 29440 29920 29840
rect 30000 29440 30080 29840
rect 30160 29440 30240 29840
rect 30320 29440 30400 29840
rect 30480 29440 30560 29840
rect 30640 29440 30720 29840
rect 30800 29440 30880 29840
rect 30960 29440 31040 29840
rect 31120 29440 31200 29840
rect 31280 29440 31360 29840
rect 31440 29440 31520 29840
rect 31600 29440 31680 29840
rect 31760 29440 31840 29840
rect 31920 29440 32000 29840
rect 32080 29440 32160 29840
rect 32240 29440 32320 29840
rect 32400 29440 32480 29840
rect 32560 29440 32640 29840
rect 32720 29440 32800 29840
rect 32880 29440 32960 29840
rect 33040 29440 33120 29840
rect 33200 29440 33280 29840
rect 33360 29440 33440 29840
rect 33520 29817 33600 29840
rect 33520 29783 33543 29817
rect 33577 29783 33600 29817
rect 33520 29497 33600 29783
rect 33520 29463 33543 29497
rect 33577 29463 33600 29497
rect 33520 29440 33600 29463
rect 33680 29817 33760 29840
rect 33680 29783 33703 29817
rect 33737 29783 33760 29817
rect 33680 29497 33760 29783
rect 33680 29463 33703 29497
rect 33737 29463 33760 29497
rect 33680 29440 33760 29463
rect 33840 29817 33920 29840
rect 33840 29783 33863 29817
rect 33897 29783 33920 29817
rect 33840 29497 33920 29783
rect 33840 29463 33863 29497
rect 33897 29463 33920 29497
rect 33840 29440 33920 29463
rect 34000 29817 34080 29840
rect 34000 29783 34023 29817
rect 34057 29783 34080 29817
rect 34000 29497 34080 29783
rect 34000 29463 34023 29497
rect 34057 29463 34080 29497
rect 34000 29440 34080 29463
rect 34160 29817 34240 29840
rect 34160 29783 34183 29817
rect 34217 29783 34240 29817
rect 34160 29497 34240 29783
rect 34160 29463 34183 29497
rect 34217 29463 34240 29497
rect 34160 29440 34240 29463
rect 34320 29817 34400 29840
rect 34320 29783 34343 29817
rect 34377 29783 34400 29817
rect 34320 29497 34400 29783
rect 34320 29463 34343 29497
rect 34377 29463 34400 29497
rect 34320 29440 34400 29463
rect 34480 29817 34560 29840
rect 34480 29783 34503 29817
rect 34537 29783 34560 29817
rect 34480 29497 34560 29783
rect 34480 29463 34503 29497
rect 34537 29463 34560 29497
rect 34480 29440 34560 29463
rect 34640 29817 34720 29840
rect 34640 29783 34663 29817
rect 34697 29783 34720 29817
rect 34640 29497 34720 29783
rect 34640 29463 34663 29497
rect 34697 29463 34720 29497
rect 34640 29440 34720 29463
rect 34800 29817 34880 29840
rect 34800 29783 34823 29817
rect 34857 29783 34880 29817
rect 34800 29497 34880 29783
rect 34800 29463 34823 29497
rect 34857 29463 34880 29497
rect 34800 29440 34880 29463
rect 34960 29817 35040 29840
rect 34960 29783 34983 29817
rect 35017 29783 35040 29817
rect 34960 29497 35040 29783
rect 34960 29463 34983 29497
rect 35017 29463 35040 29497
rect 34960 29440 35040 29463
rect 35120 29817 35200 29840
rect 35120 29783 35143 29817
rect 35177 29783 35200 29817
rect 35120 29497 35200 29783
rect 35120 29463 35143 29497
rect 35177 29463 35200 29497
rect 35120 29440 35200 29463
rect 35280 29817 35360 29840
rect 35280 29783 35303 29817
rect 35337 29783 35360 29817
rect 35280 29497 35360 29783
rect 35280 29463 35303 29497
rect 35337 29463 35360 29497
rect 35280 29440 35360 29463
rect 35440 29817 35520 29840
rect 35440 29783 35463 29817
rect 35497 29783 35520 29817
rect 35440 29497 35520 29783
rect 35440 29463 35463 29497
rect 35497 29463 35520 29497
rect 35440 29440 35520 29463
rect 35600 29817 35680 29840
rect 35600 29783 35623 29817
rect 35657 29783 35680 29817
rect 35600 29497 35680 29783
rect 35600 29463 35623 29497
rect 35657 29463 35680 29497
rect 35600 29440 35680 29463
rect 35760 29817 35840 29840
rect 35760 29783 35783 29817
rect 35817 29783 35840 29817
rect 35760 29497 35840 29783
rect 35760 29463 35783 29497
rect 35817 29463 35840 29497
rect 35760 29440 35840 29463
rect 35920 29817 36000 29840
rect 35920 29783 35943 29817
rect 35977 29783 36000 29817
rect 35920 29497 36000 29783
rect 35920 29463 35943 29497
rect 35977 29463 36000 29497
rect 35920 29440 36000 29463
rect 36080 29817 36160 29840
rect 36080 29783 36103 29817
rect 36137 29783 36160 29817
rect 36080 29497 36160 29783
rect 36080 29463 36103 29497
rect 36137 29463 36160 29497
rect 36080 29440 36160 29463
rect 36240 29817 36320 29840
rect 36240 29783 36263 29817
rect 36297 29783 36320 29817
rect 36240 29497 36320 29783
rect 36240 29463 36263 29497
rect 36297 29463 36320 29497
rect 36240 29440 36320 29463
rect 36400 29817 36480 29840
rect 36400 29783 36423 29817
rect 36457 29783 36480 29817
rect 36400 29497 36480 29783
rect 36400 29463 36423 29497
rect 36457 29463 36480 29497
rect 36400 29440 36480 29463
rect 36560 29817 36640 29840
rect 36560 29783 36583 29817
rect 36617 29783 36640 29817
rect 36560 29497 36640 29783
rect 36560 29463 36583 29497
rect 36617 29463 36640 29497
rect 36560 29440 36640 29463
rect 36720 29817 36800 29840
rect 36720 29783 36743 29817
rect 36777 29783 36800 29817
rect 36720 29497 36800 29783
rect 36720 29463 36743 29497
rect 36777 29463 36800 29497
rect 36720 29440 36800 29463
rect 36880 29817 36960 29840
rect 36880 29783 36903 29817
rect 36937 29783 36960 29817
rect 36880 29497 36960 29783
rect 36880 29463 36903 29497
rect 36937 29463 36960 29497
rect 36880 29440 36960 29463
rect 37040 29817 37120 29840
rect 37040 29783 37063 29817
rect 37097 29783 37120 29817
rect 37040 29497 37120 29783
rect 37040 29463 37063 29497
rect 37097 29463 37120 29497
rect 37040 29440 37120 29463
rect 37200 29817 37280 29840
rect 37200 29783 37223 29817
rect 37257 29783 37280 29817
rect 37200 29497 37280 29783
rect 37200 29463 37223 29497
rect 37257 29463 37280 29497
rect 37200 29440 37280 29463
rect 37360 29817 37440 29840
rect 37360 29783 37383 29817
rect 37417 29783 37440 29817
rect 37360 29497 37440 29783
rect 37360 29463 37383 29497
rect 37417 29463 37440 29497
rect 37360 29440 37440 29463
rect 37520 29817 37600 29840
rect 37520 29783 37543 29817
rect 37577 29783 37600 29817
rect 37520 29497 37600 29783
rect 37520 29463 37543 29497
rect 37577 29463 37600 29497
rect 37520 29440 37600 29463
rect 37680 29817 37760 29840
rect 37680 29783 37703 29817
rect 37737 29783 37760 29817
rect 37680 29497 37760 29783
rect 37680 29463 37703 29497
rect 37737 29463 37760 29497
rect 37680 29440 37760 29463
rect 37840 29817 37920 29840
rect 37840 29783 37863 29817
rect 37897 29783 37920 29817
rect 37840 29497 37920 29783
rect 37840 29463 37863 29497
rect 37897 29463 37920 29497
rect 37840 29440 37920 29463
rect 38000 29817 38080 29840
rect 38000 29783 38023 29817
rect 38057 29783 38080 29817
rect 38000 29497 38080 29783
rect 38000 29463 38023 29497
rect 38057 29463 38080 29497
rect 38000 29440 38080 29463
rect 38160 29817 38240 29840
rect 38160 29783 38183 29817
rect 38217 29783 38240 29817
rect 38160 29497 38240 29783
rect 38160 29463 38183 29497
rect 38217 29463 38240 29497
rect 38160 29440 38240 29463
rect 38320 29817 38400 29840
rect 38320 29783 38343 29817
rect 38377 29783 38400 29817
rect 38320 29497 38400 29783
rect 38320 29463 38343 29497
rect 38377 29463 38400 29497
rect 38320 29440 38400 29463
rect 38480 29817 38560 29840
rect 38480 29783 38503 29817
rect 38537 29783 38560 29817
rect 38480 29497 38560 29783
rect 38480 29463 38503 29497
rect 38537 29463 38560 29497
rect 38480 29440 38560 29463
rect 38640 29817 38720 29840
rect 38640 29783 38663 29817
rect 38697 29783 38720 29817
rect 38640 29497 38720 29783
rect 38640 29463 38663 29497
rect 38697 29463 38720 29497
rect 38640 29440 38720 29463
rect 38800 29817 38880 29840
rect 38800 29783 38823 29817
rect 38857 29783 38880 29817
rect 38800 29497 38880 29783
rect 38800 29463 38823 29497
rect 38857 29463 38880 29497
rect 38800 29440 38880 29463
rect 38960 29817 39040 29840
rect 38960 29783 38983 29817
rect 39017 29783 39040 29817
rect 38960 29497 39040 29783
rect 38960 29463 38983 29497
rect 39017 29463 39040 29497
rect 38960 29440 39040 29463
rect 39120 29817 39200 29840
rect 39120 29783 39143 29817
rect 39177 29783 39200 29817
rect 39120 29497 39200 29783
rect 39120 29463 39143 29497
rect 39177 29463 39200 29497
rect 39120 29440 39200 29463
rect 39280 29817 39360 29840
rect 39280 29783 39303 29817
rect 39337 29783 39360 29817
rect 39280 29497 39360 29783
rect 39280 29463 39303 29497
rect 39337 29463 39360 29497
rect 39280 29440 39360 29463
rect 39440 29817 39520 29840
rect 39440 29783 39463 29817
rect 39497 29783 39520 29817
rect 39440 29497 39520 29783
rect 39440 29463 39463 29497
rect 39497 29463 39520 29497
rect 39440 29440 39520 29463
rect 39600 29817 39680 29840
rect 39600 29783 39623 29817
rect 39657 29783 39680 29817
rect 39600 29497 39680 29783
rect 39600 29463 39623 29497
rect 39657 29463 39680 29497
rect 39600 29440 39680 29463
rect 39760 29817 39840 29840
rect 39760 29783 39783 29817
rect 39817 29783 39840 29817
rect 39760 29497 39840 29783
rect 39760 29463 39783 29497
rect 39817 29463 39840 29497
rect 39760 29440 39840 29463
rect 39920 29817 40000 29840
rect 39920 29783 39943 29817
rect 39977 29783 40000 29817
rect 39920 29497 40000 29783
rect 39920 29463 39943 29497
rect 39977 29463 40000 29497
rect 39920 29440 40000 29463
rect 40080 29817 40160 29840
rect 40080 29783 40103 29817
rect 40137 29783 40160 29817
rect 40080 29497 40160 29783
rect 40080 29463 40103 29497
rect 40137 29463 40160 29497
rect 40080 29440 40160 29463
rect 40240 29817 40320 29840
rect 40240 29783 40263 29817
rect 40297 29783 40320 29817
rect 40240 29497 40320 29783
rect 40240 29463 40263 29497
rect 40297 29463 40320 29497
rect 40240 29440 40320 29463
rect 40400 29817 40480 29840
rect 40400 29783 40423 29817
rect 40457 29783 40480 29817
rect 40400 29497 40480 29783
rect 40400 29463 40423 29497
rect 40457 29463 40480 29497
rect 40400 29440 40480 29463
rect 40560 29817 40640 29840
rect 40560 29783 40583 29817
rect 40617 29783 40640 29817
rect 40560 29497 40640 29783
rect 40560 29463 40583 29497
rect 40617 29463 40640 29497
rect 40560 29440 40640 29463
rect 40720 29817 40800 29840
rect 40720 29783 40743 29817
rect 40777 29783 40800 29817
rect 40720 29497 40800 29783
rect 40720 29463 40743 29497
rect 40777 29463 40800 29497
rect 40720 29440 40800 29463
rect 40880 29817 40960 29840
rect 40880 29783 40903 29817
rect 40937 29783 40960 29817
rect 40880 29497 40960 29783
rect 40880 29463 40903 29497
rect 40937 29463 40960 29497
rect 40880 29440 40960 29463
rect 41040 29817 41120 29840
rect 41040 29783 41063 29817
rect 41097 29783 41120 29817
rect 41040 29497 41120 29783
rect 41040 29463 41063 29497
rect 41097 29463 41120 29497
rect 41040 29440 41120 29463
rect 41200 29817 41280 29840
rect 41200 29783 41223 29817
rect 41257 29783 41280 29817
rect 41200 29497 41280 29783
rect 41200 29463 41223 29497
rect 41257 29463 41280 29497
rect 41200 29440 41280 29463
rect 41360 29817 41440 29840
rect 41360 29783 41383 29817
rect 41417 29783 41440 29817
rect 41360 29497 41440 29783
rect 41360 29463 41383 29497
rect 41417 29463 41440 29497
rect 41360 29440 41440 29463
rect 41520 29817 41600 29840
rect 41520 29783 41543 29817
rect 41577 29783 41600 29817
rect 41520 29497 41600 29783
rect 41520 29463 41543 29497
rect 41577 29463 41600 29497
rect 41520 29440 41600 29463
rect 41680 29817 41760 29840
rect 41680 29783 41703 29817
rect 41737 29783 41760 29817
rect 41680 29497 41760 29783
rect 41680 29463 41703 29497
rect 41737 29463 41760 29497
rect 41680 29440 41760 29463
rect 41840 29817 41920 29840
rect 41840 29783 41863 29817
rect 41897 29783 41920 29817
rect 41840 29497 41920 29783
rect 41840 29463 41863 29497
rect 41897 29463 41920 29497
rect 41840 29440 41920 29463
<< viali >>
rect 23 37303 57 37337
rect 23 36983 57 37017
rect 183 37303 217 37337
rect 183 36983 217 37017
rect 343 37303 377 37337
rect 343 36983 377 37017
rect 503 37303 537 37337
rect 503 36983 537 37017
rect 663 37303 697 37337
rect 663 36983 697 37017
rect 823 37303 857 37337
rect 823 36983 857 37017
rect 983 37303 1017 37337
rect 983 36983 1017 37017
rect 1143 37303 1177 37337
rect 1143 36983 1177 37017
rect 1303 37303 1337 37337
rect 1303 36983 1337 37017
rect 1463 37303 1497 37337
rect 1463 36983 1497 37017
rect 1623 37303 1657 37337
rect 1623 36983 1657 37017
rect 1783 37303 1817 37337
rect 1783 36983 1817 37017
rect 1943 37303 1977 37337
rect 1943 36983 1977 37017
rect 2103 37303 2137 37337
rect 2103 36983 2137 37017
rect 2263 37303 2297 37337
rect 2263 36983 2297 37017
rect 2423 37303 2457 37337
rect 2423 36983 2457 37017
rect 2583 37303 2617 37337
rect 2583 36983 2617 37017
rect 2743 37303 2777 37337
rect 2743 36983 2777 37017
rect 2903 37303 2937 37337
rect 2903 36983 2937 37017
rect 3063 37303 3097 37337
rect 3063 36983 3097 37017
rect 3223 37303 3257 37337
rect 3223 36983 3257 37017
rect 3383 37303 3417 37337
rect 3383 36983 3417 37017
rect 3543 37303 3577 37337
rect 3543 36983 3577 37017
rect 3703 37303 3737 37337
rect 3703 36983 3737 37017
rect 3863 37303 3897 37337
rect 3863 36983 3897 37017
rect 4023 37303 4057 37337
rect 4023 36983 4057 37017
rect 4183 37303 4217 37337
rect 4183 36983 4217 37017
rect 4343 37303 4377 37337
rect 4343 36983 4377 37017
rect 4503 37303 4537 37337
rect 4503 36983 4537 37017
rect 4663 37303 4697 37337
rect 4663 36983 4697 37017
rect 4823 37303 4857 37337
rect 4823 36983 4857 37017
rect 4983 37303 5017 37337
rect 4983 36983 5017 37017
rect 5143 37303 5177 37337
rect 5143 36983 5177 37017
rect 5303 37303 5337 37337
rect 5303 36983 5337 37017
rect 5463 37303 5497 37337
rect 5463 36983 5497 37017
rect 5623 37303 5657 37337
rect 5623 36983 5657 37017
rect 5783 37303 5817 37337
rect 5783 36983 5817 37017
rect 5943 37303 5977 37337
rect 5943 36983 5977 37017
rect 6103 37303 6137 37337
rect 6103 36983 6137 37017
rect 6263 37303 6297 37337
rect 6263 36983 6297 37017
rect 6423 37303 6457 37337
rect 6423 36983 6457 37017
rect 6583 37303 6617 37337
rect 6583 36983 6617 37017
rect 6743 37303 6777 37337
rect 6743 36983 6777 37017
rect 6903 37303 6937 37337
rect 6903 36983 6937 37017
rect 7063 37303 7097 37337
rect 7063 36983 7097 37017
rect 7223 37303 7257 37337
rect 7223 36983 7257 37017
rect 7383 37303 7417 37337
rect 7383 36983 7417 37017
rect 7543 37303 7577 37337
rect 7543 36983 7577 37017
rect 7703 37303 7737 37337
rect 7703 36983 7737 37017
rect 7863 37303 7897 37337
rect 7863 36983 7897 37017
rect 8023 37303 8057 37337
rect 8023 36983 8057 37017
rect 8183 37303 8217 37337
rect 8183 36983 8217 37017
rect 8343 37303 8377 37337
rect 8343 36983 8377 37017
rect 12503 37303 12537 37337
rect 12503 36983 12537 37017
rect 12663 37303 12697 37337
rect 12663 36983 12697 37017
rect 12823 37303 12857 37337
rect 12823 36983 12857 37017
rect 12983 37303 13017 37337
rect 12983 36983 13017 37017
rect 13143 37303 13177 37337
rect 13143 36983 13177 37017
rect 13303 37303 13337 37337
rect 13303 36983 13337 37017
rect 13463 37303 13497 37337
rect 13463 36983 13497 37017
rect 13623 37303 13657 37337
rect 13623 36983 13657 37017
rect 13783 37303 13817 37337
rect 13783 36983 13817 37017
rect 13943 37303 13977 37337
rect 13943 36983 13977 37017
rect 14103 37303 14137 37337
rect 14103 36983 14137 37017
rect 14263 37303 14297 37337
rect 14263 36983 14297 37017
rect 14423 37303 14457 37337
rect 14423 36983 14457 37017
rect 14583 37303 14617 37337
rect 14583 36983 14617 37017
rect 14743 37303 14777 37337
rect 14743 36983 14777 37017
rect 14903 37303 14937 37337
rect 14903 36983 14937 37017
rect 15063 37303 15097 37337
rect 15063 36983 15097 37017
rect 15223 37303 15257 37337
rect 15223 36983 15257 37017
rect 15383 37303 15417 37337
rect 15383 36983 15417 37017
rect 15543 37303 15577 37337
rect 15543 36983 15577 37017
rect 15703 37303 15737 37337
rect 15703 36983 15737 37017
rect 15863 37303 15897 37337
rect 15863 36983 15897 37017
rect 16023 37303 16057 37337
rect 16023 36983 16057 37017
rect 16183 37303 16217 37337
rect 16183 36983 16217 37017
rect 16343 37303 16377 37337
rect 16343 36983 16377 37017
rect 16503 37303 16537 37337
rect 16503 36983 16537 37017
rect 16663 37303 16697 37337
rect 16663 36983 16697 37017
rect 16823 37303 16857 37337
rect 16823 36983 16857 37017
rect 16983 37303 17017 37337
rect 16983 36983 17017 37017
rect 17143 37303 17177 37337
rect 17143 36983 17177 37017
rect 17303 37303 17337 37337
rect 17303 36983 17337 37017
rect 17463 37303 17497 37337
rect 17463 36983 17497 37017
rect 17623 37303 17657 37337
rect 17623 36983 17657 37017
rect 17783 37303 17817 37337
rect 17783 36983 17817 37017
rect 17943 37303 17977 37337
rect 17943 36983 17977 37017
rect 18103 37303 18137 37337
rect 18103 36983 18137 37017
rect 18263 37303 18297 37337
rect 18263 36983 18297 37017
rect 18423 37303 18457 37337
rect 18423 36983 18457 37017
rect 18583 37303 18617 37337
rect 18583 36983 18617 37017
rect 18743 37303 18777 37337
rect 18743 36983 18777 37017
rect 18903 37303 18937 37337
rect 18903 36983 18937 37017
rect 23143 37303 23177 37337
rect 23143 36983 23177 37017
rect 23303 37303 23337 37337
rect 23303 36983 23337 37017
rect 23463 37303 23497 37337
rect 23463 36983 23497 37017
rect 23623 37303 23657 37337
rect 23623 36983 23657 37017
rect 23783 37303 23817 37337
rect 23783 36983 23817 37017
rect 23943 37303 23977 37337
rect 23943 36983 23977 37017
rect 24103 37303 24137 37337
rect 24103 36983 24137 37017
rect 24263 37303 24297 37337
rect 24263 36983 24297 37017
rect 24423 37303 24457 37337
rect 24423 36983 24457 37017
rect 24583 37303 24617 37337
rect 24583 36983 24617 37017
rect 24743 37303 24777 37337
rect 24743 36983 24777 37017
rect 24903 37303 24937 37337
rect 24903 36983 24937 37017
rect 25063 37303 25097 37337
rect 25063 36983 25097 37017
rect 25223 37303 25257 37337
rect 25223 36983 25257 37017
rect 25383 37303 25417 37337
rect 25383 36983 25417 37017
rect 25543 37303 25577 37337
rect 25543 36983 25577 37017
rect 25703 37303 25737 37337
rect 25703 36983 25737 37017
rect 25863 37303 25897 37337
rect 25863 36983 25897 37017
rect 26023 37303 26057 37337
rect 26023 36983 26057 37017
rect 26183 37303 26217 37337
rect 26183 36983 26217 37017
rect 26343 37303 26377 37337
rect 26343 36983 26377 37017
rect 26503 37303 26537 37337
rect 26503 36983 26537 37017
rect 26663 37303 26697 37337
rect 26663 36983 26697 37017
rect 26823 37303 26857 37337
rect 26823 36983 26857 37017
rect 26983 37303 27017 37337
rect 26983 36983 27017 37017
rect 27143 37303 27177 37337
rect 27143 36983 27177 37017
rect 27303 37303 27337 37337
rect 27303 36983 27337 37017
rect 27463 37303 27497 37337
rect 27463 36983 27497 37017
rect 27623 37303 27657 37337
rect 27623 36983 27657 37017
rect 27783 37303 27817 37337
rect 27783 36983 27817 37017
rect 27943 37303 27977 37337
rect 27943 36983 27977 37017
rect 28103 37303 28137 37337
rect 28103 36983 28137 37017
rect 28263 37303 28297 37337
rect 28263 36983 28297 37017
rect 28423 37303 28457 37337
rect 28423 36983 28457 37017
rect 28583 37303 28617 37337
rect 28583 36983 28617 37017
rect 28743 37303 28777 37337
rect 28743 36983 28777 37017
rect 28903 37303 28937 37337
rect 28903 36983 28937 37017
rect 29063 37303 29097 37337
rect 29063 36983 29097 37017
rect 29223 37303 29257 37337
rect 29223 36983 29257 37017
rect 29383 37303 29417 37337
rect 29383 36983 29417 37017
rect 33543 37303 33577 37337
rect 33543 36983 33577 37017
rect 33703 37303 33737 37337
rect 33703 36983 33737 37017
rect 33863 37303 33897 37337
rect 33863 36983 33897 37017
rect 34023 37303 34057 37337
rect 34023 36983 34057 37017
rect 34183 37303 34217 37337
rect 34183 36983 34217 37017
rect 34343 37303 34377 37337
rect 34343 36983 34377 37017
rect 34503 37303 34537 37337
rect 34503 36983 34537 37017
rect 34663 37303 34697 37337
rect 34663 36983 34697 37017
rect 34823 37303 34857 37337
rect 34823 36983 34857 37017
rect 34983 37303 35017 37337
rect 34983 36983 35017 37017
rect 35143 37303 35177 37337
rect 35143 36983 35177 37017
rect 35303 37303 35337 37337
rect 35303 36983 35337 37017
rect 35463 37303 35497 37337
rect 35463 36983 35497 37017
rect 35623 37303 35657 37337
rect 35623 36983 35657 37017
rect 35783 37303 35817 37337
rect 35783 36983 35817 37017
rect 35943 37303 35977 37337
rect 35943 36983 35977 37017
rect 36103 37303 36137 37337
rect 36103 36983 36137 37017
rect 36263 37303 36297 37337
rect 36263 36983 36297 37017
rect 36423 37303 36457 37337
rect 36423 36983 36457 37017
rect 36583 37303 36617 37337
rect 36583 36983 36617 37017
rect 36743 37303 36777 37337
rect 36743 36983 36777 37017
rect 36903 37303 36937 37337
rect 36903 36983 36937 37017
rect 37063 37303 37097 37337
rect 37063 36983 37097 37017
rect 37223 37303 37257 37337
rect 37223 36983 37257 37017
rect 37383 37303 37417 37337
rect 37383 36983 37417 37017
rect 37543 37303 37577 37337
rect 37543 36983 37577 37017
rect 37703 37303 37737 37337
rect 37703 36983 37737 37017
rect 37863 37303 37897 37337
rect 37863 36983 37897 37017
rect 38023 37303 38057 37337
rect 38023 36983 38057 37017
rect 38183 37303 38217 37337
rect 38183 36983 38217 37017
rect 38343 37303 38377 37337
rect 38343 36983 38377 37017
rect 38503 37303 38537 37337
rect 38503 36983 38537 37017
rect 38663 37303 38697 37337
rect 38663 36983 38697 37017
rect 38823 37303 38857 37337
rect 38823 36983 38857 37017
rect 38983 37303 39017 37337
rect 38983 36983 39017 37017
rect 39143 37303 39177 37337
rect 39143 36983 39177 37017
rect 39303 37303 39337 37337
rect 39303 36983 39337 37017
rect 39463 37303 39497 37337
rect 39463 36983 39497 37017
rect 39623 37303 39657 37337
rect 39623 36983 39657 37017
rect 39783 37303 39817 37337
rect 39783 36983 39817 37017
rect 39943 37303 39977 37337
rect 39943 36983 39977 37017
rect 40103 37303 40137 37337
rect 40103 36983 40137 37017
rect 40263 37303 40297 37337
rect 40263 36983 40297 37017
rect 40423 37303 40457 37337
rect 40423 36983 40457 37017
rect 40583 37303 40617 37337
rect 40583 36983 40617 37017
rect 40743 37303 40777 37337
rect 40743 36983 40777 37017
rect 40903 37303 40937 37337
rect 40903 36983 40937 37017
rect 41063 37303 41097 37337
rect 41063 36983 41097 37017
rect 41223 37303 41257 37337
rect 41223 36983 41257 37017
rect 41383 37303 41417 37337
rect 41383 36983 41417 37017
rect 41543 37303 41577 37337
rect 41543 36983 41577 37017
rect 41703 37303 41737 37337
rect 41703 36983 41737 37017
rect 41863 37303 41897 37337
rect 41863 36983 41897 37017
rect 23 36823 57 36857
rect 23 36503 57 36537
rect 183 36823 217 36857
rect 183 36503 217 36537
rect 343 36823 377 36857
rect 343 36503 377 36537
rect 503 36823 537 36857
rect 503 36503 537 36537
rect 663 36823 697 36857
rect 663 36503 697 36537
rect 823 36823 857 36857
rect 823 36503 857 36537
rect 983 36823 1017 36857
rect 983 36503 1017 36537
rect 1143 36823 1177 36857
rect 1143 36503 1177 36537
rect 1303 36823 1337 36857
rect 1303 36503 1337 36537
rect 1463 36823 1497 36857
rect 1463 36503 1497 36537
rect 1623 36823 1657 36857
rect 1623 36503 1657 36537
rect 1783 36823 1817 36857
rect 1783 36503 1817 36537
rect 1943 36823 1977 36857
rect 1943 36503 1977 36537
rect 2103 36823 2137 36857
rect 2103 36503 2137 36537
rect 2263 36823 2297 36857
rect 2263 36503 2297 36537
rect 2423 36823 2457 36857
rect 2423 36503 2457 36537
rect 2583 36823 2617 36857
rect 2583 36503 2617 36537
rect 2743 36823 2777 36857
rect 2743 36503 2777 36537
rect 2903 36823 2937 36857
rect 2903 36503 2937 36537
rect 3063 36823 3097 36857
rect 3063 36503 3097 36537
rect 3223 36823 3257 36857
rect 3223 36503 3257 36537
rect 3383 36823 3417 36857
rect 3383 36503 3417 36537
rect 3543 36823 3577 36857
rect 3543 36503 3577 36537
rect 3703 36823 3737 36857
rect 3703 36503 3737 36537
rect 3863 36823 3897 36857
rect 3863 36503 3897 36537
rect 4023 36823 4057 36857
rect 4023 36503 4057 36537
rect 4183 36823 4217 36857
rect 4183 36503 4217 36537
rect 4343 36823 4377 36857
rect 4343 36503 4377 36537
rect 4503 36823 4537 36857
rect 4503 36503 4537 36537
rect 4663 36823 4697 36857
rect 4663 36503 4697 36537
rect 4823 36823 4857 36857
rect 4823 36503 4857 36537
rect 4983 36823 5017 36857
rect 4983 36503 5017 36537
rect 5143 36823 5177 36857
rect 5143 36503 5177 36537
rect 5303 36823 5337 36857
rect 5303 36503 5337 36537
rect 5463 36823 5497 36857
rect 5463 36503 5497 36537
rect 5623 36823 5657 36857
rect 5623 36503 5657 36537
rect 5783 36823 5817 36857
rect 5783 36503 5817 36537
rect 5943 36823 5977 36857
rect 5943 36503 5977 36537
rect 6103 36823 6137 36857
rect 6103 36503 6137 36537
rect 6263 36823 6297 36857
rect 6263 36503 6297 36537
rect 6423 36823 6457 36857
rect 6423 36503 6457 36537
rect 6583 36823 6617 36857
rect 6583 36503 6617 36537
rect 6743 36823 6777 36857
rect 6743 36503 6777 36537
rect 6903 36823 6937 36857
rect 6903 36503 6937 36537
rect 7063 36823 7097 36857
rect 7063 36503 7097 36537
rect 7223 36823 7257 36857
rect 7223 36503 7257 36537
rect 7383 36823 7417 36857
rect 7383 36503 7417 36537
rect 7543 36823 7577 36857
rect 7543 36503 7577 36537
rect 7703 36823 7737 36857
rect 7703 36503 7737 36537
rect 7863 36823 7897 36857
rect 7863 36503 7897 36537
rect 8023 36823 8057 36857
rect 8023 36503 8057 36537
rect 8183 36823 8217 36857
rect 8183 36503 8217 36537
rect 8343 36823 8377 36857
rect 8343 36503 8377 36537
rect 12503 36823 12537 36857
rect 12503 36503 12537 36537
rect 12663 36823 12697 36857
rect 12663 36503 12697 36537
rect 12823 36823 12857 36857
rect 12823 36503 12857 36537
rect 12983 36823 13017 36857
rect 12983 36503 13017 36537
rect 13143 36823 13177 36857
rect 13143 36503 13177 36537
rect 13303 36823 13337 36857
rect 13303 36503 13337 36537
rect 13463 36823 13497 36857
rect 13463 36503 13497 36537
rect 13623 36823 13657 36857
rect 13623 36503 13657 36537
rect 13783 36823 13817 36857
rect 13783 36503 13817 36537
rect 13943 36823 13977 36857
rect 13943 36503 13977 36537
rect 14103 36823 14137 36857
rect 14103 36503 14137 36537
rect 14263 36823 14297 36857
rect 14263 36503 14297 36537
rect 14423 36823 14457 36857
rect 14423 36503 14457 36537
rect 14583 36823 14617 36857
rect 14583 36503 14617 36537
rect 14743 36823 14777 36857
rect 14743 36503 14777 36537
rect 14903 36823 14937 36857
rect 14903 36503 14937 36537
rect 15063 36823 15097 36857
rect 15063 36503 15097 36537
rect 15223 36823 15257 36857
rect 15223 36503 15257 36537
rect 15383 36823 15417 36857
rect 15383 36503 15417 36537
rect 15543 36823 15577 36857
rect 15543 36503 15577 36537
rect 15703 36823 15737 36857
rect 15703 36503 15737 36537
rect 15863 36823 15897 36857
rect 15863 36503 15897 36537
rect 16023 36823 16057 36857
rect 16023 36503 16057 36537
rect 16183 36823 16217 36857
rect 16183 36503 16217 36537
rect 16343 36823 16377 36857
rect 16343 36503 16377 36537
rect 16503 36823 16537 36857
rect 16503 36503 16537 36537
rect 16663 36823 16697 36857
rect 16663 36503 16697 36537
rect 16823 36823 16857 36857
rect 16823 36503 16857 36537
rect 16983 36823 17017 36857
rect 16983 36503 17017 36537
rect 17143 36823 17177 36857
rect 17143 36503 17177 36537
rect 17303 36823 17337 36857
rect 17303 36503 17337 36537
rect 17463 36823 17497 36857
rect 17463 36503 17497 36537
rect 17623 36823 17657 36857
rect 17623 36503 17657 36537
rect 17783 36823 17817 36857
rect 17783 36503 17817 36537
rect 17943 36823 17977 36857
rect 17943 36503 17977 36537
rect 18103 36823 18137 36857
rect 18103 36503 18137 36537
rect 18263 36823 18297 36857
rect 18263 36503 18297 36537
rect 18423 36823 18457 36857
rect 18423 36503 18457 36537
rect 18583 36823 18617 36857
rect 18583 36503 18617 36537
rect 18743 36823 18777 36857
rect 18743 36503 18777 36537
rect 18903 36823 18937 36857
rect 18903 36503 18937 36537
rect 23143 36823 23177 36857
rect 23143 36503 23177 36537
rect 23303 36823 23337 36857
rect 23303 36503 23337 36537
rect 23463 36823 23497 36857
rect 23463 36503 23497 36537
rect 23623 36823 23657 36857
rect 23623 36503 23657 36537
rect 23783 36823 23817 36857
rect 23783 36503 23817 36537
rect 23943 36823 23977 36857
rect 23943 36503 23977 36537
rect 24103 36823 24137 36857
rect 24103 36503 24137 36537
rect 24263 36823 24297 36857
rect 24263 36503 24297 36537
rect 24423 36823 24457 36857
rect 24423 36503 24457 36537
rect 24583 36823 24617 36857
rect 24583 36503 24617 36537
rect 24743 36823 24777 36857
rect 24743 36503 24777 36537
rect 24903 36823 24937 36857
rect 24903 36503 24937 36537
rect 25063 36823 25097 36857
rect 25063 36503 25097 36537
rect 25223 36823 25257 36857
rect 25223 36503 25257 36537
rect 25383 36823 25417 36857
rect 25383 36503 25417 36537
rect 25543 36823 25577 36857
rect 25543 36503 25577 36537
rect 25703 36823 25737 36857
rect 25703 36503 25737 36537
rect 25863 36823 25897 36857
rect 25863 36503 25897 36537
rect 26023 36823 26057 36857
rect 26023 36503 26057 36537
rect 26183 36823 26217 36857
rect 26183 36503 26217 36537
rect 26343 36823 26377 36857
rect 26343 36503 26377 36537
rect 26503 36823 26537 36857
rect 26503 36503 26537 36537
rect 26663 36823 26697 36857
rect 26663 36503 26697 36537
rect 26823 36823 26857 36857
rect 26823 36503 26857 36537
rect 26983 36823 27017 36857
rect 26983 36503 27017 36537
rect 27143 36823 27177 36857
rect 27143 36503 27177 36537
rect 27303 36823 27337 36857
rect 27303 36503 27337 36537
rect 27463 36823 27497 36857
rect 27463 36503 27497 36537
rect 27623 36823 27657 36857
rect 27623 36503 27657 36537
rect 27783 36823 27817 36857
rect 27783 36503 27817 36537
rect 27943 36823 27977 36857
rect 27943 36503 27977 36537
rect 28103 36823 28137 36857
rect 28103 36503 28137 36537
rect 28263 36823 28297 36857
rect 28263 36503 28297 36537
rect 28423 36823 28457 36857
rect 28423 36503 28457 36537
rect 28583 36823 28617 36857
rect 28583 36503 28617 36537
rect 28743 36823 28777 36857
rect 28743 36503 28777 36537
rect 28903 36823 28937 36857
rect 28903 36503 28937 36537
rect 29063 36823 29097 36857
rect 29063 36503 29097 36537
rect 29223 36823 29257 36857
rect 29223 36503 29257 36537
rect 29383 36823 29417 36857
rect 29383 36503 29417 36537
rect 33543 36823 33577 36857
rect 33543 36503 33577 36537
rect 33703 36823 33737 36857
rect 33703 36503 33737 36537
rect 33863 36823 33897 36857
rect 33863 36503 33897 36537
rect 34023 36823 34057 36857
rect 34023 36503 34057 36537
rect 34183 36823 34217 36857
rect 34183 36503 34217 36537
rect 34343 36823 34377 36857
rect 34343 36503 34377 36537
rect 34503 36823 34537 36857
rect 34503 36503 34537 36537
rect 34663 36823 34697 36857
rect 34663 36503 34697 36537
rect 34823 36823 34857 36857
rect 34823 36503 34857 36537
rect 34983 36823 35017 36857
rect 34983 36503 35017 36537
rect 35143 36823 35177 36857
rect 35143 36503 35177 36537
rect 35303 36823 35337 36857
rect 35303 36503 35337 36537
rect 35463 36823 35497 36857
rect 35463 36503 35497 36537
rect 35623 36823 35657 36857
rect 35623 36503 35657 36537
rect 35783 36823 35817 36857
rect 35783 36503 35817 36537
rect 35943 36823 35977 36857
rect 35943 36503 35977 36537
rect 36103 36823 36137 36857
rect 36103 36503 36137 36537
rect 36263 36823 36297 36857
rect 36263 36503 36297 36537
rect 36423 36823 36457 36857
rect 36423 36503 36457 36537
rect 36583 36823 36617 36857
rect 36583 36503 36617 36537
rect 36743 36823 36777 36857
rect 36743 36503 36777 36537
rect 36903 36823 36937 36857
rect 36903 36503 36937 36537
rect 37063 36823 37097 36857
rect 37063 36503 37097 36537
rect 37223 36823 37257 36857
rect 37223 36503 37257 36537
rect 37383 36823 37417 36857
rect 37383 36503 37417 36537
rect 37543 36823 37577 36857
rect 37543 36503 37577 36537
rect 37703 36823 37737 36857
rect 37703 36503 37737 36537
rect 37863 36823 37897 36857
rect 37863 36503 37897 36537
rect 38023 36823 38057 36857
rect 38023 36503 38057 36537
rect 38183 36823 38217 36857
rect 38183 36503 38217 36537
rect 38343 36823 38377 36857
rect 38343 36503 38377 36537
rect 38503 36823 38537 36857
rect 38503 36503 38537 36537
rect 38663 36823 38697 36857
rect 38663 36503 38697 36537
rect 38823 36823 38857 36857
rect 38823 36503 38857 36537
rect 38983 36823 39017 36857
rect 38983 36503 39017 36537
rect 39143 36823 39177 36857
rect 39143 36503 39177 36537
rect 39303 36823 39337 36857
rect 39303 36503 39337 36537
rect 39463 36823 39497 36857
rect 39463 36503 39497 36537
rect 39623 36823 39657 36857
rect 39623 36503 39657 36537
rect 39783 36823 39817 36857
rect 39783 36503 39817 36537
rect 39943 36823 39977 36857
rect 39943 36503 39977 36537
rect 40103 36823 40137 36857
rect 40103 36503 40137 36537
rect 40263 36823 40297 36857
rect 40263 36503 40297 36537
rect 40423 36823 40457 36857
rect 40423 36503 40457 36537
rect 40583 36823 40617 36857
rect 40583 36503 40617 36537
rect 40743 36823 40777 36857
rect 40743 36503 40777 36537
rect 40903 36823 40937 36857
rect 40903 36503 40937 36537
rect 41063 36823 41097 36857
rect 41063 36503 41097 36537
rect 41223 36823 41257 36857
rect 41223 36503 41257 36537
rect 41383 36823 41417 36857
rect 41383 36503 41417 36537
rect 41543 36823 41577 36857
rect 41543 36503 41577 36537
rect 41703 36823 41737 36857
rect 41703 36503 41737 36537
rect 41863 36823 41897 36857
rect 41863 36503 41897 36537
rect 23 36343 57 36377
rect 23 36023 57 36057
rect 23 35703 57 35737
rect 23 35383 57 35417
rect 23 35063 57 35097
rect 23 34743 57 34777
rect 23 34423 57 34457
rect 183 36343 217 36377
rect 183 36023 217 36057
rect 183 35703 217 35737
rect 183 35383 217 35417
rect 183 35063 217 35097
rect 183 34743 217 34777
rect 183 34423 217 34457
rect 343 36343 377 36377
rect 343 36023 377 36057
rect 343 35703 377 35737
rect 343 35383 377 35417
rect 343 35063 377 35097
rect 343 34743 377 34777
rect 343 34423 377 34457
rect 503 36343 537 36377
rect 503 36023 537 36057
rect 503 35703 537 35737
rect 503 35383 537 35417
rect 503 35063 537 35097
rect 503 34743 537 34777
rect 503 34423 537 34457
rect 663 36343 697 36377
rect 663 36023 697 36057
rect 663 35703 697 35737
rect 663 35383 697 35417
rect 663 35063 697 35097
rect 663 34743 697 34777
rect 663 34423 697 34457
rect 823 36343 857 36377
rect 823 36023 857 36057
rect 823 35703 857 35737
rect 823 35383 857 35417
rect 823 35063 857 35097
rect 823 34743 857 34777
rect 823 34423 857 34457
rect 983 36343 1017 36377
rect 983 36023 1017 36057
rect 983 35703 1017 35737
rect 983 35383 1017 35417
rect 983 35063 1017 35097
rect 983 34743 1017 34777
rect 983 34423 1017 34457
rect 1143 36343 1177 36377
rect 1143 36023 1177 36057
rect 1143 35703 1177 35737
rect 1143 35383 1177 35417
rect 1143 35063 1177 35097
rect 1143 34743 1177 34777
rect 1143 34423 1177 34457
rect 1303 36343 1337 36377
rect 1303 36023 1337 36057
rect 1303 35703 1337 35737
rect 1303 35383 1337 35417
rect 1303 35063 1337 35097
rect 1303 34743 1337 34777
rect 1303 34423 1337 34457
rect 1463 36343 1497 36377
rect 1463 36023 1497 36057
rect 1463 35703 1497 35737
rect 1463 35383 1497 35417
rect 1463 35063 1497 35097
rect 1463 34743 1497 34777
rect 1463 34423 1497 34457
rect 1623 36343 1657 36377
rect 1623 36023 1657 36057
rect 1623 35703 1657 35737
rect 1623 35383 1657 35417
rect 1623 35063 1657 35097
rect 1623 34743 1657 34777
rect 1623 34423 1657 34457
rect 1783 36343 1817 36377
rect 1783 36023 1817 36057
rect 1783 35703 1817 35737
rect 1783 35383 1817 35417
rect 1783 35063 1817 35097
rect 1783 34743 1817 34777
rect 1783 34423 1817 34457
rect 1943 36343 1977 36377
rect 1943 36023 1977 36057
rect 1943 35703 1977 35737
rect 1943 35383 1977 35417
rect 1943 35063 1977 35097
rect 1943 34743 1977 34777
rect 1943 34423 1977 34457
rect 2103 36343 2137 36377
rect 2103 36023 2137 36057
rect 2103 35703 2137 35737
rect 2103 35383 2137 35417
rect 2103 35063 2137 35097
rect 2103 34743 2137 34777
rect 2103 34423 2137 34457
rect 2263 36343 2297 36377
rect 2263 36023 2297 36057
rect 2263 35703 2297 35737
rect 2263 35383 2297 35417
rect 2263 35063 2297 35097
rect 2263 34743 2297 34777
rect 2263 34423 2297 34457
rect 2423 36343 2457 36377
rect 2423 36023 2457 36057
rect 2423 35703 2457 35737
rect 2423 35383 2457 35417
rect 2423 35063 2457 35097
rect 2423 34743 2457 34777
rect 2423 34423 2457 34457
rect 2583 36343 2617 36377
rect 2583 36023 2617 36057
rect 2583 35703 2617 35737
rect 2583 35383 2617 35417
rect 2583 35063 2617 35097
rect 2583 34743 2617 34777
rect 2583 34423 2617 34457
rect 2743 36343 2777 36377
rect 2743 36023 2777 36057
rect 2743 35703 2777 35737
rect 2743 35383 2777 35417
rect 2743 35063 2777 35097
rect 2743 34743 2777 34777
rect 2743 34423 2777 34457
rect 2903 36343 2937 36377
rect 2903 36023 2937 36057
rect 2903 35703 2937 35737
rect 2903 35383 2937 35417
rect 2903 35063 2937 35097
rect 2903 34743 2937 34777
rect 2903 34423 2937 34457
rect 3063 36343 3097 36377
rect 3063 36023 3097 36057
rect 3063 35703 3097 35737
rect 3063 35383 3097 35417
rect 3063 35063 3097 35097
rect 3063 34743 3097 34777
rect 3063 34423 3097 34457
rect 3223 36343 3257 36377
rect 3223 36023 3257 36057
rect 3223 35703 3257 35737
rect 3223 35383 3257 35417
rect 3223 35063 3257 35097
rect 3223 34743 3257 34777
rect 3223 34423 3257 34457
rect 3383 36343 3417 36377
rect 3383 36023 3417 36057
rect 3383 35703 3417 35737
rect 3383 35383 3417 35417
rect 3383 35063 3417 35097
rect 3383 34743 3417 34777
rect 3383 34423 3417 34457
rect 3543 36343 3577 36377
rect 3543 36023 3577 36057
rect 3543 35703 3577 35737
rect 3543 35383 3577 35417
rect 3543 35063 3577 35097
rect 3543 34743 3577 34777
rect 3543 34423 3577 34457
rect 3703 36343 3737 36377
rect 3703 36023 3737 36057
rect 3703 35703 3737 35737
rect 3703 35383 3737 35417
rect 3703 35063 3737 35097
rect 3703 34743 3737 34777
rect 3703 34423 3737 34457
rect 3863 36343 3897 36377
rect 3863 36023 3897 36057
rect 3863 35703 3897 35737
rect 3863 35383 3897 35417
rect 3863 35063 3897 35097
rect 3863 34743 3897 34777
rect 3863 34423 3897 34457
rect 4023 36343 4057 36377
rect 4023 36023 4057 36057
rect 4023 35703 4057 35737
rect 4023 35383 4057 35417
rect 4023 35063 4057 35097
rect 4023 34743 4057 34777
rect 4023 34423 4057 34457
rect 4183 36343 4217 36377
rect 4183 36023 4217 36057
rect 4183 35703 4217 35737
rect 4183 35383 4217 35417
rect 4183 35063 4217 35097
rect 4183 34743 4217 34777
rect 4183 34423 4217 34457
rect 4343 36343 4377 36377
rect 4343 36023 4377 36057
rect 4343 35703 4377 35737
rect 4343 35383 4377 35417
rect 4343 35063 4377 35097
rect 4343 34743 4377 34777
rect 4343 34423 4377 34457
rect 4503 36343 4537 36377
rect 4503 36023 4537 36057
rect 4503 35703 4537 35737
rect 4503 35383 4537 35417
rect 4503 35063 4537 35097
rect 4503 34743 4537 34777
rect 4503 34423 4537 34457
rect 4663 36343 4697 36377
rect 4663 36023 4697 36057
rect 4663 35703 4697 35737
rect 4663 35383 4697 35417
rect 4663 35063 4697 35097
rect 4663 34743 4697 34777
rect 4663 34423 4697 34457
rect 4823 36343 4857 36377
rect 4823 36023 4857 36057
rect 4823 35703 4857 35737
rect 4823 35383 4857 35417
rect 4823 35063 4857 35097
rect 4823 34743 4857 34777
rect 4823 34423 4857 34457
rect 4983 36343 5017 36377
rect 4983 36023 5017 36057
rect 4983 35703 5017 35737
rect 4983 35383 5017 35417
rect 4983 35063 5017 35097
rect 4983 34743 5017 34777
rect 4983 34423 5017 34457
rect 5143 36343 5177 36377
rect 5143 36023 5177 36057
rect 5143 35703 5177 35737
rect 5143 35383 5177 35417
rect 5143 35063 5177 35097
rect 5143 34743 5177 34777
rect 5143 34423 5177 34457
rect 5303 36343 5337 36377
rect 5303 36023 5337 36057
rect 5303 35703 5337 35737
rect 5303 35383 5337 35417
rect 5303 35063 5337 35097
rect 5303 34743 5337 34777
rect 5303 34423 5337 34457
rect 5463 36343 5497 36377
rect 5463 36023 5497 36057
rect 5463 35703 5497 35737
rect 5463 35383 5497 35417
rect 5463 35063 5497 35097
rect 5463 34743 5497 34777
rect 5463 34423 5497 34457
rect 5623 36343 5657 36377
rect 5623 36023 5657 36057
rect 5623 35703 5657 35737
rect 5623 35383 5657 35417
rect 5623 35063 5657 35097
rect 5623 34743 5657 34777
rect 5623 34423 5657 34457
rect 5783 36343 5817 36377
rect 5783 36023 5817 36057
rect 5783 35703 5817 35737
rect 5783 35383 5817 35417
rect 5783 35063 5817 35097
rect 5783 34743 5817 34777
rect 5783 34423 5817 34457
rect 5943 36343 5977 36377
rect 5943 36023 5977 36057
rect 5943 35703 5977 35737
rect 5943 35383 5977 35417
rect 5943 35063 5977 35097
rect 5943 34743 5977 34777
rect 5943 34423 5977 34457
rect 6103 36343 6137 36377
rect 6103 36023 6137 36057
rect 6103 35703 6137 35737
rect 6103 35383 6137 35417
rect 6103 35063 6137 35097
rect 6103 34743 6137 34777
rect 6103 34423 6137 34457
rect 6263 36343 6297 36377
rect 6263 36023 6297 36057
rect 6263 35703 6297 35737
rect 6263 35383 6297 35417
rect 6263 35063 6297 35097
rect 6263 34743 6297 34777
rect 6263 34423 6297 34457
rect 6423 36343 6457 36377
rect 6423 36023 6457 36057
rect 6423 35703 6457 35737
rect 6423 35383 6457 35417
rect 6423 35063 6457 35097
rect 6423 34743 6457 34777
rect 6423 34423 6457 34457
rect 6583 36343 6617 36377
rect 6583 36023 6617 36057
rect 6583 35703 6617 35737
rect 6583 35383 6617 35417
rect 6583 35063 6617 35097
rect 6583 34743 6617 34777
rect 6583 34423 6617 34457
rect 6743 36343 6777 36377
rect 6743 36023 6777 36057
rect 6743 35703 6777 35737
rect 6743 35383 6777 35417
rect 6743 35063 6777 35097
rect 6743 34743 6777 34777
rect 6743 34423 6777 34457
rect 6903 36343 6937 36377
rect 6903 36023 6937 36057
rect 6903 35703 6937 35737
rect 6903 35383 6937 35417
rect 6903 35063 6937 35097
rect 6903 34743 6937 34777
rect 6903 34423 6937 34457
rect 7063 36343 7097 36377
rect 7063 36023 7097 36057
rect 7063 35703 7097 35737
rect 7063 35383 7097 35417
rect 7063 35063 7097 35097
rect 7063 34743 7097 34777
rect 7063 34423 7097 34457
rect 7223 36343 7257 36377
rect 7223 36023 7257 36057
rect 7223 35703 7257 35737
rect 7223 35383 7257 35417
rect 7223 35063 7257 35097
rect 7223 34743 7257 34777
rect 7223 34423 7257 34457
rect 7383 36343 7417 36377
rect 7383 36023 7417 36057
rect 7383 35703 7417 35737
rect 7383 35383 7417 35417
rect 7383 35063 7417 35097
rect 7383 34743 7417 34777
rect 7383 34423 7417 34457
rect 7543 36343 7577 36377
rect 7543 36023 7577 36057
rect 7543 35703 7577 35737
rect 7543 35383 7577 35417
rect 7543 35063 7577 35097
rect 7543 34743 7577 34777
rect 7543 34423 7577 34457
rect 7703 36343 7737 36377
rect 7703 36023 7737 36057
rect 7703 35703 7737 35737
rect 7703 35383 7737 35417
rect 7703 35063 7737 35097
rect 7703 34743 7737 34777
rect 7703 34423 7737 34457
rect 7863 36343 7897 36377
rect 7863 36023 7897 36057
rect 7863 35703 7897 35737
rect 7863 35383 7897 35417
rect 7863 35063 7897 35097
rect 7863 34743 7897 34777
rect 7863 34423 7897 34457
rect 8023 36343 8057 36377
rect 8023 36023 8057 36057
rect 8023 35703 8057 35737
rect 8023 35383 8057 35417
rect 8023 35063 8057 35097
rect 8023 34743 8057 34777
rect 8023 34423 8057 34457
rect 8183 36343 8217 36377
rect 8183 36023 8217 36057
rect 8183 35703 8217 35737
rect 8183 35383 8217 35417
rect 8183 35063 8217 35097
rect 8183 34743 8217 34777
rect 8183 34423 8217 34457
rect 8343 36343 8377 36377
rect 8343 36023 8377 36057
rect 8343 35703 8377 35737
rect 8343 35383 8377 35417
rect 8343 35063 8377 35097
rect 8343 34743 8377 34777
rect 8343 34423 8377 34457
rect 12503 36343 12537 36377
rect 12503 36023 12537 36057
rect 12503 35703 12537 35737
rect 12503 35383 12537 35417
rect 12503 35063 12537 35097
rect 12503 34743 12537 34777
rect 12503 34423 12537 34457
rect 12663 36343 12697 36377
rect 12663 36023 12697 36057
rect 12663 35703 12697 35737
rect 12663 35383 12697 35417
rect 12663 35063 12697 35097
rect 12663 34743 12697 34777
rect 12663 34423 12697 34457
rect 12823 36343 12857 36377
rect 12823 36023 12857 36057
rect 12823 35703 12857 35737
rect 12823 35383 12857 35417
rect 12823 35063 12857 35097
rect 12823 34743 12857 34777
rect 12823 34423 12857 34457
rect 12983 36343 13017 36377
rect 12983 36023 13017 36057
rect 12983 35703 13017 35737
rect 12983 35383 13017 35417
rect 12983 35063 13017 35097
rect 12983 34743 13017 34777
rect 12983 34423 13017 34457
rect 13143 36343 13177 36377
rect 13143 36023 13177 36057
rect 13143 35703 13177 35737
rect 13143 35383 13177 35417
rect 13143 35063 13177 35097
rect 13143 34743 13177 34777
rect 13143 34423 13177 34457
rect 13303 36343 13337 36377
rect 13303 36023 13337 36057
rect 13303 35703 13337 35737
rect 13303 35383 13337 35417
rect 13303 35063 13337 35097
rect 13303 34743 13337 34777
rect 13303 34423 13337 34457
rect 13463 36343 13497 36377
rect 13463 36023 13497 36057
rect 13463 35703 13497 35737
rect 13463 35383 13497 35417
rect 13463 35063 13497 35097
rect 13463 34743 13497 34777
rect 13463 34423 13497 34457
rect 13623 36343 13657 36377
rect 13623 36023 13657 36057
rect 13623 35703 13657 35737
rect 13623 35383 13657 35417
rect 13623 35063 13657 35097
rect 13623 34743 13657 34777
rect 13623 34423 13657 34457
rect 13783 36343 13817 36377
rect 13783 36023 13817 36057
rect 13783 35703 13817 35737
rect 13783 35383 13817 35417
rect 13783 35063 13817 35097
rect 13783 34743 13817 34777
rect 13783 34423 13817 34457
rect 13943 36343 13977 36377
rect 13943 36023 13977 36057
rect 13943 35703 13977 35737
rect 13943 35383 13977 35417
rect 13943 35063 13977 35097
rect 13943 34743 13977 34777
rect 13943 34423 13977 34457
rect 14103 36343 14137 36377
rect 14103 36023 14137 36057
rect 14103 35703 14137 35737
rect 14103 35383 14137 35417
rect 14103 35063 14137 35097
rect 14103 34743 14137 34777
rect 14103 34423 14137 34457
rect 14263 36343 14297 36377
rect 14263 36023 14297 36057
rect 14263 35703 14297 35737
rect 14263 35383 14297 35417
rect 14263 35063 14297 35097
rect 14263 34743 14297 34777
rect 14263 34423 14297 34457
rect 14423 36343 14457 36377
rect 14423 36023 14457 36057
rect 14423 35703 14457 35737
rect 14423 35383 14457 35417
rect 14423 35063 14457 35097
rect 14423 34743 14457 34777
rect 14423 34423 14457 34457
rect 14583 36343 14617 36377
rect 14583 36023 14617 36057
rect 14583 35703 14617 35737
rect 14583 35383 14617 35417
rect 14583 35063 14617 35097
rect 14583 34743 14617 34777
rect 14583 34423 14617 34457
rect 14743 36343 14777 36377
rect 14743 36023 14777 36057
rect 14743 35703 14777 35737
rect 14743 35383 14777 35417
rect 14743 35063 14777 35097
rect 14743 34743 14777 34777
rect 14743 34423 14777 34457
rect 14903 36343 14937 36377
rect 14903 36023 14937 36057
rect 14903 35703 14937 35737
rect 14903 35383 14937 35417
rect 14903 35063 14937 35097
rect 14903 34743 14937 34777
rect 14903 34423 14937 34457
rect 15063 36343 15097 36377
rect 15063 36023 15097 36057
rect 15063 35703 15097 35737
rect 15063 35383 15097 35417
rect 15063 35063 15097 35097
rect 15063 34743 15097 34777
rect 15063 34423 15097 34457
rect 15223 36343 15257 36377
rect 15223 36023 15257 36057
rect 15223 35703 15257 35737
rect 15223 35383 15257 35417
rect 15223 35063 15257 35097
rect 15223 34743 15257 34777
rect 15223 34423 15257 34457
rect 15383 36343 15417 36377
rect 15383 36023 15417 36057
rect 15383 35703 15417 35737
rect 15383 35383 15417 35417
rect 15383 35063 15417 35097
rect 15383 34743 15417 34777
rect 15383 34423 15417 34457
rect 15543 36343 15577 36377
rect 15543 36023 15577 36057
rect 15543 35703 15577 35737
rect 15543 35383 15577 35417
rect 15543 35063 15577 35097
rect 15543 34743 15577 34777
rect 15543 34423 15577 34457
rect 15703 36343 15737 36377
rect 15703 36023 15737 36057
rect 15703 35703 15737 35737
rect 15703 35383 15737 35417
rect 15703 35063 15737 35097
rect 15703 34743 15737 34777
rect 15703 34423 15737 34457
rect 15863 36343 15897 36377
rect 15863 36023 15897 36057
rect 15863 35703 15897 35737
rect 15863 35383 15897 35417
rect 15863 35063 15897 35097
rect 15863 34743 15897 34777
rect 15863 34423 15897 34457
rect 16023 36343 16057 36377
rect 16023 36023 16057 36057
rect 16023 35703 16057 35737
rect 16023 35383 16057 35417
rect 16023 35063 16057 35097
rect 16023 34743 16057 34777
rect 16023 34423 16057 34457
rect 16183 36343 16217 36377
rect 16183 36023 16217 36057
rect 16183 35703 16217 35737
rect 16183 35383 16217 35417
rect 16183 35063 16217 35097
rect 16183 34743 16217 34777
rect 16183 34423 16217 34457
rect 16343 36343 16377 36377
rect 16343 36023 16377 36057
rect 16343 35703 16377 35737
rect 16343 35383 16377 35417
rect 16343 35063 16377 35097
rect 16343 34743 16377 34777
rect 16343 34423 16377 34457
rect 16503 36343 16537 36377
rect 16503 36023 16537 36057
rect 16503 35703 16537 35737
rect 16503 35383 16537 35417
rect 16503 35063 16537 35097
rect 16503 34743 16537 34777
rect 16503 34423 16537 34457
rect 16663 36343 16697 36377
rect 16663 36023 16697 36057
rect 16663 35703 16697 35737
rect 16663 35383 16697 35417
rect 16663 35063 16697 35097
rect 16663 34743 16697 34777
rect 16663 34423 16697 34457
rect 16823 36343 16857 36377
rect 16823 36023 16857 36057
rect 16823 35703 16857 35737
rect 16823 35383 16857 35417
rect 16823 35063 16857 35097
rect 16823 34743 16857 34777
rect 16823 34423 16857 34457
rect 16983 36343 17017 36377
rect 16983 36023 17017 36057
rect 16983 35703 17017 35737
rect 16983 35383 17017 35417
rect 16983 35063 17017 35097
rect 16983 34743 17017 34777
rect 16983 34423 17017 34457
rect 17143 36343 17177 36377
rect 17143 36023 17177 36057
rect 17143 35703 17177 35737
rect 17143 35383 17177 35417
rect 17143 35063 17177 35097
rect 17143 34743 17177 34777
rect 17143 34423 17177 34457
rect 17303 36343 17337 36377
rect 17303 36023 17337 36057
rect 17303 35703 17337 35737
rect 17303 35383 17337 35417
rect 17303 35063 17337 35097
rect 17303 34743 17337 34777
rect 17303 34423 17337 34457
rect 17463 36343 17497 36377
rect 17463 36023 17497 36057
rect 17463 35703 17497 35737
rect 17463 35383 17497 35417
rect 17463 35063 17497 35097
rect 17463 34743 17497 34777
rect 17463 34423 17497 34457
rect 17623 36343 17657 36377
rect 17623 36023 17657 36057
rect 17623 35703 17657 35737
rect 17623 35383 17657 35417
rect 17623 35063 17657 35097
rect 17623 34743 17657 34777
rect 17623 34423 17657 34457
rect 17783 36343 17817 36377
rect 17783 36023 17817 36057
rect 17783 35703 17817 35737
rect 17783 35383 17817 35417
rect 17783 35063 17817 35097
rect 17783 34743 17817 34777
rect 17783 34423 17817 34457
rect 17943 36343 17977 36377
rect 17943 36023 17977 36057
rect 17943 35703 17977 35737
rect 17943 35383 17977 35417
rect 17943 35063 17977 35097
rect 17943 34743 17977 34777
rect 17943 34423 17977 34457
rect 18103 36343 18137 36377
rect 18103 36023 18137 36057
rect 18103 35703 18137 35737
rect 18103 35383 18137 35417
rect 18103 35063 18137 35097
rect 18103 34743 18137 34777
rect 18103 34423 18137 34457
rect 18263 36343 18297 36377
rect 18263 36023 18297 36057
rect 18263 35703 18297 35737
rect 18263 35383 18297 35417
rect 18263 35063 18297 35097
rect 18263 34743 18297 34777
rect 18263 34423 18297 34457
rect 18423 36343 18457 36377
rect 18423 36023 18457 36057
rect 18423 35703 18457 35737
rect 18423 35383 18457 35417
rect 18423 35063 18457 35097
rect 18423 34743 18457 34777
rect 18423 34423 18457 34457
rect 18583 36343 18617 36377
rect 18583 36023 18617 36057
rect 18583 35703 18617 35737
rect 18583 35383 18617 35417
rect 18583 35063 18617 35097
rect 18583 34743 18617 34777
rect 18583 34423 18617 34457
rect 18743 36343 18777 36377
rect 18743 36023 18777 36057
rect 18743 35703 18777 35737
rect 18743 35383 18777 35417
rect 18743 35063 18777 35097
rect 18743 34743 18777 34777
rect 18743 34423 18777 34457
rect 18903 36343 18937 36377
rect 18903 36023 18937 36057
rect 18903 35703 18937 35737
rect 18903 35383 18937 35417
rect 18903 35063 18937 35097
rect 18903 34743 18937 34777
rect 18903 34423 18937 34457
rect 23143 36343 23177 36377
rect 23143 36023 23177 36057
rect 23143 35703 23177 35737
rect 23143 35383 23177 35417
rect 23143 35063 23177 35097
rect 23143 34743 23177 34777
rect 23143 34423 23177 34457
rect 23303 36343 23337 36377
rect 23303 36023 23337 36057
rect 23303 35703 23337 35737
rect 23303 35383 23337 35417
rect 23303 35063 23337 35097
rect 23303 34743 23337 34777
rect 23303 34423 23337 34457
rect 23463 36343 23497 36377
rect 23463 36023 23497 36057
rect 23463 35703 23497 35737
rect 23463 35383 23497 35417
rect 23463 35063 23497 35097
rect 23463 34743 23497 34777
rect 23463 34423 23497 34457
rect 23623 36343 23657 36377
rect 23623 36023 23657 36057
rect 23623 35703 23657 35737
rect 23623 35383 23657 35417
rect 23623 35063 23657 35097
rect 23623 34743 23657 34777
rect 23623 34423 23657 34457
rect 23783 36343 23817 36377
rect 23783 36023 23817 36057
rect 23783 35703 23817 35737
rect 23783 35383 23817 35417
rect 23783 35063 23817 35097
rect 23783 34743 23817 34777
rect 23783 34423 23817 34457
rect 23943 36343 23977 36377
rect 23943 36023 23977 36057
rect 23943 35703 23977 35737
rect 23943 35383 23977 35417
rect 23943 35063 23977 35097
rect 23943 34743 23977 34777
rect 23943 34423 23977 34457
rect 24103 36343 24137 36377
rect 24103 36023 24137 36057
rect 24103 35703 24137 35737
rect 24103 35383 24137 35417
rect 24103 35063 24137 35097
rect 24103 34743 24137 34777
rect 24103 34423 24137 34457
rect 24263 36343 24297 36377
rect 24263 36023 24297 36057
rect 24263 35703 24297 35737
rect 24263 35383 24297 35417
rect 24263 35063 24297 35097
rect 24263 34743 24297 34777
rect 24263 34423 24297 34457
rect 24423 36343 24457 36377
rect 24423 36023 24457 36057
rect 24423 35703 24457 35737
rect 24423 35383 24457 35417
rect 24423 35063 24457 35097
rect 24423 34743 24457 34777
rect 24423 34423 24457 34457
rect 24583 36343 24617 36377
rect 24583 36023 24617 36057
rect 24583 35703 24617 35737
rect 24583 35383 24617 35417
rect 24583 35063 24617 35097
rect 24583 34743 24617 34777
rect 24583 34423 24617 34457
rect 24743 36343 24777 36377
rect 24743 36023 24777 36057
rect 24743 35703 24777 35737
rect 24743 35383 24777 35417
rect 24743 35063 24777 35097
rect 24743 34743 24777 34777
rect 24743 34423 24777 34457
rect 24903 36343 24937 36377
rect 24903 36023 24937 36057
rect 24903 35703 24937 35737
rect 24903 35383 24937 35417
rect 24903 35063 24937 35097
rect 24903 34743 24937 34777
rect 24903 34423 24937 34457
rect 25063 36343 25097 36377
rect 25063 36023 25097 36057
rect 25063 35703 25097 35737
rect 25063 35383 25097 35417
rect 25063 35063 25097 35097
rect 25063 34743 25097 34777
rect 25063 34423 25097 34457
rect 25223 36343 25257 36377
rect 25223 36023 25257 36057
rect 25223 35703 25257 35737
rect 25223 35383 25257 35417
rect 25223 35063 25257 35097
rect 25223 34743 25257 34777
rect 25223 34423 25257 34457
rect 25383 36343 25417 36377
rect 25383 36023 25417 36057
rect 25383 35703 25417 35737
rect 25383 35383 25417 35417
rect 25383 35063 25417 35097
rect 25383 34743 25417 34777
rect 25383 34423 25417 34457
rect 25543 36343 25577 36377
rect 25543 36023 25577 36057
rect 25543 35703 25577 35737
rect 25543 35383 25577 35417
rect 25543 35063 25577 35097
rect 25543 34743 25577 34777
rect 25543 34423 25577 34457
rect 25703 36343 25737 36377
rect 25703 36023 25737 36057
rect 25703 35703 25737 35737
rect 25703 35383 25737 35417
rect 25703 35063 25737 35097
rect 25703 34743 25737 34777
rect 25703 34423 25737 34457
rect 25863 36343 25897 36377
rect 25863 36023 25897 36057
rect 25863 35703 25897 35737
rect 25863 35383 25897 35417
rect 25863 35063 25897 35097
rect 25863 34743 25897 34777
rect 25863 34423 25897 34457
rect 26023 36343 26057 36377
rect 26023 36023 26057 36057
rect 26023 35703 26057 35737
rect 26023 35383 26057 35417
rect 26023 35063 26057 35097
rect 26023 34743 26057 34777
rect 26023 34423 26057 34457
rect 26183 36343 26217 36377
rect 26183 36023 26217 36057
rect 26183 35703 26217 35737
rect 26183 35383 26217 35417
rect 26183 35063 26217 35097
rect 26183 34743 26217 34777
rect 26183 34423 26217 34457
rect 26343 36343 26377 36377
rect 26343 36023 26377 36057
rect 26343 35703 26377 35737
rect 26343 35383 26377 35417
rect 26343 35063 26377 35097
rect 26343 34743 26377 34777
rect 26343 34423 26377 34457
rect 26503 36343 26537 36377
rect 26503 36023 26537 36057
rect 26503 35703 26537 35737
rect 26503 35383 26537 35417
rect 26503 35063 26537 35097
rect 26503 34743 26537 34777
rect 26503 34423 26537 34457
rect 26663 36343 26697 36377
rect 26663 36023 26697 36057
rect 26663 35703 26697 35737
rect 26663 35383 26697 35417
rect 26663 35063 26697 35097
rect 26663 34743 26697 34777
rect 26663 34423 26697 34457
rect 26823 36343 26857 36377
rect 26823 36023 26857 36057
rect 26823 35703 26857 35737
rect 26823 35383 26857 35417
rect 26823 35063 26857 35097
rect 26823 34743 26857 34777
rect 26823 34423 26857 34457
rect 26983 36343 27017 36377
rect 26983 36023 27017 36057
rect 26983 35703 27017 35737
rect 26983 35383 27017 35417
rect 26983 35063 27017 35097
rect 26983 34743 27017 34777
rect 26983 34423 27017 34457
rect 27143 36343 27177 36377
rect 27143 36023 27177 36057
rect 27143 35703 27177 35737
rect 27143 35383 27177 35417
rect 27143 35063 27177 35097
rect 27143 34743 27177 34777
rect 27143 34423 27177 34457
rect 27303 36343 27337 36377
rect 27303 36023 27337 36057
rect 27303 35703 27337 35737
rect 27303 35383 27337 35417
rect 27303 35063 27337 35097
rect 27303 34743 27337 34777
rect 27303 34423 27337 34457
rect 27463 36343 27497 36377
rect 27463 36023 27497 36057
rect 27463 35703 27497 35737
rect 27463 35383 27497 35417
rect 27463 35063 27497 35097
rect 27463 34743 27497 34777
rect 27463 34423 27497 34457
rect 27623 36343 27657 36377
rect 27623 36023 27657 36057
rect 27623 35703 27657 35737
rect 27623 35383 27657 35417
rect 27623 35063 27657 35097
rect 27623 34743 27657 34777
rect 27623 34423 27657 34457
rect 27783 36343 27817 36377
rect 27783 36023 27817 36057
rect 27783 35703 27817 35737
rect 27783 35383 27817 35417
rect 27783 35063 27817 35097
rect 27783 34743 27817 34777
rect 27783 34423 27817 34457
rect 27943 36343 27977 36377
rect 27943 36023 27977 36057
rect 27943 35703 27977 35737
rect 27943 35383 27977 35417
rect 27943 35063 27977 35097
rect 27943 34743 27977 34777
rect 27943 34423 27977 34457
rect 28103 36343 28137 36377
rect 28103 36023 28137 36057
rect 28103 35703 28137 35737
rect 28103 35383 28137 35417
rect 28103 35063 28137 35097
rect 28103 34743 28137 34777
rect 28103 34423 28137 34457
rect 28263 36343 28297 36377
rect 28263 36023 28297 36057
rect 28263 35703 28297 35737
rect 28263 35383 28297 35417
rect 28263 35063 28297 35097
rect 28263 34743 28297 34777
rect 28263 34423 28297 34457
rect 28423 36343 28457 36377
rect 28423 36023 28457 36057
rect 28423 35703 28457 35737
rect 28423 35383 28457 35417
rect 28423 35063 28457 35097
rect 28423 34743 28457 34777
rect 28423 34423 28457 34457
rect 28583 36343 28617 36377
rect 28583 36023 28617 36057
rect 28583 35703 28617 35737
rect 28583 35383 28617 35417
rect 28583 35063 28617 35097
rect 28583 34743 28617 34777
rect 28583 34423 28617 34457
rect 28743 36343 28777 36377
rect 28743 36023 28777 36057
rect 28743 35703 28777 35737
rect 28743 35383 28777 35417
rect 28743 35063 28777 35097
rect 28743 34743 28777 34777
rect 28743 34423 28777 34457
rect 28903 36343 28937 36377
rect 28903 36023 28937 36057
rect 28903 35703 28937 35737
rect 28903 35383 28937 35417
rect 28903 35063 28937 35097
rect 28903 34743 28937 34777
rect 28903 34423 28937 34457
rect 29063 36343 29097 36377
rect 29063 36023 29097 36057
rect 29063 35703 29097 35737
rect 29063 35383 29097 35417
rect 29063 35063 29097 35097
rect 29063 34743 29097 34777
rect 29063 34423 29097 34457
rect 29223 36343 29257 36377
rect 29223 36023 29257 36057
rect 29223 35703 29257 35737
rect 29223 35383 29257 35417
rect 29223 35063 29257 35097
rect 29223 34743 29257 34777
rect 29223 34423 29257 34457
rect 29383 36343 29417 36377
rect 29383 36023 29417 36057
rect 29383 35703 29417 35737
rect 29383 35383 29417 35417
rect 29383 35063 29417 35097
rect 29383 34743 29417 34777
rect 29383 34423 29417 34457
rect 33543 36343 33577 36377
rect 33543 36023 33577 36057
rect 33543 35703 33577 35737
rect 33543 35383 33577 35417
rect 33543 35063 33577 35097
rect 33543 34743 33577 34777
rect 33543 34423 33577 34457
rect 33703 36343 33737 36377
rect 33703 36023 33737 36057
rect 33703 35703 33737 35737
rect 33703 35383 33737 35417
rect 33703 35063 33737 35097
rect 33703 34743 33737 34777
rect 33703 34423 33737 34457
rect 33863 36343 33897 36377
rect 33863 36023 33897 36057
rect 33863 35703 33897 35737
rect 33863 35383 33897 35417
rect 33863 35063 33897 35097
rect 33863 34743 33897 34777
rect 33863 34423 33897 34457
rect 34023 36343 34057 36377
rect 34023 36023 34057 36057
rect 34023 35703 34057 35737
rect 34023 35383 34057 35417
rect 34023 35063 34057 35097
rect 34023 34743 34057 34777
rect 34023 34423 34057 34457
rect 34183 36343 34217 36377
rect 34183 36023 34217 36057
rect 34183 35703 34217 35737
rect 34183 35383 34217 35417
rect 34183 35063 34217 35097
rect 34183 34743 34217 34777
rect 34183 34423 34217 34457
rect 34343 36343 34377 36377
rect 34343 36023 34377 36057
rect 34343 35703 34377 35737
rect 34343 35383 34377 35417
rect 34343 35063 34377 35097
rect 34343 34743 34377 34777
rect 34343 34423 34377 34457
rect 34503 36343 34537 36377
rect 34503 36023 34537 36057
rect 34503 35703 34537 35737
rect 34503 35383 34537 35417
rect 34503 35063 34537 35097
rect 34503 34743 34537 34777
rect 34503 34423 34537 34457
rect 34663 36343 34697 36377
rect 34663 36023 34697 36057
rect 34663 35703 34697 35737
rect 34663 35383 34697 35417
rect 34663 35063 34697 35097
rect 34663 34743 34697 34777
rect 34663 34423 34697 34457
rect 34823 36343 34857 36377
rect 34823 36023 34857 36057
rect 34823 35703 34857 35737
rect 34823 35383 34857 35417
rect 34823 35063 34857 35097
rect 34823 34743 34857 34777
rect 34823 34423 34857 34457
rect 34983 36343 35017 36377
rect 34983 36023 35017 36057
rect 34983 35703 35017 35737
rect 34983 35383 35017 35417
rect 34983 35063 35017 35097
rect 34983 34743 35017 34777
rect 34983 34423 35017 34457
rect 35143 36343 35177 36377
rect 35143 36023 35177 36057
rect 35143 35703 35177 35737
rect 35143 35383 35177 35417
rect 35143 35063 35177 35097
rect 35143 34743 35177 34777
rect 35143 34423 35177 34457
rect 35303 36343 35337 36377
rect 35303 36023 35337 36057
rect 35303 35703 35337 35737
rect 35303 35383 35337 35417
rect 35303 35063 35337 35097
rect 35303 34743 35337 34777
rect 35303 34423 35337 34457
rect 35463 36343 35497 36377
rect 35463 36023 35497 36057
rect 35463 35703 35497 35737
rect 35463 35383 35497 35417
rect 35463 35063 35497 35097
rect 35463 34743 35497 34777
rect 35463 34423 35497 34457
rect 35623 36343 35657 36377
rect 35623 36023 35657 36057
rect 35623 35703 35657 35737
rect 35623 35383 35657 35417
rect 35623 35063 35657 35097
rect 35623 34743 35657 34777
rect 35623 34423 35657 34457
rect 35783 36343 35817 36377
rect 35783 36023 35817 36057
rect 35783 35703 35817 35737
rect 35783 35383 35817 35417
rect 35783 35063 35817 35097
rect 35783 34743 35817 34777
rect 35783 34423 35817 34457
rect 35943 36343 35977 36377
rect 35943 36023 35977 36057
rect 35943 35703 35977 35737
rect 35943 35383 35977 35417
rect 35943 35063 35977 35097
rect 35943 34743 35977 34777
rect 35943 34423 35977 34457
rect 36103 36343 36137 36377
rect 36103 36023 36137 36057
rect 36103 35703 36137 35737
rect 36103 35383 36137 35417
rect 36103 35063 36137 35097
rect 36103 34743 36137 34777
rect 36103 34423 36137 34457
rect 36263 36343 36297 36377
rect 36263 36023 36297 36057
rect 36263 35703 36297 35737
rect 36263 35383 36297 35417
rect 36263 35063 36297 35097
rect 36263 34743 36297 34777
rect 36263 34423 36297 34457
rect 36423 36343 36457 36377
rect 36423 36023 36457 36057
rect 36423 35703 36457 35737
rect 36423 35383 36457 35417
rect 36423 35063 36457 35097
rect 36423 34743 36457 34777
rect 36423 34423 36457 34457
rect 36583 36343 36617 36377
rect 36583 36023 36617 36057
rect 36583 35703 36617 35737
rect 36583 35383 36617 35417
rect 36583 35063 36617 35097
rect 36583 34743 36617 34777
rect 36583 34423 36617 34457
rect 36743 36343 36777 36377
rect 36743 36023 36777 36057
rect 36743 35703 36777 35737
rect 36743 35383 36777 35417
rect 36743 35063 36777 35097
rect 36743 34743 36777 34777
rect 36743 34423 36777 34457
rect 36903 36343 36937 36377
rect 36903 36023 36937 36057
rect 36903 35703 36937 35737
rect 36903 35383 36937 35417
rect 36903 35063 36937 35097
rect 36903 34743 36937 34777
rect 36903 34423 36937 34457
rect 37063 36343 37097 36377
rect 37063 36023 37097 36057
rect 37063 35703 37097 35737
rect 37063 35383 37097 35417
rect 37063 35063 37097 35097
rect 37063 34743 37097 34777
rect 37063 34423 37097 34457
rect 37223 36343 37257 36377
rect 37223 36023 37257 36057
rect 37223 35703 37257 35737
rect 37223 35383 37257 35417
rect 37223 35063 37257 35097
rect 37223 34743 37257 34777
rect 37223 34423 37257 34457
rect 37383 36343 37417 36377
rect 37383 36023 37417 36057
rect 37383 35703 37417 35737
rect 37383 35383 37417 35417
rect 37383 35063 37417 35097
rect 37383 34743 37417 34777
rect 37383 34423 37417 34457
rect 37543 36343 37577 36377
rect 37543 36023 37577 36057
rect 37543 35703 37577 35737
rect 37543 35383 37577 35417
rect 37543 35063 37577 35097
rect 37543 34743 37577 34777
rect 37543 34423 37577 34457
rect 37703 36343 37737 36377
rect 37703 36023 37737 36057
rect 37703 35703 37737 35737
rect 37703 35383 37737 35417
rect 37703 35063 37737 35097
rect 37703 34743 37737 34777
rect 37703 34423 37737 34457
rect 37863 36343 37897 36377
rect 37863 36023 37897 36057
rect 37863 35703 37897 35737
rect 37863 35383 37897 35417
rect 37863 35063 37897 35097
rect 37863 34743 37897 34777
rect 37863 34423 37897 34457
rect 38023 36343 38057 36377
rect 38023 36023 38057 36057
rect 38023 35703 38057 35737
rect 38023 35383 38057 35417
rect 38023 35063 38057 35097
rect 38023 34743 38057 34777
rect 38023 34423 38057 34457
rect 38183 36343 38217 36377
rect 38183 36023 38217 36057
rect 38183 35703 38217 35737
rect 38183 35383 38217 35417
rect 38183 35063 38217 35097
rect 38183 34743 38217 34777
rect 38183 34423 38217 34457
rect 38343 36343 38377 36377
rect 38343 36023 38377 36057
rect 38343 35703 38377 35737
rect 38343 35383 38377 35417
rect 38343 35063 38377 35097
rect 38343 34743 38377 34777
rect 38343 34423 38377 34457
rect 38503 36343 38537 36377
rect 38503 36023 38537 36057
rect 38503 35703 38537 35737
rect 38503 35383 38537 35417
rect 38503 35063 38537 35097
rect 38503 34743 38537 34777
rect 38503 34423 38537 34457
rect 38663 36343 38697 36377
rect 38663 36023 38697 36057
rect 38663 35703 38697 35737
rect 38663 35383 38697 35417
rect 38663 35063 38697 35097
rect 38663 34743 38697 34777
rect 38663 34423 38697 34457
rect 38823 36343 38857 36377
rect 38823 36023 38857 36057
rect 38823 35703 38857 35737
rect 38823 35383 38857 35417
rect 38823 35063 38857 35097
rect 38823 34743 38857 34777
rect 38823 34423 38857 34457
rect 38983 36343 39017 36377
rect 38983 36023 39017 36057
rect 38983 35703 39017 35737
rect 38983 35383 39017 35417
rect 38983 35063 39017 35097
rect 38983 34743 39017 34777
rect 38983 34423 39017 34457
rect 39143 36343 39177 36377
rect 39143 36023 39177 36057
rect 39143 35703 39177 35737
rect 39143 35383 39177 35417
rect 39143 35063 39177 35097
rect 39143 34743 39177 34777
rect 39143 34423 39177 34457
rect 39303 36343 39337 36377
rect 39303 36023 39337 36057
rect 39303 35703 39337 35737
rect 39303 35383 39337 35417
rect 39303 35063 39337 35097
rect 39303 34743 39337 34777
rect 39303 34423 39337 34457
rect 39463 36343 39497 36377
rect 39463 36023 39497 36057
rect 39463 35703 39497 35737
rect 39463 35383 39497 35417
rect 39463 35063 39497 35097
rect 39463 34743 39497 34777
rect 39463 34423 39497 34457
rect 39623 36343 39657 36377
rect 39623 36023 39657 36057
rect 39623 35703 39657 35737
rect 39623 35383 39657 35417
rect 39623 35063 39657 35097
rect 39623 34743 39657 34777
rect 39623 34423 39657 34457
rect 39783 36343 39817 36377
rect 39783 36023 39817 36057
rect 39783 35703 39817 35737
rect 39783 35383 39817 35417
rect 39783 35063 39817 35097
rect 39783 34743 39817 34777
rect 39783 34423 39817 34457
rect 39943 36343 39977 36377
rect 39943 36023 39977 36057
rect 39943 35703 39977 35737
rect 39943 35383 39977 35417
rect 39943 35063 39977 35097
rect 39943 34743 39977 34777
rect 39943 34423 39977 34457
rect 40103 36343 40137 36377
rect 40103 36023 40137 36057
rect 40103 35703 40137 35737
rect 40103 35383 40137 35417
rect 40103 35063 40137 35097
rect 40103 34743 40137 34777
rect 40103 34423 40137 34457
rect 40263 36343 40297 36377
rect 40263 36023 40297 36057
rect 40263 35703 40297 35737
rect 40263 35383 40297 35417
rect 40263 35063 40297 35097
rect 40263 34743 40297 34777
rect 40263 34423 40297 34457
rect 40423 36343 40457 36377
rect 40423 36023 40457 36057
rect 40423 35703 40457 35737
rect 40423 35383 40457 35417
rect 40423 35063 40457 35097
rect 40423 34743 40457 34777
rect 40423 34423 40457 34457
rect 40583 36343 40617 36377
rect 40583 36023 40617 36057
rect 40583 35703 40617 35737
rect 40583 35383 40617 35417
rect 40583 35063 40617 35097
rect 40583 34743 40617 34777
rect 40583 34423 40617 34457
rect 40743 36343 40777 36377
rect 40743 36023 40777 36057
rect 40743 35703 40777 35737
rect 40743 35383 40777 35417
rect 40743 35063 40777 35097
rect 40743 34743 40777 34777
rect 40743 34423 40777 34457
rect 40903 36343 40937 36377
rect 40903 36023 40937 36057
rect 40903 35703 40937 35737
rect 40903 35383 40937 35417
rect 40903 35063 40937 35097
rect 40903 34743 40937 34777
rect 40903 34423 40937 34457
rect 41063 36343 41097 36377
rect 41063 36023 41097 36057
rect 41063 35703 41097 35737
rect 41063 35383 41097 35417
rect 41063 35063 41097 35097
rect 41063 34743 41097 34777
rect 41063 34423 41097 34457
rect 41223 36343 41257 36377
rect 41223 36023 41257 36057
rect 41223 35703 41257 35737
rect 41223 35383 41257 35417
rect 41223 35063 41257 35097
rect 41223 34743 41257 34777
rect 41223 34423 41257 34457
rect 41383 36343 41417 36377
rect 41383 36023 41417 36057
rect 41383 35703 41417 35737
rect 41383 35383 41417 35417
rect 41383 35063 41417 35097
rect 41383 34743 41417 34777
rect 41383 34423 41417 34457
rect 41543 36343 41577 36377
rect 41543 36023 41577 36057
rect 41543 35703 41577 35737
rect 41543 35383 41577 35417
rect 41543 35063 41577 35097
rect 41543 34743 41577 34777
rect 41543 34423 41577 34457
rect 41703 36343 41737 36377
rect 41703 36023 41737 36057
rect 41703 35703 41737 35737
rect 41703 35383 41737 35417
rect 41703 35063 41737 35097
rect 41703 34743 41737 34777
rect 41703 34423 41737 34457
rect 41863 36343 41897 36377
rect 41863 36023 41897 36057
rect 41863 35703 41897 35737
rect 41863 35383 41897 35417
rect 41863 35063 41897 35097
rect 41863 34743 41897 34777
rect 41863 34423 41897 34457
rect 23 34263 57 34297
rect 23 33943 57 33977
rect 183 34263 217 34297
rect 183 33943 217 33977
rect 343 34263 377 34297
rect 343 33943 377 33977
rect 503 34263 537 34297
rect 503 33943 537 33977
rect 663 34263 697 34297
rect 663 33943 697 33977
rect 823 34263 857 34297
rect 823 33943 857 33977
rect 983 34263 1017 34297
rect 983 33943 1017 33977
rect 1143 34263 1177 34297
rect 1143 33943 1177 33977
rect 1303 34263 1337 34297
rect 1303 33943 1337 33977
rect 1463 34263 1497 34297
rect 1463 33943 1497 33977
rect 1623 34263 1657 34297
rect 1623 33943 1657 33977
rect 1783 34263 1817 34297
rect 1783 33943 1817 33977
rect 1943 34263 1977 34297
rect 1943 33943 1977 33977
rect 2103 34263 2137 34297
rect 2103 33943 2137 33977
rect 2263 34263 2297 34297
rect 2263 33943 2297 33977
rect 2423 34263 2457 34297
rect 2423 33943 2457 33977
rect 2583 34263 2617 34297
rect 2583 33943 2617 33977
rect 2743 34263 2777 34297
rect 2743 33943 2777 33977
rect 2903 34263 2937 34297
rect 2903 33943 2937 33977
rect 3063 34263 3097 34297
rect 3063 33943 3097 33977
rect 3223 34263 3257 34297
rect 3223 33943 3257 33977
rect 3383 34263 3417 34297
rect 3383 33943 3417 33977
rect 3543 34263 3577 34297
rect 3543 33943 3577 33977
rect 3703 34263 3737 34297
rect 3703 33943 3737 33977
rect 3863 34263 3897 34297
rect 3863 33943 3897 33977
rect 4023 34263 4057 34297
rect 4023 33943 4057 33977
rect 4183 34263 4217 34297
rect 4183 33943 4217 33977
rect 4343 34263 4377 34297
rect 4343 33943 4377 33977
rect 4503 34263 4537 34297
rect 4503 33943 4537 33977
rect 4663 34263 4697 34297
rect 4663 33943 4697 33977
rect 4823 34263 4857 34297
rect 4823 33943 4857 33977
rect 4983 34263 5017 34297
rect 4983 33943 5017 33977
rect 5143 34263 5177 34297
rect 5143 33943 5177 33977
rect 5303 34263 5337 34297
rect 5303 33943 5337 33977
rect 5463 34263 5497 34297
rect 5463 33943 5497 33977
rect 5623 34263 5657 34297
rect 5623 33943 5657 33977
rect 5783 34263 5817 34297
rect 5783 33943 5817 33977
rect 5943 34263 5977 34297
rect 5943 33943 5977 33977
rect 6103 34263 6137 34297
rect 6103 33943 6137 33977
rect 6263 34263 6297 34297
rect 6263 33943 6297 33977
rect 6423 34263 6457 34297
rect 6423 33943 6457 33977
rect 6583 34263 6617 34297
rect 6583 33943 6617 33977
rect 6743 34263 6777 34297
rect 6743 33943 6777 33977
rect 6903 34263 6937 34297
rect 6903 33943 6937 33977
rect 7063 34263 7097 34297
rect 7063 33943 7097 33977
rect 7223 34263 7257 34297
rect 7223 33943 7257 33977
rect 7383 34263 7417 34297
rect 7383 33943 7417 33977
rect 7543 34263 7577 34297
rect 7543 33943 7577 33977
rect 7703 34263 7737 34297
rect 7703 33943 7737 33977
rect 7863 34263 7897 34297
rect 7863 33943 7897 33977
rect 8023 34263 8057 34297
rect 8023 33943 8057 33977
rect 8183 34263 8217 34297
rect 8183 33943 8217 33977
rect 8343 34263 8377 34297
rect 8343 33943 8377 33977
rect 12503 34263 12537 34297
rect 12503 33943 12537 33977
rect 12663 34263 12697 34297
rect 12663 33943 12697 33977
rect 12823 34263 12857 34297
rect 12823 33943 12857 33977
rect 12983 34263 13017 34297
rect 12983 33943 13017 33977
rect 13143 34263 13177 34297
rect 13143 33943 13177 33977
rect 13303 34263 13337 34297
rect 13303 33943 13337 33977
rect 13463 34263 13497 34297
rect 13463 33943 13497 33977
rect 13623 34263 13657 34297
rect 13623 33943 13657 33977
rect 13783 34263 13817 34297
rect 13783 33943 13817 33977
rect 13943 34263 13977 34297
rect 13943 33943 13977 33977
rect 14103 34263 14137 34297
rect 14103 33943 14137 33977
rect 14263 34263 14297 34297
rect 14263 33943 14297 33977
rect 14423 34263 14457 34297
rect 14423 33943 14457 33977
rect 14583 34263 14617 34297
rect 14583 33943 14617 33977
rect 14743 34263 14777 34297
rect 14743 33943 14777 33977
rect 14903 34263 14937 34297
rect 14903 33943 14937 33977
rect 15063 34263 15097 34297
rect 15063 33943 15097 33977
rect 15223 34263 15257 34297
rect 15223 33943 15257 33977
rect 15383 34263 15417 34297
rect 15383 33943 15417 33977
rect 15543 34263 15577 34297
rect 15543 33943 15577 33977
rect 15703 34263 15737 34297
rect 15703 33943 15737 33977
rect 15863 34263 15897 34297
rect 15863 33943 15897 33977
rect 16023 34263 16057 34297
rect 16023 33943 16057 33977
rect 16183 34263 16217 34297
rect 16183 33943 16217 33977
rect 16343 34263 16377 34297
rect 16343 33943 16377 33977
rect 16503 34263 16537 34297
rect 16503 33943 16537 33977
rect 16663 34263 16697 34297
rect 16663 33943 16697 33977
rect 16823 34263 16857 34297
rect 16823 33943 16857 33977
rect 16983 34263 17017 34297
rect 16983 33943 17017 33977
rect 17143 34263 17177 34297
rect 17143 33943 17177 33977
rect 17303 34263 17337 34297
rect 17303 33943 17337 33977
rect 17463 34263 17497 34297
rect 17463 33943 17497 33977
rect 17623 34263 17657 34297
rect 17623 33943 17657 33977
rect 17783 34263 17817 34297
rect 17783 33943 17817 33977
rect 17943 34263 17977 34297
rect 17943 33943 17977 33977
rect 18103 34263 18137 34297
rect 18103 33943 18137 33977
rect 18263 34263 18297 34297
rect 18263 33943 18297 33977
rect 18423 34263 18457 34297
rect 18423 33943 18457 33977
rect 18583 34263 18617 34297
rect 18583 33943 18617 33977
rect 18743 34263 18777 34297
rect 18743 33943 18777 33977
rect 18903 34263 18937 34297
rect 18903 33943 18937 33977
rect 23143 34263 23177 34297
rect 23143 33943 23177 33977
rect 23303 34263 23337 34297
rect 23303 33943 23337 33977
rect 23463 34263 23497 34297
rect 23463 33943 23497 33977
rect 23623 34263 23657 34297
rect 23623 33943 23657 33977
rect 23783 34263 23817 34297
rect 23783 33943 23817 33977
rect 23943 34263 23977 34297
rect 23943 33943 23977 33977
rect 24103 34263 24137 34297
rect 24103 33943 24137 33977
rect 24263 34263 24297 34297
rect 24263 33943 24297 33977
rect 24423 34263 24457 34297
rect 24423 33943 24457 33977
rect 24583 34263 24617 34297
rect 24583 33943 24617 33977
rect 24743 34263 24777 34297
rect 24743 33943 24777 33977
rect 24903 34263 24937 34297
rect 24903 33943 24937 33977
rect 25063 34263 25097 34297
rect 25063 33943 25097 33977
rect 25223 34263 25257 34297
rect 25223 33943 25257 33977
rect 25383 34263 25417 34297
rect 25383 33943 25417 33977
rect 25543 34263 25577 34297
rect 25543 33943 25577 33977
rect 25703 34263 25737 34297
rect 25703 33943 25737 33977
rect 25863 34263 25897 34297
rect 25863 33943 25897 33977
rect 26023 34263 26057 34297
rect 26023 33943 26057 33977
rect 26183 34263 26217 34297
rect 26183 33943 26217 33977
rect 26343 34263 26377 34297
rect 26343 33943 26377 33977
rect 26503 34263 26537 34297
rect 26503 33943 26537 33977
rect 26663 34263 26697 34297
rect 26663 33943 26697 33977
rect 26823 34263 26857 34297
rect 26823 33943 26857 33977
rect 26983 34263 27017 34297
rect 26983 33943 27017 33977
rect 27143 34263 27177 34297
rect 27143 33943 27177 33977
rect 27303 34263 27337 34297
rect 27303 33943 27337 33977
rect 27463 34263 27497 34297
rect 27463 33943 27497 33977
rect 27623 34263 27657 34297
rect 27623 33943 27657 33977
rect 27783 34263 27817 34297
rect 27783 33943 27817 33977
rect 27943 34263 27977 34297
rect 27943 33943 27977 33977
rect 28103 34263 28137 34297
rect 28103 33943 28137 33977
rect 28263 34263 28297 34297
rect 28263 33943 28297 33977
rect 28423 34263 28457 34297
rect 28423 33943 28457 33977
rect 28583 34263 28617 34297
rect 28583 33943 28617 33977
rect 28743 34263 28777 34297
rect 28743 33943 28777 33977
rect 28903 34263 28937 34297
rect 28903 33943 28937 33977
rect 29063 34263 29097 34297
rect 29063 33943 29097 33977
rect 29223 34263 29257 34297
rect 29223 33943 29257 33977
rect 29383 34263 29417 34297
rect 29383 33943 29417 33977
rect 33543 34263 33577 34297
rect 33543 33943 33577 33977
rect 33703 34263 33737 34297
rect 33703 33943 33737 33977
rect 33863 34263 33897 34297
rect 33863 33943 33897 33977
rect 34023 34263 34057 34297
rect 34023 33943 34057 33977
rect 34183 34263 34217 34297
rect 34183 33943 34217 33977
rect 34343 34263 34377 34297
rect 34343 33943 34377 33977
rect 34503 34263 34537 34297
rect 34503 33943 34537 33977
rect 34663 34263 34697 34297
rect 34663 33943 34697 33977
rect 34823 34263 34857 34297
rect 34823 33943 34857 33977
rect 34983 34263 35017 34297
rect 34983 33943 35017 33977
rect 35143 34263 35177 34297
rect 35143 33943 35177 33977
rect 35303 34263 35337 34297
rect 35303 33943 35337 33977
rect 35463 34263 35497 34297
rect 35463 33943 35497 33977
rect 35623 34263 35657 34297
rect 35623 33943 35657 33977
rect 35783 34263 35817 34297
rect 35783 33943 35817 33977
rect 35943 34263 35977 34297
rect 35943 33943 35977 33977
rect 36103 34263 36137 34297
rect 36103 33943 36137 33977
rect 36263 34263 36297 34297
rect 36263 33943 36297 33977
rect 36423 34263 36457 34297
rect 36423 33943 36457 33977
rect 36583 34263 36617 34297
rect 36583 33943 36617 33977
rect 36743 34263 36777 34297
rect 36743 33943 36777 33977
rect 36903 34263 36937 34297
rect 36903 33943 36937 33977
rect 37063 34263 37097 34297
rect 37063 33943 37097 33977
rect 37223 34263 37257 34297
rect 37223 33943 37257 33977
rect 37383 34263 37417 34297
rect 37383 33943 37417 33977
rect 37543 34263 37577 34297
rect 37543 33943 37577 33977
rect 37703 34263 37737 34297
rect 37703 33943 37737 33977
rect 37863 34263 37897 34297
rect 37863 33943 37897 33977
rect 38023 34263 38057 34297
rect 38023 33943 38057 33977
rect 38183 34263 38217 34297
rect 38183 33943 38217 33977
rect 38343 34263 38377 34297
rect 38343 33943 38377 33977
rect 38503 34263 38537 34297
rect 38503 33943 38537 33977
rect 38663 34263 38697 34297
rect 38663 33943 38697 33977
rect 38823 34263 38857 34297
rect 38823 33943 38857 33977
rect 38983 34263 39017 34297
rect 38983 33943 39017 33977
rect 39143 34263 39177 34297
rect 39143 33943 39177 33977
rect 39303 34263 39337 34297
rect 39303 33943 39337 33977
rect 39463 34263 39497 34297
rect 39463 33943 39497 33977
rect 39623 34263 39657 34297
rect 39623 33943 39657 33977
rect 39783 34263 39817 34297
rect 39783 33943 39817 33977
rect 39943 34263 39977 34297
rect 39943 33943 39977 33977
rect 40103 34263 40137 34297
rect 40103 33943 40137 33977
rect 40263 34263 40297 34297
rect 40263 33943 40297 33977
rect 40423 34263 40457 34297
rect 40423 33943 40457 33977
rect 40583 34263 40617 34297
rect 40583 33943 40617 33977
rect 40743 34263 40777 34297
rect 40743 33943 40777 33977
rect 40903 34263 40937 34297
rect 40903 33943 40937 33977
rect 41063 34263 41097 34297
rect 41063 33943 41097 33977
rect 41223 34263 41257 34297
rect 41223 33943 41257 33977
rect 41383 34263 41417 34297
rect 41383 33943 41417 33977
rect 41543 34263 41577 34297
rect 41543 33943 41577 33977
rect 41703 34263 41737 34297
rect 41703 33943 41737 33977
rect 41863 34263 41897 34297
rect 41863 33943 41897 33977
rect 23 33783 57 33817
rect 23 33463 57 33497
rect 183 33783 217 33817
rect 183 33463 217 33497
rect 343 33783 377 33817
rect 343 33463 377 33497
rect 503 33783 537 33817
rect 503 33463 537 33497
rect 663 33783 697 33817
rect 663 33463 697 33497
rect 823 33783 857 33817
rect 823 33463 857 33497
rect 983 33783 1017 33817
rect 983 33463 1017 33497
rect 1143 33783 1177 33817
rect 1143 33463 1177 33497
rect 1303 33783 1337 33817
rect 1303 33463 1337 33497
rect 1463 33783 1497 33817
rect 1463 33463 1497 33497
rect 1623 33783 1657 33817
rect 1623 33463 1657 33497
rect 1783 33783 1817 33817
rect 1783 33463 1817 33497
rect 1943 33783 1977 33817
rect 1943 33463 1977 33497
rect 2103 33783 2137 33817
rect 2103 33463 2137 33497
rect 2263 33783 2297 33817
rect 2263 33463 2297 33497
rect 2423 33783 2457 33817
rect 2423 33463 2457 33497
rect 2583 33783 2617 33817
rect 2583 33463 2617 33497
rect 2743 33783 2777 33817
rect 2743 33463 2777 33497
rect 2903 33783 2937 33817
rect 2903 33463 2937 33497
rect 3063 33783 3097 33817
rect 3063 33463 3097 33497
rect 3223 33783 3257 33817
rect 3223 33463 3257 33497
rect 3383 33783 3417 33817
rect 3383 33463 3417 33497
rect 3543 33783 3577 33817
rect 3543 33463 3577 33497
rect 3703 33783 3737 33817
rect 3703 33463 3737 33497
rect 3863 33783 3897 33817
rect 3863 33463 3897 33497
rect 4023 33783 4057 33817
rect 4023 33463 4057 33497
rect 4183 33783 4217 33817
rect 4183 33463 4217 33497
rect 4343 33783 4377 33817
rect 4343 33463 4377 33497
rect 4503 33783 4537 33817
rect 4503 33463 4537 33497
rect 4663 33783 4697 33817
rect 4663 33463 4697 33497
rect 4823 33783 4857 33817
rect 4823 33463 4857 33497
rect 4983 33783 5017 33817
rect 4983 33463 5017 33497
rect 5143 33783 5177 33817
rect 5143 33463 5177 33497
rect 5303 33783 5337 33817
rect 5303 33463 5337 33497
rect 5463 33783 5497 33817
rect 5463 33463 5497 33497
rect 5623 33783 5657 33817
rect 5623 33463 5657 33497
rect 5783 33783 5817 33817
rect 5783 33463 5817 33497
rect 5943 33783 5977 33817
rect 5943 33463 5977 33497
rect 6103 33783 6137 33817
rect 6103 33463 6137 33497
rect 6263 33783 6297 33817
rect 6263 33463 6297 33497
rect 6423 33783 6457 33817
rect 6423 33463 6457 33497
rect 6583 33783 6617 33817
rect 6583 33463 6617 33497
rect 6743 33783 6777 33817
rect 6743 33463 6777 33497
rect 6903 33783 6937 33817
rect 6903 33463 6937 33497
rect 7063 33783 7097 33817
rect 7063 33463 7097 33497
rect 7223 33783 7257 33817
rect 7223 33463 7257 33497
rect 7383 33783 7417 33817
rect 7383 33463 7417 33497
rect 7543 33783 7577 33817
rect 7543 33463 7577 33497
rect 7703 33783 7737 33817
rect 7703 33463 7737 33497
rect 7863 33783 7897 33817
rect 7863 33463 7897 33497
rect 8023 33783 8057 33817
rect 8023 33463 8057 33497
rect 8183 33783 8217 33817
rect 8183 33463 8217 33497
rect 8343 33783 8377 33817
rect 8343 33463 8377 33497
rect 12503 33783 12537 33817
rect 12503 33463 12537 33497
rect 12663 33783 12697 33817
rect 12663 33463 12697 33497
rect 12823 33783 12857 33817
rect 12823 33463 12857 33497
rect 12983 33783 13017 33817
rect 12983 33463 13017 33497
rect 13143 33783 13177 33817
rect 13143 33463 13177 33497
rect 13303 33783 13337 33817
rect 13303 33463 13337 33497
rect 13463 33783 13497 33817
rect 13463 33463 13497 33497
rect 13623 33783 13657 33817
rect 13623 33463 13657 33497
rect 13783 33783 13817 33817
rect 13783 33463 13817 33497
rect 13943 33783 13977 33817
rect 13943 33463 13977 33497
rect 14103 33783 14137 33817
rect 14103 33463 14137 33497
rect 14263 33783 14297 33817
rect 14263 33463 14297 33497
rect 14423 33783 14457 33817
rect 14423 33463 14457 33497
rect 14583 33783 14617 33817
rect 14583 33463 14617 33497
rect 14743 33783 14777 33817
rect 14743 33463 14777 33497
rect 14903 33783 14937 33817
rect 14903 33463 14937 33497
rect 15063 33783 15097 33817
rect 15063 33463 15097 33497
rect 15223 33783 15257 33817
rect 15223 33463 15257 33497
rect 15383 33783 15417 33817
rect 15383 33463 15417 33497
rect 15543 33783 15577 33817
rect 15543 33463 15577 33497
rect 15703 33783 15737 33817
rect 15703 33463 15737 33497
rect 15863 33783 15897 33817
rect 15863 33463 15897 33497
rect 16023 33783 16057 33817
rect 16023 33463 16057 33497
rect 16183 33783 16217 33817
rect 16183 33463 16217 33497
rect 16343 33783 16377 33817
rect 16343 33463 16377 33497
rect 16503 33783 16537 33817
rect 16503 33463 16537 33497
rect 16663 33783 16697 33817
rect 16663 33463 16697 33497
rect 16823 33783 16857 33817
rect 16823 33463 16857 33497
rect 16983 33783 17017 33817
rect 16983 33463 17017 33497
rect 17143 33783 17177 33817
rect 17143 33463 17177 33497
rect 17303 33783 17337 33817
rect 17303 33463 17337 33497
rect 17463 33783 17497 33817
rect 17463 33463 17497 33497
rect 17623 33783 17657 33817
rect 17623 33463 17657 33497
rect 17783 33783 17817 33817
rect 17783 33463 17817 33497
rect 17943 33783 17977 33817
rect 17943 33463 17977 33497
rect 18103 33783 18137 33817
rect 18103 33463 18137 33497
rect 18263 33783 18297 33817
rect 18263 33463 18297 33497
rect 18423 33783 18457 33817
rect 18423 33463 18457 33497
rect 18583 33783 18617 33817
rect 18583 33463 18617 33497
rect 18743 33783 18777 33817
rect 18743 33463 18777 33497
rect 18903 33783 18937 33817
rect 18903 33463 18937 33497
rect 23143 33783 23177 33817
rect 23143 33463 23177 33497
rect 23303 33783 23337 33817
rect 23303 33463 23337 33497
rect 23463 33783 23497 33817
rect 23463 33463 23497 33497
rect 23623 33783 23657 33817
rect 23623 33463 23657 33497
rect 23783 33783 23817 33817
rect 23783 33463 23817 33497
rect 23943 33783 23977 33817
rect 23943 33463 23977 33497
rect 24103 33783 24137 33817
rect 24103 33463 24137 33497
rect 24263 33783 24297 33817
rect 24263 33463 24297 33497
rect 24423 33783 24457 33817
rect 24423 33463 24457 33497
rect 24583 33783 24617 33817
rect 24583 33463 24617 33497
rect 24743 33783 24777 33817
rect 24743 33463 24777 33497
rect 24903 33783 24937 33817
rect 24903 33463 24937 33497
rect 25063 33783 25097 33817
rect 25063 33463 25097 33497
rect 25223 33783 25257 33817
rect 25223 33463 25257 33497
rect 25383 33783 25417 33817
rect 25383 33463 25417 33497
rect 25543 33783 25577 33817
rect 25543 33463 25577 33497
rect 25703 33783 25737 33817
rect 25703 33463 25737 33497
rect 25863 33783 25897 33817
rect 25863 33463 25897 33497
rect 26023 33783 26057 33817
rect 26023 33463 26057 33497
rect 26183 33783 26217 33817
rect 26183 33463 26217 33497
rect 26343 33783 26377 33817
rect 26343 33463 26377 33497
rect 26503 33783 26537 33817
rect 26503 33463 26537 33497
rect 26663 33783 26697 33817
rect 26663 33463 26697 33497
rect 26823 33783 26857 33817
rect 26823 33463 26857 33497
rect 26983 33783 27017 33817
rect 26983 33463 27017 33497
rect 27143 33783 27177 33817
rect 27143 33463 27177 33497
rect 27303 33783 27337 33817
rect 27303 33463 27337 33497
rect 27463 33783 27497 33817
rect 27463 33463 27497 33497
rect 27623 33783 27657 33817
rect 27623 33463 27657 33497
rect 27783 33783 27817 33817
rect 27783 33463 27817 33497
rect 27943 33783 27977 33817
rect 27943 33463 27977 33497
rect 28103 33783 28137 33817
rect 28103 33463 28137 33497
rect 28263 33783 28297 33817
rect 28263 33463 28297 33497
rect 28423 33783 28457 33817
rect 28423 33463 28457 33497
rect 28583 33783 28617 33817
rect 28583 33463 28617 33497
rect 28743 33783 28777 33817
rect 28743 33463 28777 33497
rect 28903 33783 28937 33817
rect 28903 33463 28937 33497
rect 29063 33783 29097 33817
rect 29063 33463 29097 33497
rect 29223 33783 29257 33817
rect 29223 33463 29257 33497
rect 29383 33783 29417 33817
rect 29383 33463 29417 33497
rect 33543 33783 33577 33817
rect 33543 33463 33577 33497
rect 33703 33783 33737 33817
rect 33703 33463 33737 33497
rect 33863 33783 33897 33817
rect 33863 33463 33897 33497
rect 34023 33783 34057 33817
rect 34023 33463 34057 33497
rect 34183 33783 34217 33817
rect 34183 33463 34217 33497
rect 34343 33783 34377 33817
rect 34343 33463 34377 33497
rect 34503 33783 34537 33817
rect 34503 33463 34537 33497
rect 34663 33783 34697 33817
rect 34663 33463 34697 33497
rect 34823 33783 34857 33817
rect 34823 33463 34857 33497
rect 34983 33783 35017 33817
rect 34983 33463 35017 33497
rect 35143 33783 35177 33817
rect 35143 33463 35177 33497
rect 35303 33783 35337 33817
rect 35303 33463 35337 33497
rect 35463 33783 35497 33817
rect 35463 33463 35497 33497
rect 35623 33783 35657 33817
rect 35623 33463 35657 33497
rect 35783 33783 35817 33817
rect 35783 33463 35817 33497
rect 35943 33783 35977 33817
rect 35943 33463 35977 33497
rect 36103 33783 36137 33817
rect 36103 33463 36137 33497
rect 36263 33783 36297 33817
rect 36263 33463 36297 33497
rect 36423 33783 36457 33817
rect 36423 33463 36457 33497
rect 36583 33783 36617 33817
rect 36583 33463 36617 33497
rect 36743 33783 36777 33817
rect 36743 33463 36777 33497
rect 36903 33783 36937 33817
rect 36903 33463 36937 33497
rect 37063 33783 37097 33817
rect 37063 33463 37097 33497
rect 37223 33783 37257 33817
rect 37223 33463 37257 33497
rect 37383 33783 37417 33817
rect 37383 33463 37417 33497
rect 37543 33783 37577 33817
rect 37543 33463 37577 33497
rect 37703 33783 37737 33817
rect 37703 33463 37737 33497
rect 37863 33783 37897 33817
rect 37863 33463 37897 33497
rect 38023 33783 38057 33817
rect 38023 33463 38057 33497
rect 38183 33783 38217 33817
rect 38183 33463 38217 33497
rect 38343 33783 38377 33817
rect 38343 33463 38377 33497
rect 38503 33783 38537 33817
rect 38503 33463 38537 33497
rect 38663 33783 38697 33817
rect 38663 33463 38697 33497
rect 38823 33783 38857 33817
rect 38823 33463 38857 33497
rect 38983 33783 39017 33817
rect 38983 33463 39017 33497
rect 39143 33783 39177 33817
rect 39143 33463 39177 33497
rect 39303 33783 39337 33817
rect 39303 33463 39337 33497
rect 39463 33783 39497 33817
rect 39463 33463 39497 33497
rect 39623 33783 39657 33817
rect 39623 33463 39657 33497
rect 39783 33783 39817 33817
rect 39783 33463 39817 33497
rect 39943 33783 39977 33817
rect 39943 33463 39977 33497
rect 40103 33783 40137 33817
rect 40103 33463 40137 33497
rect 40263 33783 40297 33817
rect 40263 33463 40297 33497
rect 40423 33783 40457 33817
rect 40423 33463 40457 33497
rect 40583 33783 40617 33817
rect 40583 33463 40617 33497
rect 40743 33783 40777 33817
rect 40743 33463 40777 33497
rect 40903 33783 40937 33817
rect 40903 33463 40937 33497
rect 41063 33783 41097 33817
rect 41063 33463 41097 33497
rect 41223 33783 41257 33817
rect 41223 33463 41257 33497
rect 41383 33783 41417 33817
rect 41383 33463 41417 33497
rect 41543 33783 41577 33817
rect 41543 33463 41577 33497
rect 41703 33783 41737 33817
rect 41703 33463 41737 33497
rect 41863 33783 41897 33817
rect 41863 33463 41897 33497
rect 23 33303 57 33337
rect 23 32983 57 33017
rect 183 33303 217 33337
rect 183 32983 217 33017
rect 343 33303 377 33337
rect 343 32983 377 33017
rect 503 33303 537 33337
rect 503 32983 537 33017
rect 663 33303 697 33337
rect 663 32983 697 33017
rect 823 33303 857 33337
rect 823 32983 857 33017
rect 983 33303 1017 33337
rect 983 32983 1017 33017
rect 1143 33303 1177 33337
rect 1143 32983 1177 33017
rect 1303 33303 1337 33337
rect 1303 32983 1337 33017
rect 1463 33303 1497 33337
rect 1463 32983 1497 33017
rect 1623 33303 1657 33337
rect 1623 32983 1657 33017
rect 1783 33303 1817 33337
rect 1783 32983 1817 33017
rect 1943 33303 1977 33337
rect 1943 32983 1977 33017
rect 2103 33303 2137 33337
rect 2103 32983 2137 33017
rect 2263 33303 2297 33337
rect 2263 32983 2297 33017
rect 2423 33303 2457 33337
rect 2423 32983 2457 33017
rect 2583 33303 2617 33337
rect 2583 32983 2617 33017
rect 2743 33303 2777 33337
rect 2743 32983 2777 33017
rect 2903 33303 2937 33337
rect 2903 32983 2937 33017
rect 3063 33303 3097 33337
rect 3063 32983 3097 33017
rect 3223 33303 3257 33337
rect 3223 32983 3257 33017
rect 3383 33303 3417 33337
rect 3383 32983 3417 33017
rect 3543 33303 3577 33337
rect 3543 32983 3577 33017
rect 3703 33303 3737 33337
rect 3703 32983 3737 33017
rect 3863 33303 3897 33337
rect 3863 32983 3897 33017
rect 4023 33303 4057 33337
rect 4023 32983 4057 33017
rect 4183 33303 4217 33337
rect 4183 32983 4217 33017
rect 4343 33303 4377 33337
rect 4343 32983 4377 33017
rect 4503 33303 4537 33337
rect 4503 32983 4537 33017
rect 4663 33303 4697 33337
rect 4663 32983 4697 33017
rect 4823 33303 4857 33337
rect 4823 32983 4857 33017
rect 4983 33303 5017 33337
rect 4983 32983 5017 33017
rect 5143 33303 5177 33337
rect 5143 32983 5177 33017
rect 5303 33303 5337 33337
rect 5303 32983 5337 33017
rect 5463 33303 5497 33337
rect 5463 32983 5497 33017
rect 5623 33303 5657 33337
rect 5623 32983 5657 33017
rect 5783 33303 5817 33337
rect 5783 32983 5817 33017
rect 5943 33303 5977 33337
rect 5943 32983 5977 33017
rect 6103 33303 6137 33337
rect 6103 32983 6137 33017
rect 6263 33303 6297 33337
rect 6263 32983 6297 33017
rect 6423 33303 6457 33337
rect 6423 32983 6457 33017
rect 6583 33303 6617 33337
rect 6583 32983 6617 33017
rect 6743 33303 6777 33337
rect 6743 32983 6777 33017
rect 6903 33303 6937 33337
rect 6903 32983 6937 33017
rect 7063 33303 7097 33337
rect 7063 32983 7097 33017
rect 7223 33303 7257 33337
rect 7223 32983 7257 33017
rect 7383 33303 7417 33337
rect 7383 32983 7417 33017
rect 7543 33303 7577 33337
rect 7543 32983 7577 33017
rect 7703 33303 7737 33337
rect 7703 32983 7737 33017
rect 7863 33303 7897 33337
rect 7863 32983 7897 33017
rect 8023 33303 8057 33337
rect 8023 32983 8057 33017
rect 8183 33303 8217 33337
rect 8183 32983 8217 33017
rect 8343 33303 8377 33337
rect 8343 32983 8377 33017
rect 12503 33303 12537 33337
rect 12503 32983 12537 33017
rect 12663 33303 12697 33337
rect 12663 32983 12697 33017
rect 12823 33303 12857 33337
rect 12823 32983 12857 33017
rect 12983 33303 13017 33337
rect 12983 32983 13017 33017
rect 13143 33303 13177 33337
rect 13143 32983 13177 33017
rect 13303 33303 13337 33337
rect 13303 32983 13337 33017
rect 13463 33303 13497 33337
rect 13463 32983 13497 33017
rect 13623 33303 13657 33337
rect 13623 32983 13657 33017
rect 13783 33303 13817 33337
rect 13783 32983 13817 33017
rect 13943 33303 13977 33337
rect 13943 32983 13977 33017
rect 14103 33303 14137 33337
rect 14103 32983 14137 33017
rect 14263 33303 14297 33337
rect 14263 32983 14297 33017
rect 14423 33303 14457 33337
rect 14423 32983 14457 33017
rect 14583 33303 14617 33337
rect 14583 32983 14617 33017
rect 14743 33303 14777 33337
rect 14743 32983 14777 33017
rect 14903 33303 14937 33337
rect 14903 32983 14937 33017
rect 15063 33303 15097 33337
rect 15063 32983 15097 33017
rect 15223 33303 15257 33337
rect 15223 32983 15257 33017
rect 15383 33303 15417 33337
rect 15383 32983 15417 33017
rect 15543 33303 15577 33337
rect 15543 32983 15577 33017
rect 15703 33303 15737 33337
rect 15703 32983 15737 33017
rect 15863 33303 15897 33337
rect 15863 32983 15897 33017
rect 16023 33303 16057 33337
rect 16023 32983 16057 33017
rect 16183 33303 16217 33337
rect 16183 32983 16217 33017
rect 16343 33303 16377 33337
rect 16343 32983 16377 33017
rect 16503 33303 16537 33337
rect 16503 32983 16537 33017
rect 16663 33303 16697 33337
rect 16663 32983 16697 33017
rect 16823 33303 16857 33337
rect 16823 32983 16857 33017
rect 16983 33303 17017 33337
rect 16983 32983 17017 33017
rect 17143 33303 17177 33337
rect 17143 32983 17177 33017
rect 17303 33303 17337 33337
rect 17303 32983 17337 33017
rect 17463 33303 17497 33337
rect 17463 32983 17497 33017
rect 17623 33303 17657 33337
rect 17623 32983 17657 33017
rect 17783 33303 17817 33337
rect 17783 32983 17817 33017
rect 17943 33303 17977 33337
rect 17943 32983 17977 33017
rect 18103 33303 18137 33337
rect 18103 32983 18137 33017
rect 18263 33303 18297 33337
rect 18263 32983 18297 33017
rect 18423 33303 18457 33337
rect 18423 32983 18457 33017
rect 18583 33303 18617 33337
rect 18583 32983 18617 33017
rect 18743 33303 18777 33337
rect 18743 32983 18777 33017
rect 18903 33303 18937 33337
rect 18903 32983 18937 33017
rect 23143 33303 23177 33337
rect 23143 32983 23177 33017
rect 23303 33303 23337 33337
rect 23303 32983 23337 33017
rect 23463 33303 23497 33337
rect 23463 32983 23497 33017
rect 23623 33303 23657 33337
rect 23623 32983 23657 33017
rect 23783 33303 23817 33337
rect 23783 32983 23817 33017
rect 23943 33303 23977 33337
rect 23943 32983 23977 33017
rect 24103 33303 24137 33337
rect 24103 32983 24137 33017
rect 24263 33303 24297 33337
rect 24263 32983 24297 33017
rect 24423 33303 24457 33337
rect 24423 32983 24457 33017
rect 24583 33303 24617 33337
rect 24583 32983 24617 33017
rect 24743 33303 24777 33337
rect 24743 32983 24777 33017
rect 24903 33303 24937 33337
rect 24903 32983 24937 33017
rect 25063 33303 25097 33337
rect 25063 32983 25097 33017
rect 25223 33303 25257 33337
rect 25223 32983 25257 33017
rect 25383 33303 25417 33337
rect 25383 32983 25417 33017
rect 25543 33303 25577 33337
rect 25543 32983 25577 33017
rect 25703 33303 25737 33337
rect 25703 32983 25737 33017
rect 25863 33303 25897 33337
rect 25863 32983 25897 33017
rect 26023 33303 26057 33337
rect 26023 32983 26057 33017
rect 26183 33303 26217 33337
rect 26183 32983 26217 33017
rect 26343 33303 26377 33337
rect 26343 32983 26377 33017
rect 26503 33303 26537 33337
rect 26503 32983 26537 33017
rect 26663 33303 26697 33337
rect 26663 32983 26697 33017
rect 26823 33303 26857 33337
rect 26823 32983 26857 33017
rect 26983 33303 27017 33337
rect 26983 32983 27017 33017
rect 27143 33303 27177 33337
rect 27143 32983 27177 33017
rect 27303 33303 27337 33337
rect 27303 32983 27337 33017
rect 27463 33303 27497 33337
rect 27463 32983 27497 33017
rect 27623 33303 27657 33337
rect 27623 32983 27657 33017
rect 27783 33303 27817 33337
rect 27783 32983 27817 33017
rect 27943 33303 27977 33337
rect 27943 32983 27977 33017
rect 28103 33303 28137 33337
rect 28103 32983 28137 33017
rect 28263 33303 28297 33337
rect 28263 32983 28297 33017
rect 28423 33303 28457 33337
rect 28423 32983 28457 33017
rect 28583 33303 28617 33337
rect 28583 32983 28617 33017
rect 28743 33303 28777 33337
rect 28743 32983 28777 33017
rect 28903 33303 28937 33337
rect 28903 32983 28937 33017
rect 29063 33303 29097 33337
rect 29063 32983 29097 33017
rect 29223 33303 29257 33337
rect 29223 32983 29257 33017
rect 29383 33303 29417 33337
rect 29383 32983 29417 33017
rect 33543 33303 33577 33337
rect 33543 32983 33577 33017
rect 33703 33303 33737 33337
rect 33703 32983 33737 33017
rect 33863 33303 33897 33337
rect 33863 32983 33897 33017
rect 34023 33303 34057 33337
rect 34023 32983 34057 33017
rect 34183 33303 34217 33337
rect 34183 32983 34217 33017
rect 34343 33303 34377 33337
rect 34343 32983 34377 33017
rect 34503 33303 34537 33337
rect 34503 32983 34537 33017
rect 34663 33303 34697 33337
rect 34663 32983 34697 33017
rect 34823 33303 34857 33337
rect 34823 32983 34857 33017
rect 34983 33303 35017 33337
rect 34983 32983 35017 33017
rect 35143 33303 35177 33337
rect 35143 32983 35177 33017
rect 35303 33303 35337 33337
rect 35303 32983 35337 33017
rect 35463 33303 35497 33337
rect 35463 32983 35497 33017
rect 35623 33303 35657 33337
rect 35623 32983 35657 33017
rect 35783 33303 35817 33337
rect 35783 32983 35817 33017
rect 35943 33303 35977 33337
rect 35943 32983 35977 33017
rect 36103 33303 36137 33337
rect 36103 32983 36137 33017
rect 36263 33303 36297 33337
rect 36263 32983 36297 33017
rect 36423 33303 36457 33337
rect 36423 32983 36457 33017
rect 36583 33303 36617 33337
rect 36583 32983 36617 33017
rect 36743 33303 36777 33337
rect 36743 32983 36777 33017
rect 36903 33303 36937 33337
rect 36903 32983 36937 33017
rect 37063 33303 37097 33337
rect 37063 32983 37097 33017
rect 37223 33303 37257 33337
rect 37223 32983 37257 33017
rect 37383 33303 37417 33337
rect 37383 32983 37417 33017
rect 37543 33303 37577 33337
rect 37543 32983 37577 33017
rect 37703 33303 37737 33337
rect 37703 32983 37737 33017
rect 37863 33303 37897 33337
rect 37863 32983 37897 33017
rect 38023 33303 38057 33337
rect 38023 32983 38057 33017
rect 38183 33303 38217 33337
rect 38183 32983 38217 33017
rect 38343 33303 38377 33337
rect 38343 32983 38377 33017
rect 38503 33303 38537 33337
rect 38503 32983 38537 33017
rect 38663 33303 38697 33337
rect 38663 32983 38697 33017
rect 38823 33303 38857 33337
rect 38823 32983 38857 33017
rect 38983 33303 39017 33337
rect 38983 32983 39017 33017
rect 39143 33303 39177 33337
rect 39143 32983 39177 33017
rect 39303 33303 39337 33337
rect 39303 32983 39337 33017
rect 39463 33303 39497 33337
rect 39463 32983 39497 33017
rect 39623 33303 39657 33337
rect 39623 32983 39657 33017
rect 39783 33303 39817 33337
rect 39783 32983 39817 33017
rect 39943 33303 39977 33337
rect 39943 32983 39977 33017
rect 40103 33303 40137 33337
rect 40103 32983 40137 33017
rect 40263 33303 40297 33337
rect 40263 32983 40297 33017
rect 40423 33303 40457 33337
rect 40423 32983 40457 33017
rect 40583 33303 40617 33337
rect 40583 32983 40617 33017
rect 40743 33303 40777 33337
rect 40743 32983 40777 33017
rect 40903 33303 40937 33337
rect 40903 32983 40937 33017
rect 41063 33303 41097 33337
rect 41063 32983 41097 33017
rect 41223 33303 41257 33337
rect 41223 32983 41257 33017
rect 41383 33303 41417 33337
rect 41383 32983 41417 33017
rect 41543 33303 41577 33337
rect 41543 32983 41577 33017
rect 41703 33303 41737 33337
rect 41703 32983 41737 33017
rect 41863 33303 41897 33337
rect 41863 32983 41897 33017
rect 23 32823 57 32857
rect 23 32503 57 32537
rect 183 32823 217 32857
rect 183 32503 217 32537
rect 343 32823 377 32857
rect 343 32503 377 32537
rect 503 32823 537 32857
rect 503 32503 537 32537
rect 663 32823 697 32857
rect 663 32503 697 32537
rect 823 32823 857 32857
rect 823 32503 857 32537
rect 983 32823 1017 32857
rect 983 32503 1017 32537
rect 1143 32823 1177 32857
rect 1143 32503 1177 32537
rect 1303 32823 1337 32857
rect 1303 32503 1337 32537
rect 1463 32823 1497 32857
rect 1463 32503 1497 32537
rect 1623 32823 1657 32857
rect 1623 32503 1657 32537
rect 1783 32823 1817 32857
rect 1783 32503 1817 32537
rect 1943 32823 1977 32857
rect 1943 32503 1977 32537
rect 2103 32823 2137 32857
rect 2103 32503 2137 32537
rect 2263 32823 2297 32857
rect 2263 32503 2297 32537
rect 2423 32823 2457 32857
rect 2423 32503 2457 32537
rect 2583 32823 2617 32857
rect 2583 32503 2617 32537
rect 2743 32823 2777 32857
rect 2743 32503 2777 32537
rect 2903 32823 2937 32857
rect 2903 32503 2937 32537
rect 3063 32823 3097 32857
rect 3063 32503 3097 32537
rect 3223 32823 3257 32857
rect 3223 32503 3257 32537
rect 3383 32823 3417 32857
rect 3383 32503 3417 32537
rect 3543 32823 3577 32857
rect 3543 32503 3577 32537
rect 3703 32823 3737 32857
rect 3703 32503 3737 32537
rect 3863 32823 3897 32857
rect 3863 32503 3897 32537
rect 4023 32823 4057 32857
rect 4023 32503 4057 32537
rect 4183 32823 4217 32857
rect 4183 32503 4217 32537
rect 4343 32823 4377 32857
rect 4343 32503 4377 32537
rect 4503 32823 4537 32857
rect 4503 32503 4537 32537
rect 4663 32823 4697 32857
rect 4663 32503 4697 32537
rect 4823 32823 4857 32857
rect 4823 32503 4857 32537
rect 4983 32823 5017 32857
rect 4983 32503 5017 32537
rect 5143 32823 5177 32857
rect 5143 32503 5177 32537
rect 5303 32823 5337 32857
rect 5303 32503 5337 32537
rect 5463 32823 5497 32857
rect 5463 32503 5497 32537
rect 5623 32823 5657 32857
rect 5623 32503 5657 32537
rect 5783 32823 5817 32857
rect 5783 32503 5817 32537
rect 5943 32823 5977 32857
rect 5943 32503 5977 32537
rect 6103 32823 6137 32857
rect 6103 32503 6137 32537
rect 6263 32823 6297 32857
rect 6263 32503 6297 32537
rect 6423 32823 6457 32857
rect 6423 32503 6457 32537
rect 6583 32823 6617 32857
rect 6583 32503 6617 32537
rect 6743 32823 6777 32857
rect 6743 32503 6777 32537
rect 6903 32823 6937 32857
rect 6903 32503 6937 32537
rect 7063 32823 7097 32857
rect 7063 32503 7097 32537
rect 7223 32823 7257 32857
rect 7223 32503 7257 32537
rect 7383 32823 7417 32857
rect 7383 32503 7417 32537
rect 7543 32823 7577 32857
rect 7543 32503 7577 32537
rect 7703 32823 7737 32857
rect 7703 32503 7737 32537
rect 7863 32823 7897 32857
rect 7863 32503 7897 32537
rect 8023 32823 8057 32857
rect 8023 32503 8057 32537
rect 8183 32823 8217 32857
rect 8183 32503 8217 32537
rect 8343 32823 8377 32857
rect 8343 32503 8377 32537
rect 12503 32823 12537 32857
rect 12503 32503 12537 32537
rect 12663 32823 12697 32857
rect 12663 32503 12697 32537
rect 12823 32823 12857 32857
rect 12823 32503 12857 32537
rect 12983 32823 13017 32857
rect 12983 32503 13017 32537
rect 13143 32823 13177 32857
rect 13143 32503 13177 32537
rect 13303 32823 13337 32857
rect 13303 32503 13337 32537
rect 13463 32823 13497 32857
rect 13463 32503 13497 32537
rect 13623 32823 13657 32857
rect 13623 32503 13657 32537
rect 13783 32823 13817 32857
rect 13783 32503 13817 32537
rect 13943 32823 13977 32857
rect 13943 32503 13977 32537
rect 14103 32823 14137 32857
rect 14103 32503 14137 32537
rect 14263 32823 14297 32857
rect 14263 32503 14297 32537
rect 14423 32823 14457 32857
rect 14423 32503 14457 32537
rect 14583 32823 14617 32857
rect 14583 32503 14617 32537
rect 14743 32823 14777 32857
rect 14743 32503 14777 32537
rect 14903 32823 14937 32857
rect 14903 32503 14937 32537
rect 15063 32823 15097 32857
rect 15063 32503 15097 32537
rect 15223 32823 15257 32857
rect 15223 32503 15257 32537
rect 15383 32823 15417 32857
rect 15383 32503 15417 32537
rect 15543 32823 15577 32857
rect 15543 32503 15577 32537
rect 15703 32823 15737 32857
rect 15703 32503 15737 32537
rect 15863 32823 15897 32857
rect 15863 32503 15897 32537
rect 16023 32823 16057 32857
rect 16023 32503 16057 32537
rect 16183 32823 16217 32857
rect 16183 32503 16217 32537
rect 16343 32823 16377 32857
rect 16343 32503 16377 32537
rect 16503 32823 16537 32857
rect 16503 32503 16537 32537
rect 16663 32823 16697 32857
rect 16663 32503 16697 32537
rect 16823 32823 16857 32857
rect 16823 32503 16857 32537
rect 16983 32823 17017 32857
rect 16983 32503 17017 32537
rect 17143 32823 17177 32857
rect 17143 32503 17177 32537
rect 17303 32823 17337 32857
rect 17303 32503 17337 32537
rect 17463 32823 17497 32857
rect 17463 32503 17497 32537
rect 17623 32823 17657 32857
rect 17623 32503 17657 32537
rect 17783 32823 17817 32857
rect 17783 32503 17817 32537
rect 17943 32823 17977 32857
rect 17943 32503 17977 32537
rect 18103 32823 18137 32857
rect 18103 32503 18137 32537
rect 18263 32823 18297 32857
rect 18263 32503 18297 32537
rect 18423 32823 18457 32857
rect 18423 32503 18457 32537
rect 18583 32823 18617 32857
rect 18583 32503 18617 32537
rect 18743 32823 18777 32857
rect 18743 32503 18777 32537
rect 18903 32823 18937 32857
rect 18903 32503 18937 32537
rect 23143 32823 23177 32857
rect 23143 32503 23177 32537
rect 23303 32823 23337 32857
rect 23303 32503 23337 32537
rect 23463 32823 23497 32857
rect 23463 32503 23497 32537
rect 23623 32823 23657 32857
rect 23623 32503 23657 32537
rect 23783 32823 23817 32857
rect 23783 32503 23817 32537
rect 23943 32823 23977 32857
rect 23943 32503 23977 32537
rect 24103 32823 24137 32857
rect 24103 32503 24137 32537
rect 24263 32823 24297 32857
rect 24263 32503 24297 32537
rect 24423 32823 24457 32857
rect 24423 32503 24457 32537
rect 24583 32823 24617 32857
rect 24583 32503 24617 32537
rect 24743 32823 24777 32857
rect 24743 32503 24777 32537
rect 24903 32823 24937 32857
rect 24903 32503 24937 32537
rect 25063 32823 25097 32857
rect 25063 32503 25097 32537
rect 25223 32823 25257 32857
rect 25223 32503 25257 32537
rect 25383 32823 25417 32857
rect 25383 32503 25417 32537
rect 25543 32823 25577 32857
rect 25543 32503 25577 32537
rect 25703 32823 25737 32857
rect 25703 32503 25737 32537
rect 25863 32823 25897 32857
rect 25863 32503 25897 32537
rect 26023 32823 26057 32857
rect 26023 32503 26057 32537
rect 26183 32823 26217 32857
rect 26183 32503 26217 32537
rect 26343 32823 26377 32857
rect 26343 32503 26377 32537
rect 26503 32823 26537 32857
rect 26503 32503 26537 32537
rect 26663 32823 26697 32857
rect 26663 32503 26697 32537
rect 26823 32823 26857 32857
rect 26823 32503 26857 32537
rect 26983 32823 27017 32857
rect 26983 32503 27017 32537
rect 27143 32823 27177 32857
rect 27143 32503 27177 32537
rect 27303 32823 27337 32857
rect 27303 32503 27337 32537
rect 27463 32823 27497 32857
rect 27463 32503 27497 32537
rect 27623 32823 27657 32857
rect 27623 32503 27657 32537
rect 27783 32823 27817 32857
rect 27783 32503 27817 32537
rect 27943 32823 27977 32857
rect 27943 32503 27977 32537
rect 28103 32823 28137 32857
rect 28103 32503 28137 32537
rect 28263 32823 28297 32857
rect 28263 32503 28297 32537
rect 28423 32823 28457 32857
rect 28423 32503 28457 32537
rect 28583 32823 28617 32857
rect 28583 32503 28617 32537
rect 28743 32823 28777 32857
rect 28743 32503 28777 32537
rect 28903 32823 28937 32857
rect 28903 32503 28937 32537
rect 29063 32823 29097 32857
rect 29063 32503 29097 32537
rect 29223 32823 29257 32857
rect 29223 32503 29257 32537
rect 29383 32823 29417 32857
rect 29383 32503 29417 32537
rect 33543 32823 33577 32857
rect 33543 32503 33577 32537
rect 33703 32823 33737 32857
rect 33703 32503 33737 32537
rect 33863 32823 33897 32857
rect 33863 32503 33897 32537
rect 34023 32823 34057 32857
rect 34023 32503 34057 32537
rect 34183 32823 34217 32857
rect 34183 32503 34217 32537
rect 34343 32823 34377 32857
rect 34343 32503 34377 32537
rect 34503 32823 34537 32857
rect 34503 32503 34537 32537
rect 34663 32823 34697 32857
rect 34663 32503 34697 32537
rect 34823 32823 34857 32857
rect 34823 32503 34857 32537
rect 34983 32823 35017 32857
rect 34983 32503 35017 32537
rect 35143 32823 35177 32857
rect 35143 32503 35177 32537
rect 35303 32823 35337 32857
rect 35303 32503 35337 32537
rect 35463 32823 35497 32857
rect 35463 32503 35497 32537
rect 35623 32823 35657 32857
rect 35623 32503 35657 32537
rect 35783 32823 35817 32857
rect 35783 32503 35817 32537
rect 35943 32823 35977 32857
rect 35943 32503 35977 32537
rect 36103 32823 36137 32857
rect 36103 32503 36137 32537
rect 36263 32823 36297 32857
rect 36263 32503 36297 32537
rect 36423 32823 36457 32857
rect 36423 32503 36457 32537
rect 36583 32823 36617 32857
rect 36583 32503 36617 32537
rect 36743 32823 36777 32857
rect 36743 32503 36777 32537
rect 36903 32823 36937 32857
rect 36903 32503 36937 32537
rect 37063 32823 37097 32857
rect 37063 32503 37097 32537
rect 37223 32823 37257 32857
rect 37223 32503 37257 32537
rect 37383 32823 37417 32857
rect 37383 32503 37417 32537
rect 37543 32823 37577 32857
rect 37543 32503 37577 32537
rect 37703 32823 37737 32857
rect 37703 32503 37737 32537
rect 37863 32823 37897 32857
rect 37863 32503 37897 32537
rect 38023 32823 38057 32857
rect 38023 32503 38057 32537
rect 38183 32823 38217 32857
rect 38183 32503 38217 32537
rect 38343 32823 38377 32857
rect 38343 32503 38377 32537
rect 38503 32823 38537 32857
rect 38503 32503 38537 32537
rect 38663 32823 38697 32857
rect 38663 32503 38697 32537
rect 38823 32823 38857 32857
rect 38823 32503 38857 32537
rect 38983 32823 39017 32857
rect 38983 32503 39017 32537
rect 39143 32823 39177 32857
rect 39143 32503 39177 32537
rect 39303 32823 39337 32857
rect 39303 32503 39337 32537
rect 39463 32823 39497 32857
rect 39463 32503 39497 32537
rect 39623 32823 39657 32857
rect 39623 32503 39657 32537
rect 39783 32823 39817 32857
rect 39783 32503 39817 32537
rect 39943 32823 39977 32857
rect 39943 32503 39977 32537
rect 40103 32823 40137 32857
rect 40103 32503 40137 32537
rect 40263 32823 40297 32857
rect 40263 32503 40297 32537
rect 40423 32823 40457 32857
rect 40423 32503 40457 32537
rect 40583 32823 40617 32857
rect 40583 32503 40617 32537
rect 40743 32823 40777 32857
rect 40743 32503 40777 32537
rect 40903 32823 40937 32857
rect 40903 32503 40937 32537
rect 41063 32823 41097 32857
rect 41063 32503 41097 32537
rect 41223 32823 41257 32857
rect 41223 32503 41257 32537
rect 41383 32823 41417 32857
rect 41383 32503 41417 32537
rect 41543 32823 41577 32857
rect 41543 32503 41577 32537
rect 41703 32823 41737 32857
rect 41703 32503 41737 32537
rect 41863 32823 41897 32857
rect 41863 32503 41897 32537
rect 23 32343 57 32377
rect 23 32023 57 32057
rect 23 31703 57 31737
rect 23 31383 57 31417
rect 23 31063 57 31097
rect 23 30743 57 30777
rect 23 30423 57 30457
rect 183 32343 217 32377
rect 183 32023 217 32057
rect 183 31703 217 31737
rect 183 31383 217 31417
rect 183 31063 217 31097
rect 183 30743 217 30777
rect 183 30423 217 30457
rect 343 32343 377 32377
rect 343 32023 377 32057
rect 343 31703 377 31737
rect 343 31383 377 31417
rect 343 31063 377 31097
rect 343 30743 377 30777
rect 343 30423 377 30457
rect 503 32343 537 32377
rect 503 32023 537 32057
rect 503 31703 537 31737
rect 503 31383 537 31417
rect 503 31063 537 31097
rect 503 30743 537 30777
rect 503 30423 537 30457
rect 663 32343 697 32377
rect 663 32023 697 32057
rect 663 31703 697 31737
rect 663 31383 697 31417
rect 663 31063 697 31097
rect 663 30743 697 30777
rect 663 30423 697 30457
rect 823 32343 857 32377
rect 823 32023 857 32057
rect 823 31703 857 31737
rect 823 31383 857 31417
rect 823 31063 857 31097
rect 823 30743 857 30777
rect 823 30423 857 30457
rect 983 32343 1017 32377
rect 983 32023 1017 32057
rect 983 31703 1017 31737
rect 983 31383 1017 31417
rect 983 31063 1017 31097
rect 983 30743 1017 30777
rect 983 30423 1017 30457
rect 1143 32343 1177 32377
rect 1143 32023 1177 32057
rect 1143 31703 1177 31737
rect 1143 31383 1177 31417
rect 1143 31063 1177 31097
rect 1143 30743 1177 30777
rect 1143 30423 1177 30457
rect 1303 32343 1337 32377
rect 1303 32023 1337 32057
rect 1303 31703 1337 31737
rect 1303 31383 1337 31417
rect 1303 31063 1337 31097
rect 1303 30743 1337 30777
rect 1303 30423 1337 30457
rect 1463 32343 1497 32377
rect 1463 32023 1497 32057
rect 1463 31703 1497 31737
rect 1463 31383 1497 31417
rect 1463 31063 1497 31097
rect 1463 30743 1497 30777
rect 1463 30423 1497 30457
rect 1623 32343 1657 32377
rect 1623 32023 1657 32057
rect 1623 31703 1657 31737
rect 1623 31383 1657 31417
rect 1623 31063 1657 31097
rect 1623 30743 1657 30777
rect 1623 30423 1657 30457
rect 1783 32343 1817 32377
rect 1783 32023 1817 32057
rect 1783 31703 1817 31737
rect 1783 31383 1817 31417
rect 1783 31063 1817 31097
rect 1783 30743 1817 30777
rect 1783 30423 1817 30457
rect 1943 32343 1977 32377
rect 1943 32023 1977 32057
rect 1943 31703 1977 31737
rect 1943 31383 1977 31417
rect 1943 31063 1977 31097
rect 1943 30743 1977 30777
rect 1943 30423 1977 30457
rect 2103 32343 2137 32377
rect 2103 32023 2137 32057
rect 2103 31703 2137 31737
rect 2103 31383 2137 31417
rect 2103 31063 2137 31097
rect 2103 30743 2137 30777
rect 2103 30423 2137 30457
rect 2263 32343 2297 32377
rect 2263 32023 2297 32057
rect 2263 31703 2297 31737
rect 2263 31383 2297 31417
rect 2263 31063 2297 31097
rect 2263 30743 2297 30777
rect 2263 30423 2297 30457
rect 2423 32343 2457 32377
rect 2423 32023 2457 32057
rect 2423 31703 2457 31737
rect 2423 31383 2457 31417
rect 2423 31063 2457 31097
rect 2423 30743 2457 30777
rect 2423 30423 2457 30457
rect 2583 32343 2617 32377
rect 2583 32023 2617 32057
rect 2583 31703 2617 31737
rect 2583 31383 2617 31417
rect 2583 31063 2617 31097
rect 2583 30743 2617 30777
rect 2583 30423 2617 30457
rect 2743 32343 2777 32377
rect 2743 32023 2777 32057
rect 2743 31703 2777 31737
rect 2743 31383 2777 31417
rect 2743 31063 2777 31097
rect 2743 30743 2777 30777
rect 2743 30423 2777 30457
rect 2903 32343 2937 32377
rect 2903 32023 2937 32057
rect 2903 31703 2937 31737
rect 2903 31383 2937 31417
rect 2903 31063 2937 31097
rect 2903 30743 2937 30777
rect 2903 30423 2937 30457
rect 3063 32343 3097 32377
rect 3063 32023 3097 32057
rect 3063 31703 3097 31737
rect 3063 31383 3097 31417
rect 3063 31063 3097 31097
rect 3063 30743 3097 30777
rect 3063 30423 3097 30457
rect 3223 32343 3257 32377
rect 3223 32023 3257 32057
rect 3223 31703 3257 31737
rect 3223 31383 3257 31417
rect 3223 31063 3257 31097
rect 3223 30743 3257 30777
rect 3223 30423 3257 30457
rect 3383 32343 3417 32377
rect 3383 32023 3417 32057
rect 3383 31703 3417 31737
rect 3383 31383 3417 31417
rect 3383 31063 3417 31097
rect 3383 30743 3417 30777
rect 3383 30423 3417 30457
rect 3543 32343 3577 32377
rect 3543 32023 3577 32057
rect 3543 31703 3577 31737
rect 3543 31383 3577 31417
rect 3543 31063 3577 31097
rect 3543 30743 3577 30777
rect 3543 30423 3577 30457
rect 3703 32343 3737 32377
rect 3703 32023 3737 32057
rect 3703 31703 3737 31737
rect 3703 31383 3737 31417
rect 3703 31063 3737 31097
rect 3703 30743 3737 30777
rect 3703 30423 3737 30457
rect 3863 32343 3897 32377
rect 3863 32023 3897 32057
rect 3863 31703 3897 31737
rect 3863 31383 3897 31417
rect 3863 31063 3897 31097
rect 3863 30743 3897 30777
rect 3863 30423 3897 30457
rect 4023 32343 4057 32377
rect 4023 32023 4057 32057
rect 4023 31703 4057 31737
rect 4023 31383 4057 31417
rect 4023 31063 4057 31097
rect 4023 30743 4057 30777
rect 4023 30423 4057 30457
rect 4183 32343 4217 32377
rect 4183 32023 4217 32057
rect 4183 31703 4217 31737
rect 4183 31383 4217 31417
rect 4183 31063 4217 31097
rect 4183 30743 4217 30777
rect 4183 30423 4217 30457
rect 4343 32343 4377 32377
rect 4343 32023 4377 32057
rect 4343 31703 4377 31737
rect 4343 31383 4377 31417
rect 4343 31063 4377 31097
rect 4343 30743 4377 30777
rect 4343 30423 4377 30457
rect 4503 32343 4537 32377
rect 4503 32023 4537 32057
rect 4503 31703 4537 31737
rect 4503 31383 4537 31417
rect 4503 31063 4537 31097
rect 4503 30743 4537 30777
rect 4503 30423 4537 30457
rect 4663 32343 4697 32377
rect 4663 32023 4697 32057
rect 4663 31703 4697 31737
rect 4663 31383 4697 31417
rect 4663 31063 4697 31097
rect 4663 30743 4697 30777
rect 4663 30423 4697 30457
rect 4823 32343 4857 32377
rect 4823 32023 4857 32057
rect 4823 31703 4857 31737
rect 4823 31383 4857 31417
rect 4823 31063 4857 31097
rect 4823 30743 4857 30777
rect 4823 30423 4857 30457
rect 4983 32343 5017 32377
rect 4983 32023 5017 32057
rect 4983 31703 5017 31737
rect 4983 31383 5017 31417
rect 4983 31063 5017 31097
rect 4983 30743 5017 30777
rect 4983 30423 5017 30457
rect 5143 32343 5177 32377
rect 5143 32023 5177 32057
rect 5143 31703 5177 31737
rect 5143 31383 5177 31417
rect 5143 31063 5177 31097
rect 5143 30743 5177 30777
rect 5143 30423 5177 30457
rect 5303 32343 5337 32377
rect 5303 32023 5337 32057
rect 5303 31703 5337 31737
rect 5303 31383 5337 31417
rect 5303 31063 5337 31097
rect 5303 30743 5337 30777
rect 5303 30423 5337 30457
rect 5463 32343 5497 32377
rect 5463 32023 5497 32057
rect 5463 31703 5497 31737
rect 5463 31383 5497 31417
rect 5463 31063 5497 31097
rect 5463 30743 5497 30777
rect 5463 30423 5497 30457
rect 5623 32343 5657 32377
rect 5623 32023 5657 32057
rect 5623 31703 5657 31737
rect 5623 31383 5657 31417
rect 5623 31063 5657 31097
rect 5623 30743 5657 30777
rect 5623 30423 5657 30457
rect 5783 32343 5817 32377
rect 5783 32023 5817 32057
rect 5783 31703 5817 31737
rect 5783 31383 5817 31417
rect 5783 31063 5817 31097
rect 5783 30743 5817 30777
rect 5783 30423 5817 30457
rect 5943 32343 5977 32377
rect 5943 32023 5977 32057
rect 5943 31703 5977 31737
rect 5943 31383 5977 31417
rect 5943 31063 5977 31097
rect 5943 30743 5977 30777
rect 5943 30423 5977 30457
rect 6103 32343 6137 32377
rect 6103 32023 6137 32057
rect 6103 31703 6137 31737
rect 6103 31383 6137 31417
rect 6103 31063 6137 31097
rect 6103 30743 6137 30777
rect 6103 30423 6137 30457
rect 6263 32343 6297 32377
rect 6263 32023 6297 32057
rect 6263 31703 6297 31737
rect 6263 31383 6297 31417
rect 6263 31063 6297 31097
rect 6263 30743 6297 30777
rect 6263 30423 6297 30457
rect 6423 32343 6457 32377
rect 6423 32023 6457 32057
rect 6423 31703 6457 31737
rect 6423 31383 6457 31417
rect 6423 31063 6457 31097
rect 6423 30743 6457 30777
rect 6423 30423 6457 30457
rect 6583 32343 6617 32377
rect 6583 32023 6617 32057
rect 6583 31703 6617 31737
rect 6583 31383 6617 31417
rect 6583 31063 6617 31097
rect 6583 30743 6617 30777
rect 6583 30423 6617 30457
rect 6743 32343 6777 32377
rect 6743 32023 6777 32057
rect 6743 31703 6777 31737
rect 6743 31383 6777 31417
rect 6743 31063 6777 31097
rect 6743 30743 6777 30777
rect 6743 30423 6777 30457
rect 6903 32343 6937 32377
rect 6903 32023 6937 32057
rect 6903 31703 6937 31737
rect 6903 31383 6937 31417
rect 6903 31063 6937 31097
rect 6903 30743 6937 30777
rect 6903 30423 6937 30457
rect 7063 32343 7097 32377
rect 7063 32023 7097 32057
rect 7063 31703 7097 31737
rect 7063 31383 7097 31417
rect 7063 31063 7097 31097
rect 7063 30743 7097 30777
rect 7063 30423 7097 30457
rect 7223 32343 7257 32377
rect 7223 32023 7257 32057
rect 7223 31703 7257 31737
rect 7223 31383 7257 31417
rect 7223 31063 7257 31097
rect 7223 30743 7257 30777
rect 7223 30423 7257 30457
rect 7383 32343 7417 32377
rect 7383 32023 7417 32057
rect 7383 31703 7417 31737
rect 7383 31383 7417 31417
rect 7383 31063 7417 31097
rect 7383 30743 7417 30777
rect 7383 30423 7417 30457
rect 7543 32343 7577 32377
rect 7543 32023 7577 32057
rect 7543 31703 7577 31737
rect 7543 31383 7577 31417
rect 7543 31063 7577 31097
rect 7543 30743 7577 30777
rect 7543 30423 7577 30457
rect 7703 32343 7737 32377
rect 7703 32023 7737 32057
rect 7703 31703 7737 31737
rect 7703 31383 7737 31417
rect 7703 31063 7737 31097
rect 7703 30743 7737 30777
rect 7703 30423 7737 30457
rect 7863 32343 7897 32377
rect 7863 32023 7897 32057
rect 7863 31703 7897 31737
rect 7863 31383 7897 31417
rect 7863 31063 7897 31097
rect 7863 30743 7897 30777
rect 7863 30423 7897 30457
rect 8023 32343 8057 32377
rect 8023 32023 8057 32057
rect 8023 31703 8057 31737
rect 8023 31383 8057 31417
rect 8023 31063 8057 31097
rect 8023 30743 8057 30777
rect 8023 30423 8057 30457
rect 8183 32343 8217 32377
rect 8183 32023 8217 32057
rect 8183 31703 8217 31737
rect 8183 31383 8217 31417
rect 8183 31063 8217 31097
rect 8183 30743 8217 30777
rect 8183 30423 8217 30457
rect 8343 32343 8377 32377
rect 8343 32023 8377 32057
rect 8343 31703 8377 31737
rect 8343 31383 8377 31417
rect 8343 31063 8377 31097
rect 8343 30743 8377 30777
rect 8343 30423 8377 30457
rect 12503 32343 12537 32377
rect 12503 32023 12537 32057
rect 12503 31703 12537 31737
rect 12503 31383 12537 31417
rect 12503 31063 12537 31097
rect 12503 30743 12537 30777
rect 12503 30423 12537 30457
rect 12663 32343 12697 32377
rect 12663 32023 12697 32057
rect 12663 31703 12697 31737
rect 12663 31383 12697 31417
rect 12663 31063 12697 31097
rect 12663 30743 12697 30777
rect 12663 30423 12697 30457
rect 12823 32343 12857 32377
rect 12823 32023 12857 32057
rect 12823 31703 12857 31737
rect 12823 31383 12857 31417
rect 12823 31063 12857 31097
rect 12823 30743 12857 30777
rect 12823 30423 12857 30457
rect 12983 32343 13017 32377
rect 12983 32023 13017 32057
rect 12983 31703 13017 31737
rect 12983 31383 13017 31417
rect 12983 31063 13017 31097
rect 12983 30743 13017 30777
rect 12983 30423 13017 30457
rect 13143 32343 13177 32377
rect 13143 32023 13177 32057
rect 13143 31703 13177 31737
rect 13143 31383 13177 31417
rect 13143 31063 13177 31097
rect 13143 30743 13177 30777
rect 13143 30423 13177 30457
rect 13303 32343 13337 32377
rect 13303 32023 13337 32057
rect 13303 31703 13337 31737
rect 13303 31383 13337 31417
rect 13303 31063 13337 31097
rect 13303 30743 13337 30777
rect 13303 30423 13337 30457
rect 13463 32343 13497 32377
rect 13463 32023 13497 32057
rect 13463 31703 13497 31737
rect 13463 31383 13497 31417
rect 13463 31063 13497 31097
rect 13463 30743 13497 30777
rect 13463 30423 13497 30457
rect 13623 32343 13657 32377
rect 13623 32023 13657 32057
rect 13623 31703 13657 31737
rect 13623 31383 13657 31417
rect 13623 31063 13657 31097
rect 13623 30743 13657 30777
rect 13623 30423 13657 30457
rect 13783 32343 13817 32377
rect 13783 32023 13817 32057
rect 13783 31703 13817 31737
rect 13783 31383 13817 31417
rect 13783 31063 13817 31097
rect 13783 30743 13817 30777
rect 13783 30423 13817 30457
rect 13943 32343 13977 32377
rect 13943 32023 13977 32057
rect 13943 31703 13977 31737
rect 13943 31383 13977 31417
rect 13943 31063 13977 31097
rect 13943 30743 13977 30777
rect 13943 30423 13977 30457
rect 14103 32343 14137 32377
rect 14103 32023 14137 32057
rect 14103 31703 14137 31737
rect 14103 31383 14137 31417
rect 14103 31063 14137 31097
rect 14103 30743 14137 30777
rect 14103 30423 14137 30457
rect 14263 32343 14297 32377
rect 14263 32023 14297 32057
rect 14263 31703 14297 31737
rect 14263 31383 14297 31417
rect 14263 31063 14297 31097
rect 14263 30743 14297 30777
rect 14263 30423 14297 30457
rect 14423 32343 14457 32377
rect 14423 32023 14457 32057
rect 14423 31703 14457 31737
rect 14423 31383 14457 31417
rect 14423 31063 14457 31097
rect 14423 30743 14457 30777
rect 14423 30423 14457 30457
rect 14583 32343 14617 32377
rect 14583 32023 14617 32057
rect 14583 31703 14617 31737
rect 14583 31383 14617 31417
rect 14583 31063 14617 31097
rect 14583 30743 14617 30777
rect 14583 30423 14617 30457
rect 14743 32343 14777 32377
rect 14743 32023 14777 32057
rect 14743 31703 14777 31737
rect 14743 31383 14777 31417
rect 14743 31063 14777 31097
rect 14743 30743 14777 30777
rect 14743 30423 14777 30457
rect 14903 32343 14937 32377
rect 14903 32023 14937 32057
rect 14903 31703 14937 31737
rect 14903 31383 14937 31417
rect 14903 31063 14937 31097
rect 14903 30743 14937 30777
rect 14903 30423 14937 30457
rect 15063 32343 15097 32377
rect 15063 32023 15097 32057
rect 15063 31703 15097 31737
rect 15063 31383 15097 31417
rect 15063 31063 15097 31097
rect 15063 30743 15097 30777
rect 15063 30423 15097 30457
rect 15223 32343 15257 32377
rect 15223 32023 15257 32057
rect 15223 31703 15257 31737
rect 15223 31383 15257 31417
rect 15223 31063 15257 31097
rect 15223 30743 15257 30777
rect 15223 30423 15257 30457
rect 15383 32343 15417 32377
rect 15383 32023 15417 32057
rect 15383 31703 15417 31737
rect 15383 31383 15417 31417
rect 15383 31063 15417 31097
rect 15383 30743 15417 30777
rect 15383 30423 15417 30457
rect 15543 32343 15577 32377
rect 15543 32023 15577 32057
rect 15543 31703 15577 31737
rect 15543 31383 15577 31417
rect 15543 31063 15577 31097
rect 15543 30743 15577 30777
rect 15543 30423 15577 30457
rect 15703 32343 15737 32377
rect 15703 32023 15737 32057
rect 15703 31703 15737 31737
rect 15703 31383 15737 31417
rect 15703 31063 15737 31097
rect 15703 30743 15737 30777
rect 15703 30423 15737 30457
rect 15863 32343 15897 32377
rect 15863 32023 15897 32057
rect 15863 31703 15897 31737
rect 15863 31383 15897 31417
rect 15863 31063 15897 31097
rect 15863 30743 15897 30777
rect 15863 30423 15897 30457
rect 16023 32343 16057 32377
rect 16023 32023 16057 32057
rect 16023 31703 16057 31737
rect 16023 31383 16057 31417
rect 16023 31063 16057 31097
rect 16023 30743 16057 30777
rect 16023 30423 16057 30457
rect 16183 32343 16217 32377
rect 16183 32023 16217 32057
rect 16183 31703 16217 31737
rect 16183 31383 16217 31417
rect 16183 31063 16217 31097
rect 16183 30743 16217 30777
rect 16183 30423 16217 30457
rect 16343 32343 16377 32377
rect 16343 32023 16377 32057
rect 16343 31703 16377 31737
rect 16343 31383 16377 31417
rect 16343 31063 16377 31097
rect 16343 30743 16377 30777
rect 16343 30423 16377 30457
rect 16503 32343 16537 32377
rect 16503 32023 16537 32057
rect 16503 31703 16537 31737
rect 16503 31383 16537 31417
rect 16503 31063 16537 31097
rect 16503 30743 16537 30777
rect 16503 30423 16537 30457
rect 16663 32343 16697 32377
rect 16663 32023 16697 32057
rect 16663 31703 16697 31737
rect 16663 31383 16697 31417
rect 16663 31063 16697 31097
rect 16663 30743 16697 30777
rect 16663 30423 16697 30457
rect 16823 32343 16857 32377
rect 16823 32023 16857 32057
rect 16823 31703 16857 31737
rect 16823 31383 16857 31417
rect 16823 31063 16857 31097
rect 16823 30743 16857 30777
rect 16823 30423 16857 30457
rect 16983 32343 17017 32377
rect 16983 32023 17017 32057
rect 16983 31703 17017 31737
rect 16983 31383 17017 31417
rect 16983 31063 17017 31097
rect 16983 30743 17017 30777
rect 16983 30423 17017 30457
rect 17143 32343 17177 32377
rect 17143 32023 17177 32057
rect 17143 31703 17177 31737
rect 17143 31383 17177 31417
rect 17143 31063 17177 31097
rect 17143 30743 17177 30777
rect 17143 30423 17177 30457
rect 17303 32343 17337 32377
rect 17303 32023 17337 32057
rect 17303 31703 17337 31737
rect 17303 31383 17337 31417
rect 17303 31063 17337 31097
rect 17303 30743 17337 30777
rect 17303 30423 17337 30457
rect 17463 32343 17497 32377
rect 17463 32023 17497 32057
rect 17463 31703 17497 31737
rect 17463 31383 17497 31417
rect 17463 31063 17497 31097
rect 17463 30743 17497 30777
rect 17463 30423 17497 30457
rect 17623 32343 17657 32377
rect 17623 32023 17657 32057
rect 17623 31703 17657 31737
rect 17623 31383 17657 31417
rect 17623 31063 17657 31097
rect 17623 30743 17657 30777
rect 17623 30423 17657 30457
rect 17783 32343 17817 32377
rect 17783 32023 17817 32057
rect 17783 31703 17817 31737
rect 17783 31383 17817 31417
rect 17783 31063 17817 31097
rect 17783 30743 17817 30777
rect 17783 30423 17817 30457
rect 17943 32343 17977 32377
rect 17943 32023 17977 32057
rect 17943 31703 17977 31737
rect 17943 31383 17977 31417
rect 17943 31063 17977 31097
rect 17943 30743 17977 30777
rect 17943 30423 17977 30457
rect 18103 32343 18137 32377
rect 18103 32023 18137 32057
rect 18103 31703 18137 31737
rect 18103 31383 18137 31417
rect 18103 31063 18137 31097
rect 18103 30743 18137 30777
rect 18103 30423 18137 30457
rect 18263 32343 18297 32377
rect 18263 32023 18297 32057
rect 18263 31703 18297 31737
rect 18263 31383 18297 31417
rect 18263 31063 18297 31097
rect 18263 30743 18297 30777
rect 18263 30423 18297 30457
rect 18423 32343 18457 32377
rect 18423 32023 18457 32057
rect 18423 31703 18457 31737
rect 18423 31383 18457 31417
rect 18423 31063 18457 31097
rect 18423 30743 18457 30777
rect 18423 30423 18457 30457
rect 18583 32343 18617 32377
rect 18583 32023 18617 32057
rect 18583 31703 18617 31737
rect 18583 31383 18617 31417
rect 18583 31063 18617 31097
rect 18583 30743 18617 30777
rect 18583 30423 18617 30457
rect 18743 32343 18777 32377
rect 18743 32023 18777 32057
rect 18743 31703 18777 31737
rect 18743 31383 18777 31417
rect 18743 31063 18777 31097
rect 18743 30743 18777 30777
rect 18743 30423 18777 30457
rect 18903 32343 18937 32377
rect 18903 32023 18937 32057
rect 18903 31703 18937 31737
rect 18903 31383 18937 31417
rect 18903 31063 18937 31097
rect 18903 30743 18937 30777
rect 18903 30423 18937 30457
rect 23143 32343 23177 32377
rect 23143 32023 23177 32057
rect 23143 31703 23177 31737
rect 23143 31383 23177 31417
rect 23143 31063 23177 31097
rect 23143 30743 23177 30777
rect 23143 30423 23177 30457
rect 23303 32343 23337 32377
rect 23303 32023 23337 32057
rect 23303 31703 23337 31737
rect 23303 31383 23337 31417
rect 23303 31063 23337 31097
rect 23303 30743 23337 30777
rect 23303 30423 23337 30457
rect 23463 32343 23497 32377
rect 23463 32023 23497 32057
rect 23463 31703 23497 31737
rect 23463 31383 23497 31417
rect 23463 31063 23497 31097
rect 23463 30743 23497 30777
rect 23463 30423 23497 30457
rect 23623 32343 23657 32377
rect 23623 32023 23657 32057
rect 23623 31703 23657 31737
rect 23623 31383 23657 31417
rect 23623 31063 23657 31097
rect 23623 30743 23657 30777
rect 23623 30423 23657 30457
rect 23783 32343 23817 32377
rect 23783 32023 23817 32057
rect 23783 31703 23817 31737
rect 23783 31383 23817 31417
rect 23783 31063 23817 31097
rect 23783 30743 23817 30777
rect 23783 30423 23817 30457
rect 23943 32343 23977 32377
rect 23943 32023 23977 32057
rect 23943 31703 23977 31737
rect 23943 31383 23977 31417
rect 23943 31063 23977 31097
rect 23943 30743 23977 30777
rect 23943 30423 23977 30457
rect 24103 32343 24137 32377
rect 24103 32023 24137 32057
rect 24103 31703 24137 31737
rect 24103 31383 24137 31417
rect 24103 31063 24137 31097
rect 24103 30743 24137 30777
rect 24103 30423 24137 30457
rect 24263 32343 24297 32377
rect 24263 32023 24297 32057
rect 24263 31703 24297 31737
rect 24263 31383 24297 31417
rect 24263 31063 24297 31097
rect 24263 30743 24297 30777
rect 24263 30423 24297 30457
rect 24423 32343 24457 32377
rect 24423 32023 24457 32057
rect 24423 31703 24457 31737
rect 24423 31383 24457 31417
rect 24423 31063 24457 31097
rect 24423 30743 24457 30777
rect 24423 30423 24457 30457
rect 24583 32343 24617 32377
rect 24583 32023 24617 32057
rect 24583 31703 24617 31737
rect 24583 31383 24617 31417
rect 24583 31063 24617 31097
rect 24583 30743 24617 30777
rect 24583 30423 24617 30457
rect 24743 32343 24777 32377
rect 24743 32023 24777 32057
rect 24743 31703 24777 31737
rect 24743 31383 24777 31417
rect 24743 31063 24777 31097
rect 24743 30743 24777 30777
rect 24743 30423 24777 30457
rect 24903 32343 24937 32377
rect 24903 32023 24937 32057
rect 24903 31703 24937 31737
rect 24903 31383 24937 31417
rect 24903 31063 24937 31097
rect 24903 30743 24937 30777
rect 24903 30423 24937 30457
rect 25063 32343 25097 32377
rect 25063 32023 25097 32057
rect 25063 31703 25097 31737
rect 25063 31383 25097 31417
rect 25063 31063 25097 31097
rect 25063 30743 25097 30777
rect 25063 30423 25097 30457
rect 25223 32343 25257 32377
rect 25223 32023 25257 32057
rect 25223 31703 25257 31737
rect 25223 31383 25257 31417
rect 25223 31063 25257 31097
rect 25223 30743 25257 30777
rect 25223 30423 25257 30457
rect 25383 32343 25417 32377
rect 25383 32023 25417 32057
rect 25383 31703 25417 31737
rect 25383 31383 25417 31417
rect 25383 31063 25417 31097
rect 25383 30743 25417 30777
rect 25383 30423 25417 30457
rect 25543 32343 25577 32377
rect 25543 32023 25577 32057
rect 25543 31703 25577 31737
rect 25543 31383 25577 31417
rect 25543 31063 25577 31097
rect 25543 30743 25577 30777
rect 25543 30423 25577 30457
rect 25703 32343 25737 32377
rect 25703 32023 25737 32057
rect 25703 31703 25737 31737
rect 25703 31383 25737 31417
rect 25703 31063 25737 31097
rect 25703 30743 25737 30777
rect 25703 30423 25737 30457
rect 25863 32343 25897 32377
rect 25863 32023 25897 32057
rect 25863 31703 25897 31737
rect 25863 31383 25897 31417
rect 25863 31063 25897 31097
rect 25863 30743 25897 30777
rect 25863 30423 25897 30457
rect 26023 32343 26057 32377
rect 26023 32023 26057 32057
rect 26023 31703 26057 31737
rect 26023 31383 26057 31417
rect 26023 31063 26057 31097
rect 26023 30743 26057 30777
rect 26023 30423 26057 30457
rect 26183 32343 26217 32377
rect 26183 32023 26217 32057
rect 26183 31703 26217 31737
rect 26183 31383 26217 31417
rect 26183 31063 26217 31097
rect 26183 30743 26217 30777
rect 26183 30423 26217 30457
rect 26343 32343 26377 32377
rect 26343 32023 26377 32057
rect 26343 31703 26377 31737
rect 26343 31383 26377 31417
rect 26343 31063 26377 31097
rect 26343 30743 26377 30777
rect 26343 30423 26377 30457
rect 26503 32343 26537 32377
rect 26503 32023 26537 32057
rect 26503 31703 26537 31737
rect 26503 31383 26537 31417
rect 26503 31063 26537 31097
rect 26503 30743 26537 30777
rect 26503 30423 26537 30457
rect 26663 32343 26697 32377
rect 26663 32023 26697 32057
rect 26663 31703 26697 31737
rect 26663 31383 26697 31417
rect 26663 31063 26697 31097
rect 26663 30743 26697 30777
rect 26663 30423 26697 30457
rect 26823 32343 26857 32377
rect 26823 32023 26857 32057
rect 26823 31703 26857 31737
rect 26823 31383 26857 31417
rect 26823 31063 26857 31097
rect 26823 30743 26857 30777
rect 26823 30423 26857 30457
rect 26983 32343 27017 32377
rect 26983 32023 27017 32057
rect 26983 31703 27017 31737
rect 26983 31383 27017 31417
rect 26983 31063 27017 31097
rect 26983 30743 27017 30777
rect 26983 30423 27017 30457
rect 27143 32343 27177 32377
rect 27143 32023 27177 32057
rect 27143 31703 27177 31737
rect 27143 31383 27177 31417
rect 27143 31063 27177 31097
rect 27143 30743 27177 30777
rect 27143 30423 27177 30457
rect 27303 32343 27337 32377
rect 27303 32023 27337 32057
rect 27303 31703 27337 31737
rect 27303 31383 27337 31417
rect 27303 31063 27337 31097
rect 27303 30743 27337 30777
rect 27303 30423 27337 30457
rect 27463 32343 27497 32377
rect 27463 32023 27497 32057
rect 27463 31703 27497 31737
rect 27463 31383 27497 31417
rect 27463 31063 27497 31097
rect 27463 30743 27497 30777
rect 27463 30423 27497 30457
rect 27623 32343 27657 32377
rect 27623 32023 27657 32057
rect 27623 31703 27657 31737
rect 27623 31383 27657 31417
rect 27623 31063 27657 31097
rect 27623 30743 27657 30777
rect 27623 30423 27657 30457
rect 27783 32343 27817 32377
rect 27783 32023 27817 32057
rect 27783 31703 27817 31737
rect 27783 31383 27817 31417
rect 27783 31063 27817 31097
rect 27783 30743 27817 30777
rect 27783 30423 27817 30457
rect 27943 32343 27977 32377
rect 27943 32023 27977 32057
rect 27943 31703 27977 31737
rect 27943 31383 27977 31417
rect 27943 31063 27977 31097
rect 27943 30743 27977 30777
rect 27943 30423 27977 30457
rect 28103 32343 28137 32377
rect 28103 32023 28137 32057
rect 28103 31703 28137 31737
rect 28103 31383 28137 31417
rect 28103 31063 28137 31097
rect 28103 30743 28137 30777
rect 28103 30423 28137 30457
rect 28263 32343 28297 32377
rect 28263 32023 28297 32057
rect 28263 31703 28297 31737
rect 28263 31383 28297 31417
rect 28263 31063 28297 31097
rect 28263 30743 28297 30777
rect 28263 30423 28297 30457
rect 28423 32343 28457 32377
rect 28423 32023 28457 32057
rect 28423 31703 28457 31737
rect 28423 31383 28457 31417
rect 28423 31063 28457 31097
rect 28423 30743 28457 30777
rect 28423 30423 28457 30457
rect 28583 32343 28617 32377
rect 28583 32023 28617 32057
rect 28583 31703 28617 31737
rect 28583 31383 28617 31417
rect 28583 31063 28617 31097
rect 28583 30743 28617 30777
rect 28583 30423 28617 30457
rect 28743 32343 28777 32377
rect 28743 32023 28777 32057
rect 28743 31703 28777 31737
rect 28743 31383 28777 31417
rect 28743 31063 28777 31097
rect 28743 30743 28777 30777
rect 28743 30423 28777 30457
rect 28903 32343 28937 32377
rect 28903 32023 28937 32057
rect 28903 31703 28937 31737
rect 28903 31383 28937 31417
rect 28903 31063 28937 31097
rect 28903 30743 28937 30777
rect 28903 30423 28937 30457
rect 29063 32343 29097 32377
rect 29063 32023 29097 32057
rect 29063 31703 29097 31737
rect 29063 31383 29097 31417
rect 29063 31063 29097 31097
rect 29063 30743 29097 30777
rect 29063 30423 29097 30457
rect 29223 32343 29257 32377
rect 29223 32023 29257 32057
rect 29223 31703 29257 31737
rect 29223 31383 29257 31417
rect 29223 31063 29257 31097
rect 29223 30743 29257 30777
rect 29223 30423 29257 30457
rect 29383 32343 29417 32377
rect 29383 32023 29417 32057
rect 29383 31703 29417 31737
rect 29383 31383 29417 31417
rect 29383 31063 29417 31097
rect 29383 30743 29417 30777
rect 29383 30423 29417 30457
rect 33543 32343 33577 32377
rect 33543 32023 33577 32057
rect 33543 31703 33577 31737
rect 33543 31383 33577 31417
rect 33543 31063 33577 31097
rect 33543 30743 33577 30777
rect 33543 30423 33577 30457
rect 33703 32343 33737 32377
rect 33703 32023 33737 32057
rect 33703 31703 33737 31737
rect 33703 31383 33737 31417
rect 33703 31063 33737 31097
rect 33703 30743 33737 30777
rect 33703 30423 33737 30457
rect 33863 32343 33897 32377
rect 33863 32023 33897 32057
rect 33863 31703 33897 31737
rect 33863 31383 33897 31417
rect 33863 31063 33897 31097
rect 33863 30743 33897 30777
rect 33863 30423 33897 30457
rect 34023 32343 34057 32377
rect 34023 32023 34057 32057
rect 34023 31703 34057 31737
rect 34023 31383 34057 31417
rect 34023 31063 34057 31097
rect 34023 30743 34057 30777
rect 34023 30423 34057 30457
rect 34183 32343 34217 32377
rect 34183 32023 34217 32057
rect 34183 31703 34217 31737
rect 34183 31383 34217 31417
rect 34183 31063 34217 31097
rect 34183 30743 34217 30777
rect 34183 30423 34217 30457
rect 34343 32343 34377 32377
rect 34343 32023 34377 32057
rect 34343 31703 34377 31737
rect 34343 31383 34377 31417
rect 34343 31063 34377 31097
rect 34343 30743 34377 30777
rect 34343 30423 34377 30457
rect 34503 32343 34537 32377
rect 34503 32023 34537 32057
rect 34503 31703 34537 31737
rect 34503 31383 34537 31417
rect 34503 31063 34537 31097
rect 34503 30743 34537 30777
rect 34503 30423 34537 30457
rect 34663 32343 34697 32377
rect 34663 32023 34697 32057
rect 34663 31703 34697 31737
rect 34663 31383 34697 31417
rect 34663 31063 34697 31097
rect 34663 30743 34697 30777
rect 34663 30423 34697 30457
rect 34823 32343 34857 32377
rect 34823 32023 34857 32057
rect 34823 31703 34857 31737
rect 34823 31383 34857 31417
rect 34823 31063 34857 31097
rect 34823 30743 34857 30777
rect 34823 30423 34857 30457
rect 34983 32343 35017 32377
rect 34983 32023 35017 32057
rect 34983 31703 35017 31737
rect 34983 31383 35017 31417
rect 34983 31063 35017 31097
rect 34983 30743 35017 30777
rect 34983 30423 35017 30457
rect 35143 32343 35177 32377
rect 35143 32023 35177 32057
rect 35143 31703 35177 31737
rect 35143 31383 35177 31417
rect 35143 31063 35177 31097
rect 35143 30743 35177 30777
rect 35143 30423 35177 30457
rect 35303 32343 35337 32377
rect 35303 32023 35337 32057
rect 35303 31703 35337 31737
rect 35303 31383 35337 31417
rect 35303 31063 35337 31097
rect 35303 30743 35337 30777
rect 35303 30423 35337 30457
rect 35463 32343 35497 32377
rect 35463 32023 35497 32057
rect 35463 31703 35497 31737
rect 35463 31383 35497 31417
rect 35463 31063 35497 31097
rect 35463 30743 35497 30777
rect 35463 30423 35497 30457
rect 35623 32343 35657 32377
rect 35623 32023 35657 32057
rect 35623 31703 35657 31737
rect 35623 31383 35657 31417
rect 35623 31063 35657 31097
rect 35623 30743 35657 30777
rect 35623 30423 35657 30457
rect 35783 32343 35817 32377
rect 35783 32023 35817 32057
rect 35783 31703 35817 31737
rect 35783 31383 35817 31417
rect 35783 31063 35817 31097
rect 35783 30743 35817 30777
rect 35783 30423 35817 30457
rect 35943 32343 35977 32377
rect 35943 32023 35977 32057
rect 35943 31703 35977 31737
rect 35943 31383 35977 31417
rect 35943 31063 35977 31097
rect 35943 30743 35977 30777
rect 35943 30423 35977 30457
rect 36103 32343 36137 32377
rect 36103 32023 36137 32057
rect 36103 31703 36137 31737
rect 36103 31383 36137 31417
rect 36103 31063 36137 31097
rect 36103 30743 36137 30777
rect 36103 30423 36137 30457
rect 36263 32343 36297 32377
rect 36263 32023 36297 32057
rect 36263 31703 36297 31737
rect 36263 31383 36297 31417
rect 36263 31063 36297 31097
rect 36263 30743 36297 30777
rect 36263 30423 36297 30457
rect 36423 32343 36457 32377
rect 36423 32023 36457 32057
rect 36423 31703 36457 31737
rect 36423 31383 36457 31417
rect 36423 31063 36457 31097
rect 36423 30743 36457 30777
rect 36423 30423 36457 30457
rect 36583 32343 36617 32377
rect 36583 32023 36617 32057
rect 36583 31703 36617 31737
rect 36583 31383 36617 31417
rect 36583 31063 36617 31097
rect 36583 30743 36617 30777
rect 36583 30423 36617 30457
rect 36743 32343 36777 32377
rect 36743 32023 36777 32057
rect 36743 31703 36777 31737
rect 36743 31383 36777 31417
rect 36743 31063 36777 31097
rect 36743 30743 36777 30777
rect 36743 30423 36777 30457
rect 36903 32343 36937 32377
rect 36903 32023 36937 32057
rect 36903 31703 36937 31737
rect 36903 31383 36937 31417
rect 36903 31063 36937 31097
rect 36903 30743 36937 30777
rect 36903 30423 36937 30457
rect 37063 32343 37097 32377
rect 37063 32023 37097 32057
rect 37063 31703 37097 31737
rect 37063 31383 37097 31417
rect 37063 31063 37097 31097
rect 37063 30743 37097 30777
rect 37063 30423 37097 30457
rect 37223 32343 37257 32377
rect 37223 32023 37257 32057
rect 37223 31703 37257 31737
rect 37223 31383 37257 31417
rect 37223 31063 37257 31097
rect 37223 30743 37257 30777
rect 37223 30423 37257 30457
rect 37383 32343 37417 32377
rect 37383 32023 37417 32057
rect 37383 31703 37417 31737
rect 37383 31383 37417 31417
rect 37383 31063 37417 31097
rect 37383 30743 37417 30777
rect 37383 30423 37417 30457
rect 37543 32343 37577 32377
rect 37543 32023 37577 32057
rect 37543 31703 37577 31737
rect 37543 31383 37577 31417
rect 37543 31063 37577 31097
rect 37543 30743 37577 30777
rect 37543 30423 37577 30457
rect 37703 32343 37737 32377
rect 37703 32023 37737 32057
rect 37703 31703 37737 31737
rect 37703 31383 37737 31417
rect 37703 31063 37737 31097
rect 37703 30743 37737 30777
rect 37703 30423 37737 30457
rect 37863 32343 37897 32377
rect 37863 32023 37897 32057
rect 37863 31703 37897 31737
rect 37863 31383 37897 31417
rect 37863 31063 37897 31097
rect 37863 30743 37897 30777
rect 37863 30423 37897 30457
rect 38023 32343 38057 32377
rect 38023 32023 38057 32057
rect 38023 31703 38057 31737
rect 38023 31383 38057 31417
rect 38023 31063 38057 31097
rect 38023 30743 38057 30777
rect 38023 30423 38057 30457
rect 38183 32343 38217 32377
rect 38183 32023 38217 32057
rect 38183 31703 38217 31737
rect 38183 31383 38217 31417
rect 38183 31063 38217 31097
rect 38183 30743 38217 30777
rect 38183 30423 38217 30457
rect 38343 32343 38377 32377
rect 38343 32023 38377 32057
rect 38343 31703 38377 31737
rect 38343 31383 38377 31417
rect 38343 31063 38377 31097
rect 38343 30743 38377 30777
rect 38343 30423 38377 30457
rect 38503 32343 38537 32377
rect 38503 32023 38537 32057
rect 38503 31703 38537 31737
rect 38503 31383 38537 31417
rect 38503 31063 38537 31097
rect 38503 30743 38537 30777
rect 38503 30423 38537 30457
rect 38663 32343 38697 32377
rect 38663 32023 38697 32057
rect 38663 31703 38697 31737
rect 38663 31383 38697 31417
rect 38663 31063 38697 31097
rect 38663 30743 38697 30777
rect 38663 30423 38697 30457
rect 38823 32343 38857 32377
rect 38823 32023 38857 32057
rect 38823 31703 38857 31737
rect 38823 31383 38857 31417
rect 38823 31063 38857 31097
rect 38823 30743 38857 30777
rect 38823 30423 38857 30457
rect 38983 32343 39017 32377
rect 38983 32023 39017 32057
rect 38983 31703 39017 31737
rect 38983 31383 39017 31417
rect 38983 31063 39017 31097
rect 38983 30743 39017 30777
rect 38983 30423 39017 30457
rect 39143 32343 39177 32377
rect 39143 32023 39177 32057
rect 39143 31703 39177 31737
rect 39143 31383 39177 31417
rect 39143 31063 39177 31097
rect 39143 30743 39177 30777
rect 39143 30423 39177 30457
rect 39303 32343 39337 32377
rect 39303 32023 39337 32057
rect 39303 31703 39337 31737
rect 39303 31383 39337 31417
rect 39303 31063 39337 31097
rect 39303 30743 39337 30777
rect 39303 30423 39337 30457
rect 39463 32343 39497 32377
rect 39463 32023 39497 32057
rect 39463 31703 39497 31737
rect 39463 31383 39497 31417
rect 39463 31063 39497 31097
rect 39463 30743 39497 30777
rect 39463 30423 39497 30457
rect 39623 32343 39657 32377
rect 39623 32023 39657 32057
rect 39623 31703 39657 31737
rect 39623 31383 39657 31417
rect 39623 31063 39657 31097
rect 39623 30743 39657 30777
rect 39623 30423 39657 30457
rect 39783 32343 39817 32377
rect 39783 32023 39817 32057
rect 39783 31703 39817 31737
rect 39783 31383 39817 31417
rect 39783 31063 39817 31097
rect 39783 30743 39817 30777
rect 39783 30423 39817 30457
rect 39943 32343 39977 32377
rect 39943 32023 39977 32057
rect 39943 31703 39977 31737
rect 39943 31383 39977 31417
rect 39943 31063 39977 31097
rect 39943 30743 39977 30777
rect 39943 30423 39977 30457
rect 40103 32343 40137 32377
rect 40103 32023 40137 32057
rect 40103 31703 40137 31737
rect 40103 31383 40137 31417
rect 40103 31063 40137 31097
rect 40103 30743 40137 30777
rect 40103 30423 40137 30457
rect 40263 32343 40297 32377
rect 40263 32023 40297 32057
rect 40263 31703 40297 31737
rect 40263 31383 40297 31417
rect 40263 31063 40297 31097
rect 40263 30743 40297 30777
rect 40263 30423 40297 30457
rect 40423 32343 40457 32377
rect 40423 32023 40457 32057
rect 40423 31703 40457 31737
rect 40423 31383 40457 31417
rect 40423 31063 40457 31097
rect 40423 30743 40457 30777
rect 40423 30423 40457 30457
rect 40583 32343 40617 32377
rect 40583 32023 40617 32057
rect 40583 31703 40617 31737
rect 40583 31383 40617 31417
rect 40583 31063 40617 31097
rect 40583 30743 40617 30777
rect 40583 30423 40617 30457
rect 40743 32343 40777 32377
rect 40743 32023 40777 32057
rect 40743 31703 40777 31737
rect 40743 31383 40777 31417
rect 40743 31063 40777 31097
rect 40743 30743 40777 30777
rect 40743 30423 40777 30457
rect 40903 32343 40937 32377
rect 40903 32023 40937 32057
rect 40903 31703 40937 31737
rect 40903 31383 40937 31417
rect 40903 31063 40937 31097
rect 40903 30743 40937 30777
rect 40903 30423 40937 30457
rect 41063 32343 41097 32377
rect 41063 32023 41097 32057
rect 41063 31703 41097 31737
rect 41063 31383 41097 31417
rect 41063 31063 41097 31097
rect 41063 30743 41097 30777
rect 41063 30423 41097 30457
rect 41223 32343 41257 32377
rect 41223 32023 41257 32057
rect 41223 31703 41257 31737
rect 41223 31383 41257 31417
rect 41223 31063 41257 31097
rect 41223 30743 41257 30777
rect 41223 30423 41257 30457
rect 41383 32343 41417 32377
rect 41383 32023 41417 32057
rect 41383 31703 41417 31737
rect 41383 31383 41417 31417
rect 41383 31063 41417 31097
rect 41383 30743 41417 30777
rect 41383 30423 41417 30457
rect 41543 32343 41577 32377
rect 41543 32023 41577 32057
rect 41543 31703 41577 31737
rect 41543 31383 41577 31417
rect 41543 31063 41577 31097
rect 41543 30743 41577 30777
rect 41543 30423 41577 30457
rect 41703 32343 41737 32377
rect 41703 32023 41737 32057
rect 41703 31703 41737 31737
rect 41703 31383 41737 31417
rect 41703 31063 41737 31097
rect 41703 30743 41737 30777
rect 41703 30423 41737 30457
rect 41863 32343 41897 32377
rect 41863 32023 41897 32057
rect 41863 31703 41897 31737
rect 41863 31383 41897 31417
rect 41863 31063 41897 31097
rect 41863 30743 41897 30777
rect 41863 30423 41897 30457
rect 23 30263 57 30297
rect 23 29943 57 29977
rect 183 30263 217 30297
rect 183 29943 217 29977
rect 343 30263 377 30297
rect 343 29943 377 29977
rect 503 30263 537 30297
rect 503 29943 537 29977
rect 663 30263 697 30297
rect 663 29943 697 29977
rect 823 30263 857 30297
rect 823 29943 857 29977
rect 983 30263 1017 30297
rect 983 29943 1017 29977
rect 1143 30263 1177 30297
rect 1143 29943 1177 29977
rect 1303 30263 1337 30297
rect 1303 29943 1337 29977
rect 1463 30263 1497 30297
rect 1463 29943 1497 29977
rect 1623 30263 1657 30297
rect 1623 29943 1657 29977
rect 1783 30263 1817 30297
rect 1783 29943 1817 29977
rect 1943 30263 1977 30297
rect 1943 29943 1977 29977
rect 2103 30263 2137 30297
rect 2103 29943 2137 29977
rect 2263 30263 2297 30297
rect 2263 29943 2297 29977
rect 2423 30263 2457 30297
rect 2423 29943 2457 29977
rect 2583 30263 2617 30297
rect 2583 29943 2617 29977
rect 2743 30263 2777 30297
rect 2743 29943 2777 29977
rect 2903 30263 2937 30297
rect 2903 29943 2937 29977
rect 3063 30263 3097 30297
rect 3063 29943 3097 29977
rect 3223 30263 3257 30297
rect 3223 29943 3257 29977
rect 3383 30263 3417 30297
rect 3383 29943 3417 29977
rect 3543 30263 3577 30297
rect 3543 29943 3577 29977
rect 3703 30263 3737 30297
rect 3703 29943 3737 29977
rect 3863 30263 3897 30297
rect 3863 29943 3897 29977
rect 4023 30263 4057 30297
rect 4023 29943 4057 29977
rect 4183 30263 4217 30297
rect 4183 29943 4217 29977
rect 4343 30263 4377 30297
rect 4343 29943 4377 29977
rect 4503 30263 4537 30297
rect 4503 29943 4537 29977
rect 4663 30263 4697 30297
rect 4663 29943 4697 29977
rect 4823 30263 4857 30297
rect 4823 29943 4857 29977
rect 4983 30263 5017 30297
rect 4983 29943 5017 29977
rect 5143 30263 5177 30297
rect 5143 29943 5177 29977
rect 5303 30263 5337 30297
rect 5303 29943 5337 29977
rect 5463 30263 5497 30297
rect 5463 29943 5497 29977
rect 5623 30263 5657 30297
rect 5623 29943 5657 29977
rect 5783 30263 5817 30297
rect 5783 29943 5817 29977
rect 5943 30263 5977 30297
rect 5943 29943 5977 29977
rect 6103 30263 6137 30297
rect 6103 29943 6137 29977
rect 6263 30263 6297 30297
rect 6263 29943 6297 29977
rect 6423 30263 6457 30297
rect 6423 29943 6457 29977
rect 6583 30263 6617 30297
rect 6583 29943 6617 29977
rect 6743 30263 6777 30297
rect 6743 29943 6777 29977
rect 6903 30263 6937 30297
rect 6903 29943 6937 29977
rect 7063 30263 7097 30297
rect 7063 29943 7097 29977
rect 7223 30263 7257 30297
rect 7223 29943 7257 29977
rect 7383 30263 7417 30297
rect 7383 29943 7417 29977
rect 7543 30263 7577 30297
rect 7543 29943 7577 29977
rect 7703 30263 7737 30297
rect 7703 29943 7737 29977
rect 7863 30263 7897 30297
rect 7863 29943 7897 29977
rect 8023 30263 8057 30297
rect 8023 29943 8057 29977
rect 8183 30263 8217 30297
rect 8183 29943 8217 29977
rect 8343 30263 8377 30297
rect 8343 29943 8377 29977
rect 12503 30263 12537 30297
rect 12503 29943 12537 29977
rect 12663 30263 12697 30297
rect 12663 29943 12697 29977
rect 12823 30263 12857 30297
rect 12823 29943 12857 29977
rect 12983 30263 13017 30297
rect 12983 29943 13017 29977
rect 13143 30263 13177 30297
rect 13143 29943 13177 29977
rect 13303 30263 13337 30297
rect 13303 29943 13337 29977
rect 13463 30263 13497 30297
rect 13463 29943 13497 29977
rect 13623 30263 13657 30297
rect 13623 29943 13657 29977
rect 13783 30263 13817 30297
rect 13783 29943 13817 29977
rect 13943 30263 13977 30297
rect 13943 29943 13977 29977
rect 14103 30263 14137 30297
rect 14103 29943 14137 29977
rect 14263 30263 14297 30297
rect 14263 29943 14297 29977
rect 14423 30263 14457 30297
rect 14423 29943 14457 29977
rect 14583 30263 14617 30297
rect 14583 29943 14617 29977
rect 14743 30263 14777 30297
rect 14743 29943 14777 29977
rect 14903 30263 14937 30297
rect 14903 29943 14937 29977
rect 15063 30263 15097 30297
rect 15063 29943 15097 29977
rect 15223 30263 15257 30297
rect 15223 29943 15257 29977
rect 15383 30263 15417 30297
rect 15383 29943 15417 29977
rect 15543 30263 15577 30297
rect 15543 29943 15577 29977
rect 15703 30263 15737 30297
rect 15703 29943 15737 29977
rect 15863 30263 15897 30297
rect 15863 29943 15897 29977
rect 16023 30263 16057 30297
rect 16023 29943 16057 29977
rect 16183 30263 16217 30297
rect 16183 29943 16217 29977
rect 16343 30263 16377 30297
rect 16343 29943 16377 29977
rect 16503 30263 16537 30297
rect 16503 29943 16537 29977
rect 16663 30263 16697 30297
rect 16663 29943 16697 29977
rect 16823 30263 16857 30297
rect 16823 29943 16857 29977
rect 16983 30263 17017 30297
rect 16983 29943 17017 29977
rect 17143 30263 17177 30297
rect 17143 29943 17177 29977
rect 17303 30263 17337 30297
rect 17303 29943 17337 29977
rect 17463 30263 17497 30297
rect 17463 29943 17497 29977
rect 17623 30263 17657 30297
rect 17623 29943 17657 29977
rect 17783 30263 17817 30297
rect 17783 29943 17817 29977
rect 17943 30263 17977 30297
rect 17943 29943 17977 29977
rect 18103 30263 18137 30297
rect 18103 29943 18137 29977
rect 18263 30263 18297 30297
rect 18263 29943 18297 29977
rect 18423 30263 18457 30297
rect 18423 29943 18457 29977
rect 18583 30263 18617 30297
rect 18583 29943 18617 29977
rect 18743 30263 18777 30297
rect 18743 29943 18777 29977
rect 18903 30263 18937 30297
rect 18903 29943 18937 29977
rect 23143 30263 23177 30297
rect 23143 29943 23177 29977
rect 23303 30263 23337 30297
rect 23303 29943 23337 29977
rect 23463 30263 23497 30297
rect 23463 29943 23497 29977
rect 23623 30263 23657 30297
rect 23623 29943 23657 29977
rect 23783 30263 23817 30297
rect 23783 29943 23817 29977
rect 23943 30263 23977 30297
rect 23943 29943 23977 29977
rect 24103 30263 24137 30297
rect 24103 29943 24137 29977
rect 24263 30263 24297 30297
rect 24263 29943 24297 29977
rect 24423 30263 24457 30297
rect 24423 29943 24457 29977
rect 24583 30263 24617 30297
rect 24583 29943 24617 29977
rect 24743 30263 24777 30297
rect 24743 29943 24777 29977
rect 24903 30263 24937 30297
rect 24903 29943 24937 29977
rect 25063 30263 25097 30297
rect 25063 29943 25097 29977
rect 25223 30263 25257 30297
rect 25223 29943 25257 29977
rect 25383 30263 25417 30297
rect 25383 29943 25417 29977
rect 25543 30263 25577 30297
rect 25543 29943 25577 29977
rect 25703 30263 25737 30297
rect 25703 29943 25737 29977
rect 25863 30263 25897 30297
rect 25863 29943 25897 29977
rect 26023 30263 26057 30297
rect 26023 29943 26057 29977
rect 26183 30263 26217 30297
rect 26183 29943 26217 29977
rect 26343 30263 26377 30297
rect 26343 29943 26377 29977
rect 26503 30263 26537 30297
rect 26503 29943 26537 29977
rect 26663 30263 26697 30297
rect 26663 29943 26697 29977
rect 26823 30263 26857 30297
rect 26823 29943 26857 29977
rect 26983 30263 27017 30297
rect 26983 29943 27017 29977
rect 27143 30263 27177 30297
rect 27143 29943 27177 29977
rect 27303 30263 27337 30297
rect 27303 29943 27337 29977
rect 27463 30263 27497 30297
rect 27463 29943 27497 29977
rect 27623 30263 27657 30297
rect 27623 29943 27657 29977
rect 27783 30263 27817 30297
rect 27783 29943 27817 29977
rect 27943 30263 27977 30297
rect 27943 29943 27977 29977
rect 28103 30263 28137 30297
rect 28103 29943 28137 29977
rect 28263 30263 28297 30297
rect 28263 29943 28297 29977
rect 28423 30263 28457 30297
rect 28423 29943 28457 29977
rect 28583 30263 28617 30297
rect 28583 29943 28617 29977
rect 28743 30263 28777 30297
rect 28743 29943 28777 29977
rect 28903 30263 28937 30297
rect 28903 29943 28937 29977
rect 29063 30263 29097 30297
rect 29063 29943 29097 29977
rect 29223 30263 29257 30297
rect 29223 29943 29257 29977
rect 29383 30263 29417 30297
rect 29383 29943 29417 29977
rect 33543 30263 33577 30297
rect 33543 29943 33577 29977
rect 33703 30263 33737 30297
rect 33703 29943 33737 29977
rect 33863 30263 33897 30297
rect 33863 29943 33897 29977
rect 34023 30263 34057 30297
rect 34023 29943 34057 29977
rect 34183 30263 34217 30297
rect 34183 29943 34217 29977
rect 34343 30263 34377 30297
rect 34343 29943 34377 29977
rect 34503 30263 34537 30297
rect 34503 29943 34537 29977
rect 34663 30263 34697 30297
rect 34663 29943 34697 29977
rect 34823 30263 34857 30297
rect 34823 29943 34857 29977
rect 34983 30263 35017 30297
rect 34983 29943 35017 29977
rect 35143 30263 35177 30297
rect 35143 29943 35177 29977
rect 35303 30263 35337 30297
rect 35303 29943 35337 29977
rect 35463 30263 35497 30297
rect 35463 29943 35497 29977
rect 35623 30263 35657 30297
rect 35623 29943 35657 29977
rect 35783 30263 35817 30297
rect 35783 29943 35817 29977
rect 35943 30263 35977 30297
rect 35943 29943 35977 29977
rect 36103 30263 36137 30297
rect 36103 29943 36137 29977
rect 36263 30263 36297 30297
rect 36263 29943 36297 29977
rect 36423 30263 36457 30297
rect 36423 29943 36457 29977
rect 36583 30263 36617 30297
rect 36583 29943 36617 29977
rect 36743 30263 36777 30297
rect 36743 29943 36777 29977
rect 36903 30263 36937 30297
rect 36903 29943 36937 29977
rect 37063 30263 37097 30297
rect 37063 29943 37097 29977
rect 37223 30263 37257 30297
rect 37223 29943 37257 29977
rect 37383 30263 37417 30297
rect 37383 29943 37417 29977
rect 37543 30263 37577 30297
rect 37543 29943 37577 29977
rect 37703 30263 37737 30297
rect 37703 29943 37737 29977
rect 37863 30263 37897 30297
rect 37863 29943 37897 29977
rect 38023 30263 38057 30297
rect 38023 29943 38057 29977
rect 38183 30263 38217 30297
rect 38183 29943 38217 29977
rect 38343 30263 38377 30297
rect 38343 29943 38377 29977
rect 38503 30263 38537 30297
rect 38503 29943 38537 29977
rect 38663 30263 38697 30297
rect 38663 29943 38697 29977
rect 38823 30263 38857 30297
rect 38823 29943 38857 29977
rect 38983 30263 39017 30297
rect 38983 29943 39017 29977
rect 39143 30263 39177 30297
rect 39143 29943 39177 29977
rect 39303 30263 39337 30297
rect 39303 29943 39337 29977
rect 39463 30263 39497 30297
rect 39463 29943 39497 29977
rect 39623 30263 39657 30297
rect 39623 29943 39657 29977
rect 39783 30263 39817 30297
rect 39783 29943 39817 29977
rect 39943 30263 39977 30297
rect 39943 29943 39977 29977
rect 40103 30263 40137 30297
rect 40103 29943 40137 29977
rect 40263 30263 40297 30297
rect 40263 29943 40297 29977
rect 40423 30263 40457 30297
rect 40423 29943 40457 29977
rect 40583 30263 40617 30297
rect 40583 29943 40617 29977
rect 40743 30263 40777 30297
rect 40743 29943 40777 29977
rect 40903 30263 40937 30297
rect 40903 29943 40937 29977
rect 41063 30263 41097 30297
rect 41063 29943 41097 29977
rect 41223 30263 41257 30297
rect 41223 29943 41257 29977
rect 41383 30263 41417 30297
rect 41383 29943 41417 29977
rect 41543 30263 41577 30297
rect 41543 29943 41577 29977
rect 41703 30263 41737 30297
rect 41703 29943 41737 29977
rect 41863 30263 41897 30297
rect 41863 29943 41897 29977
rect 23 29783 57 29817
rect 23 29463 57 29497
rect 183 29783 217 29817
rect 183 29463 217 29497
rect 343 29783 377 29817
rect 343 29463 377 29497
rect 503 29783 537 29817
rect 503 29463 537 29497
rect 663 29783 697 29817
rect 663 29463 697 29497
rect 823 29783 857 29817
rect 823 29463 857 29497
rect 983 29783 1017 29817
rect 983 29463 1017 29497
rect 1143 29783 1177 29817
rect 1143 29463 1177 29497
rect 1303 29783 1337 29817
rect 1303 29463 1337 29497
rect 1463 29783 1497 29817
rect 1463 29463 1497 29497
rect 1623 29783 1657 29817
rect 1623 29463 1657 29497
rect 1783 29783 1817 29817
rect 1783 29463 1817 29497
rect 1943 29783 1977 29817
rect 1943 29463 1977 29497
rect 2103 29783 2137 29817
rect 2103 29463 2137 29497
rect 2263 29783 2297 29817
rect 2263 29463 2297 29497
rect 2423 29783 2457 29817
rect 2423 29463 2457 29497
rect 2583 29783 2617 29817
rect 2583 29463 2617 29497
rect 2743 29783 2777 29817
rect 2743 29463 2777 29497
rect 2903 29783 2937 29817
rect 2903 29463 2937 29497
rect 3063 29783 3097 29817
rect 3063 29463 3097 29497
rect 3223 29783 3257 29817
rect 3223 29463 3257 29497
rect 3383 29783 3417 29817
rect 3383 29463 3417 29497
rect 3543 29783 3577 29817
rect 3543 29463 3577 29497
rect 3703 29783 3737 29817
rect 3703 29463 3737 29497
rect 3863 29783 3897 29817
rect 3863 29463 3897 29497
rect 4023 29783 4057 29817
rect 4023 29463 4057 29497
rect 4183 29783 4217 29817
rect 4183 29463 4217 29497
rect 4343 29783 4377 29817
rect 4343 29463 4377 29497
rect 4503 29783 4537 29817
rect 4503 29463 4537 29497
rect 4663 29783 4697 29817
rect 4663 29463 4697 29497
rect 4823 29783 4857 29817
rect 4823 29463 4857 29497
rect 4983 29783 5017 29817
rect 4983 29463 5017 29497
rect 5143 29783 5177 29817
rect 5143 29463 5177 29497
rect 5303 29783 5337 29817
rect 5303 29463 5337 29497
rect 5463 29783 5497 29817
rect 5463 29463 5497 29497
rect 5623 29783 5657 29817
rect 5623 29463 5657 29497
rect 5783 29783 5817 29817
rect 5783 29463 5817 29497
rect 5943 29783 5977 29817
rect 5943 29463 5977 29497
rect 6103 29783 6137 29817
rect 6103 29463 6137 29497
rect 6263 29783 6297 29817
rect 6263 29463 6297 29497
rect 6423 29783 6457 29817
rect 6423 29463 6457 29497
rect 6583 29783 6617 29817
rect 6583 29463 6617 29497
rect 6743 29783 6777 29817
rect 6743 29463 6777 29497
rect 6903 29783 6937 29817
rect 6903 29463 6937 29497
rect 7063 29783 7097 29817
rect 7063 29463 7097 29497
rect 7223 29783 7257 29817
rect 7223 29463 7257 29497
rect 7383 29783 7417 29817
rect 7383 29463 7417 29497
rect 7543 29783 7577 29817
rect 7543 29463 7577 29497
rect 7703 29783 7737 29817
rect 7703 29463 7737 29497
rect 7863 29783 7897 29817
rect 7863 29463 7897 29497
rect 8023 29783 8057 29817
rect 8023 29463 8057 29497
rect 8183 29783 8217 29817
rect 8183 29463 8217 29497
rect 8343 29783 8377 29817
rect 8343 29463 8377 29497
rect 12503 29783 12537 29817
rect 12503 29463 12537 29497
rect 12663 29783 12697 29817
rect 12663 29463 12697 29497
rect 12823 29783 12857 29817
rect 12823 29463 12857 29497
rect 12983 29783 13017 29817
rect 12983 29463 13017 29497
rect 13143 29783 13177 29817
rect 13143 29463 13177 29497
rect 13303 29783 13337 29817
rect 13303 29463 13337 29497
rect 13463 29783 13497 29817
rect 13463 29463 13497 29497
rect 13623 29783 13657 29817
rect 13623 29463 13657 29497
rect 13783 29783 13817 29817
rect 13783 29463 13817 29497
rect 13943 29783 13977 29817
rect 13943 29463 13977 29497
rect 14103 29783 14137 29817
rect 14103 29463 14137 29497
rect 14263 29783 14297 29817
rect 14263 29463 14297 29497
rect 14423 29783 14457 29817
rect 14423 29463 14457 29497
rect 14583 29783 14617 29817
rect 14583 29463 14617 29497
rect 14743 29783 14777 29817
rect 14743 29463 14777 29497
rect 14903 29783 14937 29817
rect 14903 29463 14937 29497
rect 15063 29783 15097 29817
rect 15063 29463 15097 29497
rect 15223 29783 15257 29817
rect 15223 29463 15257 29497
rect 15383 29783 15417 29817
rect 15383 29463 15417 29497
rect 15543 29783 15577 29817
rect 15543 29463 15577 29497
rect 15703 29783 15737 29817
rect 15703 29463 15737 29497
rect 15863 29783 15897 29817
rect 15863 29463 15897 29497
rect 16023 29783 16057 29817
rect 16023 29463 16057 29497
rect 16183 29783 16217 29817
rect 16183 29463 16217 29497
rect 16343 29783 16377 29817
rect 16343 29463 16377 29497
rect 16503 29783 16537 29817
rect 16503 29463 16537 29497
rect 16663 29783 16697 29817
rect 16663 29463 16697 29497
rect 16823 29783 16857 29817
rect 16823 29463 16857 29497
rect 16983 29783 17017 29817
rect 16983 29463 17017 29497
rect 17143 29783 17177 29817
rect 17143 29463 17177 29497
rect 17303 29783 17337 29817
rect 17303 29463 17337 29497
rect 17463 29783 17497 29817
rect 17463 29463 17497 29497
rect 17623 29783 17657 29817
rect 17623 29463 17657 29497
rect 17783 29783 17817 29817
rect 17783 29463 17817 29497
rect 17943 29783 17977 29817
rect 17943 29463 17977 29497
rect 18103 29783 18137 29817
rect 18103 29463 18137 29497
rect 18263 29783 18297 29817
rect 18263 29463 18297 29497
rect 18423 29783 18457 29817
rect 18423 29463 18457 29497
rect 18583 29783 18617 29817
rect 18583 29463 18617 29497
rect 18743 29783 18777 29817
rect 18743 29463 18777 29497
rect 18903 29783 18937 29817
rect 18903 29463 18937 29497
rect 23143 29783 23177 29817
rect 23143 29463 23177 29497
rect 23303 29783 23337 29817
rect 23303 29463 23337 29497
rect 23463 29783 23497 29817
rect 23463 29463 23497 29497
rect 23623 29783 23657 29817
rect 23623 29463 23657 29497
rect 23783 29783 23817 29817
rect 23783 29463 23817 29497
rect 23943 29783 23977 29817
rect 23943 29463 23977 29497
rect 24103 29783 24137 29817
rect 24103 29463 24137 29497
rect 24263 29783 24297 29817
rect 24263 29463 24297 29497
rect 24423 29783 24457 29817
rect 24423 29463 24457 29497
rect 24583 29783 24617 29817
rect 24583 29463 24617 29497
rect 24743 29783 24777 29817
rect 24743 29463 24777 29497
rect 24903 29783 24937 29817
rect 24903 29463 24937 29497
rect 25063 29783 25097 29817
rect 25063 29463 25097 29497
rect 25223 29783 25257 29817
rect 25223 29463 25257 29497
rect 25383 29783 25417 29817
rect 25383 29463 25417 29497
rect 25543 29783 25577 29817
rect 25543 29463 25577 29497
rect 25703 29783 25737 29817
rect 25703 29463 25737 29497
rect 25863 29783 25897 29817
rect 25863 29463 25897 29497
rect 26023 29783 26057 29817
rect 26023 29463 26057 29497
rect 26183 29783 26217 29817
rect 26183 29463 26217 29497
rect 26343 29783 26377 29817
rect 26343 29463 26377 29497
rect 26503 29783 26537 29817
rect 26503 29463 26537 29497
rect 26663 29783 26697 29817
rect 26663 29463 26697 29497
rect 26823 29783 26857 29817
rect 26823 29463 26857 29497
rect 26983 29783 27017 29817
rect 26983 29463 27017 29497
rect 27143 29783 27177 29817
rect 27143 29463 27177 29497
rect 27303 29783 27337 29817
rect 27303 29463 27337 29497
rect 27463 29783 27497 29817
rect 27463 29463 27497 29497
rect 27623 29783 27657 29817
rect 27623 29463 27657 29497
rect 27783 29783 27817 29817
rect 27783 29463 27817 29497
rect 27943 29783 27977 29817
rect 27943 29463 27977 29497
rect 28103 29783 28137 29817
rect 28103 29463 28137 29497
rect 28263 29783 28297 29817
rect 28263 29463 28297 29497
rect 28423 29783 28457 29817
rect 28423 29463 28457 29497
rect 28583 29783 28617 29817
rect 28583 29463 28617 29497
rect 28743 29783 28777 29817
rect 28743 29463 28777 29497
rect 28903 29783 28937 29817
rect 28903 29463 28937 29497
rect 29063 29783 29097 29817
rect 29063 29463 29097 29497
rect 29223 29783 29257 29817
rect 29223 29463 29257 29497
rect 29383 29783 29417 29817
rect 29383 29463 29417 29497
rect 33543 29783 33577 29817
rect 33543 29463 33577 29497
rect 33703 29783 33737 29817
rect 33703 29463 33737 29497
rect 33863 29783 33897 29817
rect 33863 29463 33897 29497
rect 34023 29783 34057 29817
rect 34023 29463 34057 29497
rect 34183 29783 34217 29817
rect 34183 29463 34217 29497
rect 34343 29783 34377 29817
rect 34343 29463 34377 29497
rect 34503 29783 34537 29817
rect 34503 29463 34537 29497
rect 34663 29783 34697 29817
rect 34663 29463 34697 29497
rect 34823 29783 34857 29817
rect 34823 29463 34857 29497
rect 34983 29783 35017 29817
rect 34983 29463 35017 29497
rect 35143 29783 35177 29817
rect 35143 29463 35177 29497
rect 35303 29783 35337 29817
rect 35303 29463 35337 29497
rect 35463 29783 35497 29817
rect 35463 29463 35497 29497
rect 35623 29783 35657 29817
rect 35623 29463 35657 29497
rect 35783 29783 35817 29817
rect 35783 29463 35817 29497
rect 35943 29783 35977 29817
rect 35943 29463 35977 29497
rect 36103 29783 36137 29817
rect 36103 29463 36137 29497
rect 36263 29783 36297 29817
rect 36263 29463 36297 29497
rect 36423 29783 36457 29817
rect 36423 29463 36457 29497
rect 36583 29783 36617 29817
rect 36583 29463 36617 29497
rect 36743 29783 36777 29817
rect 36743 29463 36777 29497
rect 36903 29783 36937 29817
rect 36903 29463 36937 29497
rect 37063 29783 37097 29817
rect 37063 29463 37097 29497
rect 37223 29783 37257 29817
rect 37223 29463 37257 29497
rect 37383 29783 37417 29817
rect 37383 29463 37417 29497
rect 37543 29783 37577 29817
rect 37543 29463 37577 29497
rect 37703 29783 37737 29817
rect 37703 29463 37737 29497
rect 37863 29783 37897 29817
rect 37863 29463 37897 29497
rect 38023 29783 38057 29817
rect 38023 29463 38057 29497
rect 38183 29783 38217 29817
rect 38183 29463 38217 29497
rect 38343 29783 38377 29817
rect 38343 29463 38377 29497
rect 38503 29783 38537 29817
rect 38503 29463 38537 29497
rect 38663 29783 38697 29817
rect 38663 29463 38697 29497
rect 38823 29783 38857 29817
rect 38823 29463 38857 29497
rect 38983 29783 39017 29817
rect 38983 29463 39017 29497
rect 39143 29783 39177 29817
rect 39143 29463 39177 29497
rect 39303 29783 39337 29817
rect 39303 29463 39337 29497
rect 39463 29783 39497 29817
rect 39463 29463 39497 29497
rect 39623 29783 39657 29817
rect 39623 29463 39657 29497
rect 39783 29783 39817 29817
rect 39783 29463 39817 29497
rect 39943 29783 39977 29817
rect 39943 29463 39977 29497
rect 40103 29783 40137 29817
rect 40103 29463 40137 29497
rect 40263 29783 40297 29817
rect 40263 29463 40297 29497
rect 40423 29783 40457 29817
rect 40423 29463 40457 29497
rect 40583 29783 40617 29817
rect 40583 29463 40617 29497
rect 40743 29783 40777 29817
rect 40743 29463 40777 29497
rect 40903 29783 40937 29817
rect 40903 29463 40937 29497
rect 41063 29783 41097 29817
rect 41063 29463 41097 29497
rect 41223 29783 41257 29817
rect 41223 29463 41257 29497
rect 41383 29783 41417 29817
rect 41383 29463 41417 29497
rect 41543 29783 41577 29817
rect 41543 29463 41577 29497
rect 41703 29783 41737 29817
rect 41703 29463 41737 29497
rect 41863 29783 41897 29817
rect 41863 29463 41897 29497
<< metal1 >>
rect 0 37346 80 37360
rect 0 37294 14 37346
rect 66 37294 80 37346
rect 0 37280 80 37294
rect 160 37346 240 37360
rect 160 37294 174 37346
rect 226 37294 240 37346
rect 160 37280 240 37294
rect 320 37346 400 37360
rect 320 37294 334 37346
rect 386 37294 400 37346
rect 320 37280 400 37294
rect 480 37346 560 37360
rect 480 37294 494 37346
rect 546 37294 560 37346
rect 480 37280 560 37294
rect 640 37346 720 37360
rect 640 37294 654 37346
rect 706 37294 720 37346
rect 640 37280 720 37294
rect 800 37346 880 37360
rect 800 37294 814 37346
rect 866 37294 880 37346
rect 800 37280 880 37294
rect 960 37346 1040 37360
rect 960 37294 974 37346
rect 1026 37294 1040 37346
rect 960 37280 1040 37294
rect 1120 37346 1200 37360
rect 1120 37294 1134 37346
rect 1186 37294 1200 37346
rect 1120 37280 1200 37294
rect 1280 37346 1360 37360
rect 1280 37294 1294 37346
rect 1346 37294 1360 37346
rect 1280 37280 1360 37294
rect 1440 37346 1520 37360
rect 1440 37294 1454 37346
rect 1506 37294 1520 37346
rect 1440 37280 1520 37294
rect 1600 37346 1680 37360
rect 1600 37294 1614 37346
rect 1666 37294 1680 37346
rect 1600 37280 1680 37294
rect 1760 37346 1840 37360
rect 1760 37294 1774 37346
rect 1826 37294 1840 37346
rect 1760 37280 1840 37294
rect 1920 37346 2000 37360
rect 1920 37294 1934 37346
rect 1986 37294 2000 37346
rect 1920 37280 2000 37294
rect 2080 37346 2160 37360
rect 2080 37294 2094 37346
rect 2146 37294 2160 37346
rect 2080 37280 2160 37294
rect 2240 37346 2320 37360
rect 2240 37294 2254 37346
rect 2306 37294 2320 37346
rect 2240 37280 2320 37294
rect 2400 37346 2480 37360
rect 2400 37294 2414 37346
rect 2466 37294 2480 37346
rect 2400 37280 2480 37294
rect 2560 37346 2640 37360
rect 2560 37294 2574 37346
rect 2626 37294 2640 37346
rect 2560 37280 2640 37294
rect 2720 37346 2800 37360
rect 2720 37294 2734 37346
rect 2786 37294 2800 37346
rect 2720 37280 2800 37294
rect 2880 37346 2960 37360
rect 2880 37294 2894 37346
rect 2946 37294 2960 37346
rect 2880 37280 2960 37294
rect 3040 37346 3120 37360
rect 3040 37294 3054 37346
rect 3106 37294 3120 37346
rect 3040 37280 3120 37294
rect 3200 37346 3280 37360
rect 3200 37294 3214 37346
rect 3266 37294 3280 37346
rect 3200 37280 3280 37294
rect 3360 37346 3440 37360
rect 3360 37294 3374 37346
rect 3426 37294 3440 37346
rect 3360 37280 3440 37294
rect 3520 37346 3600 37360
rect 3520 37294 3534 37346
rect 3586 37294 3600 37346
rect 3520 37280 3600 37294
rect 3680 37346 3760 37360
rect 3680 37294 3694 37346
rect 3746 37294 3760 37346
rect 3680 37280 3760 37294
rect 3840 37346 3920 37360
rect 3840 37294 3854 37346
rect 3906 37294 3920 37346
rect 3840 37280 3920 37294
rect 4000 37346 4080 37360
rect 4000 37294 4014 37346
rect 4066 37294 4080 37346
rect 4000 37280 4080 37294
rect 4160 37346 4240 37360
rect 4160 37294 4174 37346
rect 4226 37294 4240 37346
rect 4160 37280 4240 37294
rect 4320 37346 4400 37360
rect 4320 37294 4334 37346
rect 4386 37294 4400 37346
rect 4320 37280 4400 37294
rect 4480 37346 4560 37360
rect 4480 37294 4494 37346
rect 4546 37294 4560 37346
rect 4480 37280 4560 37294
rect 4640 37346 4720 37360
rect 4640 37294 4654 37346
rect 4706 37294 4720 37346
rect 4640 37280 4720 37294
rect 4800 37346 4880 37360
rect 4800 37294 4814 37346
rect 4866 37294 4880 37346
rect 4800 37280 4880 37294
rect 4960 37346 5040 37360
rect 4960 37294 4974 37346
rect 5026 37294 5040 37346
rect 4960 37280 5040 37294
rect 5120 37346 5200 37360
rect 5120 37294 5134 37346
rect 5186 37294 5200 37346
rect 5120 37280 5200 37294
rect 5280 37346 5360 37360
rect 5280 37294 5294 37346
rect 5346 37294 5360 37346
rect 5280 37280 5360 37294
rect 5440 37346 5520 37360
rect 5440 37294 5454 37346
rect 5506 37294 5520 37346
rect 5440 37280 5520 37294
rect 5600 37346 5680 37360
rect 5600 37294 5614 37346
rect 5666 37294 5680 37346
rect 5600 37280 5680 37294
rect 5760 37346 5840 37360
rect 5760 37294 5774 37346
rect 5826 37294 5840 37346
rect 5760 37280 5840 37294
rect 5920 37346 6000 37360
rect 5920 37294 5934 37346
rect 5986 37294 6000 37346
rect 5920 37280 6000 37294
rect 6080 37346 6160 37360
rect 6080 37294 6094 37346
rect 6146 37294 6160 37346
rect 6080 37280 6160 37294
rect 6240 37346 6320 37360
rect 6240 37294 6254 37346
rect 6306 37294 6320 37346
rect 6240 37280 6320 37294
rect 6400 37346 6480 37360
rect 6400 37294 6414 37346
rect 6466 37294 6480 37346
rect 6400 37280 6480 37294
rect 6560 37346 6640 37360
rect 6560 37294 6574 37346
rect 6626 37294 6640 37346
rect 6560 37280 6640 37294
rect 6720 37346 6800 37360
rect 6720 37294 6734 37346
rect 6786 37294 6800 37346
rect 6720 37280 6800 37294
rect 6880 37346 6960 37360
rect 6880 37294 6894 37346
rect 6946 37294 6960 37346
rect 6880 37280 6960 37294
rect 7040 37346 7120 37360
rect 7040 37294 7054 37346
rect 7106 37294 7120 37346
rect 7040 37280 7120 37294
rect 7200 37346 7280 37360
rect 7200 37294 7214 37346
rect 7266 37294 7280 37346
rect 7200 37280 7280 37294
rect 7360 37346 7440 37360
rect 7360 37294 7374 37346
rect 7426 37294 7440 37346
rect 7360 37280 7440 37294
rect 7520 37346 7600 37360
rect 7520 37294 7534 37346
rect 7586 37294 7600 37346
rect 7520 37280 7600 37294
rect 7680 37346 7760 37360
rect 7680 37294 7694 37346
rect 7746 37294 7760 37346
rect 7680 37280 7760 37294
rect 7840 37346 7920 37360
rect 7840 37294 7854 37346
rect 7906 37294 7920 37346
rect 7840 37280 7920 37294
rect 8000 37346 8080 37360
rect 8000 37294 8014 37346
rect 8066 37294 8080 37346
rect 8000 37280 8080 37294
rect 8160 37346 8240 37360
rect 8160 37294 8174 37346
rect 8226 37294 8240 37346
rect 8160 37280 8240 37294
rect 8320 37346 8400 37360
rect 8320 37294 8334 37346
rect 8386 37294 8400 37346
rect 8320 37280 8400 37294
rect 12480 37346 12560 37360
rect 12480 37294 12494 37346
rect 12546 37294 12560 37346
rect 12480 37280 12560 37294
rect 12640 37346 12720 37360
rect 12640 37294 12654 37346
rect 12706 37294 12720 37346
rect 12640 37280 12720 37294
rect 12800 37346 12880 37360
rect 12800 37294 12814 37346
rect 12866 37294 12880 37346
rect 12800 37280 12880 37294
rect 12960 37346 13040 37360
rect 12960 37294 12974 37346
rect 13026 37294 13040 37346
rect 12960 37280 13040 37294
rect 13120 37346 13200 37360
rect 13120 37294 13134 37346
rect 13186 37294 13200 37346
rect 13120 37280 13200 37294
rect 13280 37346 13360 37360
rect 13280 37294 13294 37346
rect 13346 37294 13360 37346
rect 13280 37280 13360 37294
rect 13440 37346 13520 37360
rect 13440 37294 13454 37346
rect 13506 37294 13520 37346
rect 13440 37280 13520 37294
rect 13600 37346 13680 37360
rect 13600 37294 13614 37346
rect 13666 37294 13680 37346
rect 13600 37280 13680 37294
rect 13760 37346 13840 37360
rect 13760 37294 13774 37346
rect 13826 37294 13840 37346
rect 13760 37280 13840 37294
rect 13920 37346 14000 37360
rect 13920 37294 13934 37346
rect 13986 37294 14000 37346
rect 13920 37280 14000 37294
rect 14080 37346 14160 37360
rect 14080 37294 14094 37346
rect 14146 37294 14160 37346
rect 14080 37280 14160 37294
rect 14240 37346 14320 37360
rect 14240 37294 14254 37346
rect 14306 37294 14320 37346
rect 14240 37280 14320 37294
rect 14400 37346 14480 37360
rect 14400 37294 14414 37346
rect 14466 37294 14480 37346
rect 14400 37280 14480 37294
rect 14560 37346 14640 37360
rect 14560 37294 14574 37346
rect 14626 37294 14640 37346
rect 14560 37280 14640 37294
rect 14720 37346 14800 37360
rect 14720 37294 14734 37346
rect 14786 37294 14800 37346
rect 14720 37280 14800 37294
rect 14880 37346 14960 37360
rect 14880 37294 14894 37346
rect 14946 37294 14960 37346
rect 14880 37280 14960 37294
rect 15040 37346 15120 37360
rect 15040 37294 15054 37346
rect 15106 37294 15120 37346
rect 15040 37280 15120 37294
rect 15200 37346 15280 37360
rect 15200 37294 15214 37346
rect 15266 37294 15280 37346
rect 15200 37280 15280 37294
rect 15360 37346 15440 37360
rect 15360 37294 15374 37346
rect 15426 37294 15440 37346
rect 15360 37280 15440 37294
rect 15520 37346 15600 37360
rect 15520 37294 15534 37346
rect 15586 37294 15600 37346
rect 15520 37280 15600 37294
rect 15680 37346 15760 37360
rect 15680 37294 15694 37346
rect 15746 37294 15760 37346
rect 15680 37280 15760 37294
rect 15840 37346 15920 37360
rect 15840 37294 15854 37346
rect 15906 37294 15920 37346
rect 15840 37280 15920 37294
rect 16000 37346 16080 37360
rect 16000 37294 16014 37346
rect 16066 37294 16080 37346
rect 16000 37280 16080 37294
rect 16160 37346 16240 37360
rect 16160 37294 16174 37346
rect 16226 37294 16240 37346
rect 16160 37280 16240 37294
rect 16320 37346 16400 37360
rect 16320 37294 16334 37346
rect 16386 37294 16400 37346
rect 16320 37280 16400 37294
rect 16480 37346 16560 37360
rect 16480 37294 16494 37346
rect 16546 37294 16560 37346
rect 16480 37280 16560 37294
rect 16640 37346 16720 37360
rect 16640 37294 16654 37346
rect 16706 37294 16720 37346
rect 16640 37280 16720 37294
rect 16800 37346 16880 37360
rect 16800 37294 16814 37346
rect 16866 37294 16880 37346
rect 16800 37280 16880 37294
rect 16960 37346 17040 37360
rect 16960 37294 16974 37346
rect 17026 37294 17040 37346
rect 16960 37280 17040 37294
rect 17120 37346 17200 37360
rect 17120 37294 17134 37346
rect 17186 37294 17200 37346
rect 17120 37280 17200 37294
rect 17280 37346 17360 37360
rect 17280 37294 17294 37346
rect 17346 37294 17360 37346
rect 17280 37280 17360 37294
rect 17440 37346 17520 37360
rect 17440 37294 17454 37346
rect 17506 37294 17520 37346
rect 17440 37280 17520 37294
rect 17600 37346 17680 37360
rect 17600 37294 17614 37346
rect 17666 37294 17680 37346
rect 17600 37280 17680 37294
rect 17760 37346 17840 37360
rect 17760 37294 17774 37346
rect 17826 37294 17840 37346
rect 17760 37280 17840 37294
rect 17920 37346 18000 37360
rect 17920 37294 17934 37346
rect 17986 37294 18000 37346
rect 17920 37280 18000 37294
rect 18080 37346 18160 37360
rect 18080 37294 18094 37346
rect 18146 37294 18160 37346
rect 18080 37280 18160 37294
rect 18240 37346 18320 37360
rect 18240 37294 18254 37346
rect 18306 37294 18320 37346
rect 18240 37280 18320 37294
rect 18400 37346 18480 37360
rect 18400 37294 18414 37346
rect 18466 37294 18480 37346
rect 18400 37280 18480 37294
rect 18560 37346 18640 37360
rect 18560 37294 18574 37346
rect 18626 37294 18640 37346
rect 18560 37280 18640 37294
rect 18720 37346 18800 37360
rect 18720 37294 18734 37346
rect 18786 37294 18800 37346
rect 18720 37280 18800 37294
rect 18880 37346 18960 37360
rect 18880 37294 18894 37346
rect 18946 37294 18960 37346
rect 18880 37280 18960 37294
rect 23120 37346 23200 37360
rect 23120 37294 23134 37346
rect 23186 37294 23200 37346
rect 23120 37280 23200 37294
rect 23280 37346 23360 37360
rect 23280 37294 23294 37346
rect 23346 37294 23360 37346
rect 23280 37280 23360 37294
rect 23440 37346 23520 37360
rect 23440 37294 23454 37346
rect 23506 37294 23520 37346
rect 23440 37280 23520 37294
rect 23600 37346 23680 37360
rect 23600 37294 23614 37346
rect 23666 37294 23680 37346
rect 23600 37280 23680 37294
rect 23760 37346 23840 37360
rect 23760 37294 23774 37346
rect 23826 37294 23840 37346
rect 23760 37280 23840 37294
rect 23920 37346 24000 37360
rect 23920 37294 23934 37346
rect 23986 37294 24000 37346
rect 23920 37280 24000 37294
rect 24080 37346 24160 37360
rect 24080 37294 24094 37346
rect 24146 37294 24160 37346
rect 24080 37280 24160 37294
rect 24240 37346 24320 37360
rect 24240 37294 24254 37346
rect 24306 37294 24320 37346
rect 24240 37280 24320 37294
rect 24400 37346 24480 37360
rect 24400 37294 24414 37346
rect 24466 37294 24480 37346
rect 24400 37280 24480 37294
rect 24560 37346 24640 37360
rect 24560 37294 24574 37346
rect 24626 37294 24640 37346
rect 24560 37280 24640 37294
rect 24720 37346 24800 37360
rect 24720 37294 24734 37346
rect 24786 37294 24800 37346
rect 24720 37280 24800 37294
rect 24880 37346 24960 37360
rect 24880 37294 24894 37346
rect 24946 37294 24960 37346
rect 24880 37280 24960 37294
rect 25040 37346 25120 37360
rect 25040 37294 25054 37346
rect 25106 37294 25120 37346
rect 25040 37280 25120 37294
rect 25200 37346 25280 37360
rect 25200 37294 25214 37346
rect 25266 37294 25280 37346
rect 25200 37280 25280 37294
rect 25360 37346 25440 37360
rect 25360 37294 25374 37346
rect 25426 37294 25440 37346
rect 25360 37280 25440 37294
rect 25520 37346 25600 37360
rect 25520 37294 25534 37346
rect 25586 37294 25600 37346
rect 25520 37280 25600 37294
rect 25680 37346 25760 37360
rect 25680 37294 25694 37346
rect 25746 37294 25760 37346
rect 25680 37280 25760 37294
rect 25840 37346 25920 37360
rect 25840 37294 25854 37346
rect 25906 37294 25920 37346
rect 25840 37280 25920 37294
rect 26000 37346 26080 37360
rect 26000 37294 26014 37346
rect 26066 37294 26080 37346
rect 26000 37280 26080 37294
rect 26160 37346 26240 37360
rect 26160 37294 26174 37346
rect 26226 37294 26240 37346
rect 26160 37280 26240 37294
rect 26320 37346 26400 37360
rect 26320 37294 26334 37346
rect 26386 37294 26400 37346
rect 26320 37280 26400 37294
rect 26480 37346 26560 37360
rect 26480 37294 26494 37346
rect 26546 37294 26560 37346
rect 26480 37280 26560 37294
rect 26640 37346 26720 37360
rect 26640 37294 26654 37346
rect 26706 37294 26720 37346
rect 26640 37280 26720 37294
rect 26800 37346 26880 37360
rect 26800 37294 26814 37346
rect 26866 37294 26880 37346
rect 26800 37280 26880 37294
rect 26960 37346 27040 37360
rect 26960 37294 26974 37346
rect 27026 37294 27040 37346
rect 26960 37280 27040 37294
rect 27120 37346 27200 37360
rect 27120 37294 27134 37346
rect 27186 37294 27200 37346
rect 27120 37280 27200 37294
rect 27280 37346 27360 37360
rect 27280 37294 27294 37346
rect 27346 37294 27360 37346
rect 27280 37280 27360 37294
rect 27440 37346 27520 37360
rect 27440 37294 27454 37346
rect 27506 37294 27520 37346
rect 27440 37280 27520 37294
rect 27600 37346 27680 37360
rect 27600 37294 27614 37346
rect 27666 37294 27680 37346
rect 27600 37280 27680 37294
rect 27760 37346 27840 37360
rect 27760 37294 27774 37346
rect 27826 37294 27840 37346
rect 27760 37280 27840 37294
rect 27920 37346 28000 37360
rect 27920 37294 27934 37346
rect 27986 37294 28000 37346
rect 27920 37280 28000 37294
rect 28080 37346 28160 37360
rect 28080 37294 28094 37346
rect 28146 37294 28160 37346
rect 28080 37280 28160 37294
rect 28240 37346 28320 37360
rect 28240 37294 28254 37346
rect 28306 37294 28320 37346
rect 28240 37280 28320 37294
rect 28400 37346 28480 37360
rect 28400 37294 28414 37346
rect 28466 37294 28480 37346
rect 28400 37280 28480 37294
rect 28560 37346 28640 37360
rect 28560 37294 28574 37346
rect 28626 37294 28640 37346
rect 28560 37280 28640 37294
rect 28720 37346 28800 37360
rect 28720 37294 28734 37346
rect 28786 37294 28800 37346
rect 28720 37280 28800 37294
rect 28880 37346 28960 37360
rect 28880 37294 28894 37346
rect 28946 37294 28960 37346
rect 28880 37280 28960 37294
rect 29040 37346 29120 37360
rect 29040 37294 29054 37346
rect 29106 37294 29120 37346
rect 29040 37280 29120 37294
rect 29200 37346 29280 37360
rect 29200 37294 29214 37346
rect 29266 37294 29280 37346
rect 29200 37280 29280 37294
rect 29360 37346 29440 37360
rect 29360 37294 29374 37346
rect 29426 37294 29440 37346
rect 29360 37280 29440 37294
rect 33520 37346 33600 37360
rect 33520 37294 33534 37346
rect 33586 37294 33600 37346
rect 33520 37280 33600 37294
rect 33680 37346 33760 37360
rect 33680 37294 33694 37346
rect 33746 37294 33760 37346
rect 33680 37280 33760 37294
rect 33840 37346 33920 37360
rect 33840 37294 33854 37346
rect 33906 37294 33920 37346
rect 33840 37280 33920 37294
rect 34000 37346 34080 37360
rect 34000 37294 34014 37346
rect 34066 37294 34080 37346
rect 34000 37280 34080 37294
rect 34160 37346 34240 37360
rect 34160 37294 34174 37346
rect 34226 37294 34240 37346
rect 34160 37280 34240 37294
rect 34320 37346 34400 37360
rect 34320 37294 34334 37346
rect 34386 37294 34400 37346
rect 34320 37280 34400 37294
rect 34480 37346 34560 37360
rect 34480 37294 34494 37346
rect 34546 37294 34560 37346
rect 34480 37280 34560 37294
rect 34640 37346 34720 37360
rect 34640 37294 34654 37346
rect 34706 37294 34720 37346
rect 34640 37280 34720 37294
rect 34800 37346 34880 37360
rect 34800 37294 34814 37346
rect 34866 37294 34880 37346
rect 34800 37280 34880 37294
rect 34960 37346 35040 37360
rect 34960 37294 34974 37346
rect 35026 37294 35040 37346
rect 34960 37280 35040 37294
rect 35120 37346 35200 37360
rect 35120 37294 35134 37346
rect 35186 37294 35200 37346
rect 35120 37280 35200 37294
rect 35280 37346 35360 37360
rect 35280 37294 35294 37346
rect 35346 37294 35360 37346
rect 35280 37280 35360 37294
rect 35440 37346 35520 37360
rect 35440 37294 35454 37346
rect 35506 37294 35520 37346
rect 35440 37280 35520 37294
rect 35600 37346 35680 37360
rect 35600 37294 35614 37346
rect 35666 37294 35680 37346
rect 35600 37280 35680 37294
rect 35760 37346 35840 37360
rect 35760 37294 35774 37346
rect 35826 37294 35840 37346
rect 35760 37280 35840 37294
rect 35920 37346 36000 37360
rect 35920 37294 35934 37346
rect 35986 37294 36000 37346
rect 35920 37280 36000 37294
rect 36080 37346 36160 37360
rect 36080 37294 36094 37346
rect 36146 37294 36160 37346
rect 36080 37280 36160 37294
rect 36240 37346 36320 37360
rect 36240 37294 36254 37346
rect 36306 37294 36320 37346
rect 36240 37280 36320 37294
rect 36400 37346 36480 37360
rect 36400 37294 36414 37346
rect 36466 37294 36480 37346
rect 36400 37280 36480 37294
rect 36560 37346 36640 37360
rect 36560 37294 36574 37346
rect 36626 37294 36640 37346
rect 36560 37280 36640 37294
rect 36720 37346 36800 37360
rect 36720 37294 36734 37346
rect 36786 37294 36800 37346
rect 36720 37280 36800 37294
rect 36880 37346 36960 37360
rect 36880 37294 36894 37346
rect 36946 37294 36960 37346
rect 36880 37280 36960 37294
rect 37040 37346 37120 37360
rect 37040 37294 37054 37346
rect 37106 37294 37120 37346
rect 37040 37280 37120 37294
rect 37200 37346 37280 37360
rect 37200 37294 37214 37346
rect 37266 37294 37280 37346
rect 37200 37280 37280 37294
rect 37360 37346 37440 37360
rect 37360 37294 37374 37346
rect 37426 37294 37440 37346
rect 37360 37280 37440 37294
rect 37520 37346 37600 37360
rect 37520 37294 37534 37346
rect 37586 37294 37600 37346
rect 37520 37280 37600 37294
rect 37680 37346 37760 37360
rect 37680 37294 37694 37346
rect 37746 37294 37760 37346
rect 37680 37280 37760 37294
rect 37840 37346 37920 37360
rect 37840 37294 37854 37346
rect 37906 37294 37920 37346
rect 37840 37280 37920 37294
rect 38000 37346 38080 37360
rect 38000 37294 38014 37346
rect 38066 37294 38080 37346
rect 38000 37280 38080 37294
rect 38160 37346 38240 37360
rect 38160 37294 38174 37346
rect 38226 37294 38240 37346
rect 38160 37280 38240 37294
rect 38320 37346 38400 37360
rect 38320 37294 38334 37346
rect 38386 37294 38400 37346
rect 38320 37280 38400 37294
rect 38480 37346 38560 37360
rect 38480 37294 38494 37346
rect 38546 37294 38560 37346
rect 38480 37280 38560 37294
rect 38640 37346 38720 37360
rect 38640 37294 38654 37346
rect 38706 37294 38720 37346
rect 38640 37280 38720 37294
rect 38800 37346 38880 37360
rect 38800 37294 38814 37346
rect 38866 37294 38880 37346
rect 38800 37280 38880 37294
rect 38960 37346 39040 37360
rect 38960 37294 38974 37346
rect 39026 37294 39040 37346
rect 38960 37280 39040 37294
rect 39120 37346 39200 37360
rect 39120 37294 39134 37346
rect 39186 37294 39200 37346
rect 39120 37280 39200 37294
rect 39280 37346 39360 37360
rect 39280 37294 39294 37346
rect 39346 37294 39360 37346
rect 39280 37280 39360 37294
rect 39440 37346 39520 37360
rect 39440 37294 39454 37346
rect 39506 37294 39520 37346
rect 39440 37280 39520 37294
rect 39600 37346 39680 37360
rect 39600 37294 39614 37346
rect 39666 37294 39680 37346
rect 39600 37280 39680 37294
rect 39760 37346 39840 37360
rect 39760 37294 39774 37346
rect 39826 37294 39840 37346
rect 39760 37280 39840 37294
rect 39920 37346 40000 37360
rect 39920 37294 39934 37346
rect 39986 37294 40000 37346
rect 39920 37280 40000 37294
rect 40080 37346 40160 37360
rect 40080 37294 40094 37346
rect 40146 37294 40160 37346
rect 40080 37280 40160 37294
rect 40240 37346 40320 37360
rect 40240 37294 40254 37346
rect 40306 37294 40320 37346
rect 40240 37280 40320 37294
rect 40400 37346 40480 37360
rect 40400 37294 40414 37346
rect 40466 37294 40480 37346
rect 40400 37280 40480 37294
rect 40560 37346 40640 37360
rect 40560 37294 40574 37346
rect 40626 37294 40640 37346
rect 40560 37280 40640 37294
rect 40720 37346 40800 37360
rect 40720 37294 40734 37346
rect 40786 37294 40800 37346
rect 40720 37280 40800 37294
rect 40880 37346 40960 37360
rect 40880 37294 40894 37346
rect 40946 37294 40960 37346
rect 40880 37280 40960 37294
rect 41040 37346 41120 37360
rect 41040 37294 41054 37346
rect 41106 37294 41120 37346
rect 41040 37280 41120 37294
rect 41200 37346 41280 37360
rect 41200 37294 41214 37346
rect 41266 37294 41280 37346
rect 41200 37280 41280 37294
rect 41360 37346 41440 37360
rect 41360 37294 41374 37346
rect 41426 37294 41440 37346
rect 41360 37280 41440 37294
rect 41520 37346 41600 37360
rect 41520 37294 41534 37346
rect 41586 37294 41600 37346
rect 41520 37280 41600 37294
rect 41680 37346 41760 37360
rect 41680 37294 41694 37346
rect 41746 37294 41760 37346
rect 41680 37280 41760 37294
rect 41840 37346 41920 37360
rect 41840 37294 41854 37346
rect 41906 37294 41920 37346
rect 41840 37280 41920 37294
rect 0 37026 80 37040
rect 0 36974 14 37026
rect 66 36974 80 37026
rect 0 36960 80 36974
rect 160 37026 240 37040
rect 160 36974 174 37026
rect 226 36974 240 37026
rect 160 36960 240 36974
rect 320 37026 400 37040
rect 320 36974 334 37026
rect 386 36974 400 37026
rect 320 36960 400 36974
rect 480 37026 560 37040
rect 480 36974 494 37026
rect 546 36974 560 37026
rect 480 36960 560 36974
rect 640 37026 720 37040
rect 640 36974 654 37026
rect 706 36974 720 37026
rect 640 36960 720 36974
rect 800 37026 880 37040
rect 800 36974 814 37026
rect 866 36974 880 37026
rect 800 36960 880 36974
rect 960 37026 1040 37040
rect 960 36974 974 37026
rect 1026 36974 1040 37026
rect 960 36960 1040 36974
rect 1120 37026 1200 37040
rect 1120 36974 1134 37026
rect 1186 36974 1200 37026
rect 1120 36960 1200 36974
rect 1280 37026 1360 37040
rect 1280 36974 1294 37026
rect 1346 36974 1360 37026
rect 1280 36960 1360 36974
rect 1440 37026 1520 37040
rect 1440 36974 1454 37026
rect 1506 36974 1520 37026
rect 1440 36960 1520 36974
rect 1600 37026 1680 37040
rect 1600 36974 1614 37026
rect 1666 36974 1680 37026
rect 1600 36960 1680 36974
rect 1760 37026 1840 37040
rect 1760 36974 1774 37026
rect 1826 36974 1840 37026
rect 1760 36960 1840 36974
rect 1920 37026 2000 37040
rect 1920 36974 1934 37026
rect 1986 36974 2000 37026
rect 1920 36960 2000 36974
rect 2080 37026 2160 37040
rect 2080 36974 2094 37026
rect 2146 36974 2160 37026
rect 2080 36960 2160 36974
rect 2240 37026 2320 37040
rect 2240 36974 2254 37026
rect 2306 36974 2320 37026
rect 2240 36960 2320 36974
rect 2400 37026 2480 37040
rect 2400 36974 2414 37026
rect 2466 36974 2480 37026
rect 2400 36960 2480 36974
rect 2560 37026 2640 37040
rect 2560 36974 2574 37026
rect 2626 36974 2640 37026
rect 2560 36960 2640 36974
rect 2720 37026 2800 37040
rect 2720 36974 2734 37026
rect 2786 36974 2800 37026
rect 2720 36960 2800 36974
rect 2880 37026 2960 37040
rect 2880 36974 2894 37026
rect 2946 36974 2960 37026
rect 2880 36960 2960 36974
rect 3040 37026 3120 37040
rect 3040 36974 3054 37026
rect 3106 36974 3120 37026
rect 3040 36960 3120 36974
rect 3200 37026 3280 37040
rect 3200 36974 3214 37026
rect 3266 36974 3280 37026
rect 3200 36960 3280 36974
rect 3360 37026 3440 37040
rect 3360 36974 3374 37026
rect 3426 36974 3440 37026
rect 3360 36960 3440 36974
rect 3520 37026 3600 37040
rect 3520 36974 3534 37026
rect 3586 36974 3600 37026
rect 3520 36960 3600 36974
rect 3680 37026 3760 37040
rect 3680 36974 3694 37026
rect 3746 36974 3760 37026
rect 3680 36960 3760 36974
rect 3840 37026 3920 37040
rect 3840 36974 3854 37026
rect 3906 36974 3920 37026
rect 3840 36960 3920 36974
rect 4000 37026 4080 37040
rect 4000 36974 4014 37026
rect 4066 36974 4080 37026
rect 4000 36960 4080 36974
rect 4160 37026 4240 37040
rect 4160 36974 4174 37026
rect 4226 36974 4240 37026
rect 4160 36960 4240 36974
rect 4320 37026 4400 37040
rect 4320 36974 4334 37026
rect 4386 36974 4400 37026
rect 4320 36960 4400 36974
rect 4480 37026 4560 37040
rect 4480 36974 4494 37026
rect 4546 36974 4560 37026
rect 4480 36960 4560 36974
rect 4640 37026 4720 37040
rect 4640 36974 4654 37026
rect 4706 36974 4720 37026
rect 4640 36960 4720 36974
rect 4800 37026 4880 37040
rect 4800 36974 4814 37026
rect 4866 36974 4880 37026
rect 4800 36960 4880 36974
rect 4960 37026 5040 37040
rect 4960 36974 4974 37026
rect 5026 36974 5040 37026
rect 4960 36960 5040 36974
rect 5120 37026 5200 37040
rect 5120 36974 5134 37026
rect 5186 36974 5200 37026
rect 5120 36960 5200 36974
rect 5280 37026 5360 37040
rect 5280 36974 5294 37026
rect 5346 36974 5360 37026
rect 5280 36960 5360 36974
rect 5440 37026 5520 37040
rect 5440 36974 5454 37026
rect 5506 36974 5520 37026
rect 5440 36960 5520 36974
rect 5600 37026 5680 37040
rect 5600 36974 5614 37026
rect 5666 36974 5680 37026
rect 5600 36960 5680 36974
rect 5760 37026 5840 37040
rect 5760 36974 5774 37026
rect 5826 36974 5840 37026
rect 5760 36960 5840 36974
rect 5920 37026 6000 37040
rect 5920 36974 5934 37026
rect 5986 36974 6000 37026
rect 5920 36960 6000 36974
rect 6080 37026 6160 37040
rect 6080 36974 6094 37026
rect 6146 36974 6160 37026
rect 6080 36960 6160 36974
rect 6240 37026 6320 37040
rect 6240 36974 6254 37026
rect 6306 36974 6320 37026
rect 6240 36960 6320 36974
rect 6400 37026 6480 37040
rect 6400 36974 6414 37026
rect 6466 36974 6480 37026
rect 6400 36960 6480 36974
rect 6560 37026 6640 37040
rect 6560 36974 6574 37026
rect 6626 36974 6640 37026
rect 6560 36960 6640 36974
rect 6720 37026 6800 37040
rect 6720 36974 6734 37026
rect 6786 36974 6800 37026
rect 6720 36960 6800 36974
rect 6880 37026 6960 37040
rect 6880 36974 6894 37026
rect 6946 36974 6960 37026
rect 6880 36960 6960 36974
rect 7040 37026 7120 37040
rect 7040 36974 7054 37026
rect 7106 36974 7120 37026
rect 7040 36960 7120 36974
rect 7200 37026 7280 37040
rect 7200 36974 7214 37026
rect 7266 36974 7280 37026
rect 7200 36960 7280 36974
rect 7360 37026 7440 37040
rect 7360 36974 7374 37026
rect 7426 36974 7440 37026
rect 7360 36960 7440 36974
rect 7520 37026 7600 37040
rect 7520 36974 7534 37026
rect 7586 36974 7600 37026
rect 7520 36960 7600 36974
rect 7680 37026 7760 37040
rect 7680 36974 7694 37026
rect 7746 36974 7760 37026
rect 7680 36960 7760 36974
rect 7840 37026 7920 37040
rect 7840 36974 7854 37026
rect 7906 36974 7920 37026
rect 7840 36960 7920 36974
rect 8000 37026 8080 37040
rect 8000 36974 8014 37026
rect 8066 36974 8080 37026
rect 8000 36960 8080 36974
rect 8160 37026 8240 37040
rect 8160 36974 8174 37026
rect 8226 36974 8240 37026
rect 8160 36960 8240 36974
rect 8320 37026 8400 37040
rect 8320 36974 8334 37026
rect 8386 36974 8400 37026
rect 8320 36960 8400 36974
rect 12480 37026 12560 37040
rect 12480 36974 12494 37026
rect 12546 36974 12560 37026
rect 12480 36960 12560 36974
rect 12640 37026 12720 37040
rect 12640 36974 12654 37026
rect 12706 36974 12720 37026
rect 12640 36960 12720 36974
rect 12800 37026 12880 37040
rect 12800 36974 12814 37026
rect 12866 36974 12880 37026
rect 12800 36960 12880 36974
rect 12960 37026 13040 37040
rect 12960 36974 12974 37026
rect 13026 36974 13040 37026
rect 12960 36960 13040 36974
rect 13120 37026 13200 37040
rect 13120 36974 13134 37026
rect 13186 36974 13200 37026
rect 13120 36960 13200 36974
rect 13280 37026 13360 37040
rect 13280 36974 13294 37026
rect 13346 36974 13360 37026
rect 13280 36960 13360 36974
rect 13440 37026 13520 37040
rect 13440 36974 13454 37026
rect 13506 36974 13520 37026
rect 13440 36960 13520 36974
rect 13600 37026 13680 37040
rect 13600 36974 13614 37026
rect 13666 36974 13680 37026
rect 13600 36960 13680 36974
rect 13760 37026 13840 37040
rect 13760 36974 13774 37026
rect 13826 36974 13840 37026
rect 13760 36960 13840 36974
rect 13920 37026 14000 37040
rect 13920 36974 13934 37026
rect 13986 36974 14000 37026
rect 13920 36960 14000 36974
rect 14080 37026 14160 37040
rect 14080 36974 14094 37026
rect 14146 36974 14160 37026
rect 14080 36960 14160 36974
rect 14240 37026 14320 37040
rect 14240 36974 14254 37026
rect 14306 36974 14320 37026
rect 14240 36960 14320 36974
rect 14400 37026 14480 37040
rect 14400 36974 14414 37026
rect 14466 36974 14480 37026
rect 14400 36960 14480 36974
rect 14560 37026 14640 37040
rect 14560 36974 14574 37026
rect 14626 36974 14640 37026
rect 14560 36960 14640 36974
rect 14720 37026 14800 37040
rect 14720 36974 14734 37026
rect 14786 36974 14800 37026
rect 14720 36960 14800 36974
rect 14880 37026 14960 37040
rect 14880 36974 14894 37026
rect 14946 36974 14960 37026
rect 14880 36960 14960 36974
rect 15040 37026 15120 37040
rect 15040 36974 15054 37026
rect 15106 36974 15120 37026
rect 15040 36960 15120 36974
rect 15200 37026 15280 37040
rect 15200 36974 15214 37026
rect 15266 36974 15280 37026
rect 15200 36960 15280 36974
rect 15360 37026 15440 37040
rect 15360 36974 15374 37026
rect 15426 36974 15440 37026
rect 15360 36960 15440 36974
rect 15520 37026 15600 37040
rect 15520 36974 15534 37026
rect 15586 36974 15600 37026
rect 15520 36960 15600 36974
rect 15680 37026 15760 37040
rect 15680 36974 15694 37026
rect 15746 36974 15760 37026
rect 15680 36960 15760 36974
rect 15840 37026 15920 37040
rect 15840 36974 15854 37026
rect 15906 36974 15920 37026
rect 15840 36960 15920 36974
rect 16000 37026 16080 37040
rect 16000 36974 16014 37026
rect 16066 36974 16080 37026
rect 16000 36960 16080 36974
rect 16160 37026 16240 37040
rect 16160 36974 16174 37026
rect 16226 36974 16240 37026
rect 16160 36960 16240 36974
rect 16320 37026 16400 37040
rect 16320 36974 16334 37026
rect 16386 36974 16400 37026
rect 16320 36960 16400 36974
rect 16480 37026 16560 37040
rect 16480 36974 16494 37026
rect 16546 36974 16560 37026
rect 16480 36960 16560 36974
rect 16640 37026 16720 37040
rect 16640 36974 16654 37026
rect 16706 36974 16720 37026
rect 16640 36960 16720 36974
rect 16800 37026 16880 37040
rect 16800 36974 16814 37026
rect 16866 36974 16880 37026
rect 16800 36960 16880 36974
rect 16960 37026 17040 37040
rect 16960 36974 16974 37026
rect 17026 36974 17040 37026
rect 16960 36960 17040 36974
rect 17120 37026 17200 37040
rect 17120 36974 17134 37026
rect 17186 36974 17200 37026
rect 17120 36960 17200 36974
rect 17280 37026 17360 37040
rect 17280 36974 17294 37026
rect 17346 36974 17360 37026
rect 17280 36960 17360 36974
rect 17440 37026 17520 37040
rect 17440 36974 17454 37026
rect 17506 36974 17520 37026
rect 17440 36960 17520 36974
rect 17600 37026 17680 37040
rect 17600 36974 17614 37026
rect 17666 36974 17680 37026
rect 17600 36960 17680 36974
rect 17760 37026 17840 37040
rect 17760 36974 17774 37026
rect 17826 36974 17840 37026
rect 17760 36960 17840 36974
rect 17920 37026 18000 37040
rect 17920 36974 17934 37026
rect 17986 36974 18000 37026
rect 17920 36960 18000 36974
rect 18080 37026 18160 37040
rect 18080 36974 18094 37026
rect 18146 36974 18160 37026
rect 18080 36960 18160 36974
rect 18240 37026 18320 37040
rect 18240 36974 18254 37026
rect 18306 36974 18320 37026
rect 18240 36960 18320 36974
rect 18400 37026 18480 37040
rect 18400 36974 18414 37026
rect 18466 36974 18480 37026
rect 18400 36960 18480 36974
rect 18560 37026 18640 37040
rect 18560 36974 18574 37026
rect 18626 36974 18640 37026
rect 18560 36960 18640 36974
rect 18720 37026 18800 37040
rect 18720 36974 18734 37026
rect 18786 36974 18800 37026
rect 18720 36960 18800 36974
rect 18880 37026 18960 37040
rect 18880 36974 18894 37026
rect 18946 36974 18960 37026
rect 18880 36960 18960 36974
rect 23120 37026 23200 37040
rect 23120 36974 23134 37026
rect 23186 36974 23200 37026
rect 23120 36960 23200 36974
rect 23280 37026 23360 37040
rect 23280 36974 23294 37026
rect 23346 36974 23360 37026
rect 23280 36960 23360 36974
rect 23440 37026 23520 37040
rect 23440 36974 23454 37026
rect 23506 36974 23520 37026
rect 23440 36960 23520 36974
rect 23600 37026 23680 37040
rect 23600 36974 23614 37026
rect 23666 36974 23680 37026
rect 23600 36960 23680 36974
rect 23760 37026 23840 37040
rect 23760 36974 23774 37026
rect 23826 36974 23840 37026
rect 23760 36960 23840 36974
rect 23920 37026 24000 37040
rect 23920 36974 23934 37026
rect 23986 36974 24000 37026
rect 23920 36960 24000 36974
rect 24080 37026 24160 37040
rect 24080 36974 24094 37026
rect 24146 36974 24160 37026
rect 24080 36960 24160 36974
rect 24240 37026 24320 37040
rect 24240 36974 24254 37026
rect 24306 36974 24320 37026
rect 24240 36960 24320 36974
rect 24400 37026 24480 37040
rect 24400 36974 24414 37026
rect 24466 36974 24480 37026
rect 24400 36960 24480 36974
rect 24560 37026 24640 37040
rect 24560 36974 24574 37026
rect 24626 36974 24640 37026
rect 24560 36960 24640 36974
rect 24720 37026 24800 37040
rect 24720 36974 24734 37026
rect 24786 36974 24800 37026
rect 24720 36960 24800 36974
rect 24880 37026 24960 37040
rect 24880 36974 24894 37026
rect 24946 36974 24960 37026
rect 24880 36960 24960 36974
rect 25040 37026 25120 37040
rect 25040 36974 25054 37026
rect 25106 36974 25120 37026
rect 25040 36960 25120 36974
rect 25200 37026 25280 37040
rect 25200 36974 25214 37026
rect 25266 36974 25280 37026
rect 25200 36960 25280 36974
rect 25360 37026 25440 37040
rect 25360 36974 25374 37026
rect 25426 36974 25440 37026
rect 25360 36960 25440 36974
rect 25520 37026 25600 37040
rect 25520 36974 25534 37026
rect 25586 36974 25600 37026
rect 25520 36960 25600 36974
rect 25680 37026 25760 37040
rect 25680 36974 25694 37026
rect 25746 36974 25760 37026
rect 25680 36960 25760 36974
rect 25840 37026 25920 37040
rect 25840 36974 25854 37026
rect 25906 36974 25920 37026
rect 25840 36960 25920 36974
rect 26000 37026 26080 37040
rect 26000 36974 26014 37026
rect 26066 36974 26080 37026
rect 26000 36960 26080 36974
rect 26160 37026 26240 37040
rect 26160 36974 26174 37026
rect 26226 36974 26240 37026
rect 26160 36960 26240 36974
rect 26320 37026 26400 37040
rect 26320 36974 26334 37026
rect 26386 36974 26400 37026
rect 26320 36960 26400 36974
rect 26480 37026 26560 37040
rect 26480 36974 26494 37026
rect 26546 36974 26560 37026
rect 26480 36960 26560 36974
rect 26640 37026 26720 37040
rect 26640 36974 26654 37026
rect 26706 36974 26720 37026
rect 26640 36960 26720 36974
rect 26800 37026 26880 37040
rect 26800 36974 26814 37026
rect 26866 36974 26880 37026
rect 26800 36960 26880 36974
rect 26960 37026 27040 37040
rect 26960 36974 26974 37026
rect 27026 36974 27040 37026
rect 26960 36960 27040 36974
rect 27120 37026 27200 37040
rect 27120 36974 27134 37026
rect 27186 36974 27200 37026
rect 27120 36960 27200 36974
rect 27280 37026 27360 37040
rect 27280 36974 27294 37026
rect 27346 36974 27360 37026
rect 27280 36960 27360 36974
rect 27440 37026 27520 37040
rect 27440 36974 27454 37026
rect 27506 36974 27520 37026
rect 27440 36960 27520 36974
rect 27600 37026 27680 37040
rect 27600 36974 27614 37026
rect 27666 36974 27680 37026
rect 27600 36960 27680 36974
rect 27760 37026 27840 37040
rect 27760 36974 27774 37026
rect 27826 36974 27840 37026
rect 27760 36960 27840 36974
rect 27920 37026 28000 37040
rect 27920 36974 27934 37026
rect 27986 36974 28000 37026
rect 27920 36960 28000 36974
rect 28080 37026 28160 37040
rect 28080 36974 28094 37026
rect 28146 36974 28160 37026
rect 28080 36960 28160 36974
rect 28240 37026 28320 37040
rect 28240 36974 28254 37026
rect 28306 36974 28320 37026
rect 28240 36960 28320 36974
rect 28400 37026 28480 37040
rect 28400 36974 28414 37026
rect 28466 36974 28480 37026
rect 28400 36960 28480 36974
rect 28560 37026 28640 37040
rect 28560 36974 28574 37026
rect 28626 36974 28640 37026
rect 28560 36960 28640 36974
rect 28720 37026 28800 37040
rect 28720 36974 28734 37026
rect 28786 36974 28800 37026
rect 28720 36960 28800 36974
rect 28880 37026 28960 37040
rect 28880 36974 28894 37026
rect 28946 36974 28960 37026
rect 28880 36960 28960 36974
rect 29040 37026 29120 37040
rect 29040 36974 29054 37026
rect 29106 36974 29120 37026
rect 29040 36960 29120 36974
rect 29200 37026 29280 37040
rect 29200 36974 29214 37026
rect 29266 36974 29280 37026
rect 29200 36960 29280 36974
rect 29360 37026 29440 37040
rect 29360 36974 29374 37026
rect 29426 36974 29440 37026
rect 29360 36960 29440 36974
rect 33520 37026 33600 37040
rect 33520 36974 33534 37026
rect 33586 36974 33600 37026
rect 33520 36960 33600 36974
rect 33680 37026 33760 37040
rect 33680 36974 33694 37026
rect 33746 36974 33760 37026
rect 33680 36960 33760 36974
rect 33840 37026 33920 37040
rect 33840 36974 33854 37026
rect 33906 36974 33920 37026
rect 33840 36960 33920 36974
rect 34000 37026 34080 37040
rect 34000 36974 34014 37026
rect 34066 36974 34080 37026
rect 34000 36960 34080 36974
rect 34160 37026 34240 37040
rect 34160 36974 34174 37026
rect 34226 36974 34240 37026
rect 34160 36960 34240 36974
rect 34320 37026 34400 37040
rect 34320 36974 34334 37026
rect 34386 36974 34400 37026
rect 34320 36960 34400 36974
rect 34480 37026 34560 37040
rect 34480 36974 34494 37026
rect 34546 36974 34560 37026
rect 34480 36960 34560 36974
rect 34640 37026 34720 37040
rect 34640 36974 34654 37026
rect 34706 36974 34720 37026
rect 34640 36960 34720 36974
rect 34800 37026 34880 37040
rect 34800 36974 34814 37026
rect 34866 36974 34880 37026
rect 34800 36960 34880 36974
rect 34960 37026 35040 37040
rect 34960 36974 34974 37026
rect 35026 36974 35040 37026
rect 34960 36960 35040 36974
rect 35120 37026 35200 37040
rect 35120 36974 35134 37026
rect 35186 36974 35200 37026
rect 35120 36960 35200 36974
rect 35280 37026 35360 37040
rect 35280 36974 35294 37026
rect 35346 36974 35360 37026
rect 35280 36960 35360 36974
rect 35440 37026 35520 37040
rect 35440 36974 35454 37026
rect 35506 36974 35520 37026
rect 35440 36960 35520 36974
rect 35600 37026 35680 37040
rect 35600 36974 35614 37026
rect 35666 36974 35680 37026
rect 35600 36960 35680 36974
rect 35760 37026 35840 37040
rect 35760 36974 35774 37026
rect 35826 36974 35840 37026
rect 35760 36960 35840 36974
rect 35920 37026 36000 37040
rect 35920 36974 35934 37026
rect 35986 36974 36000 37026
rect 35920 36960 36000 36974
rect 36080 37026 36160 37040
rect 36080 36974 36094 37026
rect 36146 36974 36160 37026
rect 36080 36960 36160 36974
rect 36240 37026 36320 37040
rect 36240 36974 36254 37026
rect 36306 36974 36320 37026
rect 36240 36960 36320 36974
rect 36400 37026 36480 37040
rect 36400 36974 36414 37026
rect 36466 36974 36480 37026
rect 36400 36960 36480 36974
rect 36560 37026 36640 37040
rect 36560 36974 36574 37026
rect 36626 36974 36640 37026
rect 36560 36960 36640 36974
rect 36720 37026 36800 37040
rect 36720 36974 36734 37026
rect 36786 36974 36800 37026
rect 36720 36960 36800 36974
rect 36880 37026 36960 37040
rect 36880 36974 36894 37026
rect 36946 36974 36960 37026
rect 36880 36960 36960 36974
rect 37040 37026 37120 37040
rect 37040 36974 37054 37026
rect 37106 36974 37120 37026
rect 37040 36960 37120 36974
rect 37200 37026 37280 37040
rect 37200 36974 37214 37026
rect 37266 36974 37280 37026
rect 37200 36960 37280 36974
rect 37360 37026 37440 37040
rect 37360 36974 37374 37026
rect 37426 36974 37440 37026
rect 37360 36960 37440 36974
rect 37520 37026 37600 37040
rect 37520 36974 37534 37026
rect 37586 36974 37600 37026
rect 37520 36960 37600 36974
rect 37680 37026 37760 37040
rect 37680 36974 37694 37026
rect 37746 36974 37760 37026
rect 37680 36960 37760 36974
rect 37840 37026 37920 37040
rect 37840 36974 37854 37026
rect 37906 36974 37920 37026
rect 37840 36960 37920 36974
rect 38000 37026 38080 37040
rect 38000 36974 38014 37026
rect 38066 36974 38080 37026
rect 38000 36960 38080 36974
rect 38160 37026 38240 37040
rect 38160 36974 38174 37026
rect 38226 36974 38240 37026
rect 38160 36960 38240 36974
rect 38320 37026 38400 37040
rect 38320 36974 38334 37026
rect 38386 36974 38400 37026
rect 38320 36960 38400 36974
rect 38480 37026 38560 37040
rect 38480 36974 38494 37026
rect 38546 36974 38560 37026
rect 38480 36960 38560 36974
rect 38640 37026 38720 37040
rect 38640 36974 38654 37026
rect 38706 36974 38720 37026
rect 38640 36960 38720 36974
rect 38800 37026 38880 37040
rect 38800 36974 38814 37026
rect 38866 36974 38880 37026
rect 38800 36960 38880 36974
rect 38960 37026 39040 37040
rect 38960 36974 38974 37026
rect 39026 36974 39040 37026
rect 38960 36960 39040 36974
rect 39120 37026 39200 37040
rect 39120 36974 39134 37026
rect 39186 36974 39200 37026
rect 39120 36960 39200 36974
rect 39280 37026 39360 37040
rect 39280 36974 39294 37026
rect 39346 36974 39360 37026
rect 39280 36960 39360 36974
rect 39440 37026 39520 37040
rect 39440 36974 39454 37026
rect 39506 36974 39520 37026
rect 39440 36960 39520 36974
rect 39600 37026 39680 37040
rect 39600 36974 39614 37026
rect 39666 36974 39680 37026
rect 39600 36960 39680 36974
rect 39760 37026 39840 37040
rect 39760 36974 39774 37026
rect 39826 36974 39840 37026
rect 39760 36960 39840 36974
rect 39920 37026 40000 37040
rect 39920 36974 39934 37026
rect 39986 36974 40000 37026
rect 39920 36960 40000 36974
rect 40080 37026 40160 37040
rect 40080 36974 40094 37026
rect 40146 36974 40160 37026
rect 40080 36960 40160 36974
rect 40240 37026 40320 37040
rect 40240 36974 40254 37026
rect 40306 36974 40320 37026
rect 40240 36960 40320 36974
rect 40400 37026 40480 37040
rect 40400 36974 40414 37026
rect 40466 36974 40480 37026
rect 40400 36960 40480 36974
rect 40560 37026 40640 37040
rect 40560 36974 40574 37026
rect 40626 36974 40640 37026
rect 40560 36960 40640 36974
rect 40720 37026 40800 37040
rect 40720 36974 40734 37026
rect 40786 36974 40800 37026
rect 40720 36960 40800 36974
rect 40880 37026 40960 37040
rect 40880 36974 40894 37026
rect 40946 36974 40960 37026
rect 40880 36960 40960 36974
rect 41040 37026 41120 37040
rect 41040 36974 41054 37026
rect 41106 36974 41120 37026
rect 41040 36960 41120 36974
rect 41200 37026 41280 37040
rect 41200 36974 41214 37026
rect 41266 36974 41280 37026
rect 41200 36960 41280 36974
rect 41360 37026 41440 37040
rect 41360 36974 41374 37026
rect 41426 36974 41440 37026
rect 41360 36960 41440 36974
rect 41520 37026 41600 37040
rect 41520 36974 41534 37026
rect 41586 36974 41600 37026
rect 41520 36960 41600 36974
rect 41680 37026 41760 37040
rect 41680 36974 41694 37026
rect 41746 36974 41760 37026
rect 41680 36960 41760 36974
rect 41840 37026 41920 37040
rect 41840 36974 41854 37026
rect 41906 36974 41920 37026
rect 41840 36960 41920 36974
rect 0 36866 80 36880
rect 0 36814 14 36866
rect 66 36814 80 36866
rect 0 36800 80 36814
rect 160 36866 240 36880
rect 160 36814 174 36866
rect 226 36814 240 36866
rect 160 36800 240 36814
rect 320 36866 400 36880
rect 320 36814 334 36866
rect 386 36814 400 36866
rect 320 36800 400 36814
rect 480 36866 560 36880
rect 480 36814 494 36866
rect 546 36814 560 36866
rect 480 36800 560 36814
rect 640 36866 720 36880
rect 640 36814 654 36866
rect 706 36814 720 36866
rect 640 36800 720 36814
rect 800 36866 880 36880
rect 800 36814 814 36866
rect 866 36814 880 36866
rect 800 36800 880 36814
rect 960 36866 1040 36880
rect 960 36814 974 36866
rect 1026 36814 1040 36866
rect 960 36800 1040 36814
rect 1120 36866 1200 36880
rect 1120 36814 1134 36866
rect 1186 36814 1200 36866
rect 1120 36800 1200 36814
rect 1280 36866 1360 36880
rect 1280 36814 1294 36866
rect 1346 36814 1360 36866
rect 1280 36800 1360 36814
rect 1440 36866 1520 36880
rect 1440 36814 1454 36866
rect 1506 36814 1520 36866
rect 1440 36800 1520 36814
rect 1600 36866 1680 36880
rect 1600 36814 1614 36866
rect 1666 36814 1680 36866
rect 1600 36800 1680 36814
rect 1760 36866 1840 36880
rect 1760 36814 1774 36866
rect 1826 36814 1840 36866
rect 1760 36800 1840 36814
rect 1920 36866 2000 36880
rect 1920 36814 1934 36866
rect 1986 36814 2000 36866
rect 1920 36800 2000 36814
rect 2080 36866 2160 36880
rect 2080 36814 2094 36866
rect 2146 36814 2160 36866
rect 2080 36800 2160 36814
rect 2240 36866 2320 36880
rect 2240 36814 2254 36866
rect 2306 36814 2320 36866
rect 2240 36800 2320 36814
rect 2400 36866 2480 36880
rect 2400 36814 2414 36866
rect 2466 36814 2480 36866
rect 2400 36800 2480 36814
rect 2560 36866 2640 36880
rect 2560 36814 2574 36866
rect 2626 36814 2640 36866
rect 2560 36800 2640 36814
rect 2720 36866 2800 36880
rect 2720 36814 2734 36866
rect 2786 36814 2800 36866
rect 2720 36800 2800 36814
rect 2880 36866 2960 36880
rect 2880 36814 2894 36866
rect 2946 36814 2960 36866
rect 2880 36800 2960 36814
rect 3040 36866 3120 36880
rect 3040 36814 3054 36866
rect 3106 36814 3120 36866
rect 3040 36800 3120 36814
rect 3200 36866 3280 36880
rect 3200 36814 3214 36866
rect 3266 36814 3280 36866
rect 3200 36800 3280 36814
rect 3360 36866 3440 36880
rect 3360 36814 3374 36866
rect 3426 36814 3440 36866
rect 3360 36800 3440 36814
rect 3520 36866 3600 36880
rect 3520 36814 3534 36866
rect 3586 36814 3600 36866
rect 3520 36800 3600 36814
rect 3680 36866 3760 36880
rect 3680 36814 3694 36866
rect 3746 36814 3760 36866
rect 3680 36800 3760 36814
rect 3840 36866 3920 36880
rect 3840 36814 3854 36866
rect 3906 36814 3920 36866
rect 3840 36800 3920 36814
rect 4000 36866 4080 36880
rect 4000 36814 4014 36866
rect 4066 36814 4080 36866
rect 4000 36800 4080 36814
rect 4160 36866 4240 36880
rect 4160 36814 4174 36866
rect 4226 36814 4240 36866
rect 4160 36800 4240 36814
rect 4320 36866 4400 36880
rect 4320 36814 4334 36866
rect 4386 36814 4400 36866
rect 4320 36800 4400 36814
rect 4480 36866 4560 36880
rect 4480 36814 4494 36866
rect 4546 36814 4560 36866
rect 4480 36800 4560 36814
rect 4640 36866 4720 36880
rect 4640 36814 4654 36866
rect 4706 36814 4720 36866
rect 4640 36800 4720 36814
rect 4800 36866 4880 36880
rect 4800 36814 4814 36866
rect 4866 36814 4880 36866
rect 4800 36800 4880 36814
rect 4960 36866 5040 36880
rect 4960 36814 4974 36866
rect 5026 36814 5040 36866
rect 4960 36800 5040 36814
rect 5120 36866 5200 36880
rect 5120 36814 5134 36866
rect 5186 36814 5200 36866
rect 5120 36800 5200 36814
rect 5280 36866 5360 36880
rect 5280 36814 5294 36866
rect 5346 36814 5360 36866
rect 5280 36800 5360 36814
rect 5440 36866 5520 36880
rect 5440 36814 5454 36866
rect 5506 36814 5520 36866
rect 5440 36800 5520 36814
rect 5600 36866 5680 36880
rect 5600 36814 5614 36866
rect 5666 36814 5680 36866
rect 5600 36800 5680 36814
rect 5760 36866 5840 36880
rect 5760 36814 5774 36866
rect 5826 36814 5840 36866
rect 5760 36800 5840 36814
rect 5920 36866 6000 36880
rect 5920 36814 5934 36866
rect 5986 36814 6000 36866
rect 5920 36800 6000 36814
rect 6080 36866 6160 36880
rect 6080 36814 6094 36866
rect 6146 36814 6160 36866
rect 6080 36800 6160 36814
rect 6240 36866 6320 36880
rect 6240 36814 6254 36866
rect 6306 36814 6320 36866
rect 6240 36800 6320 36814
rect 6400 36866 6480 36880
rect 6400 36814 6414 36866
rect 6466 36814 6480 36866
rect 6400 36800 6480 36814
rect 6560 36866 6640 36880
rect 6560 36814 6574 36866
rect 6626 36814 6640 36866
rect 6560 36800 6640 36814
rect 6720 36866 6800 36880
rect 6720 36814 6734 36866
rect 6786 36814 6800 36866
rect 6720 36800 6800 36814
rect 6880 36866 6960 36880
rect 6880 36814 6894 36866
rect 6946 36814 6960 36866
rect 6880 36800 6960 36814
rect 7040 36866 7120 36880
rect 7040 36814 7054 36866
rect 7106 36814 7120 36866
rect 7040 36800 7120 36814
rect 7200 36866 7280 36880
rect 7200 36814 7214 36866
rect 7266 36814 7280 36866
rect 7200 36800 7280 36814
rect 7360 36866 7440 36880
rect 7360 36814 7374 36866
rect 7426 36814 7440 36866
rect 7360 36800 7440 36814
rect 7520 36866 7600 36880
rect 7520 36814 7534 36866
rect 7586 36814 7600 36866
rect 7520 36800 7600 36814
rect 7680 36866 7760 36880
rect 7680 36814 7694 36866
rect 7746 36814 7760 36866
rect 7680 36800 7760 36814
rect 7840 36866 7920 36880
rect 7840 36814 7854 36866
rect 7906 36814 7920 36866
rect 7840 36800 7920 36814
rect 8000 36866 8080 36880
rect 8000 36814 8014 36866
rect 8066 36814 8080 36866
rect 8000 36800 8080 36814
rect 8160 36866 8240 36880
rect 8160 36814 8174 36866
rect 8226 36814 8240 36866
rect 8160 36800 8240 36814
rect 8320 36866 8400 36880
rect 8320 36814 8334 36866
rect 8386 36814 8400 36866
rect 8320 36800 8400 36814
rect 12480 36866 12560 36880
rect 12480 36814 12494 36866
rect 12546 36814 12560 36866
rect 12480 36800 12560 36814
rect 12640 36866 12720 36880
rect 12640 36814 12654 36866
rect 12706 36814 12720 36866
rect 12640 36800 12720 36814
rect 12800 36866 12880 36880
rect 12800 36814 12814 36866
rect 12866 36814 12880 36866
rect 12800 36800 12880 36814
rect 12960 36866 13040 36880
rect 12960 36814 12974 36866
rect 13026 36814 13040 36866
rect 12960 36800 13040 36814
rect 13120 36866 13200 36880
rect 13120 36814 13134 36866
rect 13186 36814 13200 36866
rect 13120 36800 13200 36814
rect 13280 36866 13360 36880
rect 13280 36814 13294 36866
rect 13346 36814 13360 36866
rect 13280 36800 13360 36814
rect 13440 36866 13520 36880
rect 13440 36814 13454 36866
rect 13506 36814 13520 36866
rect 13440 36800 13520 36814
rect 13600 36866 13680 36880
rect 13600 36814 13614 36866
rect 13666 36814 13680 36866
rect 13600 36800 13680 36814
rect 13760 36866 13840 36880
rect 13760 36814 13774 36866
rect 13826 36814 13840 36866
rect 13760 36800 13840 36814
rect 13920 36866 14000 36880
rect 13920 36814 13934 36866
rect 13986 36814 14000 36866
rect 13920 36800 14000 36814
rect 14080 36866 14160 36880
rect 14080 36814 14094 36866
rect 14146 36814 14160 36866
rect 14080 36800 14160 36814
rect 14240 36866 14320 36880
rect 14240 36814 14254 36866
rect 14306 36814 14320 36866
rect 14240 36800 14320 36814
rect 14400 36866 14480 36880
rect 14400 36814 14414 36866
rect 14466 36814 14480 36866
rect 14400 36800 14480 36814
rect 14560 36866 14640 36880
rect 14560 36814 14574 36866
rect 14626 36814 14640 36866
rect 14560 36800 14640 36814
rect 14720 36866 14800 36880
rect 14720 36814 14734 36866
rect 14786 36814 14800 36866
rect 14720 36800 14800 36814
rect 14880 36866 14960 36880
rect 14880 36814 14894 36866
rect 14946 36814 14960 36866
rect 14880 36800 14960 36814
rect 15040 36866 15120 36880
rect 15040 36814 15054 36866
rect 15106 36814 15120 36866
rect 15040 36800 15120 36814
rect 15200 36866 15280 36880
rect 15200 36814 15214 36866
rect 15266 36814 15280 36866
rect 15200 36800 15280 36814
rect 15360 36866 15440 36880
rect 15360 36814 15374 36866
rect 15426 36814 15440 36866
rect 15360 36800 15440 36814
rect 15520 36866 15600 36880
rect 15520 36814 15534 36866
rect 15586 36814 15600 36866
rect 15520 36800 15600 36814
rect 15680 36866 15760 36880
rect 15680 36814 15694 36866
rect 15746 36814 15760 36866
rect 15680 36800 15760 36814
rect 15840 36866 15920 36880
rect 15840 36814 15854 36866
rect 15906 36814 15920 36866
rect 15840 36800 15920 36814
rect 16000 36866 16080 36880
rect 16000 36814 16014 36866
rect 16066 36814 16080 36866
rect 16000 36800 16080 36814
rect 16160 36866 16240 36880
rect 16160 36814 16174 36866
rect 16226 36814 16240 36866
rect 16160 36800 16240 36814
rect 16320 36866 16400 36880
rect 16320 36814 16334 36866
rect 16386 36814 16400 36866
rect 16320 36800 16400 36814
rect 16480 36866 16560 36880
rect 16480 36814 16494 36866
rect 16546 36814 16560 36866
rect 16480 36800 16560 36814
rect 16640 36866 16720 36880
rect 16640 36814 16654 36866
rect 16706 36814 16720 36866
rect 16640 36800 16720 36814
rect 16800 36866 16880 36880
rect 16800 36814 16814 36866
rect 16866 36814 16880 36866
rect 16800 36800 16880 36814
rect 16960 36866 17040 36880
rect 16960 36814 16974 36866
rect 17026 36814 17040 36866
rect 16960 36800 17040 36814
rect 17120 36866 17200 36880
rect 17120 36814 17134 36866
rect 17186 36814 17200 36866
rect 17120 36800 17200 36814
rect 17280 36866 17360 36880
rect 17280 36814 17294 36866
rect 17346 36814 17360 36866
rect 17280 36800 17360 36814
rect 17440 36866 17520 36880
rect 17440 36814 17454 36866
rect 17506 36814 17520 36866
rect 17440 36800 17520 36814
rect 17600 36866 17680 36880
rect 17600 36814 17614 36866
rect 17666 36814 17680 36866
rect 17600 36800 17680 36814
rect 17760 36866 17840 36880
rect 17760 36814 17774 36866
rect 17826 36814 17840 36866
rect 17760 36800 17840 36814
rect 17920 36866 18000 36880
rect 17920 36814 17934 36866
rect 17986 36814 18000 36866
rect 17920 36800 18000 36814
rect 18080 36866 18160 36880
rect 18080 36814 18094 36866
rect 18146 36814 18160 36866
rect 18080 36800 18160 36814
rect 18240 36866 18320 36880
rect 18240 36814 18254 36866
rect 18306 36814 18320 36866
rect 18240 36800 18320 36814
rect 18400 36866 18480 36880
rect 18400 36814 18414 36866
rect 18466 36814 18480 36866
rect 18400 36800 18480 36814
rect 18560 36866 18640 36880
rect 18560 36814 18574 36866
rect 18626 36814 18640 36866
rect 18560 36800 18640 36814
rect 18720 36866 18800 36880
rect 18720 36814 18734 36866
rect 18786 36814 18800 36866
rect 18720 36800 18800 36814
rect 18880 36866 18960 36880
rect 18880 36814 18894 36866
rect 18946 36814 18960 36866
rect 18880 36800 18960 36814
rect 23120 36866 23200 36880
rect 23120 36814 23134 36866
rect 23186 36814 23200 36866
rect 23120 36800 23200 36814
rect 23280 36866 23360 36880
rect 23280 36814 23294 36866
rect 23346 36814 23360 36866
rect 23280 36800 23360 36814
rect 23440 36866 23520 36880
rect 23440 36814 23454 36866
rect 23506 36814 23520 36866
rect 23440 36800 23520 36814
rect 23600 36866 23680 36880
rect 23600 36814 23614 36866
rect 23666 36814 23680 36866
rect 23600 36800 23680 36814
rect 23760 36866 23840 36880
rect 23760 36814 23774 36866
rect 23826 36814 23840 36866
rect 23760 36800 23840 36814
rect 23920 36866 24000 36880
rect 23920 36814 23934 36866
rect 23986 36814 24000 36866
rect 23920 36800 24000 36814
rect 24080 36866 24160 36880
rect 24080 36814 24094 36866
rect 24146 36814 24160 36866
rect 24080 36800 24160 36814
rect 24240 36866 24320 36880
rect 24240 36814 24254 36866
rect 24306 36814 24320 36866
rect 24240 36800 24320 36814
rect 24400 36866 24480 36880
rect 24400 36814 24414 36866
rect 24466 36814 24480 36866
rect 24400 36800 24480 36814
rect 24560 36866 24640 36880
rect 24560 36814 24574 36866
rect 24626 36814 24640 36866
rect 24560 36800 24640 36814
rect 24720 36866 24800 36880
rect 24720 36814 24734 36866
rect 24786 36814 24800 36866
rect 24720 36800 24800 36814
rect 24880 36866 24960 36880
rect 24880 36814 24894 36866
rect 24946 36814 24960 36866
rect 24880 36800 24960 36814
rect 25040 36866 25120 36880
rect 25040 36814 25054 36866
rect 25106 36814 25120 36866
rect 25040 36800 25120 36814
rect 25200 36866 25280 36880
rect 25200 36814 25214 36866
rect 25266 36814 25280 36866
rect 25200 36800 25280 36814
rect 25360 36866 25440 36880
rect 25360 36814 25374 36866
rect 25426 36814 25440 36866
rect 25360 36800 25440 36814
rect 25520 36866 25600 36880
rect 25520 36814 25534 36866
rect 25586 36814 25600 36866
rect 25520 36800 25600 36814
rect 25680 36866 25760 36880
rect 25680 36814 25694 36866
rect 25746 36814 25760 36866
rect 25680 36800 25760 36814
rect 25840 36866 25920 36880
rect 25840 36814 25854 36866
rect 25906 36814 25920 36866
rect 25840 36800 25920 36814
rect 26000 36866 26080 36880
rect 26000 36814 26014 36866
rect 26066 36814 26080 36866
rect 26000 36800 26080 36814
rect 26160 36866 26240 36880
rect 26160 36814 26174 36866
rect 26226 36814 26240 36866
rect 26160 36800 26240 36814
rect 26320 36866 26400 36880
rect 26320 36814 26334 36866
rect 26386 36814 26400 36866
rect 26320 36800 26400 36814
rect 26480 36866 26560 36880
rect 26480 36814 26494 36866
rect 26546 36814 26560 36866
rect 26480 36800 26560 36814
rect 26640 36866 26720 36880
rect 26640 36814 26654 36866
rect 26706 36814 26720 36866
rect 26640 36800 26720 36814
rect 26800 36866 26880 36880
rect 26800 36814 26814 36866
rect 26866 36814 26880 36866
rect 26800 36800 26880 36814
rect 26960 36866 27040 36880
rect 26960 36814 26974 36866
rect 27026 36814 27040 36866
rect 26960 36800 27040 36814
rect 27120 36866 27200 36880
rect 27120 36814 27134 36866
rect 27186 36814 27200 36866
rect 27120 36800 27200 36814
rect 27280 36866 27360 36880
rect 27280 36814 27294 36866
rect 27346 36814 27360 36866
rect 27280 36800 27360 36814
rect 27440 36866 27520 36880
rect 27440 36814 27454 36866
rect 27506 36814 27520 36866
rect 27440 36800 27520 36814
rect 27600 36866 27680 36880
rect 27600 36814 27614 36866
rect 27666 36814 27680 36866
rect 27600 36800 27680 36814
rect 27760 36866 27840 36880
rect 27760 36814 27774 36866
rect 27826 36814 27840 36866
rect 27760 36800 27840 36814
rect 27920 36866 28000 36880
rect 27920 36814 27934 36866
rect 27986 36814 28000 36866
rect 27920 36800 28000 36814
rect 28080 36866 28160 36880
rect 28080 36814 28094 36866
rect 28146 36814 28160 36866
rect 28080 36800 28160 36814
rect 28240 36866 28320 36880
rect 28240 36814 28254 36866
rect 28306 36814 28320 36866
rect 28240 36800 28320 36814
rect 28400 36866 28480 36880
rect 28400 36814 28414 36866
rect 28466 36814 28480 36866
rect 28400 36800 28480 36814
rect 28560 36866 28640 36880
rect 28560 36814 28574 36866
rect 28626 36814 28640 36866
rect 28560 36800 28640 36814
rect 28720 36866 28800 36880
rect 28720 36814 28734 36866
rect 28786 36814 28800 36866
rect 28720 36800 28800 36814
rect 28880 36866 28960 36880
rect 28880 36814 28894 36866
rect 28946 36814 28960 36866
rect 28880 36800 28960 36814
rect 29040 36866 29120 36880
rect 29040 36814 29054 36866
rect 29106 36814 29120 36866
rect 29040 36800 29120 36814
rect 29200 36866 29280 36880
rect 29200 36814 29214 36866
rect 29266 36814 29280 36866
rect 29200 36800 29280 36814
rect 29360 36866 29440 36880
rect 29360 36814 29374 36866
rect 29426 36814 29440 36866
rect 29360 36800 29440 36814
rect 33520 36866 33600 36880
rect 33520 36814 33534 36866
rect 33586 36814 33600 36866
rect 33520 36800 33600 36814
rect 33680 36866 33760 36880
rect 33680 36814 33694 36866
rect 33746 36814 33760 36866
rect 33680 36800 33760 36814
rect 33840 36866 33920 36880
rect 33840 36814 33854 36866
rect 33906 36814 33920 36866
rect 33840 36800 33920 36814
rect 34000 36866 34080 36880
rect 34000 36814 34014 36866
rect 34066 36814 34080 36866
rect 34000 36800 34080 36814
rect 34160 36866 34240 36880
rect 34160 36814 34174 36866
rect 34226 36814 34240 36866
rect 34160 36800 34240 36814
rect 34320 36866 34400 36880
rect 34320 36814 34334 36866
rect 34386 36814 34400 36866
rect 34320 36800 34400 36814
rect 34480 36866 34560 36880
rect 34480 36814 34494 36866
rect 34546 36814 34560 36866
rect 34480 36800 34560 36814
rect 34640 36866 34720 36880
rect 34640 36814 34654 36866
rect 34706 36814 34720 36866
rect 34640 36800 34720 36814
rect 34800 36866 34880 36880
rect 34800 36814 34814 36866
rect 34866 36814 34880 36866
rect 34800 36800 34880 36814
rect 34960 36866 35040 36880
rect 34960 36814 34974 36866
rect 35026 36814 35040 36866
rect 34960 36800 35040 36814
rect 35120 36866 35200 36880
rect 35120 36814 35134 36866
rect 35186 36814 35200 36866
rect 35120 36800 35200 36814
rect 35280 36866 35360 36880
rect 35280 36814 35294 36866
rect 35346 36814 35360 36866
rect 35280 36800 35360 36814
rect 35440 36866 35520 36880
rect 35440 36814 35454 36866
rect 35506 36814 35520 36866
rect 35440 36800 35520 36814
rect 35600 36866 35680 36880
rect 35600 36814 35614 36866
rect 35666 36814 35680 36866
rect 35600 36800 35680 36814
rect 35760 36866 35840 36880
rect 35760 36814 35774 36866
rect 35826 36814 35840 36866
rect 35760 36800 35840 36814
rect 35920 36866 36000 36880
rect 35920 36814 35934 36866
rect 35986 36814 36000 36866
rect 35920 36800 36000 36814
rect 36080 36866 36160 36880
rect 36080 36814 36094 36866
rect 36146 36814 36160 36866
rect 36080 36800 36160 36814
rect 36240 36866 36320 36880
rect 36240 36814 36254 36866
rect 36306 36814 36320 36866
rect 36240 36800 36320 36814
rect 36400 36866 36480 36880
rect 36400 36814 36414 36866
rect 36466 36814 36480 36866
rect 36400 36800 36480 36814
rect 36560 36866 36640 36880
rect 36560 36814 36574 36866
rect 36626 36814 36640 36866
rect 36560 36800 36640 36814
rect 36720 36866 36800 36880
rect 36720 36814 36734 36866
rect 36786 36814 36800 36866
rect 36720 36800 36800 36814
rect 36880 36866 36960 36880
rect 36880 36814 36894 36866
rect 36946 36814 36960 36866
rect 36880 36800 36960 36814
rect 37040 36866 37120 36880
rect 37040 36814 37054 36866
rect 37106 36814 37120 36866
rect 37040 36800 37120 36814
rect 37200 36866 37280 36880
rect 37200 36814 37214 36866
rect 37266 36814 37280 36866
rect 37200 36800 37280 36814
rect 37360 36866 37440 36880
rect 37360 36814 37374 36866
rect 37426 36814 37440 36866
rect 37360 36800 37440 36814
rect 37520 36866 37600 36880
rect 37520 36814 37534 36866
rect 37586 36814 37600 36866
rect 37520 36800 37600 36814
rect 37680 36866 37760 36880
rect 37680 36814 37694 36866
rect 37746 36814 37760 36866
rect 37680 36800 37760 36814
rect 37840 36866 37920 36880
rect 37840 36814 37854 36866
rect 37906 36814 37920 36866
rect 37840 36800 37920 36814
rect 38000 36866 38080 36880
rect 38000 36814 38014 36866
rect 38066 36814 38080 36866
rect 38000 36800 38080 36814
rect 38160 36866 38240 36880
rect 38160 36814 38174 36866
rect 38226 36814 38240 36866
rect 38160 36800 38240 36814
rect 38320 36866 38400 36880
rect 38320 36814 38334 36866
rect 38386 36814 38400 36866
rect 38320 36800 38400 36814
rect 38480 36866 38560 36880
rect 38480 36814 38494 36866
rect 38546 36814 38560 36866
rect 38480 36800 38560 36814
rect 38640 36866 38720 36880
rect 38640 36814 38654 36866
rect 38706 36814 38720 36866
rect 38640 36800 38720 36814
rect 38800 36866 38880 36880
rect 38800 36814 38814 36866
rect 38866 36814 38880 36866
rect 38800 36800 38880 36814
rect 38960 36866 39040 36880
rect 38960 36814 38974 36866
rect 39026 36814 39040 36866
rect 38960 36800 39040 36814
rect 39120 36866 39200 36880
rect 39120 36814 39134 36866
rect 39186 36814 39200 36866
rect 39120 36800 39200 36814
rect 39280 36866 39360 36880
rect 39280 36814 39294 36866
rect 39346 36814 39360 36866
rect 39280 36800 39360 36814
rect 39440 36866 39520 36880
rect 39440 36814 39454 36866
rect 39506 36814 39520 36866
rect 39440 36800 39520 36814
rect 39600 36866 39680 36880
rect 39600 36814 39614 36866
rect 39666 36814 39680 36866
rect 39600 36800 39680 36814
rect 39760 36866 39840 36880
rect 39760 36814 39774 36866
rect 39826 36814 39840 36866
rect 39760 36800 39840 36814
rect 39920 36866 40000 36880
rect 39920 36814 39934 36866
rect 39986 36814 40000 36866
rect 39920 36800 40000 36814
rect 40080 36866 40160 36880
rect 40080 36814 40094 36866
rect 40146 36814 40160 36866
rect 40080 36800 40160 36814
rect 40240 36866 40320 36880
rect 40240 36814 40254 36866
rect 40306 36814 40320 36866
rect 40240 36800 40320 36814
rect 40400 36866 40480 36880
rect 40400 36814 40414 36866
rect 40466 36814 40480 36866
rect 40400 36800 40480 36814
rect 40560 36866 40640 36880
rect 40560 36814 40574 36866
rect 40626 36814 40640 36866
rect 40560 36800 40640 36814
rect 40720 36866 40800 36880
rect 40720 36814 40734 36866
rect 40786 36814 40800 36866
rect 40720 36800 40800 36814
rect 40880 36866 40960 36880
rect 40880 36814 40894 36866
rect 40946 36814 40960 36866
rect 40880 36800 40960 36814
rect 41040 36866 41120 36880
rect 41040 36814 41054 36866
rect 41106 36814 41120 36866
rect 41040 36800 41120 36814
rect 41200 36866 41280 36880
rect 41200 36814 41214 36866
rect 41266 36814 41280 36866
rect 41200 36800 41280 36814
rect 41360 36866 41440 36880
rect 41360 36814 41374 36866
rect 41426 36814 41440 36866
rect 41360 36800 41440 36814
rect 41520 36866 41600 36880
rect 41520 36814 41534 36866
rect 41586 36814 41600 36866
rect 41520 36800 41600 36814
rect 41680 36866 41760 36880
rect 41680 36814 41694 36866
rect 41746 36814 41760 36866
rect 41680 36800 41760 36814
rect 41840 36866 41920 36880
rect 41840 36814 41854 36866
rect 41906 36814 41920 36866
rect 41840 36800 41920 36814
rect 0 36546 80 36560
rect 0 36494 14 36546
rect 66 36494 80 36546
rect 0 36480 80 36494
rect 160 36546 240 36560
rect 160 36494 174 36546
rect 226 36494 240 36546
rect 160 36480 240 36494
rect 320 36546 400 36560
rect 320 36494 334 36546
rect 386 36494 400 36546
rect 320 36480 400 36494
rect 480 36546 560 36560
rect 480 36494 494 36546
rect 546 36494 560 36546
rect 480 36480 560 36494
rect 640 36546 720 36560
rect 640 36494 654 36546
rect 706 36494 720 36546
rect 640 36480 720 36494
rect 800 36546 880 36560
rect 800 36494 814 36546
rect 866 36494 880 36546
rect 800 36480 880 36494
rect 960 36546 1040 36560
rect 960 36494 974 36546
rect 1026 36494 1040 36546
rect 960 36480 1040 36494
rect 1120 36546 1200 36560
rect 1120 36494 1134 36546
rect 1186 36494 1200 36546
rect 1120 36480 1200 36494
rect 1280 36546 1360 36560
rect 1280 36494 1294 36546
rect 1346 36494 1360 36546
rect 1280 36480 1360 36494
rect 1440 36546 1520 36560
rect 1440 36494 1454 36546
rect 1506 36494 1520 36546
rect 1440 36480 1520 36494
rect 1600 36546 1680 36560
rect 1600 36494 1614 36546
rect 1666 36494 1680 36546
rect 1600 36480 1680 36494
rect 1760 36546 1840 36560
rect 1760 36494 1774 36546
rect 1826 36494 1840 36546
rect 1760 36480 1840 36494
rect 1920 36546 2000 36560
rect 1920 36494 1934 36546
rect 1986 36494 2000 36546
rect 1920 36480 2000 36494
rect 2080 36546 2160 36560
rect 2080 36494 2094 36546
rect 2146 36494 2160 36546
rect 2080 36480 2160 36494
rect 2240 36546 2320 36560
rect 2240 36494 2254 36546
rect 2306 36494 2320 36546
rect 2240 36480 2320 36494
rect 2400 36546 2480 36560
rect 2400 36494 2414 36546
rect 2466 36494 2480 36546
rect 2400 36480 2480 36494
rect 2560 36546 2640 36560
rect 2560 36494 2574 36546
rect 2626 36494 2640 36546
rect 2560 36480 2640 36494
rect 2720 36546 2800 36560
rect 2720 36494 2734 36546
rect 2786 36494 2800 36546
rect 2720 36480 2800 36494
rect 2880 36546 2960 36560
rect 2880 36494 2894 36546
rect 2946 36494 2960 36546
rect 2880 36480 2960 36494
rect 3040 36546 3120 36560
rect 3040 36494 3054 36546
rect 3106 36494 3120 36546
rect 3040 36480 3120 36494
rect 3200 36546 3280 36560
rect 3200 36494 3214 36546
rect 3266 36494 3280 36546
rect 3200 36480 3280 36494
rect 3360 36546 3440 36560
rect 3360 36494 3374 36546
rect 3426 36494 3440 36546
rect 3360 36480 3440 36494
rect 3520 36546 3600 36560
rect 3520 36494 3534 36546
rect 3586 36494 3600 36546
rect 3520 36480 3600 36494
rect 3680 36546 3760 36560
rect 3680 36494 3694 36546
rect 3746 36494 3760 36546
rect 3680 36480 3760 36494
rect 3840 36546 3920 36560
rect 3840 36494 3854 36546
rect 3906 36494 3920 36546
rect 3840 36480 3920 36494
rect 4000 36546 4080 36560
rect 4000 36494 4014 36546
rect 4066 36494 4080 36546
rect 4000 36480 4080 36494
rect 4160 36546 4240 36560
rect 4160 36494 4174 36546
rect 4226 36494 4240 36546
rect 4160 36480 4240 36494
rect 4320 36546 4400 36560
rect 4320 36494 4334 36546
rect 4386 36494 4400 36546
rect 4320 36480 4400 36494
rect 4480 36546 4560 36560
rect 4480 36494 4494 36546
rect 4546 36494 4560 36546
rect 4480 36480 4560 36494
rect 4640 36546 4720 36560
rect 4640 36494 4654 36546
rect 4706 36494 4720 36546
rect 4640 36480 4720 36494
rect 4800 36546 4880 36560
rect 4800 36494 4814 36546
rect 4866 36494 4880 36546
rect 4800 36480 4880 36494
rect 4960 36546 5040 36560
rect 4960 36494 4974 36546
rect 5026 36494 5040 36546
rect 4960 36480 5040 36494
rect 5120 36546 5200 36560
rect 5120 36494 5134 36546
rect 5186 36494 5200 36546
rect 5120 36480 5200 36494
rect 5280 36546 5360 36560
rect 5280 36494 5294 36546
rect 5346 36494 5360 36546
rect 5280 36480 5360 36494
rect 5440 36546 5520 36560
rect 5440 36494 5454 36546
rect 5506 36494 5520 36546
rect 5440 36480 5520 36494
rect 5600 36546 5680 36560
rect 5600 36494 5614 36546
rect 5666 36494 5680 36546
rect 5600 36480 5680 36494
rect 5760 36546 5840 36560
rect 5760 36494 5774 36546
rect 5826 36494 5840 36546
rect 5760 36480 5840 36494
rect 5920 36546 6000 36560
rect 5920 36494 5934 36546
rect 5986 36494 6000 36546
rect 5920 36480 6000 36494
rect 6080 36546 6160 36560
rect 6080 36494 6094 36546
rect 6146 36494 6160 36546
rect 6080 36480 6160 36494
rect 6240 36546 6320 36560
rect 6240 36494 6254 36546
rect 6306 36494 6320 36546
rect 6240 36480 6320 36494
rect 6400 36546 6480 36560
rect 6400 36494 6414 36546
rect 6466 36494 6480 36546
rect 6400 36480 6480 36494
rect 6560 36546 6640 36560
rect 6560 36494 6574 36546
rect 6626 36494 6640 36546
rect 6560 36480 6640 36494
rect 6720 36546 6800 36560
rect 6720 36494 6734 36546
rect 6786 36494 6800 36546
rect 6720 36480 6800 36494
rect 6880 36546 6960 36560
rect 6880 36494 6894 36546
rect 6946 36494 6960 36546
rect 6880 36480 6960 36494
rect 7040 36546 7120 36560
rect 7040 36494 7054 36546
rect 7106 36494 7120 36546
rect 7040 36480 7120 36494
rect 7200 36546 7280 36560
rect 7200 36494 7214 36546
rect 7266 36494 7280 36546
rect 7200 36480 7280 36494
rect 7360 36546 7440 36560
rect 7360 36494 7374 36546
rect 7426 36494 7440 36546
rect 7360 36480 7440 36494
rect 7520 36546 7600 36560
rect 7520 36494 7534 36546
rect 7586 36494 7600 36546
rect 7520 36480 7600 36494
rect 7680 36546 7760 36560
rect 7680 36494 7694 36546
rect 7746 36494 7760 36546
rect 7680 36480 7760 36494
rect 7840 36546 7920 36560
rect 7840 36494 7854 36546
rect 7906 36494 7920 36546
rect 7840 36480 7920 36494
rect 8000 36546 8080 36560
rect 8000 36494 8014 36546
rect 8066 36494 8080 36546
rect 8000 36480 8080 36494
rect 8160 36546 8240 36560
rect 8160 36494 8174 36546
rect 8226 36494 8240 36546
rect 8160 36480 8240 36494
rect 8320 36546 8400 36560
rect 8320 36494 8334 36546
rect 8386 36494 8400 36546
rect 8320 36480 8400 36494
rect 12480 36546 12560 36560
rect 12480 36494 12494 36546
rect 12546 36494 12560 36546
rect 12480 36480 12560 36494
rect 12640 36546 12720 36560
rect 12640 36494 12654 36546
rect 12706 36494 12720 36546
rect 12640 36480 12720 36494
rect 12800 36546 12880 36560
rect 12800 36494 12814 36546
rect 12866 36494 12880 36546
rect 12800 36480 12880 36494
rect 12960 36546 13040 36560
rect 12960 36494 12974 36546
rect 13026 36494 13040 36546
rect 12960 36480 13040 36494
rect 13120 36546 13200 36560
rect 13120 36494 13134 36546
rect 13186 36494 13200 36546
rect 13120 36480 13200 36494
rect 13280 36546 13360 36560
rect 13280 36494 13294 36546
rect 13346 36494 13360 36546
rect 13280 36480 13360 36494
rect 13440 36546 13520 36560
rect 13440 36494 13454 36546
rect 13506 36494 13520 36546
rect 13440 36480 13520 36494
rect 13600 36546 13680 36560
rect 13600 36494 13614 36546
rect 13666 36494 13680 36546
rect 13600 36480 13680 36494
rect 13760 36546 13840 36560
rect 13760 36494 13774 36546
rect 13826 36494 13840 36546
rect 13760 36480 13840 36494
rect 13920 36546 14000 36560
rect 13920 36494 13934 36546
rect 13986 36494 14000 36546
rect 13920 36480 14000 36494
rect 14080 36546 14160 36560
rect 14080 36494 14094 36546
rect 14146 36494 14160 36546
rect 14080 36480 14160 36494
rect 14240 36546 14320 36560
rect 14240 36494 14254 36546
rect 14306 36494 14320 36546
rect 14240 36480 14320 36494
rect 14400 36546 14480 36560
rect 14400 36494 14414 36546
rect 14466 36494 14480 36546
rect 14400 36480 14480 36494
rect 14560 36546 14640 36560
rect 14560 36494 14574 36546
rect 14626 36494 14640 36546
rect 14560 36480 14640 36494
rect 14720 36546 14800 36560
rect 14720 36494 14734 36546
rect 14786 36494 14800 36546
rect 14720 36480 14800 36494
rect 14880 36546 14960 36560
rect 14880 36494 14894 36546
rect 14946 36494 14960 36546
rect 14880 36480 14960 36494
rect 15040 36546 15120 36560
rect 15040 36494 15054 36546
rect 15106 36494 15120 36546
rect 15040 36480 15120 36494
rect 15200 36546 15280 36560
rect 15200 36494 15214 36546
rect 15266 36494 15280 36546
rect 15200 36480 15280 36494
rect 15360 36546 15440 36560
rect 15360 36494 15374 36546
rect 15426 36494 15440 36546
rect 15360 36480 15440 36494
rect 15520 36546 15600 36560
rect 15520 36494 15534 36546
rect 15586 36494 15600 36546
rect 15520 36480 15600 36494
rect 15680 36546 15760 36560
rect 15680 36494 15694 36546
rect 15746 36494 15760 36546
rect 15680 36480 15760 36494
rect 15840 36546 15920 36560
rect 15840 36494 15854 36546
rect 15906 36494 15920 36546
rect 15840 36480 15920 36494
rect 16000 36546 16080 36560
rect 16000 36494 16014 36546
rect 16066 36494 16080 36546
rect 16000 36480 16080 36494
rect 16160 36546 16240 36560
rect 16160 36494 16174 36546
rect 16226 36494 16240 36546
rect 16160 36480 16240 36494
rect 16320 36546 16400 36560
rect 16320 36494 16334 36546
rect 16386 36494 16400 36546
rect 16320 36480 16400 36494
rect 16480 36546 16560 36560
rect 16480 36494 16494 36546
rect 16546 36494 16560 36546
rect 16480 36480 16560 36494
rect 16640 36546 16720 36560
rect 16640 36494 16654 36546
rect 16706 36494 16720 36546
rect 16640 36480 16720 36494
rect 16800 36546 16880 36560
rect 16800 36494 16814 36546
rect 16866 36494 16880 36546
rect 16800 36480 16880 36494
rect 16960 36546 17040 36560
rect 16960 36494 16974 36546
rect 17026 36494 17040 36546
rect 16960 36480 17040 36494
rect 17120 36546 17200 36560
rect 17120 36494 17134 36546
rect 17186 36494 17200 36546
rect 17120 36480 17200 36494
rect 17280 36546 17360 36560
rect 17280 36494 17294 36546
rect 17346 36494 17360 36546
rect 17280 36480 17360 36494
rect 17440 36546 17520 36560
rect 17440 36494 17454 36546
rect 17506 36494 17520 36546
rect 17440 36480 17520 36494
rect 17600 36546 17680 36560
rect 17600 36494 17614 36546
rect 17666 36494 17680 36546
rect 17600 36480 17680 36494
rect 17760 36546 17840 36560
rect 17760 36494 17774 36546
rect 17826 36494 17840 36546
rect 17760 36480 17840 36494
rect 17920 36546 18000 36560
rect 17920 36494 17934 36546
rect 17986 36494 18000 36546
rect 17920 36480 18000 36494
rect 18080 36546 18160 36560
rect 18080 36494 18094 36546
rect 18146 36494 18160 36546
rect 18080 36480 18160 36494
rect 18240 36546 18320 36560
rect 18240 36494 18254 36546
rect 18306 36494 18320 36546
rect 18240 36480 18320 36494
rect 18400 36546 18480 36560
rect 18400 36494 18414 36546
rect 18466 36494 18480 36546
rect 18400 36480 18480 36494
rect 18560 36546 18640 36560
rect 18560 36494 18574 36546
rect 18626 36494 18640 36546
rect 18560 36480 18640 36494
rect 18720 36546 18800 36560
rect 18720 36494 18734 36546
rect 18786 36494 18800 36546
rect 18720 36480 18800 36494
rect 18880 36546 18960 36560
rect 18880 36494 18894 36546
rect 18946 36494 18960 36546
rect 18880 36480 18960 36494
rect 23120 36546 23200 36560
rect 23120 36494 23134 36546
rect 23186 36494 23200 36546
rect 23120 36480 23200 36494
rect 23280 36546 23360 36560
rect 23280 36494 23294 36546
rect 23346 36494 23360 36546
rect 23280 36480 23360 36494
rect 23440 36546 23520 36560
rect 23440 36494 23454 36546
rect 23506 36494 23520 36546
rect 23440 36480 23520 36494
rect 23600 36546 23680 36560
rect 23600 36494 23614 36546
rect 23666 36494 23680 36546
rect 23600 36480 23680 36494
rect 23760 36546 23840 36560
rect 23760 36494 23774 36546
rect 23826 36494 23840 36546
rect 23760 36480 23840 36494
rect 23920 36546 24000 36560
rect 23920 36494 23934 36546
rect 23986 36494 24000 36546
rect 23920 36480 24000 36494
rect 24080 36546 24160 36560
rect 24080 36494 24094 36546
rect 24146 36494 24160 36546
rect 24080 36480 24160 36494
rect 24240 36546 24320 36560
rect 24240 36494 24254 36546
rect 24306 36494 24320 36546
rect 24240 36480 24320 36494
rect 24400 36546 24480 36560
rect 24400 36494 24414 36546
rect 24466 36494 24480 36546
rect 24400 36480 24480 36494
rect 24560 36546 24640 36560
rect 24560 36494 24574 36546
rect 24626 36494 24640 36546
rect 24560 36480 24640 36494
rect 24720 36546 24800 36560
rect 24720 36494 24734 36546
rect 24786 36494 24800 36546
rect 24720 36480 24800 36494
rect 24880 36546 24960 36560
rect 24880 36494 24894 36546
rect 24946 36494 24960 36546
rect 24880 36480 24960 36494
rect 25040 36546 25120 36560
rect 25040 36494 25054 36546
rect 25106 36494 25120 36546
rect 25040 36480 25120 36494
rect 25200 36546 25280 36560
rect 25200 36494 25214 36546
rect 25266 36494 25280 36546
rect 25200 36480 25280 36494
rect 25360 36546 25440 36560
rect 25360 36494 25374 36546
rect 25426 36494 25440 36546
rect 25360 36480 25440 36494
rect 25520 36546 25600 36560
rect 25520 36494 25534 36546
rect 25586 36494 25600 36546
rect 25520 36480 25600 36494
rect 25680 36546 25760 36560
rect 25680 36494 25694 36546
rect 25746 36494 25760 36546
rect 25680 36480 25760 36494
rect 25840 36546 25920 36560
rect 25840 36494 25854 36546
rect 25906 36494 25920 36546
rect 25840 36480 25920 36494
rect 26000 36546 26080 36560
rect 26000 36494 26014 36546
rect 26066 36494 26080 36546
rect 26000 36480 26080 36494
rect 26160 36546 26240 36560
rect 26160 36494 26174 36546
rect 26226 36494 26240 36546
rect 26160 36480 26240 36494
rect 26320 36546 26400 36560
rect 26320 36494 26334 36546
rect 26386 36494 26400 36546
rect 26320 36480 26400 36494
rect 26480 36546 26560 36560
rect 26480 36494 26494 36546
rect 26546 36494 26560 36546
rect 26480 36480 26560 36494
rect 26640 36546 26720 36560
rect 26640 36494 26654 36546
rect 26706 36494 26720 36546
rect 26640 36480 26720 36494
rect 26800 36546 26880 36560
rect 26800 36494 26814 36546
rect 26866 36494 26880 36546
rect 26800 36480 26880 36494
rect 26960 36546 27040 36560
rect 26960 36494 26974 36546
rect 27026 36494 27040 36546
rect 26960 36480 27040 36494
rect 27120 36546 27200 36560
rect 27120 36494 27134 36546
rect 27186 36494 27200 36546
rect 27120 36480 27200 36494
rect 27280 36546 27360 36560
rect 27280 36494 27294 36546
rect 27346 36494 27360 36546
rect 27280 36480 27360 36494
rect 27440 36546 27520 36560
rect 27440 36494 27454 36546
rect 27506 36494 27520 36546
rect 27440 36480 27520 36494
rect 27600 36546 27680 36560
rect 27600 36494 27614 36546
rect 27666 36494 27680 36546
rect 27600 36480 27680 36494
rect 27760 36546 27840 36560
rect 27760 36494 27774 36546
rect 27826 36494 27840 36546
rect 27760 36480 27840 36494
rect 27920 36546 28000 36560
rect 27920 36494 27934 36546
rect 27986 36494 28000 36546
rect 27920 36480 28000 36494
rect 28080 36546 28160 36560
rect 28080 36494 28094 36546
rect 28146 36494 28160 36546
rect 28080 36480 28160 36494
rect 28240 36546 28320 36560
rect 28240 36494 28254 36546
rect 28306 36494 28320 36546
rect 28240 36480 28320 36494
rect 28400 36546 28480 36560
rect 28400 36494 28414 36546
rect 28466 36494 28480 36546
rect 28400 36480 28480 36494
rect 28560 36546 28640 36560
rect 28560 36494 28574 36546
rect 28626 36494 28640 36546
rect 28560 36480 28640 36494
rect 28720 36546 28800 36560
rect 28720 36494 28734 36546
rect 28786 36494 28800 36546
rect 28720 36480 28800 36494
rect 28880 36546 28960 36560
rect 28880 36494 28894 36546
rect 28946 36494 28960 36546
rect 28880 36480 28960 36494
rect 29040 36546 29120 36560
rect 29040 36494 29054 36546
rect 29106 36494 29120 36546
rect 29040 36480 29120 36494
rect 29200 36546 29280 36560
rect 29200 36494 29214 36546
rect 29266 36494 29280 36546
rect 29200 36480 29280 36494
rect 29360 36546 29440 36560
rect 29360 36494 29374 36546
rect 29426 36494 29440 36546
rect 29360 36480 29440 36494
rect 33520 36546 33600 36560
rect 33520 36494 33534 36546
rect 33586 36494 33600 36546
rect 33520 36480 33600 36494
rect 33680 36546 33760 36560
rect 33680 36494 33694 36546
rect 33746 36494 33760 36546
rect 33680 36480 33760 36494
rect 33840 36546 33920 36560
rect 33840 36494 33854 36546
rect 33906 36494 33920 36546
rect 33840 36480 33920 36494
rect 34000 36546 34080 36560
rect 34000 36494 34014 36546
rect 34066 36494 34080 36546
rect 34000 36480 34080 36494
rect 34160 36546 34240 36560
rect 34160 36494 34174 36546
rect 34226 36494 34240 36546
rect 34160 36480 34240 36494
rect 34320 36546 34400 36560
rect 34320 36494 34334 36546
rect 34386 36494 34400 36546
rect 34320 36480 34400 36494
rect 34480 36546 34560 36560
rect 34480 36494 34494 36546
rect 34546 36494 34560 36546
rect 34480 36480 34560 36494
rect 34640 36546 34720 36560
rect 34640 36494 34654 36546
rect 34706 36494 34720 36546
rect 34640 36480 34720 36494
rect 34800 36546 34880 36560
rect 34800 36494 34814 36546
rect 34866 36494 34880 36546
rect 34800 36480 34880 36494
rect 34960 36546 35040 36560
rect 34960 36494 34974 36546
rect 35026 36494 35040 36546
rect 34960 36480 35040 36494
rect 35120 36546 35200 36560
rect 35120 36494 35134 36546
rect 35186 36494 35200 36546
rect 35120 36480 35200 36494
rect 35280 36546 35360 36560
rect 35280 36494 35294 36546
rect 35346 36494 35360 36546
rect 35280 36480 35360 36494
rect 35440 36546 35520 36560
rect 35440 36494 35454 36546
rect 35506 36494 35520 36546
rect 35440 36480 35520 36494
rect 35600 36546 35680 36560
rect 35600 36494 35614 36546
rect 35666 36494 35680 36546
rect 35600 36480 35680 36494
rect 35760 36546 35840 36560
rect 35760 36494 35774 36546
rect 35826 36494 35840 36546
rect 35760 36480 35840 36494
rect 35920 36546 36000 36560
rect 35920 36494 35934 36546
rect 35986 36494 36000 36546
rect 35920 36480 36000 36494
rect 36080 36546 36160 36560
rect 36080 36494 36094 36546
rect 36146 36494 36160 36546
rect 36080 36480 36160 36494
rect 36240 36546 36320 36560
rect 36240 36494 36254 36546
rect 36306 36494 36320 36546
rect 36240 36480 36320 36494
rect 36400 36546 36480 36560
rect 36400 36494 36414 36546
rect 36466 36494 36480 36546
rect 36400 36480 36480 36494
rect 36560 36546 36640 36560
rect 36560 36494 36574 36546
rect 36626 36494 36640 36546
rect 36560 36480 36640 36494
rect 36720 36546 36800 36560
rect 36720 36494 36734 36546
rect 36786 36494 36800 36546
rect 36720 36480 36800 36494
rect 36880 36546 36960 36560
rect 36880 36494 36894 36546
rect 36946 36494 36960 36546
rect 36880 36480 36960 36494
rect 37040 36546 37120 36560
rect 37040 36494 37054 36546
rect 37106 36494 37120 36546
rect 37040 36480 37120 36494
rect 37200 36546 37280 36560
rect 37200 36494 37214 36546
rect 37266 36494 37280 36546
rect 37200 36480 37280 36494
rect 37360 36546 37440 36560
rect 37360 36494 37374 36546
rect 37426 36494 37440 36546
rect 37360 36480 37440 36494
rect 37520 36546 37600 36560
rect 37520 36494 37534 36546
rect 37586 36494 37600 36546
rect 37520 36480 37600 36494
rect 37680 36546 37760 36560
rect 37680 36494 37694 36546
rect 37746 36494 37760 36546
rect 37680 36480 37760 36494
rect 37840 36546 37920 36560
rect 37840 36494 37854 36546
rect 37906 36494 37920 36546
rect 37840 36480 37920 36494
rect 38000 36546 38080 36560
rect 38000 36494 38014 36546
rect 38066 36494 38080 36546
rect 38000 36480 38080 36494
rect 38160 36546 38240 36560
rect 38160 36494 38174 36546
rect 38226 36494 38240 36546
rect 38160 36480 38240 36494
rect 38320 36546 38400 36560
rect 38320 36494 38334 36546
rect 38386 36494 38400 36546
rect 38320 36480 38400 36494
rect 38480 36546 38560 36560
rect 38480 36494 38494 36546
rect 38546 36494 38560 36546
rect 38480 36480 38560 36494
rect 38640 36546 38720 36560
rect 38640 36494 38654 36546
rect 38706 36494 38720 36546
rect 38640 36480 38720 36494
rect 38800 36546 38880 36560
rect 38800 36494 38814 36546
rect 38866 36494 38880 36546
rect 38800 36480 38880 36494
rect 38960 36546 39040 36560
rect 38960 36494 38974 36546
rect 39026 36494 39040 36546
rect 38960 36480 39040 36494
rect 39120 36546 39200 36560
rect 39120 36494 39134 36546
rect 39186 36494 39200 36546
rect 39120 36480 39200 36494
rect 39280 36546 39360 36560
rect 39280 36494 39294 36546
rect 39346 36494 39360 36546
rect 39280 36480 39360 36494
rect 39440 36546 39520 36560
rect 39440 36494 39454 36546
rect 39506 36494 39520 36546
rect 39440 36480 39520 36494
rect 39600 36546 39680 36560
rect 39600 36494 39614 36546
rect 39666 36494 39680 36546
rect 39600 36480 39680 36494
rect 39760 36546 39840 36560
rect 39760 36494 39774 36546
rect 39826 36494 39840 36546
rect 39760 36480 39840 36494
rect 39920 36546 40000 36560
rect 39920 36494 39934 36546
rect 39986 36494 40000 36546
rect 39920 36480 40000 36494
rect 40080 36546 40160 36560
rect 40080 36494 40094 36546
rect 40146 36494 40160 36546
rect 40080 36480 40160 36494
rect 40240 36546 40320 36560
rect 40240 36494 40254 36546
rect 40306 36494 40320 36546
rect 40240 36480 40320 36494
rect 40400 36546 40480 36560
rect 40400 36494 40414 36546
rect 40466 36494 40480 36546
rect 40400 36480 40480 36494
rect 40560 36546 40640 36560
rect 40560 36494 40574 36546
rect 40626 36494 40640 36546
rect 40560 36480 40640 36494
rect 40720 36546 40800 36560
rect 40720 36494 40734 36546
rect 40786 36494 40800 36546
rect 40720 36480 40800 36494
rect 40880 36546 40960 36560
rect 40880 36494 40894 36546
rect 40946 36494 40960 36546
rect 40880 36480 40960 36494
rect 41040 36546 41120 36560
rect 41040 36494 41054 36546
rect 41106 36494 41120 36546
rect 41040 36480 41120 36494
rect 41200 36546 41280 36560
rect 41200 36494 41214 36546
rect 41266 36494 41280 36546
rect 41200 36480 41280 36494
rect 41360 36546 41440 36560
rect 41360 36494 41374 36546
rect 41426 36494 41440 36546
rect 41360 36480 41440 36494
rect 41520 36546 41600 36560
rect 41520 36494 41534 36546
rect 41586 36494 41600 36546
rect 41520 36480 41600 36494
rect 41680 36546 41760 36560
rect 41680 36494 41694 36546
rect 41746 36494 41760 36546
rect 41680 36480 41760 36494
rect 41840 36546 41920 36560
rect 41840 36494 41854 36546
rect 41906 36494 41920 36546
rect 41840 36480 41920 36494
rect 0 36386 80 36400
rect 0 36334 14 36386
rect 66 36334 80 36386
rect 0 36320 80 36334
rect 160 36386 240 36400
rect 160 36334 174 36386
rect 226 36334 240 36386
rect 160 36320 240 36334
rect 320 36386 400 36400
rect 320 36334 334 36386
rect 386 36334 400 36386
rect 320 36320 400 36334
rect 480 36386 560 36400
rect 480 36334 494 36386
rect 546 36334 560 36386
rect 480 36320 560 36334
rect 640 36386 720 36400
rect 640 36334 654 36386
rect 706 36334 720 36386
rect 640 36320 720 36334
rect 800 36386 880 36400
rect 800 36334 814 36386
rect 866 36334 880 36386
rect 800 36320 880 36334
rect 960 36386 1040 36400
rect 960 36334 974 36386
rect 1026 36334 1040 36386
rect 960 36320 1040 36334
rect 1120 36386 1200 36400
rect 1120 36334 1134 36386
rect 1186 36334 1200 36386
rect 1120 36320 1200 36334
rect 1280 36386 1360 36400
rect 1280 36334 1294 36386
rect 1346 36334 1360 36386
rect 1280 36320 1360 36334
rect 1440 36386 1520 36400
rect 1440 36334 1454 36386
rect 1506 36334 1520 36386
rect 1440 36320 1520 36334
rect 1600 36386 1680 36400
rect 1600 36334 1614 36386
rect 1666 36334 1680 36386
rect 1600 36320 1680 36334
rect 1760 36386 1840 36400
rect 1760 36334 1774 36386
rect 1826 36334 1840 36386
rect 1760 36320 1840 36334
rect 1920 36386 2000 36400
rect 1920 36334 1934 36386
rect 1986 36334 2000 36386
rect 1920 36320 2000 36334
rect 2080 36386 2160 36400
rect 2080 36334 2094 36386
rect 2146 36334 2160 36386
rect 2080 36320 2160 36334
rect 2240 36386 2320 36400
rect 2240 36334 2254 36386
rect 2306 36334 2320 36386
rect 2240 36320 2320 36334
rect 2400 36386 2480 36400
rect 2400 36334 2414 36386
rect 2466 36334 2480 36386
rect 2400 36320 2480 36334
rect 2560 36386 2640 36400
rect 2560 36334 2574 36386
rect 2626 36334 2640 36386
rect 2560 36320 2640 36334
rect 2720 36386 2800 36400
rect 2720 36334 2734 36386
rect 2786 36334 2800 36386
rect 2720 36320 2800 36334
rect 2880 36386 2960 36400
rect 2880 36334 2894 36386
rect 2946 36334 2960 36386
rect 2880 36320 2960 36334
rect 3040 36386 3120 36400
rect 3040 36334 3054 36386
rect 3106 36334 3120 36386
rect 3040 36320 3120 36334
rect 3200 36386 3280 36400
rect 3200 36334 3214 36386
rect 3266 36334 3280 36386
rect 3200 36320 3280 36334
rect 3360 36386 3440 36400
rect 3360 36334 3374 36386
rect 3426 36334 3440 36386
rect 3360 36320 3440 36334
rect 3520 36386 3600 36400
rect 3520 36334 3534 36386
rect 3586 36334 3600 36386
rect 3520 36320 3600 36334
rect 3680 36386 3760 36400
rect 3680 36334 3694 36386
rect 3746 36334 3760 36386
rect 3680 36320 3760 36334
rect 3840 36386 3920 36400
rect 3840 36334 3854 36386
rect 3906 36334 3920 36386
rect 3840 36320 3920 36334
rect 4000 36386 4080 36400
rect 4000 36334 4014 36386
rect 4066 36334 4080 36386
rect 4000 36320 4080 36334
rect 4160 36386 4240 36400
rect 4160 36334 4174 36386
rect 4226 36334 4240 36386
rect 4160 36320 4240 36334
rect 4320 36386 4400 36400
rect 4320 36334 4334 36386
rect 4386 36334 4400 36386
rect 4320 36320 4400 36334
rect 4480 36386 4560 36400
rect 4480 36334 4494 36386
rect 4546 36334 4560 36386
rect 4480 36320 4560 36334
rect 4640 36386 4720 36400
rect 4640 36334 4654 36386
rect 4706 36334 4720 36386
rect 4640 36320 4720 36334
rect 4800 36386 4880 36400
rect 4800 36334 4814 36386
rect 4866 36334 4880 36386
rect 4800 36320 4880 36334
rect 4960 36386 5040 36400
rect 4960 36334 4974 36386
rect 5026 36334 5040 36386
rect 4960 36320 5040 36334
rect 5120 36386 5200 36400
rect 5120 36334 5134 36386
rect 5186 36334 5200 36386
rect 5120 36320 5200 36334
rect 5280 36386 5360 36400
rect 5280 36334 5294 36386
rect 5346 36334 5360 36386
rect 5280 36320 5360 36334
rect 5440 36386 5520 36400
rect 5440 36334 5454 36386
rect 5506 36334 5520 36386
rect 5440 36320 5520 36334
rect 5600 36386 5680 36400
rect 5600 36334 5614 36386
rect 5666 36334 5680 36386
rect 5600 36320 5680 36334
rect 5760 36386 5840 36400
rect 5760 36334 5774 36386
rect 5826 36334 5840 36386
rect 5760 36320 5840 36334
rect 5920 36386 6000 36400
rect 5920 36334 5934 36386
rect 5986 36334 6000 36386
rect 5920 36320 6000 36334
rect 6080 36386 6160 36400
rect 6080 36334 6094 36386
rect 6146 36334 6160 36386
rect 6080 36320 6160 36334
rect 6240 36386 6320 36400
rect 6240 36334 6254 36386
rect 6306 36334 6320 36386
rect 6240 36320 6320 36334
rect 6400 36386 6480 36400
rect 6400 36334 6414 36386
rect 6466 36334 6480 36386
rect 6400 36320 6480 36334
rect 6560 36386 6640 36400
rect 6560 36334 6574 36386
rect 6626 36334 6640 36386
rect 6560 36320 6640 36334
rect 6720 36386 6800 36400
rect 6720 36334 6734 36386
rect 6786 36334 6800 36386
rect 6720 36320 6800 36334
rect 6880 36386 6960 36400
rect 6880 36334 6894 36386
rect 6946 36334 6960 36386
rect 6880 36320 6960 36334
rect 7040 36386 7120 36400
rect 7040 36334 7054 36386
rect 7106 36334 7120 36386
rect 7040 36320 7120 36334
rect 7200 36386 7280 36400
rect 7200 36334 7214 36386
rect 7266 36334 7280 36386
rect 7200 36320 7280 36334
rect 7360 36386 7440 36400
rect 7360 36334 7374 36386
rect 7426 36334 7440 36386
rect 7360 36320 7440 36334
rect 7520 36386 7600 36400
rect 7520 36334 7534 36386
rect 7586 36334 7600 36386
rect 7520 36320 7600 36334
rect 7680 36386 7760 36400
rect 7680 36334 7694 36386
rect 7746 36334 7760 36386
rect 7680 36320 7760 36334
rect 7840 36386 7920 36400
rect 7840 36334 7854 36386
rect 7906 36334 7920 36386
rect 7840 36320 7920 36334
rect 8000 36386 8080 36400
rect 8000 36334 8014 36386
rect 8066 36334 8080 36386
rect 8000 36320 8080 36334
rect 8160 36386 8240 36400
rect 8160 36334 8174 36386
rect 8226 36334 8240 36386
rect 8160 36320 8240 36334
rect 8320 36386 8400 36400
rect 8320 36334 8334 36386
rect 8386 36334 8400 36386
rect 8320 36320 8400 36334
rect 12480 36386 12560 36400
rect 12480 36334 12494 36386
rect 12546 36334 12560 36386
rect 12480 36320 12560 36334
rect 12640 36386 12720 36400
rect 12640 36334 12654 36386
rect 12706 36334 12720 36386
rect 12640 36320 12720 36334
rect 12800 36386 12880 36400
rect 12800 36334 12814 36386
rect 12866 36334 12880 36386
rect 12800 36320 12880 36334
rect 12960 36386 13040 36400
rect 12960 36334 12974 36386
rect 13026 36334 13040 36386
rect 12960 36320 13040 36334
rect 13120 36386 13200 36400
rect 13120 36334 13134 36386
rect 13186 36334 13200 36386
rect 13120 36320 13200 36334
rect 13280 36386 13360 36400
rect 13280 36334 13294 36386
rect 13346 36334 13360 36386
rect 13280 36320 13360 36334
rect 13440 36386 13520 36400
rect 13440 36334 13454 36386
rect 13506 36334 13520 36386
rect 13440 36320 13520 36334
rect 13600 36386 13680 36400
rect 13600 36334 13614 36386
rect 13666 36334 13680 36386
rect 13600 36320 13680 36334
rect 13760 36386 13840 36400
rect 13760 36334 13774 36386
rect 13826 36334 13840 36386
rect 13760 36320 13840 36334
rect 13920 36386 14000 36400
rect 13920 36334 13934 36386
rect 13986 36334 14000 36386
rect 13920 36320 14000 36334
rect 14080 36386 14160 36400
rect 14080 36334 14094 36386
rect 14146 36334 14160 36386
rect 14080 36320 14160 36334
rect 14240 36386 14320 36400
rect 14240 36334 14254 36386
rect 14306 36334 14320 36386
rect 14240 36320 14320 36334
rect 14400 36386 14480 36400
rect 14400 36334 14414 36386
rect 14466 36334 14480 36386
rect 14400 36320 14480 36334
rect 14560 36386 14640 36400
rect 14560 36334 14574 36386
rect 14626 36334 14640 36386
rect 14560 36320 14640 36334
rect 14720 36386 14800 36400
rect 14720 36334 14734 36386
rect 14786 36334 14800 36386
rect 14720 36320 14800 36334
rect 14880 36386 14960 36400
rect 14880 36334 14894 36386
rect 14946 36334 14960 36386
rect 14880 36320 14960 36334
rect 15040 36386 15120 36400
rect 15040 36334 15054 36386
rect 15106 36334 15120 36386
rect 15040 36320 15120 36334
rect 15200 36386 15280 36400
rect 15200 36334 15214 36386
rect 15266 36334 15280 36386
rect 15200 36320 15280 36334
rect 15360 36386 15440 36400
rect 15360 36334 15374 36386
rect 15426 36334 15440 36386
rect 15360 36320 15440 36334
rect 15520 36386 15600 36400
rect 15520 36334 15534 36386
rect 15586 36334 15600 36386
rect 15520 36320 15600 36334
rect 15680 36386 15760 36400
rect 15680 36334 15694 36386
rect 15746 36334 15760 36386
rect 15680 36320 15760 36334
rect 15840 36386 15920 36400
rect 15840 36334 15854 36386
rect 15906 36334 15920 36386
rect 15840 36320 15920 36334
rect 16000 36386 16080 36400
rect 16000 36334 16014 36386
rect 16066 36334 16080 36386
rect 16000 36320 16080 36334
rect 16160 36386 16240 36400
rect 16160 36334 16174 36386
rect 16226 36334 16240 36386
rect 16160 36320 16240 36334
rect 16320 36386 16400 36400
rect 16320 36334 16334 36386
rect 16386 36334 16400 36386
rect 16320 36320 16400 36334
rect 16480 36386 16560 36400
rect 16480 36334 16494 36386
rect 16546 36334 16560 36386
rect 16480 36320 16560 36334
rect 16640 36386 16720 36400
rect 16640 36334 16654 36386
rect 16706 36334 16720 36386
rect 16640 36320 16720 36334
rect 16800 36386 16880 36400
rect 16800 36334 16814 36386
rect 16866 36334 16880 36386
rect 16800 36320 16880 36334
rect 16960 36386 17040 36400
rect 16960 36334 16974 36386
rect 17026 36334 17040 36386
rect 16960 36320 17040 36334
rect 17120 36386 17200 36400
rect 17120 36334 17134 36386
rect 17186 36334 17200 36386
rect 17120 36320 17200 36334
rect 17280 36386 17360 36400
rect 17280 36334 17294 36386
rect 17346 36334 17360 36386
rect 17280 36320 17360 36334
rect 17440 36386 17520 36400
rect 17440 36334 17454 36386
rect 17506 36334 17520 36386
rect 17440 36320 17520 36334
rect 17600 36386 17680 36400
rect 17600 36334 17614 36386
rect 17666 36334 17680 36386
rect 17600 36320 17680 36334
rect 17760 36386 17840 36400
rect 17760 36334 17774 36386
rect 17826 36334 17840 36386
rect 17760 36320 17840 36334
rect 17920 36386 18000 36400
rect 17920 36334 17934 36386
rect 17986 36334 18000 36386
rect 17920 36320 18000 36334
rect 18080 36386 18160 36400
rect 18080 36334 18094 36386
rect 18146 36334 18160 36386
rect 18080 36320 18160 36334
rect 18240 36386 18320 36400
rect 18240 36334 18254 36386
rect 18306 36334 18320 36386
rect 18240 36320 18320 36334
rect 18400 36386 18480 36400
rect 18400 36334 18414 36386
rect 18466 36334 18480 36386
rect 18400 36320 18480 36334
rect 18560 36386 18640 36400
rect 18560 36334 18574 36386
rect 18626 36334 18640 36386
rect 18560 36320 18640 36334
rect 18720 36386 18800 36400
rect 18720 36334 18734 36386
rect 18786 36334 18800 36386
rect 18720 36320 18800 36334
rect 18880 36386 18960 36400
rect 18880 36334 18894 36386
rect 18946 36334 18960 36386
rect 18880 36320 18960 36334
rect 23120 36386 23200 36400
rect 23120 36334 23134 36386
rect 23186 36334 23200 36386
rect 23120 36320 23200 36334
rect 23280 36386 23360 36400
rect 23280 36334 23294 36386
rect 23346 36334 23360 36386
rect 23280 36320 23360 36334
rect 23440 36386 23520 36400
rect 23440 36334 23454 36386
rect 23506 36334 23520 36386
rect 23440 36320 23520 36334
rect 23600 36386 23680 36400
rect 23600 36334 23614 36386
rect 23666 36334 23680 36386
rect 23600 36320 23680 36334
rect 23760 36386 23840 36400
rect 23760 36334 23774 36386
rect 23826 36334 23840 36386
rect 23760 36320 23840 36334
rect 23920 36386 24000 36400
rect 23920 36334 23934 36386
rect 23986 36334 24000 36386
rect 23920 36320 24000 36334
rect 24080 36386 24160 36400
rect 24080 36334 24094 36386
rect 24146 36334 24160 36386
rect 24080 36320 24160 36334
rect 24240 36386 24320 36400
rect 24240 36334 24254 36386
rect 24306 36334 24320 36386
rect 24240 36320 24320 36334
rect 24400 36386 24480 36400
rect 24400 36334 24414 36386
rect 24466 36334 24480 36386
rect 24400 36320 24480 36334
rect 24560 36386 24640 36400
rect 24560 36334 24574 36386
rect 24626 36334 24640 36386
rect 24560 36320 24640 36334
rect 24720 36386 24800 36400
rect 24720 36334 24734 36386
rect 24786 36334 24800 36386
rect 24720 36320 24800 36334
rect 24880 36386 24960 36400
rect 24880 36334 24894 36386
rect 24946 36334 24960 36386
rect 24880 36320 24960 36334
rect 25040 36386 25120 36400
rect 25040 36334 25054 36386
rect 25106 36334 25120 36386
rect 25040 36320 25120 36334
rect 25200 36386 25280 36400
rect 25200 36334 25214 36386
rect 25266 36334 25280 36386
rect 25200 36320 25280 36334
rect 25360 36386 25440 36400
rect 25360 36334 25374 36386
rect 25426 36334 25440 36386
rect 25360 36320 25440 36334
rect 25520 36386 25600 36400
rect 25520 36334 25534 36386
rect 25586 36334 25600 36386
rect 25520 36320 25600 36334
rect 25680 36386 25760 36400
rect 25680 36334 25694 36386
rect 25746 36334 25760 36386
rect 25680 36320 25760 36334
rect 25840 36386 25920 36400
rect 25840 36334 25854 36386
rect 25906 36334 25920 36386
rect 25840 36320 25920 36334
rect 26000 36386 26080 36400
rect 26000 36334 26014 36386
rect 26066 36334 26080 36386
rect 26000 36320 26080 36334
rect 26160 36386 26240 36400
rect 26160 36334 26174 36386
rect 26226 36334 26240 36386
rect 26160 36320 26240 36334
rect 26320 36386 26400 36400
rect 26320 36334 26334 36386
rect 26386 36334 26400 36386
rect 26320 36320 26400 36334
rect 26480 36386 26560 36400
rect 26480 36334 26494 36386
rect 26546 36334 26560 36386
rect 26480 36320 26560 36334
rect 26640 36386 26720 36400
rect 26640 36334 26654 36386
rect 26706 36334 26720 36386
rect 26640 36320 26720 36334
rect 26800 36386 26880 36400
rect 26800 36334 26814 36386
rect 26866 36334 26880 36386
rect 26800 36320 26880 36334
rect 26960 36386 27040 36400
rect 26960 36334 26974 36386
rect 27026 36334 27040 36386
rect 26960 36320 27040 36334
rect 27120 36386 27200 36400
rect 27120 36334 27134 36386
rect 27186 36334 27200 36386
rect 27120 36320 27200 36334
rect 27280 36386 27360 36400
rect 27280 36334 27294 36386
rect 27346 36334 27360 36386
rect 27280 36320 27360 36334
rect 27440 36386 27520 36400
rect 27440 36334 27454 36386
rect 27506 36334 27520 36386
rect 27440 36320 27520 36334
rect 27600 36386 27680 36400
rect 27600 36334 27614 36386
rect 27666 36334 27680 36386
rect 27600 36320 27680 36334
rect 27760 36386 27840 36400
rect 27760 36334 27774 36386
rect 27826 36334 27840 36386
rect 27760 36320 27840 36334
rect 27920 36386 28000 36400
rect 27920 36334 27934 36386
rect 27986 36334 28000 36386
rect 27920 36320 28000 36334
rect 28080 36386 28160 36400
rect 28080 36334 28094 36386
rect 28146 36334 28160 36386
rect 28080 36320 28160 36334
rect 28240 36386 28320 36400
rect 28240 36334 28254 36386
rect 28306 36334 28320 36386
rect 28240 36320 28320 36334
rect 28400 36386 28480 36400
rect 28400 36334 28414 36386
rect 28466 36334 28480 36386
rect 28400 36320 28480 36334
rect 28560 36386 28640 36400
rect 28560 36334 28574 36386
rect 28626 36334 28640 36386
rect 28560 36320 28640 36334
rect 28720 36386 28800 36400
rect 28720 36334 28734 36386
rect 28786 36334 28800 36386
rect 28720 36320 28800 36334
rect 28880 36386 28960 36400
rect 28880 36334 28894 36386
rect 28946 36334 28960 36386
rect 28880 36320 28960 36334
rect 29040 36386 29120 36400
rect 29040 36334 29054 36386
rect 29106 36334 29120 36386
rect 29040 36320 29120 36334
rect 29200 36386 29280 36400
rect 29200 36334 29214 36386
rect 29266 36334 29280 36386
rect 29200 36320 29280 36334
rect 29360 36386 29440 36400
rect 29360 36334 29374 36386
rect 29426 36334 29440 36386
rect 29360 36320 29440 36334
rect 33520 36386 33600 36400
rect 33520 36334 33534 36386
rect 33586 36334 33600 36386
rect 33520 36320 33600 36334
rect 33680 36386 33760 36400
rect 33680 36334 33694 36386
rect 33746 36334 33760 36386
rect 33680 36320 33760 36334
rect 33840 36386 33920 36400
rect 33840 36334 33854 36386
rect 33906 36334 33920 36386
rect 33840 36320 33920 36334
rect 34000 36386 34080 36400
rect 34000 36334 34014 36386
rect 34066 36334 34080 36386
rect 34000 36320 34080 36334
rect 34160 36386 34240 36400
rect 34160 36334 34174 36386
rect 34226 36334 34240 36386
rect 34160 36320 34240 36334
rect 34320 36386 34400 36400
rect 34320 36334 34334 36386
rect 34386 36334 34400 36386
rect 34320 36320 34400 36334
rect 34480 36386 34560 36400
rect 34480 36334 34494 36386
rect 34546 36334 34560 36386
rect 34480 36320 34560 36334
rect 34640 36386 34720 36400
rect 34640 36334 34654 36386
rect 34706 36334 34720 36386
rect 34640 36320 34720 36334
rect 34800 36386 34880 36400
rect 34800 36334 34814 36386
rect 34866 36334 34880 36386
rect 34800 36320 34880 36334
rect 34960 36386 35040 36400
rect 34960 36334 34974 36386
rect 35026 36334 35040 36386
rect 34960 36320 35040 36334
rect 35120 36386 35200 36400
rect 35120 36334 35134 36386
rect 35186 36334 35200 36386
rect 35120 36320 35200 36334
rect 35280 36386 35360 36400
rect 35280 36334 35294 36386
rect 35346 36334 35360 36386
rect 35280 36320 35360 36334
rect 35440 36386 35520 36400
rect 35440 36334 35454 36386
rect 35506 36334 35520 36386
rect 35440 36320 35520 36334
rect 35600 36386 35680 36400
rect 35600 36334 35614 36386
rect 35666 36334 35680 36386
rect 35600 36320 35680 36334
rect 35760 36386 35840 36400
rect 35760 36334 35774 36386
rect 35826 36334 35840 36386
rect 35760 36320 35840 36334
rect 35920 36386 36000 36400
rect 35920 36334 35934 36386
rect 35986 36334 36000 36386
rect 35920 36320 36000 36334
rect 36080 36386 36160 36400
rect 36080 36334 36094 36386
rect 36146 36334 36160 36386
rect 36080 36320 36160 36334
rect 36240 36386 36320 36400
rect 36240 36334 36254 36386
rect 36306 36334 36320 36386
rect 36240 36320 36320 36334
rect 36400 36386 36480 36400
rect 36400 36334 36414 36386
rect 36466 36334 36480 36386
rect 36400 36320 36480 36334
rect 36560 36386 36640 36400
rect 36560 36334 36574 36386
rect 36626 36334 36640 36386
rect 36560 36320 36640 36334
rect 36720 36386 36800 36400
rect 36720 36334 36734 36386
rect 36786 36334 36800 36386
rect 36720 36320 36800 36334
rect 36880 36386 36960 36400
rect 36880 36334 36894 36386
rect 36946 36334 36960 36386
rect 36880 36320 36960 36334
rect 37040 36386 37120 36400
rect 37040 36334 37054 36386
rect 37106 36334 37120 36386
rect 37040 36320 37120 36334
rect 37200 36386 37280 36400
rect 37200 36334 37214 36386
rect 37266 36334 37280 36386
rect 37200 36320 37280 36334
rect 37360 36386 37440 36400
rect 37360 36334 37374 36386
rect 37426 36334 37440 36386
rect 37360 36320 37440 36334
rect 37520 36386 37600 36400
rect 37520 36334 37534 36386
rect 37586 36334 37600 36386
rect 37520 36320 37600 36334
rect 37680 36386 37760 36400
rect 37680 36334 37694 36386
rect 37746 36334 37760 36386
rect 37680 36320 37760 36334
rect 37840 36386 37920 36400
rect 37840 36334 37854 36386
rect 37906 36334 37920 36386
rect 37840 36320 37920 36334
rect 38000 36386 38080 36400
rect 38000 36334 38014 36386
rect 38066 36334 38080 36386
rect 38000 36320 38080 36334
rect 38160 36386 38240 36400
rect 38160 36334 38174 36386
rect 38226 36334 38240 36386
rect 38160 36320 38240 36334
rect 38320 36386 38400 36400
rect 38320 36334 38334 36386
rect 38386 36334 38400 36386
rect 38320 36320 38400 36334
rect 38480 36386 38560 36400
rect 38480 36334 38494 36386
rect 38546 36334 38560 36386
rect 38480 36320 38560 36334
rect 38640 36386 38720 36400
rect 38640 36334 38654 36386
rect 38706 36334 38720 36386
rect 38640 36320 38720 36334
rect 38800 36386 38880 36400
rect 38800 36334 38814 36386
rect 38866 36334 38880 36386
rect 38800 36320 38880 36334
rect 38960 36386 39040 36400
rect 38960 36334 38974 36386
rect 39026 36334 39040 36386
rect 38960 36320 39040 36334
rect 39120 36386 39200 36400
rect 39120 36334 39134 36386
rect 39186 36334 39200 36386
rect 39120 36320 39200 36334
rect 39280 36386 39360 36400
rect 39280 36334 39294 36386
rect 39346 36334 39360 36386
rect 39280 36320 39360 36334
rect 39440 36386 39520 36400
rect 39440 36334 39454 36386
rect 39506 36334 39520 36386
rect 39440 36320 39520 36334
rect 39600 36386 39680 36400
rect 39600 36334 39614 36386
rect 39666 36334 39680 36386
rect 39600 36320 39680 36334
rect 39760 36386 39840 36400
rect 39760 36334 39774 36386
rect 39826 36334 39840 36386
rect 39760 36320 39840 36334
rect 39920 36386 40000 36400
rect 39920 36334 39934 36386
rect 39986 36334 40000 36386
rect 39920 36320 40000 36334
rect 40080 36386 40160 36400
rect 40080 36334 40094 36386
rect 40146 36334 40160 36386
rect 40080 36320 40160 36334
rect 40240 36386 40320 36400
rect 40240 36334 40254 36386
rect 40306 36334 40320 36386
rect 40240 36320 40320 36334
rect 40400 36386 40480 36400
rect 40400 36334 40414 36386
rect 40466 36334 40480 36386
rect 40400 36320 40480 36334
rect 40560 36386 40640 36400
rect 40560 36334 40574 36386
rect 40626 36334 40640 36386
rect 40560 36320 40640 36334
rect 40720 36386 40800 36400
rect 40720 36334 40734 36386
rect 40786 36334 40800 36386
rect 40720 36320 40800 36334
rect 40880 36386 40960 36400
rect 40880 36334 40894 36386
rect 40946 36334 40960 36386
rect 40880 36320 40960 36334
rect 41040 36386 41120 36400
rect 41040 36334 41054 36386
rect 41106 36334 41120 36386
rect 41040 36320 41120 36334
rect 41200 36386 41280 36400
rect 41200 36334 41214 36386
rect 41266 36334 41280 36386
rect 41200 36320 41280 36334
rect 41360 36386 41440 36400
rect 41360 36334 41374 36386
rect 41426 36334 41440 36386
rect 41360 36320 41440 36334
rect 41520 36386 41600 36400
rect 41520 36334 41534 36386
rect 41586 36334 41600 36386
rect 41520 36320 41600 36334
rect 41680 36386 41760 36400
rect 41680 36334 41694 36386
rect 41746 36334 41760 36386
rect 41680 36320 41760 36334
rect 41840 36386 41920 36400
rect 41840 36334 41854 36386
rect 41906 36334 41920 36386
rect 41840 36320 41920 36334
rect 0 36066 80 36080
rect 0 36014 14 36066
rect 66 36014 80 36066
rect 0 36000 80 36014
rect 160 36066 240 36080
rect 160 36014 174 36066
rect 226 36014 240 36066
rect 160 36000 240 36014
rect 320 36066 400 36080
rect 320 36014 334 36066
rect 386 36014 400 36066
rect 320 36000 400 36014
rect 480 36066 560 36080
rect 480 36014 494 36066
rect 546 36014 560 36066
rect 480 36000 560 36014
rect 640 36066 720 36080
rect 640 36014 654 36066
rect 706 36014 720 36066
rect 640 36000 720 36014
rect 800 36066 880 36080
rect 800 36014 814 36066
rect 866 36014 880 36066
rect 800 36000 880 36014
rect 960 36066 1040 36080
rect 960 36014 974 36066
rect 1026 36014 1040 36066
rect 960 36000 1040 36014
rect 1120 36066 1200 36080
rect 1120 36014 1134 36066
rect 1186 36014 1200 36066
rect 1120 36000 1200 36014
rect 1280 36066 1360 36080
rect 1280 36014 1294 36066
rect 1346 36014 1360 36066
rect 1280 36000 1360 36014
rect 1440 36066 1520 36080
rect 1440 36014 1454 36066
rect 1506 36014 1520 36066
rect 1440 36000 1520 36014
rect 1600 36066 1680 36080
rect 1600 36014 1614 36066
rect 1666 36014 1680 36066
rect 1600 36000 1680 36014
rect 1760 36066 1840 36080
rect 1760 36014 1774 36066
rect 1826 36014 1840 36066
rect 1760 36000 1840 36014
rect 1920 36066 2000 36080
rect 1920 36014 1934 36066
rect 1986 36014 2000 36066
rect 1920 36000 2000 36014
rect 2080 36066 2160 36080
rect 2080 36014 2094 36066
rect 2146 36014 2160 36066
rect 2080 36000 2160 36014
rect 2240 36066 2320 36080
rect 2240 36014 2254 36066
rect 2306 36014 2320 36066
rect 2240 36000 2320 36014
rect 2400 36066 2480 36080
rect 2400 36014 2414 36066
rect 2466 36014 2480 36066
rect 2400 36000 2480 36014
rect 2560 36066 2640 36080
rect 2560 36014 2574 36066
rect 2626 36014 2640 36066
rect 2560 36000 2640 36014
rect 2720 36066 2800 36080
rect 2720 36014 2734 36066
rect 2786 36014 2800 36066
rect 2720 36000 2800 36014
rect 2880 36066 2960 36080
rect 2880 36014 2894 36066
rect 2946 36014 2960 36066
rect 2880 36000 2960 36014
rect 3040 36066 3120 36080
rect 3040 36014 3054 36066
rect 3106 36014 3120 36066
rect 3040 36000 3120 36014
rect 3200 36066 3280 36080
rect 3200 36014 3214 36066
rect 3266 36014 3280 36066
rect 3200 36000 3280 36014
rect 3360 36066 3440 36080
rect 3360 36014 3374 36066
rect 3426 36014 3440 36066
rect 3360 36000 3440 36014
rect 3520 36066 3600 36080
rect 3520 36014 3534 36066
rect 3586 36014 3600 36066
rect 3520 36000 3600 36014
rect 3680 36066 3760 36080
rect 3680 36014 3694 36066
rect 3746 36014 3760 36066
rect 3680 36000 3760 36014
rect 3840 36066 3920 36080
rect 3840 36014 3854 36066
rect 3906 36014 3920 36066
rect 3840 36000 3920 36014
rect 4000 36066 4080 36080
rect 4000 36014 4014 36066
rect 4066 36014 4080 36066
rect 4000 36000 4080 36014
rect 4160 36066 4240 36080
rect 4160 36014 4174 36066
rect 4226 36014 4240 36066
rect 4160 36000 4240 36014
rect 4320 36066 4400 36080
rect 4320 36014 4334 36066
rect 4386 36014 4400 36066
rect 4320 36000 4400 36014
rect 4480 36066 4560 36080
rect 4480 36014 4494 36066
rect 4546 36014 4560 36066
rect 4480 36000 4560 36014
rect 4640 36066 4720 36080
rect 4640 36014 4654 36066
rect 4706 36014 4720 36066
rect 4640 36000 4720 36014
rect 4800 36066 4880 36080
rect 4800 36014 4814 36066
rect 4866 36014 4880 36066
rect 4800 36000 4880 36014
rect 4960 36066 5040 36080
rect 4960 36014 4974 36066
rect 5026 36014 5040 36066
rect 4960 36000 5040 36014
rect 5120 36066 5200 36080
rect 5120 36014 5134 36066
rect 5186 36014 5200 36066
rect 5120 36000 5200 36014
rect 5280 36066 5360 36080
rect 5280 36014 5294 36066
rect 5346 36014 5360 36066
rect 5280 36000 5360 36014
rect 5440 36066 5520 36080
rect 5440 36014 5454 36066
rect 5506 36014 5520 36066
rect 5440 36000 5520 36014
rect 5600 36066 5680 36080
rect 5600 36014 5614 36066
rect 5666 36014 5680 36066
rect 5600 36000 5680 36014
rect 5760 36066 5840 36080
rect 5760 36014 5774 36066
rect 5826 36014 5840 36066
rect 5760 36000 5840 36014
rect 5920 36066 6000 36080
rect 5920 36014 5934 36066
rect 5986 36014 6000 36066
rect 5920 36000 6000 36014
rect 6080 36066 6160 36080
rect 6080 36014 6094 36066
rect 6146 36014 6160 36066
rect 6080 36000 6160 36014
rect 6240 36066 6320 36080
rect 6240 36014 6254 36066
rect 6306 36014 6320 36066
rect 6240 36000 6320 36014
rect 6400 36066 6480 36080
rect 6400 36014 6414 36066
rect 6466 36014 6480 36066
rect 6400 36000 6480 36014
rect 6560 36066 6640 36080
rect 6560 36014 6574 36066
rect 6626 36014 6640 36066
rect 6560 36000 6640 36014
rect 6720 36066 6800 36080
rect 6720 36014 6734 36066
rect 6786 36014 6800 36066
rect 6720 36000 6800 36014
rect 6880 36066 6960 36080
rect 6880 36014 6894 36066
rect 6946 36014 6960 36066
rect 6880 36000 6960 36014
rect 7040 36066 7120 36080
rect 7040 36014 7054 36066
rect 7106 36014 7120 36066
rect 7040 36000 7120 36014
rect 7200 36066 7280 36080
rect 7200 36014 7214 36066
rect 7266 36014 7280 36066
rect 7200 36000 7280 36014
rect 7360 36066 7440 36080
rect 7360 36014 7374 36066
rect 7426 36014 7440 36066
rect 7360 36000 7440 36014
rect 7520 36066 7600 36080
rect 7520 36014 7534 36066
rect 7586 36014 7600 36066
rect 7520 36000 7600 36014
rect 7680 36066 7760 36080
rect 7680 36014 7694 36066
rect 7746 36014 7760 36066
rect 7680 36000 7760 36014
rect 7840 36066 7920 36080
rect 7840 36014 7854 36066
rect 7906 36014 7920 36066
rect 7840 36000 7920 36014
rect 8000 36066 8080 36080
rect 8000 36014 8014 36066
rect 8066 36014 8080 36066
rect 8000 36000 8080 36014
rect 8160 36066 8240 36080
rect 8160 36014 8174 36066
rect 8226 36014 8240 36066
rect 8160 36000 8240 36014
rect 8320 36066 8400 36080
rect 8320 36014 8334 36066
rect 8386 36014 8400 36066
rect 8320 36000 8400 36014
rect 12480 36066 12560 36080
rect 12480 36014 12494 36066
rect 12546 36014 12560 36066
rect 12480 36000 12560 36014
rect 12640 36066 12720 36080
rect 12640 36014 12654 36066
rect 12706 36014 12720 36066
rect 12640 36000 12720 36014
rect 12800 36066 12880 36080
rect 12800 36014 12814 36066
rect 12866 36014 12880 36066
rect 12800 36000 12880 36014
rect 12960 36066 13040 36080
rect 12960 36014 12974 36066
rect 13026 36014 13040 36066
rect 12960 36000 13040 36014
rect 13120 36066 13200 36080
rect 13120 36014 13134 36066
rect 13186 36014 13200 36066
rect 13120 36000 13200 36014
rect 13280 36066 13360 36080
rect 13280 36014 13294 36066
rect 13346 36014 13360 36066
rect 13280 36000 13360 36014
rect 13440 36066 13520 36080
rect 13440 36014 13454 36066
rect 13506 36014 13520 36066
rect 13440 36000 13520 36014
rect 13600 36066 13680 36080
rect 13600 36014 13614 36066
rect 13666 36014 13680 36066
rect 13600 36000 13680 36014
rect 13760 36066 13840 36080
rect 13760 36014 13774 36066
rect 13826 36014 13840 36066
rect 13760 36000 13840 36014
rect 13920 36066 14000 36080
rect 13920 36014 13934 36066
rect 13986 36014 14000 36066
rect 13920 36000 14000 36014
rect 14080 36066 14160 36080
rect 14080 36014 14094 36066
rect 14146 36014 14160 36066
rect 14080 36000 14160 36014
rect 14240 36066 14320 36080
rect 14240 36014 14254 36066
rect 14306 36014 14320 36066
rect 14240 36000 14320 36014
rect 14400 36066 14480 36080
rect 14400 36014 14414 36066
rect 14466 36014 14480 36066
rect 14400 36000 14480 36014
rect 14560 36066 14640 36080
rect 14560 36014 14574 36066
rect 14626 36014 14640 36066
rect 14560 36000 14640 36014
rect 14720 36066 14800 36080
rect 14720 36014 14734 36066
rect 14786 36014 14800 36066
rect 14720 36000 14800 36014
rect 14880 36066 14960 36080
rect 14880 36014 14894 36066
rect 14946 36014 14960 36066
rect 14880 36000 14960 36014
rect 15040 36066 15120 36080
rect 15040 36014 15054 36066
rect 15106 36014 15120 36066
rect 15040 36000 15120 36014
rect 15200 36066 15280 36080
rect 15200 36014 15214 36066
rect 15266 36014 15280 36066
rect 15200 36000 15280 36014
rect 15360 36066 15440 36080
rect 15360 36014 15374 36066
rect 15426 36014 15440 36066
rect 15360 36000 15440 36014
rect 15520 36066 15600 36080
rect 15520 36014 15534 36066
rect 15586 36014 15600 36066
rect 15520 36000 15600 36014
rect 15680 36066 15760 36080
rect 15680 36014 15694 36066
rect 15746 36014 15760 36066
rect 15680 36000 15760 36014
rect 15840 36066 15920 36080
rect 15840 36014 15854 36066
rect 15906 36014 15920 36066
rect 15840 36000 15920 36014
rect 16000 36066 16080 36080
rect 16000 36014 16014 36066
rect 16066 36014 16080 36066
rect 16000 36000 16080 36014
rect 16160 36066 16240 36080
rect 16160 36014 16174 36066
rect 16226 36014 16240 36066
rect 16160 36000 16240 36014
rect 16320 36066 16400 36080
rect 16320 36014 16334 36066
rect 16386 36014 16400 36066
rect 16320 36000 16400 36014
rect 16480 36066 16560 36080
rect 16480 36014 16494 36066
rect 16546 36014 16560 36066
rect 16480 36000 16560 36014
rect 16640 36066 16720 36080
rect 16640 36014 16654 36066
rect 16706 36014 16720 36066
rect 16640 36000 16720 36014
rect 16800 36066 16880 36080
rect 16800 36014 16814 36066
rect 16866 36014 16880 36066
rect 16800 36000 16880 36014
rect 16960 36066 17040 36080
rect 16960 36014 16974 36066
rect 17026 36014 17040 36066
rect 16960 36000 17040 36014
rect 17120 36066 17200 36080
rect 17120 36014 17134 36066
rect 17186 36014 17200 36066
rect 17120 36000 17200 36014
rect 17280 36066 17360 36080
rect 17280 36014 17294 36066
rect 17346 36014 17360 36066
rect 17280 36000 17360 36014
rect 17440 36066 17520 36080
rect 17440 36014 17454 36066
rect 17506 36014 17520 36066
rect 17440 36000 17520 36014
rect 17600 36066 17680 36080
rect 17600 36014 17614 36066
rect 17666 36014 17680 36066
rect 17600 36000 17680 36014
rect 17760 36066 17840 36080
rect 17760 36014 17774 36066
rect 17826 36014 17840 36066
rect 17760 36000 17840 36014
rect 17920 36066 18000 36080
rect 17920 36014 17934 36066
rect 17986 36014 18000 36066
rect 17920 36000 18000 36014
rect 18080 36066 18160 36080
rect 18080 36014 18094 36066
rect 18146 36014 18160 36066
rect 18080 36000 18160 36014
rect 18240 36066 18320 36080
rect 18240 36014 18254 36066
rect 18306 36014 18320 36066
rect 18240 36000 18320 36014
rect 18400 36066 18480 36080
rect 18400 36014 18414 36066
rect 18466 36014 18480 36066
rect 18400 36000 18480 36014
rect 18560 36066 18640 36080
rect 18560 36014 18574 36066
rect 18626 36014 18640 36066
rect 18560 36000 18640 36014
rect 18720 36066 18800 36080
rect 18720 36014 18734 36066
rect 18786 36014 18800 36066
rect 18720 36000 18800 36014
rect 18880 36066 18960 36080
rect 18880 36014 18894 36066
rect 18946 36014 18960 36066
rect 18880 36000 18960 36014
rect 23120 36066 23200 36080
rect 23120 36014 23134 36066
rect 23186 36014 23200 36066
rect 23120 36000 23200 36014
rect 23280 36066 23360 36080
rect 23280 36014 23294 36066
rect 23346 36014 23360 36066
rect 23280 36000 23360 36014
rect 23440 36066 23520 36080
rect 23440 36014 23454 36066
rect 23506 36014 23520 36066
rect 23440 36000 23520 36014
rect 23600 36066 23680 36080
rect 23600 36014 23614 36066
rect 23666 36014 23680 36066
rect 23600 36000 23680 36014
rect 23760 36066 23840 36080
rect 23760 36014 23774 36066
rect 23826 36014 23840 36066
rect 23760 36000 23840 36014
rect 23920 36066 24000 36080
rect 23920 36014 23934 36066
rect 23986 36014 24000 36066
rect 23920 36000 24000 36014
rect 24080 36066 24160 36080
rect 24080 36014 24094 36066
rect 24146 36014 24160 36066
rect 24080 36000 24160 36014
rect 24240 36066 24320 36080
rect 24240 36014 24254 36066
rect 24306 36014 24320 36066
rect 24240 36000 24320 36014
rect 24400 36066 24480 36080
rect 24400 36014 24414 36066
rect 24466 36014 24480 36066
rect 24400 36000 24480 36014
rect 24560 36066 24640 36080
rect 24560 36014 24574 36066
rect 24626 36014 24640 36066
rect 24560 36000 24640 36014
rect 24720 36066 24800 36080
rect 24720 36014 24734 36066
rect 24786 36014 24800 36066
rect 24720 36000 24800 36014
rect 24880 36066 24960 36080
rect 24880 36014 24894 36066
rect 24946 36014 24960 36066
rect 24880 36000 24960 36014
rect 25040 36066 25120 36080
rect 25040 36014 25054 36066
rect 25106 36014 25120 36066
rect 25040 36000 25120 36014
rect 25200 36066 25280 36080
rect 25200 36014 25214 36066
rect 25266 36014 25280 36066
rect 25200 36000 25280 36014
rect 25360 36066 25440 36080
rect 25360 36014 25374 36066
rect 25426 36014 25440 36066
rect 25360 36000 25440 36014
rect 25520 36066 25600 36080
rect 25520 36014 25534 36066
rect 25586 36014 25600 36066
rect 25520 36000 25600 36014
rect 25680 36066 25760 36080
rect 25680 36014 25694 36066
rect 25746 36014 25760 36066
rect 25680 36000 25760 36014
rect 25840 36066 25920 36080
rect 25840 36014 25854 36066
rect 25906 36014 25920 36066
rect 25840 36000 25920 36014
rect 26000 36066 26080 36080
rect 26000 36014 26014 36066
rect 26066 36014 26080 36066
rect 26000 36000 26080 36014
rect 26160 36066 26240 36080
rect 26160 36014 26174 36066
rect 26226 36014 26240 36066
rect 26160 36000 26240 36014
rect 26320 36066 26400 36080
rect 26320 36014 26334 36066
rect 26386 36014 26400 36066
rect 26320 36000 26400 36014
rect 26480 36066 26560 36080
rect 26480 36014 26494 36066
rect 26546 36014 26560 36066
rect 26480 36000 26560 36014
rect 26640 36066 26720 36080
rect 26640 36014 26654 36066
rect 26706 36014 26720 36066
rect 26640 36000 26720 36014
rect 26800 36066 26880 36080
rect 26800 36014 26814 36066
rect 26866 36014 26880 36066
rect 26800 36000 26880 36014
rect 26960 36066 27040 36080
rect 26960 36014 26974 36066
rect 27026 36014 27040 36066
rect 26960 36000 27040 36014
rect 27120 36066 27200 36080
rect 27120 36014 27134 36066
rect 27186 36014 27200 36066
rect 27120 36000 27200 36014
rect 27280 36066 27360 36080
rect 27280 36014 27294 36066
rect 27346 36014 27360 36066
rect 27280 36000 27360 36014
rect 27440 36066 27520 36080
rect 27440 36014 27454 36066
rect 27506 36014 27520 36066
rect 27440 36000 27520 36014
rect 27600 36066 27680 36080
rect 27600 36014 27614 36066
rect 27666 36014 27680 36066
rect 27600 36000 27680 36014
rect 27760 36066 27840 36080
rect 27760 36014 27774 36066
rect 27826 36014 27840 36066
rect 27760 36000 27840 36014
rect 27920 36066 28000 36080
rect 27920 36014 27934 36066
rect 27986 36014 28000 36066
rect 27920 36000 28000 36014
rect 28080 36066 28160 36080
rect 28080 36014 28094 36066
rect 28146 36014 28160 36066
rect 28080 36000 28160 36014
rect 28240 36066 28320 36080
rect 28240 36014 28254 36066
rect 28306 36014 28320 36066
rect 28240 36000 28320 36014
rect 28400 36066 28480 36080
rect 28400 36014 28414 36066
rect 28466 36014 28480 36066
rect 28400 36000 28480 36014
rect 28560 36066 28640 36080
rect 28560 36014 28574 36066
rect 28626 36014 28640 36066
rect 28560 36000 28640 36014
rect 28720 36066 28800 36080
rect 28720 36014 28734 36066
rect 28786 36014 28800 36066
rect 28720 36000 28800 36014
rect 28880 36066 28960 36080
rect 28880 36014 28894 36066
rect 28946 36014 28960 36066
rect 28880 36000 28960 36014
rect 29040 36066 29120 36080
rect 29040 36014 29054 36066
rect 29106 36014 29120 36066
rect 29040 36000 29120 36014
rect 29200 36066 29280 36080
rect 29200 36014 29214 36066
rect 29266 36014 29280 36066
rect 29200 36000 29280 36014
rect 29360 36066 29440 36080
rect 29360 36014 29374 36066
rect 29426 36014 29440 36066
rect 29360 36000 29440 36014
rect 33520 36066 33600 36080
rect 33520 36014 33534 36066
rect 33586 36014 33600 36066
rect 33520 36000 33600 36014
rect 33680 36066 33760 36080
rect 33680 36014 33694 36066
rect 33746 36014 33760 36066
rect 33680 36000 33760 36014
rect 33840 36066 33920 36080
rect 33840 36014 33854 36066
rect 33906 36014 33920 36066
rect 33840 36000 33920 36014
rect 34000 36066 34080 36080
rect 34000 36014 34014 36066
rect 34066 36014 34080 36066
rect 34000 36000 34080 36014
rect 34160 36066 34240 36080
rect 34160 36014 34174 36066
rect 34226 36014 34240 36066
rect 34160 36000 34240 36014
rect 34320 36066 34400 36080
rect 34320 36014 34334 36066
rect 34386 36014 34400 36066
rect 34320 36000 34400 36014
rect 34480 36066 34560 36080
rect 34480 36014 34494 36066
rect 34546 36014 34560 36066
rect 34480 36000 34560 36014
rect 34640 36066 34720 36080
rect 34640 36014 34654 36066
rect 34706 36014 34720 36066
rect 34640 36000 34720 36014
rect 34800 36066 34880 36080
rect 34800 36014 34814 36066
rect 34866 36014 34880 36066
rect 34800 36000 34880 36014
rect 34960 36066 35040 36080
rect 34960 36014 34974 36066
rect 35026 36014 35040 36066
rect 34960 36000 35040 36014
rect 35120 36066 35200 36080
rect 35120 36014 35134 36066
rect 35186 36014 35200 36066
rect 35120 36000 35200 36014
rect 35280 36066 35360 36080
rect 35280 36014 35294 36066
rect 35346 36014 35360 36066
rect 35280 36000 35360 36014
rect 35440 36066 35520 36080
rect 35440 36014 35454 36066
rect 35506 36014 35520 36066
rect 35440 36000 35520 36014
rect 35600 36066 35680 36080
rect 35600 36014 35614 36066
rect 35666 36014 35680 36066
rect 35600 36000 35680 36014
rect 35760 36066 35840 36080
rect 35760 36014 35774 36066
rect 35826 36014 35840 36066
rect 35760 36000 35840 36014
rect 35920 36066 36000 36080
rect 35920 36014 35934 36066
rect 35986 36014 36000 36066
rect 35920 36000 36000 36014
rect 36080 36066 36160 36080
rect 36080 36014 36094 36066
rect 36146 36014 36160 36066
rect 36080 36000 36160 36014
rect 36240 36066 36320 36080
rect 36240 36014 36254 36066
rect 36306 36014 36320 36066
rect 36240 36000 36320 36014
rect 36400 36066 36480 36080
rect 36400 36014 36414 36066
rect 36466 36014 36480 36066
rect 36400 36000 36480 36014
rect 36560 36066 36640 36080
rect 36560 36014 36574 36066
rect 36626 36014 36640 36066
rect 36560 36000 36640 36014
rect 36720 36066 36800 36080
rect 36720 36014 36734 36066
rect 36786 36014 36800 36066
rect 36720 36000 36800 36014
rect 36880 36066 36960 36080
rect 36880 36014 36894 36066
rect 36946 36014 36960 36066
rect 36880 36000 36960 36014
rect 37040 36066 37120 36080
rect 37040 36014 37054 36066
rect 37106 36014 37120 36066
rect 37040 36000 37120 36014
rect 37200 36066 37280 36080
rect 37200 36014 37214 36066
rect 37266 36014 37280 36066
rect 37200 36000 37280 36014
rect 37360 36066 37440 36080
rect 37360 36014 37374 36066
rect 37426 36014 37440 36066
rect 37360 36000 37440 36014
rect 37520 36066 37600 36080
rect 37520 36014 37534 36066
rect 37586 36014 37600 36066
rect 37520 36000 37600 36014
rect 37680 36066 37760 36080
rect 37680 36014 37694 36066
rect 37746 36014 37760 36066
rect 37680 36000 37760 36014
rect 37840 36066 37920 36080
rect 37840 36014 37854 36066
rect 37906 36014 37920 36066
rect 37840 36000 37920 36014
rect 38000 36066 38080 36080
rect 38000 36014 38014 36066
rect 38066 36014 38080 36066
rect 38000 36000 38080 36014
rect 38160 36066 38240 36080
rect 38160 36014 38174 36066
rect 38226 36014 38240 36066
rect 38160 36000 38240 36014
rect 38320 36066 38400 36080
rect 38320 36014 38334 36066
rect 38386 36014 38400 36066
rect 38320 36000 38400 36014
rect 38480 36066 38560 36080
rect 38480 36014 38494 36066
rect 38546 36014 38560 36066
rect 38480 36000 38560 36014
rect 38640 36066 38720 36080
rect 38640 36014 38654 36066
rect 38706 36014 38720 36066
rect 38640 36000 38720 36014
rect 38800 36066 38880 36080
rect 38800 36014 38814 36066
rect 38866 36014 38880 36066
rect 38800 36000 38880 36014
rect 38960 36066 39040 36080
rect 38960 36014 38974 36066
rect 39026 36014 39040 36066
rect 38960 36000 39040 36014
rect 39120 36066 39200 36080
rect 39120 36014 39134 36066
rect 39186 36014 39200 36066
rect 39120 36000 39200 36014
rect 39280 36066 39360 36080
rect 39280 36014 39294 36066
rect 39346 36014 39360 36066
rect 39280 36000 39360 36014
rect 39440 36066 39520 36080
rect 39440 36014 39454 36066
rect 39506 36014 39520 36066
rect 39440 36000 39520 36014
rect 39600 36066 39680 36080
rect 39600 36014 39614 36066
rect 39666 36014 39680 36066
rect 39600 36000 39680 36014
rect 39760 36066 39840 36080
rect 39760 36014 39774 36066
rect 39826 36014 39840 36066
rect 39760 36000 39840 36014
rect 39920 36066 40000 36080
rect 39920 36014 39934 36066
rect 39986 36014 40000 36066
rect 39920 36000 40000 36014
rect 40080 36066 40160 36080
rect 40080 36014 40094 36066
rect 40146 36014 40160 36066
rect 40080 36000 40160 36014
rect 40240 36066 40320 36080
rect 40240 36014 40254 36066
rect 40306 36014 40320 36066
rect 40240 36000 40320 36014
rect 40400 36066 40480 36080
rect 40400 36014 40414 36066
rect 40466 36014 40480 36066
rect 40400 36000 40480 36014
rect 40560 36066 40640 36080
rect 40560 36014 40574 36066
rect 40626 36014 40640 36066
rect 40560 36000 40640 36014
rect 40720 36066 40800 36080
rect 40720 36014 40734 36066
rect 40786 36014 40800 36066
rect 40720 36000 40800 36014
rect 40880 36066 40960 36080
rect 40880 36014 40894 36066
rect 40946 36014 40960 36066
rect 40880 36000 40960 36014
rect 41040 36066 41120 36080
rect 41040 36014 41054 36066
rect 41106 36014 41120 36066
rect 41040 36000 41120 36014
rect 41200 36066 41280 36080
rect 41200 36014 41214 36066
rect 41266 36014 41280 36066
rect 41200 36000 41280 36014
rect 41360 36066 41440 36080
rect 41360 36014 41374 36066
rect 41426 36014 41440 36066
rect 41360 36000 41440 36014
rect 41520 36066 41600 36080
rect 41520 36014 41534 36066
rect 41586 36014 41600 36066
rect 41520 36000 41600 36014
rect 41680 36066 41760 36080
rect 41680 36014 41694 36066
rect 41746 36014 41760 36066
rect 41680 36000 41760 36014
rect 41840 36066 41920 36080
rect 41840 36014 41854 36066
rect 41906 36014 41920 36066
rect 41840 36000 41920 36014
rect 0 35746 80 35760
rect 0 35694 14 35746
rect 66 35694 80 35746
rect 0 35680 80 35694
rect 160 35746 240 35760
rect 160 35694 174 35746
rect 226 35694 240 35746
rect 160 35680 240 35694
rect 320 35746 400 35760
rect 320 35694 334 35746
rect 386 35694 400 35746
rect 320 35680 400 35694
rect 480 35746 560 35760
rect 480 35694 494 35746
rect 546 35694 560 35746
rect 480 35680 560 35694
rect 640 35746 720 35760
rect 640 35694 654 35746
rect 706 35694 720 35746
rect 640 35680 720 35694
rect 800 35746 880 35760
rect 800 35694 814 35746
rect 866 35694 880 35746
rect 800 35680 880 35694
rect 960 35746 1040 35760
rect 960 35694 974 35746
rect 1026 35694 1040 35746
rect 960 35680 1040 35694
rect 1120 35746 1200 35760
rect 1120 35694 1134 35746
rect 1186 35694 1200 35746
rect 1120 35680 1200 35694
rect 1280 35746 1360 35760
rect 1280 35694 1294 35746
rect 1346 35694 1360 35746
rect 1280 35680 1360 35694
rect 1440 35746 1520 35760
rect 1440 35694 1454 35746
rect 1506 35694 1520 35746
rect 1440 35680 1520 35694
rect 1600 35746 1680 35760
rect 1600 35694 1614 35746
rect 1666 35694 1680 35746
rect 1600 35680 1680 35694
rect 1760 35746 1840 35760
rect 1760 35694 1774 35746
rect 1826 35694 1840 35746
rect 1760 35680 1840 35694
rect 1920 35746 2000 35760
rect 1920 35694 1934 35746
rect 1986 35694 2000 35746
rect 1920 35680 2000 35694
rect 2080 35746 2160 35760
rect 2080 35694 2094 35746
rect 2146 35694 2160 35746
rect 2080 35680 2160 35694
rect 2240 35746 2320 35760
rect 2240 35694 2254 35746
rect 2306 35694 2320 35746
rect 2240 35680 2320 35694
rect 2400 35746 2480 35760
rect 2400 35694 2414 35746
rect 2466 35694 2480 35746
rect 2400 35680 2480 35694
rect 2560 35746 2640 35760
rect 2560 35694 2574 35746
rect 2626 35694 2640 35746
rect 2560 35680 2640 35694
rect 2720 35746 2800 35760
rect 2720 35694 2734 35746
rect 2786 35694 2800 35746
rect 2720 35680 2800 35694
rect 2880 35746 2960 35760
rect 2880 35694 2894 35746
rect 2946 35694 2960 35746
rect 2880 35680 2960 35694
rect 3040 35746 3120 35760
rect 3040 35694 3054 35746
rect 3106 35694 3120 35746
rect 3040 35680 3120 35694
rect 3200 35746 3280 35760
rect 3200 35694 3214 35746
rect 3266 35694 3280 35746
rect 3200 35680 3280 35694
rect 3360 35746 3440 35760
rect 3360 35694 3374 35746
rect 3426 35694 3440 35746
rect 3360 35680 3440 35694
rect 3520 35746 3600 35760
rect 3520 35694 3534 35746
rect 3586 35694 3600 35746
rect 3520 35680 3600 35694
rect 3680 35746 3760 35760
rect 3680 35694 3694 35746
rect 3746 35694 3760 35746
rect 3680 35680 3760 35694
rect 3840 35746 3920 35760
rect 3840 35694 3854 35746
rect 3906 35694 3920 35746
rect 3840 35680 3920 35694
rect 4000 35746 4080 35760
rect 4000 35694 4014 35746
rect 4066 35694 4080 35746
rect 4000 35680 4080 35694
rect 4160 35746 4240 35760
rect 4160 35694 4174 35746
rect 4226 35694 4240 35746
rect 4160 35680 4240 35694
rect 4320 35746 4400 35760
rect 4320 35694 4334 35746
rect 4386 35694 4400 35746
rect 4320 35680 4400 35694
rect 4480 35746 4560 35760
rect 4480 35694 4494 35746
rect 4546 35694 4560 35746
rect 4480 35680 4560 35694
rect 4640 35746 4720 35760
rect 4640 35694 4654 35746
rect 4706 35694 4720 35746
rect 4640 35680 4720 35694
rect 4800 35746 4880 35760
rect 4800 35694 4814 35746
rect 4866 35694 4880 35746
rect 4800 35680 4880 35694
rect 4960 35746 5040 35760
rect 4960 35694 4974 35746
rect 5026 35694 5040 35746
rect 4960 35680 5040 35694
rect 5120 35746 5200 35760
rect 5120 35694 5134 35746
rect 5186 35694 5200 35746
rect 5120 35680 5200 35694
rect 5280 35746 5360 35760
rect 5280 35694 5294 35746
rect 5346 35694 5360 35746
rect 5280 35680 5360 35694
rect 5440 35746 5520 35760
rect 5440 35694 5454 35746
rect 5506 35694 5520 35746
rect 5440 35680 5520 35694
rect 5600 35746 5680 35760
rect 5600 35694 5614 35746
rect 5666 35694 5680 35746
rect 5600 35680 5680 35694
rect 5760 35746 5840 35760
rect 5760 35694 5774 35746
rect 5826 35694 5840 35746
rect 5760 35680 5840 35694
rect 5920 35746 6000 35760
rect 5920 35694 5934 35746
rect 5986 35694 6000 35746
rect 5920 35680 6000 35694
rect 6080 35746 6160 35760
rect 6080 35694 6094 35746
rect 6146 35694 6160 35746
rect 6080 35680 6160 35694
rect 6240 35746 6320 35760
rect 6240 35694 6254 35746
rect 6306 35694 6320 35746
rect 6240 35680 6320 35694
rect 6400 35746 6480 35760
rect 6400 35694 6414 35746
rect 6466 35694 6480 35746
rect 6400 35680 6480 35694
rect 6560 35746 6640 35760
rect 6560 35694 6574 35746
rect 6626 35694 6640 35746
rect 6560 35680 6640 35694
rect 6720 35746 6800 35760
rect 6720 35694 6734 35746
rect 6786 35694 6800 35746
rect 6720 35680 6800 35694
rect 6880 35746 6960 35760
rect 6880 35694 6894 35746
rect 6946 35694 6960 35746
rect 6880 35680 6960 35694
rect 7040 35746 7120 35760
rect 7040 35694 7054 35746
rect 7106 35694 7120 35746
rect 7040 35680 7120 35694
rect 7200 35746 7280 35760
rect 7200 35694 7214 35746
rect 7266 35694 7280 35746
rect 7200 35680 7280 35694
rect 7360 35746 7440 35760
rect 7360 35694 7374 35746
rect 7426 35694 7440 35746
rect 7360 35680 7440 35694
rect 7520 35746 7600 35760
rect 7520 35694 7534 35746
rect 7586 35694 7600 35746
rect 7520 35680 7600 35694
rect 7680 35746 7760 35760
rect 7680 35694 7694 35746
rect 7746 35694 7760 35746
rect 7680 35680 7760 35694
rect 7840 35746 7920 35760
rect 7840 35694 7854 35746
rect 7906 35694 7920 35746
rect 7840 35680 7920 35694
rect 8000 35746 8080 35760
rect 8000 35694 8014 35746
rect 8066 35694 8080 35746
rect 8000 35680 8080 35694
rect 8160 35746 8240 35760
rect 8160 35694 8174 35746
rect 8226 35694 8240 35746
rect 8160 35680 8240 35694
rect 8320 35746 8400 35760
rect 8320 35694 8334 35746
rect 8386 35694 8400 35746
rect 8320 35680 8400 35694
rect 12480 35746 12560 35760
rect 12480 35694 12494 35746
rect 12546 35694 12560 35746
rect 12480 35680 12560 35694
rect 12640 35746 12720 35760
rect 12640 35694 12654 35746
rect 12706 35694 12720 35746
rect 12640 35680 12720 35694
rect 12800 35746 12880 35760
rect 12800 35694 12814 35746
rect 12866 35694 12880 35746
rect 12800 35680 12880 35694
rect 12960 35746 13040 35760
rect 12960 35694 12974 35746
rect 13026 35694 13040 35746
rect 12960 35680 13040 35694
rect 13120 35746 13200 35760
rect 13120 35694 13134 35746
rect 13186 35694 13200 35746
rect 13120 35680 13200 35694
rect 13280 35746 13360 35760
rect 13280 35694 13294 35746
rect 13346 35694 13360 35746
rect 13280 35680 13360 35694
rect 13440 35746 13520 35760
rect 13440 35694 13454 35746
rect 13506 35694 13520 35746
rect 13440 35680 13520 35694
rect 13600 35746 13680 35760
rect 13600 35694 13614 35746
rect 13666 35694 13680 35746
rect 13600 35680 13680 35694
rect 13760 35746 13840 35760
rect 13760 35694 13774 35746
rect 13826 35694 13840 35746
rect 13760 35680 13840 35694
rect 13920 35746 14000 35760
rect 13920 35694 13934 35746
rect 13986 35694 14000 35746
rect 13920 35680 14000 35694
rect 14080 35746 14160 35760
rect 14080 35694 14094 35746
rect 14146 35694 14160 35746
rect 14080 35680 14160 35694
rect 14240 35746 14320 35760
rect 14240 35694 14254 35746
rect 14306 35694 14320 35746
rect 14240 35680 14320 35694
rect 14400 35746 14480 35760
rect 14400 35694 14414 35746
rect 14466 35694 14480 35746
rect 14400 35680 14480 35694
rect 14560 35746 14640 35760
rect 14560 35694 14574 35746
rect 14626 35694 14640 35746
rect 14560 35680 14640 35694
rect 14720 35746 14800 35760
rect 14720 35694 14734 35746
rect 14786 35694 14800 35746
rect 14720 35680 14800 35694
rect 14880 35746 14960 35760
rect 14880 35694 14894 35746
rect 14946 35694 14960 35746
rect 14880 35680 14960 35694
rect 15040 35746 15120 35760
rect 15040 35694 15054 35746
rect 15106 35694 15120 35746
rect 15040 35680 15120 35694
rect 15200 35746 15280 35760
rect 15200 35694 15214 35746
rect 15266 35694 15280 35746
rect 15200 35680 15280 35694
rect 15360 35746 15440 35760
rect 15360 35694 15374 35746
rect 15426 35694 15440 35746
rect 15360 35680 15440 35694
rect 15520 35746 15600 35760
rect 15520 35694 15534 35746
rect 15586 35694 15600 35746
rect 15520 35680 15600 35694
rect 15680 35746 15760 35760
rect 15680 35694 15694 35746
rect 15746 35694 15760 35746
rect 15680 35680 15760 35694
rect 15840 35746 15920 35760
rect 15840 35694 15854 35746
rect 15906 35694 15920 35746
rect 15840 35680 15920 35694
rect 16000 35746 16080 35760
rect 16000 35694 16014 35746
rect 16066 35694 16080 35746
rect 16000 35680 16080 35694
rect 16160 35746 16240 35760
rect 16160 35694 16174 35746
rect 16226 35694 16240 35746
rect 16160 35680 16240 35694
rect 16320 35746 16400 35760
rect 16320 35694 16334 35746
rect 16386 35694 16400 35746
rect 16320 35680 16400 35694
rect 16480 35746 16560 35760
rect 16480 35694 16494 35746
rect 16546 35694 16560 35746
rect 16480 35680 16560 35694
rect 16640 35746 16720 35760
rect 16640 35694 16654 35746
rect 16706 35694 16720 35746
rect 16640 35680 16720 35694
rect 16800 35746 16880 35760
rect 16800 35694 16814 35746
rect 16866 35694 16880 35746
rect 16800 35680 16880 35694
rect 16960 35746 17040 35760
rect 16960 35694 16974 35746
rect 17026 35694 17040 35746
rect 16960 35680 17040 35694
rect 17120 35746 17200 35760
rect 17120 35694 17134 35746
rect 17186 35694 17200 35746
rect 17120 35680 17200 35694
rect 17280 35746 17360 35760
rect 17280 35694 17294 35746
rect 17346 35694 17360 35746
rect 17280 35680 17360 35694
rect 17440 35746 17520 35760
rect 17440 35694 17454 35746
rect 17506 35694 17520 35746
rect 17440 35680 17520 35694
rect 17600 35746 17680 35760
rect 17600 35694 17614 35746
rect 17666 35694 17680 35746
rect 17600 35680 17680 35694
rect 17760 35746 17840 35760
rect 17760 35694 17774 35746
rect 17826 35694 17840 35746
rect 17760 35680 17840 35694
rect 17920 35746 18000 35760
rect 17920 35694 17934 35746
rect 17986 35694 18000 35746
rect 17920 35680 18000 35694
rect 18080 35746 18160 35760
rect 18080 35694 18094 35746
rect 18146 35694 18160 35746
rect 18080 35680 18160 35694
rect 18240 35746 18320 35760
rect 18240 35694 18254 35746
rect 18306 35694 18320 35746
rect 18240 35680 18320 35694
rect 18400 35746 18480 35760
rect 18400 35694 18414 35746
rect 18466 35694 18480 35746
rect 18400 35680 18480 35694
rect 18560 35746 18640 35760
rect 18560 35694 18574 35746
rect 18626 35694 18640 35746
rect 18560 35680 18640 35694
rect 18720 35746 18800 35760
rect 18720 35694 18734 35746
rect 18786 35694 18800 35746
rect 18720 35680 18800 35694
rect 18880 35746 18960 35760
rect 18880 35694 18894 35746
rect 18946 35694 18960 35746
rect 18880 35680 18960 35694
rect 23120 35746 23200 35760
rect 23120 35694 23134 35746
rect 23186 35694 23200 35746
rect 23120 35680 23200 35694
rect 23280 35746 23360 35760
rect 23280 35694 23294 35746
rect 23346 35694 23360 35746
rect 23280 35680 23360 35694
rect 23440 35746 23520 35760
rect 23440 35694 23454 35746
rect 23506 35694 23520 35746
rect 23440 35680 23520 35694
rect 23600 35746 23680 35760
rect 23600 35694 23614 35746
rect 23666 35694 23680 35746
rect 23600 35680 23680 35694
rect 23760 35746 23840 35760
rect 23760 35694 23774 35746
rect 23826 35694 23840 35746
rect 23760 35680 23840 35694
rect 23920 35746 24000 35760
rect 23920 35694 23934 35746
rect 23986 35694 24000 35746
rect 23920 35680 24000 35694
rect 24080 35746 24160 35760
rect 24080 35694 24094 35746
rect 24146 35694 24160 35746
rect 24080 35680 24160 35694
rect 24240 35746 24320 35760
rect 24240 35694 24254 35746
rect 24306 35694 24320 35746
rect 24240 35680 24320 35694
rect 24400 35746 24480 35760
rect 24400 35694 24414 35746
rect 24466 35694 24480 35746
rect 24400 35680 24480 35694
rect 24560 35746 24640 35760
rect 24560 35694 24574 35746
rect 24626 35694 24640 35746
rect 24560 35680 24640 35694
rect 24720 35746 24800 35760
rect 24720 35694 24734 35746
rect 24786 35694 24800 35746
rect 24720 35680 24800 35694
rect 24880 35746 24960 35760
rect 24880 35694 24894 35746
rect 24946 35694 24960 35746
rect 24880 35680 24960 35694
rect 25040 35746 25120 35760
rect 25040 35694 25054 35746
rect 25106 35694 25120 35746
rect 25040 35680 25120 35694
rect 25200 35746 25280 35760
rect 25200 35694 25214 35746
rect 25266 35694 25280 35746
rect 25200 35680 25280 35694
rect 25360 35746 25440 35760
rect 25360 35694 25374 35746
rect 25426 35694 25440 35746
rect 25360 35680 25440 35694
rect 25520 35746 25600 35760
rect 25520 35694 25534 35746
rect 25586 35694 25600 35746
rect 25520 35680 25600 35694
rect 25680 35746 25760 35760
rect 25680 35694 25694 35746
rect 25746 35694 25760 35746
rect 25680 35680 25760 35694
rect 25840 35746 25920 35760
rect 25840 35694 25854 35746
rect 25906 35694 25920 35746
rect 25840 35680 25920 35694
rect 26000 35746 26080 35760
rect 26000 35694 26014 35746
rect 26066 35694 26080 35746
rect 26000 35680 26080 35694
rect 26160 35746 26240 35760
rect 26160 35694 26174 35746
rect 26226 35694 26240 35746
rect 26160 35680 26240 35694
rect 26320 35746 26400 35760
rect 26320 35694 26334 35746
rect 26386 35694 26400 35746
rect 26320 35680 26400 35694
rect 26480 35746 26560 35760
rect 26480 35694 26494 35746
rect 26546 35694 26560 35746
rect 26480 35680 26560 35694
rect 26640 35746 26720 35760
rect 26640 35694 26654 35746
rect 26706 35694 26720 35746
rect 26640 35680 26720 35694
rect 26800 35746 26880 35760
rect 26800 35694 26814 35746
rect 26866 35694 26880 35746
rect 26800 35680 26880 35694
rect 26960 35746 27040 35760
rect 26960 35694 26974 35746
rect 27026 35694 27040 35746
rect 26960 35680 27040 35694
rect 27120 35746 27200 35760
rect 27120 35694 27134 35746
rect 27186 35694 27200 35746
rect 27120 35680 27200 35694
rect 27280 35746 27360 35760
rect 27280 35694 27294 35746
rect 27346 35694 27360 35746
rect 27280 35680 27360 35694
rect 27440 35746 27520 35760
rect 27440 35694 27454 35746
rect 27506 35694 27520 35746
rect 27440 35680 27520 35694
rect 27600 35746 27680 35760
rect 27600 35694 27614 35746
rect 27666 35694 27680 35746
rect 27600 35680 27680 35694
rect 27760 35746 27840 35760
rect 27760 35694 27774 35746
rect 27826 35694 27840 35746
rect 27760 35680 27840 35694
rect 27920 35746 28000 35760
rect 27920 35694 27934 35746
rect 27986 35694 28000 35746
rect 27920 35680 28000 35694
rect 28080 35746 28160 35760
rect 28080 35694 28094 35746
rect 28146 35694 28160 35746
rect 28080 35680 28160 35694
rect 28240 35746 28320 35760
rect 28240 35694 28254 35746
rect 28306 35694 28320 35746
rect 28240 35680 28320 35694
rect 28400 35746 28480 35760
rect 28400 35694 28414 35746
rect 28466 35694 28480 35746
rect 28400 35680 28480 35694
rect 28560 35746 28640 35760
rect 28560 35694 28574 35746
rect 28626 35694 28640 35746
rect 28560 35680 28640 35694
rect 28720 35746 28800 35760
rect 28720 35694 28734 35746
rect 28786 35694 28800 35746
rect 28720 35680 28800 35694
rect 28880 35746 28960 35760
rect 28880 35694 28894 35746
rect 28946 35694 28960 35746
rect 28880 35680 28960 35694
rect 29040 35746 29120 35760
rect 29040 35694 29054 35746
rect 29106 35694 29120 35746
rect 29040 35680 29120 35694
rect 29200 35746 29280 35760
rect 29200 35694 29214 35746
rect 29266 35694 29280 35746
rect 29200 35680 29280 35694
rect 29360 35746 29440 35760
rect 29360 35694 29374 35746
rect 29426 35694 29440 35746
rect 29360 35680 29440 35694
rect 33520 35746 33600 35760
rect 33520 35694 33534 35746
rect 33586 35694 33600 35746
rect 33520 35680 33600 35694
rect 33680 35746 33760 35760
rect 33680 35694 33694 35746
rect 33746 35694 33760 35746
rect 33680 35680 33760 35694
rect 33840 35746 33920 35760
rect 33840 35694 33854 35746
rect 33906 35694 33920 35746
rect 33840 35680 33920 35694
rect 34000 35746 34080 35760
rect 34000 35694 34014 35746
rect 34066 35694 34080 35746
rect 34000 35680 34080 35694
rect 34160 35746 34240 35760
rect 34160 35694 34174 35746
rect 34226 35694 34240 35746
rect 34160 35680 34240 35694
rect 34320 35746 34400 35760
rect 34320 35694 34334 35746
rect 34386 35694 34400 35746
rect 34320 35680 34400 35694
rect 34480 35746 34560 35760
rect 34480 35694 34494 35746
rect 34546 35694 34560 35746
rect 34480 35680 34560 35694
rect 34640 35746 34720 35760
rect 34640 35694 34654 35746
rect 34706 35694 34720 35746
rect 34640 35680 34720 35694
rect 34800 35746 34880 35760
rect 34800 35694 34814 35746
rect 34866 35694 34880 35746
rect 34800 35680 34880 35694
rect 34960 35746 35040 35760
rect 34960 35694 34974 35746
rect 35026 35694 35040 35746
rect 34960 35680 35040 35694
rect 35120 35746 35200 35760
rect 35120 35694 35134 35746
rect 35186 35694 35200 35746
rect 35120 35680 35200 35694
rect 35280 35746 35360 35760
rect 35280 35694 35294 35746
rect 35346 35694 35360 35746
rect 35280 35680 35360 35694
rect 35440 35746 35520 35760
rect 35440 35694 35454 35746
rect 35506 35694 35520 35746
rect 35440 35680 35520 35694
rect 35600 35746 35680 35760
rect 35600 35694 35614 35746
rect 35666 35694 35680 35746
rect 35600 35680 35680 35694
rect 35760 35746 35840 35760
rect 35760 35694 35774 35746
rect 35826 35694 35840 35746
rect 35760 35680 35840 35694
rect 35920 35746 36000 35760
rect 35920 35694 35934 35746
rect 35986 35694 36000 35746
rect 35920 35680 36000 35694
rect 36080 35746 36160 35760
rect 36080 35694 36094 35746
rect 36146 35694 36160 35746
rect 36080 35680 36160 35694
rect 36240 35746 36320 35760
rect 36240 35694 36254 35746
rect 36306 35694 36320 35746
rect 36240 35680 36320 35694
rect 36400 35746 36480 35760
rect 36400 35694 36414 35746
rect 36466 35694 36480 35746
rect 36400 35680 36480 35694
rect 36560 35746 36640 35760
rect 36560 35694 36574 35746
rect 36626 35694 36640 35746
rect 36560 35680 36640 35694
rect 36720 35746 36800 35760
rect 36720 35694 36734 35746
rect 36786 35694 36800 35746
rect 36720 35680 36800 35694
rect 36880 35746 36960 35760
rect 36880 35694 36894 35746
rect 36946 35694 36960 35746
rect 36880 35680 36960 35694
rect 37040 35746 37120 35760
rect 37040 35694 37054 35746
rect 37106 35694 37120 35746
rect 37040 35680 37120 35694
rect 37200 35746 37280 35760
rect 37200 35694 37214 35746
rect 37266 35694 37280 35746
rect 37200 35680 37280 35694
rect 37360 35746 37440 35760
rect 37360 35694 37374 35746
rect 37426 35694 37440 35746
rect 37360 35680 37440 35694
rect 37520 35746 37600 35760
rect 37520 35694 37534 35746
rect 37586 35694 37600 35746
rect 37520 35680 37600 35694
rect 37680 35746 37760 35760
rect 37680 35694 37694 35746
rect 37746 35694 37760 35746
rect 37680 35680 37760 35694
rect 37840 35746 37920 35760
rect 37840 35694 37854 35746
rect 37906 35694 37920 35746
rect 37840 35680 37920 35694
rect 38000 35746 38080 35760
rect 38000 35694 38014 35746
rect 38066 35694 38080 35746
rect 38000 35680 38080 35694
rect 38160 35746 38240 35760
rect 38160 35694 38174 35746
rect 38226 35694 38240 35746
rect 38160 35680 38240 35694
rect 38320 35746 38400 35760
rect 38320 35694 38334 35746
rect 38386 35694 38400 35746
rect 38320 35680 38400 35694
rect 38480 35746 38560 35760
rect 38480 35694 38494 35746
rect 38546 35694 38560 35746
rect 38480 35680 38560 35694
rect 38640 35746 38720 35760
rect 38640 35694 38654 35746
rect 38706 35694 38720 35746
rect 38640 35680 38720 35694
rect 38800 35746 38880 35760
rect 38800 35694 38814 35746
rect 38866 35694 38880 35746
rect 38800 35680 38880 35694
rect 38960 35746 39040 35760
rect 38960 35694 38974 35746
rect 39026 35694 39040 35746
rect 38960 35680 39040 35694
rect 39120 35746 39200 35760
rect 39120 35694 39134 35746
rect 39186 35694 39200 35746
rect 39120 35680 39200 35694
rect 39280 35746 39360 35760
rect 39280 35694 39294 35746
rect 39346 35694 39360 35746
rect 39280 35680 39360 35694
rect 39440 35746 39520 35760
rect 39440 35694 39454 35746
rect 39506 35694 39520 35746
rect 39440 35680 39520 35694
rect 39600 35746 39680 35760
rect 39600 35694 39614 35746
rect 39666 35694 39680 35746
rect 39600 35680 39680 35694
rect 39760 35746 39840 35760
rect 39760 35694 39774 35746
rect 39826 35694 39840 35746
rect 39760 35680 39840 35694
rect 39920 35746 40000 35760
rect 39920 35694 39934 35746
rect 39986 35694 40000 35746
rect 39920 35680 40000 35694
rect 40080 35746 40160 35760
rect 40080 35694 40094 35746
rect 40146 35694 40160 35746
rect 40080 35680 40160 35694
rect 40240 35746 40320 35760
rect 40240 35694 40254 35746
rect 40306 35694 40320 35746
rect 40240 35680 40320 35694
rect 40400 35746 40480 35760
rect 40400 35694 40414 35746
rect 40466 35694 40480 35746
rect 40400 35680 40480 35694
rect 40560 35746 40640 35760
rect 40560 35694 40574 35746
rect 40626 35694 40640 35746
rect 40560 35680 40640 35694
rect 40720 35746 40800 35760
rect 40720 35694 40734 35746
rect 40786 35694 40800 35746
rect 40720 35680 40800 35694
rect 40880 35746 40960 35760
rect 40880 35694 40894 35746
rect 40946 35694 40960 35746
rect 40880 35680 40960 35694
rect 41040 35746 41120 35760
rect 41040 35694 41054 35746
rect 41106 35694 41120 35746
rect 41040 35680 41120 35694
rect 41200 35746 41280 35760
rect 41200 35694 41214 35746
rect 41266 35694 41280 35746
rect 41200 35680 41280 35694
rect 41360 35746 41440 35760
rect 41360 35694 41374 35746
rect 41426 35694 41440 35746
rect 41360 35680 41440 35694
rect 41520 35746 41600 35760
rect 41520 35694 41534 35746
rect 41586 35694 41600 35746
rect 41520 35680 41600 35694
rect 41680 35746 41760 35760
rect 41680 35694 41694 35746
rect 41746 35694 41760 35746
rect 41680 35680 41760 35694
rect 41840 35746 41920 35760
rect 41840 35694 41854 35746
rect 41906 35694 41920 35746
rect 41840 35680 41920 35694
rect 0 35426 80 35440
rect 0 35374 14 35426
rect 66 35374 80 35426
rect 0 35360 80 35374
rect 160 35426 240 35440
rect 160 35374 174 35426
rect 226 35374 240 35426
rect 160 35360 240 35374
rect 320 35426 400 35440
rect 320 35374 334 35426
rect 386 35374 400 35426
rect 320 35360 400 35374
rect 480 35426 560 35440
rect 480 35374 494 35426
rect 546 35374 560 35426
rect 480 35360 560 35374
rect 640 35426 720 35440
rect 640 35374 654 35426
rect 706 35374 720 35426
rect 640 35360 720 35374
rect 800 35426 880 35440
rect 800 35374 814 35426
rect 866 35374 880 35426
rect 800 35360 880 35374
rect 960 35426 1040 35440
rect 960 35374 974 35426
rect 1026 35374 1040 35426
rect 960 35360 1040 35374
rect 1120 35426 1200 35440
rect 1120 35374 1134 35426
rect 1186 35374 1200 35426
rect 1120 35360 1200 35374
rect 1280 35426 1360 35440
rect 1280 35374 1294 35426
rect 1346 35374 1360 35426
rect 1280 35360 1360 35374
rect 1440 35426 1520 35440
rect 1440 35374 1454 35426
rect 1506 35374 1520 35426
rect 1440 35360 1520 35374
rect 1600 35426 1680 35440
rect 1600 35374 1614 35426
rect 1666 35374 1680 35426
rect 1600 35360 1680 35374
rect 1760 35426 1840 35440
rect 1760 35374 1774 35426
rect 1826 35374 1840 35426
rect 1760 35360 1840 35374
rect 1920 35426 2000 35440
rect 1920 35374 1934 35426
rect 1986 35374 2000 35426
rect 1920 35360 2000 35374
rect 2080 35426 2160 35440
rect 2080 35374 2094 35426
rect 2146 35374 2160 35426
rect 2080 35360 2160 35374
rect 2240 35426 2320 35440
rect 2240 35374 2254 35426
rect 2306 35374 2320 35426
rect 2240 35360 2320 35374
rect 2400 35426 2480 35440
rect 2400 35374 2414 35426
rect 2466 35374 2480 35426
rect 2400 35360 2480 35374
rect 2560 35426 2640 35440
rect 2560 35374 2574 35426
rect 2626 35374 2640 35426
rect 2560 35360 2640 35374
rect 2720 35426 2800 35440
rect 2720 35374 2734 35426
rect 2786 35374 2800 35426
rect 2720 35360 2800 35374
rect 2880 35426 2960 35440
rect 2880 35374 2894 35426
rect 2946 35374 2960 35426
rect 2880 35360 2960 35374
rect 3040 35426 3120 35440
rect 3040 35374 3054 35426
rect 3106 35374 3120 35426
rect 3040 35360 3120 35374
rect 3200 35426 3280 35440
rect 3200 35374 3214 35426
rect 3266 35374 3280 35426
rect 3200 35360 3280 35374
rect 3360 35426 3440 35440
rect 3360 35374 3374 35426
rect 3426 35374 3440 35426
rect 3360 35360 3440 35374
rect 3520 35426 3600 35440
rect 3520 35374 3534 35426
rect 3586 35374 3600 35426
rect 3520 35360 3600 35374
rect 3680 35426 3760 35440
rect 3680 35374 3694 35426
rect 3746 35374 3760 35426
rect 3680 35360 3760 35374
rect 3840 35426 3920 35440
rect 3840 35374 3854 35426
rect 3906 35374 3920 35426
rect 3840 35360 3920 35374
rect 4000 35426 4080 35440
rect 4000 35374 4014 35426
rect 4066 35374 4080 35426
rect 4000 35360 4080 35374
rect 4160 35426 4240 35440
rect 4160 35374 4174 35426
rect 4226 35374 4240 35426
rect 4160 35360 4240 35374
rect 4320 35426 4400 35440
rect 4320 35374 4334 35426
rect 4386 35374 4400 35426
rect 4320 35360 4400 35374
rect 4480 35426 4560 35440
rect 4480 35374 4494 35426
rect 4546 35374 4560 35426
rect 4480 35360 4560 35374
rect 4640 35426 4720 35440
rect 4640 35374 4654 35426
rect 4706 35374 4720 35426
rect 4640 35360 4720 35374
rect 4800 35426 4880 35440
rect 4800 35374 4814 35426
rect 4866 35374 4880 35426
rect 4800 35360 4880 35374
rect 4960 35426 5040 35440
rect 4960 35374 4974 35426
rect 5026 35374 5040 35426
rect 4960 35360 5040 35374
rect 5120 35426 5200 35440
rect 5120 35374 5134 35426
rect 5186 35374 5200 35426
rect 5120 35360 5200 35374
rect 5280 35426 5360 35440
rect 5280 35374 5294 35426
rect 5346 35374 5360 35426
rect 5280 35360 5360 35374
rect 5440 35426 5520 35440
rect 5440 35374 5454 35426
rect 5506 35374 5520 35426
rect 5440 35360 5520 35374
rect 5600 35426 5680 35440
rect 5600 35374 5614 35426
rect 5666 35374 5680 35426
rect 5600 35360 5680 35374
rect 5760 35426 5840 35440
rect 5760 35374 5774 35426
rect 5826 35374 5840 35426
rect 5760 35360 5840 35374
rect 5920 35426 6000 35440
rect 5920 35374 5934 35426
rect 5986 35374 6000 35426
rect 5920 35360 6000 35374
rect 6080 35426 6160 35440
rect 6080 35374 6094 35426
rect 6146 35374 6160 35426
rect 6080 35360 6160 35374
rect 6240 35426 6320 35440
rect 6240 35374 6254 35426
rect 6306 35374 6320 35426
rect 6240 35360 6320 35374
rect 6400 35426 6480 35440
rect 6400 35374 6414 35426
rect 6466 35374 6480 35426
rect 6400 35360 6480 35374
rect 6560 35426 6640 35440
rect 6560 35374 6574 35426
rect 6626 35374 6640 35426
rect 6560 35360 6640 35374
rect 6720 35426 6800 35440
rect 6720 35374 6734 35426
rect 6786 35374 6800 35426
rect 6720 35360 6800 35374
rect 6880 35426 6960 35440
rect 6880 35374 6894 35426
rect 6946 35374 6960 35426
rect 6880 35360 6960 35374
rect 7040 35426 7120 35440
rect 7040 35374 7054 35426
rect 7106 35374 7120 35426
rect 7040 35360 7120 35374
rect 7200 35426 7280 35440
rect 7200 35374 7214 35426
rect 7266 35374 7280 35426
rect 7200 35360 7280 35374
rect 7360 35426 7440 35440
rect 7360 35374 7374 35426
rect 7426 35374 7440 35426
rect 7360 35360 7440 35374
rect 7520 35426 7600 35440
rect 7520 35374 7534 35426
rect 7586 35374 7600 35426
rect 7520 35360 7600 35374
rect 7680 35426 7760 35440
rect 7680 35374 7694 35426
rect 7746 35374 7760 35426
rect 7680 35360 7760 35374
rect 7840 35426 7920 35440
rect 7840 35374 7854 35426
rect 7906 35374 7920 35426
rect 7840 35360 7920 35374
rect 8000 35426 8080 35440
rect 8000 35374 8014 35426
rect 8066 35374 8080 35426
rect 8000 35360 8080 35374
rect 8160 35426 8240 35440
rect 8160 35374 8174 35426
rect 8226 35374 8240 35426
rect 8160 35360 8240 35374
rect 8320 35426 8400 35440
rect 8320 35374 8334 35426
rect 8386 35374 8400 35426
rect 8320 35360 8400 35374
rect 12480 35426 12560 35440
rect 12480 35374 12494 35426
rect 12546 35374 12560 35426
rect 12480 35360 12560 35374
rect 12640 35426 12720 35440
rect 12640 35374 12654 35426
rect 12706 35374 12720 35426
rect 12640 35360 12720 35374
rect 12800 35426 12880 35440
rect 12800 35374 12814 35426
rect 12866 35374 12880 35426
rect 12800 35360 12880 35374
rect 12960 35426 13040 35440
rect 12960 35374 12974 35426
rect 13026 35374 13040 35426
rect 12960 35360 13040 35374
rect 13120 35426 13200 35440
rect 13120 35374 13134 35426
rect 13186 35374 13200 35426
rect 13120 35360 13200 35374
rect 13280 35426 13360 35440
rect 13280 35374 13294 35426
rect 13346 35374 13360 35426
rect 13280 35360 13360 35374
rect 13440 35426 13520 35440
rect 13440 35374 13454 35426
rect 13506 35374 13520 35426
rect 13440 35360 13520 35374
rect 13600 35426 13680 35440
rect 13600 35374 13614 35426
rect 13666 35374 13680 35426
rect 13600 35360 13680 35374
rect 13760 35426 13840 35440
rect 13760 35374 13774 35426
rect 13826 35374 13840 35426
rect 13760 35360 13840 35374
rect 13920 35426 14000 35440
rect 13920 35374 13934 35426
rect 13986 35374 14000 35426
rect 13920 35360 14000 35374
rect 14080 35426 14160 35440
rect 14080 35374 14094 35426
rect 14146 35374 14160 35426
rect 14080 35360 14160 35374
rect 14240 35426 14320 35440
rect 14240 35374 14254 35426
rect 14306 35374 14320 35426
rect 14240 35360 14320 35374
rect 14400 35426 14480 35440
rect 14400 35374 14414 35426
rect 14466 35374 14480 35426
rect 14400 35360 14480 35374
rect 14560 35426 14640 35440
rect 14560 35374 14574 35426
rect 14626 35374 14640 35426
rect 14560 35360 14640 35374
rect 14720 35426 14800 35440
rect 14720 35374 14734 35426
rect 14786 35374 14800 35426
rect 14720 35360 14800 35374
rect 14880 35426 14960 35440
rect 14880 35374 14894 35426
rect 14946 35374 14960 35426
rect 14880 35360 14960 35374
rect 15040 35426 15120 35440
rect 15040 35374 15054 35426
rect 15106 35374 15120 35426
rect 15040 35360 15120 35374
rect 15200 35426 15280 35440
rect 15200 35374 15214 35426
rect 15266 35374 15280 35426
rect 15200 35360 15280 35374
rect 15360 35426 15440 35440
rect 15360 35374 15374 35426
rect 15426 35374 15440 35426
rect 15360 35360 15440 35374
rect 15520 35426 15600 35440
rect 15520 35374 15534 35426
rect 15586 35374 15600 35426
rect 15520 35360 15600 35374
rect 15680 35426 15760 35440
rect 15680 35374 15694 35426
rect 15746 35374 15760 35426
rect 15680 35360 15760 35374
rect 15840 35426 15920 35440
rect 15840 35374 15854 35426
rect 15906 35374 15920 35426
rect 15840 35360 15920 35374
rect 16000 35426 16080 35440
rect 16000 35374 16014 35426
rect 16066 35374 16080 35426
rect 16000 35360 16080 35374
rect 16160 35426 16240 35440
rect 16160 35374 16174 35426
rect 16226 35374 16240 35426
rect 16160 35360 16240 35374
rect 16320 35426 16400 35440
rect 16320 35374 16334 35426
rect 16386 35374 16400 35426
rect 16320 35360 16400 35374
rect 16480 35426 16560 35440
rect 16480 35374 16494 35426
rect 16546 35374 16560 35426
rect 16480 35360 16560 35374
rect 16640 35426 16720 35440
rect 16640 35374 16654 35426
rect 16706 35374 16720 35426
rect 16640 35360 16720 35374
rect 16800 35426 16880 35440
rect 16800 35374 16814 35426
rect 16866 35374 16880 35426
rect 16800 35360 16880 35374
rect 16960 35426 17040 35440
rect 16960 35374 16974 35426
rect 17026 35374 17040 35426
rect 16960 35360 17040 35374
rect 17120 35426 17200 35440
rect 17120 35374 17134 35426
rect 17186 35374 17200 35426
rect 17120 35360 17200 35374
rect 17280 35426 17360 35440
rect 17280 35374 17294 35426
rect 17346 35374 17360 35426
rect 17280 35360 17360 35374
rect 17440 35426 17520 35440
rect 17440 35374 17454 35426
rect 17506 35374 17520 35426
rect 17440 35360 17520 35374
rect 17600 35426 17680 35440
rect 17600 35374 17614 35426
rect 17666 35374 17680 35426
rect 17600 35360 17680 35374
rect 17760 35426 17840 35440
rect 17760 35374 17774 35426
rect 17826 35374 17840 35426
rect 17760 35360 17840 35374
rect 17920 35426 18000 35440
rect 17920 35374 17934 35426
rect 17986 35374 18000 35426
rect 17920 35360 18000 35374
rect 18080 35426 18160 35440
rect 18080 35374 18094 35426
rect 18146 35374 18160 35426
rect 18080 35360 18160 35374
rect 18240 35426 18320 35440
rect 18240 35374 18254 35426
rect 18306 35374 18320 35426
rect 18240 35360 18320 35374
rect 18400 35426 18480 35440
rect 18400 35374 18414 35426
rect 18466 35374 18480 35426
rect 18400 35360 18480 35374
rect 18560 35426 18640 35440
rect 18560 35374 18574 35426
rect 18626 35374 18640 35426
rect 18560 35360 18640 35374
rect 18720 35426 18800 35440
rect 18720 35374 18734 35426
rect 18786 35374 18800 35426
rect 18720 35360 18800 35374
rect 18880 35426 18960 35440
rect 18880 35374 18894 35426
rect 18946 35374 18960 35426
rect 18880 35360 18960 35374
rect 23120 35426 23200 35440
rect 23120 35374 23134 35426
rect 23186 35374 23200 35426
rect 23120 35360 23200 35374
rect 23280 35426 23360 35440
rect 23280 35374 23294 35426
rect 23346 35374 23360 35426
rect 23280 35360 23360 35374
rect 23440 35426 23520 35440
rect 23440 35374 23454 35426
rect 23506 35374 23520 35426
rect 23440 35360 23520 35374
rect 23600 35426 23680 35440
rect 23600 35374 23614 35426
rect 23666 35374 23680 35426
rect 23600 35360 23680 35374
rect 23760 35426 23840 35440
rect 23760 35374 23774 35426
rect 23826 35374 23840 35426
rect 23760 35360 23840 35374
rect 23920 35426 24000 35440
rect 23920 35374 23934 35426
rect 23986 35374 24000 35426
rect 23920 35360 24000 35374
rect 24080 35426 24160 35440
rect 24080 35374 24094 35426
rect 24146 35374 24160 35426
rect 24080 35360 24160 35374
rect 24240 35426 24320 35440
rect 24240 35374 24254 35426
rect 24306 35374 24320 35426
rect 24240 35360 24320 35374
rect 24400 35426 24480 35440
rect 24400 35374 24414 35426
rect 24466 35374 24480 35426
rect 24400 35360 24480 35374
rect 24560 35426 24640 35440
rect 24560 35374 24574 35426
rect 24626 35374 24640 35426
rect 24560 35360 24640 35374
rect 24720 35426 24800 35440
rect 24720 35374 24734 35426
rect 24786 35374 24800 35426
rect 24720 35360 24800 35374
rect 24880 35426 24960 35440
rect 24880 35374 24894 35426
rect 24946 35374 24960 35426
rect 24880 35360 24960 35374
rect 25040 35426 25120 35440
rect 25040 35374 25054 35426
rect 25106 35374 25120 35426
rect 25040 35360 25120 35374
rect 25200 35426 25280 35440
rect 25200 35374 25214 35426
rect 25266 35374 25280 35426
rect 25200 35360 25280 35374
rect 25360 35426 25440 35440
rect 25360 35374 25374 35426
rect 25426 35374 25440 35426
rect 25360 35360 25440 35374
rect 25520 35426 25600 35440
rect 25520 35374 25534 35426
rect 25586 35374 25600 35426
rect 25520 35360 25600 35374
rect 25680 35426 25760 35440
rect 25680 35374 25694 35426
rect 25746 35374 25760 35426
rect 25680 35360 25760 35374
rect 25840 35426 25920 35440
rect 25840 35374 25854 35426
rect 25906 35374 25920 35426
rect 25840 35360 25920 35374
rect 26000 35426 26080 35440
rect 26000 35374 26014 35426
rect 26066 35374 26080 35426
rect 26000 35360 26080 35374
rect 26160 35426 26240 35440
rect 26160 35374 26174 35426
rect 26226 35374 26240 35426
rect 26160 35360 26240 35374
rect 26320 35426 26400 35440
rect 26320 35374 26334 35426
rect 26386 35374 26400 35426
rect 26320 35360 26400 35374
rect 26480 35426 26560 35440
rect 26480 35374 26494 35426
rect 26546 35374 26560 35426
rect 26480 35360 26560 35374
rect 26640 35426 26720 35440
rect 26640 35374 26654 35426
rect 26706 35374 26720 35426
rect 26640 35360 26720 35374
rect 26800 35426 26880 35440
rect 26800 35374 26814 35426
rect 26866 35374 26880 35426
rect 26800 35360 26880 35374
rect 26960 35426 27040 35440
rect 26960 35374 26974 35426
rect 27026 35374 27040 35426
rect 26960 35360 27040 35374
rect 27120 35426 27200 35440
rect 27120 35374 27134 35426
rect 27186 35374 27200 35426
rect 27120 35360 27200 35374
rect 27280 35426 27360 35440
rect 27280 35374 27294 35426
rect 27346 35374 27360 35426
rect 27280 35360 27360 35374
rect 27440 35426 27520 35440
rect 27440 35374 27454 35426
rect 27506 35374 27520 35426
rect 27440 35360 27520 35374
rect 27600 35426 27680 35440
rect 27600 35374 27614 35426
rect 27666 35374 27680 35426
rect 27600 35360 27680 35374
rect 27760 35426 27840 35440
rect 27760 35374 27774 35426
rect 27826 35374 27840 35426
rect 27760 35360 27840 35374
rect 27920 35426 28000 35440
rect 27920 35374 27934 35426
rect 27986 35374 28000 35426
rect 27920 35360 28000 35374
rect 28080 35426 28160 35440
rect 28080 35374 28094 35426
rect 28146 35374 28160 35426
rect 28080 35360 28160 35374
rect 28240 35426 28320 35440
rect 28240 35374 28254 35426
rect 28306 35374 28320 35426
rect 28240 35360 28320 35374
rect 28400 35426 28480 35440
rect 28400 35374 28414 35426
rect 28466 35374 28480 35426
rect 28400 35360 28480 35374
rect 28560 35426 28640 35440
rect 28560 35374 28574 35426
rect 28626 35374 28640 35426
rect 28560 35360 28640 35374
rect 28720 35426 28800 35440
rect 28720 35374 28734 35426
rect 28786 35374 28800 35426
rect 28720 35360 28800 35374
rect 28880 35426 28960 35440
rect 28880 35374 28894 35426
rect 28946 35374 28960 35426
rect 28880 35360 28960 35374
rect 29040 35426 29120 35440
rect 29040 35374 29054 35426
rect 29106 35374 29120 35426
rect 29040 35360 29120 35374
rect 29200 35426 29280 35440
rect 29200 35374 29214 35426
rect 29266 35374 29280 35426
rect 29200 35360 29280 35374
rect 29360 35426 29440 35440
rect 29360 35374 29374 35426
rect 29426 35374 29440 35426
rect 29360 35360 29440 35374
rect 33520 35426 33600 35440
rect 33520 35374 33534 35426
rect 33586 35374 33600 35426
rect 33520 35360 33600 35374
rect 33680 35426 33760 35440
rect 33680 35374 33694 35426
rect 33746 35374 33760 35426
rect 33680 35360 33760 35374
rect 33840 35426 33920 35440
rect 33840 35374 33854 35426
rect 33906 35374 33920 35426
rect 33840 35360 33920 35374
rect 34000 35426 34080 35440
rect 34000 35374 34014 35426
rect 34066 35374 34080 35426
rect 34000 35360 34080 35374
rect 34160 35426 34240 35440
rect 34160 35374 34174 35426
rect 34226 35374 34240 35426
rect 34160 35360 34240 35374
rect 34320 35426 34400 35440
rect 34320 35374 34334 35426
rect 34386 35374 34400 35426
rect 34320 35360 34400 35374
rect 34480 35426 34560 35440
rect 34480 35374 34494 35426
rect 34546 35374 34560 35426
rect 34480 35360 34560 35374
rect 34640 35426 34720 35440
rect 34640 35374 34654 35426
rect 34706 35374 34720 35426
rect 34640 35360 34720 35374
rect 34800 35426 34880 35440
rect 34800 35374 34814 35426
rect 34866 35374 34880 35426
rect 34800 35360 34880 35374
rect 34960 35426 35040 35440
rect 34960 35374 34974 35426
rect 35026 35374 35040 35426
rect 34960 35360 35040 35374
rect 35120 35426 35200 35440
rect 35120 35374 35134 35426
rect 35186 35374 35200 35426
rect 35120 35360 35200 35374
rect 35280 35426 35360 35440
rect 35280 35374 35294 35426
rect 35346 35374 35360 35426
rect 35280 35360 35360 35374
rect 35440 35426 35520 35440
rect 35440 35374 35454 35426
rect 35506 35374 35520 35426
rect 35440 35360 35520 35374
rect 35600 35426 35680 35440
rect 35600 35374 35614 35426
rect 35666 35374 35680 35426
rect 35600 35360 35680 35374
rect 35760 35426 35840 35440
rect 35760 35374 35774 35426
rect 35826 35374 35840 35426
rect 35760 35360 35840 35374
rect 35920 35426 36000 35440
rect 35920 35374 35934 35426
rect 35986 35374 36000 35426
rect 35920 35360 36000 35374
rect 36080 35426 36160 35440
rect 36080 35374 36094 35426
rect 36146 35374 36160 35426
rect 36080 35360 36160 35374
rect 36240 35426 36320 35440
rect 36240 35374 36254 35426
rect 36306 35374 36320 35426
rect 36240 35360 36320 35374
rect 36400 35426 36480 35440
rect 36400 35374 36414 35426
rect 36466 35374 36480 35426
rect 36400 35360 36480 35374
rect 36560 35426 36640 35440
rect 36560 35374 36574 35426
rect 36626 35374 36640 35426
rect 36560 35360 36640 35374
rect 36720 35426 36800 35440
rect 36720 35374 36734 35426
rect 36786 35374 36800 35426
rect 36720 35360 36800 35374
rect 36880 35426 36960 35440
rect 36880 35374 36894 35426
rect 36946 35374 36960 35426
rect 36880 35360 36960 35374
rect 37040 35426 37120 35440
rect 37040 35374 37054 35426
rect 37106 35374 37120 35426
rect 37040 35360 37120 35374
rect 37200 35426 37280 35440
rect 37200 35374 37214 35426
rect 37266 35374 37280 35426
rect 37200 35360 37280 35374
rect 37360 35426 37440 35440
rect 37360 35374 37374 35426
rect 37426 35374 37440 35426
rect 37360 35360 37440 35374
rect 37520 35426 37600 35440
rect 37520 35374 37534 35426
rect 37586 35374 37600 35426
rect 37520 35360 37600 35374
rect 37680 35426 37760 35440
rect 37680 35374 37694 35426
rect 37746 35374 37760 35426
rect 37680 35360 37760 35374
rect 37840 35426 37920 35440
rect 37840 35374 37854 35426
rect 37906 35374 37920 35426
rect 37840 35360 37920 35374
rect 38000 35426 38080 35440
rect 38000 35374 38014 35426
rect 38066 35374 38080 35426
rect 38000 35360 38080 35374
rect 38160 35426 38240 35440
rect 38160 35374 38174 35426
rect 38226 35374 38240 35426
rect 38160 35360 38240 35374
rect 38320 35426 38400 35440
rect 38320 35374 38334 35426
rect 38386 35374 38400 35426
rect 38320 35360 38400 35374
rect 38480 35426 38560 35440
rect 38480 35374 38494 35426
rect 38546 35374 38560 35426
rect 38480 35360 38560 35374
rect 38640 35426 38720 35440
rect 38640 35374 38654 35426
rect 38706 35374 38720 35426
rect 38640 35360 38720 35374
rect 38800 35426 38880 35440
rect 38800 35374 38814 35426
rect 38866 35374 38880 35426
rect 38800 35360 38880 35374
rect 38960 35426 39040 35440
rect 38960 35374 38974 35426
rect 39026 35374 39040 35426
rect 38960 35360 39040 35374
rect 39120 35426 39200 35440
rect 39120 35374 39134 35426
rect 39186 35374 39200 35426
rect 39120 35360 39200 35374
rect 39280 35426 39360 35440
rect 39280 35374 39294 35426
rect 39346 35374 39360 35426
rect 39280 35360 39360 35374
rect 39440 35426 39520 35440
rect 39440 35374 39454 35426
rect 39506 35374 39520 35426
rect 39440 35360 39520 35374
rect 39600 35426 39680 35440
rect 39600 35374 39614 35426
rect 39666 35374 39680 35426
rect 39600 35360 39680 35374
rect 39760 35426 39840 35440
rect 39760 35374 39774 35426
rect 39826 35374 39840 35426
rect 39760 35360 39840 35374
rect 39920 35426 40000 35440
rect 39920 35374 39934 35426
rect 39986 35374 40000 35426
rect 39920 35360 40000 35374
rect 40080 35426 40160 35440
rect 40080 35374 40094 35426
rect 40146 35374 40160 35426
rect 40080 35360 40160 35374
rect 40240 35426 40320 35440
rect 40240 35374 40254 35426
rect 40306 35374 40320 35426
rect 40240 35360 40320 35374
rect 40400 35426 40480 35440
rect 40400 35374 40414 35426
rect 40466 35374 40480 35426
rect 40400 35360 40480 35374
rect 40560 35426 40640 35440
rect 40560 35374 40574 35426
rect 40626 35374 40640 35426
rect 40560 35360 40640 35374
rect 40720 35426 40800 35440
rect 40720 35374 40734 35426
rect 40786 35374 40800 35426
rect 40720 35360 40800 35374
rect 40880 35426 40960 35440
rect 40880 35374 40894 35426
rect 40946 35374 40960 35426
rect 40880 35360 40960 35374
rect 41040 35426 41120 35440
rect 41040 35374 41054 35426
rect 41106 35374 41120 35426
rect 41040 35360 41120 35374
rect 41200 35426 41280 35440
rect 41200 35374 41214 35426
rect 41266 35374 41280 35426
rect 41200 35360 41280 35374
rect 41360 35426 41440 35440
rect 41360 35374 41374 35426
rect 41426 35374 41440 35426
rect 41360 35360 41440 35374
rect 41520 35426 41600 35440
rect 41520 35374 41534 35426
rect 41586 35374 41600 35426
rect 41520 35360 41600 35374
rect 41680 35426 41760 35440
rect 41680 35374 41694 35426
rect 41746 35374 41760 35426
rect 41680 35360 41760 35374
rect 41840 35426 41920 35440
rect 41840 35374 41854 35426
rect 41906 35374 41920 35426
rect 41840 35360 41920 35374
rect 0 35106 80 35120
rect 0 35054 14 35106
rect 66 35054 80 35106
rect 0 35040 80 35054
rect 160 35106 240 35120
rect 160 35054 174 35106
rect 226 35054 240 35106
rect 160 35040 240 35054
rect 320 35106 400 35120
rect 320 35054 334 35106
rect 386 35054 400 35106
rect 320 35040 400 35054
rect 480 35106 560 35120
rect 480 35054 494 35106
rect 546 35054 560 35106
rect 480 35040 560 35054
rect 640 35106 720 35120
rect 640 35054 654 35106
rect 706 35054 720 35106
rect 640 35040 720 35054
rect 800 35106 880 35120
rect 800 35054 814 35106
rect 866 35054 880 35106
rect 800 35040 880 35054
rect 960 35106 1040 35120
rect 960 35054 974 35106
rect 1026 35054 1040 35106
rect 960 35040 1040 35054
rect 1120 35106 1200 35120
rect 1120 35054 1134 35106
rect 1186 35054 1200 35106
rect 1120 35040 1200 35054
rect 1280 35106 1360 35120
rect 1280 35054 1294 35106
rect 1346 35054 1360 35106
rect 1280 35040 1360 35054
rect 1440 35106 1520 35120
rect 1440 35054 1454 35106
rect 1506 35054 1520 35106
rect 1440 35040 1520 35054
rect 1600 35106 1680 35120
rect 1600 35054 1614 35106
rect 1666 35054 1680 35106
rect 1600 35040 1680 35054
rect 1760 35106 1840 35120
rect 1760 35054 1774 35106
rect 1826 35054 1840 35106
rect 1760 35040 1840 35054
rect 1920 35106 2000 35120
rect 1920 35054 1934 35106
rect 1986 35054 2000 35106
rect 1920 35040 2000 35054
rect 2080 35106 2160 35120
rect 2080 35054 2094 35106
rect 2146 35054 2160 35106
rect 2080 35040 2160 35054
rect 2240 35106 2320 35120
rect 2240 35054 2254 35106
rect 2306 35054 2320 35106
rect 2240 35040 2320 35054
rect 2400 35106 2480 35120
rect 2400 35054 2414 35106
rect 2466 35054 2480 35106
rect 2400 35040 2480 35054
rect 2560 35106 2640 35120
rect 2560 35054 2574 35106
rect 2626 35054 2640 35106
rect 2560 35040 2640 35054
rect 2720 35106 2800 35120
rect 2720 35054 2734 35106
rect 2786 35054 2800 35106
rect 2720 35040 2800 35054
rect 2880 35106 2960 35120
rect 2880 35054 2894 35106
rect 2946 35054 2960 35106
rect 2880 35040 2960 35054
rect 3040 35106 3120 35120
rect 3040 35054 3054 35106
rect 3106 35054 3120 35106
rect 3040 35040 3120 35054
rect 3200 35106 3280 35120
rect 3200 35054 3214 35106
rect 3266 35054 3280 35106
rect 3200 35040 3280 35054
rect 3360 35106 3440 35120
rect 3360 35054 3374 35106
rect 3426 35054 3440 35106
rect 3360 35040 3440 35054
rect 3520 35106 3600 35120
rect 3520 35054 3534 35106
rect 3586 35054 3600 35106
rect 3520 35040 3600 35054
rect 3680 35106 3760 35120
rect 3680 35054 3694 35106
rect 3746 35054 3760 35106
rect 3680 35040 3760 35054
rect 3840 35106 3920 35120
rect 3840 35054 3854 35106
rect 3906 35054 3920 35106
rect 3840 35040 3920 35054
rect 4000 35106 4080 35120
rect 4000 35054 4014 35106
rect 4066 35054 4080 35106
rect 4000 35040 4080 35054
rect 4160 35106 4240 35120
rect 4160 35054 4174 35106
rect 4226 35054 4240 35106
rect 4160 35040 4240 35054
rect 4320 35106 4400 35120
rect 4320 35054 4334 35106
rect 4386 35054 4400 35106
rect 4320 35040 4400 35054
rect 4480 35106 4560 35120
rect 4480 35054 4494 35106
rect 4546 35054 4560 35106
rect 4480 35040 4560 35054
rect 4640 35106 4720 35120
rect 4640 35054 4654 35106
rect 4706 35054 4720 35106
rect 4640 35040 4720 35054
rect 4800 35106 4880 35120
rect 4800 35054 4814 35106
rect 4866 35054 4880 35106
rect 4800 35040 4880 35054
rect 4960 35106 5040 35120
rect 4960 35054 4974 35106
rect 5026 35054 5040 35106
rect 4960 35040 5040 35054
rect 5120 35106 5200 35120
rect 5120 35054 5134 35106
rect 5186 35054 5200 35106
rect 5120 35040 5200 35054
rect 5280 35106 5360 35120
rect 5280 35054 5294 35106
rect 5346 35054 5360 35106
rect 5280 35040 5360 35054
rect 5440 35106 5520 35120
rect 5440 35054 5454 35106
rect 5506 35054 5520 35106
rect 5440 35040 5520 35054
rect 5600 35106 5680 35120
rect 5600 35054 5614 35106
rect 5666 35054 5680 35106
rect 5600 35040 5680 35054
rect 5760 35106 5840 35120
rect 5760 35054 5774 35106
rect 5826 35054 5840 35106
rect 5760 35040 5840 35054
rect 5920 35106 6000 35120
rect 5920 35054 5934 35106
rect 5986 35054 6000 35106
rect 5920 35040 6000 35054
rect 6080 35106 6160 35120
rect 6080 35054 6094 35106
rect 6146 35054 6160 35106
rect 6080 35040 6160 35054
rect 6240 35106 6320 35120
rect 6240 35054 6254 35106
rect 6306 35054 6320 35106
rect 6240 35040 6320 35054
rect 6400 35106 6480 35120
rect 6400 35054 6414 35106
rect 6466 35054 6480 35106
rect 6400 35040 6480 35054
rect 6560 35106 6640 35120
rect 6560 35054 6574 35106
rect 6626 35054 6640 35106
rect 6560 35040 6640 35054
rect 6720 35106 6800 35120
rect 6720 35054 6734 35106
rect 6786 35054 6800 35106
rect 6720 35040 6800 35054
rect 6880 35106 6960 35120
rect 6880 35054 6894 35106
rect 6946 35054 6960 35106
rect 6880 35040 6960 35054
rect 7040 35106 7120 35120
rect 7040 35054 7054 35106
rect 7106 35054 7120 35106
rect 7040 35040 7120 35054
rect 7200 35106 7280 35120
rect 7200 35054 7214 35106
rect 7266 35054 7280 35106
rect 7200 35040 7280 35054
rect 7360 35106 7440 35120
rect 7360 35054 7374 35106
rect 7426 35054 7440 35106
rect 7360 35040 7440 35054
rect 7520 35106 7600 35120
rect 7520 35054 7534 35106
rect 7586 35054 7600 35106
rect 7520 35040 7600 35054
rect 7680 35106 7760 35120
rect 7680 35054 7694 35106
rect 7746 35054 7760 35106
rect 7680 35040 7760 35054
rect 7840 35106 7920 35120
rect 7840 35054 7854 35106
rect 7906 35054 7920 35106
rect 7840 35040 7920 35054
rect 8000 35106 8080 35120
rect 8000 35054 8014 35106
rect 8066 35054 8080 35106
rect 8000 35040 8080 35054
rect 8160 35106 8240 35120
rect 8160 35054 8174 35106
rect 8226 35054 8240 35106
rect 8160 35040 8240 35054
rect 8320 35106 8400 35120
rect 8320 35054 8334 35106
rect 8386 35054 8400 35106
rect 8320 35040 8400 35054
rect 12480 35106 12560 35120
rect 12480 35054 12494 35106
rect 12546 35054 12560 35106
rect 12480 35040 12560 35054
rect 12640 35106 12720 35120
rect 12640 35054 12654 35106
rect 12706 35054 12720 35106
rect 12640 35040 12720 35054
rect 12800 35106 12880 35120
rect 12800 35054 12814 35106
rect 12866 35054 12880 35106
rect 12800 35040 12880 35054
rect 12960 35106 13040 35120
rect 12960 35054 12974 35106
rect 13026 35054 13040 35106
rect 12960 35040 13040 35054
rect 13120 35106 13200 35120
rect 13120 35054 13134 35106
rect 13186 35054 13200 35106
rect 13120 35040 13200 35054
rect 13280 35106 13360 35120
rect 13280 35054 13294 35106
rect 13346 35054 13360 35106
rect 13280 35040 13360 35054
rect 13440 35106 13520 35120
rect 13440 35054 13454 35106
rect 13506 35054 13520 35106
rect 13440 35040 13520 35054
rect 13600 35106 13680 35120
rect 13600 35054 13614 35106
rect 13666 35054 13680 35106
rect 13600 35040 13680 35054
rect 13760 35106 13840 35120
rect 13760 35054 13774 35106
rect 13826 35054 13840 35106
rect 13760 35040 13840 35054
rect 13920 35106 14000 35120
rect 13920 35054 13934 35106
rect 13986 35054 14000 35106
rect 13920 35040 14000 35054
rect 14080 35106 14160 35120
rect 14080 35054 14094 35106
rect 14146 35054 14160 35106
rect 14080 35040 14160 35054
rect 14240 35106 14320 35120
rect 14240 35054 14254 35106
rect 14306 35054 14320 35106
rect 14240 35040 14320 35054
rect 14400 35106 14480 35120
rect 14400 35054 14414 35106
rect 14466 35054 14480 35106
rect 14400 35040 14480 35054
rect 14560 35106 14640 35120
rect 14560 35054 14574 35106
rect 14626 35054 14640 35106
rect 14560 35040 14640 35054
rect 14720 35106 14800 35120
rect 14720 35054 14734 35106
rect 14786 35054 14800 35106
rect 14720 35040 14800 35054
rect 14880 35106 14960 35120
rect 14880 35054 14894 35106
rect 14946 35054 14960 35106
rect 14880 35040 14960 35054
rect 15040 35106 15120 35120
rect 15040 35054 15054 35106
rect 15106 35054 15120 35106
rect 15040 35040 15120 35054
rect 15200 35106 15280 35120
rect 15200 35054 15214 35106
rect 15266 35054 15280 35106
rect 15200 35040 15280 35054
rect 15360 35106 15440 35120
rect 15360 35054 15374 35106
rect 15426 35054 15440 35106
rect 15360 35040 15440 35054
rect 15520 35106 15600 35120
rect 15520 35054 15534 35106
rect 15586 35054 15600 35106
rect 15520 35040 15600 35054
rect 15680 35106 15760 35120
rect 15680 35054 15694 35106
rect 15746 35054 15760 35106
rect 15680 35040 15760 35054
rect 15840 35106 15920 35120
rect 15840 35054 15854 35106
rect 15906 35054 15920 35106
rect 15840 35040 15920 35054
rect 16000 35106 16080 35120
rect 16000 35054 16014 35106
rect 16066 35054 16080 35106
rect 16000 35040 16080 35054
rect 16160 35106 16240 35120
rect 16160 35054 16174 35106
rect 16226 35054 16240 35106
rect 16160 35040 16240 35054
rect 16320 35106 16400 35120
rect 16320 35054 16334 35106
rect 16386 35054 16400 35106
rect 16320 35040 16400 35054
rect 16480 35106 16560 35120
rect 16480 35054 16494 35106
rect 16546 35054 16560 35106
rect 16480 35040 16560 35054
rect 16640 35106 16720 35120
rect 16640 35054 16654 35106
rect 16706 35054 16720 35106
rect 16640 35040 16720 35054
rect 16800 35106 16880 35120
rect 16800 35054 16814 35106
rect 16866 35054 16880 35106
rect 16800 35040 16880 35054
rect 16960 35106 17040 35120
rect 16960 35054 16974 35106
rect 17026 35054 17040 35106
rect 16960 35040 17040 35054
rect 17120 35106 17200 35120
rect 17120 35054 17134 35106
rect 17186 35054 17200 35106
rect 17120 35040 17200 35054
rect 17280 35106 17360 35120
rect 17280 35054 17294 35106
rect 17346 35054 17360 35106
rect 17280 35040 17360 35054
rect 17440 35106 17520 35120
rect 17440 35054 17454 35106
rect 17506 35054 17520 35106
rect 17440 35040 17520 35054
rect 17600 35106 17680 35120
rect 17600 35054 17614 35106
rect 17666 35054 17680 35106
rect 17600 35040 17680 35054
rect 17760 35106 17840 35120
rect 17760 35054 17774 35106
rect 17826 35054 17840 35106
rect 17760 35040 17840 35054
rect 17920 35106 18000 35120
rect 17920 35054 17934 35106
rect 17986 35054 18000 35106
rect 17920 35040 18000 35054
rect 18080 35106 18160 35120
rect 18080 35054 18094 35106
rect 18146 35054 18160 35106
rect 18080 35040 18160 35054
rect 18240 35106 18320 35120
rect 18240 35054 18254 35106
rect 18306 35054 18320 35106
rect 18240 35040 18320 35054
rect 18400 35106 18480 35120
rect 18400 35054 18414 35106
rect 18466 35054 18480 35106
rect 18400 35040 18480 35054
rect 18560 35106 18640 35120
rect 18560 35054 18574 35106
rect 18626 35054 18640 35106
rect 18560 35040 18640 35054
rect 18720 35106 18800 35120
rect 18720 35054 18734 35106
rect 18786 35054 18800 35106
rect 18720 35040 18800 35054
rect 18880 35106 18960 35120
rect 18880 35054 18894 35106
rect 18946 35054 18960 35106
rect 18880 35040 18960 35054
rect 23120 35106 23200 35120
rect 23120 35054 23134 35106
rect 23186 35054 23200 35106
rect 23120 35040 23200 35054
rect 23280 35106 23360 35120
rect 23280 35054 23294 35106
rect 23346 35054 23360 35106
rect 23280 35040 23360 35054
rect 23440 35106 23520 35120
rect 23440 35054 23454 35106
rect 23506 35054 23520 35106
rect 23440 35040 23520 35054
rect 23600 35106 23680 35120
rect 23600 35054 23614 35106
rect 23666 35054 23680 35106
rect 23600 35040 23680 35054
rect 23760 35106 23840 35120
rect 23760 35054 23774 35106
rect 23826 35054 23840 35106
rect 23760 35040 23840 35054
rect 23920 35106 24000 35120
rect 23920 35054 23934 35106
rect 23986 35054 24000 35106
rect 23920 35040 24000 35054
rect 24080 35106 24160 35120
rect 24080 35054 24094 35106
rect 24146 35054 24160 35106
rect 24080 35040 24160 35054
rect 24240 35106 24320 35120
rect 24240 35054 24254 35106
rect 24306 35054 24320 35106
rect 24240 35040 24320 35054
rect 24400 35106 24480 35120
rect 24400 35054 24414 35106
rect 24466 35054 24480 35106
rect 24400 35040 24480 35054
rect 24560 35106 24640 35120
rect 24560 35054 24574 35106
rect 24626 35054 24640 35106
rect 24560 35040 24640 35054
rect 24720 35106 24800 35120
rect 24720 35054 24734 35106
rect 24786 35054 24800 35106
rect 24720 35040 24800 35054
rect 24880 35106 24960 35120
rect 24880 35054 24894 35106
rect 24946 35054 24960 35106
rect 24880 35040 24960 35054
rect 25040 35106 25120 35120
rect 25040 35054 25054 35106
rect 25106 35054 25120 35106
rect 25040 35040 25120 35054
rect 25200 35106 25280 35120
rect 25200 35054 25214 35106
rect 25266 35054 25280 35106
rect 25200 35040 25280 35054
rect 25360 35106 25440 35120
rect 25360 35054 25374 35106
rect 25426 35054 25440 35106
rect 25360 35040 25440 35054
rect 25520 35106 25600 35120
rect 25520 35054 25534 35106
rect 25586 35054 25600 35106
rect 25520 35040 25600 35054
rect 25680 35106 25760 35120
rect 25680 35054 25694 35106
rect 25746 35054 25760 35106
rect 25680 35040 25760 35054
rect 25840 35106 25920 35120
rect 25840 35054 25854 35106
rect 25906 35054 25920 35106
rect 25840 35040 25920 35054
rect 26000 35106 26080 35120
rect 26000 35054 26014 35106
rect 26066 35054 26080 35106
rect 26000 35040 26080 35054
rect 26160 35106 26240 35120
rect 26160 35054 26174 35106
rect 26226 35054 26240 35106
rect 26160 35040 26240 35054
rect 26320 35106 26400 35120
rect 26320 35054 26334 35106
rect 26386 35054 26400 35106
rect 26320 35040 26400 35054
rect 26480 35106 26560 35120
rect 26480 35054 26494 35106
rect 26546 35054 26560 35106
rect 26480 35040 26560 35054
rect 26640 35106 26720 35120
rect 26640 35054 26654 35106
rect 26706 35054 26720 35106
rect 26640 35040 26720 35054
rect 26800 35106 26880 35120
rect 26800 35054 26814 35106
rect 26866 35054 26880 35106
rect 26800 35040 26880 35054
rect 26960 35106 27040 35120
rect 26960 35054 26974 35106
rect 27026 35054 27040 35106
rect 26960 35040 27040 35054
rect 27120 35106 27200 35120
rect 27120 35054 27134 35106
rect 27186 35054 27200 35106
rect 27120 35040 27200 35054
rect 27280 35106 27360 35120
rect 27280 35054 27294 35106
rect 27346 35054 27360 35106
rect 27280 35040 27360 35054
rect 27440 35106 27520 35120
rect 27440 35054 27454 35106
rect 27506 35054 27520 35106
rect 27440 35040 27520 35054
rect 27600 35106 27680 35120
rect 27600 35054 27614 35106
rect 27666 35054 27680 35106
rect 27600 35040 27680 35054
rect 27760 35106 27840 35120
rect 27760 35054 27774 35106
rect 27826 35054 27840 35106
rect 27760 35040 27840 35054
rect 27920 35106 28000 35120
rect 27920 35054 27934 35106
rect 27986 35054 28000 35106
rect 27920 35040 28000 35054
rect 28080 35106 28160 35120
rect 28080 35054 28094 35106
rect 28146 35054 28160 35106
rect 28080 35040 28160 35054
rect 28240 35106 28320 35120
rect 28240 35054 28254 35106
rect 28306 35054 28320 35106
rect 28240 35040 28320 35054
rect 28400 35106 28480 35120
rect 28400 35054 28414 35106
rect 28466 35054 28480 35106
rect 28400 35040 28480 35054
rect 28560 35106 28640 35120
rect 28560 35054 28574 35106
rect 28626 35054 28640 35106
rect 28560 35040 28640 35054
rect 28720 35106 28800 35120
rect 28720 35054 28734 35106
rect 28786 35054 28800 35106
rect 28720 35040 28800 35054
rect 28880 35106 28960 35120
rect 28880 35054 28894 35106
rect 28946 35054 28960 35106
rect 28880 35040 28960 35054
rect 29040 35106 29120 35120
rect 29040 35054 29054 35106
rect 29106 35054 29120 35106
rect 29040 35040 29120 35054
rect 29200 35106 29280 35120
rect 29200 35054 29214 35106
rect 29266 35054 29280 35106
rect 29200 35040 29280 35054
rect 29360 35106 29440 35120
rect 29360 35054 29374 35106
rect 29426 35054 29440 35106
rect 29360 35040 29440 35054
rect 33520 35106 33600 35120
rect 33520 35054 33534 35106
rect 33586 35054 33600 35106
rect 33520 35040 33600 35054
rect 33680 35106 33760 35120
rect 33680 35054 33694 35106
rect 33746 35054 33760 35106
rect 33680 35040 33760 35054
rect 33840 35106 33920 35120
rect 33840 35054 33854 35106
rect 33906 35054 33920 35106
rect 33840 35040 33920 35054
rect 34000 35106 34080 35120
rect 34000 35054 34014 35106
rect 34066 35054 34080 35106
rect 34000 35040 34080 35054
rect 34160 35106 34240 35120
rect 34160 35054 34174 35106
rect 34226 35054 34240 35106
rect 34160 35040 34240 35054
rect 34320 35106 34400 35120
rect 34320 35054 34334 35106
rect 34386 35054 34400 35106
rect 34320 35040 34400 35054
rect 34480 35106 34560 35120
rect 34480 35054 34494 35106
rect 34546 35054 34560 35106
rect 34480 35040 34560 35054
rect 34640 35106 34720 35120
rect 34640 35054 34654 35106
rect 34706 35054 34720 35106
rect 34640 35040 34720 35054
rect 34800 35106 34880 35120
rect 34800 35054 34814 35106
rect 34866 35054 34880 35106
rect 34800 35040 34880 35054
rect 34960 35106 35040 35120
rect 34960 35054 34974 35106
rect 35026 35054 35040 35106
rect 34960 35040 35040 35054
rect 35120 35106 35200 35120
rect 35120 35054 35134 35106
rect 35186 35054 35200 35106
rect 35120 35040 35200 35054
rect 35280 35106 35360 35120
rect 35280 35054 35294 35106
rect 35346 35054 35360 35106
rect 35280 35040 35360 35054
rect 35440 35106 35520 35120
rect 35440 35054 35454 35106
rect 35506 35054 35520 35106
rect 35440 35040 35520 35054
rect 35600 35106 35680 35120
rect 35600 35054 35614 35106
rect 35666 35054 35680 35106
rect 35600 35040 35680 35054
rect 35760 35106 35840 35120
rect 35760 35054 35774 35106
rect 35826 35054 35840 35106
rect 35760 35040 35840 35054
rect 35920 35106 36000 35120
rect 35920 35054 35934 35106
rect 35986 35054 36000 35106
rect 35920 35040 36000 35054
rect 36080 35106 36160 35120
rect 36080 35054 36094 35106
rect 36146 35054 36160 35106
rect 36080 35040 36160 35054
rect 36240 35106 36320 35120
rect 36240 35054 36254 35106
rect 36306 35054 36320 35106
rect 36240 35040 36320 35054
rect 36400 35106 36480 35120
rect 36400 35054 36414 35106
rect 36466 35054 36480 35106
rect 36400 35040 36480 35054
rect 36560 35106 36640 35120
rect 36560 35054 36574 35106
rect 36626 35054 36640 35106
rect 36560 35040 36640 35054
rect 36720 35106 36800 35120
rect 36720 35054 36734 35106
rect 36786 35054 36800 35106
rect 36720 35040 36800 35054
rect 36880 35106 36960 35120
rect 36880 35054 36894 35106
rect 36946 35054 36960 35106
rect 36880 35040 36960 35054
rect 37040 35106 37120 35120
rect 37040 35054 37054 35106
rect 37106 35054 37120 35106
rect 37040 35040 37120 35054
rect 37200 35106 37280 35120
rect 37200 35054 37214 35106
rect 37266 35054 37280 35106
rect 37200 35040 37280 35054
rect 37360 35106 37440 35120
rect 37360 35054 37374 35106
rect 37426 35054 37440 35106
rect 37360 35040 37440 35054
rect 37520 35106 37600 35120
rect 37520 35054 37534 35106
rect 37586 35054 37600 35106
rect 37520 35040 37600 35054
rect 37680 35106 37760 35120
rect 37680 35054 37694 35106
rect 37746 35054 37760 35106
rect 37680 35040 37760 35054
rect 37840 35106 37920 35120
rect 37840 35054 37854 35106
rect 37906 35054 37920 35106
rect 37840 35040 37920 35054
rect 38000 35106 38080 35120
rect 38000 35054 38014 35106
rect 38066 35054 38080 35106
rect 38000 35040 38080 35054
rect 38160 35106 38240 35120
rect 38160 35054 38174 35106
rect 38226 35054 38240 35106
rect 38160 35040 38240 35054
rect 38320 35106 38400 35120
rect 38320 35054 38334 35106
rect 38386 35054 38400 35106
rect 38320 35040 38400 35054
rect 38480 35106 38560 35120
rect 38480 35054 38494 35106
rect 38546 35054 38560 35106
rect 38480 35040 38560 35054
rect 38640 35106 38720 35120
rect 38640 35054 38654 35106
rect 38706 35054 38720 35106
rect 38640 35040 38720 35054
rect 38800 35106 38880 35120
rect 38800 35054 38814 35106
rect 38866 35054 38880 35106
rect 38800 35040 38880 35054
rect 38960 35106 39040 35120
rect 38960 35054 38974 35106
rect 39026 35054 39040 35106
rect 38960 35040 39040 35054
rect 39120 35106 39200 35120
rect 39120 35054 39134 35106
rect 39186 35054 39200 35106
rect 39120 35040 39200 35054
rect 39280 35106 39360 35120
rect 39280 35054 39294 35106
rect 39346 35054 39360 35106
rect 39280 35040 39360 35054
rect 39440 35106 39520 35120
rect 39440 35054 39454 35106
rect 39506 35054 39520 35106
rect 39440 35040 39520 35054
rect 39600 35106 39680 35120
rect 39600 35054 39614 35106
rect 39666 35054 39680 35106
rect 39600 35040 39680 35054
rect 39760 35106 39840 35120
rect 39760 35054 39774 35106
rect 39826 35054 39840 35106
rect 39760 35040 39840 35054
rect 39920 35106 40000 35120
rect 39920 35054 39934 35106
rect 39986 35054 40000 35106
rect 39920 35040 40000 35054
rect 40080 35106 40160 35120
rect 40080 35054 40094 35106
rect 40146 35054 40160 35106
rect 40080 35040 40160 35054
rect 40240 35106 40320 35120
rect 40240 35054 40254 35106
rect 40306 35054 40320 35106
rect 40240 35040 40320 35054
rect 40400 35106 40480 35120
rect 40400 35054 40414 35106
rect 40466 35054 40480 35106
rect 40400 35040 40480 35054
rect 40560 35106 40640 35120
rect 40560 35054 40574 35106
rect 40626 35054 40640 35106
rect 40560 35040 40640 35054
rect 40720 35106 40800 35120
rect 40720 35054 40734 35106
rect 40786 35054 40800 35106
rect 40720 35040 40800 35054
rect 40880 35106 40960 35120
rect 40880 35054 40894 35106
rect 40946 35054 40960 35106
rect 40880 35040 40960 35054
rect 41040 35106 41120 35120
rect 41040 35054 41054 35106
rect 41106 35054 41120 35106
rect 41040 35040 41120 35054
rect 41200 35106 41280 35120
rect 41200 35054 41214 35106
rect 41266 35054 41280 35106
rect 41200 35040 41280 35054
rect 41360 35106 41440 35120
rect 41360 35054 41374 35106
rect 41426 35054 41440 35106
rect 41360 35040 41440 35054
rect 41520 35106 41600 35120
rect 41520 35054 41534 35106
rect 41586 35054 41600 35106
rect 41520 35040 41600 35054
rect 41680 35106 41760 35120
rect 41680 35054 41694 35106
rect 41746 35054 41760 35106
rect 41680 35040 41760 35054
rect 41840 35106 41920 35120
rect 41840 35054 41854 35106
rect 41906 35054 41920 35106
rect 41840 35040 41920 35054
rect 0 34786 80 34800
rect 0 34734 14 34786
rect 66 34734 80 34786
rect 0 34720 80 34734
rect 160 34786 240 34800
rect 160 34734 174 34786
rect 226 34734 240 34786
rect 160 34720 240 34734
rect 320 34786 400 34800
rect 320 34734 334 34786
rect 386 34734 400 34786
rect 320 34720 400 34734
rect 480 34786 560 34800
rect 480 34734 494 34786
rect 546 34734 560 34786
rect 480 34720 560 34734
rect 640 34786 720 34800
rect 640 34734 654 34786
rect 706 34734 720 34786
rect 640 34720 720 34734
rect 800 34786 880 34800
rect 800 34734 814 34786
rect 866 34734 880 34786
rect 800 34720 880 34734
rect 960 34786 1040 34800
rect 960 34734 974 34786
rect 1026 34734 1040 34786
rect 960 34720 1040 34734
rect 1120 34786 1200 34800
rect 1120 34734 1134 34786
rect 1186 34734 1200 34786
rect 1120 34720 1200 34734
rect 1280 34786 1360 34800
rect 1280 34734 1294 34786
rect 1346 34734 1360 34786
rect 1280 34720 1360 34734
rect 1440 34786 1520 34800
rect 1440 34734 1454 34786
rect 1506 34734 1520 34786
rect 1440 34720 1520 34734
rect 1600 34786 1680 34800
rect 1600 34734 1614 34786
rect 1666 34734 1680 34786
rect 1600 34720 1680 34734
rect 1760 34786 1840 34800
rect 1760 34734 1774 34786
rect 1826 34734 1840 34786
rect 1760 34720 1840 34734
rect 1920 34786 2000 34800
rect 1920 34734 1934 34786
rect 1986 34734 2000 34786
rect 1920 34720 2000 34734
rect 2080 34786 2160 34800
rect 2080 34734 2094 34786
rect 2146 34734 2160 34786
rect 2080 34720 2160 34734
rect 2240 34786 2320 34800
rect 2240 34734 2254 34786
rect 2306 34734 2320 34786
rect 2240 34720 2320 34734
rect 2400 34786 2480 34800
rect 2400 34734 2414 34786
rect 2466 34734 2480 34786
rect 2400 34720 2480 34734
rect 2560 34786 2640 34800
rect 2560 34734 2574 34786
rect 2626 34734 2640 34786
rect 2560 34720 2640 34734
rect 2720 34786 2800 34800
rect 2720 34734 2734 34786
rect 2786 34734 2800 34786
rect 2720 34720 2800 34734
rect 2880 34786 2960 34800
rect 2880 34734 2894 34786
rect 2946 34734 2960 34786
rect 2880 34720 2960 34734
rect 3040 34786 3120 34800
rect 3040 34734 3054 34786
rect 3106 34734 3120 34786
rect 3040 34720 3120 34734
rect 3200 34786 3280 34800
rect 3200 34734 3214 34786
rect 3266 34734 3280 34786
rect 3200 34720 3280 34734
rect 3360 34786 3440 34800
rect 3360 34734 3374 34786
rect 3426 34734 3440 34786
rect 3360 34720 3440 34734
rect 3520 34786 3600 34800
rect 3520 34734 3534 34786
rect 3586 34734 3600 34786
rect 3520 34720 3600 34734
rect 3680 34786 3760 34800
rect 3680 34734 3694 34786
rect 3746 34734 3760 34786
rect 3680 34720 3760 34734
rect 3840 34786 3920 34800
rect 3840 34734 3854 34786
rect 3906 34734 3920 34786
rect 3840 34720 3920 34734
rect 4000 34786 4080 34800
rect 4000 34734 4014 34786
rect 4066 34734 4080 34786
rect 4000 34720 4080 34734
rect 4160 34786 4240 34800
rect 4160 34734 4174 34786
rect 4226 34734 4240 34786
rect 4160 34720 4240 34734
rect 4320 34786 4400 34800
rect 4320 34734 4334 34786
rect 4386 34734 4400 34786
rect 4320 34720 4400 34734
rect 4480 34786 4560 34800
rect 4480 34734 4494 34786
rect 4546 34734 4560 34786
rect 4480 34720 4560 34734
rect 4640 34786 4720 34800
rect 4640 34734 4654 34786
rect 4706 34734 4720 34786
rect 4640 34720 4720 34734
rect 4800 34786 4880 34800
rect 4800 34734 4814 34786
rect 4866 34734 4880 34786
rect 4800 34720 4880 34734
rect 4960 34786 5040 34800
rect 4960 34734 4974 34786
rect 5026 34734 5040 34786
rect 4960 34720 5040 34734
rect 5120 34786 5200 34800
rect 5120 34734 5134 34786
rect 5186 34734 5200 34786
rect 5120 34720 5200 34734
rect 5280 34786 5360 34800
rect 5280 34734 5294 34786
rect 5346 34734 5360 34786
rect 5280 34720 5360 34734
rect 5440 34786 5520 34800
rect 5440 34734 5454 34786
rect 5506 34734 5520 34786
rect 5440 34720 5520 34734
rect 5600 34786 5680 34800
rect 5600 34734 5614 34786
rect 5666 34734 5680 34786
rect 5600 34720 5680 34734
rect 5760 34786 5840 34800
rect 5760 34734 5774 34786
rect 5826 34734 5840 34786
rect 5760 34720 5840 34734
rect 5920 34786 6000 34800
rect 5920 34734 5934 34786
rect 5986 34734 6000 34786
rect 5920 34720 6000 34734
rect 6080 34786 6160 34800
rect 6080 34734 6094 34786
rect 6146 34734 6160 34786
rect 6080 34720 6160 34734
rect 6240 34786 6320 34800
rect 6240 34734 6254 34786
rect 6306 34734 6320 34786
rect 6240 34720 6320 34734
rect 6400 34786 6480 34800
rect 6400 34734 6414 34786
rect 6466 34734 6480 34786
rect 6400 34720 6480 34734
rect 6560 34786 6640 34800
rect 6560 34734 6574 34786
rect 6626 34734 6640 34786
rect 6560 34720 6640 34734
rect 6720 34786 6800 34800
rect 6720 34734 6734 34786
rect 6786 34734 6800 34786
rect 6720 34720 6800 34734
rect 6880 34786 6960 34800
rect 6880 34734 6894 34786
rect 6946 34734 6960 34786
rect 6880 34720 6960 34734
rect 7040 34786 7120 34800
rect 7040 34734 7054 34786
rect 7106 34734 7120 34786
rect 7040 34720 7120 34734
rect 7200 34786 7280 34800
rect 7200 34734 7214 34786
rect 7266 34734 7280 34786
rect 7200 34720 7280 34734
rect 7360 34786 7440 34800
rect 7360 34734 7374 34786
rect 7426 34734 7440 34786
rect 7360 34720 7440 34734
rect 7520 34786 7600 34800
rect 7520 34734 7534 34786
rect 7586 34734 7600 34786
rect 7520 34720 7600 34734
rect 7680 34786 7760 34800
rect 7680 34734 7694 34786
rect 7746 34734 7760 34786
rect 7680 34720 7760 34734
rect 7840 34786 7920 34800
rect 7840 34734 7854 34786
rect 7906 34734 7920 34786
rect 7840 34720 7920 34734
rect 8000 34786 8080 34800
rect 8000 34734 8014 34786
rect 8066 34734 8080 34786
rect 8000 34720 8080 34734
rect 8160 34786 8240 34800
rect 8160 34734 8174 34786
rect 8226 34734 8240 34786
rect 8160 34720 8240 34734
rect 8320 34786 8400 34800
rect 8320 34734 8334 34786
rect 8386 34734 8400 34786
rect 8320 34720 8400 34734
rect 12480 34786 12560 34800
rect 12480 34734 12494 34786
rect 12546 34734 12560 34786
rect 12480 34720 12560 34734
rect 12640 34786 12720 34800
rect 12640 34734 12654 34786
rect 12706 34734 12720 34786
rect 12640 34720 12720 34734
rect 12800 34786 12880 34800
rect 12800 34734 12814 34786
rect 12866 34734 12880 34786
rect 12800 34720 12880 34734
rect 12960 34786 13040 34800
rect 12960 34734 12974 34786
rect 13026 34734 13040 34786
rect 12960 34720 13040 34734
rect 13120 34786 13200 34800
rect 13120 34734 13134 34786
rect 13186 34734 13200 34786
rect 13120 34720 13200 34734
rect 13280 34786 13360 34800
rect 13280 34734 13294 34786
rect 13346 34734 13360 34786
rect 13280 34720 13360 34734
rect 13440 34786 13520 34800
rect 13440 34734 13454 34786
rect 13506 34734 13520 34786
rect 13440 34720 13520 34734
rect 13600 34786 13680 34800
rect 13600 34734 13614 34786
rect 13666 34734 13680 34786
rect 13600 34720 13680 34734
rect 13760 34786 13840 34800
rect 13760 34734 13774 34786
rect 13826 34734 13840 34786
rect 13760 34720 13840 34734
rect 13920 34786 14000 34800
rect 13920 34734 13934 34786
rect 13986 34734 14000 34786
rect 13920 34720 14000 34734
rect 14080 34786 14160 34800
rect 14080 34734 14094 34786
rect 14146 34734 14160 34786
rect 14080 34720 14160 34734
rect 14240 34786 14320 34800
rect 14240 34734 14254 34786
rect 14306 34734 14320 34786
rect 14240 34720 14320 34734
rect 14400 34786 14480 34800
rect 14400 34734 14414 34786
rect 14466 34734 14480 34786
rect 14400 34720 14480 34734
rect 14560 34786 14640 34800
rect 14560 34734 14574 34786
rect 14626 34734 14640 34786
rect 14560 34720 14640 34734
rect 14720 34786 14800 34800
rect 14720 34734 14734 34786
rect 14786 34734 14800 34786
rect 14720 34720 14800 34734
rect 14880 34786 14960 34800
rect 14880 34734 14894 34786
rect 14946 34734 14960 34786
rect 14880 34720 14960 34734
rect 15040 34786 15120 34800
rect 15040 34734 15054 34786
rect 15106 34734 15120 34786
rect 15040 34720 15120 34734
rect 15200 34786 15280 34800
rect 15200 34734 15214 34786
rect 15266 34734 15280 34786
rect 15200 34720 15280 34734
rect 15360 34786 15440 34800
rect 15360 34734 15374 34786
rect 15426 34734 15440 34786
rect 15360 34720 15440 34734
rect 15520 34786 15600 34800
rect 15520 34734 15534 34786
rect 15586 34734 15600 34786
rect 15520 34720 15600 34734
rect 15680 34786 15760 34800
rect 15680 34734 15694 34786
rect 15746 34734 15760 34786
rect 15680 34720 15760 34734
rect 15840 34786 15920 34800
rect 15840 34734 15854 34786
rect 15906 34734 15920 34786
rect 15840 34720 15920 34734
rect 16000 34786 16080 34800
rect 16000 34734 16014 34786
rect 16066 34734 16080 34786
rect 16000 34720 16080 34734
rect 16160 34786 16240 34800
rect 16160 34734 16174 34786
rect 16226 34734 16240 34786
rect 16160 34720 16240 34734
rect 16320 34786 16400 34800
rect 16320 34734 16334 34786
rect 16386 34734 16400 34786
rect 16320 34720 16400 34734
rect 16480 34786 16560 34800
rect 16480 34734 16494 34786
rect 16546 34734 16560 34786
rect 16480 34720 16560 34734
rect 16640 34786 16720 34800
rect 16640 34734 16654 34786
rect 16706 34734 16720 34786
rect 16640 34720 16720 34734
rect 16800 34786 16880 34800
rect 16800 34734 16814 34786
rect 16866 34734 16880 34786
rect 16800 34720 16880 34734
rect 16960 34786 17040 34800
rect 16960 34734 16974 34786
rect 17026 34734 17040 34786
rect 16960 34720 17040 34734
rect 17120 34786 17200 34800
rect 17120 34734 17134 34786
rect 17186 34734 17200 34786
rect 17120 34720 17200 34734
rect 17280 34786 17360 34800
rect 17280 34734 17294 34786
rect 17346 34734 17360 34786
rect 17280 34720 17360 34734
rect 17440 34786 17520 34800
rect 17440 34734 17454 34786
rect 17506 34734 17520 34786
rect 17440 34720 17520 34734
rect 17600 34786 17680 34800
rect 17600 34734 17614 34786
rect 17666 34734 17680 34786
rect 17600 34720 17680 34734
rect 17760 34786 17840 34800
rect 17760 34734 17774 34786
rect 17826 34734 17840 34786
rect 17760 34720 17840 34734
rect 17920 34786 18000 34800
rect 17920 34734 17934 34786
rect 17986 34734 18000 34786
rect 17920 34720 18000 34734
rect 18080 34786 18160 34800
rect 18080 34734 18094 34786
rect 18146 34734 18160 34786
rect 18080 34720 18160 34734
rect 18240 34786 18320 34800
rect 18240 34734 18254 34786
rect 18306 34734 18320 34786
rect 18240 34720 18320 34734
rect 18400 34786 18480 34800
rect 18400 34734 18414 34786
rect 18466 34734 18480 34786
rect 18400 34720 18480 34734
rect 18560 34786 18640 34800
rect 18560 34734 18574 34786
rect 18626 34734 18640 34786
rect 18560 34720 18640 34734
rect 18720 34786 18800 34800
rect 18720 34734 18734 34786
rect 18786 34734 18800 34786
rect 18720 34720 18800 34734
rect 18880 34786 18960 34800
rect 18880 34734 18894 34786
rect 18946 34734 18960 34786
rect 18880 34720 18960 34734
rect 23120 34786 23200 34800
rect 23120 34734 23134 34786
rect 23186 34734 23200 34786
rect 23120 34720 23200 34734
rect 23280 34786 23360 34800
rect 23280 34734 23294 34786
rect 23346 34734 23360 34786
rect 23280 34720 23360 34734
rect 23440 34786 23520 34800
rect 23440 34734 23454 34786
rect 23506 34734 23520 34786
rect 23440 34720 23520 34734
rect 23600 34786 23680 34800
rect 23600 34734 23614 34786
rect 23666 34734 23680 34786
rect 23600 34720 23680 34734
rect 23760 34786 23840 34800
rect 23760 34734 23774 34786
rect 23826 34734 23840 34786
rect 23760 34720 23840 34734
rect 23920 34786 24000 34800
rect 23920 34734 23934 34786
rect 23986 34734 24000 34786
rect 23920 34720 24000 34734
rect 24080 34786 24160 34800
rect 24080 34734 24094 34786
rect 24146 34734 24160 34786
rect 24080 34720 24160 34734
rect 24240 34786 24320 34800
rect 24240 34734 24254 34786
rect 24306 34734 24320 34786
rect 24240 34720 24320 34734
rect 24400 34786 24480 34800
rect 24400 34734 24414 34786
rect 24466 34734 24480 34786
rect 24400 34720 24480 34734
rect 24560 34786 24640 34800
rect 24560 34734 24574 34786
rect 24626 34734 24640 34786
rect 24560 34720 24640 34734
rect 24720 34786 24800 34800
rect 24720 34734 24734 34786
rect 24786 34734 24800 34786
rect 24720 34720 24800 34734
rect 24880 34786 24960 34800
rect 24880 34734 24894 34786
rect 24946 34734 24960 34786
rect 24880 34720 24960 34734
rect 25040 34786 25120 34800
rect 25040 34734 25054 34786
rect 25106 34734 25120 34786
rect 25040 34720 25120 34734
rect 25200 34786 25280 34800
rect 25200 34734 25214 34786
rect 25266 34734 25280 34786
rect 25200 34720 25280 34734
rect 25360 34786 25440 34800
rect 25360 34734 25374 34786
rect 25426 34734 25440 34786
rect 25360 34720 25440 34734
rect 25520 34786 25600 34800
rect 25520 34734 25534 34786
rect 25586 34734 25600 34786
rect 25520 34720 25600 34734
rect 25680 34786 25760 34800
rect 25680 34734 25694 34786
rect 25746 34734 25760 34786
rect 25680 34720 25760 34734
rect 25840 34786 25920 34800
rect 25840 34734 25854 34786
rect 25906 34734 25920 34786
rect 25840 34720 25920 34734
rect 26000 34786 26080 34800
rect 26000 34734 26014 34786
rect 26066 34734 26080 34786
rect 26000 34720 26080 34734
rect 26160 34786 26240 34800
rect 26160 34734 26174 34786
rect 26226 34734 26240 34786
rect 26160 34720 26240 34734
rect 26320 34786 26400 34800
rect 26320 34734 26334 34786
rect 26386 34734 26400 34786
rect 26320 34720 26400 34734
rect 26480 34786 26560 34800
rect 26480 34734 26494 34786
rect 26546 34734 26560 34786
rect 26480 34720 26560 34734
rect 26640 34786 26720 34800
rect 26640 34734 26654 34786
rect 26706 34734 26720 34786
rect 26640 34720 26720 34734
rect 26800 34786 26880 34800
rect 26800 34734 26814 34786
rect 26866 34734 26880 34786
rect 26800 34720 26880 34734
rect 26960 34786 27040 34800
rect 26960 34734 26974 34786
rect 27026 34734 27040 34786
rect 26960 34720 27040 34734
rect 27120 34786 27200 34800
rect 27120 34734 27134 34786
rect 27186 34734 27200 34786
rect 27120 34720 27200 34734
rect 27280 34786 27360 34800
rect 27280 34734 27294 34786
rect 27346 34734 27360 34786
rect 27280 34720 27360 34734
rect 27440 34786 27520 34800
rect 27440 34734 27454 34786
rect 27506 34734 27520 34786
rect 27440 34720 27520 34734
rect 27600 34786 27680 34800
rect 27600 34734 27614 34786
rect 27666 34734 27680 34786
rect 27600 34720 27680 34734
rect 27760 34786 27840 34800
rect 27760 34734 27774 34786
rect 27826 34734 27840 34786
rect 27760 34720 27840 34734
rect 27920 34786 28000 34800
rect 27920 34734 27934 34786
rect 27986 34734 28000 34786
rect 27920 34720 28000 34734
rect 28080 34786 28160 34800
rect 28080 34734 28094 34786
rect 28146 34734 28160 34786
rect 28080 34720 28160 34734
rect 28240 34786 28320 34800
rect 28240 34734 28254 34786
rect 28306 34734 28320 34786
rect 28240 34720 28320 34734
rect 28400 34786 28480 34800
rect 28400 34734 28414 34786
rect 28466 34734 28480 34786
rect 28400 34720 28480 34734
rect 28560 34786 28640 34800
rect 28560 34734 28574 34786
rect 28626 34734 28640 34786
rect 28560 34720 28640 34734
rect 28720 34786 28800 34800
rect 28720 34734 28734 34786
rect 28786 34734 28800 34786
rect 28720 34720 28800 34734
rect 28880 34786 28960 34800
rect 28880 34734 28894 34786
rect 28946 34734 28960 34786
rect 28880 34720 28960 34734
rect 29040 34786 29120 34800
rect 29040 34734 29054 34786
rect 29106 34734 29120 34786
rect 29040 34720 29120 34734
rect 29200 34786 29280 34800
rect 29200 34734 29214 34786
rect 29266 34734 29280 34786
rect 29200 34720 29280 34734
rect 29360 34786 29440 34800
rect 29360 34734 29374 34786
rect 29426 34734 29440 34786
rect 29360 34720 29440 34734
rect 33520 34786 33600 34800
rect 33520 34734 33534 34786
rect 33586 34734 33600 34786
rect 33520 34720 33600 34734
rect 33680 34786 33760 34800
rect 33680 34734 33694 34786
rect 33746 34734 33760 34786
rect 33680 34720 33760 34734
rect 33840 34786 33920 34800
rect 33840 34734 33854 34786
rect 33906 34734 33920 34786
rect 33840 34720 33920 34734
rect 34000 34786 34080 34800
rect 34000 34734 34014 34786
rect 34066 34734 34080 34786
rect 34000 34720 34080 34734
rect 34160 34786 34240 34800
rect 34160 34734 34174 34786
rect 34226 34734 34240 34786
rect 34160 34720 34240 34734
rect 34320 34786 34400 34800
rect 34320 34734 34334 34786
rect 34386 34734 34400 34786
rect 34320 34720 34400 34734
rect 34480 34786 34560 34800
rect 34480 34734 34494 34786
rect 34546 34734 34560 34786
rect 34480 34720 34560 34734
rect 34640 34786 34720 34800
rect 34640 34734 34654 34786
rect 34706 34734 34720 34786
rect 34640 34720 34720 34734
rect 34800 34786 34880 34800
rect 34800 34734 34814 34786
rect 34866 34734 34880 34786
rect 34800 34720 34880 34734
rect 34960 34786 35040 34800
rect 34960 34734 34974 34786
rect 35026 34734 35040 34786
rect 34960 34720 35040 34734
rect 35120 34786 35200 34800
rect 35120 34734 35134 34786
rect 35186 34734 35200 34786
rect 35120 34720 35200 34734
rect 35280 34786 35360 34800
rect 35280 34734 35294 34786
rect 35346 34734 35360 34786
rect 35280 34720 35360 34734
rect 35440 34786 35520 34800
rect 35440 34734 35454 34786
rect 35506 34734 35520 34786
rect 35440 34720 35520 34734
rect 35600 34786 35680 34800
rect 35600 34734 35614 34786
rect 35666 34734 35680 34786
rect 35600 34720 35680 34734
rect 35760 34786 35840 34800
rect 35760 34734 35774 34786
rect 35826 34734 35840 34786
rect 35760 34720 35840 34734
rect 35920 34786 36000 34800
rect 35920 34734 35934 34786
rect 35986 34734 36000 34786
rect 35920 34720 36000 34734
rect 36080 34786 36160 34800
rect 36080 34734 36094 34786
rect 36146 34734 36160 34786
rect 36080 34720 36160 34734
rect 36240 34786 36320 34800
rect 36240 34734 36254 34786
rect 36306 34734 36320 34786
rect 36240 34720 36320 34734
rect 36400 34786 36480 34800
rect 36400 34734 36414 34786
rect 36466 34734 36480 34786
rect 36400 34720 36480 34734
rect 36560 34786 36640 34800
rect 36560 34734 36574 34786
rect 36626 34734 36640 34786
rect 36560 34720 36640 34734
rect 36720 34786 36800 34800
rect 36720 34734 36734 34786
rect 36786 34734 36800 34786
rect 36720 34720 36800 34734
rect 36880 34786 36960 34800
rect 36880 34734 36894 34786
rect 36946 34734 36960 34786
rect 36880 34720 36960 34734
rect 37040 34786 37120 34800
rect 37040 34734 37054 34786
rect 37106 34734 37120 34786
rect 37040 34720 37120 34734
rect 37200 34786 37280 34800
rect 37200 34734 37214 34786
rect 37266 34734 37280 34786
rect 37200 34720 37280 34734
rect 37360 34786 37440 34800
rect 37360 34734 37374 34786
rect 37426 34734 37440 34786
rect 37360 34720 37440 34734
rect 37520 34786 37600 34800
rect 37520 34734 37534 34786
rect 37586 34734 37600 34786
rect 37520 34720 37600 34734
rect 37680 34786 37760 34800
rect 37680 34734 37694 34786
rect 37746 34734 37760 34786
rect 37680 34720 37760 34734
rect 37840 34786 37920 34800
rect 37840 34734 37854 34786
rect 37906 34734 37920 34786
rect 37840 34720 37920 34734
rect 38000 34786 38080 34800
rect 38000 34734 38014 34786
rect 38066 34734 38080 34786
rect 38000 34720 38080 34734
rect 38160 34786 38240 34800
rect 38160 34734 38174 34786
rect 38226 34734 38240 34786
rect 38160 34720 38240 34734
rect 38320 34786 38400 34800
rect 38320 34734 38334 34786
rect 38386 34734 38400 34786
rect 38320 34720 38400 34734
rect 38480 34786 38560 34800
rect 38480 34734 38494 34786
rect 38546 34734 38560 34786
rect 38480 34720 38560 34734
rect 38640 34786 38720 34800
rect 38640 34734 38654 34786
rect 38706 34734 38720 34786
rect 38640 34720 38720 34734
rect 38800 34786 38880 34800
rect 38800 34734 38814 34786
rect 38866 34734 38880 34786
rect 38800 34720 38880 34734
rect 38960 34786 39040 34800
rect 38960 34734 38974 34786
rect 39026 34734 39040 34786
rect 38960 34720 39040 34734
rect 39120 34786 39200 34800
rect 39120 34734 39134 34786
rect 39186 34734 39200 34786
rect 39120 34720 39200 34734
rect 39280 34786 39360 34800
rect 39280 34734 39294 34786
rect 39346 34734 39360 34786
rect 39280 34720 39360 34734
rect 39440 34786 39520 34800
rect 39440 34734 39454 34786
rect 39506 34734 39520 34786
rect 39440 34720 39520 34734
rect 39600 34786 39680 34800
rect 39600 34734 39614 34786
rect 39666 34734 39680 34786
rect 39600 34720 39680 34734
rect 39760 34786 39840 34800
rect 39760 34734 39774 34786
rect 39826 34734 39840 34786
rect 39760 34720 39840 34734
rect 39920 34786 40000 34800
rect 39920 34734 39934 34786
rect 39986 34734 40000 34786
rect 39920 34720 40000 34734
rect 40080 34786 40160 34800
rect 40080 34734 40094 34786
rect 40146 34734 40160 34786
rect 40080 34720 40160 34734
rect 40240 34786 40320 34800
rect 40240 34734 40254 34786
rect 40306 34734 40320 34786
rect 40240 34720 40320 34734
rect 40400 34786 40480 34800
rect 40400 34734 40414 34786
rect 40466 34734 40480 34786
rect 40400 34720 40480 34734
rect 40560 34786 40640 34800
rect 40560 34734 40574 34786
rect 40626 34734 40640 34786
rect 40560 34720 40640 34734
rect 40720 34786 40800 34800
rect 40720 34734 40734 34786
rect 40786 34734 40800 34786
rect 40720 34720 40800 34734
rect 40880 34786 40960 34800
rect 40880 34734 40894 34786
rect 40946 34734 40960 34786
rect 40880 34720 40960 34734
rect 41040 34786 41120 34800
rect 41040 34734 41054 34786
rect 41106 34734 41120 34786
rect 41040 34720 41120 34734
rect 41200 34786 41280 34800
rect 41200 34734 41214 34786
rect 41266 34734 41280 34786
rect 41200 34720 41280 34734
rect 41360 34786 41440 34800
rect 41360 34734 41374 34786
rect 41426 34734 41440 34786
rect 41360 34720 41440 34734
rect 41520 34786 41600 34800
rect 41520 34734 41534 34786
rect 41586 34734 41600 34786
rect 41520 34720 41600 34734
rect 41680 34786 41760 34800
rect 41680 34734 41694 34786
rect 41746 34734 41760 34786
rect 41680 34720 41760 34734
rect 41840 34786 41920 34800
rect 41840 34734 41854 34786
rect 41906 34734 41920 34786
rect 41840 34720 41920 34734
rect 0 34466 80 34480
rect 0 34414 14 34466
rect 66 34414 80 34466
rect 0 34400 80 34414
rect 160 34466 240 34480
rect 160 34414 174 34466
rect 226 34414 240 34466
rect 160 34400 240 34414
rect 320 34466 400 34480
rect 320 34414 334 34466
rect 386 34414 400 34466
rect 320 34400 400 34414
rect 480 34466 560 34480
rect 480 34414 494 34466
rect 546 34414 560 34466
rect 480 34400 560 34414
rect 640 34466 720 34480
rect 640 34414 654 34466
rect 706 34414 720 34466
rect 640 34400 720 34414
rect 800 34466 880 34480
rect 800 34414 814 34466
rect 866 34414 880 34466
rect 800 34400 880 34414
rect 960 34466 1040 34480
rect 960 34414 974 34466
rect 1026 34414 1040 34466
rect 960 34400 1040 34414
rect 1120 34466 1200 34480
rect 1120 34414 1134 34466
rect 1186 34414 1200 34466
rect 1120 34400 1200 34414
rect 1280 34466 1360 34480
rect 1280 34414 1294 34466
rect 1346 34414 1360 34466
rect 1280 34400 1360 34414
rect 1440 34466 1520 34480
rect 1440 34414 1454 34466
rect 1506 34414 1520 34466
rect 1440 34400 1520 34414
rect 1600 34466 1680 34480
rect 1600 34414 1614 34466
rect 1666 34414 1680 34466
rect 1600 34400 1680 34414
rect 1760 34466 1840 34480
rect 1760 34414 1774 34466
rect 1826 34414 1840 34466
rect 1760 34400 1840 34414
rect 1920 34466 2000 34480
rect 1920 34414 1934 34466
rect 1986 34414 2000 34466
rect 1920 34400 2000 34414
rect 2080 34466 2160 34480
rect 2080 34414 2094 34466
rect 2146 34414 2160 34466
rect 2080 34400 2160 34414
rect 2240 34466 2320 34480
rect 2240 34414 2254 34466
rect 2306 34414 2320 34466
rect 2240 34400 2320 34414
rect 2400 34466 2480 34480
rect 2400 34414 2414 34466
rect 2466 34414 2480 34466
rect 2400 34400 2480 34414
rect 2560 34466 2640 34480
rect 2560 34414 2574 34466
rect 2626 34414 2640 34466
rect 2560 34400 2640 34414
rect 2720 34466 2800 34480
rect 2720 34414 2734 34466
rect 2786 34414 2800 34466
rect 2720 34400 2800 34414
rect 2880 34466 2960 34480
rect 2880 34414 2894 34466
rect 2946 34414 2960 34466
rect 2880 34400 2960 34414
rect 3040 34466 3120 34480
rect 3040 34414 3054 34466
rect 3106 34414 3120 34466
rect 3040 34400 3120 34414
rect 3200 34466 3280 34480
rect 3200 34414 3214 34466
rect 3266 34414 3280 34466
rect 3200 34400 3280 34414
rect 3360 34466 3440 34480
rect 3360 34414 3374 34466
rect 3426 34414 3440 34466
rect 3360 34400 3440 34414
rect 3520 34466 3600 34480
rect 3520 34414 3534 34466
rect 3586 34414 3600 34466
rect 3520 34400 3600 34414
rect 3680 34466 3760 34480
rect 3680 34414 3694 34466
rect 3746 34414 3760 34466
rect 3680 34400 3760 34414
rect 3840 34466 3920 34480
rect 3840 34414 3854 34466
rect 3906 34414 3920 34466
rect 3840 34400 3920 34414
rect 4000 34466 4080 34480
rect 4000 34414 4014 34466
rect 4066 34414 4080 34466
rect 4000 34400 4080 34414
rect 4160 34466 4240 34480
rect 4160 34414 4174 34466
rect 4226 34414 4240 34466
rect 4160 34400 4240 34414
rect 4320 34466 4400 34480
rect 4320 34414 4334 34466
rect 4386 34414 4400 34466
rect 4320 34400 4400 34414
rect 4480 34466 4560 34480
rect 4480 34414 4494 34466
rect 4546 34414 4560 34466
rect 4480 34400 4560 34414
rect 4640 34466 4720 34480
rect 4640 34414 4654 34466
rect 4706 34414 4720 34466
rect 4640 34400 4720 34414
rect 4800 34466 4880 34480
rect 4800 34414 4814 34466
rect 4866 34414 4880 34466
rect 4800 34400 4880 34414
rect 4960 34466 5040 34480
rect 4960 34414 4974 34466
rect 5026 34414 5040 34466
rect 4960 34400 5040 34414
rect 5120 34466 5200 34480
rect 5120 34414 5134 34466
rect 5186 34414 5200 34466
rect 5120 34400 5200 34414
rect 5280 34466 5360 34480
rect 5280 34414 5294 34466
rect 5346 34414 5360 34466
rect 5280 34400 5360 34414
rect 5440 34466 5520 34480
rect 5440 34414 5454 34466
rect 5506 34414 5520 34466
rect 5440 34400 5520 34414
rect 5600 34466 5680 34480
rect 5600 34414 5614 34466
rect 5666 34414 5680 34466
rect 5600 34400 5680 34414
rect 5760 34466 5840 34480
rect 5760 34414 5774 34466
rect 5826 34414 5840 34466
rect 5760 34400 5840 34414
rect 5920 34466 6000 34480
rect 5920 34414 5934 34466
rect 5986 34414 6000 34466
rect 5920 34400 6000 34414
rect 6080 34466 6160 34480
rect 6080 34414 6094 34466
rect 6146 34414 6160 34466
rect 6080 34400 6160 34414
rect 6240 34466 6320 34480
rect 6240 34414 6254 34466
rect 6306 34414 6320 34466
rect 6240 34400 6320 34414
rect 6400 34466 6480 34480
rect 6400 34414 6414 34466
rect 6466 34414 6480 34466
rect 6400 34400 6480 34414
rect 6560 34466 6640 34480
rect 6560 34414 6574 34466
rect 6626 34414 6640 34466
rect 6560 34400 6640 34414
rect 6720 34466 6800 34480
rect 6720 34414 6734 34466
rect 6786 34414 6800 34466
rect 6720 34400 6800 34414
rect 6880 34466 6960 34480
rect 6880 34414 6894 34466
rect 6946 34414 6960 34466
rect 6880 34400 6960 34414
rect 7040 34466 7120 34480
rect 7040 34414 7054 34466
rect 7106 34414 7120 34466
rect 7040 34400 7120 34414
rect 7200 34466 7280 34480
rect 7200 34414 7214 34466
rect 7266 34414 7280 34466
rect 7200 34400 7280 34414
rect 7360 34466 7440 34480
rect 7360 34414 7374 34466
rect 7426 34414 7440 34466
rect 7360 34400 7440 34414
rect 7520 34466 7600 34480
rect 7520 34414 7534 34466
rect 7586 34414 7600 34466
rect 7520 34400 7600 34414
rect 7680 34466 7760 34480
rect 7680 34414 7694 34466
rect 7746 34414 7760 34466
rect 7680 34400 7760 34414
rect 7840 34466 7920 34480
rect 7840 34414 7854 34466
rect 7906 34414 7920 34466
rect 7840 34400 7920 34414
rect 8000 34466 8080 34480
rect 8000 34414 8014 34466
rect 8066 34414 8080 34466
rect 8000 34400 8080 34414
rect 8160 34466 8240 34480
rect 8160 34414 8174 34466
rect 8226 34414 8240 34466
rect 8160 34400 8240 34414
rect 8320 34466 8400 34480
rect 8320 34414 8334 34466
rect 8386 34414 8400 34466
rect 8320 34400 8400 34414
rect 12480 34466 12560 34480
rect 12480 34414 12494 34466
rect 12546 34414 12560 34466
rect 12480 34400 12560 34414
rect 12640 34466 12720 34480
rect 12640 34414 12654 34466
rect 12706 34414 12720 34466
rect 12640 34400 12720 34414
rect 12800 34466 12880 34480
rect 12800 34414 12814 34466
rect 12866 34414 12880 34466
rect 12800 34400 12880 34414
rect 12960 34466 13040 34480
rect 12960 34414 12974 34466
rect 13026 34414 13040 34466
rect 12960 34400 13040 34414
rect 13120 34466 13200 34480
rect 13120 34414 13134 34466
rect 13186 34414 13200 34466
rect 13120 34400 13200 34414
rect 13280 34466 13360 34480
rect 13280 34414 13294 34466
rect 13346 34414 13360 34466
rect 13280 34400 13360 34414
rect 13440 34466 13520 34480
rect 13440 34414 13454 34466
rect 13506 34414 13520 34466
rect 13440 34400 13520 34414
rect 13600 34466 13680 34480
rect 13600 34414 13614 34466
rect 13666 34414 13680 34466
rect 13600 34400 13680 34414
rect 13760 34466 13840 34480
rect 13760 34414 13774 34466
rect 13826 34414 13840 34466
rect 13760 34400 13840 34414
rect 13920 34466 14000 34480
rect 13920 34414 13934 34466
rect 13986 34414 14000 34466
rect 13920 34400 14000 34414
rect 14080 34466 14160 34480
rect 14080 34414 14094 34466
rect 14146 34414 14160 34466
rect 14080 34400 14160 34414
rect 14240 34466 14320 34480
rect 14240 34414 14254 34466
rect 14306 34414 14320 34466
rect 14240 34400 14320 34414
rect 14400 34466 14480 34480
rect 14400 34414 14414 34466
rect 14466 34414 14480 34466
rect 14400 34400 14480 34414
rect 14560 34466 14640 34480
rect 14560 34414 14574 34466
rect 14626 34414 14640 34466
rect 14560 34400 14640 34414
rect 14720 34466 14800 34480
rect 14720 34414 14734 34466
rect 14786 34414 14800 34466
rect 14720 34400 14800 34414
rect 14880 34466 14960 34480
rect 14880 34414 14894 34466
rect 14946 34414 14960 34466
rect 14880 34400 14960 34414
rect 15040 34466 15120 34480
rect 15040 34414 15054 34466
rect 15106 34414 15120 34466
rect 15040 34400 15120 34414
rect 15200 34466 15280 34480
rect 15200 34414 15214 34466
rect 15266 34414 15280 34466
rect 15200 34400 15280 34414
rect 15360 34466 15440 34480
rect 15360 34414 15374 34466
rect 15426 34414 15440 34466
rect 15360 34400 15440 34414
rect 15520 34466 15600 34480
rect 15520 34414 15534 34466
rect 15586 34414 15600 34466
rect 15520 34400 15600 34414
rect 15680 34466 15760 34480
rect 15680 34414 15694 34466
rect 15746 34414 15760 34466
rect 15680 34400 15760 34414
rect 15840 34466 15920 34480
rect 15840 34414 15854 34466
rect 15906 34414 15920 34466
rect 15840 34400 15920 34414
rect 16000 34466 16080 34480
rect 16000 34414 16014 34466
rect 16066 34414 16080 34466
rect 16000 34400 16080 34414
rect 16160 34466 16240 34480
rect 16160 34414 16174 34466
rect 16226 34414 16240 34466
rect 16160 34400 16240 34414
rect 16320 34466 16400 34480
rect 16320 34414 16334 34466
rect 16386 34414 16400 34466
rect 16320 34400 16400 34414
rect 16480 34466 16560 34480
rect 16480 34414 16494 34466
rect 16546 34414 16560 34466
rect 16480 34400 16560 34414
rect 16640 34466 16720 34480
rect 16640 34414 16654 34466
rect 16706 34414 16720 34466
rect 16640 34400 16720 34414
rect 16800 34466 16880 34480
rect 16800 34414 16814 34466
rect 16866 34414 16880 34466
rect 16800 34400 16880 34414
rect 16960 34466 17040 34480
rect 16960 34414 16974 34466
rect 17026 34414 17040 34466
rect 16960 34400 17040 34414
rect 17120 34466 17200 34480
rect 17120 34414 17134 34466
rect 17186 34414 17200 34466
rect 17120 34400 17200 34414
rect 17280 34466 17360 34480
rect 17280 34414 17294 34466
rect 17346 34414 17360 34466
rect 17280 34400 17360 34414
rect 17440 34466 17520 34480
rect 17440 34414 17454 34466
rect 17506 34414 17520 34466
rect 17440 34400 17520 34414
rect 17600 34466 17680 34480
rect 17600 34414 17614 34466
rect 17666 34414 17680 34466
rect 17600 34400 17680 34414
rect 17760 34466 17840 34480
rect 17760 34414 17774 34466
rect 17826 34414 17840 34466
rect 17760 34400 17840 34414
rect 17920 34466 18000 34480
rect 17920 34414 17934 34466
rect 17986 34414 18000 34466
rect 17920 34400 18000 34414
rect 18080 34466 18160 34480
rect 18080 34414 18094 34466
rect 18146 34414 18160 34466
rect 18080 34400 18160 34414
rect 18240 34466 18320 34480
rect 18240 34414 18254 34466
rect 18306 34414 18320 34466
rect 18240 34400 18320 34414
rect 18400 34466 18480 34480
rect 18400 34414 18414 34466
rect 18466 34414 18480 34466
rect 18400 34400 18480 34414
rect 18560 34466 18640 34480
rect 18560 34414 18574 34466
rect 18626 34414 18640 34466
rect 18560 34400 18640 34414
rect 18720 34466 18800 34480
rect 18720 34414 18734 34466
rect 18786 34414 18800 34466
rect 18720 34400 18800 34414
rect 18880 34466 18960 34480
rect 18880 34414 18894 34466
rect 18946 34414 18960 34466
rect 18880 34400 18960 34414
rect 23120 34466 23200 34480
rect 23120 34414 23134 34466
rect 23186 34414 23200 34466
rect 23120 34400 23200 34414
rect 23280 34466 23360 34480
rect 23280 34414 23294 34466
rect 23346 34414 23360 34466
rect 23280 34400 23360 34414
rect 23440 34466 23520 34480
rect 23440 34414 23454 34466
rect 23506 34414 23520 34466
rect 23440 34400 23520 34414
rect 23600 34466 23680 34480
rect 23600 34414 23614 34466
rect 23666 34414 23680 34466
rect 23600 34400 23680 34414
rect 23760 34466 23840 34480
rect 23760 34414 23774 34466
rect 23826 34414 23840 34466
rect 23760 34400 23840 34414
rect 23920 34466 24000 34480
rect 23920 34414 23934 34466
rect 23986 34414 24000 34466
rect 23920 34400 24000 34414
rect 24080 34466 24160 34480
rect 24080 34414 24094 34466
rect 24146 34414 24160 34466
rect 24080 34400 24160 34414
rect 24240 34466 24320 34480
rect 24240 34414 24254 34466
rect 24306 34414 24320 34466
rect 24240 34400 24320 34414
rect 24400 34466 24480 34480
rect 24400 34414 24414 34466
rect 24466 34414 24480 34466
rect 24400 34400 24480 34414
rect 24560 34466 24640 34480
rect 24560 34414 24574 34466
rect 24626 34414 24640 34466
rect 24560 34400 24640 34414
rect 24720 34466 24800 34480
rect 24720 34414 24734 34466
rect 24786 34414 24800 34466
rect 24720 34400 24800 34414
rect 24880 34466 24960 34480
rect 24880 34414 24894 34466
rect 24946 34414 24960 34466
rect 24880 34400 24960 34414
rect 25040 34466 25120 34480
rect 25040 34414 25054 34466
rect 25106 34414 25120 34466
rect 25040 34400 25120 34414
rect 25200 34466 25280 34480
rect 25200 34414 25214 34466
rect 25266 34414 25280 34466
rect 25200 34400 25280 34414
rect 25360 34466 25440 34480
rect 25360 34414 25374 34466
rect 25426 34414 25440 34466
rect 25360 34400 25440 34414
rect 25520 34466 25600 34480
rect 25520 34414 25534 34466
rect 25586 34414 25600 34466
rect 25520 34400 25600 34414
rect 25680 34466 25760 34480
rect 25680 34414 25694 34466
rect 25746 34414 25760 34466
rect 25680 34400 25760 34414
rect 25840 34466 25920 34480
rect 25840 34414 25854 34466
rect 25906 34414 25920 34466
rect 25840 34400 25920 34414
rect 26000 34466 26080 34480
rect 26000 34414 26014 34466
rect 26066 34414 26080 34466
rect 26000 34400 26080 34414
rect 26160 34466 26240 34480
rect 26160 34414 26174 34466
rect 26226 34414 26240 34466
rect 26160 34400 26240 34414
rect 26320 34466 26400 34480
rect 26320 34414 26334 34466
rect 26386 34414 26400 34466
rect 26320 34400 26400 34414
rect 26480 34466 26560 34480
rect 26480 34414 26494 34466
rect 26546 34414 26560 34466
rect 26480 34400 26560 34414
rect 26640 34466 26720 34480
rect 26640 34414 26654 34466
rect 26706 34414 26720 34466
rect 26640 34400 26720 34414
rect 26800 34466 26880 34480
rect 26800 34414 26814 34466
rect 26866 34414 26880 34466
rect 26800 34400 26880 34414
rect 26960 34466 27040 34480
rect 26960 34414 26974 34466
rect 27026 34414 27040 34466
rect 26960 34400 27040 34414
rect 27120 34466 27200 34480
rect 27120 34414 27134 34466
rect 27186 34414 27200 34466
rect 27120 34400 27200 34414
rect 27280 34466 27360 34480
rect 27280 34414 27294 34466
rect 27346 34414 27360 34466
rect 27280 34400 27360 34414
rect 27440 34466 27520 34480
rect 27440 34414 27454 34466
rect 27506 34414 27520 34466
rect 27440 34400 27520 34414
rect 27600 34466 27680 34480
rect 27600 34414 27614 34466
rect 27666 34414 27680 34466
rect 27600 34400 27680 34414
rect 27760 34466 27840 34480
rect 27760 34414 27774 34466
rect 27826 34414 27840 34466
rect 27760 34400 27840 34414
rect 27920 34466 28000 34480
rect 27920 34414 27934 34466
rect 27986 34414 28000 34466
rect 27920 34400 28000 34414
rect 28080 34466 28160 34480
rect 28080 34414 28094 34466
rect 28146 34414 28160 34466
rect 28080 34400 28160 34414
rect 28240 34466 28320 34480
rect 28240 34414 28254 34466
rect 28306 34414 28320 34466
rect 28240 34400 28320 34414
rect 28400 34466 28480 34480
rect 28400 34414 28414 34466
rect 28466 34414 28480 34466
rect 28400 34400 28480 34414
rect 28560 34466 28640 34480
rect 28560 34414 28574 34466
rect 28626 34414 28640 34466
rect 28560 34400 28640 34414
rect 28720 34466 28800 34480
rect 28720 34414 28734 34466
rect 28786 34414 28800 34466
rect 28720 34400 28800 34414
rect 28880 34466 28960 34480
rect 28880 34414 28894 34466
rect 28946 34414 28960 34466
rect 28880 34400 28960 34414
rect 29040 34466 29120 34480
rect 29040 34414 29054 34466
rect 29106 34414 29120 34466
rect 29040 34400 29120 34414
rect 29200 34466 29280 34480
rect 29200 34414 29214 34466
rect 29266 34414 29280 34466
rect 29200 34400 29280 34414
rect 29360 34466 29440 34480
rect 29360 34414 29374 34466
rect 29426 34414 29440 34466
rect 29360 34400 29440 34414
rect 33520 34466 33600 34480
rect 33520 34414 33534 34466
rect 33586 34414 33600 34466
rect 33520 34400 33600 34414
rect 33680 34466 33760 34480
rect 33680 34414 33694 34466
rect 33746 34414 33760 34466
rect 33680 34400 33760 34414
rect 33840 34466 33920 34480
rect 33840 34414 33854 34466
rect 33906 34414 33920 34466
rect 33840 34400 33920 34414
rect 34000 34466 34080 34480
rect 34000 34414 34014 34466
rect 34066 34414 34080 34466
rect 34000 34400 34080 34414
rect 34160 34466 34240 34480
rect 34160 34414 34174 34466
rect 34226 34414 34240 34466
rect 34160 34400 34240 34414
rect 34320 34466 34400 34480
rect 34320 34414 34334 34466
rect 34386 34414 34400 34466
rect 34320 34400 34400 34414
rect 34480 34466 34560 34480
rect 34480 34414 34494 34466
rect 34546 34414 34560 34466
rect 34480 34400 34560 34414
rect 34640 34466 34720 34480
rect 34640 34414 34654 34466
rect 34706 34414 34720 34466
rect 34640 34400 34720 34414
rect 34800 34466 34880 34480
rect 34800 34414 34814 34466
rect 34866 34414 34880 34466
rect 34800 34400 34880 34414
rect 34960 34466 35040 34480
rect 34960 34414 34974 34466
rect 35026 34414 35040 34466
rect 34960 34400 35040 34414
rect 35120 34466 35200 34480
rect 35120 34414 35134 34466
rect 35186 34414 35200 34466
rect 35120 34400 35200 34414
rect 35280 34466 35360 34480
rect 35280 34414 35294 34466
rect 35346 34414 35360 34466
rect 35280 34400 35360 34414
rect 35440 34466 35520 34480
rect 35440 34414 35454 34466
rect 35506 34414 35520 34466
rect 35440 34400 35520 34414
rect 35600 34466 35680 34480
rect 35600 34414 35614 34466
rect 35666 34414 35680 34466
rect 35600 34400 35680 34414
rect 35760 34466 35840 34480
rect 35760 34414 35774 34466
rect 35826 34414 35840 34466
rect 35760 34400 35840 34414
rect 35920 34466 36000 34480
rect 35920 34414 35934 34466
rect 35986 34414 36000 34466
rect 35920 34400 36000 34414
rect 36080 34466 36160 34480
rect 36080 34414 36094 34466
rect 36146 34414 36160 34466
rect 36080 34400 36160 34414
rect 36240 34466 36320 34480
rect 36240 34414 36254 34466
rect 36306 34414 36320 34466
rect 36240 34400 36320 34414
rect 36400 34466 36480 34480
rect 36400 34414 36414 34466
rect 36466 34414 36480 34466
rect 36400 34400 36480 34414
rect 36560 34466 36640 34480
rect 36560 34414 36574 34466
rect 36626 34414 36640 34466
rect 36560 34400 36640 34414
rect 36720 34466 36800 34480
rect 36720 34414 36734 34466
rect 36786 34414 36800 34466
rect 36720 34400 36800 34414
rect 36880 34466 36960 34480
rect 36880 34414 36894 34466
rect 36946 34414 36960 34466
rect 36880 34400 36960 34414
rect 37040 34466 37120 34480
rect 37040 34414 37054 34466
rect 37106 34414 37120 34466
rect 37040 34400 37120 34414
rect 37200 34466 37280 34480
rect 37200 34414 37214 34466
rect 37266 34414 37280 34466
rect 37200 34400 37280 34414
rect 37360 34466 37440 34480
rect 37360 34414 37374 34466
rect 37426 34414 37440 34466
rect 37360 34400 37440 34414
rect 37520 34466 37600 34480
rect 37520 34414 37534 34466
rect 37586 34414 37600 34466
rect 37520 34400 37600 34414
rect 37680 34466 37760 34480
rect 37680 34414 37694 34466
rect 37746 34414 37760 34466
rect 37680 34400 37760 34414
rect 37840 34466 37920 34480
rect 37840 34414 37854 34466
rect 37906 34414 37920 34466
rect 37840 34400 37920 34414
rect 38000 34466 38080 34480
rect 38000 34414 38014 34466
rect 38066 34414 38080 34466
rect 38000 34400 38080 34414
rect 38160 34466 38240 34480
rect 38160 34414 38174 34466
rect 38226 34414 38240 34466
rect 38160 34400 38240 34414
rect 38320 34466 38400 34480
rect 38320 34414 38334 34466
rect 38386 34414 38400 34466
rect 38320 34400 38400 34414
rect 38480 34466 38560 34480
rect 38480 34414 38494 34466
rect 38546 34414 38560 34466
rect 38480 34400 38560 34414
rect 38640 34466 38720 34480
rect 38640 34414 38654 34466
rect 38706 34414 38720 34466
rect 38640 34400 38720 34414
rect 38800 34466 38880 34480
rect 38800 34414 38814 34466
rect 38866 34414 38880 34466
rect 38800 34400 38880 34414
rect 38960 34466 39040 34480
rect 38960 34414 38974 34466
rect 39026 34414 39040 34466
rect 38960 34400 39040 34414
rect 39120 34466 39200 34480
rect 39120 34414 39134 34466
rect 39186 34414 39200 34466
rect 39120 34400 39200 34414
rect 39280 34466 39360 34480
rect 39280 34414 39294 34466
rect 39346 34414 39360 34466
rect 39280 34400 39360 34414
rect 39440 34466 39520 34480
rect 39440 34414 39454 34466
rect 39506 34414 39520 34466
rect 39440 34400 39520 34414
rect 39600 34466 39680 34480
rect 39600 34414 39614 34466
rect 39666 34414 39680 34466
rect 39600 34400 39680 34414
rect 39760 34466 39840 34480
rect 39760 34414 39774 34466
rect 39826 34414 39840 34466
rect 39760 34400 39840 34414
rect 39920 34466 40000 34480
rect 39920 34414 39934 34466
rect 39986 34414 40000 34466
rect 39920 34400 40000 34414
rect 40080 34466 40160 34480
rect 40080 34414 40094 34466
rect 40146 34414 40160 34466
rect 40080 34400 40160 34414
rect 40240 34466 40320 34480
rect 40240 34414 40254 34466
rect 40306 34414 40320 34466
rect 40240 34400 40320 34414
rect 40400 34466 40480 34480
rect 40400 34414 40414 34466
rect 40466 34414 40480 34466
rect 40400 34400 40480 34414
rect 40560 34466 40640 34480
rect 40560 34414 40574 34466
rect 40626 34414 40640 34466
rect 40560 34400 40640 34414
rect 40720 34466 40800 34480
rect 40720 34414 40734 34466
rect 40786 34414 40800 34466
rect 40720 34400 40800 34414
rect 40880 34466 40960 34480
rect 40880 34414 40894 34466
rect 40946 34414 40960 34466
rect 40880 34400 40960 34414
rect 41040 34466 41120 34480
rect 41040 34414 41054 34466
rect 41106 34414 41120 34466
rect 41040 34400 41120 34414
rect 41200 34466 41280 34480
rect 41200 34414 41214 34466
rect 41266 34414 41280 34466
rect 41200 34400 41280 34414
rect 41360 34466 41440 34480
rect 41360 34414 41374 34466
rect 41426 34414 41440 34466
rect 41360 34400 41440 34414
rect 41520 34466 41600 34480
rect 41520 34414 41534 34466
rect 41586 34414 41600 34466
rect 41520 34400 41600 34414
rect 41680 34466 41760 34480
rect 41680 34414 41694 34466
rect 41746 34414 41760 34466
rect 41680 34400 41760 34414
rect 41840 34466 41920 34480
rect 41840 34414 41854 34466
rect 41906 34414 41920 34466
rect 41840 34400 41920 34414
rect 0 34306 80 34320
rect 0 34254 14 34306
rect 66 34254 80 34306
rect 0 34240 80 34254
rect 160 34306 240 34320
rect 160 34254 174 34306
rect 226 34254 240 34306
rect 160 34240 240 34254
rect 320 34306 400 34320
rect 320 34254 334 34306
rect 386 34254 400 34306
rect 320 34240 400 34254
rect 480 34306 560 34320
rect 480 34254 494 34306
rect 546 34254 560 34306
rect 480 34240 560 34254
rect 640 34306 720 34320
rect 640 34254 654 34306
rect 706 34254 720 34306
rect 640 34240 720 34254
rect 800 34306 880 34320
rect 800 34254 814 34306
rect 866 34254 880 34306
rect 800 34240 880 34254
rect 960 34306 1040 34320
rect 960 34254 974 34306
rect 1026 34254 1040 34306
rect 960 34240 1040 34254
rect 1120 34306 1200 34320
rect 1120 34254 1134 34306
rect 1186 34254 1200 34306
rect 1120 34240 1200 34254
rect 1280 34306 1360 34320
rect 1280 34254 1294 34306
rect 1346 34254 1360 34306
rect 1280 34240 1360 34254
rect 1440 34306 1520 34320
rect 1440 34254 1454 34306
rect 1506 34254 1520 34306
rect 1440 34240 1520 34254
rect 1600 34306 1680 34320
rect 1600 34254 1614 34306
rect 1666 34254 1680 34306
rect 1600 34240 1680 34254
rect 1760 34306 1840 34320
rect 1760 34254 1774 34306
rect 1826 34254 1840 34306
rect 1760 34240 1840 34254
rect 1920 34306 2000 34320
rect 1920 34254 1934 34306
rect 1986 34254 2000 34306
rect 1920 34240 2000 34254
rect 2080 34306 2160 34320
rect 2080 34254 2094 34306
rect 2146 34254 2160 34306
rect 2080 34240 2160 34254
rect 2240 34306 2320 34320
rect 2240 34254 2254 34306
rect 2306 34254 2320 34306
rect 2240 34240 2320 34254
rect 2400 34306 2480 34320
rect 2400 34254 2414 34306
rect 2466 34254 2480 34306
rect 2400 34240 2480 34254
rect 2560 34306 2640 34320
rect 2560 34254 2574 34306
rect 2626 34254 2640 34306
rect 2560 34240 2640 34254
rect 2720 34306 2800 34320
rect 2720 34254 2734 34306
rect 2786 34254 2800 34306
rect 2720 34240 2800 34254
rect 2880 34306 2960 34320
rect 2880 34254 2894 34306
rect 2946 34254 2960 34306
rect 2880 34240 2960 34254
rect 3040 34306 3120 34320
rect 3040 34254 3054 34306
rect 3106 34254 3120 34306
rect 3040 34240 3120 34254
rect 3200 34306 3280 34320
rect 3200 34254 3214 34306
rect 3266 34254 3280 34306
rect 3200 34240 3280 34254
rect 3360 34306 3440 34320
rect 3360 34254 3374 34306
rect 3426 34254 3440 34306
rect 3360 34240 3440 34254
rect 3520 34306 3600 34320
rect 3520 34254 3534 34306
rect 3586 34254 3600 34306
rect 3520 34240 3600 34254
rect 3680 34306 3760 34320
rect 3680 34254 3694 34306
rect 3746 34254 3760 34306
rect 3680 34240 3760 34254
rect 3840 34306 3920 34320
rect 3840 34254 3854 34306
rect 3906 34254 3920 34306
rect 3840 34240 3920 34254
rect 4000 34306 4080 34320
rect 4000 34254 4014 34306
rect 4066 34254 4080 34306
rect 4000 34240 4080 34254
rect 4160 34306 4240 34320
rect 4160 34254 4174 34306
rect 4226 34254 4240 34306
rect 4160 34240 4240 34254
rect 4320 34306 4400 34320
rect 4320 34254 4334 34306
rect 4386 34254 4400 34306
rect 4320 34240 4400 34254
rect 4480 34306 4560 34320
rect 4480 34254 4494 34306
rect 4546 34254 4560 34306
rect 4480 34240 4560 34254
rect 4640 34306 4720 34320
rect 4640 34254 4654 34306
rect 4706 34254 4720 34306
rect 4640 34240 4720 34254
rect 4800 34306 4880 34320
rect 4800 34254 4814 34306
rect 4866 34254 4880 34306
rect 4800 34240 4880 34254
rect 4960 34306 5040 34320
rect 4960 34254 4974 34306
rect 5026 34254 5040 34306
rect 4960 34240 5040 34254
rect 5120 34306 5200 34320
rect 5120 34254 5134 34306
rect 5186 34254 5200 34306
rect 5120 34240 5200 34254
rect 5280 34306 5360 34320
rect 5280 34254 5294 34306
rect 5346 34254 5360 34306
rect 5280 34240 5360 34254
rect 5440 34306 5520 34320
rect 5440 34254 5454 34306
rect 5506 34254 5520 34306
rect 5440 34240 5520 34254
rect 5600 34306 5680 34320
rect 5600 34254 5614 34306
rect 5666 34254 5680 34306
rect 5600 34240 5680 34254
rect 5760 34306 5840 34320
rect 5760 34254 5774 34306
rect 5826 34254 5840 34306
rect 5760 34240 5840 34254
rect 5920 34306 6000 34320
rect 5920 34254 5934 34306
rect 5986 34254 6000 34306
rect 5920 34240 6000 34254
rect 6080 34306 6160 34320
rect 6080 34254 6094 34306
rect 6146 34254 6160 34306
rect 6080 34240 6160 34254
rect 6240 34306 6320 34320
rect 6240 34254 6254 34306
rect 6306 34254 6320 34306
rect 6240 34240 6320 34254
rect 6400 34306 6480 34320
rect 6400 34254 6414 34306
rect 6466 34254 6480 34306
rect 6400 34240 6480 34254
rect 6560 34306 6640 34320
rect 6560 34254 6574 34306
rect 6626 34254 6640 34306
rect 6560 34240 6640 34254
rect 6720 34306 6800 34320
rect 6720 34254 6734 34306
rect 6786 34254 6800 34306
rect 6720 34240 6800 34254
rect 6880 34306 6960 34320
rect 6880 34254 6894 34306
rect 6946 34254 6960 34306
rect 6880 34240 6960 34254
rect 7040 34306 7120 34320
rect 7040 34254 7054 34306
rect 7106 34254 7120 34306
rect 7040 34240 7120 34254
rect 7200 34306 7280 34320
rect 7200 34254 7214 34306
rect 7266 34254 7280 34306
rect 7200 34240 7280 34254
rect 7360 34306 7440 34320
rect 7360 34254 7374 34306
rect 7426 34254 7440 34306
rect 7360 34240 7440 34254
rect 7520 34306 7600 34320
rect 7520 34254 7534 34306
rect 7586 34254 7600 34306
rect 7520 34240 7600 34254
rect 7680 34306 7760 34320
rect 7680 34254 7694 34306
rect 7746 34254 7760 34306
rect 7680 34240 7760 34254
rect 7840 34306 7920 34320
rect 7840 34254 7854 34306
rect 7906 34254 7920 34306
rect 7840 34240 7920 34254
rect 8000 34306 8080 34320
rect 8000 34254 8014 34306
rect 8066 34254 8080 34306
rect 8000 34240 8080 34254
rect 8160 34306 8240 34320
rect 8160 34254 8174 34306
rect 8226 34254 8240 34306
rect 8160 34240 8240 34254
rect 8320 34306 8400 34320
rect 8320 34254 8334 34306
rect 8386 34254 8400 34306
rect 8320 34240 8400 34254
rect 12480 34306 12560 34320
rect 12480 34254 12494 34306
rect 12546 34254 12560 34306
rect 12480 34240 12560 34254
rect 12640 34306 12720 34320
rect 12640 34254 12654 34306
rect 12706 34254 12720 34306
rect 12640 34240 12720 34254
rect 12800 34306 12880 34320
rect 12800 34254 12814 34306
rect 12866 34254 12880 34306
rect 12800 34240 12880 34254
rect 12960 34306 13040 34320
rect 12960 34254 12974 34306
rect 13026 34254 13040 34306
rect 12960 34240 13040 34254
rect 13120 34306 13200 34320
rect 13120 34254 13134 34306
rect 13186 34254 13200 34306
rect 13120 34240 13200 34254
rect 13280 34306 13360 34320
rect 13280 34254 13294 34306
rect 13346 34254 13360 34306
rect 13280 34240 13360 34254
rect 13440 34306 13520 34320
rect 13440 34254 13454 34306
rect 13506 34254 13520 34306
rect 13440 34240 13520 34254
rect 13600 34306 13680 34320
rect 13600 34254 13614 34306
rect 13666 34254 13680 34306
rect 13600 34240 13680 34254
rect 13760 34306 13840 34320
rect 13760 34254 13774 34306
rect 13826 34254 13840 34306
rect 13760 34240 13840 34254
rect 13920 34306 14000 34320
rect 13920 34254 13934 34306
rect 13986 34254 14000 34306
rect 13920 34240 14000 34254
rect 14080 34306 14160 34320
rect 14080 34254 14094 34306
rect 14146 34254 14160 34306
rect 14080 34240 14160 34254
rect 14240 34306 14320 34320
rect 14240 34254 14254 34306
rect 14306 34254 14320 34306
rect 14240 34240 14320 34254
rect 14400 34306 14480 34320
rect 14400 34254 14414 34306
rect 14466 34254 14480 34306
rect 14400 34240 14480 34254
rect 14560 34306 14640 34320
rect 14560 34254 14574 34306
rect 14626 34254 14640 34306
rect 14560 34240 14640 34254
rect 14720 34306 14800 34320
rect 14720 34254 14734 34306
rect 14786 34254 14800 34306
rect 14720 34240 14800 34254
rect 14880 34306 14960 34320
rect 14880 34254 14894 34306
rect 14946 34254 14960 34306
rect 14880 34240 14960 34254
rect 15040 34306 15120 34320
rect 15040 34254 15054 34306
rect 15106 34254 15120 34306
rect 15040 34240 15120 34254
rect 15200 34306 15280 34320
rect 15200 34254 15214 34306
rect 15266 34254 15280 34306
rect 15200 34240 15280 34254
rect 15360 34306 15440 34320
rect 15360 34254 15374 34306
rect 15426 34254 15440 34306
rect 15360 34240 15440 34254
rect 15520 34306 15600 34320
rect 15520 34254 15534 34306
rect 15586 34254 15600 34306
rect 15520 34240 15600 34254
rect 15680 34306 15760 34320
rect 15680 34254 15694 34306
rect 15746 34254 15760 34306
rect 15680 34240 15760 34254
rect 15840 34306 15920 34320
rect 15840 34254 15854 34306
rect 15906 34254 15920 34306
rect 15840 34240 15920 34254
rect 16000 34306 16080 34320
rect 16000 34254 16014 34306
rect 16066 34254 16080 34306
rect 16000 34240 16080 34254
rect 16160 34306 16240 34320
rect 16160 34254 16174 34306
rect 16226 34254 16240 34306
rect 16160 34240 16240 34254
rect 16320 34306 16400 34320
rect 16320 34254 16334 34306
rect 16386 34254 16400 34306
rect 16320 34240 16400 34254
rect 16480 34306 16560 34320
rect 16480 34254 16494 34306
rect 16546 34254 16560 34306
rect 16480 34240 16560 34254
rect 16640 34306 16720 34320
rect 16640 34254 16654 34306
rect 16706 34254 16720 34306
rect 16640 34240 16720 34254
rect 16800 34306 16880 34320
rect 16800 34254 16814 34306
rect 16866 34254 16880 34306
rect 16800 34240 16880 34254
rect 16960 34306 17040 34320
rect 16960 34254 16974 34306
rect 17026 34254 17040 34306
rect 16960 34240 17040 34254
rect 17120 34306 17200 34320
rect 17120 34254 17134 34306
rect 17186 34254 17200 34306
rect 17120 34240 17200 34254
rect 17280 34306 17360 34320
rect 17280 34254 17294 34306
rect 17346 34254 17360 34306
rect 17280 34240 17360 34254
rect 17440 34306 17520 34320
rect 17440 34254 17454 34306
rect 17506 34254 17520 34306
rect 17440 34240 17520 34254
rect 17600 34306 17680 34320
rect 17600 34254 17614 34306
rect 17666 34254 17680 34306
rect 17600 34240 17680 34254
rect 17760 34306 17840 34320
rect 17760 34254 17774 34306
rect 17826 34254 17840 34306
rect 17760 34240 17840 34254
rect 17920 34306 18000 34320
rect 17920 34254 17934 34306
rect 17986 34254 18000 34306
rect 17920 34240 18000 34254
rect 18080 34306 18160 34320
rect 18080 34254 18094 34306
rect 18146 34254 18160 34306
rect 18080 34240 18160 34254
rect 18240 34306 18320 34320
rect 18240 34254 18254 34306
rect 18306 34254 18320 34306
rect 18240 34240 18320 34254
rect 18400 34306 18480 34320
rect 18400 34254 18414 34306
rect 18466 34254 18480 34306
rect 18400 34240 18480 34254
rect 18560 34306 18640 34320
rect 18560 34254 18574 34306
rect 18626 34254 18640 34306
rect 18560 34240 18640 34254
rect 18720 34306 18800 34320
rect 18720 34254 18734 34306
rect 18786 34254 18800 34306
rect 18720 34240 18800 34254
rect 18880 34306 18960 34320
rect 18880 34254 18894 34306
rect 18946 34254 18960 34306
rect 18880 34240 18960 34254
rect 23120 34306 23200 34320
rect 23120 34254 23134 34306
rect 23186 34254 23200 34306
rect 23120 34240 23200 34254
rect 23280 34306 23360 34320
rect 23280 34254 23294 34306
rect 23346 34254 23360 34306
rect 23280 34240 23360 34254
rect 23440 34306 23520 34320
rect 23440 34254 23454 34306
rect 23506 34254 23520 34306
rect 23440 34240 23520 34254
rect 23600 34306 23680 34320
rect 23600 34254 23614 34306
rect 23666 34254 23680 34306
rect 23600 34240 23680 34254
rect 23760 34306 23840 34320
rect 23760 34254 23774 34306
rect 23826 34254 23840 34306
rect 23760 34240 23840 34254
rect 23920 34306 24000 34320
rect 23920 34254 23934 34306
rect 23986 34254 24000 34306
rect 23920 34240 24000 34254
rect 24080 34306 24160 34320
rect 24080 34254 24094 34306
rect 24146 34254 24160 34306
rect 24080 34240 24160 34254
rect 24240 34306 24320 34320
rect 24240 34254 24254 34306
rect 24306 34254 24320 34306
rect 24240 34240 24320 34254
rect 24400 34306 24480 34320
rect 24400 34254 24414 34306
rect 24466 34254 24480 34306
rect 24400 34240 24480 34254
rect 24560 34306 24640 34320
rect 24560 34254 24574 34306
rect 24626 34254 24640 34306
rect 24560 34240 24640 34254
rect 24720 34306 24800 34320
rect 24720 34254 24734 34306
rect 24786 34254 24800 34306
rect 24720 34240 24800 34254
rect 24880 34306 24960 34320
rect 24880 34254 24894 34306
rect 24946 34254 24960 34306
rect 24880 34240 24960 34254
rect 25040 34306 25120 34320
rect 25040 34254 25054 34306
rect 25106 34254 25120 34306
rect 25040 34240 25120 34254
rect 25200 34306 25280 34320
rect 25200 34254 25214 34306
rect 25266 34254 25280 34306
rect 25200 34240 25280 34254
rect 25360 34306 25440 34320
rect 25360 34254 25374 34306
rect 25426 34254 25440 34306
rect 25360 34240 25440 34254
rect 25520 34306 25600 34320
rect 25520 34254 25534 34306
rect 25586 34254 25600 34306
rect 25520 34240 25600 34254
rect 25680 34306 25760 34320
rect 25680 34254 25694 34306
rect 25746 34254 25760 34306
rect 25680 34240 25760 34254
rect 25840 34306 25920 34320
rect 25840 34254 25854 34306
rect 25906 34254 25920 34306
rect 25840 34240 25920 34254
rect 26000 34306 26080 34320
rect 26000 34254 26014 34306
rect 26066 34254 26080 34306
rect 26000 34240 26080 34254
rect 26160 34306 26240 34320
rect 26160 34254 26174 34306
rect 26226 34254 26240 34306
rect 26160 34240 26240 34254
rect 26320 34306 26400 34320
rect 26320 34254 26334 34306
rect 26386 34254 26400 34306
rect 26320 34240 26400 34254
rect 26480 34306 26560 34320
rect 26480 34254 26494 34306
rect 26546 34254 26560 34306
rect 26480 34240 26560 34254
rect 26640 34306 26720 34320
rect 26640 34254 26654 34306
rect 26706 34254 26720 34306
rect 26640 34240 26720 34254
rect 26800 34306 26880 34320
rect 26800 34254 26814 34306
rect 26866 34254 26880 34306
rect 26800 34240 26880 34254
rect 26960 34306 27040 34320
rect 26960 34254 26974 34306
rect 27026 34254 27040 34306
rect 26960 34240 27040 34254
rect 27120 34306 27200 34320
rect 27120 34254 27134 34306
rect 27186 34254 27200 34306
rect 27120 34240 27200 34254
rect 27280 34306 27360 34320
rect 27280 34254 27294 34306
rect 27346 34254 27360 34306
rect 27280 34240 27360 34254
rect 27440 34306 27520 34320
rect 27440 34254 27454 34306
rect 27506 34254 27520 34306
rect 27440 34240 27520 34254
rect 27600 34306 27680 34320
rect 27600 34254 27614 34306
rect 27666 34254 27680 34306
rect 27600 34240 27680 34254
rect 27760 34306 27840 34320
rect 27760 34254 27774 34306
rect 27826 34254 27840 34306
rect 27760 34240 27840 34254
rect 27920 34306 28000 34320
rect 27920 34254 27934 34306
rect 27986 34254 28000 34306
rect 27920 34240 28000 34254
rect 28080 34306 28160 34320
rect 28080 34254 28094 34306
rect 28146 34254 28160 34306
rect 28080 34240 28160 34254
rect 28240 34306 28320 34320
rect 28240 34254 28254 34306
rect 28306 34254 28320 34306
rect 28240 34240 28320 34254
rect 28400 34306 28480 34320
rect 28400 34254 28414 34306
rect 28466 34254 28480 34306
rect 28400 34240 28480 34254
rect 28560 34306 28640 34320
rect 28560 34254 28574 34306
rect 28626 34254 28640 34306
rect 28560 34240 28640 34254
rect 28720 34306 28800 34320
rect 28720 34254 28734 34306
rect 28786 34254 28800 34306
rect 28720 34240 28800 34254
rect 28880 34306 28960 34320
rect 28880 34254 28894 34306
rect 28946 34254 28960 34306
rect 28880 34240 28960 34254
rect 29040 34306 29120 34320
rect 29040 34254 29054 34306
rect 29106 34254 29120 34306
rect 29040 34240 29120 34254
rect 29200 34306 29280 34320
rect 29200 34254 29214 34306
rect 29266 34254 29280 34306
rect 29200 34240 29280 34254
rect 29360 34306 29440 34320
rect 29360 34254 29374 34306
rect 29426 34254 29440 34306
rect 29360 34240 29440 34254
rect 33520 34306 33600 34320
rect 33520 34254 33534 34306
rect 33586 34254 33600 34306
rect 33520 34240 33600 34254
rect 33680 34306 33760 34320
rect 33680 34254 33694 34306
rect 33746 34254 33760 34306
rect 33680 34240 33760 34254
rect 33840 34306 33920 34320
rect 33840 34254 33854 34306
rect 33906 34254 33920 34306
rect 33840 34240 33920 34254
rect 34000 34306 34080 34320
rect 34000 34254 34014 34306
rect 34066 34254 34080 34306
rect 34000 34240 34080 34254
rect 34160 34306 34240 34320
rect 34160 34254 34174 34306
rect 34226 34254 34240 34306
rect 34160 34240 34240 34254
rect 34320 34306 34400 34320
rect 34320 34254 34334 34306
rect 34386 34254 34400 34306
rect 34320 34240 34400 34254
rect 34480 34306 34560 34320
rect 34480 34254 34494 34306
rect 34546 34254 34560 34306
rect 34480 34240 34560 34254
rect 34640 34306 34720 34320
rect 34640 34254 34654 34306
rect 34706 34254 34720 34306
rect 34640 34240 34720 34254
rect 34800 34306 34880 34320
rect 34800 34254 34814 34306
rect 34866 34254 34880 34306
rect 34800 34240 34880 34254
rect 34960 34306 35040 34320
rect 34960 34254 34974 34306
rect 35026 34254 35040 34306
rect 34960 34240 35040 34254
rect 35120 34306 35200 34320
rect 35120 34254 35134 34306
rect 35186 34254 35200 34306
rect 35120 34240 35200 34254
rect 35280 34306 35360 34320
rect 35280 34254 35294 34306
rect 35346 34254 35360 34306
rect 35280 34240 35360 34254
rect 35440 34306 35520 34320
rect 35440 34254 35454 34306
rect 35506 34254 35520 34306
rect 35440 34240 35520 34254
rect 35600 34306 35680 34320
rect 35600 34254 35614 34306
rect 35666 34254 35680 34306
rect 35600 34240 35680 34254
rect 35760 34306 35840 34320
rect 35760 34254 35774 34306
rect 35826 34254 35840 34306
rect 35760 34240 35840 34254
rect 35920 34306 36000 34320
rect 35920 34254 35934 34306
rect 35986 34254 36000 34306
rect 35920 34240 36000 34254
rect 36080 34306 36160 34320
rect 36080 34254 36094 34306
rect 36146 34254 36160 34306
rect 36080 34240 36160 34254
rect 36240 34306 36320 34320
rect 36240 34254 36254 34306
rect 36306 34254 36320 34306
rect 36240 34240 36320 34254
rect 36400 34306 36480 34320
rect 36400 34254 36414 34306
rect 36466 34254 36480 34306
rect 36400 34240 36480 34254
rect 36560 34306 36640 34320
rect 36560 34254 36574 34306
rect 36626 34254 36640 34306
rect 36560 34240 36640 34254
rect 36720 34306 36800 34320
rect 36720 34254 36734 34306
rect 36786 34254 36800 34306
rect 36720 34240 36800 34254
rect 36880 34306 36960 34320
rect 36880 34254 36894 34306
rect 36946 34254 36960 34306
rect 36880 34240 36960 34254
rect 37040 34306 37120 34320
rect 37040 34254 37054 34306
rect 37106 34254 37120 34306
rect 37040 34240 37120 34254
rect 37200 34306 37280 34320
rect 37200 34254 37214 34306
rect 37266 34254 37280 34306
rect 37200 34240 37280 34254
rect 37360 34306 37440 34320
rect 37360 34254 37374 34306
rect 37426 34254 37440 34306
rect 37360 34240 37440 34254
rect 37520 34306 37600 34320
rect 37520 34254 37534 34306
rect 37586 34254 37600 34306
rect 37520 34240 37600 34254
rect 37680 34306 37760 34320
rect 37680 34254 37694 34306
rect 37746 34254 37760 34306
rect 37680 34240 37760 34254
rect 37840 34306 37920 34320
rect 37840 34254 37854 34306
rect 37906 34254 37920 34306
rect 37840 34240 37920 34254
rect 38000 34306 38080 34320
rect 38000 34254 38014 34306
rect 38066 34254 38080 34306
rect 38000 34240 38080 34254
rect 38160 34306 38240 34320
rect 38160 34254 38174 34306
rect 38226 34254 38240 34306
rect 38160 34240 38240 34254
rect 38320 34306 38400 34320
rect 38320 34254 38334 34306
rect 38386 34254 38400 34306
rect 38320 34240 38400 34254
rect 38480 34306 38560 34320
rect 38480 34254 38494 34306
rect 38546 34254 38560 34306
rect 38480 34240 38560 34254
rect 38640 34306 38720 34320
rect 38640 34254 38654 34306
rect 38706 34254 38720 34306
rect 38640 34240 38720 34254
rect 38800 34306 38880 34320
rect 38800 34254 38814 34306
rect 38866 34254 38880 34306
rect 38800 34240 38880 34254
rect 38960 34306 39040 34320
rect 38960 34254 38974 34306
rect 39026 34254 39040 34306
rect 38960 34240 39040 34254
rect 39120 34306 39200 34320
rect 39120 34254 39134 34306
rect 39186 34254 39200 34306
rect 39120 34240 39200 34254
rect 39280 34306 39360 34320
rect 39280 34254 39294 34306
rect 39346 34254 39360 34306
rect 39280 34240 39360 34254
rect 39440 34306 39520 34320
rect 39440 34254 39454 34306
rect 39506 34254 39520 34306
rect 39440 34240 39520 34254
rect 39600 34306 39680 34320
rect 39600 34254 39614 34306
rect 39666 34254 39680 34306
rect 39600 34240 39680 34254
rect 39760 34306 39840 34320
rect 39760 34254 39774 34306
rect 39826 34254 39840 34306
rect 39760 34240 39840 34254
rect 39920 34306 40000 34320
rect 39920 34254 39934 34306
rect 39986 34254 40000 34306
rect 39920 34240 40000 34254
rect 40080 34306 40160 34320
rect 40080 34254 40094 34306
rect 40146 34254 40160 34306
rect 40080 34240 40160 34254
rect 40240 34306 40320 34320
rect 40240 34254 40254 34306
rect 40306 34254 40320 34306
rect 40240 34240 40320 34254
rect 40400 34306 40480 34320
rect 40400 34254 40414 34306
rect 40466 34254 40480 34306
rect 40400 34240 40480 34254
rect 40560 34306 40640 34320
rect 40560 34254 40574 34306
rect 40626 34254 40640 34306
rect 40560 34240 40640 34254
rect 40720 34306 40800 34320
rect 40720 34254 40734 34306
rect 40786 34254 40800 34306
rect 40720 34240 40800 34254
rect 40880 34306 40960 34320
rect 40880 34254 40894 34306
rect 40946 34254 40960 34306
rect 40880 34240 40960 34254
rect 41040 34306 41120 34320
rect 41040 34254 41054 34306
rect 41106 34254 41120 34306
rect 41040 34240 41120 34254
rect 41200 34306 41280 34320
rect 41200 34254 41214 34306
rect 41266 34254 41280 34306
rect 41200 34240 41280 34254
rect 41360 34306 41440 34320
rect 41360 34254 41374 34306
rect 41426 34254 41440 34306
rect 41360 34240 41440 34254
rect 41520 34306 41600 34320
rect 41520 34254 41534 34306
rect 41586 34254 41600 34306
rect 41520 34240 41600 34254
rect 41680 34306 41760 34320
rect 41680 34254 41694 34306
rect 41746 34254 41760 34306
rect 41680 34240 41760 34254
rect 41840 34306 41920 34320
rect 41840 34254 41854 34306
rect 41906 34254 41920 34306
rect 41840 34240 41920 34254
rect 0 33986 80 34000
rect 0 33934 14 33986
rect 66 33934 80 33986
rect 0 33920 80 33934
rect 160 33986 240 34000
rect 160 33934 174 33986
rect 226 33934 240 33986
rect 160 33920 240 33934
rect 320 33986 400 34000
rect 320 33934 334 33986
rect 386 33934 400 33986
rect 320 33920 400 33934
rect 480 33986 560 34000
rect 480 33934 494 33986
rect 546 33934 560 33986
rect 480 33920 560 33934
rect 640 33986 720 34000
rect 640 33934 654 33986
rect 706 33934 720 33986
rect 640 33920 720 33934
rect 800 33986 880 34000
rect 800 33934 814 33986
rect 866 33934 880 33986
rect 800 33920 880 33934
rect 960 33986 1040 34000
rect 960 33934 974 33986
rect 1026 33934 1040 33986
rect 960 33920 1040 33934
rect 1120 33986 1200 34000
rect 1120 33934 1134 33986
rect 1186 33934 1200 33986
rect 1120 33920 1200 33934
rect 1280 33986 1360 34000
rect 1280 33934 1294 33986
rect 1346 33934 1360 33986
rect 1280 33920 1360 33934
rect 1440 33986 1520 34000
rect 1440 33934 1454 33986
rect 1506 33934 1520 33986
rect 1440 33920 1520 33934
rect 1600 33986 1680 34000
rect 1600 33934 1614 33986
rect 1666 33934 1680 33986
rect 1600 33920 1680 33934
rect 1760 33986 1840 34000
rect 1760 33934 1774 33986
rect 1826 33934 1840 33986
rect 1760 33920 1840 33934
rect 1920 33986 2000 34000
rect 1920 33934 1934 33986
rect 1986 33934 2000 33986
rect 1920 33920 2000 33934
rect 2080 33986 2160 34000
rect 2080 33934 2094 33986
rect 2146 33934 2160 33986
rect 2080 33920 2160 33934
rect 2240 33986 2320 34000
rect 2240 33934 2254 33986
rect 2306 33934 2320 33986
rect 2240 33920 2320 33934
rect 2400 33986 2480 34000
rect 2400 33934 2414 33986
rect 2466 33934 2480 33986
rect 2400 33920 2480 33934
rect 2560 33986 2640 34000
rect 2560 33934 2574 33986
rect 2626 33934 2640 33986
rect 2560 33920 2640 33934
rect 2720 33986 2800 34000
rect 2720 33934 2734 33986
rect 2786 33934 2800 33986
rect 2720 33920 2800 33934
rect 2880 33986 2960 34000
rect 2880 33934 2894 33986
rect 2946 33934 2960 33986
rect 2880 33920 2960 33934
rect 3040 33986 3120 34000
rect 3040 33934 3054 33986
rect 3106 33934 3120 33986
rect 3040 33920 3120 33934
rect 3200 33986 3280 34000
rect 3200 33934 3214 33986
rect 3266 33934 3280 33986
rect 3200 33920 3280 33934
rect 3360 33986 3440 34000
rect 3360 33934 3374 33986
rect 3426 33934 3440 33986
rect 3360 33920 3440 33934
rect 3520 33986 3600 34000
rect 3520 33934 3534 33986
rect 3586 33934 3600 33986
rect 3520 33920 3600 33934
rect 3680 33986 3760 34000
rect 3680 33934 3694 33986
rect 3746 33934 3760 33986
rect 3680 33920 3760 33934
rect 3840 33986 3920 34000
rect 3840 33934 3854 33986
rect 3906 33934 3920 33986
rect 3840 33920 3920 33934
rect 4000 33986 4080 34000
rect 4000 33934 4014 33986
rect 4066 33934 4080 33986
rect 4000 33920 4080 33934
rect 4160 33986 4240 34000
rect 4160 33934 4174 33986
rect 4226 33934 4240 33986
rect 4160 33920 4240 33934
rect 4320 33986 4400 34000
rect 4320 33934 4334 33986
rect 4386 33934 4400 33986
rect 4320 33920 4400 33934
rect 4480 33986 4560 34000
rect 4480 33934 4494 33986
rect 4546 33934 4560 33986
rect 4480 33920 4560 33934
rect 4640 33986 4720 34000
rect 4640 33934 4654 33986
rect 4706 33934 4720 33986
rect 4640 33920 4720 33934
rect 4800 33986 4880 34000
rect 4800 33934 4814 33986
rect 4866 33934 4880 33986
rect 4800 33920 4880 33934
rect 4960 33986 5040 34000
rect 4960 33934 4974 33986
rect 5026 33934 5040 33986
rect 4960 33920 5040 33934
rect 5120 33986 5200 34000
rect 5120 33934 5134 33986
rect 5186 33934 5200 33986
rect 5120 33920 5200 33934
rect 5280 33986 5360 34000
rect 5280 33934 5294 33986
rect 5346 33934 5360 33986
rect 5280 33920 5360 33934
rect 5440 33986 5520 34000
rect 5440 33934 5454 33986
rect 5506 33934 5520 33986
rect 5440 33920 5520 33934
rect 5600 33986 5680 34000
rect 5600 33934 5614 33986
rect 5666 33934 5680 33986
rect 5600 33920 5680 33934
rect 5760 33986 5840 34000
rect 5760 33934 5774 33986
rect 5826 33934 5840 33986
rect 5760 33920 5840 33934
rect 5920 33986 6000 34000
rect 5920 33934 5934 33986
rect 5986 33934 6000 33986
rect 5920 33920 6000 33934
rect 6080 33986 6160 34000
rect 6080 33934 6094 33986
rect 6146 33934 6160 33986
rect 6080 33920 6160 33934
rect 6240 33986 6320 34000
rect 6240 33934 6254 33986
rect 6306 33934 6320 33986
rect 6240 33920 6320 33934
rect 6400 33986 6480 34000
rect 6400 33934 6414 33986
rect 6466 33934 6480 33986
rect 6400 33920 6480 33934
rect 6560 33986 6640 34000
rect 6560 33934 6574 33986
rect 6626 33934 6640 33986
rect 6560 33920 6640 33934
rect 6720 33986 6800 34000
rect 6720 33934 6734 33986
rect 6786 33934 6800 33986
rect 6720 33920 6800 33934
rect 6880 33986 6960 34000
rect 6880 33934 6894 33986
rect 6946 33934 6960 33986
rect 6880 33920 6960 33934
rect 7040 33986 7120 34000
rect 7040 33934 7054 33986
rect 7106 33934 7120 33986
rect 7040 33920 7120 33934
rect 7200 33986 7280 34000
rect 7200 33934 7214 33986
rect 7266 33934 7280 33986
rect 7200 33920 7280 33934
rect 7360 33986 7440 34000
rect 7360 33934 7374 33986
rect 7426 33934 7440 33986
rect 7360 33920 7440 33934
rect 7520 33986 7600 34000
rect 7520 33934 7534 33986
rect 7586 33934 7600 33986
rect 7520 33920 7600 33934
rect 7680 33986 7760 34000
rect 7680 33934 7694 33986
rect 7746 33934 7760 33986
rect 7680 33920 7760 33934
rect 7840 33986 7920 34000
rect 7840 33934 7854 33986
rect 7906 33934 7920 33986
rect 7840 33920 7920 33934
rect 8000 33986 8080 34000
rect 8000 33934 8014 33986
rect 8066 33934 8080 33986
rect 8000 33920 8080 33934
rect 8160 33986 8240 34000
rect 8160 33934 8174 33986
rect 8226 33934 8240 33986
rect 8160 33920 8240 33934
rect 8320 33986 8400 34000
rect 8320 33934 8334 33986
rect 8386 33934 8400 33986
rect 8320 33920 8400 33934
rect 12480 33986 12560 34000
rect 12480 33934 12494 33986
rect 12546 33934 12560 33986
rect 12480 33920 12560 33934
rect 12640 33986 12720 34000
rect 12640 33934 12654 33986
rect 12706 33934 12720 33986
rect 12640 33920 12720 33934
rect 12800 33986 12880 34000
rect 12800 33934 12814 33986
rect 12866 33934 12880 33986
rect 12800 33920 12880 33934
rect 12960 33986 13040 34000
rect 12960 33934 12974 33986
rect 13026 33934 13040 33986
rect 12960 33920 13040 33934
rect 13120 33986 13200 34000
rect 13120 33934 13134 33986
rect 13186 33934 13200 33986
rect 13120 33920 13200 33934
rect 13280 33986 13360 34000
rect 13280 33934 13294 33986
rect 13346 33934 13360 33986
rect 13280 33920 13360 33934
rect 13440 33986 13520 34000
rect 13440 33934 13454 33986
rect 13506 33934 13520 33986
rect 13440 33920 13520 33934
rect 13600 33986 13680 34000
rect 13600 33934 13614 33986
rect 13666 33934 13680 33986
rect 13600 33920 13680 33934
rect 13760 33986 13840 34000
rect 13760 33934 13774 33986
rect 13826 33934 13840 33986
rect 13760 33920 13840 33934
rect 13920 33986 14000 34000
rect 13920 33934 13934 33986
rect 13986 33934 14000 33986
rect 13920 33920 14000 33934
rect 14080 33986 14160 34000
rect 14080 33934 14094 33986
rect 14146 33934 14160 33986
rect 14080 33920 14160 33934
rect 14240 33986 14320 34000
rect 14240 33934 14254 33986
rect 14306 33934 14320 33986
rect 14240 33920 14320 33934
rect 14400 33986 14480 34000
rect 14400 33934 14414 33986
rect 14466 33934 14480 33986
rect 14400 33920 14480 33934
rect 14560 33986 14640 34000
rect 14560 33934 14574 33986
rect 14626 33934 14640 33986
rect 14560 33920 14640 33934
rect 14720 33986 14800 34000
rect 14720 33934 14734 33986
rect 14786 33934 14800 33986
rect 14720 33920 14800 33934
rect 14880 33986 14960 34000
rect 14880 33934 14894 33986
rect 14946 33934 14960 33986
rect 14880 33920 14960 33934
rect 15040 33986 15120 34000
rect 15040 33934 15054 33986
rect 15106 33934 15120 33986
rect 15040 33920 15120 33934
rect 15200 33986 15280 34000
rect 15200 33934 15214 33986
rect 15266 33934 15280 33986
rect 15200 33920 15280 33934
rect 15360 33986 15440 34000
rect 15360 33934 15374 33986
rect 15426 33934 15440 33986
rect 15360 33920 15440 33934
rect 15520 33986 15600 34000
rect 15520 33934 15534 33986
rect 15586 33934 15600 33986
rect 15520 33920 15600 33934
rect 15680 33986 15760 34000
rect 15680 33934 15694 33986
rect 15746 33934 15760 33986
rect 15680 33920 15760 33934
rect 15840 33986 15920 34000
rect 15840 33934 15854 33986
rect 15906 33934 15920 33986
rect 15840 33920 15920 33934
rect 16000 33986 16080 34000
rect 16000 33934 16014 33986
rect 16066 33934 16080 33986
rect 16000 33920 16080 33934
rect 16160 33986 16240 34000
rect 16160 33934 16174 33986
rect 16226 33934 16240 33986
rect 16160 33920 16240 33934
rect 16320 33986 16400 34000
rect 16320 33934 16334 33986
rect 16386 33934 16400 33986
rect 16320 33920 16400 33934
rect 16480 33986 16560 34000
rect 16480 33934 16494 33986
rect 16546 33934 16560 33986
rect 16480 33920 16560 33934
rect 16640 33986 16720 34000
rect 16640 33934 16654 33986
rect 16706 33934 16720 33986
rect 16640 33920 16720 33934
rect 16800 33986 16880 34000
rect 16800 33934 16814 33986
rect 16866 33934 16880 33986
rect 16800 33920 16880 33934
rect 16960 33986 17040 34000
rect 16960 33934 16974 33986
rect 17026 33934 17040 33986
rect 16960 33920 17040 33934
rect 17120 33986 17200 34000
rect 17120 33934 17134 33986
rect 17186 33934 17200 33986
rect 17120 33920 17200 33934
rect 17280 33986 17360 34000
rect 17280 33934 17294 33986
rect 17346 33934 17360 33986
rect 17280 33920 17360 33934
rect 17440 33986 17520 34000
rect 17440 33934 17454 33986
rect 17506 33934 17520 33986
rect 17440 33920 17520 33934
rect 17600 33986 17680 34000
rect 17600 33934 17614 33986
rect 17666 33934 17680 33986
rect 17600 33920 17680 33934
rect 17760 33986 17840 34000
rect 17760 33934 17774 33986
rect 17826 33934 17840 33986
rect 17760 33920 17840 33934
rect 17920 33986 18000 34000
rect 17920 33934 17934 33986
rect 17986 33934 18000 33986
rect 17920 33920 18000 33934
rect 18080 33986 18160 34000
rect 18080 33934 18094 33986
rect 18146 33934 18160 33986
rect 18080 33920 18160 33934
rect 18240 33986 18320 34000
rect 18240 33934 18254 33986
rect 18306 33934 18320 33986
rect 18240 33920 18320 33934
rect 18400 33986 18480 34000
rect 18400 33934 18414 33986
rect 18466 33934 18480 33986
rect 18400 33920 18480 33934
rect 18560 33986 18640 34000
rect 18560 33934 18574 33986
rect 18626 33934 18640 33986
rect 18560 33920 18640 33934
rect 18720 33986 18800 34000
rect 18720 33934 18734 33986
rect 18786 33934 18800 33986
rect 18720 33920 18800 33934
rect 18880 33986 18960 34000
rect 18880 33934 18894 33986
rect 18946 33934 18960 33986
rect 18880 33920 18960 33934
rect 23120 33986 23200 34000
rect 23120 33934 23134 33986
rect 23186 33934 23200 33986
rect 23120 33920 23200 33934
rect 23280 33986 23360 34000
rect 23280 33934 23294 33986
rect 23346 33934 23360 33986
rect 23280 33920 23360 33934
rect 23440 33986 23520 34000
rect 23440 33934 23454 33986
rect 23506 33934 23520 33986
rect 23440 33920 23520 33934
rect 23600 33986 23680 34000
rect 23600 33934 23614 33986
rect 23666 33934 23680 33986
rect 23600 33920 23680 33934
rect 23760 33986 23840 34000
rect 23760 33934 23774 33986
rect 23826 33934 23840 33986
rect 23760 33920 23840 33934
rect 23920 33986 24000 34000
rect 23920 33934 23934 33986
rect 23986 33934 24000 33986
rect 23920 33920 24000 33934
rect 24080 33986 24160 34000
rect 24080 33934 24094 33986
rect 24146 33934 24160 33986
rect 24080 33920 24160 33934
rect 24240 33986 24320 34000
rect 24240 33934 24254 33986
rect 24306 33934 24320 33986
rect 24240 33920 24320 33934
rect 24400 33986 24480 34000
rect 24400 33934 24414 33986
rect 24466 33934 24480 33986
rect 24400 33920 24480 33934
rect 24560 33986 24640 34000
rect 24560 33934 24574 33986
rect 24626 33934 24640 33986
rect 24560 33920 24640 33934
rect 24720 33986 24800 34000
rect 24720 33934 24734 33986
rect 24786 33934 24800 33986
rect 24720 33920 24800 33934
rect 24880 33986 24960 34000
rect 24880 33934 24894 33986
rect 24946 33934 24960 33986
rect 24880 33920 24960 33934
rect 25040 33986 25120 34000
rect 25040 33934 25054 33986
rect 25106 33934 25120 33986
rect 25040 33920 25120 33934
rect 25200 33986 25280 34000
rect 25200 33934 25214 33986
rect 25266 33934 25280 33986
rect 25200 33920 25280 33934
rect 25360 33986 25440 34000
rect 25360 33934 25374 33986
rect 25426 33934 25440 33986
rect 25360 33920 25440 33934
rect 25520 33986 25600 34000
rect 25520 33934 25534 33986
rect 25586 33934 25600 33986
rect 25520 33920 25600 33934
rect 25680 33986 25760 34000
rect 25680 33934 25694 33986
rect 25746 33934 25760 33986
rect 25680 33920 25760 33934
rect 25840 33986 25920 34000
rect 25840 33934 25854 33986
rect 25906 33934 25920 33986
rect 25840 33920 25920 33934
rect 26000 33986 26080 34000
rect 26000 33934 26014 33986
rect 26066 33934 26080 33986
rect 26000 33920 26080 33934
rect 26160 33986 26240 34000
rect 26160 33934 26174 33986
rect 26226 33934 26240 33986
rect 26160 33920 26240 33934
rect 26320 33986 26400 34000
rect 26320 33934 26334 33986
rect 26386 33934 26400 33986
rect 26320 33920 26400 33934
rect 26480 33986 26560 34000
rect 26480 33934 26494 33986
rect 26546 33934 26560 33986
rect 26480 33920 26560 33934
rect 26640 33986 26720 34000
rect 26640 33934 26654 33986
rect 26706 33934 26720 33986
rect 26640 33920 26720 33934
rect 26800 33986 26880 34000
rect 26800 33934 26814 33986
rect 26866 33934 26880 33986
rect 26800 33920 26880 33934
rect 26960 33986 27040 34000
rect 26960 33934 26974 33986
rect 27026 33934 27040 33986
rect 26960 33920 27040 33934
rect 27120 33986 27200 34000
rect 27120 33934 27134 33986
rect 27186 33934 27200 33986
rect 27120 33920 27200 33934
rect 27280 33986 27360 34000
rect 27280 33934 27294 33986
rect 27346 33934 27360 33986
rect 27280 33920 27360 33934
rect 27440 33986 27520 34000
rect 27440 33934 27454 33986
rect 27506 33934 27520 33986
rect 27440 33920 27520 33934
rect 27600 33986 27680 34000
rect 27600 33934 27614 33986
rect 27666 33934 27680 33986
rect 27600 33920 27680 33934
rect 27760 33986 27840 34000
rect 27760 33934 27774 33986
rect 27826 33934 27840 33986
rect 27760 33920 27840 33934
rect 27920 33986 28000 34000
rect 27920 33934 27934 33986
rect 27986 33934 28000 33986
rect 27920 33920 28000 33934
rect 28080 33986 28160 34000
rect 28080 33934 28094 33986
rect 28146 33934 28160 33986
rect 28080 33920 28160 33934
rect 28240 33986 28320 34000
rect 28240 33934 28254 33986
rect 28306 33934 28320 33986
rect 28240 33920 28320 33934
rect 28400 33986 28480 34000
rect 28400 33934 28414 33986
rect 28466 33934 28480 33986
rect 28400 33920 28480 33934
rect 28560 33986 28640 34000
rect 28560 33934 28574 33986
rect 28626 33934 28640 33986
rect 28560 33920 28640 33934
rect 28720 33986 28800 34000
rect 28720 33934 28734 33986
rect 28786 33934 28800 33986
rect 28720 33920 28800 33934
rect 28880 33986 28960 34000
rect 28880 33934 28894 33986
rect 28946 33934 28960 33986
rect 28880 33920 28960 33934
rect 29040 33986 29120 34000
rect 29040 33934 29054 33986
rect 29106 33934 29120 33986
rect 29040 33920 29120 33934
rect 29200 33986 29280 34000
rect 29200 33934 29214 33986
rect 29266 33934 29280 33986
rect 29200 33920 29280 33934
rect 29360 33986 29440 34000
rect 29360 33934 29374 33986
rect 29426 33934 29440 33986
rect 29360 33920 29440 33934
rect 33520 33986 33600 34000
rect 33520 33934 33534 33986
rect 33586 33934 33600 33986
rect 33520 33920 33600 33934
rect 33680 33986 33760 34000
rect 33680 33934 33694 33986
rect 33746 33934 33760 33986
rect 33680 33920 33760 33934
rect 33840 33986 33920 34000
rect 33840 33934 33854 33986
rect 33906 33934 33920 33986
rect 33840 33920 33920 33934
rect 34000 33986 34080 34000
rect 34000 33934 34014 33986
rect 34066 33934 34080 33986
rect 34000 33920 34080 33934
rect 34160 33986 34240 34000
rect 34160 33934 34174 33986
rect 34226 33934 34240 33986
rect 34160 33920 34240 33934
rect 34320 33986 34400 34000
rect 34320 33934 34334 33986
rect 34386 33934 34400 33986
rect 34320 33920 34400 33934
rect 34480 33986 34560 34000
rect 34480 33934 34494 33986
rect 34546 33934 34560 33986
rect 34480 33920 34560 33934
rect 34640 33986 34720 34000
rect 34640 33934 34654 33986
rect 34706 33934 34720 33986
rect 34640 33920 34720 33934
rect 34800 33986 34880 34000
rect 34800 33934 34814 33986
rect 34866 33934 34880 33986
rect 34800 33920 34880 33934
rect 34960 33986 35040 34000
rect 34960 33934 34974 33986
rect 35026 33934 35040 33986
rect 34960 33920 35040 33934
rect 35120 33986 35200 34000
rect 35120 33934 35134 33986
rect 35186 33934 35200 33986
rect 35120 33920 35200 33934
rect 35280 33986 35360 34000
rect 35280 33934 35294 33986
rect 35346 33934 35360 33986
rect 35280 33920 35360 33934
rect 35440 33986 35520 34000
rect 35440 33934 35454 33986
rect 35506 33934 35520 33986
rect 35440 33920 35520 33934
rect 35600 33986 35680 34000
rect 35600 33934 35614 33986
rect 35666 33934 35680 33986
rect 35600 33920 35680 33934
rect 35760 33986 35840 34000
rect 35760 33934 35774 33986
rect 35826 33934 35840 33986
rect 35760 33920 35840 33934
rect 35920 33986 36000 34000
rect 35920 33934 35934 33986
rect 35986 33934 36000 33986
rect 35920 33920 36000 33934
rect 36080 33986 36160 34000
rect 36080 33934 36094 33986
rect 36146 33934 36160 33986
rect 36080 33920 36160 33934
rect 36240 33986 36320 34000
rect 36240 33934 36254 33986
rect 36306 33934 36320 33986
rect 36240 33920 36320 33934
rect 36400 33986 36480 34000
rect 36400 33934 36414 33986
rect 36466 33934 36480 33986
rect 36400 33920 36480 33934
rect 36560 33986 36640 34000
rect 36560 33934 36574 33986
rect 36626 33934 36640 33986
rect 36560 33920 36640 33934
rect 36720 33986 36800 34000
rect 36720 33934 36734 33986
rect 36786 33934 36800 33986
rect 36720 33920 36800 33934
rect 36880 33986 36960 34000
rect 36880 33934 36894 33986
rect 36946 33934 36960 33986
rect 36880 33920 36960 33934
rect 37040 33986 37120 34000
rect 37040 33934 37054 33986
rect 37106 33934 37120 33986
rect 37040 33920 37120 33934
rect 37200 33986 37280 34000
rect 37200 33934 37214 33986
rect 37266 33934 37280 33986
rect 37200 33920 37280 33934
rect 37360 33986 37440 34000
rect 37360 33934 37374 33986
rect 37426 33934 37440 33986
rect 37360 33920 37440 33934
rect 37520 33986 37600 34000
rect 37520 33934 37534 33986
rect 37586 33934 37600 33986
rect 37520 33920 37600 33934
rect 37680 33986 37760 34000
rect 37680 33934 37694 33986
rect 37746 33934 37760 33986
rect 37680 33920 37760 33934
rect 37840 33986 37920 34000
rect 37840 33934 37854 33986
rect 37906 33934 37920 33986
rect 37840 33920 37920 33934
rect 38000 33986 38080 34000
rect 38000 33934 38014 33986
rect 38066 33934 38080 33986
rect 38000 33920 38080 33934
rect 38160 33986 38240 34000
rect 38160 33934 38174 33986
rect 38226 33934 38240 33986
rect 38160 33920 38240 33934
rect 38320 33986 38400 34000
rect 38320 33934 38334 33986
rect 38386 33934 38400 33986
rect 38320 33920 38400 33934
rect 38480 33986 38560 34000
rect 38480 33934 38494 33986
rect 38546 33934 38560 33986
rect 38480 33920 38560 33934
rect 38640 33986 38720 34000
rect 38640 33934 38654 33986
rect 38706 33934 38720 33986
rect 38640 33920 38720 33934
rect 38800 33986 38880 34000
rect 38800 33934 38814 33986
rect 38866 33934 38880 33986
rect 38800 33920 38880 33934
rect 38960 33986 39040 34000
rect 38960 33934 38974 33986
rect 39026 33934 39040 33986
rect 38960 33920 39040 33934
rect 39120 33986 39200 34000
rect 39120 33934 39134 33986
rect 39186 33934 39200 33986
rect 39120 33920 39200 33934
rect 39280 33986 39360 34000
rect 39280 33934 39294 33986
rect 39346 33934 39360 33986
rect 39280 33920 39360 33934
rect 39440 33986 39520 34000
rect 39440 33934 39454 33986
rect 39506 33934 39520 33986
rect 39440 33920 39520 33934
rect 39600 33986 39680 34000
rect 39600 33934 39614 33986
rect 39666 33934 39680 33986
rect 39600 33920 39680 33934
rect 39760 33986 39840 34000
rect 39760 33934 39774 33986
rect 39826 33934 39840 33986
rect 39760 33920 39840 33934
rect 39920 33986 40000 34000
rect 39920 33934 39934 33986
rect 39986 33934 40000 33986
rect 39920 33920 40000 33934
rect 40080 33986 40160 34000
rect 40080 33934 40094 33986
rect 40146 33934 40160 33986
rect 40080 33920 40160 33934
rect 40240 33986 40320 34000
rect 40240 33934 40254 33986
rect 40306 33934 40320 33986
rect 40240 33920 40320 33934
rect 40400 33986 40480 34000
rect 40400 33934 40414 33986
rect 40466 33934 40480 33986
rect 40400 33920 40480 33934
rect 40560 33986 40640 34000
rect 40560 33934 40574 33986
rect 40626 33934 40640 33986
rect 40560 33920 40640 33934
rect 40720 33986 40800 34000
rect 40720 33934 40734 33986
rect 40786 33934 40800 33986
rect 40720 33920 40800 33934
rect 40880 33986 40960 34000
rect 40880 33934 40894 33986
rect 40946 33934 40960 33986
rect 40880 33920 40960 33934
rect 41040 33986 41120 34000
rect 41040 33934 41054 33986
rect 41106 33934 41120 33986
rect 41040 33920 41120 33934
rect 41200 33986 41280 34000
rect 41200 33934 41214 33986
rect 41266 33934 41280 33986
rect 41200 33920 41280 33934
rect 41360 33986 41440 34000
rect 41360 33934 41374 33986
rect 41426 33934 41440 33986
rect 41360 33920 41440 33934
rect 41520 33986 41600 34000
rect 41520 33934 41534 33986
rect 41586 33934 41600 33986
rect 41520 33920 41600 33934
rect 41680 33986 41760 34000
rect 41680 33934 41694 33986
rect 41746 33934 41760 33986
rect 41680 33920 41760 33934
rect 41840 33986 41920 34000
rect 41840 33934 41854 33986
rect 41906 33934 41920 33986
rect 41840 33920 41920 33934
rect 0 33826 80 33840
rect 0 33774 14 33826
rect 66 33774 80 33826
rect 0 33760 80 33774
rect 160 33826 240 33840
rect 160 33774 174 33826
rect 226 33774 240 33826
rect 160 33760 240 33774
rect 320 33826 400 33840
rect 320 33774 334 33826
rect 386 33774 400 33826
rect 320 33760 400 33774
rect 480 33826 560 33840
rect 480 33774 494 33826
rect 546 33774 560 33826
rect 480 33760 560 33774
rect 640 33826 720 33840
rect 640 33774 654 33826
rect 706 33774 720 33826
rect 640 33760 720 33774
rect 800 33826 880 33840
rect 800 33774 814 33826
rect 866 33774 880 33826
rect 800 33760 880 33774
rect 960 33826 1040 33840
rect 960 33774 974 33826
rect 1026 33774 1040 33826
rect 960 33760 1040 33774
rect 1120 33826 1200 33840
rect 1120 33774 1134 33826
rect 1186 33774 1200 33826
rect 1120 33760 1200 33774
rect 1280 33826 1360 33840
rect 1280 33774 1294 33826
rect 1346 33774 1360 33826
rect 1280 33760 1360 33774
rect 1440 33826 1520 33840
rect 1440 33774 1454 33826
rect 1506 33774 1520 33826
rect 1440 33760 1520 33774
rect 1600 33826 1680 33840
rect 1600 33774 1614 33826
rect 1666 33774 1680 33826
rect 1600 33760 1680 33774
rect 1760 33826 1840 33840
rect 1760 33774 1774 33826
rect 1826 33774 1840 33826
rect 1760 33760 1840 33774
rect 1920 33826 2000 33840
rect 1920 33774 1934 33826
rect 1986 33774 2000 33826
rect 1920 33760 2000 33774
rect 2080 33826 2160 33840
rect 2080 33774 2094 33826
rect 2146 33774 2160 33826
rect 2080 33760 2160 33774
rect 2240 33826 2320 33840
rect 2240 33774 2254 33826
rect 2306 33774 2320 33826
rect 2240 33760 2320 33774
rect 2400 33826 2480 33840
rect 2400 33774 2414 33826
rect 2466 33774 2480 33826
rect 2400 33760 2480 33774
rect 2560 33826 2640 33840
rect 2560 33774 2574 33826
rect 2626 33774 2640 33826
rect 2560 33760 2640 33774
rect 2720 33826 2800 33840
rect 2720 33774 2734 33826
rect 2786 33774 2800 33826
rect 2720 33760 2800 33774
rect 2880 33826 2960 33840
rect 2880 33774 2894 33826
rect 2946 33774 2960 33826
rect 2880 33760 2960 33774
rect 3040 33826 3120 33840
rect 3040 33774 3054 33826
rect 3106 33774 3120 33826
rect 3040 33760 3120 33774
rect 3200 33826 3280 33840
rect 3200 33774 3214 33826
rect 3266 33774 3280 33826
rect 3200 33760 3280 33774
rect 3360 33826 3440 33840
rect 3360 33774 3374 33826
rect 3426 33774 3440 33826
rect 3360 33760 3440 33774
rect 3520 33826 3600 33840
rect 3520 33774 3534 33826
rect 3586 33774 3600 33826
rect 3520 33760 3600 33774
rect 3680 33826 3760 33840
rect 3680 33774 3694 33826
rect 3746 33774 3760 33826
rect 3680 33760 3760 33774
rect 3840 33826 3920 33840
rect 3840 33774 3854 33826
rect 3906 33774 3920 33826
rect 3840 33760 3920 33774
rect 4000 33826 4080 33840
rect 4000 33774 4014 33826
rect 4066 33774 4080 33826
rect 4000 33760 4080 33774
rect 4160 33826 4240 33840
rect 4160 33774 4174 33826
rect 4226 33774 4240 33826
rect 4160 33760 4240 33774
rect 4320 33826 4400 33840
rect 4320 33774 4334 33826
rect 4386 33774 4400 33826
rect 4320 33760 4400 33774
rect 4480 33826 4560 33840
rect 4480 33774 4494 33826
rect 4546 33774 4560 33826
rect 4480 33760 4560 33774
rect 4640 33826 4720 33840
rect 4640 33774 4654 33826
rect 4706 33774 4720 33826
rect 4640 33760 4720 33774
rect 4800 33826 4880 33840
rect 4800 33774 4814 33826
rect 4866 33774 4880 33826
rect 4800 33760 4880 33774
rect 4960 33826 5040 33840
rect 4960 33774 4974 33826
rect 5026 33774 5040 33826
rect 4960 33760 5040 33774
rect 5120 33826 5200 33840
rect 5120 33774 5134 33826
rect 5186 33774 5200 33826
rect 5120 33760 5200 33774
rect 5280 33826 5360 33840
rect 5280 33774 5294 33826
rect 5346 33774 5360 33826
rect 5280 33760 5360 33774
rect 5440 33826 5520 33840
rect 5440 33774 5454 33826
rect 5506 33774 5520 33826
rect 5440 33760 5520 33774
rect 5600 33826 5680 33840
rect 5600 33774 5614 33826
rect 5666 33774 5680 33826
rect 5600 33760 5680 33774
rect 5760 33826 5840 33840
rect 5760 33774 5774 33826
rect 5826 33774 5840 33826
rect 5760 33760 5840 33774
rect 5920 33826 6000 33840
rect 5920 33774 5934 33826
rect 5986 33774 6000 33826
rect 5920 33760 6000 33774
rect 6080 33826 6160 33840
rect 6080 33774 6094 33826
rect 6146 33774 6160 33826
rect 6080 33760 6160 33774
rect 6240 33826 6320 33840
rect 6240 33774 6254 33826
rect 6306 33774 6320 33826
rect 6240 33760 6320 33774
rect 6400 33826 6480 33840
rect 6400 33774 6414 33826
rect 6466 33774 6480 33826
rect 6400 33760 6480 33774
rect 6560 33826 6640 33840
rect 6560 33774 6574 33826
rect 6626 33774 6640 33826
rect 6560 33760 6640 33774
rect 6720 33826 6800 33840
rect 6720 33774 6734 33826
rect 6786 33774 6800 33826
rect 6720 33760 6800 33774
rect 6880 33826 6960 33840
rect 6880 33774 6894 33826
rect 6946 33774 6960 33826
rect 6880 33760 6960 33774
rect 7040 33826 7120 33840
rect 7040 33774 7054 33826
rect 7106 33774 7120 33826
rect 7040 33760 7120 33774
rect 7200 33826 7280 33840
rect 7200 33774 7214 33826
rect 7266 33774 7280 33826
rect 7200 33760 7280 33774
rect 7360 33826 7440 33840
rect 7360 33774 7374 33826
rect 7426 33774 7440 33826
rect 7360 33760 7440 33774
rect 7520 33826 7600 33840
rect 7520 33774 7534 33826
rect 7586 33774 7600 33826
rect 7520 33760 7600 33774
rect 7680 33826 7760 33840
rect 7680 33774 7694 33826
rect 7746 33774 7760 33826
rect 7680 33760 7760 33774
rect 7840 33826 7920 33840
rect 7840 33774 7854 33826
rect 7906 33774 7920 33826
rect 7840 33760 7920 33774
rect 8000 33826 8080 33840
rect 8000 33774 8014 33826
rect 8066 33774 8080 33826
rect 8000 33760 8080 33774
rect 8160 33826 8240 33840
rect 8160 33774 8174 33826
rect 8226 33774 8240 33826
rect 8160 33760 8240 33774
rect 8320 33826 8400 33840
rect 8320 33774 8334 33826
rect 8386 33774 8400 33826
rect 8320 33760 8400 33774
rect 12480 33826 12560 33840
rect 12480 33774 12494 33826
rect 12546 33774 12560 33826
rect 12480 33760 12560 33774
rect 12640 33826 12720 33840
rect 12640 33774 12654 33826
rect 12706 33774 12720 33826
rect 12640 33760 12720 33774
rect 12800 33826 12880 33840
rect 12800 33774 12814 33826
rect 12866 33774 12880 33826
rect 12800 33760 12880 33774
rect 12960 33826 13040 33840
rect 12960 33774 12974 33826
rect 13026 33774 13040 33826
rect 12960 33760 13040 33774
rect 13120 33826 13200 33840
rect 13120 33774 13134 33826
rect 13186 33774 13200 33826
rect 13120 33760 13200 33774
rect 13280 33826 13360 33840
rect 13280 33774 13294 33826
rect 13346 33774 13360 33826
rect 13280 33760 13360 33774
rect 13440 33826 13520 33840
rect 13440 33774 13454 33826
rect 13506 33774 13520 33826
rect 13440 33760 13520 33774
rect 13600 33826 13680 33840
rect 13600 33774 13614 33826
rect 13666 33774 13680 33826
rect 13600 33760 13680 33774
rect 13760 33826 13840 33840
rect 13760 33774 13774 33826
rect 13826 33774 13840 33826
rect 13760 33760 13840 33774
rect 13920 33826 14000 33840
rect 13920 33774 13934 33826
rect 13986 33774 14000 33826
rect 13920 33760 14000 33774
rect 14080 33826 14160 33840
rect 14080 33774 14094 33826
rect 14146 33774 14160 33826
rect 14080 33760 14160 33774
rect 14240 33826 14320 33840
rect 14240 33774 14254 33826
rect 14306 33774 14320 33826
rect 14240 33760 14320 33774
rect 14400 33826 14480 33840
rect 14400 33774 14414 33826
rect 14466 33774 14480 33826
rect 14400 33760 14480 33774
rect 14560 33826 14640 33840
rect 14560 33774 14574 33826
rect 14626 33774 14640 33826
rect 14560 33760 14640 33774
rect 14720 33826 14800 33840
rect 14720 33774 14734 33826
rect 14786 33774 14800 33826
rect 14720 33760 14800 33774
rect 14880 33826 14960 33840
rect 14880 33774 14894 33826
rect 14946 33774 14960 33826
rect 14880 33760 14960 33774
rect 15040 33826 15120 33840
rect 15040 33774 15054 33826
rect 15106 33774 15120 33826
rect 15040 33760 15120 33774
rect 15200 33826 15280 33840
rect 15200 33774 15214 33826
rect 15266 33774 15280 33826
rect 15200 33760 15280 33774
rect 15360 33826 15440 33840
rect 15360 33774 15374 33826
rect 15426 33774 15440 33826
rect 15360 33760 15440 33774
rect 15520 33826 15600 33840
rect 15520 33774 15534 33826
rect 15586 33774 15600 33826
rect 15520 33760 15600 33774
rect 15680 33826 15760 33840
rect 15680 33774 15694 33826
rect 15746 33774 15760 33826
rect 15680 33760 15760 33774
rect 15840 33826 15920 33840
rect 15840 33774 15854 33826
rect 15906 33774 15920 33826
rect 15840 33760 15920 33774
rect 16000 33826 16080 33840
rect 16000 33774 16014 33826
rect 16066 33774 16080 33826
rect 16000 33760 16080 33774
rect 16160 33826 16240 33840
rect 16160 33774 16174 33826
rect 16226 33774 16240 33826
rect 16160 33760 16240 33774
rect 16320 33826 16400 33840
rect 16320 33774 16334 33826
rect 16386 33774 16400 33826
rect 16320 33760 16400 33774
rect 16480 33826 16560 33840
rect 16480 33774 16494 33826
rect 16546 33774 16560 33826
rect 16480 33760 16560 33774
rect 16640 33826 16720 33840
rect 16640 33774 16654 33826
rect 16706 33774 16720 33826
rect 16640 33760 16720 33774
rect 16800 33826 16880 33840
rect 16800 33774 16814 33826
rect 16866 33774 16880 33826
rect 16800 33760 16880 33774
rect 16960 33826 17040 33840
rect 16960 33774 16974 33826
rect 17026 33774 17040 33826
rect 16960 33760 17040 33774
rect 17120 33826 17200 33840
rect 17120 33774 17134 33826
rect 17186 33774 17200 33826
rect 17120 33760 17200 33774
rect 17280 33826 17360 33840
rect 17280 33774 17294 33826
rect 17346 33774 17360 33826
rect 17280 33760 17360 33774
rect 17440 33826 17520 33840
rect 17440 33774 17454 33826
rect 17506 33774 17520 33826
rect 17440 33760 17520 33774
rect 17600 33826 17680 33840
rect 17600 33774 17614 33826
rect 17666 33774 17680 33826
rect 17600 33760 17680 33774
rect 17760 33826 17840 33840
rect 17760 33774 17774 33826
rect 17826 33774 17840 33826
rect 17760 33760 17840 33774
rect 17920 33826 18000 33840
rect 17920 33774 17934 33826
rect 17986 33774 18000 33826
rect 17920 33760 18000 33774
rect 18080 33826 18160 33840
rect 18080 33774 18094 33826
rect 18146 33774 18160 33826
rect 18080 33760 18160 33774
rect 18240 33826 18320 33840
rect 18240 33774 18254 33826
rect 18306 33774 18320 33826
rect 18240 33760 18320 33774
rect 18400 33826 18480 33840
rect 18400 33774 18414 33826
rect 18466 33774 18480 33826
rect 18400 33760 18480 33774
rect 18560 33826 18640 33840
rect 18560 33774 18574 33826
rect 18626 33774 18640 33826
rect 18560 33760 18640 33774
rect 18720 33826 18800 33840
rect 18720 33774 18734 33826
rect 18786 33774 18800 33826
rect 18720 33760 18800 33774
rect 18880 33826 18960 33840
rect 18880 33774 18894 33826
rect 18946 33774 18960 33826
rect 18880 33760 18960 33774
rect 23120 33826 23200 33840
rect 23120 33774 23134 33826
rect 23186 33774 23200 33826
rect 23120 33760 23200 33774
rect 23280 33826 23360 33840
rect 23280 33774 23294 33826
rect 23346 33774 23360 33826
rect 23280 33760 23360 33774
rect 23440 33826 23520 33840
rect 23440 33774 23454 33826
rect 23506 33774 23520 33826
rect 23440 33760 23520 33774
rect 23600 33826 23680 33840
rect 23600 33774 23614 33826
rect 23666 33774 23680 33826
rect 23600 33760 23680 33774
rect 23760 33826 23840 33840
rect 23760 33774 23774 33826
rect 23826 33774 23840 33826
rect 23760 33760 23840 33774
rect 23920 33826 24000 33840
rect 23920 33774 23934 33826
rect 23986 33774 24000 33826
rect 23920 33760 24000 33774
rect 24080 33826 24160 33840
rect 24080 33774 24094 33826
rect 24146 33774 24160 33826
rect 24080 33760 24160 33774
rect 24240 33826 24320 33840
rect 24240 33774 24254 33826
rect 24306 33774 24320 33826
rect 24240 33760 24320 33774
rect 24400 33826 24480 33840
rect 24400 33774 24414 33826
rect 24466 33774 24480 33826
rect 24400 33760 24480 33774
rect 24560 33826 24640 33840
rect 24560 33774 24574 33826
rect 24626 33774 24640 33826
rect 24560 33760 24640 33774
rect 24720 33826 24800 33840
rect 24720 33774 24734 33826
rect 24786 33774 24800 33826
rect 24720 33760 24800 33774
rect 24880 33826 24960 33840
rect 24880 33774 24894 33826
rect 24946 33774 24960 33826
rect 24880 33760 24960 33774
rect 25040 33826 25120 33840
rect 25040 33774 25054 33826
rect 25106 33774 25120 33826
rect 25040 33760 25120 33774
rect 25200 33826 25280 33840
rect 25200 33774 25214 33826
rect 25266 33774 25280 33826
rect 25200 33760 25280 33774
rect 25360 33826 25440 33840
rect 25360 33774 25374 33826
rect 25426 33774 25440 33826
rect 25360 33760 25440 33774
rect 25520 33826 25600 33840
rect 25520 33774 25534 33826
rect 25586 33774 25600 33826
rect 25520 33760 25600 33774
rect 25680 33826 25760 33840
rect 25680 33774 25694 33826
rect 25746 33774 25760 33826
rect 25680 33760 25760 33774
rect 25840 33826 25920 33840
rect 25840 33774 25854 33826
rect 25906 33774 25920 33826
rect 25840 33760 25920 33774
rect 26000 33826 26080 33840
rect 26000 33774 26014 33826
rect 26066 33774 26080 33826
rect 26000 33760 26080 33774
rect 26160 33826 26240 33840
rect 26160 33774 26174 33826
rect 26226 33774 26240 33826
rect 26160 33760 26240 33774
rect 26320 33826 26400 33840
rect 26320 33774 26334 33826
rect 26386 33774 26400 33826
rect 26320 33760 26400 33774
rect 26480 33826 26560 33840
rect 26480 33774 26494 33826
rect 26546 33774 26560 33826
rect 26480 33760 26560 33774
rect 26640 33826 26720 33840
rect 26640 33774 26654 33826
rect 26706 33774 26720 33826
rect 26640 33760 26720 33774
rect 26800 33826 26880 33840
rect 26800 33774 26814 33826
rect 26866 33774 26880 33826
rect 26800 33760 26880 33774
rect 26960 33826 27040 33840
rect 26960 33774 26974 33826
rect 27026 33774 27040 33826
rect 26960 33760 27040 33774
rect 27120 33826 27200 33840
rect 27120 33774 27134 33826
rect 27186 33774 27200 33826
rect 27120 33760 27200 33774
rect 27280 33826 27360 33840
rect 27280 33774 27294 33826
rect 27346 33774 27360 33826
rect 27280 33760 27360 33774
rect 27440 33826 27520 33840
rect 27440 33774 27454 33826
rect 27506 33774 27520 33826
rect 27440 33760 27520 33774
rect 27600 33826 27680 33840
rect 27600 33774 27614 33826
rect 27666 33774 27680 33826
rect 27600 33760 27680 33774
rect 27760 33826 27840 33840
rect 27760 33774 27774 33826
rect 27826 33774 27840 33826
rect 27760 33760 27840 33774
rect 27920 33826 28000 33840
rect 27920 33774 27934 33826
rect 27986 33774 28000 33826
rect 27920 33760 28000 33774
rect 28080 33826 28160 33840
rect 28080 33774 28094 33826
rect 28146 33774 28160 33826
rect 28080 33760 28160 33774
rect 28240 33826 28320 33840
rect 28240 33774 28254 33826
rect 28306 33774 28320 33826
rect 28240 33760 28320 33774
rect 28400 33826 28480 33840
rect 28400 33774 28414 33826
rect 28466 33774 28480 33826
rect 28400 33760 28480 33774
rect 28560 33826 28640 33840
rect 28560 33774 28574 33826
rect 28626 33774 28640 33826
rect 28560 33760 28640 33774
rect 28720 33826 28800 33840
rect 28720 33774 28734 33826
rect 28786 33774 28800 33826
rect 28720 33760 28800 33774
rect 28880 33826 28960 33840
rect 28880 33774 28894 33826
rect 28946 33774 28960 33826
rect 28880 33760 28960 33774
rect 29040 33826 29120 33840
rect 29040 33774 29054 33826
rect 29106 33774 29120 33826
rect 29040 33760 29120 33774
rect 29200 33826 29280 33840
rect 29200 33774 29214 33826
rect 29266 33774 29280 33826
rect 29200 33760 29280 33774
rect 29360 33826 29440 33840
rect 29360 33774 29374 33826
rect 29426 33774 29440 33826
rect 29360 33760 29440 33774
rect 33520 33826 33600 33840
rect 33520 33774 33534 33826
rect 33586 33774 33600 33826
rect 33520 33760 33600 33774
rect 33680 33826 33760 33840
rect 33680 33774 33694 33826
rect 33746 33774 33760 33826
rect 33680 33760 33760 33774
rect 33840 33826 33920 33840
rect 33840 33774 33854 33826
rect 33906 33774 33920 33826
rect 33840 33760 33920 33774
rect 34000 33826 34080 33840
rect 34000 33774 34014 33826
rect 34066 33774 34080 33826
rect 34000 33760 34080 33774
rect 34160 33826 34240 33840
rect 34160 33774 34174 33826
rect 34226 33774 34240 33826
rect 34160 33760 34240 33774
rect 34320 33826 34400 33840
rect 34320 33774 34334 33826
rect 34386 33774 34400 33826
rect 34320 33760 34400 33774
rect 34480 33826 34560 33840
rect 34480 33774 34494 33826
rect 34546 33774 34560 33826
rect 34480 33760 34560 33774
rect 34640 33826 34720 33840
rect 34640 33774 34654 33826
rect 34706 33774 34720 33826
rect 34640 33760 34720 33774
rect 34800 33826 34880 33840
rect 34800 33774 34814 33826
rect 34866 33774 34880 33826
rect 34800 33760 34880 33774
rect 34960 33826 35040 33840
rect 34960 33774 34974 33826
rect 35026 33774 35040 33826
rect 34960 33760 35040 33774
rect 35120 33826 35200 33840
rect 35120 33774 35134 33826
rect 35186 33774 35200 33826
rect 35120 33760 35200 33774
rect 35280 33826 35360 33840
rect 35280 33774 35294 33826
rect 35346 33774 35360 33826
rect 35280 33760 35360 33774
rect 35440 33826 35520 33840
rect 35440 33774 35454 33826
rect 35506 33774 35520 33826
rect 35440 33760 35520 33774
rect 35600 33826 35680 33840
rect 35600 33774 35614 33826
rect 35666 33774 35680 33826
rect 35600 33760 35680 33774
rect 35760 33826 35840 33840
rect 35760 33774 35774 33826
rect 35826 33774 35840 33826
rect 35760 33760 35840 33774
rect 35920 33826 36000 33840
rect 35920 33774 35934 33826
rect 35986 33774 36000 33826
rect 35920 33760 36000 33774
rect 36080 33826 36160 33840
rect 36080 33774 36094 33826
rect 36146 33774 36160 33826
rect 36080 33760 36160 33774
rect 36240 33826 36320 33840
rect 36240 33774 36254 33826
rect 36306 33774 36320 33826
rect 36240 33760 36320 33774
rect 36400 33826 36480 33840
rect 36400 33774 36414 33826
rect 36466 33774 36480 33826
rect 36400 33760 36480 33774
rect 36560 33826 36640 33840
rect 36560 33774 36574 33826
rect 36626 33774 36640 33826
rect 36560 33760 36640 33774
rect 36720 33826 36800 33840
rect 36720 33774 36734 33826
rect 36786 33774 36800 33826
rect 36720 33760 36800 33774
rect 36880 33826 36960 33840
rect 36880 33774 36894 33826
rect 36946 33774 36960 33826
rect 36880 33760 36960 33774
rect 37040 33826 37120 33840
rect 37040 33774 37054 33826
rect 37106 33774 37120 33826
rect 37040 33760 37120 33774
rect 37200 33826 37280 33840
rect 37200 33774 37214 33826
rect 37266 33774 37280 33826
rect 37200 33760 37280 33774
rect 37360 33826 37440 33840
rect 37360 33774 37374 33826
rect 37426 33774 37440 33826
rect 37360 33760 37440 33774
rect 37520 33826 37600 33840
rect 37520 33774 37534 33826
rect 37586 33774 37600 33826
rect 37520 33760 37600 33774
rect 37680 33826 37760 33840
rect 37680 33774 37694 33826
rect 37746 33774 37760 33826
rect 37680 33760 37760 33774
rect 37840 33826 37920 33840
rect 37840 33774 37854 33826
rect 37906 33774 37920 33826
rect 37840 33760 37920 33774
rect 38000 33826 38080 33840
rect 38000 33774 38014 33826
rect 38066 33774 38080 33826
rect 38000 33760 38080 33774
rect 38160 33826 38240 33840
rect 38160 33774 38174 33826
rect 38226 33774 38240 33826
rect 38160 33760 38240 33774
rect 38320 33826 38400 33840
rect 38320 33774 38334 33826
rect 38386 33774 38400 33826
rect 38320 33760 38400 33774
rect 38480 33826 38560 33840
rect 38480 33774 38494 33826
rect 38546 33774 38560 33826
rect 38480 33760 38560 33774
rect 38640 33826 38720 33840
rect 38640 33774 38654 33826
rect 38706 33774 38720 33826
rect 38640 33760 38720 33774
rect 38800 33826 38880 33840
rect 38800 33774 38814 33826
rect 38866 33774 38880 33826
rect 38800 33760 38880 33774
rect 38960 33826 39040 33840
rect 38960 33774 38974 33826
rect 39026 33774 39040 33826
rect 38960 33760 39040 33774
rect 39120 33826 39200 33840
rect 39120 33774 39134 33826
rect 39186 33774 39200 33826
rect 39120 33760 39200 33774
rect 39280 33826 39360 33840
rect 39280 33774 39294 33826
rect 39346 33774 39360 33826
rect 39280 33760 39360 33774
rect 39440 33826 39520 33840
rect 39440 33774 39454 33826
rect 39506 33774 39520 33826
rect 39440 33760 39520 33774
rect 39600 33826 39680 33840
rect 39600 33774 39614 33826
rect 39666 33774 39680 33826
rect 39600 33760 39680 33774
rect 39760 33826 39840 33840
rect 39760 33774 39774 33826
rect 39826 33774 39840 33826
rect 39760 33760 39840 33774
rect 39920 33826 40000 33840
rect 39920 33774 39934 33826
rect 39986 33774 40000 33826
rect 39920 33760 40000 33774
rect 40080 33826 40160 33840
rect 40080 33774 40094 33826
rect 40146 33774 40160 33826
rect 40080 33760 40160 33774
rect 40240 33826 40320 33840
rect 40240 33774 40254 33826
rect 40306 33774 40320 33826
rect 40240 33760 40320 33774
rect 40400 33826 40480 33840
rect 40400 33774 40414 33826
rect 40466 33774 40480 33826
rect 40400 33760 40480 33774
rect 40560 33826 40640 33840
rect 40560 33774 40574 33826
rect 40626 33774 40640 33826
rect 40560 33760 40640 33774
rect 40720 33826 40800 33840
rect 40720 33774 40734 33826
rect 40786 33774 40800 33826
rect 40720 33760 40800 33774
rect 40880 33826 40960 33840
rect 40880 33774 40894 33826
rect 40946 33774 40960 33826
rect 40880 33760 40960 33774
rect 41040 33826 41120 33840
rect 41040 33774 41054 33826
rect 41106 33774 41120 33826
rect 41040 33760 41120 33774
rect 41200 33826 41280 33840
rect 41200 33774 41214 33826
rect 41266 33774 41280 33826
rect 41200 33760 41280 33774
rect 41360 33826 41440 33840
rect 41360 33774 41374 33826
rect 41426 33774 41440 33826
rect 41360 33760 41440 33774
rect 41520 33826 41600 33840
rect 41520 33774 41534 33826
rect 41586 33774 41600 33826
rect 41520 33760 41600 33774
rect 41680 33826 41760 33840
rect 41680 33774 41694 33826
rect 41746 33774 41760 33826
rect 41680 33760 41760 33774
rect 41840 33826 41920 33840
rect 41840 33774 41854 33826
rect 41906 33774 41920 33826
rect 41840 33760 41920 33774
rect 0 33506 80 33520
rect 0 33454 14 33506
rect 66 33454 80 33506
rect 0 33440 80 33454
rect 160 33506 240 33520
rect 160 33454 174 33506
rect 226 33454 240 33506
rect 160 33440 240 33454
rect 320 33506 400 33520
rect 320 33454 334 33506
rect 386 33454 400 33506
rect 320 33440 400 33454
rect 480 33506 560 33520
rect 480 33454 494 33506
rect 546 33454 560 33506
rect 480 33440 560 33454
rect 640 33506 720 33520
rect 640 33454 654 33506
rect 706 33454 720 33506
rect 640 33440 720 33454
rect 800 33506 880 33520
rect 800 33454 814 33506
rect 866 33454 880 33506
rect 800 33440 880 33454
rect 960 33506 1040 33520
rect 960 33454 974 33506
rect 1026 33454 1040 33506
rect 960 33440 1040 33454
rect 1120 33506 1200 33520
rect 1120 33454 1134 33506
rect 1186 33454 1200 33506
rect 1120 33440 1200 33454
rect 1280 33506 1360 33520
rect 1280 33454 1294 33506
rect 1346 33454 1360 33506
rect 1280 33440 1360 33454
rect 1440 33506 1520 33520
rect 1440 33454 1454 33506
rect 1506 33454 1520 33506
rect 1440 33440 1520 33454
rect 1600 33506 1680 33520
rect 1600 33454 1614 33506
rect 1666 33454 1680 33506
rect 1600 33440 1680 33454
rect 1760 33506 1840 33520
rect 1760 33454 1774 33506
rect 1826 33454 1840 33506
rect 1760 33440 1840 33454
rect 1920 33506 2000 33520
rect 1920 33454 1934 33506
rect 1986 33454 2000 33506
rect 1920 33440 2000 33454
rect 2080 33506 2160 33520
rect 2080 33454 2094 33506
rect 2146 33454 2160 33506
rect 2080 33440 2160 33454
rect 2240 33506 2320 33520
rect 2240 33454 2254 33506
rect 2306 33454 2320 33506
rect 2240 33440 2320 33454
rect 2400 33506 2480 33520
rect 2400 33454 2414 33506
rect 2466 33454 2480 33506
rect 2400 33440 2480 33454
rect 2560 33506 2640 33520
rect 2560 33454 2574 33506
rect 2626 33454 2640 33506
rect 2560 33440 2640 33454
rect 2720 33506 2800 33520
rect 2720 33454 2734 33506
rect 2786 33454 2800 33506
rect 2720 33440 2800 33454
rect 2880 33506 2960 33520
rect 2880 33454 2894 33506
rect 2946 33454 2960 33506
rect 2880 33440 2960 33454
rect 3040 33506 3120 33520
rect 3040 33454 3054 33506
rect 3106 33454 3120 33506
rect 3040 33440 3120 33454
rect 3200 33506 3280 33520
rect 3200 33454 3214 33506
rect 3266 33454 3280 33506
rect 3200 33440 3280 33454
rect 3360 33506 3440 33520
rect 3360 33454 3374 33506
rect 3426 33454 3440 33506
rect 3360 33440 3440 33454
rect 3520 33506 3600 33520
rect 3520 33454 3534 33506
rect 3586 33454 3600 33506
rect 3520 33440 3600 33454
rect 3680 33506 3760 33520
rect 3680 33454 3694 33506
rect 3746 33454 3760 33506
rect 3680 33440 3760 33454
rect 3840 33506 3920 33520
rect 3840 33454 3854 33506
rect 3906 33454 3920 33506
rect 3840 33440 3920 33454
rect 4000 33506 4080 33520
rect 4000 33454 4014 33506
rect 4066 33454 4080 33506
rect 4000 33440 4080 33454
rect 4160 33506 4240 33520
rect 4160 33454 4174 33506
rect 4226 33454 4240 33506
rect 4160 33440 4240 33454
rect 4320 33506 4400 33520
rect 4320 33454 4334 33506
rect 4386 33454 4400 33506
rect 4320 33440 4400 33454
rect 4480 33506 4560 33520
rect 4480 33454 4494 33506
rect 4546 33454 4560 33506
rect 4480 33440 4560 33454
rect 4640 33506 4720 33520
rect 4640 33454 4654 33506
rect 4706 33454 4720 33506
rect 4640 33440 4720 33454
rect 4800 33506 4880 33520
rect 4800 33454 4814 33506
rect 4866 33454 4880 33506
rect 4800 33440 4880 33454
rect 4960 33506 5040 33520
rect 4960 33454 4974 33506
rect 5026 33454 5040 33506
rect 4960 33440 5040 33454
rect 5120 33506 5200 33520
rect 5120 33454 5134 33506
rect 5186 33454 5200 33506
rect 5120 33440 5200 33454
rect 5280 33506 5360 33520
rect 5280 33454 5294 33506
rect 5346 33454 5360 33506
rect 5280 33440 5360 33454
rect 5440 33506 5520 33520
rect 5440 33454 5454 33506
rect 5506 33454 5520 33506
rect 5440 33440 5520 33454
rect 5600 33506 5680 33520
rect 5600 33454 5614 33506
rect 5666 33454 5680 33506
rect 5600 33440 5680 33454
rect 5760 33506 5840 33520
rect 5760 33454 5774 33506
rect 5826 33454 5840 33506
rect 5760 33440 5840 33454
rect 5920 33506 6000 33520
rect 5920 33454 5934 33506
rect 5986 33454 6000 33506
rect 5920 33440 6000 33454
rect 6080 33506 6160 33520
rect 6080 33454 6094 33506
rect 6146 33454 6160 33506
rect 6080 33440 6160 33454
rect 6240 33506 6320 33520
rect 6240 33454 6254 33506
rect 6306 33454 6320 33506
rect 6240 33440 6320 33454
rect 6400 33506 6480 33520
rect 6400 33454 6414 33506
rect 6466 33454 6480 33506
rect 6400 33440 6480 33454
rect 6560 33506 6640 33520
rect 6560 33454 6574 33506
rect 6626 33454 6640 33506
rect 6560 33440 6640 33454
rect 6720 33506 6800 33520
rect 6720 33454 6734 33506
rect 6786 33454 6800 33506
rect 6720 33440 6800 33454
rect 6880 33506 6960 33520
rect 6880 33454 6894 33506
rect 6946 33454 6960 33506
rect 6880 33440 6960 33454
rect 7040 33506 7120 33520
rect 7040 33454 7054 33506
rect 7106 33454 7120 33506
rect 7040 33440 7120 33454
rect 7200 33506 7280 33520
rect 7200 33454 7214 33506
rect 7266 33454 7280 33506
rect 7200 33440 7280 33454
rect 7360 33506 7440 33520
rect 7360 33454 7374 33506
rect 7426 33454 7440 33506
rect 7360 33440 7440 33454
rect 7520 33506 7600 33520
rect 7520 33454 7534 33506
rect 7586 33454 7600 33506
rect 7520 33440 7600 33454
rect 7680 33506 7760 33520
rect 7680 33454 7694 33506
rect 7746 33454 7760 33506
rect 7680 33440 7760 33454
rect 7840 33506 7920 33520
rect 7840 33454 7854 33506
rect 7906 33454 7920 33506
rect 7840 33440 7920 33454
rect 8000 33506 8080 33520
rect 8000 33454 8014 33506
rect 8066 33454 8080 33506
rect 8000 33440 8080 33454
rect 8160 33506 8240 33520
rect 8160 33454 8174 33506
rect 8226 33454 8240 33506
rect 8160 33440 8240 33454
rect 8320 33506 8400 33520
rect 8320 33454 8334 33506
rect 8386 33454 8400 33506
rect 8320 33440 8400 33454
rect 12480 33506 12560 33520
rect 12480 33454 12494 33506
rect 12546 33454 12560 33506
rect 12480 33440 12560 33454
rect 12640 33506 12720 33520
rect 12640 33454 12654 33506
rect 12706 33454 12720 33506
rect 12640 33440 12720 33454
rect 12800 33506 12880 33520
rect 12800 33454 12814 33506
rect 12866 33454 12880 33506
rect 12800 33440 12880 33454
rect 12960 33506 13040 33520
rect 12960 33454 12974 33506
rect 13026 33454 13040 33506
rect 12960 33440 13040 33454
rect 13120 33506 13200 33520
rect 13120 33454 13134 33506
rect 13186 33454 13200 33506
rect 13120 33440 13200 33454
rect 13280 33506 13360 33520
rect 13280 33454 13294 33506
rect 13346 33454 13360 33506
rect 13280 33440 13360 33454
rect 13440 33506 13520 33520
rect 13440 33454 13454 33506
rect 13506 33454 13520 33506
rect 13440 33440 13520 33454
rect 13600 33506 13680 33520
rect 13600 33454 13614 33506
rect 13666 33454 13680 33506
rect 13600 33440 13680 33454
rect 13760 33506 13840 33520
rect 13760 33454 13774 33506
rect 13826 33454 13840 33506
rect 13760 33440 13840 33454
rect 13920 33506 14000 33520
rect 13920 33454 13934 33506
rect 13986 33454 14000 33506
rect 13920 33440 14000 33454
rect 14080 33506 14160 33520
rect 14080 33454 14094 33506
rect 14146 33454 14160 33506
rect 14080 33440 14160 33454
rect 14240 33506 14320 33520
rect 14240 33454 14254 33506
rect 14306 33454 14320 33506
rect 14240 33440 14320 33454
rect 14400 33506 14480 33520
rect 14400 33454 14414 33506
rect 14466 33454 14480 33506
rect 14400 33440 14480 33454
rect 14560 33506 14640 33520
rect 14560 33454 14574 33506
rect 14626 33454 14640 33506
rect 14560 33440 14640 33454
rect 14720 33506 14800 33520
rect 14720 33454 14734 33506
rect 14786 33454 14800 33506
rect 14720 33440 14800 33454
rect 14880 33506 14960 33520
rect 14880 33454 14894 33506
rect 14946 33454 14960 33506
rect 14880 33440 14960 33454
rect 15040 33506 15120 33520
rect 15040 33454 15054 33506
rect 15106 33454 15120 33506
rect 15040 33440 15120 33454
rect 15200 33506 15280 33520
rect 15200 33454 15214 33506
rect 15266 33454 15280 33506
rect 15200 33440 15280 33454
rect 15360 33506 15440 33520
rect 15360 33454 15374 33506
rect 15426 33454 15440 33506
rect 15360 33440 15440 33454
rect 15520 33506 15600 33520
rect 15520 33454 15534 33506
rect 15586 33454 15600 33506
rect 15520 33440 15600 33454
rect 15680 33506 15760 33520
rect 15680 33454 15694 33506
rect 15746 33454 15760 33506
rect 15680 33440 15760 33454
rect 15840 33506 15920 33520
rect 15840 33454 15854 33506
rect 15906 33454 15920 33506
rect 15840 33440 15920 33454
rect 16000 33506 16080 33520
rect 16000 33454 16014 33506
rect 16066 33454 16080 33506
rect 16000 33440 16080 33454
rect 16160 33506 16240 33520
rect 16160 33454 16174 33506
rect 16226 33454 16240 33506
rect 16160 33440 16240 33454
rect 16320 33506 16400 33520
rect 16320 33454 16334 33506
rect 16386 33454 16400 33506
rect 16320 33440 16400 33454
rect 16480 33506 16560 33520
rect 16480 33454 16494 33506
rect 16546 33454 16560 33506
rect 16480 33440 16560 33454
rect 16640 33506 16720 33520
rect 16640 33454 16654 33506
rect 16706 33454 16720 33506
rect 16640 33440 16720 33454
rect 16800 33506 16880 33520
rect 16800 33454 16814 33506
rect 16866 33454 16880 33506
rect 16800 33440 16880 33454
rect 16960 33506 17040 33520
rect 16960 33454 16974 33506
rect 17026 33454 17040 33506
rect 16960 33440 17040 33454
rect 17120 33506 17200 33520
rect 17120 33454 17134 33506
rect 17186 33454 17200 33506
rect 17120 33440 17200 33454
rect 17280 33506 17360 33520
rect 17280 33454 17294 33506
rect 17346 33454 17360 33506
rect 17280 33440 17360 33454
rect 17440 33506 17520 33520
rect 17440 33454 17454 33506
rect 17506 33454 17520 33506
rect 17440 33440 17520 33454
rect 17600 33506 17680 33520
rect 17600 33454 17614 33506
rect 17666 33454 17680 33506
rect 17600 33440 17680 33454
rect 17760 33506 17840 33520
rect 17760 33454 17774 33506
rect 17826 33454 17840 33506
rect 17760 33440 17840 33454
rect 17920 33506 18000 33520
rect 17920 33454 17934 33506
rect 17986 33454 18000 33506
rect 17920 33440 18000 33454
rect 18080 33506 18160 33520
rect 18080 33454 18094 33506
rect 18146 33454 18160 33506
rect 18080 33440 18160 33454
rect 18240 33506 18320 33520
rect 18240 33454 18254 33506
rect 18306 33454 18320 33506
rect 18240 33440 18320 33454
rect 18400 33506 18480 33520
rect 18400 33454 18414 33506
rect 18466 33454 18480 33506
rect 18400 33440 18480 33454
rect 18560 33506 18640 33520
rect 18560 33454 18574 33506
rect 18626 33454 18640 33506
rect 18560 33440 18640 33454
rect 18720 33506 18800 33520
rect 18720 33454 18734 33506
rect 18786 33454 18800 33506
rect 18720 33440 18800 33454
rect 18880 33506 18960 33520
rect 18880 33454 18894 33506
rect 18946 33454 18960 33506
rect 18880 33440 18960 33454
rect 23120 33506 23200 33520
rect 23120 33454 23134 33506
rect 23186 33454 23200 33506
rect 23120 33440 23200 33454
rect 23280 33506 23360 33520
rect 23280 33454 23294 33506
rect 23346 33454 23360 33506
rect 23280 33440 23360 33454
rect 23440 33506 23520 33520
rect 23440 33454 23454 33506
rect 23506 33454 23520 33506
rect 23440 33440 23520 33454
rect 23600 33506 23680 33520
rect 23600 33454 23614 33506
rect 23666 33454 23680 33506
rect 23600 33440 23680 33454
rect 23760 33506 23840 33520
rect 23760 33454 23774 33506
rect 23826 33454 23840 33506
rect 23760 33440 23840 33454
rect 23920 33506 24000 33520
rect 23920 33454 23934 33506
rect 23986 33454 24000 33506
rect 23920 33440 24000 33454
rect 24080 33506 24160 33520
rect 24080 33454 24094 33506
rect 24146 33454 24160 33506
rect 24080 33440 24160 33454
rect 24240 33506 24320 33520
rect 24240 33454 24254 33506
rect 24306 33454 24320 33506
rect 24240 33440 24320 33454
rect 24400 33506 24480 33520
rect 24400 33454 24414 33506
rect 24466 33454 24480 33506
rect 24400 33440 24480 33454
rect 24560 33506 24640 33520
rect 24560 33454 24574 33506
rect 24626 33454 24640 33506
rect 24560 33440 24640 33454
rect 24720 33506 24800 33520
rect 24720 33454 24734 33506
rect 24786 33454 24800 33506
rect 24720 33440 24800 33454
rect 24880 33506 24960 33520
rect 24880 33454 24894 33506
rect 24946 33454 24960 33506
rect 24880 33440 24960 33454
rect 25040 33506 25120 33520
rect 25040 33454 25054 33506
rect 25106 33454 25120 33506
rect 25040 33440 25120 33454
rect 25200 33506 25280 33520
rect 25200 33454 25214 33506
rect 25266 33454 25280 33506
rect 25200 33440 25280 33454
rect 25360 33506 25440 33520
rect 25360 33454 25374 33506
rect 25426 33454 25440 33506
rect 25360 33440 25440 33454
rect 25520 33506 25600 33520
rect 25520 33454 25534 33506
rect 25586 33454 25600 33506
rect 25520 33440 25600 33454
rect 25680 33506 25760 33520
rect 25680 33454 25694 33506
rect 25746 33454 25760 33506
rect 25680 33440 25760 33454
rect 25840 33506 25920 33520
rect 25840 33454 25854 33506
rect 25906 33454 25920 33506
rect 25840 33440 25920 33454
rect 26000 33506 26080 33520
rect 26000 33454 26014 33506
rect 26066 33454 26080 33506
rect 26000 33440 26080 33454
rect 26160 33506 26240 33520
rect 26160 33454 26174 33506
rect 26226 33454 26240 33506
rect 26160 33440 26240 33454
rect 26320 33506 26400 33520
rect 26320 33454 26334 33506
rect 26386 33454 26400 33506
rect 26320 33440 26400 33454
rect 26480 33506 26560 33520
rect 26480 33454 26494 33506
rect 26546 33454 26560 33506
rect 26480 33440 26560 33454
rect 26640 33506 26720 33520
rect 26640 33454 26654 33506
rect 26706 33454 26720 33506
rect 26640 33440 26720 33454
rect 26800 33506 26880 33520
rect 26800 33454 26814 33506
rect 26866 33454 26880 33506
rect 26800 33440 26880 33454
rect 26960 33506 27040 33520
rect 26960 33454 26974 33506
rect 27026 33454 27040 33506
rect 26960 33440 27040 33454
rect 27120 33506 27200 33520
rect 27120 33454 27134 33506
rect 27186 33454 27200 33506
rect 27120 33440 27200 33454
rect 27280 33506 27360 33520
rect 27280 33454 27294 33506
rect 27346 33454 27360 33506
rect 27280 33440 27360 33454
rect 27440 33506 27520 33520
rect 27440 33454 27454 33506
rect 27506 33454 27520 33506
rect 27440 33440 27520 33454
rect 27600 33506 27680 33520
rect 27600 33454 27614 33506
rect 27666 33454 27680 33506
rect 27600 33440 27680 33454
rect 27760 33506 27840 33520
rect 27760 33454 27774 33506
rect 27826 33454 27840 33506
rect 27760 33440 27840 33454
rect 27920 33506 28000 33520
rect 27920 33454 27934 33506
rect 27986 33454 28000 33506
rect 27920 33440 28000 33454
rect 28080 33506 28160 33520
rect 28080 33454 28094 33506
rect 28146 33454 28160 33506
rect 28080 33440 28160 33454
rect 28240 33506 28320 33520
rect 28240 33454 28254 33506
rect 28306 33454 28320 33506
rect 28240 33440 28320 33454
rect 28400 33506 28480 33520
rect 28400 33454 28414 33506
rect 28466 33454 28480 33506
rect 28400 33440 28480 33454
rect 28560 33506 28640 33520
rect 28560 33454 28574 33506
rect 28626 33454 28640 33506
rect 28560 33440 28640 33454
rect 28720 33506 28800 33520
rect 28720 33454 28734 33506
rect 28786 33454 28800 33506
rect 28720 33440 28800 33454
rect 28880 33506 28960 33520
rect 28880 33454 28894 33506
rect 28946 33454 28960 33506
rect 28880 33440 28960 33454
rect 29040 33506 29120 33520
rect 29040 33454 29054 33506
rect 29106 33454 29120 33506
rect 29040 33440 29120 33454
rect 29200 33506 29280 33520
rect 29200 33454 29214 33506
rect 29266 33454 29280 33506
rect 29200 33440 29280 33454
rect 29360 33506 29440 33520
rect 29360 33454 29374 33506
rect 29426 33454 29440 33506
rect 29360 33440 29440 33454
rect 33520 33506 33600 33520
rect 33520 33454 33534 33506
rect 33586 33454 33600 33506
rect 33520 33440 33600 33454
rect 33680 33506 33760 33520
rect 33680 33454 33694 33506
rect 33746 33454 33760 33506
rect 33680 33440 33760 33454
rect 33840 33506 33920 33520
rect 33840 33454 33854 33506
rect 33906 33454 33920 33506
rect 33840 33440 33920 33454
rect 34000 33506 34080 33520
rect 34000 33454 34014 33506
rect 34066 33454 34080 33506
rect 34000 33440 34080 33454
rect 34160 33506 34240 33520
rect 34160 33454 34174 33506
rect 34226 33454 34240 33506
rect 34160 33440 34240 33454
rect 34320 33506 34400 33520
rect 34320 33454 34334 33506
rect 34386 33454 34400 33506
rect 34320 33440 34400 33454
rect 34480 33506 34560 33520
rect 34480 33454 34494 33506
rect 34546 33454 34560 33506
rect 34480 33440 34560 33454
rect 34640 33506 34720 33520
rect 34640 33454 34654 33506
rect 34706 33454 34720 33506
rect 34640 33440 34720 33454
rect 34800 33506 34880 33520
rect 34800 33454 34814 33506
rect 34866 33454 34880 33506
rect 34800 33440 34880 33454
rect 34960 33506 35040 33520
rect 34960 33454 34974 33506
rect 35026 33454 35040 33506
rect 34960 33440 35040 33454
rect 35120 33506 35200 33520
rect 35120 33454 35134 33506
rect 35186 33454 35200 33506
rect 35120 33440 35200 33454
rect 35280 33506 35360 33520
rect 35280 33454 35294 33506
rect 35346 33454 35360 33506
rect 35280 33440 35360 33454
rect 35440 33506 35520 33520
rect 35440 33454 35454 33506
rect 35506 33454 35520 33506
rect 35440 33440 35520 33454
rect 35600 33506 35680 33520
rect 35600 33454 35614 33506
rect 35666 33454 35680 33506
rect 35600 33440 35680 33454
rect 35760 33506 35840 33520
rect 35760 33454 35774 33506
rect 35826 33454 35840 33506
rect 35760 33440 35840 33454
rect 35920 33506 36000 33520
rect 35920 33454 35934 33506
rect 35986 33454 36000 33506
rect 35920 33440 36000 33454
rect 36080 33506 36160 33520
rect 36080 33454 36094 33506
rect 36146 33454 36160 33506
rect 36080 33440 36160 33454
rect 36240 33506 36320 33520
rect 36240 33454 36254 33506
rect 36306 33454 36320 33506
rect 36240 33440 36320 33454
rect 36400 33506 36480 33520
rect 36400 33454 36414 33506
rect 36466 33454 36480 33506
rect 36400 33440 36480 33454
rect 36560 33506 36640 33520
rect 36560 33454 36574 33506
rect 36626 33454 36640 33506
rect 36560 33440 36640 33454
rect 36720 33506 36800 33520
rect 36720 33454 36734 33506
rect 36786 33454 36800 33506
rect 36720 33440 36800 33454
rect 36880 33506 36960 33520
rect 36880 33454 36894 33506
rect 36946 33454 36960 33506
rect 36880 33440 36960 33454
rect 37040 33506 37120 33520
rect 37040 33454 37054 33506
rect 37106 33454 37120 33506
rect 37040 33440 37120 33454
rect 37200 33506 37280 33520
rect 37200 33454 37214 33506
rect 37266 33454 37280 33506
rect 37200 33440 37280 33454
rect 37360 33506 37440 33520
rect 37360 33454 37374 33506
rect 37426 33454 37440 33506
rect 37360 33440 37440 33454
rect 37520 33506 37600 33520
rect 37520 33454 37534 33506
rect 37586 33454 37600 33506
rect 37520 33440 37600 33454
rect 37680 33506 37760 33520
rect 37680 33454 37694 33506
rect 37746 33454 37760 33506
rect 37680 33440 37760 33454
rect 37840 33506 37920 33520
rect 37840 33454 37854 33506
rect 37906 33454 37920 33506
rect 37840 33440 37920 33454
rect 38000 33506 38080 33520
rect 38000 33454 38014 33506
rect 38066 33454 38080 33506
rect 38000 33440 38080 33454
rect 38160 33506 38240 33520
rect 38160 33454 38174 33506
rect 38226 33454 38240 33506
rect 38160 33440 38240 33454
rect 38320 33506 38400 33520
rect 38320 33454 38334 33506
rect 38386 33454 38400 33506
rect 38320 33440 38400 33454
rect 38480 33506 38560 33520
rect 38480 33454 38494 33506
rect 38546 33454 38560 33506
rect 38480 33440 38560 33454
rect 38640 33506 38720 33520
rect 38640 33454 38654 33506
rect 38706 33454 38720 33506
rect 38640 33440 38720 33454
rect 38800 33506 38880 33520
rect 38800 33454 38814 33506
rect 38866 33454 38880 33506
rect 38800 33440 38880 33454
rect 38960 33506 39040 33520
rect 38960 33454 38974 33506
rect 39026 33454 39040 33506
rect 38960 33440 39040 33454
rect 39120 33506 39200 33520
rect 39120 33454 39134 33506
rect 39186 33454 39200 33506
rect 39120 33440 39200 33454
rect 39280 33506 39360 33520
rect 39280 33454 39294 33506
rect 39346 33454 39360 33506
rect 39280 33440 39360 33454
rect 39440 33506 39520 33520
rect 39440 33454 39454 33506
rect 39506 33454 39520 33506
rect 39440 33440 39520 33454
rect 39600 33506 39680 33520
rect 39600 33454 39614 33506
rect 39666 33454 39680 33506
rect 39600 33440 39680 33454
rect 39760 33506 39840 33520
rect 39760 33454 39774 33506
rect 39826 33454 39840 33506
rect 39760 33440 39840 33454
rect 39920 33506 40000 33520
rect 39920 33454 39934 33506
rect 39986 33454 40000 33506
rect 39920 33440 40000 33454
rect 40080 33506 40160 33520
rect 40080 33454 40094 33506
rect 40146 33454 40160 33506
rect 40080 33440 40160 33454
rect 40240 33506 40320 33520
rect 40240 33454 40254 33506
rect 40306 33454 40320 33506
rect 40240 33440 40320 33454
rect 40400 33506 40480 33520
rect 40400 33454 40414 33506
rect 40466 33454 40480 33506
rect 40400 33440 40480 33454
rect 40560 33506 40640 33520
rect 40560 33454 40574 33506
rect 40626 33454 40640 33506
rect 40560 33440 40640 33454
rect 40720 33506 40800 33520
rect 40720 33454 40734 33506
rect 40786 33454 40800 33506
rect 40720 33440 40800 33454
rect 40880 33506 40960 33520
rect 40880 33454 40894 33506
rect 40946 33454 40960 33506
rect 40880 33440 40960 33454
rect 41040 33506 41120 33520
rect 41040 33454 41054 33506
rect 41106 33454 41120 33506
rect 41040 33440 41120 33454
rect 41200 33506 41280 33520
rect 41200 33454 41214 33506
rect 41266 33454 41280 33506
rect 41200 33440 41280 33454
rect 41360 33506 41440 33520
rect 41360 33454 41374 33506
rect 41426 33454 41440 33506
rect 41360 33440 41440 33454
rect 41520 33506 41600 33520
rect 41520 33454 41534 33506
rect 41586 33454 41600 33506
rect 41520 33440 41600 33454
rect 41680 33506 41760 33520
rect 41680 33454 41694 33506
rect 41746 33454 41760 33506
rect 41680 33440 41760 33454
rect 41840 33506 41920 33520
rect 41840 33454 41854 33506
rect 41906 33454 41920 33506
rect 41840 33440 41920 33454
rect 0 33346 80 33360
rect 0 33294 14 33346
rect 66 33294 80 33346
rect 0 33280 80 33294
rect 160 33346 240 33360
rect 160 33294 174 33346
rect 226 33294 240 33346
rect 160 33280 240 33294
rect 320 33346 400 33360
rect 320 33294 334 33346
rect 386 33294 400 33346
rect 320 33280 400 33294
rect 480 33346 560 33360
rect 480 33294 494 33346
rect 546 33294 560 33346
rect 480 33280 560 33294
rect 640 33346 720 33360
rect 640 33294 654 33346
rect 706 33294 720 33346
rect 640 33280 720 33294
rect 800 33346 880 33360
rect 800 33294 814 33346
rect 866 33294 880 33346
rect 800 33280 880 33294
rect 960 33346 1040 33360
rect 960 33294 974 33346
rect 1026 33294 1040 33346
rect 960 33280 1040 33294
rect 1120 33346 1200 33360
rect 1120 33294 1134 33346
rect 1186 33294 1200 33346
rect 1120 33280 1200 33294
rect 1280 33346 1360 33360
rect 1280 33294 1294 33346
rect 1346 33294 1360 33346
rect 1280 33280 1360 33294
rect 1440 33346 1520 33360
rect 1440 33294 1454 33346
rect 1506 33294 1520 33346
rect 1440 33280 1520 33294
rect 1600 33346 1680 33360
rect 1600 33294 1614 33346
rect 1666 33294 1680 33346
rect 1600 33280 1680 33294
rect 1760 33346 1840 33360
rect 1760 33294 1774 33346
rect 1826 33294 1840 33346
rect 1760 33280 1840 33294
rect 1920 33346 2000 33360
rect 1920 33294 1934 33346
rect 1986 33294 2000 33346
rect 1920 33280 2000 33294
rect 2080 33346 2160 33360
rect 2080 33294 2094 33346
rect 2146 33294 2160 33346
rect 2080 33280 2160 33294
rect 2240 33346 2320 33360
rect 2240 33294 2254 33346
rect 2306 33294 2320 33346
rect 2240 33280 2320 33294
rect 2400 33346 2480 33360
rect 2400 33294 2414 33346
rect 2466 33294 2480 33346
rect 2400 33280 2480 33294
rect 2560 33346 2640 33360
rect 2560 33294 2574 33346
rect 2626 33294 2640 33346
rect 2560 33280 2640 33294
rect 2720 33346 2800 33360
rect 2720 33294 2734 33346
rect 2786 33294 2800 33346
rect 2720 33280 2800 33294
rect 2880 33346 2960 33360
rect 2880 33294 2894 33346
rect 2946 33294 2960 33346
rect 2880 33280 2960 33294
rect 3040 33346 3120 33360
rect 3040 33294 3054 33346
rect 3106 33294 3120 33346
rect 3040 33280 3120 33294
rect 3200 33346 3280 33360
rect 3200 33294 3214 33346
rect 3266 33294 3280 33346
rect 3200 33280 3280 33294
rect 3360 33346 3440 33360
rect 3360 33294 3374 33346
rect 3426 33294 3440 33346
rect 3360 33280 3440 33294
rect 3520 33346 3600 33360
rect 3520 33294 3534 33346
rect 3586 33294 3600 33346
rect 3520 33280 3600 33294
rect 3680 33346 3760 33360
rect 3680 33294 3694 33346
rect 3746 33294 3760 33346
rect 3680 33280 3760 33294
rect 3840 33346 3920 33360
rect 3840 33294 3854 33346
rect 3906 33294 3920 33346
rect 3840 33280 3920 33294
rect 4000 33346 4080 33360
rect 4000 33294 4014 33346
rect 4066 33294 4080 33346
rect 4000 33280 4080 33294
rect 4160 33346 4240 33360
rect 4160 33294 4174 33346
rect 4226 33294 4240 33346
rect 4160 33280 4240 33294
rect 4320 33346 4400 33360
rect 4320 33294 4334 33346
rect 4386 33294 4400 33346
rect 4320 33280 4400 33294
rect 4480 33346 4560 33360
rect 4480 33294 4494 33346
rect 4546 33294 4560 33346
rect 4480 33280 4560 33294
rect 4640 33346 4720 33360
rect 4640 33294 4654 33346
rect 4706 33294 4720 33346
rect 4640 33280 4720 33294
rect 4800 33346 4880 33360
rect 4800 33294 4814 33346
rect 4866 33294 4880 33346
rect 4800 33280 4880 33294
rect 4960 33346 5040 33360
rect 4960 33294 4974 33346
rect 5026 33294 5040 33346
rect 4960 33280 5040 33294
rect 5120 33346 5200 33360
rect 5120 33294 5134 33346
rect 5186 33294 5200 33346
rect 5120 33280 5200 33294
rect 5280 33346 5360 33360
rect 5280 33294 5294 33346
rect 5346 33294 5360 33346
rect 5280 33280 5360 33294
rect 5440 33346 5520 33360
rect 5440 33294 5454 33346
rect 5506 33294 5520 33346
rect 5440 33280 5520 33294
rect 5600 33346 5680 33360
rect 5600 33294 5614 33346
rect 5666 33294 5680 33346
rect 5600 33280 5680 33294
rect 5760 33346 5840 33360
rect 5760 33294 5774 33346
rect 5826 33294 5840 33346
rect 5760 33280 5840 33294
rect 5920 33346 6000 33360
rect 5920 33294 5934 33346
rect 5986 33294 6000 33346
rect 5920 33280 6000 33294
rect 6080 33346 6160 33360
rect 6080 33294 6094 33346
rect 6146 33294 6160 33346
rect 6080 33280 6160 33294
rect 6240 33346 6320 33360
rect 6240 33294 6254 33346
rect 6306 33294 6320 33346
rect 6240 33280 6320 33294
rect 6400 33346 6480 33360
rect 6400 33294 6414 33346
rect 6466 33294 6480 33346
rect 6400 33280 6480 33294
rect 6560 33346 6640 33360
rect 6560 33294 6574 33346
rect 6626 33294 6640 33346
rect 6560 33280 6640 33294
rect 6720 33346 6800 33360
rect 6720 33294 6734 33346
rect 6786 33294 6800 33346
rect 6720 33280 6800 33294
rect 6880 33346 6960 33360
rect 6880 33294 6894 33346
rect 6946 33294 6960 33346
rect 6880 33280 6960 33294
rect 7040 33346 7120 33360
rect 7040 33294 7054 33346
rect 7106 33294 7120 33346
rect 7040 33280 7120 33294
rect 7200 33346 7280 33360
rect 7200 33294 7214 33346
rect 7266 33294 7280 33346
rect 7200 33280 7280 33294
rect 7360 33346 7440 33360
rect 7360 33294 7374 33346
rect 7426 33294 7440 33346
rect 7360 33280 7440 33294
rect 7520 33346 7600 33360
rect 7520 33294 7534 33346
rect 7586 33294 7600 33346
rect 7520 33280 7600 33294
rect 7680 33346 7760 33360
rect 7680 33294 7694 33346
rect 7746 33294 7760 33346
rect 7680 33280 7760 33294
rect 7840 33346 7920 33360
rect 7840 33294 7854 33346
rect 7906 33294 7920 33346
rect 7840 33280 7920 33294
rect 8000 33346 8080 33360
rect 8000 33294 8014 33346
rect 8066 33294 8080 33346
rect 8000 33280 8080 33294
rect 8160 33346 8240 33360
rect 8160 33294 8174 33346
rect 8226 33294 8240 33346
rect 8160 33280 8240 33294
rect 8320 33346 8400 33360
rect 8320 33294 8334 33346
rect 8386 33294 8400 33346
rect 8320 33280 8400 33294
rect 12480 33346 12560 33360
rect 12480 33294 12494 33346
rect 12546 33294 12560 33346
rect 12480 33280 12560 33294
rect 12640 33346 12720 33360
rect 12640 33294 12654 33346
rect 12706 33294 12720 33346
rect 12640 33280 12720 33294
rect 12800 33346 12880 33360
rect 12800 33294 12814 33346
rect 12866 33294 12880 33346
rect 12800 33280 12880 33294
rect 12960 33346 13040 33360
rect 12960 33294 12974 33346
rect 13026 33294 13040 33346
rect 12960 33280 13040 33294
rect 13120 33346 13200 33360
rect 13120 33294 13134 33346
rect 13186 33294 13200 33346
rect 13120 33280 13200 33294
rect 13280 33346 13360 33360
rect 13280 33294 13294 33346
rect 13346 33294 13360 33346
rect 13280 33280 13360 33294
rect 13440 33346 13520 33360
rect 13440 33294 13454 33346
rect 13506 33294 13520 33346
rect 13440 33280 13520 33294
rect 13600 33346 13680 33360
rect 13600 33294 13614 33346
rect 13666 33294 13680 33346
rect 13600 33280 13680 33294
rect 13760 33346 13840 33360
rect 13760 33294 13774 33346
rect 13826 33294 13840 33346
rect 13760 33280 13840 33294
rect 13920 33346 14000 33360
rect 13920 33294 13934 33346
rect 13986 33294 14000 33346
rect 13920 33280 14000 33294
rect 14080 33346 14160 33360
rect 14080 33294 14094 33346
rect 14146 33294 14160 33346
rect 14080 33280 14160 33294
rect 14240 33346 14320 33360
rect 14240 33294 14254 33346
rect 14306 33294 14320 33346
rect 14240 33280 14320 33294
rect 14400 33346 14480 33360
rect 14400 33294 14414 33346
rect 14466 33294 14480 33346
rect 14400 33280 14480 33294
rect 14560 33346 14640 33360
rect 14560 33294 14574 33346
rect 14626 33294 14640 33346
rect 14560 33280 14640 33294
rect 14720 33346 14800 33360
rect 14720 33294 14734 33346
rect 14786 33294 14800 33346
rect 14720 33280 14800 33294
rect 14880 33346 14960 33360
rect 14880 33294 14894 33346
rect 14946 33294 14960 33346
rect 14880 33280 14960 33294
rect 15040 33346 15120 33360
rect 15040 33294 15054 33346
rect 15106 33294 15120 33346
rect 15040 33280 15120 33294
rect 15200 33346 15280 33360
rect 15200 33294 15214 33346
rect 15266 33294 15280 33346
rect 15200 33280 15280 33294
rect 15360 33346 15440 33360
rect 15360 33294 15374 33346
rect 15426 33294 15440 33346
rect 15360 33280 15440 33294
rect 15520 33346 15600 33360
rect 15520 33294 15534 33346
rect 15586 33294 15600 33346
rect 15520 33280 15600 33294
rect 15680 33346 15760 33360
rect 15680 33294 15694 33346
rect 15746 33294 15760 33346
rect 15680 33280 15760 33294
rect 15840 33346 15920 33360
rect 15840 33294 15854 33346
rect 15906 33294 15920 33346
rect 15840 33280 15920 33294
rect 16000 33346 16080 33360
rect 16000 33294 16014 33346
rect 16066 33294 16080 33346
rect 16000 33280 16080 33294
rect 16160 33346 16240 33360
rect 16160 33294 16174 33346
rect 16226 33294 16240 33346
rect 16160 33280 16240 33294
rect 16320 33346 16400 33360
rect 16320 33294 16334 33346
rect 16386 33294 16400 33346
rect 16320 33280 16400 33294
rect 16480 33346 16560 33360
rect 16480 33294 16494 33346
rect 16546 33294 16560 33346
rect 16480 33280 16560 33294
rect 16640 33346 16720 33360
rect 16640 33294 16654 33346
rect 16706 33294 16720 33346
rect 16640 33280 16720 33294
rect 16800 33346 16880 33360
rect 16800 33294 16814 33346
rect 16866 33294 16880 33346
rect 16800 33280 16880 33294
rect 16960 33346 17040 33360
rect 16960 33294 16974 33346
rect 17026 33294 17040 33346
rect 16960 33280 17040 33294
rect 17120 33346 17200 33360
rect 17120 33294 17134 33346
rect 17186 33294 17200 33346
rect 17120 33280 17200 33294
rect 17280 33346 17360 33360
rect 17280 33294 17294 33346
rect 17346 33294 17360 33346
rect 17280 33280 17360 33294
rect 17440 33346 17520 33360
rect 17440 33294 17454 33346
rect 17506 33294 17520 33346
rect 17440 33280 17520 33294
rect 17600 33346 17680 33360
rect 17600 33294 17614 33346
rect 17666 33294 17680 33346
rect 17600 33280 17680 33294
rect 17760 33346 17840 33360
rect 17760 33294 17774 33346
rect 17826 33294 17840 33346
rect 17760 33280 17840 33294
rect 17920 33346 18000 33360
rect 17920 33294 17934 33346
rect 17986 33294 18000 33346
rect 17920 33280 18000 33294
rect 18080 33346 18160 33360
rect 18080 33294 18094 33346
rect 18146 33294 18160 33346
rect 18080 33280 18160 33294
rect 18240 33346 18320 33360
rect 18240 33294 18254 33346
rect 18306 33294 18320 33346
rect 18240 33280 18320 33294
rect 18400 33346 18480 33360
rect 18400 33294 18414 33346
rect 18466 33294 18480 33346
rect 18400 33280 18480 33294
rect 18560 33346 18640 33360
rect 18560 33294 18574 33346
rect 18626 33294 18640 33346
rect 18560 33280 18640 33294
rect 18720 33346 18800 33360
rect 18720 33294 18734 33346
rect 18786 33294 18800 33346
rect 18720 33280 18800 33294
rect 18880 33346 18960 33360
rect 18880 33294 18894 33346
rect 18946 33294 18960 33346
rect 18880 33280 18960 33294
rect 23120 33346 23200 33360
rect 23120 33294 23134 33346
rect 23186 33294 23200 33346
rect 23120 33280 23200 33294
rect 23280 33346 23360 33360
rect 23280 33294 23294 33346
rect 23346 33294 23360 33346
rect 23280 33280 23360 33294
rect 23440 33346 23520 33360
rect 23440 33294 23454 33346
rect 23506 33294 23520 33346
rect 23440 33280 23520 33294
rect 23600 33346 23680 33360
rect 23600 33294 23614 33346
rect 23666 33294 23680 33346
rect 23600 33280 23680 33294
rect 23760 33346 23840 33360
rect 23760 33294 23774 33346
rect 23826 33294 23840 33346
rect 23760 33280 23840 33294
rect 23920 33346 24000 33360
rect 23920 33294 23934 33346
rect 23986 33294 24000 33346
rect 23920 33280 24000 33294
rect 24080 33346 24160 33360
rect 24080 33294 24094 33346
rect 24146 33294 24160 33346
rect 24080 33280 24160 33294
rect 24240 33346 24320 33360
rect 24240 33294 24254 33346
rect 24306 33294 24320 33346
rect 24240 33280 24320 33294
rect 24400 33346 24480 33360
rect 24400 33294 24414 33346
rect 24466 33294 24480 33346
rect 24400 33280 24480 33294
rect 24560 33346 24640 33360
rect 24560 33294 24574 33346
rect 24626 33294 24640 33346
rect 24560 33280 24640 33294
rect 24720 33346 24800 33360
rect 24720 33294 24734 33346
rect 24786 33294 24800 33346
rect 24720 33280 24800 33294
rect 24880 33346 24960 33360
rect 24880 33294 24894 33346
rect 24946 33294 24960 33346
rect 24880 33280 24960 33294
rect 25040 33346 25120 33360
rect 25040 33294 25054 33346
rect 25106 33294 25120 33346
rect 25040 33280 25120 33294
rect 25200 33346 25280 33360
rect 25200 33294 25214 33346
rect 25266 33294 25280 33346
rect 25200 33280 25280 33294
rect 25360 33346 25440 33360
rect 25360 33294 25374 33346
rect 25426 33294 25440 33346
rect 25360 33280 25440 33294
rect 25520 33346 25600 33360
rect 25520 33294 25534 33346
rect 25586 33294 25600 33346
rect 25520 33280 25600 33294
rect 25680 33346 25760 33360
rect 25680 33294 25694 33346
rect 25746 33294 25760 33346
rect 25680 33280 25760 33294
rect 25840 33346 25920 33360
rect 25840 33294 25854 33346
rect 25906 33294 25920 33346
rect 25840 33280 25920 33294
rect 26000 33346 26080 33360
rect 26000 33294 26014 33346
rect 26066 33294 26080 33346
rect 26000 33280 26080 33294
rect 26160 33346 26240 33360
rect 26160 33294 26174 33346
rect 26226 33294 26240 33346
rect 26160 33280 26240 33294
rect 26320 33346 26400 33360
rect 26320 33294 26334 33346
rect 26386 33294 26400 33346
rect 26320 33280 26400 33294
rect 26480 33346 26560 33360
rect 26480 33294 26494 33346
rect 26546 33294 26560 33346
rect 26480 33280 26560 33294
rect 26640 33346 26720 33360
rect 26640 33294 26654 33346
rect 26706 33294 26720 33346
rect 26640 33280 26720 33294
rect 26800 33346 26880 33360
rect 26800 33294 26814 33346
rect 26866 33294 26880 33346
rect 26800 33280 26880 33294
rect 26960 33346 27040 33360
rect 26960 33294 26974 33346
rect 27026 33294 27040 33346
rect 26960 33280 27040 33294
rect 27120 33346 27200 33360
rect 27120 33294 27134 33346
rect 27186 33294 27200 33346
rect 27120 33280 27200 33294
rect 27280 33346 27360 33360
rect 27280 33294 27294 33346
rect 27346 33294 27360 33346
rect 27280 33280 27360 33294
rect 27440 33346 27520 33360
rect 27440 33294 27454 33346
rect 27506 33294 27520 33346
rect 27440 33280 27520 33294
rect 27600 33346 27680 33360
rect 27600 33294 27614 33346
rect 27666 33294 27680 33346
rect 27600 33280 27680 33294
rect 27760 33346 27840 33360
rect 27760 33294 27774 33346
rect 27826 33294 27840 33346
rect 27760 33280 27840 33294
rect 27920 33346 28000 33360
rect 27920 33294 27934 33346
rect 27986 33294 28000 33346
rect 27920 33280 28000 33294
rect 28080 33346 28160 33360
rect 28080 33294 28094 33346
rect 28146 33294 28160 33346
rect 28080 33280 28160 33294
rect 28240 33346 28320 33360
rect 28240 33294 28254 33346
rect 28306 33294 28320 33346
rect 28240 33280 28320 33294
rect 28400 33346 28480 33360
rect 28400 33294 28414 33346
rect 28466 33294 28480 33346
rect 28400 33280 28480 33294
rect 28560 33346 28640 33360
rect 28560 33294 28574 33346
rect 28626 33294 28640 33346
rect 28560 33280 28640 33294
rect 28720 33346 28800 33360
rect 28720 33294 28734 33346
rect 28786 33294 28800 33346
rect 28720 33280 28800 33294
rect 28880 33346 28960 33360
rect 28880 33294 28894 33346
rect 28946 33294 28960 33346
rect 28880 33280 28960 33294
rect 29040 33346 29120 33360
rect 29040 33294 29054 33346
rect 29106 33294 29120 33346
rect 29040 33280 29120 33294
rect 29200 33346 29280 33360
rect 29200 33294 29214 33346
rect 29266 33294 29280 33346
rect 29200 33280 29280 33294
rect 29360 33346 29440 33360
rect 29360 33294 29374 33346
rect 29426 33294 29440 33346
rect 29360 33280 29440 33294
rect 33520 33346 33600 33360
rect 33520 33294 33534 33346
rect 33586 33294 33600 33346
rect 33520 33280 33600 33294
rect 33680 33346 33760 33360
rect 33680 33294 33694 33346
rect 33746 33294 33760 33346
rect 33680 33280 33760 33294
rect 33840 33346 33920 33360
rect 33840 33294 33854 33346
rect 33906 33294 33920 33346
rect 33840 33280 33920 33294
rect 34000 33346 34080 33360
rect 34000 33294 34014 33346
rect 34066 33294 34080 33346
rect 34000 33280 34080 33294
rect 34160 33346 34240 33360
rect 34160 33294 34174 33346
rect 34226 33294 34240 33346
rect 34160 33280 34240 33294
rect 34320 33346 34400 33360
rect 34320 33294 34334 33346
rect 34386 33294 34400 33346
rect 34320 33280 34400 33294
rect 34480 33346 34560 33360
rect 34480 33294 34494 33346
rect 34546 33294 34560 33346
rect 34480 33280 34560 33294
rect 34640 33346 34720 33360
rect 34640 33294 34654 33346
rect 34706 33294 34720 33346
rect 34640 33280 34720 33294
rect 34800 33346 34880 33360
rect 34800 33294 34814 33346
rect 34866 33294 34880 33346
rect 34800 33280 34880 33294
rect 34960 33346 35040 33360
rect 34960 33294 34974 33346
rect 35026 33294 35040 33346
rect 34960 33280 35040 33294
rect 35120 33346 35200 33360
rect 35120 33294 35134 33346
rect 35186 33294 35200 33346
rect 35120 33280 35200 33294
rect 35280 33346 35360 33360
rect 35280 33294 35294 33346
rect 35346 33294 35360 33346
rect 35280 33280 35360 33294
rect 35440 33346 35520 33360
rect 35440 33294 35454 33346
rect 35506 33294 35520 33346
rect 35440 33280 35520 33294
rect 35600 33346 35680 33360
rect 35600 33294 35614 33346
rect 35666 33294 35680 33346
rect 35600 33280 35680 33294
rect 35760 33346 35840 33360
rect 35760 33294 35774 33346
rect 35826 33294 35840 33346
rect 35760 33280 35840 33294
rect 35920 33346 36000 33360
rect 35920 33294 35934 33346
rect 35986 33294 36000 33346
rect 35920 33280 36000 33294
rect 36080 33346 36160 33360
rect 36080 33294 36094 33346
rect 36146 33294 36160 33346
rect 36080 33280 36160 33294
rect 36240 33346 36320 33360
rect 36240 33294 36254 33346
rect 36306 33294 36320 33346
rect 36240 33280 36320 33294
rect 36400 33346 36480 33360
rect 36400 33294 36414 33346
rect 36466 33294 36480 33346
rect 36400 33280 36480 33294
rect 36560 33346 36640 33360
rect 36560 33294 36574 33346
rect 36626 33294 36640 33346
rect 36560 33280 36640 33294
rect 36720 33346 36800 33360
rect 36720 33294 36734 33346
rect 36786 33294 36800 33346
rect 36720 33280 36800 33294
rect 36880 33346 36960 33360
rect 36880 33294 36894 33346
rect 36946 33294 36960 33346
rect 36880 33280 36960 33294
rect 37040 33346 37120 33360
rect 37040 33294 37054 33346
rect 37106 33294 37120 33346
rect 37040 33280 37120 33294
rect 37200 33346 37280 33360
rect 37200 33294 37214 33346
rect 37266 33294 37280 33346
rect 37200 33280 37280 33294
rect 37360 33346 37440 33360
rect 37360 33294 37374 33346
rect 37426 33294 37440 33346
rect 37360 33280 37440 33294
rect 37520 33346 37600 33360
rect 37520 33294 37534 33346
rect 37586 33294 37600 33346
rect 37520 33280 37600 33294
rect 37680 33346 37760 33360
rect 37680 33294 37694 33346
rect 37746 33294 37760 33346
rect 37680 33280 37760 33294
rect 37840 33346 37920 33360
rect 37840 33294 37854 33346
rect 37906 33294 37920 33346
rect 37840 33280 37920 33294
rect 38000 33346 38080 33360
rect 38000 33294 38014 33346
rect 38066 33294 38080 33346
rect 38000 33280 38080 33294
rect 38160 33346 38240 33360
rect 38160 33294 38174 33346
rect 38226 33294 38240 33346
rect 38160 33280 38240 33294
rect 38320 33346 38400 33360
rect 38320 33294 38334 33346
rect 38386 33294 38400 33346
rect 38320 33280 38400 33294
rect 38480 33346 38560 33360
rect 38480 33294 38494 33346
rect 38546 33294 38560 33346
rect 38480 33280 38560 33294
rect 38640 33346 38720 33360
rect 38640 33294 38654 33346
rect 38706 33294 38720 33346
rect 38640 33280 38720 33294
rect 38800 33346 38880 33360
rect 38800 33294 38814 33346
rect 38866 33294 38880 33346
rect 38800 33280 38880 33294
rect 38960 33346 39040 33360
rect 38960 33294 38974 33346
rect 39026 33294 39040 33346
rect 38960 33280 39040 33294
rect 39120 33346 39200 33360
rect 39120 33294 39134 33346
rect 39186 33294 39200 33346
rect 39120 33280 39200 33294
rect 39280 33346 39360 33360
rect 39280 33294 39294 33346
rect 39346 33294 39360 33346
rect 39280 33280 39360 33294
rect 39440 33346 39520 33360
rect 39440 33294 39454 33346
rect 39506 33294 39520 33346
rect 39440 33280 39520 33294
rect 39600 33346 39680 33360
rect 39600 33294 39614 33346
rect 39666 33294 39680 33346
rect 39600 33280 39680 33294
rect 39760 33346 39840 33360
rect 39760 33294 39774 33346
rect 39826 33294 39840 33346
rect 39760 33280 39840 33294
rect 39920 33346 40000 33360
rect 39920 33294 39934 33346
rect 39986 33294 40000 33346
rect 39920 33280 40000 33294
rect 40080 33346 40160 33360
rect 40080 33294 40094 33346
rect 40146 33294 40160 33346
rect 40080 33280 40160 33294
rect 40240 33346 40320 33360
rect 40240 33294 40254 33346
rect 40306 33294 40320 33346
rect 40240 33280 40320 33294
rect 40400 33346 40480 33360
rect 40400 33294 40414 33346
rect 40466 33294 40480 33346
rect 40400 33280 40480 33294
rect 40560 33346 40640 33360
rect 40560 33294 40574 33346
rect 40626 33294 40640 33346
rect 40560 33280 40640 33294
rect 40720 33346 40800 33360
rect 40720 33294 40734 33346
rect 40786 33294 40800 33346
rect 40720 33280 40800 33294
rect 40880 33346 40960 33360
rect 40880 33294 40894 33346
rect 40946 33294 40960 33346
rect 40880 33280 40960 33294
rect 41040 33346 41120 33360
rect 41040 33294 41054 33346
rect 41106 33294 41120 33346
rect 41040 33280 41120 33294
rect 41200 33346 41280 33360
rect 41200 33294 41214 33346
rect 41266 33294 41280 33346
rect 41200 33280 41280 33294
rect 41360 33346 41440 33360
rect 41360 33294 41374 33346
rect 41426 33294 41440 33346
rect 41360 33280 41440 33294
rect 41520 33346 41600 33360
rect 41520 33294 41534 33346
rect 41586 33294 41600 33346
rect 41520 33280 41600 33294
rect 41680 33346 41760 33360
rect 41680 33294 41694 33346
rect 41746 33294 41760 33346
rect 41680 33280 41760 33294
rect 41840 33346 41920 33360
rect 41840 33294 41854 33346
rect 41906 33294 41920 33346
rect 41840 33280 41920 33294
rect 0 33026 80 33040
rect 0 32974 14 33026
rect 66 32974 80 33026
rect 0 32960 80 32974
rect 160 33026 240 33040
rect 160 32974 174 33026
rect 226 32974 240 33026
rect 160 32960 240 32974
rect 320 33026 400 33040
rect 320 32974 334 33026
rect 386 32974 400 33026
rect 320 32960 400 32974
rect 480 33026 560 33040
rect 480 32974 494 33026
rect 546 32974 560 33026
rect 480 32960 560 32974
rect 640 33026 720 33040
rect 640 32974 654 33026
rect 706 32974 720 33026
rect 640 32960 720 32974
rect 800 33026 880 33040
rect 800 32974 814 33026
rect 866 32974 880 33026
rect 800 32960 880 32974
rect 960 33026 1040 33040
rect 960 32974 974 33026
rect 1026 32974 1040 33026
rect 960 32960 1040 32974
rect 1120 33026 1200 33040
rect 1120 32974 1134 33026
rect 1186 32974 1200 33026
rect 1120 32960 1200 32974
rect 1280 33026 1360 33040
rect 1280 32974 1294 33026
rect 1346 32974 1360 33026
rect 1280 32960 1360 32974
rect 1440 33026 1520 33040
rect 1440 32974 1454 33026
rect 1506 32974 1520 33026
rect 1440 32960 1520 32974
rect 1600 33026 1680 33040
rect 1600 32974 1614 33026
rect 1666 32974 1680 33026
rect 1600 32960 1680 32974
rect 1760 33026 1840 33040
rect 1760 32974 1774 33026
rect 1826 32974 1840 33026
rect 1760 32960 1840 32974
rect 1920 33026 2000 33040
rect 1920 32974 1934 33026
rect 1986 32974 2000 33026
rect 1920 32960 2000 32974
rect 2080 33026 2160 33040
rect 2080 32974 2094 33026
rect 2146 32974 2160 33026
rect 2080 32960 2160 32974
rect 2240 33026 2320 33040
rect 2240 32974 2254 33026
rect 2306 32974 2320 33026
rect 2240 32960 2320 32974
rect 2400 33026 2480 33040
rect 2400 32974 2414 33026
rect 2466 32974 2480 33026
rect 2400 32960 2480 32974
rect 2560 33026 2640 33040
rect 2560 32974 2574 33026
rect 2626 32974 2640 33026
rect 2560 32960 2640 32974
rect 2720 33026 2800 33040
rect 2720 32974 2734 33026
rect 2786 32974 2800 33026
rect 2720 32960 2800 32974
rect 2880 33026 2960 33040
rect 2880 32974 2894 33026
rect 2946 32974 2960 33026
rect 2880 32960 2960 32974
rect 3040 33026 3120 33040
rect 3040 32974 3054 33026
rect 3106 32974 3120 33026
rect 3040 32960 3120 32974
rect 3200 33026 3280 33040
rect 3200 32974 3214 33026
rect 3266 32974 3280 33026
rect 3200 32960 3280 32974
rect 3360 33026 3440 33040
rect 3360 32974 3374 33026
rect 3426 32974 3440 33026
rect 3360 32960 3440 32974
rect 3520 33026 3600 33040
rect 3520 32974 3534 33026
rect 3586 32974 3600 33026
rect 3520 32960 3600 32974
rect 3680 33026 3760 33040
rect 3680 32974 3694 33026
rect 3746 32974 3760 33026
rect 3680 32960 3760 32974
rect 3840 33026 3920 33040
rect 3840 32974 3854 33026
rect 3906 32974 3920 33026
rect 3840 32960 3920 32974
rect 4000 33026 4080 33040
rect 4000 32974 4014 33026
rect 4066 32974 4080 33026
rect 4000 32960 4080 32974
rect 4160 33026 4240 33040
rect 4160 32974 4174 33026
rect 4226 32974 4240 33026
rect 4160 32960 4240 32974
rect 4320 33026 4400 33040
rect 4320 32974 4334 33026
rect 4386 32974 4400 33026
rect 4320 32960 4400 32974
rect 4480 33026 4560 33040
rect 4480 32974 4494 33026
rect 4546 32974 4560 33026
rect 4480 32960 4560 32974
rect 4640 33026 4720 33040
rect 4640 32974 4654 33026
rect 4706 32974 4720 33026
rect 4640 32960 4720 32974
rect 4800 33026 4880 33040
rect 4800 32974 4814 33026
rect 4866 32974 4880 33026
rect 4800 32960 4880 32974
rect 4960 33026 5040 33040
rect 4960 32974 4974 33026
rect 5026 32974 5040 33026
rect 4960 32960 5040 32974
rect 5120 33026 5200 33040
rect 5120 32974 5134 33026
rect 5186 32974 5200 33026
rect 5120 32960 5200 32974
rect 5280 33026 5360 33040
rect 5280 32974 5294 33026
rect 5346 32974 5360 33026
rect 5280 32960 5360 32974
rect 5440 33026 5520 33040
rect 5440 32974 5454 33026
rect 5506 32974 5520 33026
rect 5440 32960 5520 32974
rect 5600 33026 5680 33040
rect 5600 32974 5614 33026
rect 5666 32974 5680 33026
rect 5600 32960 5680 32974
rect 5760 33026 5840 33040
rect 5760 32974 5774 33026
rect 5826 32974 5840 33026
rect 5760 32960 5840 32974
rect 5920 33026 6000 33040
rect 5920 32974 5934 33026
rect 5986 32974 6000 33026
rect 5920 32960 6000 32974
rect 6080 33026 6160 33040
rect 6080 32974 6094 33026
rect 6146 32974 6160 33026
rect 6080 32960 6160 32974
rect 6240 33026 6320 33040
rect 6240 32974 6254 33026
rect 6306 32974 6320 33026
rect 6240 32960 6320 32974
rect 6400 33026 6480 33040
rect 6400 32974 6414 33026
rect 6466 32974 6480 33026
rect 6400 32960 6480 32974
rect 6560 33026 6640 33040
rect 6560 32974 6574 33026
rect 6626 32974 6640 33026
rect 6560 32960 6640 32974
rect 6720 33026 6800 33040
rect 6720 32974 6734 33026
rect 6786 32974 6800 33026
rect 6720 32960 6800 32974
rect 6880 33026 6960 33040
rect 6880 32974 6894 33026
rect 6946 32974 6960 33026
rect 6880 32960 6960 32974
rect 7040 33026 7120 33040
rect 7040 32974 7054 33026
rect 7106 32974 7120 33026
rect 7040 32960 7120 32974
rect 7200 33026 7280 33040
rect 7200 32974 7214 33026
rect 7266 32974 7280 33026
rect 7200 32960 7280 32974
rect 7360 33026 7440 33040
rect 7360 32974 7374 33026
rect 7426 32974 7440 33026
rect 7360 32960 7440 32974
rect 7520 33026 7600 33040
rect 7520 32974 7534 33026
rect 7586 32974 7600 33026
rect 7520 32960 7600 32974
rect 7680 33026 7760 33040
rect 7680 32974 7694 33026
rect 7746 32974 7760 33026
rect 7680 32960 7760 32974
rect 7840 33026 7920 33040
rect 7840 32974 7854 33026
rect 7906 32974 7920 33026
rect 7840 32960 7920 32974
rect 8000 33026 8080 33040
rect 8000 32974 8014 33026
rect 8066 32974 8080 33026
rect 8000 32960 8080 32974
rect 8160 33026 8240 33040
rect 8160 32974 8174 33026
rect 8226 32974 8240 33026
rect 8160 32960 8240 32974
rect 8320 33026 8400 33040
rect 8320 32974 8334 33026
rect 8386 32974 8400 33026
rect 8320 32960 8400 32974
rect 12480 33026 12560 33040
rect 12480 32974 12494 33026
rect 12546 32974 12560 33026
rect 12480 32960 12560 32974
rect 12640 33026 12720 33040
rect 12640 32974 12654 33026
rect 12706 32974 12720 33026
rect 12640 32960 12720 32974
rect 12800 33026 12880 33040
rect 12800 32974 12814 33026
rect 12866 32974 12880 33026
rect 12800 32960 12880 32974
rect 12960 33026 13040 33040
rect 12960 32974 12974 33026
rect 13026 32974 13040 33026
rect 12960 32960 13040 32974
rect 13120 33026 13200 33040
rect 13120 32974 13134 33026
rect 13186 32974 13200 33026
rect 13120 32960 13200 32974
rect 13280 33026 13360 33040
rect 13280 32974 13294 33026
rect 13346 32974 13360 33026
rect 13280 32960 13360 32974
rect 13440 33026 13520 33040
rect 13440 32974 13454 33026
rect 13506 32974 13520 33026
rect 13440 32960 13520 32974
rect 13600 33026 13680 33040
rect 13600 32974 13614 33026
rect 13666 32974 13680 33026
rect 13600 32960 13680 32974
rect 13760 33026 13840 33040
rect 13760 32974 13774 33026
rect 13826 32974 13840 33026
rect 13760 32960 13840 32974
rect 13920 33026 14000 33040
rect 13920 32974 13934 33026
rect 13986 32974 14000 33026
rect 13920 32960 14000 32974
rect 14080 33026 14160 33040
rect 14080 32974 14094 33026
rect 14146 32974 14160 33026
rect 14080 32960 14160 32974
rect 14240 33026 14320 33040
rect 14240 32974 14254 33026
rect 14306 32974 14320 33026
rect 14240 32960 14320 32974
rect 14400 33026 14480 33040
rect 14400 32974 14414 33026
rect 14466 32974 14480 33026
rect 14400 32960 14480 32974
rect 14560 33026 14640 33040
rect 14560 32974 14574 33026
rect 14626 32974 14640 33026
rect 14560 32960 14640 32974
rect 14720 33026 14800 33040
rect 14720 32974 14734 33026
rect 14786 32974 14800 33026
rect 14720 32960 14800 32974
rect 14880 33026 14960 33040
rect 14880 32974 14894 33026
rect 14946 32974 14960 33026
rect 14880 32960 14960 32974
rect 15040 33026 15120 33040
rect 15040 32974 15054 33026
rect 15106 32974 15120 33026
rect 15040 32960 15120 32974
rect 15200 33026 15280 33040
rect 15200 32974 15214 33026
rect 15266 32974 15280 33026
rect 15200 32960 15280 32974
rect 15360 33026 15440 33040
rect 15360 32974 15374 33026
rect 15426 32974 15440 33026
rect 15360 32960 15440 32974
rect 15520 33026 15600 33040
rect 15520 32974 15534 33026
rect 15586 32974 15600 33026
rect 15520 32960 15600 32974
rect 15680 33026 15760 33040
rect 15680 32974 15694 33026
rect 15746 32974 15760 33026
rect 15680 32960 15760 32974
rect 15840 33026 15920 33040
rect 15840 32974 15854 33026
rect 15906 32974 15920 33026
rect 15840 32960 15920 32974
rect 16000 33026 16080 33040
rect 16000 32974 16014 33026
rect 16066 32974 16080 33026
rect 16000 32960 16080 32974
rect 16160 33026 16240 33040
rect 16160 32974 16174 33026
rect 16226 32974 16240 33026
rect 16160 32960 16240 32974
rect 16320 33026 16400 33040
rect 16320 32974 16334 33026
rect 16386 32974 16400 33026
rect 16320 32960 16400 32974
rect 16480 33026 16560 33040
rect 16480 32974 16494 33026
rect 16546 32974 16560 33026
rect 16480 32960 16560 32974
rect 16640 33026 16720 33040
rect 16640 32974 16654 33026
rect 16706 32974 16720 33026
rect 16640 32960 16720 32974
rect 16800 33026 16880 33040
rect 16800 32974 16814 33026
rect 16866 32974 16880 33026
rect 16800 32960 16880 32974
rect 16960 33026 17040 33040
rect 16960 32974 16974 33026
rect 17026 32974 17040 33026
rect 16960 32960 17040 32974
rect 17120 33026 17200 33040
rect 17120 32974 17134 33026
rect 17186 32974 17200 33026
rect 17120 32960 17200 32974
rect 17280 33026 17360 33040
rect 17280 32974 17294 33026
rect 17346 32974 17360 33026
rect 17280 32960 17360 32974
rect 17440 33026 17520 33040
rect 17440 32974 17454 33026
rect 17506 32974 17520 33026
rect 17440 32960 17520 32974
rect 17600 33026 17680 33040
rect 17600 32974 17614 33026
rect 17666 32974 17680 33026
rect 17600 32960 17680 32974
rect 17760 33026 17840 33040
rect 17760 32974 17774 33026
rect 17826 32974 17840 33026
rect 17760 32960 17840 32974
rect 17920 33026 18000 33040
rect 17920 32974 17934 33026
rect 17986 32974 18000 33026
rect 17920 32960 18000 32974
rect 18080 33026 18160 33040
rect 18080 32974 18094 33026
rect 18146 32974 18160 33026
rect 18080 32960 18160 32974
rect 18240 33026 18320 33040
rect 18240 32974 18254 33026
rect 18306 32974 18320 33026
rect 18240 32960 18320 32974
rect 18400 33026 18480 33040
rect 18400 32974 18414 33026
rect 18466 32974 18480 33026
rect 18400 32960 18480 32974
rect 18560 33026 18640 33040
rect 18560 32974 18574 33026
rect 18626 32974 18640 33026
rect 18560 32960 18640 32974
rect 18720 33026 18800 33040
rect 18720 32974 18734 33026
rect 18786 32974 18800 33026
rect 18720 32960 18800 32974
rect 18880 33026 18960 33040
rect 18880 32974 18894 33026
rect 18946 32974 18960 33026
rect 18880 32960 18960 32974
rect 23120 33026 23200 33040
rect 23120 32974 23134 33026
rect 23186 32974 23200 33026
rect 23120 32960 23200 32974
rect 23280 33026 23360 33040
rect 23280 32974 23294 33026
rect 23346 32974 23360 33026
rect 23280 32960 23360 32974
rect 23440 33026 23520 33040
rect 23440 32974 23454 33026
rect 23506 32974 23520 33026
rect 23440 32960 23520 32974
rect 23600 33026 23680 33040
rect 23600 32974 23614 33026
rect 23666 32974 23680 33026
rect 23600 32960 23680 32974
rect 23760 33026 23840 33040
rect 23760 32974 23774 33026
rect 23826 32974 23840 33026
rect 23760 32960 23840 32974
rect 23920 33026 24000 33040
rect 23920 32974 23934 33026
rect 23986 32974 24000 33026
rect 23920 32960 24000 32974
rect 24080 33026 24160 33040
rect 24080 32974 24094 33026
rect 24146 32974 24160 33026
rect 24080 32960 24160 32974
rect 24240 33026 24320 33040
rect 24240 32974 24254 33026
rect 24306 32974 24320 33026
rect 24240 32960 24320 32974
rect 24400 33026 24480 33040
rect 24400 32974 24414 33026
rect 24466 32974 24480 33026
rect 24400 32960 24480 32974
rect 24560 33026 24640 33040
rect 24560 32974 24574 33026
rect 24626 32974 24640 33026
rect 24560 32960 24640 32974
rect 24720 33026 24800 33040
rect 24720 32974 24734 33026
rect 24786 32974 24800 33026
rect 24720 32960 24800 32974
rect 24880 33026 24960 33040
rect 24880 32974 24894 33026
rect 24946 32974 24960 33026
rect 24880 32960 24960 32974
rect 25040 33026 25120 33040
rect 25040 32974 25054 33026
rect 25106 32974 25120 33026
rect 25040 32960 25120 32974
rect 25200 33026 25280 33040
rect 25200 32974 25214 33026
rect 25266 32974 25280 33026
rect 25200 32960 25280 32974
rect 25360 33026 25440 33040
rect 25360 32974 25374 33026
rect 25426 32974 25440 33026
rect 25360 32960 25440 32974
rect 25520 33026 25600 33040
rect 25520 32974 25534 33026
rect 25586 32974 25600 33026
rect 25520 32960 25600 32974
rect 25680 33026 25760 33040
rect 25680 32974 25694 33026
rect 25746 32974 25760 33026
rect 25680 32960 25760 32974
rect 25840 33026 25920 33040
rect 25840 32974 25854 33026
rect 25906 32974 25920 33026
rect 25840 32960 25920 32974
rect 26000 33026 26080 33040
rect 26000 32974 26014 33026
rect 26066 32974 26080 33026
rect 26000 32960 26080 32974
rect 26160 33026 26240 33040
rect 26160 32974 26174 33026
rect 26226 32974 26240 33026
rect 26160 32960 26240 32974
rect 26320 33026 26400 33040
rect 26320 32974 26334 33026
rect 26386 32974 26400 33026
rect 26320 32960 26400 32974
rect 26480 33026 26560 33040
rect 26480 32974 26494 33026
rect 26546 32974 26560 33026
rect 26480 32960 26560 32974
rect 26640 33026 26720 33040
rect 26640 32974 26654 33026
rect 26706 32974 26720 33026
rect 26640 32960 26720 32974
rect 26800 33026 26880 33040
rect 26800 32974 26814 33026
rect 26866 32974 26880 33026
rect 26800 32960 26880 32974
rect 26960 33026 27040 33040
rect 26960 32974 26974 33026
rect 27026 32974 27040 33026
rect 26960 32960 27040 32974
rect 27120 33026 27200 33040
rect 27120 32974 27134 33026
rect 27186 32974 27200 33026
rect 27120 32960 27200 32974
rect 27280 33026 27360 33040
rect 27280 32974 27294 33026
rect 27346 32974 27360 33026
rect 27280 32960 27360 32974
rect 27440 33026 27520 33040
rect 27440 32974 27454 33026
rect 27506 32974 27520 33026
rect 27440 32960 27520 32974
rect 27600 33026 27680 33040
rect 27600 32974 27614 33026
rect 27666 32974 27680 33026
rect 27600 32960 27680 32974
rect 27760 33026 27840 33040
rect 27760 32974 27774 33026
rect 27826 32974 27840 33026
rect 27760 32960 27840 32974
rect 27920 33026 28000 33040
rect 27920 32974 27934 33026
rect 27986 32974 28000 33026
rect 27920 32960 28000 32974
rect 28080 33026 28160 33040
rect 28080 32974 28094 33026
rect 28146 32974 28160 33026
rect 28080 32960 28160 32974
rect 28240 33026 28320 33040
rect 28240 32974 28254 33026
rect 28306 32974 28320 33026
rect 28240 32960 28320 32974
rect 28400 33026 28480 33040
rect 28400 32974 28414 33026
rect 28466 32974 28480 33026
rect 28400 32960 28480 32974
rect 28560 33026 28640 33040
rect 28560 32974 28574 33026
rect 28626 32974 28640 33026
rect 28560 32960 28640 32974
rect 28720 33026 28800 33040
rect 28720 32974 28734 33026
rect 28786 32974 28800 33026
rect 28720 32960 28800 32974
rect 28880 33026 28960 33040
rect 28880 32974 28894 33026
rect 28946 32974 28960 33026
rect 28880 32960 28960 32974
rect 29040 33026 29120 33040
rect 29040 32974 29054 33026
rect 29106 32974 29120 33026
rect 29040 32960 29120 32974
rect 29200 33026 29280 33040
rect 29200 32974 29214 33026
rect 29266 32974 29280 33026
rect 29200 32960 29280 32974
rect 29360 33026 29440 33040
rect 29360 32974 29374 33026
rect 29426 32974 29440 33026
rect 29360 32960 29440 32974
rect 33520 33026 33600 33040
rect 33520 32974 33534 33026
rect 33586 32974 33600 33026
rect 33520 32960 33600 32974
rect 33680 33026 33760 33040
rect 33680 32974 33694 33026
rect 33746 32974 33760 33026
rect 33680 32960 33760 32974
rect 33840 33026 33920 33040
rect 33840 32974 33854 33026
rect 33906 32974 33920 33026
rect 33840 32960 33920 32974
rect 34000 33026 34080 33040
rect 34000 32974 34014 33026
rect 34066 32974 34080 33026
rect 34000 32960 34080 32974
rect 34160 33026 34240 33040
rect 34160 32974 34174 33026
rect 34226 32974 34240 33026
rect 34160 32960 34240 32974
rect 34320 33026 34400 33040
rect 34320 32974 34334 33026
rect 34386 32974 34400 33026
rect 34320 32960 34400 32974
rect 34480 33026 34560 33040
rect 34480 32974 34494 33026
rect 34546 32974 34560 33026
rect 34480 32960 34560 32974
rect 34640 33026 34720 33040
rect 34640 32974 34654 33026
rect 34706 32974 34720 33026
rect 34640 32960 34720 32974
rect 34800 33026 34880 33040
rect 34800 32974 34814 33026
rect 34866 32974 34880 33026
rect 34800 32960 34880 32974
rect 34960 33026 35040 33040
rect 34960 32974 34974 33026
rect 35026 32974 35040 33026
rect 34960 32960 35040 32974
rect 35120 33026 35200 33040
rect 35120 32974 35134 33026
rect 35186 32974 35200 33026
rect 35120 32960 35200 32974
rect 35280 33026 35360 33040
rect 35280 32974 35294 33026
rect 35346 32974 35360 33026
rect 35280 32960 35360 32974
rect 35440 33026 35520 33040
rect 35440 32974 35454 33026
rect 35506 32974 35520 33026
rect 35440 32960 35520 32974
rect 35600 33026 35680 33040
rect 35600 32974 35614 33026
rect 35666 32974 35680 33026
rect 35600 32960 35680 32974
rect 35760 33026 35840 33040
rect 35760 32974 35774 33026
rect 35826 32974 35840 33026
rect 35760 32960 35840 32974
rect 35920 33026 36000 33040
rect 35920 32974 35934 33026
rect 35986 32974 36000 33026
rect 35920 32960 36000 32974
rect 36080 33026 36160 33040
rect 36080 32974 36094 33026
rect 36146 32974 36160 33026
rect 36080 32960 36160 32974
rect 36240 33026 36320 33040
rect 36240 32974 36254 33026
rect 36306 32974 36320 33026
rect 36240 32960 36320 32974
rect 36400 33026 36480 33040
rect 36400 32974 36414 33026
rect 36466 32974 36480 33026
rect 36400 32960 36480 32974
rect 36560 33026 36640 33040
rect 36560 32974 36574 33026
rect 36626 32974 36640 33026
rect 36560 32960 36640 32974
rect 36720 33026 36800 33040
rect 36720 32974 36734 33026
rect 36786 32974 36800 33026
rect 36720 32960 36800 32974
rect 36880 33026 36960 33040
rect 36880 32974 36894 33026
rect 36946 32974 36960 33026
rect 36880 32960 36960 32974
rect 37040 33026 37120 33040
rect 37040 32974 37054 33026
rect 37106 32974 37120 33026
rect 37040 32960 37120 32974
rect 37200 33026 37280 33040
rect 37200 32974 37214 33026
rect 37266 32974 37280 33026
rect 37200 32960 37280 32974
rect 37360 33026 37440 33040
rect 37360 32974 37374 33026
rect 37426 32974 37440 33026
rect 37360 32960 37440 32974
rect 37520 33026 37600 33040
rect 37520 32974 37534 33026
rect 37586 32974 37600 33026
rect 37520 32960 37600 32974
rect 37680 33026 37760 33040
rect 37680 32974 37694 33026
rect 37746 32974 37760 33026
rect 37680 32960 37760 32974
rect 37840 33026 37920 33040
rect 37840 32974 37854 33026
rect 37906 32974 37920 33026
rect 37840 32960 37920 32974
rect 38000 33026 38080 33040
rect 38000 32974 38014 33026
rect 38066 32974 38080 33026
rect 38000 32960 38080 32974
rect 38160 33026 38240 33040
rect 38160 32974 38174 33026
rect 38226 32974 38240 33026
rect 38160 32960 38240 32974
rect 38320 33026 38400 33040
rect 38320 32974 38334 33026
rect 38386 32974 38400 33026
rect 38320 32960 38400 32974
rect 38480 33026 38560 33040
rect 38480 32974 38494 33026
rect 38546 32974 38560 33026
rect 38480 32960 38560 32974
rect 38640 33026 38720 33040
rect 38640 32974 38654 33026
rect 38706 32974 38720 33026
rect 38640 32960 38720 32974
rect 38800 33026 38880 33040
rect 38800 32974 38814 33026
rect 38866 32974 38880 33026
rect 38800 32960 38880 32974
rect 38960 33026 39040 33040
rect 38960 32974 38974 33026
rect 39026 32974 39040 33026
rect 38960 32960 39040 32974
rect 39120 33026 39200 33040
rect 39120 32974 39134 33026
rect 39186 32974 39200 33026
rect 39120 32960 39200 32974
rect 39280 33026 39360 33040
rect 39280 32974 39294 33026
rect 39346 32974 39360 33026
rect 39280 32960 39360 32974
rect 39440 33026 39520 33040
rect 39440 32974 39454 33026
rect 39506 32974 39520 33026
rect 39440 32960 39520 32974
rect 39600 33026 39680 33040
rect 39600 32974 39614 33026
rect 39666 32974 39680 33026
rect 39600 32960 39680 32974
rect 39760 33026 39840 33040
rect 39760 32974 39774 33026
rect 39826 32974 39840 33026
rect 39760 32960 39840 32974
rect 39920 33026 40000 33040
rect 39920 32974 39934 33026
rect 39986 32974 40000 33026
rect 39920 32960 40000 32974
rect 40080 33026 40160 33040
rect 40080 32974 40094 33026
rect 40146 32974 40160 33026
rect 40080 32960 40160 32974
rect 40240 33026 40320 33040
rect 40240 32974 40254 33026
rect 40306 32974 40320 33026
rect 40240 32960 40320 32974
rect 40400 33026 40480 33040
rect 40400 32974 40414 33026
rect 40466 32974 40480 33026
rect 40400 32960 40480 32974
rect 40560 33026 40640 33040
rect 40560 32974 40574 33026
rect 40626 32974 40640 33026
rect 40560 32960 40640 32974
rect 40720 33026 40800 33040
rect 40720 32974 40734 33026
rect 40786 32974 40800 33026
rect 40720 32960 40800 32974
rect 40880 33026 40960 33040
rect 40880 32974 40894 33026
rect 40946 32974 40960 33026
rect 40880 32960 40960 32974
rect 41040 33026 41120 33040
rect 41040 32974 41054 33026
rect 41106 32974 41120 33026
rect 41040 32960 41120 32974
rect 41200 33026 41280 33040
rect 41200 32974 41214 33026
rect 41266 32974 41280 33026
rect 41200 32960 41280 32974
rect 41360 33026 41440 33040
rect 41360 32974 41374 33026
rect 41426 32974 41440 33026
rect 41360 32960 41440 32974
rect 41520 33026 41600 33040
rect 41520 32974 41534 33026
rect 41586 32974 41600 33026
rect 41520 32960 41600 32974
rect 41680 33026 41760 33040
rect 41680 32974 41694 33026
rect 41746 32974 41760 33026
rect 41680 32960 41760 32974
rect 41840 33026 41920 33040
rect 41840 32974 41854 33026
rect 41906 32974 41920 33026
rect 41840 32960 41920 32974
rect 0 32866 80 32880
rect 0 32814 14 32866
rect 66 32814 80 32866
rect 0 32800 80 32814
rect 160 32866 240 32880
rect 160 32814 174 32866
rect 226 32814 240 32866
rect 160 32800 240 32814
rect 320 32866 400 32880
rect 320 32814 334 32866
rect 386 32814 400 32866
rect 320 32800 400 32814
rect 480 32866 560 32880
rect 480 32814 494 32866
rect 546 32814 560 32866
rect 480 32800 560 32814
rect 640 32866 720 32880
rect 640 32814 654 32866
rect 706 32814 720 32866
rect 640 32800 720 32814
rect 800 32866 880 32880
rect 800 32814 814 32866
rect 866 32814 880 32866
rect 800 32800 880 32814
rect 960 32866 1040 32880
rect 960 32814 974 32866
rect 1026 32814 1040 32866
rect 960 32800 1040 32814
rect 1120 32866 1200 32880
rect 1120 32814 1134 32866
rect 1186 32814 1200 32866
rect 1120 32800 1200 32814
rect 1280 32866 1360 32880
rect 1280 32814 1294 32866
rect 1346 32814 1360 32866
rect 1280 32800 1360 32814
rect 1440 32866 1520 32880
rect 1440 32814 1454 32866
rect 1506 32814 1520 32866
rect 1440 32800 1520 32814
rect 1600 32866 1680 32880
rect 1600 32814 1614 32866
rect 1666 32814 1680 32866
rect 1600 32800 1680 32814
rect 1760 32866 1840 32880
rect 1760 32814 1774 32866
rect 1826 32814 1840 32866
rect 1760 32800 1840 32814
rect 1920 32866 2000 32880
rect 1920 32814 1934 32866
rect 1986 32814 2000 32866
rect 1920 32800 2000 32814
rect 2080 32866 2160 32880
rect 2080 32814 2094 32866
rect 2146 32814 2160 32866
rect 2080 32800 2160 32814
rect 2240 32866 2320 32880
rect 2240 32814 2254 32866
rect 2306 32814 2320 32866
rect 2240 32800 2320 32814
rect 2400 32866 2480 32880
rect 2400 32814 2414 32866
rect 2466 32814 2480 32866
rect 2400 32800 2480 32814
rect 2560 32866 2640 32880
rect 2560 32814 2574 32866
rect 2626 32814 2640 32866
rect 2560 32800 2640 32814
rect 2720 32866 2800 32880
rect 2720 32814 2734 32866
rect 2786 32814 2800 32866
rect 2720 32800 2800 32814
rect 2880 32866 2960 32880
rect 2880 32814 2894 32866
rect 2946 32814 2960 32866
rect 2880 32800 2960 32814
rect 3040 32866 3120 32880
rect 3040 32814 3054 32866
rect 3106 32814 3120 32866
rect 3040 32800 3120 32814
rect 3200 32866 3280 32880
rect 3200 32814 3214 32866
rect 3266 32814 3280 32866
rect 3200 32800 3280 32814
rect 3360 32866 3440 32880
rect 3360 32814 3374 32866
rect 3426 32814 3440 32866
rect 3360 32800 3440 32814
rect 3520 32866 3600 32880
rect 3520 32814 3534 32866
rect 3586 32814 3600 32866
rect 3520 32800 3600 32814
rect 3680 32866 3760 32880
rect 3680 32814 3694 32866
rect 3746 32814 3760 32866
rect 3680 32800 3760 32814
rect 3840 32866 3920 32880
rect 3840 32814 3854 32866
rect 3906 32814 3920 32866
rect 3840 32800 3920 32814
rect 4000 32866 4080 32880
rect 4000 32814 4014 32866
rect 4066 32814 4080 32866
rect 4000 32800 4080 32814
rect 4160 32866 4240 32880
rect 4160 32814 4174 32866
rect 4226 32814 4240 32866
rect 4160 32800 4240 32814
rect 4320 32866 4400 32880
rect 4320 32814 4334 32866
rect 4386 32814 4400 32866
rect 4320 32800 4400 32814
rect 4480 32866 4560 32880
rect 4480 32814 4494 32866
rect 4546 32814 4560 32866
rect 4480 32800 4560 32814
rect 4640 32866 4720 32880
rect 4640 32814 4654 32866
rect 4706 32814 4720 32866
rect 4640 32800 4720 32814
rect 4800 32866 4880 32880
rect 4800 32814 4814 32866
rect 4866 32814 4880 32866
rect 4800 32800 4880 32814
rect 4960 32866 5040 32880
rect 4960 32814 4974 32866
rect 5026 32814 5040 32866
rect 4960 32800 5040 32814
rect 5120 32866 5200 32880
rect 5120 32814 5134 32866
rect 5186 32814 5200 32866
rect 5120 32800 5200 32814
rect 5280 32866 5360 32880
rect 5280 32814 5294 32866
rect 5346 32814 5360 32866
rect 5280 32800 5360 32814
rect 5440 32866 5520 32880
rect 5440 32814 5454 32866
rect 5506 32814 5520 32866
rect 5440 32800 5520 32814
rect 5600 32866 5680 32880
rect 5600 32814 5614 32866
rect 5666 32814 5680 32866
rect 5600 32800 5680 32814
rect 5760 32866 5840 32880
rect 5760 32814 5774 32866
rect 5826 32814 5840 32866
rect 5760 32800 5840 32814
rect 5920 32866 6000 32880
rect 5920 32814 5934 32866
rect 5986 32814 6000 32866
rect 5920 32800 6000 32814
rect 6080 32866 6160 32880
rect 6080 32814 6094 32866
rect 6146 32814 6160 32866
rect 6080 32800 6160 32814
rect 6240 32866 6320 32880
rect 6240 32814 6254 32866
rect 6306 32814 6320 32866
rect 6240 32800 6320 32814
rect 6400 32866 6480 32880
rect 6400 32814 6414 32866
rect 6466 32814 6480 32866
rect 6400 32800 6480 32814
rect 6560 32866 6640 32880
rect 6560 32814 6574 32866
rect 6626 32814 6640 32866
rect 6560 32800 6640 32814
rect 6720 32866 6800 32880
rect 6720 32814 6734 32866
rect 6786 32814 6800 32866
rect 6720 32800 6800 32814
rect 6880 32866 6960 32880
rect 6880 32814 6894 32866
rect 6946 32814 6960 32866
rect 6880 32800 6960 32814
rect 7040 32866 7120 32880
rect 7040 32814 7054 32866
rect 7106 32814 7120 32866
rect 7040 32800 7120 32814
rect 7200 32866 7280 32880
rect 7200 32814 7214 32866
rect 7266 32814 7280 32866
rect 7200 32800 7280 32814
rect 7360 32866 7440 32880
rect 7360 32814 7374 32866
rect 7426 32814 7440 32866
rect 7360 32800 7440 32814
rect 7520 32866 7600 32880
rect 7520 32814 7534 32866
rect 7586 32814 7600 32866
rect 7520 32800 7600 32814
rect 7680 32866 7760 32880
rect 7680 32814 7694 32866
rect 7746 32814 7760 32866
rect 7680 32800 7760 32814
rect 7840 32866 7920 32880
rect 7840 32814 7854 32866
rect 7906 32814 7920 32866
rect 7840 32800 7920 32814
rect 8000 32866 8080 32880
rect 8000 32814 8014 32866
rect 8066 32814 8080 32866
rect 8000 32800 8080 32814
rect 8160 32866 8240 32880
rect 8160 32814 8174 32866
rect 8226 32814 8240 32866
rect 8160 32800 8240 32814
rect 8320 32866 8400 32880
rect 8320 32814 8334 32866
rect 8386 32814 8400 32866
rect 8320 32800 8400 32814
rect 12480 32866 12560 32880
rect 12480 32814 12494 32866
rect 12546 32814 12560 32866
rect 12480 32800 12560 32814
rect 12640 32866 12720 32880
rect 12640 32814 12654 32866
rect 12706 32814 12720 32866
rect 12640 32800 12720 32814
rect 12800 32866 12880 32880
rect 12800 32814 12814 32866
rect 12866 32814 12880 32866
rect 12800 32800 12880 32814
rect 12960 32866 13040 32880
rect 12960 32814 12974 32866
rect 13026 32814 13040 32866
rect 12960 32800 13040 32814
rect 13120 32866 13200 32880
rect 13120 32814 13134 32866
rect 13186 32814 13200 32866
rect 13120 32800 13200 32814
rect 13280 32866 13360 32880
rect 13280 32814 13294 32866
rect 13346 32814 13360 32866
rect 13280 32800 13360 32814
rect 13440 32866 13520 32880
rect 13440 32814 13454 32866
rect 13506 32814 13520 32866
rect 13440 32800 13520 32814
rect 13600 32866 13680 32880
rect 13600 32814 13614 32866
rect 13666 32814 13680 32866
rect 13600 32800 13680 32814
rect 13760 32866 13840 32880
rect 13760 32814 13774 32866
rect 13826 32814 13840 32866
rect 13760 32800 13840 32814
rect 13920 32866 14000 32880
rect 13920 32814 13934 32866
rect 13986 32814 14000 32866
rect 13920 32800 14000 32814
rect 14080 32866 14160 32880
rect 14080 32814 14094 32866
rect 14146 32814 14160 32866
rect 14080 32800 14160 32814
rect 14240 32866 14320 32880
rect 14240 32814 14254 32866
rect 14306 32814 14320 32866
rect 14240 32800 14320 32814
rect 14400 32866 14480 32880
rect 14400 32814 14414 32866
rect 14466 32814 14480 32866
rect 14400 32800 14480 32814
rect 14560 32866 14640 32880
rect 14560 32814 14574 32866
rect 14626 32814 14640 32866
rect 14560 32800 14640 32814
rect 14720 32866 14800 32880
rect 14720 32814 14734 32866
rect 14786 32814 14800 32866
rect 14720 32800 14800 32814
rect 14880 32866 14960 32880
rect 14880 32814 14894 32866
rect 14946 32814 14960 32866
rect 14880 32800 14960 32814
rect 15040 32866 15120 32880
rect 15040 32814 15054 32866
rect 15106 32814 15120 32866
rect 15040 32800 15120 32814
rect 15200 32866 15280 32880
rect 15200 32814 15214 32866
rect 15266 32814 15280 32866
rect 15200 32800 15280 32814
rect 15360 32866 15440 32880
rect 15360 32814 15374 32866
rect 15426 32814 15440 32866
rect 15360 32800 15440 32814
rect 15520 32866 15600 32880
rect 15520 32814 15534 32866
rect 15586 32814 15600 32866
rect 15520 32800 15600 32814
rect 15680 32866 15760 32880
rect 15680 32814 15694 32866
rect 15746 32814 15760 32866
rect 15680 32800 15760 32814
rect 15840 32866 15920 32880
rect 15840 32814 15854 32866
rect 15906 32814 15920 32866
rect 15840 32800 15920 32814
rect 16000 32866 16080 32880
rect 16000 32814 16014 32866
rect 16066 32814 16080 32866
rect 16000 32800 16080 32814
rect 16160 32866 16240 32880
rect 16160 32814 16174 32866
rect 16226 32814 16240 32866
rect 16160 32800 16240 32814
rect 16320 32866 16400 32880
rect 16320 32814 16334 32866
rect 16386 32814 16400 32866
rect 16320 32800 16400 32814
rect 16480 32866 16560 32880
rect 16480 32814 16494 32866
rect 16546 32814 16560 32866
rect 16480 32800 16560 32814
rect 16640 32866 16720 32880
rect 16640 32814 16654 32866
rect 16706 32814 16720 32866
rect 16640 32800 16720 32814
rect 16800 32866 16880 32880
rect 16800 32814 16814 32866
rect 16866 32814 16880 32866
rect 16800 32800 16880 32814
rect 16960 32866 17040 32880
rect 16960 32814 16974 32866
rect 17026 32814 17040 32866
rect 16960 32800 17040 32814
rect 17120 32866 17200 32880
rect 17120 32814 17134 32866
rect 17186 32814 17200 32866
rect 17120 32800 17200 32814
rect 17280 32866 17360 32880
rect 17280 32814 17294 32866
rect 17346 32814 17360 32866
rect 17280 32800 17360 32814
rect 17440 32866 17520 32880
rect 17440 32814 17454 32866
rect 17506 32814 17520 32866
rect 17440 32800 17520 32814
rect 17600 32866 17680 32880
rect 17600 32814 17614 32866
rect 17666 32814 17680 32866
rect 17600 32800 17680 32814
rect 17760 32866 17840 32880
rect 17760 32814 17774 32866
rect 17826 32814 17840 32866
rect 17760 32800 17840 32814
rect 17920 32866 18000 32880
rect 17920 32814 17934 32866
rect 17986 32814 18000 32866
rect 17920 32800 18000 32814
rect 18080 32866 18160 32880
rect 18080 32814 18094 32866
rect 18146 32814 18160 32866
rect 18080 32800 18160 32814
rect 18240 32866 18320 32880
rect 18240 32814 18254 32866
rect 18306 32814 18320 32866
rect 18240 32800 18320 32814
rect 18400 32866 18480 32880
rect 18400 32814 18414 32866
rect 18466 32814 18480 32866
rect 18400 32800 18480 32814
rect 18560 32866 18640 32880
rect 18560 32814 18574 32866
rect 18626 32814 18640 32866
rect 18560 32800 18640 32814
rect 18720 32866 18800 32880
rect 18720 32814 18734 32866
rect 18786 32814 18800 32866
rect 18720 32800 18800 32814
rect 18880 32866 18960 32880
rect 18880 32814 18894 32866
rect 18946 32814 18960 32866
rect 18880 32800 18960 32814
rect 23120 32866 23200 32880
rect 23120 32814 23134 32866
rect 23186 32814 23200 32866
rect 23120 32800 23200 32814
rect 23280 32866 23360 32880
rect 23280 32814 23294 32866
rect 23346 32814 23360 32866
rect 23280 32800 23360 32814
rect 23440 32866 23520 32880
rect 23440 32814 23454 32866
rect 23506 32814 23520 32866
rect 23440 32800 23520 32814
rect 23600 32866 23680 32880
rect 23600 32814 23614 32866
rect 23666 32814 23680 32866
rect 23600 32800 23680 32814
rect 23760 32866 23840 32880
rect 23760 32814 23774 32866
rect 23826 32814 23840 32866
rect 23760 32800 23840 32814
rect 23920 32866 24000 32880
rect 23920 32814 23934 32866
rect 23986 32814 24000 32866
rect 23920 32800 24000 32814
rect 24080 32866 24160 32880
rect 24080 32814 24094 32866
rect 24146 32814 24160 32866
rect 24080 32800 24160 32814
rect 24240 32866 24320 32880
rect 24240 32814 24254 32866
rect 24306 32814 24320 32866
rect 24240 32800 24320 32814
rect 24400 32866 24480 32880
rect 24400 32814 24414 32866
rect 24466 32814 24480 32866
rect 24400 32800 24480 32814
rect 24560 32866 24640 32880
rect 24560 32814 24574 32866
rect 24626 32814 24640 32866
rect 24560 32800 24640 32814
rect 24720 32866 24800 32880
rect 24720 32814 24734 32866
rect 24786 32814 24800 32866
rect 24720 32800 24800 32814
rect 24880 32866 24960 32880
rect 24880 32814 24894 32866
rect 24946 32814 24960 32866
rect 24880 32800 24960 32814
rect 25040 32866 25120 32880
rect 25040 32814 25054 32866
rect 25106 32814 25120 32866
rect 25040 32800 25120 32814
rect 25200 32866 25280 32880
rect 25200 32814 25214 32866
rect 25266 32814 25280 32866
rect 25200 32800 25280 32814
rect 25360 32866 25440 32880
rect 25360 32814 25374 32866
rect 25426 32814 25440 32866
rect 25360 32800 25440 32814
rect 25520 32866 25600 32880
rect 25520 32814 25534 32866
rect 25586 32814 25600 32866
rect 25520 32800 25600 32814
rect 25680 32866 25760 32880
rect 25680 32814 25694 32866
rect 25746 32814 25760 32866
rect 25680 32800 25760 32814
rect 25840 32866 25920 32880
rect 25840 32814 25854 32866
rect 25906 32814 25920 32866
rect 25840 32800 25920 32814
rect 26000 32866 26080 32880
rect 26000 32814 26014 32866
rect 26066 32814 26080 32866
rect 26000 32800 26080 32814
rect 26160 32866 26240 32880
rect 26160 32814 26174 32866
rect 26226 32814 26240 32866
rect 26160 32800 26240 32814
rect 26320 32866 26400 32880
rect 26320 32814 26334 32866
rect 26386 32814 26400 32866
rect 26320 32800 26400 32814
rect 26480 32866 26560 32880
rect 26480 32814 26494 32866
rect 26546 32814 26560 32866
rect 26480 32800 26560 32814
rect 26640 32866 26720 32880
rect 26640 32814 26654 32866
rect 26706 32814 26720 32866
rect 26640 32800 26720 32814
rect 26800 32866 26880 32880
rect 26800 32814 26814 32866
rect 26866 32814 26880 32866
rect 26800 32800 26880 32814
rect 26960 32866 27040 32880
rect 26960 32814 26974 32866
rect 27026 32814 27040 32866
rect 26960 32800 27040 32814
rect 27120 32866 27200 32880
rect 27120 32814 27134 32866
rect 27186 32814 27200 32866
rect 27120 32800 27200 32814
rect 27280 32866 27360 32880
rect 27280 32814 27294 32866
rect 27346 32814 27360 32866
rect 27280 32800 27360 32814
rect 27440 32866 27520 32880
rect 27440 32814 27454 32866
rect 27506 32814 27520 32866
rect 27440 32800 27520 32814
rect 27600 32866 27680 32880
rect 27600 32814 27614 32866
rect 27666 32814 27680 32866
rect 27600 32800 27680 32814
rect 27760 32866 27840 32880
rect 27760 32814 27774 32866
rect 27826 32814 27840 32866
rect 27760 32800 27840 32814
rect 27920 32866 28000 32880
rect 27920 32814 27934 32866
rect 27986 32814 28000 32866
rect 27920 32800 28000 32814
rect 28080 32866 28160 32880
rect 28080 32814 28094 32866
rect 28146 32814 28160 32866
rect 28080 32800 28160 32814
rect 28240 32866 28320 32880
rect 28240 32814 28254 32866
rect 28306 32814 28320 32866
rect 28240 32800 28320 32814
rect 28400 32866 28480 32880
rect 28400 32814 28414 32866
rect 28466 32814 28480 32866
rect 28400 32800 28480 32814
rect 28560 32866 28640 32880
rect 28560 32814 28574 32866
rect 28626 32814 28640 32866
rect 28560 32800 28640 32814
rect 28720 32866 28800 32880
rect 28720 32814 28734 32866
rect 28786 32814 28800 32866
rect 28720 32800 28800 32814
rect 28880 32866 28960 32880
rect 28880 32814 28894 32866
rect 28946 32814 28960 32866
rect 28880 32800 28960 32814
rect 29040 32866 29120 32880
rect 29040 32814 29054 32866
rect 29106 32814 29120 32866
rect 29040 32800 29120 32814
rect 29200 32866 29280 32880
rect 29200 32814 29214 32866
rect 29266 32814 29280 32866
rect 29200 32800 29280 32814
rect 29360 32866 29440 32880
rect 29360 32814 29374 32866
rect 29426 32814 29440 32866
rect 29360 32800 29440 32814
rect 33520 32866 33600 32880
rect 33520 32814 33534 32866
rect 33586 32814 33600 32866
rect 33520 32800 33600 32814
rect 33680 32866 33760 32880
rect 33680 32814 33694 32866
rect 33746 32814 33760 32866
rect 33680 32800 33760 32814
rect 33840 32866 33920 32880
rect 33840 32814 33854 32866
rect 33906 32814 33920 32866
rect 33840 32800 33920 32814
rect 34000 32866 34080 32880
rect 34000 32814 34014 32866
rect 34066 32814 34080 32866
rect 34000 32800 34080 32814
rect 34160 32866 34240 32880
rect 34160 32814 34174 32866
rect 34226 32814 34240 32866
rect 34160 32800 34240 32814
rect 34320 32866 34400 32880
rect 34320 32814 34334 32866
rect 34386 32814 34400 32866
rect 34320 32800 34400 32814
rect 34480 32866 34560 32880
rect 34480 32814 34494 32866
rect 34546 32814 34560 32866
rect 34480 32800 34560 32814
rect 34640 32866 34720 32880
rect 34640 32814 34654 32866
rect 34706 32814 34720 32866
rect 34640 32800 34720 32814
rect 34800 32866 34880 32880
rect 34800 32814 34814 32866
rect 34866 32814 34880 32866
rect 34800 32800 34880 32814
rect 34960 32866 35040 32880
rect 34960 32814 34974 32866
rect 35026 32814 35040 32866
rect 34960 32800 35040 32814
rect 35120 32866 35200 32880
rect 35120 32814 35134 32866
rect 35186 32814 35200 32866
rect 35120 32800 35200 32814
rect 35280 32866 35360 32880
rect 35280 32814 35294 32866
rect 35346 32814 35360 32866
rect 35280 32800 35360 32814
rect 35440 32866 35520 32880
rect 35440 32814 35454 32866
rect 35506 32814 35520 32866
rect 35440 32800 35520 32814
rect 35600 32866 35680 32880
rect 35600 32814 35614 32866
rect 35666 32814 35680 32866
rect 35600 32800 35680 32814
rect 35760 32866 35840 32880
rect 35760 32814 35774 32866
rect 35826 32814 35840 32866
rect 35760 32800 35840 32814
rect 35920 32866 36000 32880
rect 35920 32814 35934 32866
rect 35986 32814 36000 32866
rect 35920 32800 36000 32814
rect 36080 32866 36160 32880
rect 36080 32814 36094 32866
rect 36146 32814 36160 32866
rect 36080 32800 36160 32814
rect 36240 32866 36320 32880
rect 36240 32814 36254 32866
rect 36306 32814 36320 32866
rect 36240 32800 36320 32814
rect 36400 32866 36480 32880
rect 36400 32814 36414 32866
rect 36466 32814 36480 32866
rect 36400 32800 36480 32814
rect 36560 32866 36640 32880
rect 36560 32814 36574 32866
rect 36626 32814 36640 32866
rect 36560 32800 36640 32814
rect 36720 32866 36800 32880
rect 36720 32814 36734 32866
rect 36786 32814 36800 32866
rect 36720 32800 36800 32814
rect 36880 32866 36960 32880
rect 36880 32814 36894 32866
rect 36946 32814 36960 32866
rect 36880 32800 36960 32814
rect 37040 32866 37120 32880
rect 37040 32814 37054 32866
rect 37106 32814 37120 32866
rect 37040 32800 37120 32814
rect 37200 32866 37280 32880
rect 37200 32814 37214 32866
rect 37266 32814 37280 32866
rect 37200 32800 37280 32814
rect 37360 32866 37440 32880
rect 37360 32814 37374 32866
rect 37426 32814 37440 32866
rect 37360 32800 37440 32814
rect 37520 32866 37600 32880
rect 37520 32814 37534 32866
rect 37586 32814 37600 32866
rect 37520 32800 37600 32814
rect 37680 32866 37760 32880
rect 37680 32814 37694 32866
rect 37746 32814 37760 32866
rect 37680 32800 37760 32814
rect 37840 32866 37920 32880
rect 37840 32814 37854 32866
rect 37906 32814 37920 32866
rect 37840 32800 37920 32814
rect 38000 32866 38080 32880
rect 38000 32814 38014 32866
rect 38066 32814 38080 32866
rect 38000 32800 38080 32814
rect 38160 32866 38240 32880
rect 38160 32814 38174 32866
rect 38226 32814 38240 32866
rect 38160 32800 38240 32814
rect 38320 32866 38400 32880
rect 38320 32814 38334 32866
rect 38386 32814 38400 32866
rect 38320 32800 38400 32814
rect 38480 32866 38560 32880
rect 38480 32814 38494 32866
rect 38546 32814 38560 32866
rect 38480 32800 38560 32814
rect 38640 32866 38720 32880
rect 38640 32814 38654 32866
rect 38706 32814 38720 32866
rect 38640 32800 38720 32814
rect 38800 32866 38880 32880
rect 38800 32814 38814 32866
rect 38866 32814 38880 32866
rect 38800 32800 38880 32814
rect 38960 32866 39040 32880
rect 38960 32814 38974 32866
rect 39026 32814 39040 32866
rect 38960 32800 39040 32814
rect 39120 32866 39200 32880
rect 39120 32814 39134 32866
rect 39186 32814 39200 32866
rect 39120 32800 39200 32814
rect 39280 32866 39360 32880
rect 39280 32814 39294 32866
rect 39346 32814 39360 32866
rect 39280 32800 39360 32814
rect 39440 32866 39520 32880
rect 39440 32814 39454 32866
rect 39506 32814 39520 32866
rect 39440 32800 39520 32814
rect 39600 32866 39680 32880
rect 39600 32814 39614 32866
rect 39666 32814 39680 32866
rect 39600 32800 39680 32814
rect 39760 32866 39840 32880
rect 39760 32814 39774 32866
rect 39826 32814 39840 32866
rect 39760 32800 39840 32814
rect 39920 32866 40000 32880
rect 39920 32814 39934 32866
rect 39986 32814 40000 32866
rect 39920 32800 40000 32814
rect 40080 32866 40160 32880
rect 40080 32814 40094 32866
rect 40146 32814 40160 32866
rect 40080 32800 40160 32814
rect 40240 32866 40320 32880
rect 40240 32814 40254 32866
rect 40306 32814 40320 32866
rect 40240 32800 40320 32814
rect 40400 32866 40480 32880
rect 40400 32814 40414 32866
rect 40466 32814 40480 32866
rect 40400 32800 40480 32814
rect 40560 32866 40640 32880
rect 40560 32814 40574 32866
rect 40626 32814 40640 32866
rect 40560 32800 40640 32814
rect 40720 32866 40800 32880
rect 40720 32814 40734 32866
rect 40786 32814 40800 32866
rect 40720 32800 40800 32814
rect 40880 32866 40960 32880
rect 40880 32814 40894 32866
rect 40946 32814 40960 32866
rect 40880 32800 40960 32814
rect 41040 32866 41120 32880
rect 41040 32814 41054 32866
rect 41106 32814 41120 32866
rect 41040 32800 41120 32814
rect 41200 32866 41280 32880
rect 41200 32814 41214 32866
rect 41266 32814 41280 32866
rect 41200 32800 41280 32814
rect 41360 32866 41440 32880
rect 41360 32814 41374 32866
rect 41426 32814 41440 32866
rect 41360 32800 41440 32814
rect 41520 32866 41600 32880
rect 41520 32814 41534 32866
rect 41586 32814 41600 32866
rect 41520 32800 41600 32814
rect 41680 32866 41760 32880
rect 41680 32814 41694 32866
rect 41746 32814 41760 32866
rect 41680 32800 41760 32814
rect 41840 32866 41920 32880
rect 41840 32814 41854 32866
rect 41906 32814 41920 32866
rect 41840 32800 41920 32814
rect 0 32546 80 32560
rect 0 32494 14 32546
rect 66 32494 80 32546
rect 0 32480 80 32494
rect 160 32546 240 32560
rect 160 32494 174 32546
rect 226 32494 240 32546
rect 160 32480 240 32494
rect 320 32546 400 32560
rect 320 32494 334 32546
rect 386 32494 400 32546
rect 320 32480 400 32494
rect 480 32546 560 32560
rect 480 32494 494 32546
rect 546 32494 560 32546
rect 480 32480 560 32494
rect 640 32546 720 32560
rect 640 32494 654 32546
rect 706 32494 720 32546
rect 640 32480 720 32494
rect 800 32546 880 32560
rect 800 32494 814 32546
rect 866 32494 880 32546
rect 800 32480 880 32494
rect 960 32546 1040 32560
rect 960 32494 974 32546
rect 1026 32494 1040 32546
rect 960 32480 1040 32494
rect 1120 32546 1200 32560
rect 1120 32494 1134 32546
rect 1186 32494 1200 32546
rect 1120 32480 1200 32494
rect 1280 32546 1360 32560
rect 1280 32494 1294 32546
rect 1346 32494 1360 32546
rect 1280 32480 1360 32494
rect 1440 32546 1520 32560
rect 1440 32494 1454 32546
rect 1506 32494 1520 32546
rect 1440 32480 1520 32494
rect 1600 32546 1680 32560
rect 1600 32494 1614 32546
rect 1666 32494 1680 32546
rect 1600 32480 1680 32494
rect 1760 32546 1840 32560
rect 1760 32494 1774 32546
rect 1826 32494 1840 32546
rect 1760 32480 1840 32494
rect 1920 32546 2000 32560
rect 1920 32494 1934 32546
rect 1986 32494 2000 32546
rect 1920 32480 2000 32494
rect 2080 32546 2160 32560
rect 2080 32494 2094 32546
rect 2146 32494 2160 32546
rect 2080 32480 2160 32494
rect 2240 32546 2320 32560
rect 2240 32494 2254 32546
rect 2306 32494 2320 32546
rect 2240 32480 2320 32494
rect 2400 32546 2480 32560
rect 2400 32494 2414 32546
rect 2466 32494 2480 32546
rect 2400 32480 2480 32494
rect 2560 32546 2640 32560
rect 2560 32494 2574 32546
rect 2626 32494 2640 32546
rect 2560 32480 2640 32494
rect 2720 32546 2800 32560
rect 2720 32494 2734 32546
rect 2786 32494 2800 32546
rect 2720 32480 2800 32494
rect 2880 32546 2960 32560
rect 2880 32494 2894 32546
rect 2946 32494 2960 32546
rect 2880 32480 2960 32494
rect 3040 32546 3120 32560
rect 3040 32494 3054 32546
rect 3106 32494 3120 32546
rect 3040 32480 3120 32494
rect 3200 32546 3280 32560
rect 3200 32494 3214 32546
rect 3266 32494 3280 32546
rect 3200 32480 3280 32494
rect 3360 32546 3440 32560
rect 3360 32494 3374 32546
rect 3426 32494 3440 32546
rect 3360 32480 3440 32494
rect 3520 32546 3600 32560
rect 3520 32494 3534 32546
rect 3586 32494 3600 32546
rect 3520 32480 3600 32494
rect 3680 32546 3760 32560
rect 3680 32494 3694 32546
rect 3746 32494 3760 32546
rect 3680 32480 3760 32494
rect 3840 32546 3920 32560
rect 3840 32494 3854 32546
rect 3906 32494 3920 32546
rect 3840 32480 3920 32494
rect 4000 32546 4080 32560
rect 4000 32494 4014 32546
rect 4066 32494 4080 32546
rect 4000 32480 4080 32494
rect 4160 32546 4240 32560
rect 4160 32494 4174 32546
rect 4226 32494 4240 32546
rect 4160 32480 4240 32494
rect 4320 32546 4400 32560
rect 4320 32494 4334 32546
rect 4386 32494 4400 32546
rect 4320 32480 4400 32494
rect 4480 32546 4560 32560
rect 4480 32494 4494 32546
rect 4546 32494 4560 32546
rect 4480 32480 4560 32494
rect 4640 32546 4720 32560
rect 4640 32494 4654 32546
rect 4706 32494 4720 32546
rect 4640 32480 4720 32494
rect 4800 32546 4880 32560
rect 4800 32494 4814 32546
rect 4866 32494 4880 32546
rect 4800 32480 4880 32494
rect 4960 32546 5040 32560
rect 4960 32494 4974 32546
rect 5026 32494 5040 32546
rect 4960 32480 5040 32494
rect 5120 32546 5200 32560
rect 5120 32494 5134 32546
rect 5186 32494 5200 32546
rect 5120 32480 5200 32494
rect 5280 32546 5360 32560
rect 5280 32494 5294 32546
rect 5346 32494 5360 32546
rect 5280 32480 5360 32494
rect 5440 32546 5520 32560
rect 5440 32494 5454 32546
rect 5506 32494 5520 32546
rect 5440 32480 5520 32494
rect 5600 32546 5680 32560
rect 5600 32494 5614 32546
rect 5666 32494 5680 32546
rect 5600 32480 5680 32494
rect 5760 32546 5840 32560
rect 5760 32494 5774 32546
rect 5826 32494 5840 32546
rect 5760 32480 5840 32494
rect 5920 32546 6000 32560
rect 5920 32494 5934 32546
rect 5986 32494 6000 32546
rect 5920 32480 6000 32494
rect 6080 32546 6160 32560
rect 6080 32494 6094 32546
rect 6146 32494 6160 32546
rect 6080 32480 6160 32494
rect 6240 32546 6320 32560
rect 6240 32494 6254 32546
rect 6306 32494 6320 32546
rect 6240 32480 6320 32494
rect 6400 32546 6480 32560
rect 6400 32494 6414 32546
rect 6466 32494 6480 32546
rect 6400 32480 6480 32494
rect 6560 32546 6640 32560
rect 6560 32494 6574 32546
rect 6626 32494 6640 32546
rect 6560 32480 6640 32494
rect 6720 32546 6800 32560
rect 6720 32494 6734 32546
rect 6786 32494 6800 32546
rect 6720 32480 6800 32494
rect 6880 32546 6960 32560
rect 6880 32494 6894 32546
rect 6946 32494 6960 32546
rect 6880 32480 6960 32494
rect 7040 32546 7120 32560
rect 7040 32494 7054 32546
rect 7106 32494 7120 32546
rect 7040 32480 7120 32494
rect 7200 32546 7280 32560
rect 7200 32494 7214 32546
rect 7266 32494 7280 32546
rect 7200 32480 7280 32494
rect 7360 32546 7440 32560
rect 7360 32494 7374 32546
rect 7426 32494 7440 32546
rect 7360 32480 7440 32494
rect 7520 32546 7600 32560
rect 7520 32494 7534 32546
rect 7586 32494 7600 32546
rect 7520 32480 7600 32494
rect 7680 32546 7760 32560
rect 7680 32494 7694 32546
rect 7746 32494 7760 32546
rect 7680 32480 7760 32494
rect 7840 32546 7920 32560
rect 7840 32494 7854 32546
rect 7906 32494 7920 32546
rect 7840 32480 7920 32494
rect 8000 32546 8080 32560
rect 8000 32494 8014 32546
rect 8066 32494 8080 32546
rect 8000 32480 8080 32494
rect 8160 32546 8240 32560
rect 8160 32494 8174 32546
rect 8226 32494 8240 32546
rect 8160 32480 8240 32494
rect 8320 32546 8400 32560
rect 8320 32494 8334 32546
rect 8386 32494 8400 32546
rect 8320 32480 8400 32494
rect 12480 32546 12560 32560
rect 12480 32494 12494 32546
rect 12546 32494 12560 32546
rect 12480 32480 12560 32494
rect 12640 32546 12720 32560
rect 12640 32494 12654 32546
rect 12706 32494 12720 32546
rect 12640 32480 12720 32494
rect 12800 32546 12880 32560
rect 12800 32494 12814 32546
rect 12866 32494 12880 32546
rect 12800 32480 12880 32494
rect 12960 32546 13040 32560
rect 12960 32494 12974 32546
rect 13026 32494 13040 32546
rect 12960 32480 13040 32494
rect 13120 32546 13200 32560
rect 13120 32494 13134 32546
rect 13186 32494 13200 32546
rect 13120 32480 13200 32494
rect 13280 32546 13360 32560
rect 13280 32494 13294 32546
rect 13346 32494 13360 32546
rect 13280 32480 13360 32494
rect 13440 32546 13520 32560
rect 13440 32494 13454 32546
rect 13506 32494 13520 32546
rect 13440 32480 13520 32494
rect 13600 32546 13680 32560
rect 13600 32494 13614 32546
rect 13666 32494 13680 32546
rect 13600 32480 13680 32494
rect 13760 32546 13840 32560
rect 13760 32494 13774 32546
rect 13826 32494 13840 32546
rect 13760 32480 13840 32494
rect 13920 32546 14000 32560
rect 13920 32494 13934 32546
rect 13986 32494 14000 32546
rect 13920 32480 14000 32494
rect 14080 32546 14160 32560
rect 14080 32494 14094 32546
rect 14146 32494 14160 32546
rect 14080 32480 14160 32494
rect 14240 32546 14320 32560
rect 14240 32494 14254 32546
rect 14306 32494 14320 32546
rect 14240 32480 14320 32494
rect 14400 32546 14480 32560
rect 14400 32494 14414 32546
rect 14466 32494 14480 32546
rect 14400 32480 14480 32494
rect 14560 32546 14640 32560
rect 14560 32494 14574 32546
rect 14626 32494 14640 32546
rect 14560 32480 14640 32494
rect 14720 32546 14800 32560
rect 14720 32494 14734 32546
rect 14786 32494 14800 32546
rect 14720 32480 14800 32494
rect 14880 32546 14960 32560
rect 14880 32494 14894 32546
rect 14946 32494 14960 32546
rect 14880 32480 14960 32494
rect 15040 32546 15120 32560
rect 15040 32494 15054 32546
rect 15106 32494 15120 32546
rect 15040 32480 15120 32494
rect 15200 32546 15280 32560
rect 15200 32494 15214 32546
rect 15266 32494 15280 32546
rect 15200 32480 15280 32494
rect 15360 32546 15440 32560
rect 15360 32494 15374 32546
rect 15426 32494 15440 32546
rect 15360 32480 15440 32494
rect 15520 32546 15600 32560
rect 15520 32494 15534 32546
rect 15586 32494 15600 32546
rect 15520 32480 15600 32494
rect 15680 32546 15760 32560
rect 15680 32494 15694 32546
rect 15746 32494 15760 32546
rect 15680 32480 15760 32494
rect 15840 32546 15920 32560
rect 15840 32494 15854 32546
rect 15906 32494 15920 32546
rect 15840 32480 15920 32494
rect 16000 32546 16080 32560
rect 16000 32494 16014 32546
rect 16066 32494 16080 32546
rect 16000 32480 16080 32494
rect 16160 32546 16240 32560
rect 16160 32494 16174 32546
rect 16226 32494 16240 32546
rect 16160 32480 16240 32494
rect 16320 32546 16400 32560
rect 16320 32494 16334 32546
rect 16386 32494 16400 32546
rect 16320 32480 16400 32494
rect 16480 32546 16560 32560
rect 16480 32494 16494 32546
rect 16546 32494 16560 32546
rect 16480 32480 16560 32494
rect 16640 32546 16720 32560
rect 16640 32494 16654 32546
rect 16706 32494 16720 32546
rect 16640 32480 16720 32494
rect 16800 32546 16880 32560
rect 16800 32494 16814 32546
rect 16866 32494 16880 32546
rect 16800 32480 16880 32494
rect 16960 32546 17040 32560
rect 16960 32494 16974 32546
rect 17026 32494 17040 32546
rect 16960 32480 17040 32494
rect 17120 32546 17200 32560
rect 17120 32494 17134 32546
rect 17186 32494 17200 32546
rect 17120 32480 17200 32494
rect 17280 32546 17360 32560
rect 17280 32494 17294 32546
rect 17346 32494 17360 32546
rect 17280 32480 17360 32494
rect 17440 32546 17520 32560
rect 17440 32494 17454 32546
rect 17506 32494 17520 32546
rect 17440 32480 17520 32494
rect 17600 32546 17680 32560
rect 17600 32494 17614 32546
rect 17666 32494 17680 32546
rect 17600 32480 17680 32494
rect 17760 32546 17840 32560
rect 17760 32494 17774 32546
rect 17826 32494 17840 32546
rect 17760 32480 17840 32494
rect 17920 32546 18000 32560
rect 17920 32494 17934 32546
rect 17986 32494 18000 32546
rect 17920 32480 18000 32494
rect 18080 32546 18160 32560
rect 18080 32494 18094 32546
rect 18146 32494 18160 32546
rect 18080 32480 18160 32494
rect 18240 32546 18320 32560
rect 18240 32494 18254 32546
rect 18306 32494 18320 32546
rect 18240 32480 18320 32494
rect 18400 32546 18480 32560
rect 18400 32494 18414 32546
rect 18466 32494 18480 32546
rect 18400 32480 18480 32494
rect 18560 32546 18640 32560
rect 18560 32494 18574 32546
rect 18626 32494 18640 32546
rect 18560 32480 18640 32494
rect 18720 32546 18800 32560
rect 18720 32494 18734 32546
rect 18786 32494 18800 32546
rect 18720 32480 18800 32494
rect 18880 32546 18960 32560
rect 18880 32494 18894 32546
rect 18946 32494 18960 32546
rect 18880 32480 18960 32494
rect 23120 32546 23200 32560
rect 23120 32494 23134 32546
rect 23186 32494 23200 32546
rect 23120 32480 23200 32494
rect 23280 32546 23360 32560
rect 23280 32494 23294 32546
rect 23346 32494 23360 32546
rect 23280 32480 23360 32494
rect 23440 32546 23520 32560
rect 23440 32494 23454 32546
rect 23506 32494 23520 32546
rect 23440 32480 23520 32494
rect 23600 32546 23680 32560
rect 23600 32494 23614 32546
rect 23666 32494 23680 32546
rect 23600 32480 23680 32494
rect 23760 32546 23840 32560
rect 23760 32494 23774 32546
rect 23826 32494 23840 32546
rect 23760 32480 23840 32494
rect 23920 32546 24000 32560
rect 23920 32494 23934 32546
rect 23986 32494 24000 32546
rect 23920 32480 24000 32494
rect 24080 32546 24160 32560
rect 24080 32494 24094 32546
rect 24146 32494 24160 32546
rect 24080 32480 24160 32494
rect 24240 32546 24320 32560
rect 24240 32494 24254 32546
rect 24306 32494 24320 32546
rect 24240 32480 24320 32494
rect 24400 32546 24480 32560
rect 24400 32494 24414 32546
rect 24466 32494 24480 32546
rect 24400 32480 24480 32494
rect 24560 32546 24640 32560
rect 24560 32494 24574 32546
rect 24626 32494 24640 32546
rect 24560 32480 24640 32494
rect 24720 32546 24800 32560
rect 24720 32494 24734 32546
rect 24786 32494 24800 32546
rect 24720 32480 24800 32494
rect 24880 32546 24960 32560
rect 24880 32494 24894 32546
rect 24946 32494 24960 32546
rect 24880 32480 24960 32494
rect 25040 32546 25120 32560
rect 25040 32494 25054 32546
rect 25106 32494 25120 32546
rect 25040 32480 25120 32494
rect 25200 32546 25280 32560
rect 25200 32494 25214 32546
rect 25266 32494 25280 32546
rect 25200 32480 25280 32494
rect 25360 32546 25440 32560
rect 25360 32494 25374 32546
rect 25426 32494 25440 32546
rect 25360 32480 25440 32494
rect 25520 32546 25600 32560
rect 25520 32494 25534 32546
rect 25586 32494 25600 32546
rect 25520 32480 25600 32494
rect 25680 32546 25760 32560
rect 25680 32494 25694 32546
rect 25746 32494 25760 32546
rect 25680 32480 25760 32494
rect 25840 32546 25920 32560
rect 25840 32494 25854 32546
rect 25906 32494 25920 32546
rect 25840 32480 25920 32494
rect 26000 32546 26080 32560
rect 26000 32494 26014 32546
rect 26066 32494 26080 32546
rect 26000 32480 26080 32494
rect 26160 32546 26240 32560
rect 26160 32494 26174 32546
rect 26226 32494 26240 32546
rect 26160 32480 26240 32494
rect 26320 32546 26400 32560
rect 26320 32494 26334 32546
rect 26386 32494 26400 32546
rect 26320 32480 26400 32494
rect 26480 32546 26560 32560
rect 26480 32494 26494 32546
rect 26546 32494 26560 32546
rect 26480 32480 26560 32494
rect 26640 32546 26720 32560
rect 26640 32494 26654 32546
rect 26706 32494 26720 32546
rect 26640 32480 26720 32494
rect 26800 32546 26880 32560
rect 26800 32494 26814 32546
rect 26866 32494 26880 32546
rect 26800 32480 26880 32494
rect 26960 32546 27040 32560
rect 26960 32494 26974 32546
rect 27026 32494 27040 32546
rect 26960 32480 27040 32494
rect 27120 32546 27200 32560
rect 27120 32494 27134 32546
rect 27186 32494 27200 32546
rect 27120 32480 27200 32494
rect 27280 32546 27360 32560
rect 27280 32494 27294 32546
rect 27346 32494 27360 32546
rect 27280 32480 27360 32494
rect 27440 32546 27520 32560
rect 27440 32494 27454 32546
rect 27506 32494 27520 32546
rect 27440 32480 27520 32494
rect 27600 32546 27680 32560
rect 27600 32494 27614 32546
rect 27666 32494 27680 32546
rect 27600 32480 27680 32494
rect 27760 32546 27840 32560
rect 27760 32494 27774 32546
rect 27826 32494 27840 32546
rect 27760 32480 27840 32494
rect 27920 32546 28000 32560
rect 27920 32494 27934 32546
rect 27986 32494 28000 32546
rect 27920 32480 28000 32494
rect 28080 32546 28160 32560
rect 28080 32494 28094 32546
rect 28146 32494 28160 32546
rect 28080 32480 28160 32494
rect 28240 32546 28320 32560
rect 28240 32494 28254 32546
rect 28306 32494 28320 32546
rect 28240 32480 28320 32494
rect 28400 32546 28480 32560
rect 28400 32494 28414 32546
rect 28466 32494 28480 32546
rect 28400 32480 28480 32494
rect 28560 32546 28640 32560
rect 28560 32494 28574 32546
rect 28626 32494 28640 32546
rect 28560 32480 28640 32494
rect 28720 32546 28800 32560
rect 28720 32494 28734 32546
rect 28786 32494 28800 32546
rect 28720 32480 28800 32494
rect 28880 32546 28960 32560
rect 28880 32494 28894 32546
rect 28946 32494 28960 32546
rect 28880 32480 28960 32494
rect 29040 32546 29120 32560
rect 29040 32494 29054 32546
rect 29106 32494 29120 32546
rect 29040 32480 29120 32494
rect 29200 32546 29280 32560
rect 29200 32494 29214 32546
rect 29266 32494 29280 32546
rect 29200 32480 29280 32494
rect 29360 32546 29440 32560
rect 29360 32494 29374 32546
rect 29426 32494 29440 32546
rect 29360 32480 29440 32494
rect 33520 32546 33600 32560
rect 33520 32494 33534 32546
rect 33586 32494 33600 32546
rect 33520 32480 33600 32494
rect 33680 32546 33760 32560
rect 33680 32494 33694 32546
rect 33746 32494 33760 32546
rect 33680 32480 33760 32494
rect 33840 32546 33920 32560
rect 33840 32494 33854 32546
rect 33906 32494 33920 32546
rect 33840 32480 33920 32494
rect 34000 32546 34080 32560
rect 34000 32494 34014 32546
rect 34066 32494 34080 32546
rect 34000 32480 34080 32494
rect 34160 32546 34240 32560
rect 34160 32494 34174 32546
rect 34226 32494 34240 32546
rect 34160 32480 34240 32494
rect 34320 32546 34400 32560
rect 34320 32494 34334 32546
rect 34386 32494 34400 32546
rect 34320 32480 34400 32494
rect 34480 32546 34560 32560
rect 34480 32494 34494 32546
rect 34546 32494 34560 32546
rect 34480 32480 34560 32494
rect 34640 32546 34720 32560
rect 34640 32494 34654 32546
rect 34706 32494 34720 32546
rect 34640 32480 34720 32494
rect 34800 32546 34880 32560
rect 34800 32494 34814 32546
rect 34866 32494 34880 32546
rect 34800 32480 34880 32494
rect 34960 32546 35040 32560
rect 34960 32494 34974 32546
rect 35026 32494 35040 32546
rect 34960 32480 35040 32494
rect 35120 32546 35200 32560
rect 35120 32494 35134 32546
rect 35186 32494 35200 32546
rect 35120 32480 35200 32494
rect 35280 32546 35360 32560
rect 35280 32494 35294 32546
rect 35346 32494 35360 32546
rect 35280 32480 35360 32494
rect 35440 32546 35520 32560
rect 35440 32494 35454 32546
rect 35506 32494 35520 32546
rect 35440 32480 35520 32494
rect 35600 32546 35680 32560
rect 35600 32494 35614 32546
rect 35666 32494 35680 32546
rect 35600 32480 35680 32494
rect 35760 32546 35840 32560
rect 35760 32494 35774 32546
rect 35826 32494 35840 32546
rect 35760 32480 35840 32494
rect 35920 32546 36000 32560
rect 35920 32494 35934 32546
rect 35986 32494 36000 32546
rect 35920 32480 36000 32494
rect 36080 32546 36160 32560
rect 36080 32494 36094 32546
rect 36146 32494 36160 32546
rect 36080 32480 36160 32494
rect 36240 32546 36320 32560
rect 36240 32494 36254 32546
rect 36306 32494 36320 32546
rect 36240 32480 36320 32494
rect 36400 32546 36480 32560
rect 36400 32494 36414 32546
rect 36466 32494 36480 32546
rect 36400 32480 36480 32494
rect 36560 32546 36640 32560
rect 36560 32494 36574 32546
rect 36626 32494 36640 32546
rect 36560 32480 36640 32494
rect 36720 32546 36800 32560
rect 36720 32494 36734 32546
rect 36786 32494 36800 32546
rect 36720 32480 36800 32494
rect 36880 32546 36960 32560
rect 36880 32494 36894 32546
rect 36946 32494 36960 32546
rect 36880 32480 36960 32494
rect 37040 32546 37120 32560
rect 37040 32494 37054 32546
rect 37106 32494 37120 32546
rect 37040 32480 37120 32494
rect 37200 32546 37280 32560
rect 37200 32494 37214 32546
rect 37266 32494 37280 32546
rect 37200 32480 37280 32494
rect 37360 32546 37440 32560
rect 37360 32494 37374 32546
rect 37426 32494 37440 32546
rect 37360 32480 37440 32494
rect 37520 32546 37600 32560
rect 37520 32494 37534 32546
rect 37586 32494 37600 32546
rect 37520 32480 37600 32494
rect 37680 32546 37760 32560
rect 37680 32494 37694 32546
rect 37746 32494 37760 32546
rect 37680 32480 37760 32494
rect 37840 32546 37920 32560
rect 37840 32494 37854 32546
rect 37906 32494 37920 32546
rect 37840 32480 37920 32494
rect 38000 32546 38080 32560
rect 38000 32494 38014 32546
rect 38066 32494 38080 32546
rect 38000 32480 38080 32494
rect 38160 32546 38240 32560
rect 38160 32494 38174 32546
rect 38226 32494 38240 32546
rect 38160 32480 38240 32494
rect 38320 32546 38400 32560
rect 38320 32494 38334 32546
rect 38386 32494 38400 32546
rect 38320 32480 38400 32494
rect 38480 32546 38560 32560
rect 38480 32494 38494 32546
rect 38546 32494 38560 32546
rect 38480 32480 38560 32494
rect 38640 32546 38720 32560
rect 38640 32494 38654 32546
rect 38706 32494 38720 32546
rect 38640 32480 38720 32494
rect 38800 32546 38880 32560
rect 38800 32494 38814 32546
rect 38866 32494 38880 32546
rect 38800 32480 38880 32494
rect 38960 32546 39040 32560
rect 38960 32494 38974 32546
rect 39026 32494 39040 32546
rect 38960 32480 39040 32494
rect 39120 32546 39200 32560
rect 39120 32494 39134 32546
rect 39186 32494 39200 32546
rect 39120 32480 39200 32494
rect 39280 32546 39360 32560
rect 39280 32494 39294 32546
rect 39346 32494 39360 32546
rect 39280 32480 39360 32494
rect 39440 32546 39520 32560
rect 39440 32494 39454 32546
rect 39506 32494 39520 32546
rect 39440 32480 39520 32494
rect 39600 32546 39680 32560
rect 39600 32494 39614 32546
rect 39666 32494 39680 32546
rect 39600 32480 39680 32494
rect 39760 32546 39840 32560
rect 39760 32494 39774 32546
rect 39826 32494 39840 32546
rect 39760 32480 39840 32494
rect 39920 32546 40000 32560
rect 39920 32494 39934 32546
rect 39986 32494 40000 32546
rect 39920 32480 40000 32494
rect 40080 32546 40160 32560
rect 40080 32494 40094 32546
rect 40146 32494 40160 32546
rect 40080 32480 40160 32494
rect 40240 32546 40320 32560
rect 40240 32494 40254 32546
rect 40306 32494 40320 32546
rect 40240 32480 40320 32494
rect 40400 32546 40480 32560
rect 40400 32494 40414 32546
rect 40466 32494 40480 32546
rect 40400 32480 40480 32494
rect 40560 32546 40640 32560
rect 40560 32494 40574 32546
rect 40626 32494 40640 32546
rect 40560 32480 40640 32494
rect 40720 32546 40800 32560
rect 40720 32494 40734 32546
rect 40786 32494 40800 32546
rect 40720 32480 40800 32494
rect 40880 32546 40960 32560
rect 40880 32494 40894 32546
rect 40946 32494 40960 32546
rect 40880 32480 40960 32494
rect 41040 32546 41120 32560
rect 41040 32494 41054 32546
rect 41106 32494 41120 32546
rect 41040 32480 41120 32494
rect 41200 32546 41280 32560
rect 41200 32494 41214 32546
rect 41266 32494 41280 32546
rect 41200 32480 41280 32494
rect 41360 32546 41440 32560
rect 41360 32494 41374 32546
rect 41426 32494 41440 32546
rect 41360 32480 41440 32494
rect 41520 32546 41600 32560
rect 41520 32494 41534 32546
rect 41586 32494 41600 32546
rect 41520 32480 41600 32494
rect 41680 32546 41760 32560
rect 41680 32494 41694 32546
rect 41746 32494 41760 32546
rect 41680 32480 41760 32494
rect 41840 32546 41920 32560
rect 41840 32494 41854 32546
rect 41906 32494 41920 32546
rect 41840 32480 41920 32494
rect 0 32386 80 32400
rect 0 32334 14 32386
rect 66 32334 80 32386
rect 0 32320 80 32334
rect 160 32386 240 32400
rect 160 32334 174 32386
rect 226 32334 240 32386
rect 160 32320 240 32334
rect 320 32386 400 32400
rect 320 32334 334 32386
rect 386 32334 400 32386
rect 320 32320 400 32334
rect 480 32386 560 32400
rect 480 32334 494 32386
rect 546 32334 560 32386
rect 480 32320 560 32334
rect 640 32386 720 32400
rect 640 32334 654 32386
rect 706 32334 720 32386
rect 640 32320 720 32334
rect 800 32386 880 32400
rect 800 32334 814 32386
rect 866 32334 880 32386
rect 800 32320 880 32334
rect 960 32386 1040 32400
rect 960 32334 974 32386
rect 1026 32334 1040 32386
rect 960 32320 1040 32334
rect 1120 32386 1200 32400
rect 1120 32334 1134 32386
rect 1186 32334 1200 32386
rect 1120 32320 1200 32334
rect 1280 32386 1360 32400
rect 1280 32334 1294 32386
rect 1346 32334 1360 32386
rect 1280 32320 1360 32334
rect 1440 32386 1520 32400
rect 1440 32334 1454 32386
rect 1506 32334 1520 32386
rect 1440 32320 1520 32334
rect 1600 32386 1680 32400
rect 1600 32334 1614 32386
rect 1666 32334 1680 32386
rect 1600 32320 1680 32334
rect 1760 32386 1840 32400
rect 1760 32334 1774 32386
rect 1826 32334 1840 32386
rect 1760 32320 1840 32334
rect 1920 32386 2000 32400
rect 1920 32334 1934 32386
rect 1986 32334 2000 32386
rect 1920 32320 2000 32334
rect 2080 32386 2160 32400
rect 2080 32334 2094 32386
rect 2146 32334 2160 32386
rect 2080 32320 2160 32334
rect 2240 32386 2320 32400
rect 2240 32334 2254 32386
rect 2306 32334 2320 32386
rect 2240 32320 2320 32334
rect 2400 32386 2480 32400
rect 2400 32334 2414 32386
rect 2466 32334 2480 32386
rect 2400 32320 2480 32334
rect 2560 32386 2640 32400
rect 2560 32334 2574 32386
rect 2626 32334 2640 32386
rect 2560 32320 2640 32334
rect 2720 32386 2800 32400
rect 2720 32334 2734 32386
rect 2786 32334 2800 32386
rect 2720 32320 2800 32334
rect 2880 32386 2960 32400
rect 2880 32334 2894 32386
rect 2946 32334 2960 32386
rect 2880 32320 2960 32334
rect 3040 32386 3120 32400
rect 3040 32334 3054 32386
rect 3106 32334 3120 32386
rect 3040 32320 3120 32334
rect 3200 32386 3280 32400
rect 3200 32334 3214 32386
rect 3266 32334 3280 32386
rect 3200 32320 3280 32334
rect 3360 32386 3440 32400
rect 3360 32334 3374 32386
rect 3426 32334 3440 32386
rect 3360 32320 3440 32334
rect 3520 32386 3600 32400
rect 3520 32334 3534 32386
rect 3586 32334 3600 32386
rect 3520 32320 3600 32334
rect 3680 32386 3760 32400
rect 3680 32334 3694 32386
rect 3746 32334 3760 32386
rect 3680 32320 3760 32334
rect 3840 32386 3920 32400
rect 3840 32334 3854 32386
rect 3906 32334 3920 32386
rect 3840 32320 3920 32334
rect 4000 32386 4080 32400
rect 4000 32334 4014 32386
rect 4066 32334 4080 32386
rect 4000 32320 4080 32334
rect 4160 32386 4240 32400
rect 4160 32334 4174 32386
rect 4226 32334 4240 32386
rect 4160 32320 4240 32334
rect 4320 32386 4400 32400
rect 4320 32334 4334 32386
rect 4386 32334 4400 32386
rect 4320 32320 4400 32334
rect 4480 32386 4560 32400
rect 4480 32334 4494 32386
rect 4546 32334 4560 32386
rect 4480 32320 4560 32334
rect 4640 32386 4720 32400
rect 4640 32334 4654 32386
rect 4706 32334 4720 32386
rect 4640 32320 4720 32334
rect 4800 32386 4880 32400
rect 4800 32334 4814 32386
rect 4866 32334 4880 32386
rect 4800 32320 4880 32334
rect 4960 32386 5040 32400
rect 4960 32334 4974 32386
rect 5026 32334 5040 32386
rect 4960 32320 5040 32334
rect 5120 32386 5200 32400
rect 5120 32334 5134 32386
rect 5186 32334 5200 32386
rect 5120 32320 5200 32334
rect 5280 32386 5360 32400
rect 5280 32334 5294 32386
rect 5346 32334 5360 32386
rect 5280 32320 5360 32334
rect 5440 32386 5520 32400
rect 5440 32334 5454 32386
rect 5506 32334 5520 32386
rect 5440 32320 5520 32334
rect 5600 32386 5680 32400
rect 5600 32334 5614 32386
rect 5666 32334 5680 32386
rect 5600 32320 5680 32334
rect 5760 32386 5840 32400
rect 5760 32334 5774 32386
rect 5826 32334 5840 32386
rect 5760 32320 5840 32334
rect 5920 32386 6000 32400
rect 5920 32334 5934 32386
rect 5986 32334 6000 32386
rect 5920 32320 6000 32334
rect 6080 32386 6160 32400
rect 6080 32334 6094 32386
rect 6146 32334 6160 32386
rect 6080 32320 6160 32334
rect 6240 32386 6320 32400
rect 6240 32334 6254 32386
rect 6306 32334 6320 32386
rect 6240 32320 6320 32334
rect 6400 32386 6480 32400
rect 6400 32334 6414 32386
rect 6466 32334 6480 32386
rect 6400 32320 6480 32334
rect 6560 32386 6640 32400
rect 6560 32334 6574 32386
rect 6626 32334 6640 32386
rect 6560 32320 6640 32334
rect 6720 32386 6800 32400
rect 6720 32334 6734 32386
rect 6786 32334 6800 32386
rect 6720 32320 6800 32334
rect 6880 32386 6960 32400
rect 6880 32334 6894 32386
rect 6946 32334 6960 32386
rect 6880 32320 6960 32334
rect 7040 32386 7120 32400
rect 7040 32334 7054 32386
rect 7106 32334 7120 32386
rect 7040 32320 7120 32334
rect 7200 32386 7280 32400
rect 7200 32334 7214 32386
rect 7266 32334 7280 32386
rect 7200 32320 7280 32334
rect 7360 32386 7440 32400
rect 7360 32334 7374 32386
rect 7426 32334 7440 32386
rect 7360 32320 7440 32334
rect 7520 32386 7600 32400
rect 7520 32334 7534 32386
rect 7586 32334 7600 32386
rect 7520 32320 7600 32334
rect 7680 32386 7760 32400
rect 7680 32334 7694 32386
rect 7746 32334 7760 32386
rect 7680 32320 7760 32334
rect 7840 32386 7920 32400
rect 7840 32334 7854 32386
rect 7906 32334 7920 32386
rect 7840 32320 7920 32334
rect 8000 32386 8080 32400
rect 8000 32334 8014 32386
rect 8066 32334 8080 32386
rect 8000 32320 8080 32334
rect 8160 32386 8240 32400
rect 8160 32334 8174 32386
rect 8226 32334 8240 32386
rect 8160 32320 8240 32334
rect 8320 32386 8400 32400
rect 8320 32334 8334 32386
rect 8386 32334 8400 32386
rect 8320 32320 8400 32334
rect 12480 32386 12560 32400
rect 12480 32334 12494 32386
rect 12546 32334 12560 32386
rect 12480 32320 12560 32334
rect 12640 32386 12720 32400
rect 12640 32334 12654 32386
rect 12706 32334 12720 32386
rect 12640 32320 12720 32334
rect 12800 32386 12880 32400
rect 12800 32334 12814 32386
rect 12866 32334 12880 32386
rect 12800 32320 12880 32334
rect 12960 32386 13040 32400
rect 12960 32334 12974 32386
rect 13026 32334 13040 32386
rect 12960 32320 13040 32334
rect 13120 32386 13200 32400
rect 13120 32334 13134 32386
rect 13186 32334 13200 32386
rect 13120 32320 13200 32334
rect 13280 32386 13360 32400
rect 13280 32334 13294 32386
rect 13346 32334 13360 32386
rect 13280 32320 13360 32334
rect 13440 32386 13520 32400
rect 13440 32334 13454 32386
rect 13506 32334 13520 32386
rect 13440 32320 13520 32334
rect 13600 32386 13680 32400
rect 13600 32334 13614 32386
rect 13666 32334 13680 32386
rect 13600 32320 13680 32334
rect 13760 32386 13840 32400
rect 13760 32334 13774 32386
rect 13826 32334 13840 32386
rect 13760 32320 13840 32334
rect 13920 32386 14000 32400
rect 13920 32334 13934 32386
rect 13986 32334 14000 32386
rect 13920 32320 14000 32334
rect 14080 32386 14160 32400
rect 14080 32334 14094 32386
rect 14146 32334 14160 32386
rect 14080 32320 14160 32334
rect 14240 32386 14320 32400
rect 14240 32334 14254 32386
rect 14306 32334 14320 32386
rect 14240 32320 14320 32334
rect 14400 32386 14480 32400
rect 14400 32334 14414 32386
rect 14466 32334 14480 32386
rect 14400 32320 14480 32334
rect 14560 32386 14640 32400
rect 14560 32334 14574 32386
rect 14626 32334 14640 32386
rect 14560 32320 14640 32334
rect 14720 32386 14800 32400
rect 14720 32334 14734 32386
rect 14786 32334 14800 32386
rect 14720 32320 14800 32334
rect 14880 32386 14960 32400
rect 14880 32334 14894 32386
rect 14946 32334 14960 32386
rect 14880 32320 14960 32334
rect 15040 32386 15120 32400
rect 15040 32334 15054 32386
rect 15106 32334 15120 32386
rect 15040 32320 15120 32334
rect 15200 32386 15280 32400
rect 15200 32334 15214 32386
rect 15266 32334 15280 32386
rect 15200 32320 15280 32334
rect 15360 32386 15440 32400
rect 15360 32334 15374 32386
rect 15426 32334 15440 32386
rect 15360 32320 15440 32334
rect 15520 32386 15600 32400
rect 15520 32334 15534 32386
rect 15586 32334 15600 32386
rect 15520 32320 15600 32334
rect 15680 32386 15760 32400
rect 15680 32334 15694 32386
rect 15746 32334 15760 32386
rect 15680 32320 15760 32334
rect 15840 32386 15920 32400
rect 15840 32334 15854 32386
rect 15906 32334 15920 32386
rect 15840 32320 15920 32334
rect 16000 32386 16080 32400
rect 16000 32334 16014 32386
rect 16066 32334 16080 32386
rect 16000 32320 16080 32334
rect 16160 32386 16240 32400
rect 16160 32334 16174 32386
rect 16226 32334 16240 32386
rect 16160 32320 16240 32334
rect 16320 32386 16400 32400
rect 16320 32334 16334 32386
rect 16386 32334 16400 32386
rect 16320 32320 16400 32334
rect 16480 32386 16560 32400
rect 16480 32334 16494 32386
rect 16546 32334 16560 32386
rect 16480 32320 16560 32334
rect 16640 32386 16720 32400
rect 16640 32334 16654 32386
rect 16706 32334 16720 32386
rect 16640 32320 16720 32334
rect 16800 32386 16880 32400
rect 16800 32334 16814 32386
rect 16866 32334 16880 32386
rect 16800 32320 16880 32334
rect 16960 32386 17040 32400
rect 16960 32334 16974 32386
rect 17026 32334 17040 32386
rect 16960 32320 17040 32334
rect 17120 32386 17200 32400
rect 17120 32334 17134 32386
rect 17186 32334 17200 32386
rect 17120 32320 17200 32334
rect 17280 32386 17360 32400
rect 17280 32334 17294 32386
rect 17346 32334 17360 32386
rect 17280 32320 17360 32334
rect 17440 32386 17520 32400
rect 17440 32334 17454 32386
rect 17506 32334 17520 32386
rect 17440 32320 17520 32334
rect 17600 32386 17680 32400
rect 17600 32334 17614 32386
rect 17666 32334 17680 32386
rect 17600 32320 17680 32334
rect 17760 32386 17840 32400
rect 17760 32334 17774 32386
rect 17826 32334 17840 32386
rect 17760 32320 17840 32334
rect 17920 32386 18000 32400
rect 17920 32334 17934 32386
rect 17986 32334 18000 32386
rect 17920 32320 18000 32334
rect 18080 32386 18160 32400
rect 18080 32334 18094 32386
rect 18146 32334 18160 32386
rect 18080 32320 18160 32334
rect 18240 32386 18320 32400
rect 18240 32334 18254 32386
rect 18306 32334 18320 32386
rect 18240 32320 18320 32334
rect 18400 32386 18480 32400
rect 18400 32334 18414 32386
rect 18466 32334 18480 32386
rect 18400 32320 18480 32334
rect 18560 32386 18640 32400
rect 18560 32334 18574 32386
rect 18626 32334 18640 32386
rect 18560 32320 18640 32334
rect 18720 32386 18800 32400
rect 18720 32334 18734 32386
rect 18786 32334 18800 32386
rect 18720 32320 18800 32334
rect 18880 32386 18960 32400
rect 18880 32334 18894 32386
rect 18946 32334 18960 32386
rect 18880 32320 18960 32334
rect 23120 32386 23200 32400
rect 23120 32334 23134 32386
rect 23186 32334 23200 32386
rect 23120 32320 23200 32334
rect 23280 32386 23360 32400
rect 23280 32334 23294 32386
rect 23346 32334 23360 32386
rect 23280 32320 23360 32334
rect 23440 32386 23520 32400
rect 23440 32334 23454 32386
rect 23506 32334 23520 32386
rect 23440 32320 23520 32334
rect 23600 32386 23680 32400
rect 23600 32334 23614 32386
rect 23666 32334 23680 32386
rect 23600 32320 23680 32334
rect 23760 32386 23840 32400
rect 23760 32334 23774 32386
rect 23826 32334 23840 32386
rect 23760 32320 23840 32334
rect 23920 32386 24000 32400
rect 23920 32334 23934 32386
rect 23986 32334 24000 32386
rect 23920 32320 24000 32334
rect 24080 32386 24160 32400
rect 24080 32334 24094 32386
rect 24146 32334 24160 32386
rect 24080 32320 24160 32334
rect 24240 32386 24320 32400
rect 24240 32334 24254 32386
rect 24306 32334 24320 32386
rect 24240 32320 24320 32334
rect 24400 32386 24480 32400
rect 24400 32334 24414 32386
rect 24466 32334 24480 32386
rect 24400 32320 24480 32334
rect 24560 32386 24640 32400
rect 24560 32334 24574 32386
rect 24626 32334 24640 32386
rect 24560 32320 24640 32334
rect 24720 32386 24800 32400
rect 24720 32334 24734 32386
rect 24786 32334 24800 32386
rect 24720 32320 24800 32334
rect 24880 32386 24960 32400
rect 24880 32334 24894 32386
rect 24946 32334 24960 32386
rect 24880 32320 24960 32334
rect 25040 32386 25120 32400
rect 25040 32334 25054 32386
rect 25106 32334 25120 32386
rect 25040 32320 25120 32334
rect 25200 32386 25280 32400
rect 25200 32334 25214 32386
rect 25266 32334 25280 32386
rect 25200 32320 25280 32334
rect 25360 32386 25440 32400
rect 25360 32334 25374 32386
rect 25426 32334 25440 32386
rect 25360 32320 25440 32334
rect 25520 32386 25600 32400
rect 25520 32334 25534 32386
rect 25586 32334 25600 32386
rect 25520 32320 25600 32334
rect 25680 32386 25760 32400
rect 25680 32334 25694 32386
rect 25746 32334 25760 32386
rect 25680 32320 25760 32334
rect 25840 32386 25920 32400
rect 25840 32334 25854 32386
rect 25906 32334 25920 32386
rect 25840 32320 25920 32334
rect 26000 32386 26080 32400
rect 26000 32334 26014 32386
rect 26066 32334 26080 32386
rect 26000 32320 26080 32334
rect 26160 32386 26240 32400
rect 26160 32334 26174 32386
rect 26226 32334 26240 32386
rect 26160 32320 26240 32334
rect 26320 32386 26400 32400
rect 26320 32334 26334 32386
rect 26386 32334 26400 32386
rect 26320 32320 26400 32334
rect 26480 32386 26560 32400
rect 26480 32334 26494 32386
rect 26546 32334 26560 32386
rect 26480 32320 26560 32334
rect 26640 32386 26720 32400
rect 26640 32334 26654 32386
rect 26706 32334 26720 32386
rect 26640 32320 26720 32334
rect 26800 32386 26880 32400
rect 26800 32334 26814 32386
rect 26866 32334 26880 32386
rect 26800 32320 26880 32334
rect 26960 32386 27040 32400
rect 26960 32334 26974 32386
rect 27026 32334 27040 32386
rect 26960 32320 27040 32334
rect 27120 32386 27200 32400
rect 27120 32334 27134 32386
rect 27186 32334 27200 32386
rect 27120 32320 27200 32334
rect 27280 32386 27360 32400
rect 27280 32334 27294 32386
rect 27346 32334 27360 32386
rect 27280 32320 27360 32334
rect 27440 32386 27520 32400
rect 27440 32334 27454 32386
rect 27506 32334 27520 32386
rect 27440 32320 27520 32334
rect 27600 32386 27680 32400
rect 27600 32334 27614 32386
rect 27666 32334 27680 32386
rect 27600 32320 27680 32334
rect 27760 32386 27840 32400
rect 27760 32334 27774 32386
rect 27826 32334 27840 32386
rect 27760 32320 27840 32334
rect 27920 32386 28000 32400
rect 27920 32334 27934 32386
rect 27986 32334 28000 32386
rect 27920 32320 28000 32334
rect 28080 32386 28160 32400
rect 28080 32334 28094 32386
rect 28146 32334 28160 32386
rect 28080 32320 28160 32334
rect 28240 32386 28320 32400
rect 28240 32334 28254 32386
rect 28306 32334 28320 32386
rect 28240 32320 28320 32334
rect 28400 32386 28480 32400
rect 28400 32334 28414 32386
rect 28466 32334 28480 32386
rect 28400 32320 28480 32334
rect 28560 32386 28640 32400
rect 28560 32334 28574 32386
rect 28626 32334 28640 32386
rect 28560 32320 28640 32334
rect 28720 32386 28800 32400
rect 28720 32334 28734 32386
rect 28786 32334 28800 32386
rect 28720 32320 28800 32334
rect 28880 32386 28960 32400
rect 28880 32334 28894 32386
rect 28946 32334 28960 32386
rect 28880 32320 28960 32334
rect 29040 32386 29120 32400
rect 29040 32334 29054 32386
rect 29106 32334 29120 32386
rect 29040 32320 29120 32334
rect 29200 32386 29280 32400
rect 29200 32334 29214 32386
rect 29266 32334 29280 32386
rect 29200 32320 29280 32334
rect 29360 32386 29440 32400
rect 29360 32334 29374 32386
rect 29426 32334 29440 32386
rect 29360 32320 29440 32334
rect 33520 32386 33600 32400
rect 33520 32334 33534 32386
rect 33586 32334 33600 32386
rect 33520 32320 33600 32334
rect 33680 32386 33760 32400
rect 33680 32334 33694 32386
rect 33746 32334 33760 32386
rect 33680 32320 33760 32334
rect 33840 32386 33920 32400
rect 33840 32334 33854 32386
rect 33906 32334 33920 32386
rect 33840 32320 33920 32334
rect 34000 32386 34080 32400
rect 34000 32334 34014 32386
rect 34066 32334 34080 32386
rect 34000 32320 34080 32334
rect 34160 32386 34240 32400
rect 34160 32334 34174 32386
rect 34226 32334 34240 32386
rect 34160 32320 34240 32334
rect 34320 32386 34400 32400
rect 34320 32334 34334 32386
rect 34386 32334 34400 32386
rect 34320 32320 34400 32334
rect 34480 32386 34560 32400
rect 34480 32334 34494 32386
rect 34546 32334 34560 32386
rect 34480 32320 34560 32334
rect 34640 32386 34720 32400
rect 34640 32334 34654 32386
rect 34706 32334 34720 32386
rect 34640 32320 34720 32334
rect 34800 32386 34880 32400
rect 34800 32334 34814 32386
rect 34866 32334 34880 32386
rect 34800 32320 34880 32334
rect 34960 32386 35040 32400
rect 34960 32334 34974 32386
rect 35026 32334 35040 32386
rect 34960 32320 35040 32334
rect 35120 32386 35200 32400
rect 35120 32334 35134 32386
rect 35186 32334 35200 32386
rect 35120 32320 35200 32334
rect 35280 32386 35360 32400
rect 35280 32334 35294 32386
rect 35346 32334 35360 32386
rect 35280 32320 35360 32334
rect 35440 32386 35520 32400
rect 35440 32334 35454 32386
rect 35506 32334 35520 32386
rect 35440 32320 35520 32334
rect 35600 32386 35680 32400
rect 35600 32334 35614 32386
rect 35666 32334 35680 32386
rect 35600 32320 35680 32334
rect 35760 32386 35840 32400
rect 35760 32334 35774 32386
rect 35826 32334 35840 32386
rect 35760 32320 35840 32334
rect 35920 32386 36000 32400
rect 35920 32334 35934 32386
rect 35986 32334 36000 32386
rect 35920 32320 36000 32334
rect 36080 32386 36160 32400
rect 36080 32334 36094 32386
rect 36146 32334 36160 32386
rect 36080 32320 36160 32334
rect 36240 32386 36320 32400
rect 36240 32334 36254 32386
rect 36306 32334 36320 32386
rect 36240 32320 36320 32334
rect 36400 32386 36480 32400
rect 36400 32334 36414 32386
rect 36466 32334 36480 32386
rect 36400 32320 36480 32334
rect 36560 32386 36640 32400
rect 36560 32334 36574 32386
rect 36626 32334 36640 32386
rect 36560 32320 36640 32334
rect 36720 32386 36800 32400
rect 36720 32334 36734 32386
rect 36786 32334 36800 32386
rect 36720 32320 36800 32334
rect 36880 32386 36960 32400
rect 36880 32334 36894 32386
rect 36946 32334 36960 32386
rect 36880 32320 36960 32334
rect 37040 32386 37120 32400
rect 37040 32334 37054 32386
rect 37106 32334 37120 32386
rect 37040 32320 37120 32334
rect 37200 32386 37280 32400
rect 37200 32334 37214 32386
rect 37266 32334 37280 32386
rect 37200 32320 37280 32334
rect 37360 32386 37440 32400
rect 37360 32334 37374 32386
rect 37426 32334 37440 32386
rect 37360 32320 37440 32334
rect 37520 32386 37600 32400
rect 37520 32334 37534 32386
rect 37586 32334 37600 32386
rect 37520 32320 37600 32334
rect 37680 32386 37760 32400
rect 37680 32334 37694 32386
rect 37746 32334 37760 32386
rect 37680 32320 37760 32334
rect 37840 32386 37920 32400
rect 37840 32334 37854 32386
rect 37906 32334 37920 32386
rect 37840 32320 37920 32334
rect 38000 32386 38080 32400
rect 38000 32334 38014 32386
rect 38066 32334 38080 32386
rect 38000 32320 38080 32334
rect 38160 32386 38240 32400
rect 38160 32334 38174 32386
rect 38226 32334 38240 32386
rect 38160 32320 38240 32334
rect 38320 32386 38400 32400
rect 38320 32334 38334 32386
rect 38386 32334 38400 32386
rect 38320 32320 38400 32334
rect 38480 32386 38560 32400
rect 38480 32334 38494 32386
rect 38546 32334 38560 32386
rect 38480 32320 38560 32334
rect 38640 32386 38720 32400
rect 38640 32334 38654 32386
rect 38706 32334 38720 32386
rect 38640 32320 38720 32334
rect 38800 32386 38880 32400
rect 38800 32334 38814 32386
rect 38866 32334 38880 32386
rect 38800 32320 38880 32334
rect 38960 32386 39040 32400
rect 38960 32334 38974 32386
rect 39026 32334 39040 32386
rect 38960 32320 39040 32334
rect 39120 32386 39200 32400
rect 39120 32334 39134 32386
rect 39186 32334 39200 32386
rect 39120 32320 39200 32334
rect 39280 32386 39360 32400
rect 39280 32334 39294 32386
rect 39346 32334 39360 32386
rect 39280 32320 39360 32334
rect 39440 32386 39520 32400
rect 39440 32334 39454 32386
rect 39506 32334 39520 32386
rect 39440 32320 39520 32334
rect 39600 32386 39680 32400
rect 39600 32334 39614 32386
rect 39666 32334 39680 32386
rect 39600 32320 39680 32334
rect 39760 32386 39840 32400
rect 39760 32334 39774 32386
rect 39826 32334 39840 32386
rect 39760 32320 39840 32334
rect 39920 32386 40000 32400
rect 39920 32334 39934 32386
rect 39986 32334 40000 32386
rect 39920 32320 40000 32334
rect 40080 32386 40160 32400
rect 40080 32334 40094 32386
rect 40146 32334 40160 32386
rect 40080 32320 40160 32334
rect 40240 32386 40320 32400
rect 40240 32334 40254 32386
rect 40306 32334 40320 32386
rect 40240 32320 40320 32334
rect 40400 32386 40480 32400
rect 40400 32334 40414 32386
rect 40466 32334 40480 32386
rect 40400 32320 40480 32334
rect 40560 32386 40640 32400
rect 40560 32334 40574 32386
rect 40626 32334 40640 32386
rect 40560 32320 40640 32334
rect 40720 32386 40800 32400
rect 40720 32334 40734 32386
rect 40786 32334 40800 32386
rect 40720 32320 40800 32334
rect 40880 32386 40960 32400
rect 40880 32334 40894 32386
rect 40946 32334 40960 32386
rect 40880 32320 40960 32334
rect 41040 32386 41120 32400
rect 41040 32334 41054 32386
rect 41106 32334 41120 32386
rect 41040 32320 41120 32334
rect 41200 32386 41280 32400
rect 41200 32334 41214 32386
rect 41266 32334 41280 32386
rect 41200 32320 41280 32334
rect 41360 32386 41440 32400
rect 41360 32334 41374 32386
rect 41426 32334 41440 32386
rect 41360 32320 41440 32334
rect 41520 32386 41600 32400
rect 41520 32334 41534 32386
rect 41586 32334 41600 32386
rect 41520 32320 41600 32334
rect 41680 32386 41760 32400
rect 41680 32334 41694 32386
rect 41746 32334 41760 32386
rect 41680 32320 41760 32334
rect 41840 32386 41920 32400
rect 41840 32334 41854 32386
rect 41906 32334 41920 32386
rect 41840 32320 41920 32334
rect 0 32066 80 32080
rect 0 32014 14 32066
rect 66 32014 80 32066
rect 0 32000 80 32014
rect 160 32066 240 32080
rect 160 32014 174 32066
rect 226 32014 240 32066
rect 160 32000 240 32014
rect 320 32066 400 32080
rect 320 32014 334 32066
rect 386 32014 400 32066
rect 320 32000 400 32014
rect 480 32066 560 32080
rect 480 32014 494 32066
rect 546 32014 560 32066
rect 480 32000 560 32014
rect 640 32066 720 32080
rect 640 32014 654 32066
rect 706 32014 720 32066
rect 640 32000 720 32014
rect 800 32066 880 32080
rect 800 32014 814 32066
rect 866 32014 880 32066
rect 800 32000 880 32014
rect 960 32066 1040 32080
rect 960 32014 974 32066
rect 1026 32014 1040 32066
rect 960 32000 1040 32014
rect 1120 32066 1200 32080
rect 1120 32014 1134 32066
rect 1186 32014 1200 32066
rect 1120 32000 1200 32014
rect 1280 32066 1360 32080
rect 1280 32014 1294 32066
rect 1346 32014 1360 32066
rect 1280 32000 1360 32014
rect 1440 32066 1520 32080
rect 1440 32014 1454 32066
rect 1506 32014 1520 32066
rect 1440 32000 1520 32014
rect 1600 32066 1680 32080
rect 1600 32014 1614 32066
rect 1666 32014 1680 32066
rect 1600 32000 1680 32014
rect 1760 32066 1840 32080
rect 1760 32014 1774 32066
rect 1826 32014 1840 32066
rect 1760 32000 1840 32014
rect 1920 32066 2000 32080
rect 1920 32014 1934 32066
rect 1986 32014 2000 32066
rect 1920 32000 2000 32014
rect 2080 32066 2160 32080
rect 2080 32014 2094 32066
rect 2146 32014 2160 32066
rect 2080 32000 2160 32014
rect 2240 32066 2320 32080
rect 2240 32014 2254 32066
rect 2306 32014 2320 32066
rect 2240 32000 2320 32014
rect 2400 32066 2480 32080
rect 2400 32014 2414 32066
rect 2466 32014 2480 32066
rect 2400 32000 2480 32014
rect 2560 32066 2640 32080
rect 2560 32014 2574 32066
rect 2626 32014 2640 32066
rect 2560 32000 2640 32014
rect 2720 32066 2800 32080
rect 2720 32014 2734 32066
rect 2786 32014 2800 32066
rect 2720 32000 2800 32014
rect 2880 32066 2960 32080
rect 2880 32014 2894 32066
rect 2946 32014 2960 32066
rect 2880 32000 2960 32014
rect 3040 32066 3120 32080
rect 3040 32014 3054 32066
rect 3106 32014 3120 32066
rect 3040 32000 3120 32014
rect 3200 32066 3280 32080
rect 3200 32014 3214 32066
rect 3266 32014 3280 32066
rect 3200 32000 3280 32014
rect 3360 32066 3440 32080
rect 3360 32014 3374 32066
rect 3426 32014 3440 32066
rect 3360 32000 3440 32014
rect 3520 32066 3600 32080
rect 3520 32014 3534 32066
rect 3586 32014 3600 32066
rect 3520 32000 3600 32014
rect 3680 32066 3760 32080
rect 3680 32014 3694 32066
rect 3746 32014 3760 32066
rect 3680 32000 3760 32014
rect 3840 32066 3920 32080
rect 3840 32014 3854 32066
rect 3906 32014 3920 32066
rect 3840 32000 3920 32014
rect 4000 32066 4080 32080
rect 4000 32014 4014 32066
rect 4066 32014 4080 32066
rect 4000 32000 4080 32014
rect 4160 32066 4240 32080
rect 4160 32014 4174 32066
rect 4226 32014 4240 32066
rect 4160 32000 4240 32014
rect 4320 32066 4400 32080
rect 4320 32014 4334 32066
rect 4386 32014 4400 32066
rect 4320 32000 4400 32014
rect 4480 32066 4560 32080
rect 4480 32014 4494 32066
rect 4546 32014 4560 32066
rect 4480 32000 4560 32014
rect 4640 32066 4720 32080
rect 4640 32014 4654 32066
rect 4706 32014 4720 32066
rect 4640 32000 4720 32014
rect 4800 32066 4880 32080
rect 4800 32014 4814 32066
rect 4866 32014 4880 32066
rect 4800 32000 4880 32014
rect 4960 32066 5040 32080
rect 4960 32014 4974 32066
rect 5026 32014 5040 32066
rect 4960 32000 5040 32014
rect 5120 32066 5200 32080
rect 5120 32014 5134 32066
rect 5186 32014 5200 32066
rect 5120 32000 5200 32014
rect 5280 32066 5360 32080
rect 5280 32014 5294 32066
rect 5346 32014 5360 32066
rect 5280 32000 5360 32014
rect 5440 32066 5520 32080
rect 5440 32014 5454 32066
rect 5506 32014 5520 32066
rect 5440 32000 5520 32014
rect 5600 32066 5680 32080
rect 5600 32014 5614 32066
rect 5666 32014 5680 32066
rect 5600 32000 5680 32014
rect 5760 32066 5840 32080
rect 5760 32014 5774 32066
rect 5826 32014 5840 32066
rect 5760 32000 5840 32014
rect 5920 32066 6000 32080
rect 5920 32014 5934 32066
rect 5986 32014 6000 32066
rect 5920 32000 6000 32014
rect 6080 32066 6160 32080
rect 6080 32014 6094 32066
rect 6146 32014 6160 32066
rect 6080 32000 6160 32014
rect 6240 32066 6320 32080
rect 6240 32014 6254 32066
rect 6306 32014 6320 32066
rect 6240 32000 6320 32014
rect 6400 32066 6480 32080
rect 6400 32014 6414 32066
rect 6466 32014 6480 32066
rect 6400 32000 6480 32014
rect 6560 32066 6640 32080
rect 6560 32014 6574 32066
rect 6626 32014 6640 32066
rect 6560 32000 6640 32014
rect 6720 32066 6800 32080
rect 6720 32014 6734 32066
rect 6786 32014 6800 32066
rect 6720 32000 6800 32014
rect 6880 32066 6960 32080
rect 6880 32014 6894 32066
rect 6946 32014 6960 32066
rect 6880 32000 6960 32014
rect 7040 32066 7120 32080
rect 7040 32014 7054 32066
rect 7106 32014 7120 32066
rect 7040 32000 7120 32014
rect 7200 32066 7280 32080
rect 7200 32014 7214 32066
rect 7266 32014 7280 32066
rect 7200 32000 7280 32014
rect 7360 32066 7440 32080
rect 7360 32014 7374 32066
rect 7426 32014 7440 32066
rect 7360 32000 7440 32014
rect 7520 32066 7600 32080
rect 7520 32014 7534 32066
rect 7586 32014 7600 32066
rect 7520 32000 7600 32014
rect 7680 32066 7760 32080
rect 7680 32014 7694 32066
rect 7746 32014 7760 32066
rect 7680 32000 7760 32014
rect 7840 32066 7920 32080
rect 7840 32014 7854 32066
rect 7906 32014 7920 32066
rect 7840 32000 7920 32014
rect 8000 32066 8080 32080
rect 8000 32014 8014 32066
rect 8066 32014 8080 32066
rect 8000 32000 8080 32014
rect 8160 32066 8240 32080
rect 8160 32014 8174 32066
rect 8226 32014 8240 32066
rect 8160 32000 8240 32014
rect 8320 32066 8400 32080
rect 8320 32014 8334 32066
rect 8386 32014 8400 32066
rect 8320 32000 8400 32014
rect 12480 32066 12560 32080
rect 12480 32014 12494 32066
rect 12546 32014 12560 32066
rect 12480 32000 12560 32014
rect 12640 32066 12720 32080
rect 12640 32014 12654 32066
rect 12706 32014 12720 32066
rect 12640 32000 12720 32014
rect 12800 32066 12880 32080
rect 12800 32014 12814 32066
rect 12866 32014 12880 32066
rect 12800 32000 12880 32014
rect 12960 32066 13040 32080
rect 12960 32014 12974 32066
rect 13026 32014 13040 32066
rect 12960 32000 13040 32014
rect 13120 32066 13200 32080
rect 13120 32014 13134 32066
rect 13186 32014 13200 32066
rect 13120 32000 13200 32014
rect 13280 32066 13360 32080
rect 13280 32014 13294 32066
rect 13346 32014 13360 32066
rect 13280 32000 13360 32014
rect 13440 32066 13520 32080
rect 13440 32014 13454 32066
rect 13506 32014 13520 32066
rect 13440 32000 13520 32014
rect 13600 32066 13680 32080
rect 13600 32014 13614 32066
rect 13666 32014 13680 32066
rect 13600 32000 13680 32014
rect 13760 32066 13840 32080
rect 13760 32014 13774 32066
rect 13826 32014 13840 32066
rect 13760 32000 13840 32014
rect 13920 32066 14000 32080
rect 13920 32014 13934 32066
rect 13986 32014 14000 32066
rect 13920 32000 14000 32014
rect 14080 32066 14160 32080
rect 14080 32014 14094 32066
rect 14146 32014 14160 32066
rect 14080 32000 14160 32014
rect 14240 32066 14320 32080
rect 14240 32014 14254 32066
rect 14306 32014 14320 32066
rect 14240 32000 14320 32014
rect 14400 32066 14480 32080
rect 14400 32014 14414 32066
rect 14466 32014 14480 32066
rect 14400 32000 14480 32014
rect 14560 32066 14640 32080
rect 14560 32014 14574 32066
rect 14626 32014 14640 32066
rect 14560 32000 14640 32014
rect 14720 32066 14800 32080
rect 14720 32014 14734 32066
rect 14786 32014 14800 32066
rect 14720 32000 14800 32014
rect 14880 32066 14960 32080
rect 14880 32014 14894 32066
rect 14946 32014 14960 32066
rect 14880 32000 14960 32014
rect 15040 32066 15120 32080
rect 15040 32014 15054 32066
rect 15106 32014 15120 32066
rect 15040 32000 15120 32014
rect 15200 32066 15280 32080
rect 15200 32014 15214 32066
rect 15266 32014 15280 32066
rect 15200 32000 15280 32014
rect 15360 32066 15440 32080
rect 15360 32014 15374 32066
rect 15426 32014 15440 32066
rect 15360 32000 15440 32014
rect 15520 32066 15600 32080
rect 15520 32014 15534 32066
rect 15586 32014 15600 32066
rect 15520 32000 15600 32014
rect 15680 32066 15760 32080
rect 15680 32014 15694 32066
rect 15746 32014 15760 32066
rect 15680 32000 15760 32014
rect 15840 32066 15920 32080
rect 15840 32014 15854 32066
rect 15906 32014 15920 32066
rect 15840 32000 15920 32014
rect 16000 32066 16080 32080
rect 16000 32014 16014 32066
rect 16066 32014 16080 32066
rect 16000 32000 16080 32014
rect 16160 32066 16240 32080
rect 16160 32014 16174 32066
rect 16226 32014 16240 32066
rect 16160 32000 16240 32014
rect 16320 32066 16400 32080
rect 16320 32014 16334 32066
rect 16386 32014 16400 32066
rect 16320 32000 16400 32014
rect 16480 32066 16560 32080
rect 16480 32014 16494 32066
rect 16546 32014 16560 32066
rect 16480 32000 16560 32014
rect 16640 32066 16720 32080
rect 16640 32014 16654 32066
rect 16706 32014 16720 32066
rect 16640 32000 16720 32014
rect 16800 32066 16880 32080
rect 16800 32014 16814 32066
rect 16866 32014 16880 32066
rect 16800 32000 16880 32014
rect 16960 32066 17040 32080
rect 16960 32014 16974 32066
rect 17026 32014 17040 32066
rect 16960 32000 17040 32014
rect 17120 32066 17200 32080
rect 17120 32014 17134 32066
rect 17186 32014 17200 32066
rect 17120 32000 17200 32014
rect 17280 32066 17360 32080
rect 17280 32014 17294 32066
rect 17346 32014 17360 32066
rect 17280 32000 17360 32014
rect 17440 32066 17520 32080
rect 17440 32014 17454 32066
rect 17506 32014 17520 32066
rect 17440 32000 17520 32014
rect 17600 32066 17680 32080
rect 17600 32014 17614 32066
rect 17666 32014 17680 32066
rect 17600 32000 17680 32014
rect 17760 32066 17840 32080
rect 17760 32014 17774 32066
rect 17826 32014 17840 32066
rect 17760 32000 17840 32014
rect 17920 32066 18000 32080
rect 17920 32014 17934 32066
rect 17986 32014 18000 32066
rect 17920 32000 18000 32014
rect 18080 32066 18160 32080
rect 18080 32014 18094 32066
rect 18146 32014 18160 32066
rect 18080 32000 18160 32014
rect 18240 32066 18320 32080
rect 18240 32014 18254 32066
rect 18306 32014 18320 32066
rect 18240 32000 18320 32014
rect 18400 32066 18480 32080
rect 18400 32014 18414 32066
rect 18466 32014 18480 32066
rect 18400 32000 18480 32014
rect 18560 32066 18640 32080
rect 18560 32014 18574 32066
rect 18626 32014 18640 32066
rect 18560 32000 18640 32014
rect 18720 32066 18800 32080
rect 18720 32014 18734 32066
rect 18786 32014 18800 32066
rect 18720 32000 18800 32014
rect 18880 32066 18960 32080
rect 18880 32014 18894 32066
rect 18946 32014 18960 32066
rect 18880 32000 18960 32014
rect 23120 32066 23200 32080
rect 23120 32014 23134 32066
rect 23186 32014 23200 32066
rect 23120 32000 23200 32014
rect 23280 32066 23360 32080
rect 23280 32014 23294 32066
rect 23346 32014 23360 32066
rect 23280 32000 23360 32014
rect 23440 32066 23520 32080
rect 23440 32014 23454 32066
rect 23506 32014 23520 32066
rect 23440 32000 23520 32014
rect 23600 32066 23680 32080
rect 23600 32014 23614 32066
rect 23666 32014 23680 32066
rect 23600 32000 23680 32014
rect 23760 32066 23840 32080
rect 23760 32014 23774 32066
rect 23826 32014 23840 32066
rect 23760 32000 23840 32014
rect 23920 32066 24000 32080
rect 23920 32014 23934 32066
rect 23986 32014 24000 32066
rect 23920 32000 24000 32014
rect 24080 32066 24160 32080
rect 24080 32014 24094 32066
rect 24146 32014 24160 32066
rect 24080 32000 24160 32014
rect 24240 32066 24320 32080
rect 24240 32014 24254 32066
rect 24306 32014 24320 32066
rect 24240 32000 24320 32014
rect 24400 32066 24480 32080
rect 24400 32014 24414 32066
rect 24466 32014 24480 32066
rect 24400 32000 24480 32014
rect 24560 32066 24640 32080
rect 24560 32014 24574 32066
rect 24626 32014 24640 32066
rect 24560 32000 24640 32014
rect 24720 32066 24800 32080
rect 24720 32014 24734 32066
rect 24786 32014 24800 32066
rect 24720 32000 24800 32014
rect 24880 32066 24960 32080
rect 24880 32014 24894 32066
rect 24946 32014 24960 32066
rect 24880 32000 24960 32014
rect 25040 32066 25120 32080
rect 25040 32014 25054 32066
rect 25106 32014 25120 32066
rect 25040 32000 25120 32014
rect 25200 32066 25280 32080
rect 25200 32014 25214 32066
rect 25266 32014 25280 32066
rect 25200 32000 25280 32014
rect 25360 32066 25440 32080
rect 25360 32014 25374 32066
rect 25426 32014 25440 32066
rect 25360 32000 25440 32014
rect 25520 32066 25600 32080
rect 25520 32014 25534 32066
rect 25586 32014 25600 32066
rect 25520 32000 25600 32014
rect 25680 32066 25760 32080
rect 25680 32014 25694 32066
rect 25746 32014 25760 32066
rect 25680 32000 25760 32014
rect 25840 32066 25920 32080
rect 25840 32014 25854 32066
rect 25906 32014 25920 32066
rect 25840 32000 25920 32014
rect 26000 32066 26080 32080
rect 26000 32014 26014 32066
rect 26066 32014 26080 32066
rect 26000 32000 26080 32014
rect 26160 32066 26240 32080
rect 26160 32014 26174 32066
rect 26226 32014 26240 32066
rect 26160 32000 26240 32014
rect 26320 32066 26400 32080
rect 26320 32014 26334 32066
rect 26386 32014 26400 32066
rect 26320 32000 26400 32014
rect 26480 32066 26560 32080
rect 26480 32014 26494 32066
rect 26546 32014 26560 32066
rect 26480 32000 26560 32014
rect 26640 32066 26720 32080
rect 26640 32014 26654 32066
rect 26706 32014 26720 32066
rect 26640 32000 26720 32014
rect 26800 32066 26880 32080
rect 26800 32014 26814 32066
rect 26866 32014 26880 32066
rect 26800 32000 26880 32014
rect 26960 32066 27040 32080
rect 26960 32014 26974 32066
rect 27026 32014 27040 32066
rect 26960 32000 27040 32014
rect 27120 32066 27200 32080
rect 27120 32014 27134 32066
rect 27186 32014 27200 32066
rect 27120 32000 27200 32014
rect 27280 32066 27360 32080
rect 27280 32014 27294 32066
rect 27346 32014 27360 32066
rect 27280 32000 27360 32014
rect 27440 32066 27520 32080
rect 27440 32014 27454 32066
rect 27506 32014 27520 32066
rect 27440 32000 27520 32014
rect 27600 32066 27680 32080
rect 27600 32014 27614 32066
rect 27666 32014 27680 32066
rect 27600 32000 27680 32014
rect 27760 32066 27840 32080
rect 27760 32014 27774 32066
rect 27826 32014 27840 32066
rect 27760 32000 27840 32014
rect 27920 32066 28000 32080
rect 27920 32014 27934 32066
rect 27986 32014 28000 32066
rect 27920 32000 28000 32014
rect 28080 32066 28160 32080
rect 28080 32014 28094 32066
rect 28146 32014 28160 32066
rect 28080 32000 28160 32014
rect 28240 32066 28320 32080
rect 28240 32014 28254 32066
rect 28306 32014 28320 32066
rect 28240 32000 28320 32014
rect 28400 32066 28480 32080
rect 28400 32014 28414 32066
rect 28466 32014 28480 32066
rect 28400 32000 28480 32014
rect 28560 32066 28640 32080
rect 28560 32014 28574 32066
rect 28626 32014 28640 32066
rect 28560 32000 28640 32014
rect 28720 32066 28800 32080
rect 28720 32014 28734 32066
rect 28786 32014 28800 32066
rect 28720 32000 28800 32014
rect 28880 32066 28960 32080
rect 28880 32014 28894 32066
rect 28946 32014 28960 32066
rect 28880 32000 28960 32014
rect 29040 32066 29120 32080
rect 29040 32014 29054 32066
rect 29106 32014 29120 32066
rect 29040 32000 29120 32014
rect 29200 32066 29280 32080
rect 29200 32014 29214 32066
rect 29266 32014 29280 32066
rect 29200 32000 29280 32014
rect 29360 32066 29440 32080
rect 29360 32014 29374 32066
rect 29426 32014 29440 32066
rect 29360 32000 29440 32014
rect 33520 32066 33600 32080
rect 33520 32014 33534 32066
rect 33586 32014 33600 32066
rect 33520 32000 33600 32014
rect 33680 32066 33760 32080
rect 33680 32014 33694 32066
rect 33746 32014 33760 32066
rect 33680 32000 33760 32014
rect 33840 32066 33920 32080
rect 33840 32014 33854 32066
rect 33906 32014 33920 32066
rect 33840 32000 33920 32014
rect 34000 32066 34080 32080
rect 34000 32014 34014 32066
rect 34066 32014 34080 32066
rect 34000 32000 34080 32014
rect 34160 32066 34240 32080
rect 34160 32014 34174 32066
rect 34226 32014 34240 32066
rect 34160 32000 34240 32014
rect 34320 32066 34400 32080
rect 34320 32014 34334 32066
rect 34386 32014 34400 32066
rect 34320 32000 34400 32014
rect 34480 32066 34560 32080
rect 34480 32014 34494 32066
rect 34546 32014 34560 32066
rect 34480 32000 34560 32014
rect 34640 32066 34720 32080
rect 34640 32014 34654 32066
rect 34706 32014 34720 32066
rect 34640 32000 34720 32014
rect 34800 32066 34880 32080
rect 34800 32014 34814 32066
rect 34866 32014 34880 32066
rect 34800 32000 34880 32014
rect 34960 32066 35040 32080
rect 34960 32014 34974 32066
rect 35026 32014 35040 32066
rect 34960 32000 35040 32014
rect 35120 32066 35200 32080
rect 35120 32014 35134 32066
rect 35186 32014 35200 32066
rect 35120 32000 35200 32014
rect 35280 32066 35360 32080
rect 35280 32014 35294 32066
rect 35346 32014 35360 32066
rect 35280 32000 35360 32014
rect 35440 32066 35520 32080
rect 35440 32014 35454 32066
rect 35506 32014 35520 32066
rect 35440 32000 35520 32014
rect 35600 32066 35680 32080
rect 35600 32014 35614 32066
rect 35666 32014 35680 32066
rect 35600 32000 35680 32014
rect 35760 32066 35840 32080
rect 35760 32014 35774 32066
rect 35826 32014 35840 32066
rect 35760 32000 35840 32014
rect 35920 32066 36000 32080
rect 35920 32014 35934 32066
rect 35986 32014 36000 32066
rect 35920 32000 36000 32014
rect 36080 32066 36160 32080
rect 36080 32014 36094 32066
rect 36146 32014 36160 32066
rect 36080 32000 36160 32014
rect 36240 32066 36320 32080
rect 36240 32014 36254 32066
rect 36306 32014 36320 32066
rect 36240 32000 36320 32014
rect 36400 32066 36480 32080
rect 36400 32014 36414 32066
rect 36466 32014 36480 32066
rect 36400 32000 36480 32014
rect 36560 32066 36640 32080
rect 36560 32014 36574 32066
rect 36626 32014 36640 32066
rect 36560 32000 36640 32014
rect 36720 32066 36800 32080
rect 36720 32014 36734 32066
rect 36786 32014 36800 32066
rect 36720 32000 36800 32014
rect 36880 32066 36960 32080
rect 36880 32014 36894 32066
rect 36946 32014 36960 32066
rect 36880 32000 36960 32014
rect 37040 32066 37120 32080
rect 37040 32014 37054 32066
rect 37106 32014 37120 32066
rect 37040 32000 37120 32014
rect 37200 32066 37280 32080
rect 37200 32014 37214 32066
rect 37266 32014 37280 32066
rect 37200 32000 37280 32014
rect 37360 32066 37440 32080
rect 37360 32014 37374 32066
rect 37426 32014 37440 32066
rect 37360 32000 37440 32014
rect 37520 32066 37600 32080
rect 37520 32014 37534 32066
rect 37586 32014 37600 32066
rect 37520 32000 37600 32014
rect 37680 32066 37760 32080
rect 37680 32014 37694 32066
rect 37746 32014 37760 32066
rect 37680 32000 37760 32014
rect 37840 32066 37920 32080
rect 37840 32014 37854 32066
rect 37906 32014 37920 32066
rect 37840 32000 37920 32014
rect 38000 32066 38080 32080
rect 38000 32014 38014 32066
rect 38066 32014 38080 32066
rect 38000 32000 38080 32014
rect 38160 32066 38240 32080
rect 38160 32014 38174 32066
rect 38226 32014 38240 32066
rect 38160 32000 38240 32014
rect 38320 32066 38400 32080
rect 38320 32014 38334 32066
rect 38386 32014 38400 32066
rect 38320 32000 38400 32014
rect 38480 32066 38560 32080
rect 38480 32014 38494 32066
rect 38546 32014 38560 32066
rect 38480 32000 38560 32014
rect 38640 32066 38720 32080
rect 38640 32014 38654 32066
rect 38706 32014 38720 32066
rect 38640 32000 38720 32014
rect 38800 32066 38880 32080
rect 38800 32014 38814 32066
rect 38866 32014 38880 32066
rect 38800 32000 38880 32014
rect 38960 32066 39040 32080
rect 38960 32014 38974 32066
rect 39026 32014 39040 32066
rect 38960 32000 39040 32014
rect 39120 32066 39200 32080
rect 39120 32014 39134 32066
rect 39186 32014 39200 32066
rect 39120 32000 39200 32014
rect 39280 32066 39360 32080
rect 39280 32014 39294 32066
rect 39346 32014 39360 32066
rect 39280 32000 39360 32014
rect 39440 32066 39520 32080
rect 39440 32014 39454 32066
rect 39506 32014 39520 32066
rect 39440 32000 39520 32014
rect 39600 32066 39680 32080
rect 39600 32014 39614 32066
rect 39666 32014 39680 32066
rect 39600 32000 39680 32014
rect 39760 32066 39840 32080
rect 39760 32014 39774 32066
rect 39826 32014 39840 32066
rect 39760 32000 39840 32014
rect 39920 32066 40000 32080
rect 39920 32014 39934 32066
rect 39986 32014 40000 32066
rect 39920 32000 40000 32014
rect 40080 32066 40160 32080
rect 40080 32014 40094 32066
rect 40146 32014 40160 32066
rect 40080 32000 40160 32014
rect 40240 32066 40320 32080
rect 40240 32014 40254 32066
rect 40306 32014 40320 32066
rect 40240 32000 40320 32014
rect 40400 32066 40480 32080
rect 40400 32014 40414 32066
rect 40466 32014 40480 32066
rect 40400 32000 40480 32014
rect 40560 32066 40640 32080
rect 40560 32014 40574 32066
rect 40626 32014 40640 32066
rect 40560 32000 40640 32014
rect 40720 32066 40800 32080
rect 40720 32014 40734 32066
rect 40786 32014 40800 32066
rect 40720 32000 40800 32014
rect 40880 32066 40960 32080
rect 40880 32014 40894 32066
rect 40946 32014 40960 32066
rect 40880 32000 40960 32014
rect 41040 32066 41120 32080
rect 41040 32014 41054 32066
rect 41106 32014 41120 32066
rect 41040 32000 41120 32014
rect 41200 32066 41280 32080
rect 41200 32014 41214 32066
rect 41266 32014 41280 32066
rect 41200 32000 41280 32014
rect 41360 32066 41440 32080
rect 41360 32014 41374 32066
rect 41426 32014 41440 32066
rect 41360 32000 41440 32014
rect 41520 32066 41600 32080
rect 41520 32014 41534 32066
rect 41586 32014 41600 32066
rect 41520 32000 41600 32014
rect 41680 32066 41760 32080
rect 41680 32014 41694 32066
rect 41746 32014 41760 32066
rect 41680 32000 41760 32014
rect 41840 32066 41920 32080
rect 41840 32014 41854 32066
rect 41906 32014 41920 32066
rect 41840 32000 41920 32014
rect 0 31746 80 31760
rect 0 31694 14 31746
rect 66 31694 80 31746
rect 0 31680 80 31694
rect 160 31746 240 31760
rect 160 31694 174 31746
rect 226 31694 240 31746
rect 160 31680 240 31694
rect 320 31746 400 31760
rect 320 31694 334 31746
rect 386 31694 400 31746
rect 320 31680 400 31694
rect 480 31746 560 31760
rect 480 31694 494 31746
rect 546 31694 560 31746
rect 480 31680 560 31694
rect 640 31746 720 31760
rect 640 31694 654 31746
rect 706 31694 720 31746
rect 640 31680 720 31694
rect 800 31746 880 31760
rect 800 31694 814 31746
rect 866 31694 880 31746
rect 800 31680 880 31694
rect 960 31746 1040 31760
rect 960 31694 974 31746
rect 1026 31694 1040 31746
rect 960 31680 1040 31694
rect 1120 31746 1200 31760
rect 1120 31694 1134 31746
rect 1186 31694 1200 31746
rect 1120 31680 1200 31694
rect 1280 31746 1360 31760
rect 1280 31694 1294 31746
rect 1346 31694 1360 31746
rect 1280 31680 1360 31694
rect 1440 31746 1520 31760
rect 1440 31694 1454 31746
rect 1506 31694 1520 31746
rect 1440 31680 1520 31694
rect 1600 31746 1680 31760
rect 1600 31694 1614 31746
rect 1666 31694 1680 31746
rect 1600 31680 1680 31694
rect 1760 31746 1840 31760
rect 1760 31694 1774 31746
rect 1826 31694 1840 31746
rect 1760 31680 1840 31694
rect 1920 31746 2000 31760
rect 1920 31694 1934 31746
rect 1986 31694 2000 31746
rect 1920 31680 2000 31694
rect 2080 31746 2160 31760
rect 2080 31694 2094 31746
rect 2146 31694 2160 31746
rect 2080 31680 2160 31694
rect 2240 31746 2320 31760
rect 2240 31694 2254 31746
rect 2306 31694 2320 31746
rect 2240 31680 2320 31694
rect 2400 31746 2480 31760
rect 2400 31694 2414 31746
rect 2466 31694 2480 31746
rect 2400 31680 2480 31694
rect 2560 31746 2640 31760
rect 2560 31694 2574 31746
rect 2626 31694 2640 31746
rect 2560 31680 2640 31694
rect 2720 31746 2800 31760
rect 2720 31694 2734 31746
rect 2786 31694 2800 31746
rect 2720 31680 2800 31694
rect 2880 31746 2960 31760
rect 2880 31694 2894 31746
rect 2946 31694 2960 31746
rect 2880 31680 2960 31694
rect 3040 31746 3120 31760
rect 3040 31694 3054 31746
rect 3106 31694 3120 31746
rect 3040 31680 3120 31694
rect 3200 31746 3280 31760
rect 3200 31694 3214 31746
rect 3266 31694 3280 31746
rect 3200 31680 3280 31694
rect 3360 31746 3440 31760
rect 3360 31694 3374 31746
rect 3426 31694 3440 31746
rect 3360 31680 3440 31694
rect 3520 31746 3600 31760
rect 3520 31694 3534 31746
rect 3586 31694 3600 31746
rect 3520 31680 3600 31694
rect 3680 31746 3760 31760
rect 3680 31694 3694 31746
rect 3746 31694 3760 31746
rect 3680 31680 3760 31694
rect 3840 31746 3920 31760
rect 3840 31694 3854 31746
rect 3906 31694 3920 31746
rect 3840 31680 3920 31694
rect 4000 31746 4080 31760
rect 4000 31694 4014 31746
rect 4066 31694 4080 31746
rect 4000 31680 4080 31694
rect 4160 31746 4240 31760
rect 4160 31694 4174 31746
rect 4226 31694 4240 31746
rect 4160 31680 4240 31694
rect 4320 31746 4400 31760
rect 4320 31694 4334 31746
rect 4386 31694 4400 31746
rect 4320 31680 4400 31694
rect 4480 31746 4560 31760
rect 4480 31694 4494 31746
rect 4546 31694 4560 31746
rect 4480 31680 4560 31694
rect 4640 31746 4720 31760
rect 4640 31694 4654 31746
rect 4706 31694 4720 31746
rect 4640 31680 4720 31694
rect 4800 31746 4880 31760
rect 4800 31694 4814 31746
rect 4866 31694 4880 31746
rect 4800 31680 4880 31694
rect 4960 31746 5040 31760
rect 4960 31694 4974 31746
rect 5026 31694 5040 31746
rect 4960 31680 5040 31694
rect 5120 31746 5200 31760
rect 5120 31694 5134 31746
rect 5186 31694 5200 31746
rect 5120 31680 5200 31694
rect 5280 31746 5360 31760
rect 5280 31694 5294 31746
rect 5346 31694 5360 31746
rect 5280 31680 5360 31694
rect 5440 31746 5520 31760
rect 5440 31694 5454 31746
rect 5506 31694 5520 31746
rect 5440 31680 5520 31694
rect 5600 31746 5680 31760
rect 5600 31694 5614 31746
rect 5666 31694 5680 31746
rect 5600 31680 5680 31694
rect 5760 31746 5840 31760
rect 5760 31694 5774 31746
rect 5826 31694 5840 31746
rect 5760 31680 5840 31694
rect 5920 31746 6000 31760
rect 5920 31694 5934 31746
rect 5986 31694 6000 31746
rect 5920 31680 6000 31694
rect 6080 31746 6160 31760
rect 6080 31694 6094 31746
rect 6146 31694 6160 31746
rect 6080 31680 6160 31694
rect 6240 31746 6320 31760
rect 6240 31694 6254 31746
rect 6306 31694 6320 31746
rect 6240 31680 6320 31694
rect 6400 31746 6480 31760
rect 6400 31694 6414 31746
rect 6466 31694 6480 31746
rect 6400 31680 6480 31694
rect 6560 31746 6640 31760
rect 6560 31694 6574 31746
rect 6626 31694 6640 31746
rect 6560 31680 6640 31694
rect 6720 31746 6800 31760
rect 6720 31694 6734 31746
rect 6786 31694 6800 31746
rect 6720 31680 6800 31694
rect 6880 31746 6960 31760
rect 6880 31694 6894 31746
rect 6946 31694 6960 31746
rect 6880 31680 6960 31694
rect 7040 31746 7120 31760
rect 7040 31694 7054 31746
rect 7106 31694 7120 31746
rect 7040 31680 7120 31694
rect 7200 31746 7280 31760
rect 7200 31694 7214 31746
rect 7266 31694 7280 31746
rect 7200 31680 7280 31694
rect 7360 31746 7440 31760
rect 7360 31694 7374 31746
rect 7426 31694 7440 31746
rect 7360 31680 7440 31694
rect 7520 31746 7600 31760
rect 7520 31694 7534 31746
rect 7586 31694 7600 31746
rect 7520 31680 7600 31694
rect 7680 31746 7760 31760
rect 7680 31694 7694 31746
rect 7746 31694 7760 31746
rect 7680 31680 7760 31694
rect 7840 31746 7920 31760
rect 7840 31694 7854 31746
rect 7906 31694 7920 31746
rect 7840 31680 7920 31694
rect 8000 31746 8080 31760
rect 8000 31694 8014 31746
rect 8066 31694 8080 31746
rect 8000 31680 8080 31694
rect 8160 31746 8240 31760
rect 8160 31694 8174 31746
rect 8226 31694 8240 31746
rect 8160 31680 8240 31694
rect 8320 31746 8400 31760
rect 8320 31694 8334 31746
rect 8386 31694 8400 31746
rect 8320 31680 8400 31694
rect 12480 31746 12560 31760
rect 12480 31694 12494 31746
rect 12546 31694 12560 31746
rect 12480 31680 12560 31694
rect 12640 31746 12720 31760
rect 12640 31694 12654 31746
rect 12706 31694 12720 31746
rect 12640 31680 12720 31694
rect 12800 31746 12880 31760
rect 12800 31694 12814 31746
rect 12866 31694 12880 31746
rect 12800 31680 12880 31694
rect 12960 31746 13040 31760
rect 12960 31694 12974 31746
rect 13026 31694 13040 31746
rect 12960 31680 13040 31694
rect 13120 31746 13200 31760
rect 13120 31694 13134 31746
rect 13186 31694 13200 31746
rect 13120 31680 13200 31694
rect 13280 31746 13360 31760
rect 13280 31694 13294 31746
rect 13346 31694 13360 31746
rect 13280 31680 13360 31694
rect 13440 31746 13520 31760
rect 13440 31694 13454 31746
rect 13506 31694 13520 31746
rect 13440 31680 13520 31694
rect 13600 31746 13680 31760
rect 13600 31694 13614 31746
rect 13666 31694 13680 31746
rect 13600 31680 13680 31694
rect 13760 31746 13840 31760
rect 13760 31694 13774 31746
rect 13826 31694 13840 31746
rect 13760 31680 13840 31694
rect 13920 31746 14000 31760
rect 13920 31694 13934 31746
rect 13986 31694 14000 31746
rect 13920 31680 14000 31694
rect 14080 31746 14160 31760
rect 14080 31694 14094 31746
rect 14146 31694 14160 31746
rect 14080 31680 14160 31694
rect 14240 31746 14320 31760
rect 14240 31694 14254 31746
rect 14306 31694 14320 31746
rect 14240 31680 14320 31694
rect 14400 31746 14480 31760
rect 14400 31694 14414 31746
rect 14466 31694 14480 31746
rect 14400 31680 14480 31694
rect 14560 31746 14640 31760
rect 14560 31694 14574 31746
rect 14626 31694 14640 31746
rect 14560 31680 14640 31694
rect 14720 31746 14800 31760
rect 14720 31694 14734 31746
rect 14786 31694 14800 31746
rect 14720 31680 14800 31694
rect 14880 31746 14960 31760
rect 14880 31694 14894 31746
rect 14946 31694 14960 31746
rect 14880 31680 14960 31694
rect 15040 31746 15120 31760
rect 15040 31694 15054 31746
rect 15106 31694 15120 31746
rect 15040 31680 15120 31694
rect 15200 31746 15280 31760
rect 15200 31694 15214 31746
rect 15266 31694 15280 31746
rect 15200 31680 15280 31694
rect 15360 31746 15440 31760
rect 15360 31694 15374 31746
rect 15426 31694 15440 31746
rect 15360 31680 15440 31694
rect 15520 31746 15600 31760
rect 15520 31694 15534 31746
rect 15586 31694 15600 31746
rect 15520 31680 15600 31694
rect 15680 31746 15760 31760
rect 15680 31694 15694 31746
rect 15746 31694 15760 31746
rect 15680 31680 15760 31694
rect 15840 31746 15920 31760
rect 15840 31694 15854 31746
rect 15906 31694 15920 31746
rect 15840 31680 15920 31694
rect 16000 31746 16080 31760
rect 16000 31694 16014 31746
rect 16066 31694 16080 31746
rect 16000 31680 16080 31694
rect 16160 31746 16240 31760
rect 16160 31694 16174 31746
rect 16226 31694 16240 31746
rect 16160 31680 16240 31694
rect 16320 31746 16400 31760
rect 16320 31694 16334 31746
rect 16386 31694 16400 31746
rect 16320 31680 16400 31694
rect 16480 31746 16560 31760
rect 16480 31694 16494 31746
rect 16546 31694 16560 31746
rect 16480 31680 16560 31694
rect 16640 31746 16720 31760
rect 16640 31694 16654 31746
rect 16706 31694 16720 31746
rect 16640 31680 16720 31694
rect 16800 31746 16880 31760
rect 16800 31694 16814 31746
rect 16866 31694 16880 31746
rect 16800 31680 16880 31694
rect 16960 31746 17040 31760
rect 16960 31694 16974 31746
rect 17026 31694 17040 31746
rect 16960 31680 17040 31694
rect 17120 31746 17200 31760
rect 17120 31694 17134 31746
rect 17186 31694 17200 31746
rect 17120 31680 17200 31694
rect 17280 31746 17360 31760
rect 17280 31694 17294 31746
rect 17346 31694 17360 31746
rect 17280 31680 17360 31694
rect 17440 31746 17520 31760
rect 17440 31694 17454 31746
rect 17506 31694 17520 31746
rect 17440 31680 17520 31694
rect 17600 31746 17680 31760
rect 17600 31694 17614 31746
rect 17666 31694 17680 31746
rect 17600 31680 17680 31694
rect 17760 31746 17840 31760
rect 17760 31694 17774 31746
rect 17826 31694 17840 31746
rect 17760 31680 17840 31694
rect 17920 31746 18000 31760
rect 17920 31694 17934 31746
rect 17986 31694 18000 31746
rect 17920 31680 18000 31694
rect 18080 31746 18160 31760
rect 18080 31694 18094 31746
rect 18146 31694 18160 31746
rect 18080 31680 18160 31694
rect 18240 31746 18320 31760
rect 18240 31694 18254 31746
rect 18306 31694 18320 31746
rect 18240 31680 18320 31694
rect 18400 31746 18480 31760
rect 18400 31694 18414 31746
rect 18466 31694 18480 31746
rect 18400 31680 18480 31694
rect 18560 31746 18640 31760
rect 18560 31694 18574 31746
rect 18626 31694 18640 31746
rect 18560 31680 18640 31694
rect 18720 31746 18800 31760
rect 18720 31694 18734 31746
rect 18786 31694 18800 31746
rect 18720 31680 18800 31694
rect 18880 31746 18960 31760
rect 18880 31694 18894 31746
rect 18946 31694 18960 31746
rect 18880 31680 18960 31694
rect 23120 31746 23200 31760
rect 23120 31694 23134 31746
rect 23186 31694 23200 31746
rect 23120 31680 23200 31694
rect 23280 31746 23360 31760
rect 23280 31694 23294 31746
rect 23346 31694 23360 31746
rect 23280 31680 23360 31694
rect 23440 31746 23520 31760
rect 23440 31694 23454 31746
rect 23506 31694 23520 31746
rect 23440 31680 23520 31694
rect 23600 31746 23680 31760
rect 23600 31694 23614 31746
rect 23666 31694 23680 31746
rect 23600 31680 23680 31694
rect 23760 31746 23840 31760
rect 23760 31694 23774 31746
rect 23826 31694 23840 31746
rect 23760 31680 23840 31694
rect 23920 31746 24000 31760
rect 23920 31694 23934 31746
rect 23986 31694 24000 31746
rect 23920 31680 24000 31694
rect 24080 31746 24160 31760
rect 24080 31694 24094 31746
rect 24146 31694 24160 31746
rect 24080 31680 24160 31694
rect 24240 31746 24320 31760
rect 24240 31694 24254 31746
rect 24306 31694 24320 31746
rect 24240 31680 24320 31694
rect 24400 31746 24480 31760
rect 24400 31694 24414 31746
rect 24466 31694 24480 31746
rect 24400 31680 24480 31694
rect 24560 31746 24640 31760
rect 24560 31694 24574 31746
rect 24626 31694 24640 31746
rect 24560 31680 24640 31694
rect 24720 31746 24800 31760
rect 24720 31694 24734 31746
rect 24786 31694 24800 31746
rect 24720 31680 24800 31694
rect 24880 31746 24960 31760
rect 24880 31694 24894 31746
rect 24946 31694 24960 31746
rect 24880 31680 24960 31694
rect 25040 31746 25120 31760
rect 25040 31694 25054 31746
rect 25106 31694 25120 31746
rect 25040 31680 25120 31694
rect 25200 31746 25280 31760
rect 25200 31694 25214 31746
rect 25266 31694 25280 31746
rect 25200 31680 25280 31694
rect 25360 31746 25440 31760
rect 25360 31694 25374 31746
rect 25426 31694 25440 31746
rect 25360 31680 25440 31694
rect 25520 31746 25600 31760
rect 25520 31694 25534 31746
rect 25586 31694 25600 31746
rect 25520 31680 25600 31694
rect 25680 31746 25760 31760
rect 25680 31694 25694 31746
rect 25746 31694 25760 31746
rect 25680 31680 25760 31694
rect 25840 31746 25920 31760
rect 25840 31694 25854 31746
rect 25906 31694 25920 31746
rect 25840 31680 25920 31694
rect 26000 31746 26080 31760
rect 26000 31694 26014 31746
rect 26066 31694 26080 31746
rect 26000 31680 26080 31694
rect 26160 31746 26240 31760
rect 26160 31694 26174 31746
rect 26226 31694 26240 31746
rect 26160 31680 26240 31694
rect 26320 31746 26400 31760
rect 26320 31694 26334 31746
rect 26386 31694 26400 31746
rect 26320 31680 26400 31694
rect 26480 31746 26560 31760
rect 26480 31694 26494 31746
rect 26546 31694 26560 31746
rect 26480 31680 26560 31694
rect 26640 31746 26720 31760
rect 26640 31694 26654 31746
rect 26706 31694 26720 31746
rect 26640 31680 26720 31694
rect 26800 31746 26880 31760
rect 26800 31694 26814 31746
rect 26866 31694 26880 31746
rect 26800 31680 26880 31694
rect 26960 31746 27040 31760
rect 26960 31694 26974 31746
rect 27026 31694 27040 31746
rect 26960 31680 27040 31694
rect 27120 31746 27200 31760
rect 27120 31694 27134 31746
rect 27186 31694 27200 31746
rect 27120 31680 27200 31694
rect 27280 31746 27360 31760
rect 27280 31694 27294 31746
rect 27346 31694 27360 31746
rect 27280 31680 27360 31694
rect 27440 31746 27520 31760
rect 27440 31694 27454 31746
rect 27506 31694 27520 31746
rect 27440 31680 27520 31694
rect 27600 31746 27680 31760
rect 27600 31694 27614 31746
rect 27666 31694 27680 31746
rect 27600 31680 27680 31694
rect 27760 31746 27840 31760
rect 27760 31694 27774 31746
rect 27826 31694 27840 31746
rect 27760 31680 27840 31694
rect 27920 31746 28000 31760
rect 27920 31694 27934 31746
rect 27986 31694 28000 31746
rect 27920 31680 28000 31694
rect 28080 31746 28160 31760
rect 28080 31694 28094 31746
rect 28146 31694 28160 31746
rect 28080 31680 28160 31694
rect 28240 31746 28320 31760
rect 28240 31694 28254 31746
rect 28306 31694 28320 31746
rect 28240 31680 28320 31694
rect 28400 31746 28480 31760
rect 28400 31694 28414 31746
rect 28466 31694 28480 31746
rect 28400 31680 28480 31694
rect 28560 31746 28640 31760
rect 28560 31694 28574 31746
rect 28626 31694 28640 31746
rect 28560 31680 28640 31694
rect 28720 31746 28800 31760
rect 28720 31694 28734 31746
rect 28786 31694 28800 31746
rect 28720 31680 28800 31694
rect 28880 31746 28960 31760
rect 28880 31694 28894 31746
rect 28946 31694 28960 31746
rect 28880 31680 28960 31694
rect 29040 31746 29120 31760
rect 29040 31694 29054 31746
rect 29106 31694 29120 31746
rect 29040 31680 29120 31694
rect 29200 31746 29280 31760
rect 29200 31694 29214 31746
rect 29266 31694 29280 31746
rect 29200 31680 29280 31694
rect 29360 31746 29440 31760
rect 29360 31694 29374 31746
rect 29426 31694 29440 31746
rect 29360 31680 29440 31694
rect 33520 31746 33600 31760
rect 33520 31694 33534 31746
rect 33586 31694 33600 31746
rect 33520 31680 33600 31694
rect 33680 31746 33760 31760
rect 33680 31694 33694 31746
rect 33746 31694 33760 31746
rect 33680 31680 33760 31694
rect 33840 31746 33920 31760
rect 33840 31694 33854 31746
rect 33906 31694 33920 31746
rect 33840 31680 33920 31694
rect 34000 31746 34080 31760
rect 34000 31694 34014 31746
rect 34066 31694 34080 31746
rect 34000 31680 34080 31694
rect 34160 31746 34240 31760
rect 34160 31694 34174 31746
rect 34226 31694 34240 31746
rect 34160 31680 34240 31694
rect 34320 31746 34400 31760
rect 34320 31694 34334 31746
rect 34386 31694 34400 31746
rect 34320 31680 34400 31694
rect 34480 31746 34560 31760
rect 34480 31694 34494 31746
rect 34546 31694 34560 31746
rect 34480 31680 34560 31694
rect 34640 31746 34720 31760
rect 34640 31694 34654 31746
rect 34706 31694 34720 31746
rect 34640 31680 34720 31694
rect 34800 31746 34880 31760
rect 34800 31694 34814 31746
rect 34866 31694 34880 31746
rect 34800 31680 34880 31694
rect 34960 31746 35040 31760
rect 34960 31694 34974 31746
rect 35026 31694 35040 31746
rect 34960 31680 35040 31694
rect 35120 31746 35200 31760
rect 35120 31694 35134 31746
rect 35186 31694 35200 31746
rect 35120 31680 35200 31694
rect 35280 31746 35360 31760
rect 35280 31694 35294 31746
rect 35346 31694 35360 31746
rect 35280 31680 35360 31694
rect 35440 31746 35520 31760
rect 35440 31694 35454 31746
rect 35506 31694 35520 31746
rect 35440 31680 35520 31694
rect 35600 31746 35680 31760
rect 35600 31694 35614 31746
rect 35666 31694 35680 31746
rect 35600 31680 35680 31694
rect 35760 31746 35840 31760
rect 35760 31694 35774 31746
rect 35826 31694 35840 31746
rect 35760 31680 35840 31694
rect 35920 31746 36000 31760
rect 35920 31694 35934 31746
rect 35986 31694 36000 31746
rect 35920 31680 36000 31694
rect 36080 31746 36160 31760
rect 36080 31694 36094 31746
rect 36146 31694 36160 31746
rect 36080 31680 36160 31694
rect 36240 31746 36320 31760
rect 36240 31694 36254 31746
rect 36306 31694 36320 31746
rect 36240 31680 36320 31694
rect 36400 31746 36480 31760
rect 36400 31694 36414 31746
rect 36466 31694 36480 31746
rect 36400 31680 36480 31694
rect 36560 31746 36640 31760
rect 36560 31694 36574 31746
rect 36626 31694 36640 31746
rect 36560 31680 36640 31694
rect 36720 31746 36800 31760
rect 36720 31694 36734 31746
rect 36786 31694 36800 31746
rect 36720 31680 36800 31694
rect 36880 31746 36960 31760
rect 36880 31694 36894 31746
rect 36946 31694 36960 31746
rect 36880 31680 36960 31694
rect 37040 31746 37120 31760
rect 37040 31694 37054 31746
rect 37106 31694 37120 31746
rect 37040 31680 37120 31694
rect 37200 31746 37280 31760
rect 37200 31694 37214 31746
rect 37266 31694 37280 31746
rect 37200 31680 37280 31694
rect 37360 31746 37440 31760
rect 37360 31694 37374 31746
rect 37426 31694 37440 31746
rect 37360 31680 37440 31694
rect 37520 31746 37600 31760
rect 37520 31694 37534 31746
rect 37586 31694 37600 31746
rect 37520 31680 37600 31694
rect 37680 31746 37760 31760
rect 37680 31694 37694 31746
rect 37746 31694 37760 31746
rect 37680 31680 37760 31694
rect 37840 31746 37920 31760
rect 37840 31694 37854 31746
rect 37906 31694 37920 31746
rect 37840 31680 37920 31694
rect 38000 31746 38080 31760
rect 38000 31694 38014 31746
rect 38066 31694 38080 31746
rect 38000 31680 38080 31694
rect 38160 31746 38240 31760
rect 38160 31694 38174 31746
rect 38226 31694 38240 31746
rect 38160 31680 38240 31694
rect 38320 31746 38400 31760
rect 38320 31694 38334 31746
rect 38386 31694 38400 31746
rect 38320 31680 38400 31694
rect 38480 31746 38560 31760
rect 38480 31694 38494 31746
rect 38546 31694 38560 31746
rect 38480 31680 38560 31694
rect 38640 31746 38720 31760
rect 38640 31694 38654 31746
rect 38706 31694 38720 31746
rect 38640 31680 38720 31694
rect 38800 31746 38880 31760
rect 38800 31694 38814 31746
rect 38866 31694 38880 31746
rect 38800 31680 38880 31694
rect 38960 31746 39040 31760
rect 38960 31694 38974 31746
rect 39026 31694 39040 31746
rect 38960 31680 39040 31694
rect 39120 31746 39200 31760
rect 39120 31694 39134 31746
rect 39186 31694 39200 31746
rect 39120 31680 39200 31694
rect 39280 31746 39360 31760
rect 39280 31694 39294 31746
rect 39346 31694 39360 31746
rect 39280 31680 39360 31694
rect 39440 31746 39520 31760
rect 39440 31694 39454 31746
rect 39506 31694 39520 31746
rect 39440 31680 39520 31694
rect 39600 31746 39680 31760
rect 39600 31694 39614 31746
rect 39666 31694 39680 31746
rect 39600 31680 39680 31694
rect 39760 31746 39840 31760
rect 39760 31694 39774 31746
rect 39826 31694 39840 31746
rect 39760 31680 39840 31694
rect 39920 31746 40000 31760
rect 39920 31694 39934 31746
rect 39986 31694 40000 31746
rect 39920 31680 40000 31694
rect 40080 31746 40160 31760
rect 40080 31694 40094 31746
rect 40146 31694 40160 31746
rect 40080 31680 40160 31694
rect 40240 31746 40320 31760
rect 40240 31694 40254 31746
rect 40306 31694 40320 31746
rect 40240 31680 40320 31694
rect 40400 31746 40480 31760
rect 40400 31694 40414 31746
rect 40466 31694 40480 31746
rect 40400 31680 40480 31694
rect 40560 31746 40640 31760
rect 40560 31694 40574 31746
rect 40626 31694 40640 31746
rect 40560 31680 40640 31694
rect 40720 31746 40800 31760
rect 40720 31694 40734 31746
rect 40786 31694 40800 31746
rect 40720 31680 40800 31694
rect 40880 31746 40960 31760
rect 40880 31694 40894 31746
rect 40946 31694 40960 31746
rect 40880 31680 40960 31694
rect 41040 31746 41120 31760
rect 41040 31694 41054 31746
rect 41106 31694 41120 31746
rect 41040 31680 41120 31694
rect 41200 31746 41280 31760
rect 41200 31694 41214 31746
rect 41266 31694 41280 31746
rect 41200 31680 41280 31694
rect 41360 31746 41440 31760
rect 41360 31694 41374 31746
rect 41426 31694 41440 31746
rect 41360 31680 41440 31694
rect 41520 31746 41600 31760
rect 41520 31694 41534 31746
rect 41586 31694 41600 31746
rect 41520 31680 41600 31694
rect 41680 31746 41760 31760
rect 41680 31694 41694 31746
rect 41746 31694 41760 31746
rect 41680 31680 41760 31694
rect 41840 31746 41920 31760
rect 41840 31694 41854 31746
rect 41906 31694 41920 31746
rect 41840 31680 41920 31694
rect 0 31426 80 31440
rect 0 31374 14 31426
rect 66 31374 80 31426
rect 0 31360 80 31374
rect 160 31426 240 31440
rect 160 31374 174 31426
rect 226 31374 240 31426
rect 160 31360 240 31374
rect 320 31426 400 31440
rect 320 31374 334 31426
rect 386 31374 400 31426
rect 320 31360 400 31374
rect 480 31426 560 31440
rect 480 31374 494 31426
rect 546 31374 560 31426
rect 480 31360 560 31374
rect 640 31426 720 31440
rect 640 31374 654 31426
rect 706 31374 720 31426
rect 640 31360 720 31374
rect 800 31426 880 31440
rect 800 31374 814 31426
rect 866 31374 880 31426
rect 800 31360 880 31374
rect 960 31426 1040 31440
rect 960 31374 974 31426
rect 1026 31374 1040 31426
rect 960 31360 1040 31374
rect 1120 31426 1200 31440
rect 1120 31374 1134 31426
rect 1186 31374 1200 31426
rect 1120 31360 1200 31374
rect 1280 31426 1360 31440
rect 1280 31374 1294 31426
rect 1346 31374 1360 31426
rect 1280 31360 1360 31374
rect 1440 31426 1520 31440
rect 1440 31374 1454 31426
rect 1506 31374 1520 31426
rect 1440 31360 1520 31374
rect 1600 31426 1680 31440
rect 1600 31374 1614 31426
rect 1666 31374 1680 31426
rect 1600 31360 1680 31374
rect 1760 31426 1840 31440
rect 1760 31374 1774 31426
rect 1826 31374 1840 31426
rect 1760 31360 1840 31374
rect 1920 31426 2000 31440
rect 1920 31374 1934 31426
rect 1986 31374 2000 31426
rect 1920 31360 2000 31374
rect 2080 31426 2160 31440
rect 2080 31374 2094 31426
rect 2146 31374 2160 31426
rect 2080 31360 2160 31374
rect 2240 31426 2320 31440
rect 2240 31374 2254 31426
rect 2306 31374 2320 31426
rect 2240 31360 2320 31374
rect 2400 31426 2480 31440
rect 2400 31374 2414 31426
rect 2466 31374 2480 31426
rect 2400 31360 2480 31374
rect 2560 31426 2640 31440
rect 2560 31374 2574 31426
rect 2626 31374 2640 31426
rect 2560 31360 2640 31374
rect 2720 31426 2800 31440
rect 2720 31374 2734 31426
rect 2786 31374 2800 31426
rect 2720 31360 2800 31374
rect 2880 31426 2960 31440
rect 2880 31374 2894 31426
rect 2946 31374 2960 31426
rect 2880 31360 2960 31374
rect 3040 31426 3120 31440
rect 3040 31374 3054 31426
rect 3106 31374 3120 31426
rect 3040 31360 3120 31374
rect 3200 31426 3280 31440
rect 3200 31374 3214 31426
rect 3266 31374 3280 31426
rect 3200 31360 3280 31374
rect 3360 31426 3440 31440
rect 3360 31374 3374 31426
rect 3426 31374 3440 31426
rect 3360 31360 3440 31374
rect 3520 31426 3600 31440
rect 3520 31374 3534 31426
rect 3586 31374 3600 31426
rect 3520 31360 3600 31374
rect 3680 31426 3760 31440
rect 3680 31374 3694 31426
rect 3746 31374 3760 31426
rect 3680 31360 3760 31374
rect 3840 31426 3920 31440
rect 3840 31374 3854 31426
rect 3906 31374 3920 31426
rect 3840 31360 3920 31374
rect 4000 31426 4080 31440
rect 4000 31374 4014 31426
rect 4066 31374 4080 31426
rect 4000 31360 4080 31374
rect 4160 31426 4240 31440
rect 4160 31374 4174 31426
rect 4226 31374 4240 31426
rect 4160 31360 4240 31374
rect 4320 31426 4400 31440
rect 4320 31374 4334 31426
rect 4386 31374 4400 31426
rect 4320 31360 4400 31374
rect 4480 31426 4560 31440
rect 4480 31374 4494 31426
rect 4546 31374 4560 31426
rect 4480 31360 4560 31374
rect 4640 31426 4720 31440
rect 4640 31374 4654 31426
rect 4706 31374 4720 31426
rect 4640 31360 4720 31374
rect 4800 31426 4880 31440
rect 4800 31374 4814 31426
rect 4866 31374 4880 31426
rect 4800 31360 4880 31374
rect 4960 31426 5040 31440
rect 4960 31374 4974 31426
rect 5026 31374 5040 31426
rect 4960 31360 5040 31374
rect 5120 31426 5200 31440
rect 5120 31374 5134 31426
rect 5186 31374 5200 31426
rect 5120 31360 5200 31374
rect 5280 31426 5360 31440
rect 5280 31374 5294 31426
rect 5346 31374 5360 31426
rect 5280 31360 5360 31374
rect 5440 31426 5520 31440
rect 5440 31374 5454 31426
rect 5506 31374 5520 31426
rect 5440 31360 5520 31374
rect 5600 31426 5680 31440
rect 5600 31374 5614 31426
rect 5666 31374 5680 31426
rect 5600 31360 5680 31374
rect 5760 31426 5840 31440
rect 5760 31374 5774 31426
rect 5826 31374 5840 31426
rect 5760 31360 5840 31374
rect 5920 31426 6000 31440
rect 5920 31374 5934 31426
rect 5986 31374 6000 31426
rect 5920 31360 6000 31374
rect 6080 31426 6160 31440
rect 6080 31374 6094 31426
rect 6146 31374 6160 31426
rect 6080 31360 6160 31374
rect 6240 31426 6320 31440
rect 6240 31374 6254 31426
rect 6306 31374 6320 31426
rect 6240 31360 6320 31374
rect 6400 31426 6480 31440
rect 6400 31374 6414 31426
rect 6466 31374 6480 31426
rect 6400 31360 6480 31374
rect 6560 31426 6640 31440
rect 6560 31374 6574 31426
rect 6626 31374 6640 31426
rect 6560 31360 6640 31374
rect 6720 31426 6800 31440
rect 6720 31374 6734 31426
rect 6786 31374 6800 31426
rect 6720 31360 6800 31374
rect 6880 31426 6960 31440
rect 6880 31374 6894 31426
rect 6946 31374 6960 31426
rect 6880 31360 6960 31374
rect 7040 31426 7120 31440
rect 7040 31374 7054 31426
rect 7106 31374 7120 31426
rect 7040 31360 7120 31374
rect 7200 31426 7280 31440
rect 7200 31374 7214 31426
rect 7266 31374 7280 31426
rect 7200 31360 7280 31374
rect 7360 31426 7440 31440
rect 7360 31374 7374 31426
rect 7426 31374 7440 31426
rect 7360 31360 7440 31374
rect 7520 31426 7600 31440
rect 7520 31374 7534 31426
rect 7586 31374 7600 31426
rect 7520 31360 7600 31374
rect 7680 31426 7760 31440
rect 7680 31374 7694 31426
rect 7746 31374 7760 31426
rect 7680 31360 7760 31374
rect 7840 31426 7920 31440
rect 7840 31374 7854 31426
rect 7906 31374 7920 31426
rect 7840 31360 7920 31374
rect 8000 31426 8080 31440
rect 8000 31374 8014 31426
rect 8066 31374 8080 31426
rect 8000 31360 8080 31374
rect 8160 31426 8240 31440
rect 8160 31374 8174 31426
rect 8226 31374 8240 31426
rect 8160 31360 8240 31374
rect 8320 31426 8400 31440
rect 8320 31374 8334 31426
rect 8386 31374 8400 31426
rect 8320 31360 8400 31374
rect 12480 31426 12560 31440
rect 12480 31374 12494 31426
rect 12546 31374 12560 31426
rect 12480 31360 12560 31374
rect 12640 31426 12720 31440
rect 12640 31374 12654 31426
rect 12706 31374 12720 31426
rect 12640 31360 12720 31374
rect 12800 31426 12880 31440
rect 12800 31374 12814 31426
rect 12866 31374 12880 31426
rect 12800 31360 12880 31374
rect 12960 31426 13040 31440
rect 12960 31374 12974 31426
rect 13026 31374 13040 31426
rect 12960 31360 13040 31374
rect 13120 31426 13200 31440
rect 13120 31374 13134 31426
rect 13186 31374 13200 31426
rect 13120 31360 13200 31374
rect 13280 31426 13360 31440
rect 13280 31374 13294 31426
rect 13346 31374 13360 31426
rect 13280 31360 13360 31374
rect 13440 31426 13520 31440
rect 13440 31374 13454 31426
rect 13506 31374 13520 31426
rect 13440 31360 13520 31374
rect 13600 31426 13680 31440
rect 13600 31374 13614 31426
rect 13666 31374 13680 31426
rect 13600 31360 13680 31374
rect 13760 31426 13840 31440
rect 13760 31374 13774 31426
rect 13826 31374 13840 31426
rect 13760 31360 13840 31374
rect 13920 31426 14000 31440
rect 13920 31374 13934 31426
rect 13986 31374 14000 31426
rect 13920 31360 14000 31374
rect 14080 31426 14160 31440
rect 14080 31374 14094 31426
rect 14146 31374 14160 31426
rect 14080 31360 14160 31374
rect 14240 31426 14320 31440
rect 14240 31374 14254 31426
rect 14306 31374 14320 31426
rect 14240 31360 14320 31374
rect 14400 31426 14480 31440
rect 14400 31374 14414 31426
rect 14466 31374 14480 31426
rect 14400 31360 14480 31374
rect 14560 31426 14640 31440
rect 14560 31374 14574 31426
rect 14626 31374 14640 31426
rect 14560 31360 14640 31374
rect 14720 31426 14800 31440
rect 14720 31374 14734 31426
rect 14786 31374 14800 31426
rect 14720 31360 14800 31374
rect 14880 31426 14960 31440
rect 14880 31374 14894 31426
rect 14946 31374 14960 31426
rect 14880 31360 14960 31374
rect 15040 31426 15120 31440
rect 15040 31374 15054 31426
rect 15106 31374 15120 31426
rect 15040 31360 15120 31374
rect 15200 31426 15280 31440
rect 15200 31374 15214 31426
rect 15266 31374 15280 31426
rect 15200 31360 15280 31374
rect 15360 31426 15440 31440
rect 15360 31374 15374 31426
rect 15426 31374 15440 31426
rect 15360 31360 15440 31374
rect 15520 31426 15600 31440
rect 15520 31374 15534 31426
rect 15586 31374 15600 31426
rect 15520 31360 15600 31374
rect 15680 31426 15760 31440
rect 15680 31374 15694 31426
rect 15746 31374 15760 31426
rect 15680 31360 15760 31374
rect 15840 31426 15920 31440
rect 15840 31374 15854 31426
rect 15906 31374 15920 31426
rect 15840 31360 15920 31374
rect 16000 31426 16080 31440
rect 16000 31374 16014 31426
rect 16066 31374 16080 31426
rect 16000 31360 16080 31374
rect 16160 31426 16240 31440
rect 16160 31374 16174 31426
rect 16226 31374 16240 31426
rect 16160 31360 16240 31374
rect 16320 31426 16400 31440
rect 16320 31374 16334 31426
rect 16386 31374 16400 31426
rect 16320 31360 16400 31374
rect 16480 31426 16560 31440
rect 16480 31374 16494 31426
rect 16546 31374 16560 31426
rect 16480 31360 16560 31374
rect 16640 31426 16720 31440
rect 16640 31374 16654 31426
rect 16706 31374 16720 31426
rect 16640 31360 16720 31374
rect 16800 31426 16880 31440
rect 16800 31374 16814 31426
rect 16866 31374 16880 31426
rect 16800 31360 16880 31374
rect 16960 31426 17040 31440
rect 16960 31374 16974 31426
rect 17026 31374 17040 31426
rect 16960 31360 17040 31374
rect 17120 31426 17200 31440
rect 17120 31374 17134 31426
rect 17186 31374 17200 31426
rect 17120 31360 17200 31374
rect 17280 31426 17360 31440
rect 17280 31374 17294 31426
rect 17346 31374 17360 31426
rect 17280 31360 17360 31374
rect 17440 31426 17520 31440
rect 17440 31374 17454 31426
rect 17506 31374 17520 31426
rect 17440 31360 17520 31374
rect 17600 31426 17680 31440
rect 17600 31374 17614 31426
rect 17666 31374 17680 31426
rect 17600 31360 17680 31374
rect 17760 31426 17840 31440
rect 17760 31374 17774 31426
rect 17826 31374 17840 31426
rect 17760 31360 17840 31374
rect 17920 31426 18000 31440
rect 17920 31374 17934 31426
rect 17986 31374 18000 31426
rect 17920 31360 18000 31374
rect 18080 31426 18160 31440
rect 18080 31374 18094 31426
rect 18146 31374 18160 31426
rect 18080 31360 18160 31374
rect 18240 31426 18320 31440
rect 18240 31374 18254 31426
rect 18306 31374 18320 31426
rect 18240 31360 18320 31374
rect 18400 31426 18480 31440
rect 18400 31374 18414 31426
rect 18466 31374 18480 31426
rect 18400 31360 18480 31374
rect 18560 31426 18640 31440
rect 18560 31374 18574 31426
rect 18626 31374 18640 31426
rect 18560 31360 18640 31374
rect 18720 31426 18800 31440
rect 18720 31374 18734 31426
rect 18786 31374 18800 31426
rect 18720 31360 18800 31374
rect 18880 31426 18960 31440
rect 18880 31374 18894 31426
rect 18946 31374 18960 31426
rect 18880 31360 18960 31374
rect 23120 31426 23200 31440
rect 23120 31374 23134 31426
rect 23186 31374 23200 31426
rect 23120 31360 23200 31374
rect 23280 31426 23360 31440
rect 23280 31374 23294 31426
rect 23346 31374 23360 31426
rect 23280 31360 23360 31374
rect 23440 31426 23520 31440
rect 23440 31374 23454 31426
rect 23506 31374 23520 31426
rect 23440 31360 23520 31374
rect 23600 31426 23680 31440
rect 23600 31374 23614 31426
rect 23666 31374 23680 31426
rect 23600 31360 23680 31374
rect 23760 31426 23840 31440
rect 23760 31374 23774 31426
rect 23826 31374 23840 31426
rect 23760 31360 23840 31374
rect 23920 31426 24000 31440
rect 23920 31374 23934 31426
rect 23986 31374 24000 31426
rect 23920 31360 24000 31374
rect 24080 31426 24160 31440
rect 24080 31374 24094 31426
rect 24146 31374 24160 31426
rect 24080 31360 24160 31374
rect 24240 31426 24320 31440
rect 24240 31374 24254 31426
rect 24306 31374 24320 31426
rect 24240 31360 24320 31374
rect 24400 31426 24480 31440
rect 24400 31374 24414 31426
rect 24466 31374 24480 31426
rect 24400 31360 24480 31374
rect 24560 31426 24640 31440
rect 24560 31374 24574 31426
rect 24626 31374 24640 31426
rect 24560 31360 24640 31374
rect 24720 31426 24800 31440
rect 24720 31374 24734 31426
rect 24786 31374 24800 31426
rect 24720 31360 24800 31374
rect 24880 31426 24960 31440
rect 24880 31374 24894 31426
rect 24946 31374 24960 31426
rect 24880 31360 24960 31374
rect 25040 31426 25120 31440
rect 25040 31374 25054 31426
rect 25106 31374 25120 31426
rect 25040 31360 25120 31374
rect 25200 31426 25280 31440
rect 25200 31374 25214 31426
rect 25266 31374 25280 31426
rect 25200 31360 25280 31374
rect 25360 31426 25440 31440
rect 25360 31374 25374 31426
rect 25426 31374 25440 31426
rect 25360 31360 25440 31374
rect 25520 31426 25600 31440
rect 25520 31374 25534 31426
rect 25586 31374 25600 31426
rect 25520 31360 25600 31374
rect 25680 31426 25760 31440
rect 25680 31374 25694 31426
rect 25746 31374 25760 31426
rect 25680 31360 25760 31374
rect 25840 31426 25920 31440
rect 25840 31374 25854 31426
rect 25906 31374 25920 31426
rect 25840 31360 25920 31374
rect 26000 31426 26080 31440
rect 26000 31374 26014 31426
rect 26066 31374 26080 31426
rect 26000 31360 26080 31374
rect 26160 31426 26240 31440
rect 26160 31374 26174 31426
rect 26226 31374 26240 31426
rect 26160 31360 26240 31374
rect 26320 31426 26400 31440
rect 26320 31374 26334 31426
rect 26386 31374 26400 31426
rect 26320 31360 26400 31374
rect 26480 31426 26560 31440
rect 26480 31374 26494 31426
rect 26546 31374 26560 31426
rect 26480 31360 26560 31374
rect 26640 31426 26720 31440
rect 26640 31374 26654 31426
rect 26706 31374 26720 31426
rect 26640 31360 26720 31374
rect 26800 31426 26880 31440
rect 26800 31374 26814 31426
rect 26866 31374 26880 31426
rect 26800 31360 26880 31374
rect 26960 31426 27040 31440
rect 26960 31374 26974 31426
rect 27026 31374 27040 31426
rect 26960 31360 27040 31374
rect 27120 31426 27200 31440
rect 27120 31374 27134 31426
rect 27186 31374 27200 31426
rect 27120 31360 27200 31374
rect 27280 31426 27360 31440
rect 27280 31374 27294 31426
rect 27346 31374 27360 31426
rect 27280 31360 27360 31374
rect 27440 31426 27520 31440
rect 27440 31374 27454 31426
rect 27506 31374 27520 31426
rect 27440 31360 27520 31374
rect 27600 31426 27680 31440
rect 27600 31374 27614 31426
rect 27666 31374 27680 31426
rect 27600 31360 27680 31374
rect 27760 31426 27840 31440
rect 27760 31374 27774 31426
rect 27826 31374 27840 31426
rect 27760 31360 27840 31374
rect 27920 31426 28000 31440
rect 27920 31374 27934 31426
rect 27986 31374 28000 31426
rect 27920 31360 28000 31374
rect 28080 31426 28160 31440
rect 28080 31374 28094 31426
rect 28146 31374 28160 31426
rect 28080 31360 28160 31374
rect 28240 31426 28320 31440
rect 28240 31374 28254 31426
rect 28306 31374 28320 31426
rect 28240 31360 28320 31374
rect 28400 31426 28480 31440
rect 28400 31374 28414 31426
rect 28466 31374 28480 31426
rect 28400 31360 28480 31374
rect 28560 31426 28640 31440
rect 28560 31374 28574 31426
rect 28626 31374 28640 31426
rect 28560 31360 28640 31374
rect 28720 31426 28800 31440
rect 28720 31374 28734 31426
rect 28786 31374 28800 31426
rect 28720 31360 28800 31374
rect 28880 31426 28960 31440
rect 28880 31374 28894 31426
rect 28946 31374 28960 31426
rect 28880 31360 28960 31374
rect 29040 31426 29120 31440
rect 29040 31374 29054 31426
rect 29106 31374 29120 31426
rect 29040 31360 29120 31374
rect 29200 31426 29280 31440
rect 29200 31374 29214 31426
rect 29266 31374 29280 31426
rect 29200 31360 29280 31374
rect 29360 31426 29440 31440
rect 29360 31374 29374 31426
rect 29426 31374 29440 31426
rect 29360 31360 29440 31374
rect 33520 31426 33600 31440
rect 33520 31374 33534 31426
rect 33586 31374 33600 31426
rect 33520 31360 33600 31374
rect 33680 31426 33760 31440
rect 33680 31374 33694 31426
rect 33746 31374 33760 31426
rect 33680 31360 33760 31374
rect 33840 31426 33920 31440
rect 33840 31374 33854 31426
rect 33906 31374 33920 31426
rect 33840 31360 33920 31374
rect 34000 31426 34080 31440
rect 34000 31374 34014 31426
rect 34066 31374 34080 31426
rect 34000 31360 34080 31374
rect 34160 31426 34240 31440
rect 34160 31374 34174 31426
rect 34226 31374 34240 31426
rect 34160 31360 34240 31374
rect 34320 31426 34400 31440
rect 34320 31374 34334 31426
rect 34386 31374 34400 31426
rect 34320 31360 34400 31374
rect 34480 31426 34560 31440
rect 34480 31374 34494 31426
rect 34546 31374 34560 31426
rect 34480 31360 34560 31374
rect 34640 31426 34720 31440
rect 34640 31374 34654 31426
rect 34706 31374 34720 31426
rect 34640 31360 34720 31374
rect 34800 31426 34880 31440
rect 34800 31374 34814 31426
rect 34866 31374 34880 31426
rect 34800 31360 34880 31374
rect 34960 31426 35040 31440
rect 34960 31374 34974 31426
rect 35026 31374 35040 31426
rect 34960 31360 35040 31374
rect 35120 31426 35200 31440
rect 35120 31374 35134 31426
rect 35186 31374 35200 31426
rect 35120 31360 35200 31374
rect 35280 31426 35360 31440
rect 35280 31374 35294 31426
rect 35346 31374 35360 31426
rect 35280 31360 35360 31374
rect 35440 31426 35520 31440
rect 35440 31374 35454 31426
rect 35506 31374 35520 31426
rect 35440 31360 35520 31374
rect 35600 31426 35680 31440
rect 35600 31374 35614 31426
rect 35666 31374 35680 31426
rect 35600 31360 35680 31374
rect 35760 31426 35840 31440
rect 35760 31374 35774 31426
rect 35826 31374 35840 31426
rect 35760 31360 35840 31374
rect 35920 31426 36000 31440
rect 35920 31374 35934 31426
rect 35986 31374 36000 31426
rect 35920 31360 36000 31374
rect 36080 31426 36160 31440
rect 36080 31374 36094 31426
rect 36146 31374 36160 31426
rect 36080 31360 36160 31374
rect 36240 31426 36320 31440
rect 36240 31374 36254 31426
rect 36306 31374 36320 31426
rect 36240 31360 36320 31374
rect 36400 31426 36480 31440
rect 36400 31374 36414 31426
rect 36466 31374 36480 31426
rect 36400 31360 36480 31374
rect 36560 31426 36640 31440
rect 36560 31374 36574 31426
rect 36626 31374 36640 31426
rect 36560 31360 36640 31374
rect 36720 31426 36800 31440
rect 36720 31374 36734 31426
rect 36786 31374 36800 31426
rect 36720 31360 36800 31374
rect 36880 31426 36960 31440
rect 36880 31374 36894 31426
rect 36946 31374 36960 31426
rect 36880 31360 36960 31374
rect 37040 31426 37120 31440
rect 37040 31374 37054 31426
rect 37106 31374 37120 31426
rect 37040 31360 37120 31374
rect 37200 31426 37280 31440
rect 37200 31374 37214 31426
rect 37266 31374 37280 31426
rect 37200 31360 37280 31374
rect 37360 31426 37440 31440
rect 37360 31374 37374 31426
rect 37426 31374 37440 31426
rect 37360 31360 37440 31374
rect 37520 31426 37600 31440
rect 37520 31374 37534 31426
rect 37586 31374 37600 31426
rect 37520 31360 37600 31374
rect 37680 31426 37760 31440
rect 37680 31374 37694 31426
rect 37746 31374 37760 31426
rect 37680 31360 37760 31374
rect 37840 31426 37920 31440
rect 37840 31374 37854 31426
rect 37906 31374 37920 31426
rect 37840 31360 37920 31374
rect 38000 31426 38080 31440
rect 38000 31374 38014 31426
rect 38066 31374 38080 31426
rect 38000 31360 38080 31374
rect 38160 31426 38240 31440
rect 38160 31374 38174 31426
rect 38226 31374 38240 31426
rect 38160 31360 38240 31374
rect 38320 31426 38400 31440
rect 38320 31374 38334 31426
rect 38386 31374 38400 31426
rect 38320 31360 38400 31374
rect 38480 31426 38560 31440
rect 38480 31374 38494 31426
rect 38546 31374 38560 31426
rect 38480 31360 38560 31374
rect 38640 31426 38720 31440
rect 38640 31374 38654 31426
rect 38706 31374 38720 31426
rect 38640 31360 38720 31374
rect 38800 31426 38880 31440
rect 38800 31374 38814 31426
rect 38866 31374 38880 31426
rect 38800 31360 38880 31374
rect 38960 31426 39040 31440
rect 38960 31374 38974 31426
rect 39026 31374 39040 31426
rect 38960 31360 39040 31374
rect 39120 31426 39200 31440
rect 39120 31374 39134 31426
rect 39186 31374 39200 31426
rect 39120 31360 39200 31374
rect 39280 31426 39360 31440
rect 39280 31374 39294 31426
rect 39346 31374 39360 31426
rect 39280 31360 39360 31374
rect 39440 31426 39520 31440
rect 39440 31374 39454 31426
rect 39506 31374 39520 31426
rect 39440 31360 39520 31374
rect 39600 31426 39680 31440
rect 39600 31374 39614 31426
rect 39666 31374 39680 31426
rect 39600 31360 39680 31374
rect 39760 31426 39840 31440
rect 39760 31374 39774 31426
rect 39826 31374 39840 31426
rect 39760 31360 39840 31374
rect 39920 31426 40000 31440
rect 39920 31374 39934 31426
rect 39986 31374 40000 31426
rect 39920 31360 40000 31374
rect 40080 31426 40160 31440
rect 40080 31374 40094 31426
rect 40146 31374 40160 31426
rect 40080 31360 40160 31374
rect 40240 31426 40320 31440
rect 40240 31374 40254 31426
rect 40306 31374 40320 31426
rect 40240 31360 40320 31374
rect 40400 31426 40480 31440
rect 40400 31374 40414 31426
rect 40466 31374 40480 31426
rect 40400 31360 40480 31374
rect 40560 31426 40640 31440
rect 40560 31374 40574 31426
rect 40626 31374 40640 31426
rect 40560 31360 40640 31374
rect 40720 31426 40800 31440
rect 40720 31374 40734 31426
rect 40786 31374 40800 31426
rect 40720 31360 40800 31374
rect 40880 31426 40960 31440
rect 40880 31374 40894 31426
rect 40946 31374 40960 31426
rect 40880 31360 40960 31374
rect 41040 31426 41120 31440
rect 41040 31374 41054 31426
rect 41106 31374 41120 31426
rect 41040 31360 41120 31374
rect 41200 31426 41280 31440
rect 41200 31374 41214 31426
rect 41266 31374 41280 31426
rect 41200 31360 41280 31374
rect 41360 31426 41440 31440
rect 41360 31374 41374 31426
rect 41426 31374 41440 31426
rect 41360 31360 41440 31374
rect 41520 31426 41600 31440
rect 41520 31374 41534 31426
rect 41586 31374 41600 31426
rect 41520 31360 41600 31374
rect 41680 31426 41760 31440
rect 41680 31374 41694 31426
rect 41746 31374 41760 31426
rect 41680 31360 41760 31374
rect 41840 31426 41920 31440
rect 41840 31374 41854 31426
rect 41906 31374 41920 31426
rect 41840 31360 41920 31374
rect 0 31106 80 31120
rect 0 31054 14 31106
rect 66 31054 80 31106
rect 0 31040 80 31054
rect 160 31106 240 31120
rect 160 31054 174 31106
rect 226 31054 240 31106
rect 160 31040 240 31054
rect 320 31106 400 31120
rect 320 31054 334 31106
rect 386 31054 400 31106
rect 320 31040 400 31054
rect 480 31106 560 31120
rect 480 31054 494 31106
rect 546 31054 560 31106
rect 480 31040 560 31054
rect 640 31106 720 31120
rect 640 31054 654 31106
rect 706 31054 720 31106
rect 640 31040 720 31054
rect 800 31106 880 31120
rect 800 31054 814 31106
rect 866 31054 880 31106
rect 800 31040 880 31054
rect 960 31106 1040 31120
rect 960 31054 974 31106
rect 1026 31054 1040 31106
rect 960 31040 1040 31054
rect 1120 31106 1200 31120
rect 1120 31054 1134 31106
rect 1186 31054 1200 31106
rect 1120 31040 1200 31054
rect 1280 31106 1360 31120
rect 1280 31054 1294 31106
rect 1346 31054 1360 31106
rect 1280 31040 1360 31054
rect 1440 31106 1520 31120
rect 1440 31054 1454 31106
rect 1506 31054 1520 31106
rect 1440 31040 1520 31054
rect 1600 31106 1680 31120
rect 1600 31054 1614 31106
rect 1666 31054 1680 31106
rect 1600 31040 1680 31054
rect 1760 31106 1840 31120
rect 1760 31054 1774 31106
rect 1826 31054 1840 31106
rect 1760 31040 1840 31054
rect 1920 31106 2000 31120
rect 1920 31054 1934 31106
rect 1986 31054 2000 31106
rect 1920 31040 2000 31054
rect 2080 31106 2160 31120
rect 2080 31054 2094 31106
rect 2146 31054 2160 31106
rect 2080 31040 2160 31054
rect 2240 31106 2320 31120
rect 2240 31054 2254 31106
rect 2306 31054 2320 31106
rect 2240 31040 2320 31054
rect 2400 31106 2480 31120
rect 2400 31054 2414 31106
rect 2466 31054 2480 31106
rect 2400 31040 2480 31054
rect 2560 31106 2640 31120
rect 2560 31054 2574 31106
rect 2626 31054 2640 31106
rect 2560 31040 2640 31054
rect 2720 31106 2800 31120
rect 2720 31054 2734 31106
rect 2786 31054 2800 31106
rect 2720 31040 2800 31054
rect 2880 31106 2960 31120
rect 2880 31054 2894 31106
rect 2946 31054 2960 31106
rect 2880 31040 2960 31054
rect 3040 31106 3120 31120
rect 3040 31054 3054 31106
rect 3106 31054 3120 31106
rect 3040 31040 3120 31054
rect 3200 31106 3280 31120
rect 3200 31054 3214 31106
rect 3266 31054 3280 31106
rect 3200 31040 3280 31054
rect 3360 31106 3440 31120
rect 3360 31054 3374 31106
rect 3426 31054 3440 31106
rect 3360 31040 3440 31054
rect 3520 31106 3600 31120
rect 3520 31054 3534 31106
rect 3586 31054 3600 31106
rect 3520 31040 3600 31054
rect 3680 31106 3760 31120
rect 3680 31054 3694 31106
rect 3746 31054 3760 31106
rect 3680 31040 3760 31054
rect 3840 31106 3920 31120
rect 3840 31054 3854 31106
rect 3906 31054 3920 31106
rect 3840 31040 3920 31054
rect 4000 31106 4080 31120
rect 4000 31054 4014 31106
rect 4066 31054 4080 31106
rect 4000 31040 4080 31054
rect 4160 31106 4240 31120
rect 4160 31054 4174 31106
rect 4226 31054 4240 31106
rect 4160 31040 4240 31054
rect 4320 31106 4400 31120
rect 4320 31054 4334 31106
rect 4386 31054 4400 31106
rect 4320 31040 4400 31054
rect 4480 31106 4560 31120
rect 4480 31054 4494 31106
rect 4546 31054 4560 31106
rect 4480 31040 4560 31054
rect 4640 31106 4720 31120
rect 4640 31054 4654 31106
rect 4706 31054 4720 31106
rect 4640 31040 4720 31054
rect 4800 31106 4880 31120
rect 4800 31054 4814 31106
rect 4866 31054 4880 31106
rect 4800 31040 4880 31054
rect 4960 31106 5040 31120
rect 4960 31054 4974 31106
rect 5026 31054 5040 31106
rect 4960 31040 5040 31054
rect 5120 31106 5200 31120
rect 5120 31054 5134 31106
rect 5186 31054 5200 31106
rect 5120 31040 5200 31054
rect 5280 31106 5360 31120
rect 5280 31054 5294 31106
rect 5346 31054 5360 31106
rect 5280 31040 5360 31054
rect 5440 31106 5520 31120
rect 5440 31054 5454 31106
rect 5506 31054 5520 31106
rect 5440 31040 5520 31054
rect 5600 31106 5680 31120
rect 5600 31054 5614 31106
rect 5666 31054 5680 31106
rect 5600 31040 5680 31054
rect 5760 31106 5840 31120
rect 5760 31054 5774 31106
rect 5826 31054 5840 31106
rect 5760 31040 5840 31054
rect 5920 31106 6000 31120
rect 5920 31054 5934 31106
rect 5986 31054 6000 31106
rect 5920 31040 6000 31054
rect 6080 31106 6160 31120
rect 6080 31054 6094 31106
rect 6146 31054 6160 31106
rect 6080 31040 6160 31054
rect 6240 31106 6320 31120
rect 6240 31054 6254 31106
rect 6306 31054 6320 31106
rect 6240 31040 6320 31054
rect 6400 31106 6480 31120
rect 6400 31054 6414 31106
rect 6466 31054 6480 31106
rect 6400 31040 6480 31054
rect 6560 31106 6640 31120
rect 6560 31054 6574 31106
rect 6626 31054 6640 31106
rect 6560 31040 6640 31054
rect 6720 31106 6800 31120
rect 6720 31054 6734 31106
rect 6786 31054 6800 31106
rect 6720 31040 6800 31054
rect 6880 31106 6960 31120
rect 6880 31054 6894 31106
rect 6946 31054 6960 31106
rect 6880 31040 6960 31054
rect 7040 31106 7120 31120
rect 7040 31054 7054 31106
rect 7106 31054 7120 31106
rect 7040 31040 7120 31054
rect 7200 31106 7280 31120
rect 7200 31054 7214 31106
rect 7266 31054 7280 31106
rect 7200 31040 7280 31054
rect 7360 31106 7440 31120
rect 7360 31054 7374 31106
rect 7426 31054 7440 31106
rect 7360 31040 7440 31054
rect 7520 31106 7600 31120
rect 7520 31054 7534 31106
rect 7586 31054 7600 31106
rect 7520 31040 7600 31054
rect 7680 31106 7760 31120
rect 7680 31054 7694 31106
rect 7746 31054 7760 31106
rect 7680 31040 7760 31054
rect 7840 31106 7920 31120
rect 7840 31054 7854 31106
rect 7906 31054 7920 31106
rect 7840 31040 7920 31054
rect 8000 31106 8080 31120
rect 8000 31054 8014 31106
rect 8066 31054 8080 31106
rect 8000 31040 8080 31054
rect 8160 31106 8240 31120
rect 8160 31054 8174 31106
rect 8226 31054 8240 31106
rect 8160 31040 8240 31054
rect 8320 31106 8400 31120
rect 8320 31054 8334 31106
rect 8386 31054 8400 31106
rect 8320 31040 8400 31054
rect 12480 31106 12560 31120
rect 12480 31054 12494 31106
rect 12546 31054 12560 31106
rect 12480 31040 12560 31054
rect 12640 31106 12720 31120
rect 12640 31054 12654 31106
rect 12706 31054 12720 31106
rect 12640 31040 12720 31054
rect 12800 31106 12880 31120
rect 12800 31054 12814 31106
rect 12866 31054 12880 31106
rect 12800 31040 12880 31054
rect 12960 31106 13040 31120
rect 12960 31054 12974 31106
rect 13026 31054 13040 31106
rect 12960 31040 13040 31054
rect 13120 31106 13200 31120
rect 13120 31054 13134 31106
rect 13186 31054 13200 31106
rect 13120 31040 13200 31054
rect 13280 31106 13360 31120
rect 13280 31054 13294 31106
rect 13346 31054 13360 31106
rect 13280 31040 13360 31054
rect 13440 31106 13520 31120
rect 13440 31054 13454 31106
rect 13506 31054 13520 31106
rect 13440 31040 13520 31054
rect 13600 31106 13680 31120
rect 13600 31054 13614 31106
rect 13666 31054 13680 31106
rect 13600 31040 13680 31054
rect 13760 31106 13840 31120
rect 13760 31054 13774 31106
rect 13826 31054 13840 31106
rect 13760 31040 13840 31054
rect 13920 31106 14000 31120
rect 13920 31054 13934 31106
rect 13986 31054 14000 31106
rect 13920 31040 14000 31054
rect 14080 31106 14160 31120
rect 14080 31054 14094 31106
rect 14146 31054 14160 31106
rect 14080 31040 14160 31054
rect 14240 31106 14320 31120
rect 14240 31054 14254 31106
rect 14306 31054 14320 31106
rect 14240 31040 14320 31054
rect 14400 31106 14480 31120
rect 14400 31054 14414 31106
rect 14466 31054 14480 31106
rect 14400 31040 14480 31054
rect 14560 31106 14640 31120
rect 14560 31054 14574 31106
rect 14626 31054 14640 31106
rect 14560 31040 14640 31054
rect 14720 31106 14800 31120
rect 14720 31054 14734 31106
rect 14786 31054 14800 31106
rect 14720 31040 14800 31054
rect 14880 31106 14960 31120
rect 14880 31054 14894 31106
rect 14946 31054 14960 31106
rect 14880 31040 14960 31054
rect 15040 31106 15120 31120
rect 15040 31054 15054 31106
rect 15106 31054 15120 31106
rect 15040 31040 15120 31054
rect 15200 31106 15280 31120
rect 15200 31054 15214 31106
rect 15266 31054 15280 31106
rect 15200 31040 15280 31054
rect 15360 31106 15440 31120
rect 15360 31054 15374 31106
rect 15426 31054 15440 31106
rect 15360 31040 15440 31054
rect 15520 31106 15600 31120
rect 15520 31054 15534 31106
rect 15586 31054 15600 31106
rect 15520 31040 15600 31054
rect 15680 31106 15760 31120
rect 15680 31054 15694 31106
rect 15746 31054 15760 31106
rect 15680 31040 15760 31054
rect 15840 31106 15920 31120
rect 15840 31054 15854 31106
rect 15906 31054 15920 31106
rect 15840 31040 15920 31054
rect 16000 31106 16080 31120
rect 16000 31054 16014 31106
rect 16066 31054 16080 31106
rect 16000 31040 16080 31054
rect 16160 31106 16240 31120
rect 16160 31054 16174 31106
rect 16226 31054 16240 31106
rect 16160 31040 16240 31054
rect 16320 31106 16400 31120
rect 16320 31054 16334 31106
rect 16386 31054 16400 31106
rect 16320 31040 16400 31054
rect 16480 31106 16560 31120
rect 16480 31054 16494 31106
rect 16546 31054 16560 31106
rect 16480 31040 16560 31054
rect 16640 31106 16720 31120
rect 16640 31054 16654 31106
rect 16706 31054 16720 31106
rect 16640 31040 16720 31054
rect 16800 31106 16880 31120
rect 16800 31054 16814 31106
rect 16866 31054 16880 31106
rect 16800 31040 16880 31054
rect 16960 31106 17040 31120
rect 16960 31054 16974 31106
rect 17026 31054 17040 31106
rect 16960 31040 17040 31054
rect 17120 31106 17200 31120
rect 17120 31054 17134 31106
rect 17186 31054 17200 31106
rect 17120 31040 17200 31054
rect 17280 31106 17360 31120
rect 17280 31054 17294 31106
rect 17346 31054 17360 31106
rect 17280 31040 17360 31054
rect 17440 31106 17520 31120
rect 17440 31054 17454 31106
rect 17506 31054 17520 31106
rect 17440 31040 17520 31054
rect 17600 31106 17680 31120
rect 17600 31054 17614 31106
rect 17666 31054 17680 31106
rect 17600 31040 17680 31054
rect 17760 31106 17840 31120
rect 17760 31054 17774 31106
rect 17826 31054 17840 31106
rect 17760 31040 17840 31054
rect 17920 31106 18000 31120
rect 17920 31054 17934 31106
rect 17986 31054 18000 31106
rect 17920 31040 18000 31054
rect 18080 31106 18160 31120
rect 18080 31054 18094 31106
rect 18146 31054 18160 31106
rect 18080 31040 18160 31054
rect 18240 31106 18320 31120
rect 18240 31054 18254 31106
rect 18306 31054 18320 31106
rect 18240 31040 18320 31054
rect 18400 31106 18480 31120
rect 18400 31054 18414 31106
rect 18466 31054 18480 31106
rect 18400 31040 18480 31054
rect 18560 31106 18640 31120
rect 18560 31054 18574 31106
rect 18626 31054 18640 31106
rect 18560 31040 18640 31054
rect 18720 31106 18800 31120
rect 18720 31054 18734 31106
rect 18786 31054 18800 31106
rect 18720 31040 18800 31054
rect 18880 31106 18960 31120
rect 18880 31054 18894 31106
rect 18946 31054 18960 31106
rect 18880 31040 18960 31054
rect 23120 31106 23200 31120
rect 23120 31054 23134 31106
rect 23186 31054 23200 31106
rect 23120 31040 23200 31054
rect 23280 31106 23360 31120
rect 23280 31054 23294 31106
rect 23346 31054 23360 31106
rect 23280 31040 23360 31054
rect 23440 31106 23520 31120
rect 23440 31054 23454 31106
rect 23506 31054 23520 31106
rect 23440 31040 23520 31054
rect 23600 31106 23680 31120
rect 23600 31054 23614 31106
rect 23666 31054 23680 31106
rect 23600 31040 23680 31054
rect 23760 31106 23840 31120
rect 23760 31054 23774 31106
rect 23826 31054 23840 31106
rect 23760 31040 23840 31054
rect 23920 31106 24000 31120
rect 23920 31054 23934 31106
rect 23986 31054 24000 31106
rect 23920 31040 24000 31054
rect 24080 31106 24160 31120
rect 24080 31054 24094 31106
rect 24146 31054 24160 31106
rect 24080 31040 24160 31054
rect 24240 31106 24320 31120
rect 24240 31054 24254 31106
rect 24306 31054 24320 31106
rect 24240 31040 24320 31054
rect 24400 31106 24480 31120
rect 24400 31054 24414 31106
rect 24466 31054 24480 31106
rect 24400 31040 24480 31054
rect 24560 31106 24640 31120
rect 24560 31054 24574 31106
rect 24626 31054 24640 31106
rect 24560 31040 24640 31054
rect 24720 31106 24800 31120
rect 24720 31054 24734 31106
rect 24786 31054 24800 31106
rect 24720 31040 24800 31054
rect 24880 31106 24960 31120
rect 24880 31054 24894 31106
rect 24946 31054 24960 31106
rect 24880 31040 24960 31054
rect 25040 31106 25120 31120
rect 25040 31054 25054 31106
rect 25106 31054 25120 31106
rect 25040 31040 25120 31054
rect 25200 31106 25280 31120
rect 25200 31054 25214 31106
rect 25266 31054 25280 31106
rect 25200 31040 25280 31054
rect 25360 31106 25440 31120
rect 25360 31054 25374 31106
rect 25426 31054 25440 31106
rect 25360 31040 25440 31054
rect 25520 31106 25600 31120
rect 25520 31054 25534 31106
rect 25586 31054 25600 31106
rect 25520 31040 25600 31054
rect 25680 31106 25760 31120
rect 25680 31054 25694 31106
rect 25746 31054 25760 31106
rect 25680 31040 25760 31054
rect 25840 31106 25920 31120
rect 25840 31054 25854 31106
rect 25906 31054 25920 31106
rect 25840 31040 25920 31054
rect 26000 31106 26080 31120
rect 26000 31054 26014 31106
rect 26066 31054 26080 31106
rect 26000 31040 26080 31054
rect 26160 31106 26240 31120
rect 26160 31054 26174 31106
rect 26226 31054 26240 31106
rect 26160 31040 26240 31054
rect 26320 31106 26400 31120
rect 26320 31054 26334 31106
rect 26386 31054 26400 31106
rect 26320 31040 26400 31054
rect 26480 31106 26560 31120
rect 26480 31054 26494 31106
rect 26546 31054 26560 31106
rect 26480 31040 26560 31054
rect 26640 31106 26720 31120
rect 26640 31054 26654 31106
rect 26706 31054 26720 31106
rect 26640 31040 26720 31054
rect 26800 31106 26880 31120
rect 26800 31054 26814 31106
rect 26866 31054 26880 31106
rect 26800 31040 26880 31054
rect 26960 31106 27040 31120
rect 26960 31054 26974 31106
rect 27026 31054 27040 31106
rect 26960 31040 27040 31054
rect 27120 31106 27200 31120
rect 27120 31054 27134 31106
rect 27186 31054 27200 31106
rect 27120 31040 27200 31054
rect 27280 31106 27360 31120
rect 27280 31054 27294 31106
rect 27346 31054 27360 31106
rect 27280 31040 27360 31054
rect 27440 31106 27520 31120
rect 27440 31054 27454 31106
rect 27506 31054 27520 31106
rect 27440 31040 27520 31054
rect 27600 31106 27680 31120
rect 27600 31054 27614 31106
rect 27666 31054 27680 31106
rect 27600 31040 27680 31054
rect 27760 31106 27840 31120
rect 27760 31054 27774 31106
rect 27826 31054 27840 31106
rect 27760 31040 27840 31054
rect 27920 31106 28000 31120
rect 27920 31054 27934 31106
rect 27986 31054 28000 31106
rect 27920 31040 28000 31054
rect 28080 31106 28160 31120
rect 28080 31054 28094 31106
rect 28146 31054 28160 31106
rect 28080 31040 28160 31054
rect 28240 31106 28320 31120
rect 28240 31054 28254 31106
rect 28306 31054 28320 31106
rect 28240 31040 28320 31054
rect 28400 31106 28480 31120
rect 28400 31054 28414 31106
rect 28466 31054 28480 31106
rect 28400 31040 28480 31054
rect 28560 31106 28640 31120
rect 28560 31054 28574 31106
rect 28626 31054 28640 31106
rect 28560 31040 28640 31054
rect 28720 31106 28800 31120
rect 28720 31054 28734 31106
rect 28786 31054 28800 31106
rect 28720 31040 28800 31054
rect 28880 31106 28960 31120
rect 28880 31054 28894 31106
rect 28946 31054 28960 31106
rect 28880 31040 28960 31054
rect 29040 31106 29120 31120
rect 29040 31054 29054 31106
rect 29106 31054 29120 31106
rect 29040 31040 29120 31054
rect 29200 31106 29280 31120
rect 29200 31054 29214 31106
rect 29266 31054 29280 31106
rect 29200 31040 29280 31054
rect 29360 31106 29440 31120
rect 29360 31054 29374 31106
rect 29426 31054 29440 31106
rect 29360 31040 29440 31054
rect 33520 31106 33600 31120
rect 33520 31054 33534 31106
rect 33586 31054 33600 31106
rect 33520 31040 33600 31054
rect 33680 31106 33760 31120
rect 33680 31054 33694 31106
rect 33746 31054 33760 31106
rect 33680 31040 33760 31054
rect 33840 31106 33920 31120
rect 33840 31054 33854 31106
rect 33906 31054 33920 31106
rect 33840 31040 33920 31054
rect 34000 31106 34080 31120
rect 34000 31054 34014 31106
rect 34066 31054 34080 31106
rect 34000 31040 34080 31054
rect 34160 31106 34240 31120
rect 34160 31054 34174 31106
rect 34226 31054 34240 31106
rect 34160 31040 34240 31054
rect 34320 31106 34400 31120
rect 34320 31054 34334 31106
rect 34386 31054 34400 31106
rect 34320 31040 34400 31054
rect 34480 31106 34560 31120
rect 34480 31054 34494 31106
rect 34546 31054 34560 31106
rect 34480 31040 34560 31054
rect 34640 31106 34720 31120
rect 34640 31054 34654 31106
rect 34706 31054 34720 31106
rect 34640 31040 34720 31054
rect 34800 31106 34880 31120
rect 34800 31054 34814 31106
rect 34866 31054 34880 31106
rect 34800 31040 34880 31054
rect 34960 31106 35040 31120
rect 34960 31054 34974 31106
rect 35026 31054 35040 31106
rect 34960 31040 35040 31054
rect 35120 31106 35200 31120
rect 35120 31054 35134 31106
rect 35186 31054 35200 31106
rect 35120 31040 35200 31054
rect 35280 31106 35360 31120
rect 35280 31054 35294 31106
rect 35346 31054 35360 31106
rect 35280 31040 35360 31054
rect 35440 31106 35520 31120
rect 35440 31054 35454 31106
rect 35506 31054 35520 31106
rect 35440 31040 35520 31054
rect 35600 31106 35680 31120
rect 35600 31054 35614 31106
rect 35666 31054 35680 31106
rect 35600 31040 35680 31054
rect 35760 31106 35840 31120
rect 35760 31054 35774 31106
rect 35826 31054 35840 31106
rect 35760 31040 35840 31054
rect 35920 31106 36000 31120
rect 35920 31054 35934 31106
rect 35986 31054 36000 31106
rect 35920 31040 36000 31054
rect 36080 31106 36160 31120
rect 36080 31054 36094 31106
rect 36146 31054 36160 31106
rect 36080 31040 36160 31054
rect 36240 31106 36320 31120
rect 36240 31054 36254 31106
rect 36306 31054 36320 31106
rect 36240 31040 36320 31054
rect 36400 31106 36480 31120
rect 36400 31054 36414 31106
rect 36466 31054 36480 31106
rect 36400 31040 36480 31054
rect 36560 31106 36640 31120
rect 36560 31054 36574 31106
rect 36626 31054 36640 31106
rect 36560 31040 36640 31054
rect 36720 31106 36800 31120
rect 36720 31054 36734 31106
rect 36786 31054 36800 31106
rect 36720 31040 36800 31054
rect 36880 31106 36960 31120
rect 36880 31054 36894 31106
rect 36946 31054 36960 31106
rect 36880 31040 36960 31054
rect 37040 31106 37120 31120
rect 37040 31054 37054 31106
rect 37106 31054 37120 31106
rect 37040 31040 37120 31054
rect 37200 31106 37280 31120
rect 37200 31054 37214 31106
rect 37266 31054 37280 31106
rect 37200 31040 37280 31054
rect 37360 31106 37440 31120
rect 37360 31054 37374 31106
rect 37426 31054 37440 31106
rect 37360 31040 37440 31054
rect 37520 31106 37600 31120
rect 37520 31054 37534 31106
rect 37586 31054 37600 31106
rect 37520 31040 37600 31054
rect 37680 31106 37760 31120
rect 37680 31054 37694 31106
rect 37746 31054 37760 31106
rect 37680 31040 37760 31054
rect 37840 31106 37920 31120
rect 37840 31054 37854 31106
rect 37906 31054 37920 31106
rect 37840 31040 37920 31054
rect 38000 31106 38080 31120
rect 38000 31054 38014 31106
rect 38066 31054 38080 31106
rect 38000 31040 38080 31054
rect 38160 31106 38240 31120
rect 38160 31054 38174 31106
rect 38226 31054 38240 31106
rect 38160 31040 38240 31054
rect 38320 31106 38400 31120
rect 38320 31054 38334 31106
rect 38386 31054 38400 31106
rect 38320 31040 38400 31054
rect 38480 31106 38560 31120
rect 38480 31054 38494 31106
rect 38546 31054 38560 31106
rect 38480 31040 38560 31054
rect 38640 31106 38720 31120
rect 38640 31054 38654 31106
rect 38706 31054 38720 31106
rect 38640 31040 38720 31054
rect 38800 31106 38880 31120
rect 38800 31054 38814 31106
rect 38866 31054 38880 31106
rect 38800 31040 38880 31054
rect 38960 31106 39040 31120
rect 38960 31054 38974 31106
rect 39026 31054 39040 31106
rect 38960 31040 39040 31054
rect 39120 31106 39200 31120
rect 39120 31054 39134 31106
rect 39186 31054 39200 31106
rect 39120 31040 39200 31054
rect 39280 31106 39360 31120
rect 39280 31054 39294 31106
rect 39346 31054 39360 31106
rect 39280 31040 39360 31054
rect 39440 31106 39520 31120
rect 39440 31054 39454 31106
rect 39506 31054 39520 31106
rect 39440 31040 39520 31054
rect 39600 31106 39680 31120
rect 39600 31054 39614 31106
rect 39666 31054 39680 31106
rect 39600 31040 39680 31054
rect 39760 31106 39840 31120
rect 39760 31054 39774 31106
rect 39826 31054 39840 31106
rect 39760 31040 39840 31054
rect 39920 31106 40000 31120
rect 39920 31054 39934 31106
rect 39986 31054 40000 31106
rect 39920 31040 40000 31054
rect 40080 31106 40160 31120
rect 40080 31054 40094 31106
rect 40146 31054 40160 31106
rect 40080 31040 40160 31054
rect 40240 31106 40320 31120
rect 40240 31054 40254 31106
rect 40306 31054 40320 31106
rect 40240 31040 40320 31054
rect 40400 31106 40480 31120
rect 40400 31054 40414 31106
rect 40466 31054 40480 31106
rect 40400 31040 40480 31054
rect 40560 31106 40640 31120
rect 40560 31054 40574 31106
rect 40626 31054 40640 31106
rect 40560 31040 40640 31054
rect 40720 31106 40800 31120
rect 40720 31054 40734 31106
rect 40786 31054 40800 31106
rect 40720 31040 40800 31054
rect 40880 31106 40960 31120
rect 40880 31054 40894 31106
rect 40946 31054 40960 31106
rect 40880 31040 40960 31054
rect 41040 31106 41120 31120
rect 41040 31054 41054 31106
rect 41106 31054 41120 31106
rect 41040 31040 41120 31054
rect 41200 31106 41280 31120
rect 41200 31054 41214 31106
rect 41266 31054 41280 31106
rect 41200 31040 41280 31054
rect 41360 31106 41440 31120
rect 41360 31054 41374 31106
rect 41426 31054 41440 31106
rect 41360 31040 41440 31054
rect 41520 31106 41600 31120
rect 41520 31054 41534 31106
rect 41586 31054 41600 31106
rect 41520 31040 41600 31054
rect 41680 31106 41760 31120
rect 41680 31054 41694 31106
rect 41746 31054 41760 31106
rect 41680 31040 41760 31054
rect 41840 31106 41920 31120
rect 41840 31054 41854 31106
rect 41906 31054 41920 31106
rect 41840 31040 41920 31054
rect 0 30786 80 30800
rect 0 30734 14 30786
rect 66 30734 80 30786
rect 0 30720 80 30734
rect 160 30786 240 30800
rect 160 30734 174 30786
rect 226 30734 240 30786
rect 160 30720 240 30734
rect 320 30786 400 30800
rect 320 30734 334 30786
rect 386 30734 400 30786
rect 320 30720 400 30734
rect 480 30786 560 30800
rect 480 30734 494 30786
rect 546 30734 560 30786
rect 480 30720 560 30734
rect 640 30786 720 30800
rect 640 30734 654 30786
rect 706 30734 720 30786
rect 640 30720 720 30734
rect 800 30786 880 30800
rect 800 30734 814 30786
rect 866 30734 880 30786
rect 800 30720 880 30734
rect 960 30786 1040 30800
rect 960 30734 974 30786
rect 1026 30734 1040 30786
rect 960 30720 1040 30734
rect 1120 30786 1200 30800
rect 1120 30734 1134 30786
rect 1186 30734 1200 30786
rect 1120 30720 1200 30734
rect 1280 30786 1360 30800
rect 1280 30734 1294 30786
rect 1346 30734 1360 30786
rect 1280 30720 1360 30734
rect 1440 30786 1520 30800
rect 1440 30734 1454 30786
rect 1506 30734 1520 30786
rect 1440 30720 1520 30734
rect 1600 30786 1680 30800
rect 1600 30734 1614 30786
rect 1666 30734 1680 30786
rect 1600 30720 1680 30734
rect 1760 30786 1840 30800
rect 1760 30734 1774 30786
rect 1826 30734 1840 30786
rect 1760 30720 1840 30734
rect 1920 30786 2000 30800
rect 1920 30734 1934 30786
rect 1986 30734 2000 30786
rect 1920 30720 2000 30734
rect 2080 30786 2160 30800
rect 2080 30734 2094 30786
rect 2146 30734 2160 30786
rect 2080 30720 2160 30734
rect 2240 30786 2320 30800
rect 2240 30734 2254 30786
rect 2306 30734 2320 30786
rect 2240 30720 2320 30734
rect 2400 30786 2480 30800
rect 2400 30734 2414 30786
rect 2466 30734 2480 30786
rect 2400 30720 2480 30734
rect 2560 30786 2640 30800
rect 2560 30734 2574 30786
rect 2626 30734 2640 30786
rect 2560 30720 2640 30734
rect 2720 30786 2800 30800
rect 2720 30734 2734 30786
rect 2786 30734 2800 30786
rect 2720 30720 2800 30734
rect 2880 30786 2960 30800
rect 2880 30734 2894 30786
rect 2946 30734 2960 30786
rect 2880 30720 2960 30734
rect 3040 30786 3120 30800
rect 3040 30734 3054 30786
rect 3106 30734 3120 30786
rect 3040 30720 3120 30734
rect 3200 30786 3280 30800
rect 3200 30734 3214 30786
rect 3266 30734 3280 30786
rect 3200 30720 3280 30734
rect 3360 30786 3440 30800
rect 3360 30734 3374 30786
rect 3426 30734 3440 30786
rect 3360 30720 3440 30734
rect 3520 30786 3600 30800
rect 3520 30734 3534 30786
rect 3586 30734 3600 30786
rect 3520 30720 3600 30734
rect 3680 30786 3760 30800
rect 3680 30734 3694 30786
rect 3746 30734 3760 30786
rect 3680 30720 3760 30734
rect 3840 30786 3920 30800
rect 3840 30734 3854 30786
rect 3906 30734 3920 30786
rect 3840 30720 3920 30734
rect 4000 30786 4080 30800
rect 4000 30734 4014 30786
rect 4066 30734 4080 30786
rect 4000 30720 4080 30734
rect 4160 30786 4240 30800
rect 4160 30734 4174 30786
rect 4226 30734 4240 30786
rect 4160 30720 4240 30734
rect 4320 30786 4400 30800
rect 4320 30734 4334 30786
rect 4386 30734 4400 30786
rect 4320 30720 4400 30734
rect 4480 30786 4560 30800
rect 4480 30734 4494 30786
rect 4546 30734 4560 30786
rect 4480 30720 4560 30734
rect 4640 30786 4720 30800
rect 4640 30734 4654 30786
rect 4706 30734 4720 30786
rect 4640 30720 4720 30734
rect 4800 30786 4880 30800
rect 4800 30734 4814 30786
rect 4866 30734 4880 30786
rect 4800 30720 4880 30734
rect 4960 30786 5040 30800
rect 4960 30734 4974 30786
rect 5026 30734 5040 30786
rect 4960 30720 5040 30734
rect 5120 30786 5200 30800
rect 5120 30734 5134 30786
rect 5186 30734 5200 30786
rect 5120 30720 5200 30734
rect 5280 30786 5360 30800
rect 5280 30734 5294 30786
rect 5346 30734 5360 30786
rect 5280 30720 5360 30734
rect 5440 30786 5520 30800
rect 5440 30734 5454 30786
rect 5506 30734 5520 30786
rect 5440 30720 5520 30734
rect 5600 30786 5680 30800
rect 5600 30734 5614 30786
rect 5666 30734 5680 30786
rect 5600 30720 5680 30734
rect 5760 30786 5840 30800
rect 5760 30734 5774 30786
rect 5826 30734 5840 30786
rect 5760 30720 5840 30734
rect 5920 30786 6000 30800
rect 5920 30734 5934 30786
rect 5986 30734 6000 30786
rect 5920 30720 6000 30734
rect 6080 30786 6160 30800
rect 6080 30734 6094 30786
rect 6146 30734 6160 30786
rect 6080 30720 6160 30734
rect 6240 30786 6320 30800
rect 6240 30734 6254 30786
rect 6306 30734 6320 30786
rect 6240 30720 6320 30734
rect 6400 30786 6480 30800
rect 6400 30734 6414 30786
rect 6466 30734 6480 30786
rect 6400 30720 6480 30734
rect 6560 30786 6640 30800
rect 6560 30734 6574 30786
rect 6626 30734 6640 30786
rect 6560 30720 6640 30734
rect 6720 30786 6800 30800
rect 6720 30734 6734 30786
rect 6786 30734 6800 30786
rect 6720 30720 6800 30734
rect 6880 30786 6960 30800
rect 6880 30734 6894 30786
rect 6946 30734 6960 30786
rect 6880 30720 6960 30734
rect 7040 30786 7120 30800
rect 7040 30734 7054 30786
rect 7106 30734 7120 30786
rect 7040 30720 7120 30734
rect 7200 30786 7280 30800
rect 7200 30734 7214 30786
rect 7266 30734 7280 30786
rect 7200 30720 7280 30734
rect 7360 30786 7440 30800
rect 7360 30734 7374 30786
rect 7426 30734 7440 30786
rect 7360 30720 7440 30734
rect 7520 30786 7600 30800
rect 7520 30734 7534 30786
rect 7586 30734 7600 30786
rect 7520 30720 7600 30734
rect 7680 30786 7760 30800
rect 7680 30734 7694 30786
rect 7746 30734 7760 30786
rect 7680 30720 7760 30734
rect 7840 30786 7920 30800
rect 7840 30734 7854 30786
rect 7906 30734 7920 30786
rect 7840 30720 7920 30734
rect 8000 30786 8080 30800
rect 8000 30734 8014 30786
rect 8066 30734 8080 30786
rect 8000 30720 8080 30734
rect 8160 30786 8240 30800
rect 8160 30734 8174 30786
rect 8226 30734 8240 30786
rect 8160 30720 8240 30734
rect 8320 30786 8400 30800
rect 8320 30734 8334 30786
rect 8386 30734 8400 30786
rect 8320 30720 8400 30734
rect 12480 30786 12560 30800
rect 12480 30734 12494 30786
rect 12546 30734 12560 30786
rect 12480 30720 12560 30734
rect 12640 30786 12720 30800
rect 12640 30734 12654 30786
rect 12706 30734 12720 30786
rect 12640 30720 12720 30734
rect 12800 30786 12880 30800
rect 12800 30734 12814 30786
rect 12866 30734 12880 30786
rect 12800 30720 12880 30734
rect 12960 30786 13040 30800
rect 12960 30734 12974 30786
rect 13026 30734 13040 30786
rect 12960 30720 13040 30734
rect 13120 30786 13200 30800
rect 13120 30734 13134 30786
rect 13186 30734 13200 30786
rect 13120 30720 13200 30734
rect 13280 30786 13360 30800
rect 13280 30734 13294 30786
rect 13346 30734 13360 30786
rect 13280 30720 13360 30734
rect 13440 30786 13520 30800
rect 13440 30734 13454 30786
rect 13506 30734 13520 30786
rect 13440 30720 13520 30734
rect 13600 30786 13680 30800
rect 13600 30734 13614 30786
rect 13666 30734 13680 30786
rect 13600 30720 13680 30734
rect 13760 30786 13840 30800
rect 13760 30734 13774 30786
rect 13826 30734 13840 30786
rect 13760 30720 13840 30734
rect 13920 30786 14000 30800
rect 13920 30734 13934 30786
rect 13986 30734 14000 30786
rect 13920 30720 14000 30734
rect 14080 30786 14160 30800
rect 14080 30734 14094 30786
rect 14146 30734 14160 30786
rect 14080 30720 14160 30734
rect 14240 30786 14320 30800
rect 14240 30734 14254 30786
rect 14306 30734 14320 30786
rect 14240 30720 14320 30734
rect 14400 30786 14480 30800
rect 14400 30734 14414 30786
rect 14466 30734 14480 30786
rect 14400 30720 14480 30734
rect 14560 30786 14640 30800
rect 14560 30734 14574 30786
rect 14626 30734 14640 30786
rect 14560 30720 14640 30734
rect 14720 30786 14800 30800
rect 14720 30734 14734 30786
rect 14786 30734 14800 30786
rect 14720 30720 14800 30734
rect 14880 30786 14960 30800
rect 14880 30734 14894 30786
rect 14946 30734 14960 30786
rect 14880 30720 14960 30734
rect 15040 30786 15120 30800
rect 15040 30734 15054 30786
rect 15106 30734 15120 30786
rect 15040 30720 15120 30734
rect 15200 30786 15280 30800
rect 15200 30734 15214 30786
rect 15266 30734 15280 30786
rect 15200 30720 15280 30734
rect 15360 30786 15440 30800
rect 15360 30734 15374 30786
rect 15426 30734 15440 30786
rect 15360 30720 15440 30734
rect 15520 30786 15600 30800
rect 15520 30734 15534 30786
rect 15586 30734 15600 30786
rect 15520 30720 15600 30734
rect 15680 30786 15760 30800
rect 15680 30734 15694 30786
rect 15746 30734 15760 30786
rect 15680 30720 15760 30734
rect 15840 30786 15920 30800
rect 15840 30734 15854 30786
rect 15906 30734 15920 30786
rect 15840 30720 15920 30734
rect 16000 30786 16080 30800
rect 16000 30734 16014 30786
rect 16066 30734 16080 30786
rect 16000 30720 16080 30734
rect 16160 30786 16240 30800
rect 16160 30734 16174 30786
rect 16226 30734 16240 30786
rect 16160 30720 16240 30734
rect 16320 30786 16400 30800
rect 16320 30734 16334 30786
rect 16386 30734 16400 30786
rect 16320 30720 16400 30734
rect 16480 30786 16560 30800
rect 16480 30734 16494 30786
rect 16546 30734 16560 30786
rect 16480 30720 16560 30734
rect 16640 30786 16720 30800
rect 16640 30734 16654 30786
rect 16706 30734 16720 30786
rect 16640 30720 16720 30734
rect 16800 30786 16880 30800
rect 16800 30734 16814 30786
rect 16866 30734 16880 30786
rect 16800 30720 16880 30734
rect 16960 30786 17040 30800
rect 16960 30734 16974 30786
rect 17026 30734 17040 30786
rect 16960 30720 17040 30734
rect 17120 30786 17200 30800
rect 17120 30734 17134 30786
rect 17186 30734 17200 30786
rect 17120 30720 17200 30734
rect 17280 30786 17360 30800
rect 17280 30734 17294 30786
rect 17346 30734 17360 30786
rect 17280 30720 17360 30734
rect 17440 30786 17520 30800
rect 17440 30734 17454 30786
rect 17506 30734 17520 30786
rect 17440 30720 17520 30734
rect 17600 30786 17680 30800
rect 17600 30734 17614 30786
rect 17666 30734 17680 30786
rect 17600 30720 17680 30734
rect 17760 30786 17840 30800
rect 17760 30734 17774 30786
rect 17826 30734 17840 30786
rect 17760 30720 17840 30734
rect 17920 30786 18000 30800
rect 17920 30734 17934 30786
rect 17986 30734 18000 30786
rect 17920 30720 18000 30734
rect 18080 30786 18160 30800
rect 18080 30734 18094 30786
rect 18146 30734 18160 30786
rect 18080 30720 18160 30734
rect 18240 30786 18320 30800
rect 18240 30734 18254 30786
rect 18306 30734 18320 30786
rect 18240 30720 18320 30734
rect 18400 30786 18480 30800
rect 18400 30734 18414 30786
rect 18466 30734 18480 30786
rect 18400 30720 18480 30734
rect 18560 30786 18640 30800
rect 18560 30734 18574 30786
rect 18626 30734 18640 30786
rect 18560 30720 18640 30734
rect 18720 30786 18800 30800
rect 18720 30734 18734 30786
rect 18786 30734 18800 30786
rect 18720 30720 18800 30734
rect 18880 30786 18960 30800
rect 18880 30734 18894 30786
rect 18946 30734 18960 30786
rect 18880 30720 18960 30734
rect 23120 30786 23200 30800
rect 23120 30734 23134 30786
rect 23186 30734 23200 30786
rect 23120 30720 23200 30734
rect 23280 30786 23360 30800
rect 23280 30734 23294 30786
rect 23346 30734 23360 30786
rect 23280 30720 23360 30734
rect 23440 30786 23520 30800
rect 23440 30734 23454 30786
rect 23506 30734 23520 30786
rect 23440 30720 23520 30734
rect 23600 30786 23680 30800
rect 23600 30734 23614 30786
rect 23666 30734 23680 30786
rect 23600 30720 23680 30734
rect 23760 30786 23840 30800
rect 23760 30734 23774 30786
rect 23826 30734 23840 30786
rect 23760 30720 23840 30734
rect 23920 30786 24000 30800
rect 23920 30734 23934 30786
rect 23986 30734 24000 30786
rect 23920 30720 24000 30734
rect 24080 30786 24160 30800
rect 24080 30734 24094 30786
rect 24146 30734 24160 30786
rect 24080 30720 24160 30734
rect 24240 30786 24320 30800
rect 24240 30734 24254 30786
rect 24306 30734 24320 30786
rect 24240 30720 24320 30734
rect 24400 30786 24480 30800
rect 24400 30734 24414 30786
rect 24466 30734 24480 30786
rect 24400 30720 24480 30734
rect 24560 30786 24640 30800
rect 24560 30734 24574 30786
rect 24626 30734 24640 30786
rect 24560 30720 24640 30734
rect 24720 30786 24800 30800
rect 24720 30734 24734 30786
rect 24786 30734 24800 30786
rect 24720 30720 24800 30734
rect 24880 30786 24960 30800
rect 24880 30734 24894 30786
rect 24946 30734 24960 30786
rect 24880 30720 24960 30734
rect 25040 30786 25120 30800
rect 25040 30734 25054 30786
rect 25106 30734 25120 30786
rect 25040 30720 25120 30734
rect 25200 30786 25280 30800
rect 25200 30734 25214 30786
rect 25266 30734 25280 30786
rect 25200 30720 25280 30734
rect 25360 30786 25440 30800
rect 25360 30734 25374 30786
rect 25426 30734 25440 30786
rect 25360 30720 25440 30734
rect 25520 30786 25600 30800
rect 25520 30734 25534 30786
rect 25586 30734 25600 30786
rect 25520 30720 25600 30734
rect 25680 30786 25760 30800
rect 25680 30734 25694 30786
rect 25746 30734 25760 30786
rect 25680 30720 25760 30734
rect 25840 30786 25920 30800
rect 25840 30734 25854 30786
rect 25906 30734 25920 30786
rect 25840 30720 25920 30734
rect 26000 30786 26080 30800
rect 26000 30734 26014 30786
rect 26066 30734 26080 30786
rect 26000 30720 26080 30734
rect 26160 30786 26240 30800
rect 26160 30734 26174 30786
rect 26226 30734 26240 30786
rect 26160 30720 26240 30734
rect 26320 30786 26400 30800
rect 26320 30734 26334 30786
rect 26386 30734 26400 30786
rect 26320 30720 26400 30734
rect 26480 30786 26560 30800
rect 26480 30734 26494 30786
rect 26546 30734 26560 30786
rect 26480 30720 26560 30734
rect 26640 30786 26720 30800
rect 26640 30734 26654 30786
rect 26706 30734 26720 30786
rect 26640 30720 26720 30734
rect 26800 30786 26880 30800
rect 26800 30734 26814 30786
rect 26866 30734 26880 30786
rect 26800 30720 26880 30734
rect 26960 30786 27040 30800
rect 26960 30734 26974 30786
rect 27026 30734 27040 30786
rect 26960 30720 27040 30734
rect 27120 30786 27200 30800
rect 27120 30734 27134 30786
rect 27186 30734 27200 30786
rect 27120 30720 27200 30734
rect 27280 30786 27360 30800
rect 27280 30734 27294 30786
rect 27346 30734 27360 30786
rect 27280 30720 27360 30734
rect 27440 30786 27520 30800
rect 27440 30734 27454 30786
rect 27506 30734 27520 30786
rect 27440 30720 27520 30734
rect 27600 30786 27680 30800
rect 27600 30734 27614 30786
rect 27666 30734 27680 30786
rect 27600 30720 27680 30734
rect 27760 30786 27840 30800
rect 27760 30734 27774 30786
rect 27826 30734 27840 30786
rect 27760 30720 27840 30734
rect 27920 30786 28000 30800
rect 27920 30734 27934 30786
rect 27986 30734 28000 30786
rect 27920 30720 28000 30734
rect 28080 30786 28160 30800
rect 28080 30734 28094 30786
rect 28146 30734 28160 30786
rect 28080 30720 28160 30734
rect 28240 30786 28320 30800
rect 28240 30734 28254 30786
rect 28306 30734 28320 30786
rect 28240 30720 28320 30734
rect 28400 30786 28480 30800
rect 28400 30734 28414 30786
rect 28466 30734 28480 30786
rect 28400 30720 28480 30734
rect 28560 30786 28640 30800
rect 28560 30734 28574 30786
rect 28626 30734 28640 30786
rect 28560 30720 28640 30734
rect 28720 30786 28800 30800
rect 28720 30734 28734 30786
rect 28786 30734 28800 30786
rect 28720 30720 28800 30734
rect 28880 30786 28960 30800
rect 28880 30734 28894 30786
rect 28946 30734 28960 30786
rect 28880 30720 28960 30734
rect 29040 30786 29120 30800
rect 29040 30734 29054 30786
rect 29106 30734 29120 30786
rect 29040 30720 29120 30734
rect 29200 30786 29280 30800
rect 29200 30734 29214 30786
rect 29266 30734 29280 30786
rect 29200 30720 29280 30734
rect 29360 30786 29440 30800
rect 29360 30734 29374 30786
rect 29426 30734 29440 30786
rect 29360 30720 29440 30734
rect 33520 30786 33600 30800
rect 33520 30734 33534 30786
rect 33586 30734 33600 30786
rect 33520 30720 33600 30734
rect 33680 30786 33760 30800
rect 33680 30734 33694 30786
rect 33746 30734 33760 30786
rect 33680 30720 33760 30734
rect 33840 30786 33920 30800
rect 33840 30734 33854 30786
rect 33906 30734 33920 30786
rect 33840 30720 33920 30734
rect 34000 30786 34080 30800
rect 34000 30734 34014 30786
rect 34066 30734 34080 30786
rect 34000 30720 34080 30734
rect 34160 30786 34240 30800
rect 34160 30734 34174 30786
rect 34226 30734 34240 30786
rect 34160 30720 34240 30734
rect 34320 30786 34400 30800
rect 34320 30734 34334 30786
rect 34386 30734 34400 30786
rect 34320 30720 34400 30734
rect 34480 30786 34560 30800
rect 34480 30734 34494 30786
rect 34546 30734 34560 30786
rect 34480 30720 34560 30734
rect 34640 30786 34720 30800
rect 34640 30734 34654 30786
rect 34706 30734 34720 30786
rect 34640 30720 34720 30734
rect 34800 30786 34880 30800
rect 34800 30734 34814 30786
rect 34866 30734 34880 30786
rect 34800 30720 34880 30734
rect 34960 30786 35040 30800
rect 34960 30734 34974 30786
rect 35026 30734 35040 30786
rect 34960 30720 35040 30734
rect 35120 30786 35200 30800
rect 35120 30734 35134 30786
rect 35186 30734 35200 30786
rect 35120 30720 35200 30734
rect 35280 30786 35360 30800
rect 35280 30734 35294 30786
rect 35346 30734 35360 30786
rect 35280 30720 35360 30734
rect 35440 30786 35520 30800
rect 35440 30734 35454 30786
rect 35506 30734 35520 30786
rect 35440 30720 35520 30734
rect 35600 30786 35680 30800
rect 35600 30734 35614 30786
rect 35666 30734 35680 30786
rect 35600 30720 35680 30734
rect 35760 30786 35840 30800
rect 35760 30734 35774 30786
rect 35826 30734 35840 30786
rect 35760 30720 35840 30734
rect 35920 30786 36000 30800
rect 35920 30734 35934 30786
rect 35986 30734 36000 30786
rect 35920 30720 36000 30734
rect 36080 30786 36160 30800
rect 36080 30734 36094 30786
rect 36146 30734 36160 30786
rect 36080 30720 36160 30734
rect 36240 30786 36320 30800
rect 36240 30734 36254 30786
rect 36306 30734 36320 30786
rect 36240 30720 36320 30734
rect 36400 30786 36480 30800
rect 36400 30734 36414 30786
rect 36466 30734 36480 30786
rect 36400 30720 36480 30734
rect 36560 30786 36640 30800
rect 36560 30734 36574 30786
rect 36626 30734 36640 30786
rect 36560 30720 36640 30734
rect 36720 30786 36800 30800
rect 36720 30734 36734 30786
rect 36786 30734 36800 30786
rect 36720 30720 36800 30734
rect 36880 30786 36960 30800
rect 36880 30734 36894 30786
rect 36946 30734 36960 30786
rect 36880 30720 36960 30734
rect 37040 30786 37120 30800
rect 37040 30734 37054 30786
rect 37106 30734 37120 30786
rect 37040 30720 37120 30734
rect 37200 30786 37280 30800
rect 37200 30734 37214 30786
rect 37266 30734 37280 30786
rect 37200 30720 37280 30734
rect 37360 30786 37440 30800
rect 37360 30734 37374 30786
rect 37426 30734 37440 30786
rect 37360 30720 37440 30734
rect 37520 30786 37600 30800
rect 37520 30734 37534 30786
rect 37586 30734 37600 30786
rect 37520 30720 37600 30734
rect 37680 30786 37760 30800
rect 37680 30734 37694 30786
rect 37746 30734 37760 30786
rect 37680 30720 37760 30734
rect 37840 30786 37920 30800
rect 37840 30734 37854 30786
rect 37906 30734 37920 30786
rect 37840 30720 37920 30734
rect 38000 30786 38080 30800
rect 38000 30734 38014 30786
rect 38066 30734 38080 30786
rect 38000 30720 38080 30734
rect 38160 30786 38240 30800
rect 38160 30734 38174 30786
rect 38226 30734 38240 30786
rect 38160 30720 38240 30734
rect 38320 30786 38400 30800
rect 38320 30734 38334 30786
rect 38386 30734 38400 30786
rect 38320 30720 38400 30734
rect 38480 30786 38560 30800
rect 38480 30734 38494 30786
rect 38546 30734 38560 30786
rect 38480 30720 38560 30734
rect 38640 30786 38720 30800
rect 38640 30734 38654 30786
rect 38706 30734 38720 30786
rect 38640 30720 38720 30734
rect 38800 30786 38880 30800
rect 38800 30734 38814 30786
rect 38866 30734 38880 30786
rect 38800 30720 38880 30734
rect 38960 30786 39040 30800
rect 38960 30734 38974 30786
rect 39026 30734 39040 30786
rect 38960 30720 39040 30734
rect 39120 30786 39200 30800
rect 39120 30734 39134 30786
rect 39186 30734 39200 30786
rect 39120 30720 39200 30734
rect 39280 30786 39360 30800
rect 39280 30734 39294 30786
rect 39346 30734 39360 30786
rect 39280 30720 39360 30734
rect 39440 30786 39520 30800
rect 39440 30734 39454 30786
rect 39506 30734 39520 30786
rect 39440 30720 39520 30734
rect 39600 30786 39680 30800
rect 39600 30734 39614 30786
rect 39666 30734 39680 30786
rect 39600 30720 39680 30734
rect 39760 30786 39840 30800
rect 39760 30734 39774 30786
rect 39826 30734 39840 30786
rect 39760 30720 39840 30734
rect 39920 30786 40000 30800
rect 39920 30734 39934 30786
rect 39986 30734 40000 30786
rect 39920 30720 40000 30734
rect 40080 30786 40160 30800
rect 40080 30734 40094 30786
rect 40146 30734 40160 30786
rect 40080 30720 40160 30734
rect 40240 30786 40320 30800
rect 40240 30734 40254 30786
rect 40306 30734 40320 30786
rect 40240 30720 40320 30734
rect 40400 30786 40480 30800
rect 40400 30734 40414 30786
rect 40466 30734 40480 30786
rect 40400 30720 40480 30734
rect 40560 30786 40640 30800
rect 40560 30734 40574 30786
rect 40626 30734 40640 30786
rect 40560 30720 40640 30734
rect 40720 30786 40800 30800
rect 40720 30734 40734 30786
rect 40786 30734 40800 30786
rect 40720 30720 40800 30734
rect 40880 30786 40960 30800
rect 40880 30734 40894 30786
rect 40946 30734 40960 30786
rect 40880 30720 40960 30734
rect 41040 30786 41120 30800
rect 41040 30734 41054 30786
rect 41106 30734 41120 30786
rect 41040 30720 41120 30734
rect 41200 30786 41280 30800
rect 41200 30734 41214 30786
rect 41266 30734 41280 30786
rect 41200 30720 41280 30734
rect 41360 30786 41440 30800
rect 41360 30734 41374 30786
rect 41426 30734 41440 30786
rect 41360 30720 41440 30734
rect 41520 30786 41600 30800
rect 41520 30734 41534 30786
rect 41586 30734 41600 30786
rect 41520 30720 41600 30734
rect 41680 30786 41760 30800
rect 41680 30734 41694 30786
rect 41746 30734 41760 30786
rect 41680 30720 41760 30734
rect 41840 30786 41920 30800
rect 41840 30734 41854 30786
rect 41906 30734 41920 30786
rect 41840 30720 41920 30734
rect 0 30466 80 30480
rect 0 30414 14 30466
rect 66 30414 80 30466
rect 0 30400 80 30414
rect 160 30466 240 30480
rect 160 30414 174 30466
rect 226 30414 240 30466
rect 160 30400 240 30414
rect 320 30466 400 30480
rect 320 30414 334 30466
rect 386 30414 400 30466
rect 320 30400 400 30414
rect 480 30466 560 30480
rect 480 30414 494 30466
rect 546 30414 560 30466
rect 480 30400 560 30414
rect 640 30466 720 30480
rect 640 30414 654 30466
rect 706 30414 720 30466
rect 640 30400 720 30414
rect 800 30466 880 30480
rect 800 30414 814 30466
rect 866 30414 880 30466
rect 800 30400 880 30414
rect 960 30466 1040 30480
rect 960 30414 974 30466
rect 1026 30414 1040 30466
rect 960 30400 1040 30414
rect 1120 30466 1200 30480
rect 1120 30414 1134 30466
rect 1186 30414 1200 30466
rect 1120 30400 1200 30414
rect 1280 30466 1360 30480
rect 1280 30414 1294 30466
rect 1346 30414 1360 30466
rect 1280 30400 1360 30414
rect 1440 30466 1520 30480
rect 1440 30414 1454 30466
rect 1506 30414 1520 30466
rect 1440 30400 1520 30414
rect 1600 30466 1680 30480
rect 1600 30414 1614 30466
rect 1666 30414 1680 30466
rect 1600 30400 1680 30414
rect 1760 30466 1840 30480
rect 1760 30414 1774 30466
rect 1826 30414 1840 30466
rect 1760 30400 1840 30414
rect 1920 30466 2000 30480
rect 1920 30414 1934 30466
rect 1986 30414 2000 30466
rect 1920 30400 2000 30414
rect 2080 30466 2160 30480
rect 2080 30414 2094 30466
rect 2146 30414 2160 30466
rect 2080 30400 2160 30414
rect 2240 30466 2320 30480
rect 2240 30414 2254 30466
rect 2306 30414 2320 30466
rect 2240 30400 2320 30414
rect 2400 30466 2480 30480
rect 2400 30414 2414 30466
rect 2466 30414 2480 30466
rect 2400 30400 2480 30414
rect 2560 30466 2640 30480
rect 2560 30414 2574 30466
rect 2626 30414 2640 30466
rect 2560 30400 2640 30414
rect 2720 30466 2800 30480
rect 2720 30414 2734 30466
rect 2786 30414 2800 30466
rect 2720 30400 2800 30414
rect 2880 30466 2960 30480
rect 2880 30414 2894 30466
rect 2946 30414 2960 30466
rect 2880 30400 2960 30414
rect 3040 30466 3120 30480
rect 3040 30414 3054 30466
rect 3106 30414 3120 30466
rect 3040 30400 3120 30414
rect 3200 30466 3280 30480
rect 3200 30414 3214 30466
rect 3266 30414 3280 30466
rect 3200 30400 3280 30414
rect 3360 30466 3440 30480
rect 3360 30414 3374 30466
rect 3426 30414 3440 30466
rect 3360 30400 3440 30414
rect 3520 30466 3600 30480
rect 3520 30414 3534 30466
rect 3586 30414 3600 30466
rect 3520 30400 3600 30414
rect 3680 30466 3760 30480
rect 3680 30414 3694 30466
rect 3746 30414 3760 30466
rect 3680 30400 3760 30414
rect 3840 30466 3920 30480
rect 3840 30414 3854 30466
rect 3906 30414 3920 30466
rect 3840 30400 3920 30414
rect 4000 30466 4080 30480
rect 4000 30414 4014 30466
rect 4066 30414 4080 30466
rect 4000 30400 4080 30414
rect 4160 30466 4240 30480
rect 4160 30414 4174 30466
rect 4226 30414 4240 30466
rect 4160 30400 4240 30414
rect 4320 30466 4400 30480
rect 4320 30414 4334 30466
rect 4386 30414 4400 30466
rect 4320 30400 4400 30414
rect 4480 30466 4560 30480
rect 4480 30414 4494 30466
rect 4546 30414 4560 30466
rect 4480 30400 4560 30414
rect 4640 30466 4720 30480
rect 4640 30414 4654 30466
rect 4706 30414 4720 30466
rect 4640 30400 4720 30414
rect 4800 30466 4880 30480
rect 4800 30414 4814 30466
rect 4866 30414 4880 30466
rect 4800 30400 4880 30414
rect 4960 30466 5040 30480
rect 4960 30414 4974 30466
rect 5026 30414 5040 30466
rect 4960 30400 5040 30414
rect 5120 30466 5200 30480
rect 5120 30414 5134 30466
rect 5186 30414 5200 30466
rect 5120 30400 5200 30414
rect 5280 30466 5360 30480
rect 5280 30414 5294 30466
rect 5346 30414 5360 30466
rect 5280 30400 5360 30414
rect 5440 30466 5520 30480
rect 5440 30414 5454 30466
rect 5506 30414 5520 30466
rect 5440 30400 5520 30414
rect 5600 30466 5680 30480
rect 5600 30414 5614 30466
rect 5666 30414 5680 30466
rect 5600 30400 5680 30414
rect 5760 30466 5840 30480
rect 5760 30414 5774 30466
rect 5826 30414 5840 30466
rect 5760 30400 5840 30414
rect 5920 30466 6000 30480
rect 5920 30414 5934 30466
rect 5986 30414 6000 30466
rect 5920 30400 6000 30414
rect 6080 30466 6160 30480
rect 6080 30414 6094 30466
rect 6146 30414 6160 30466
rect 6080 30400 6160 30414
rect 6240 30466 6320 30480
rect 6240 30414 6254 30466
rect 6306 30414 6320 30466
rect 6240 30400 6320 30414
rect 6400 30466 6480 30480
rect 6400 30414 6414 30466
rect 6466 30414 6480 30466
rect 6400 30400 6480 30414
rect 6560 30466 6640 30480
rect 6560 30414 6574 30466
rect 6626 30414 6640 30466
rect 6560 30400 6640 30414
rect 6720 30466 6800 30480
rect 6720 30414 6734 30466
rect 6786 30414 6800 30466
rect 6720 30400 6800 30414
rect 6880 30466 6960 30480
rect 6880 30414 6894 30466
rect 6946 30414 6960 30466
rect 6880 30400 6960 30414
rect 7040 30466 7120 30480
rect 7040 30414 7054 30466
rect 7106 30414 7120 30466
rect 7040 30400 7120 30414
rect 7200 30466 7280 30480
rect 7200 30414 7214 30466
rect 7266 30414 7280 30466
rect 7200 30400 7280 30414
rect 7360 30466 7440 30480
rect 7360 30414 7374 30466
rect 7426 30414 7440 30466
rect 7360 30400 7440 30414
rect 7520 30466 7600 30480
rect 7520 30414 7534 30466
rect 7586 30414 7600 30466
rect 7520 30400 7600 30414
rect 7680 30466 7760 30480
rect 7680 30414 7694 30466
rect 7746 30414 7760 30466
rect 7680 30400 7760 30414
rect 7840 30466 7920 30480
rect 7840 30414 7854 30466
rect 7906 30414 7920 30466
rect 7840 30400 7920 30414
rect 8000 30466 8080 30480
rect 8000 30414 8014 30466
rect 8066 30414 8080 30466
rect 8000 30400 8080 30414
rect 8160 30466 8240 30480
rect 8160 30414 8174 30466
rect 8226 30414 8240 30466
rect 8160 30400 8240 30414
rect 8320 30466 8400 30480
rect 8320 30414 8334 30466
rect 8386 30414 8400 30466
rect 8320 30400 8400 30414
rect 12480 30466 12560 30480
rect 12480 30414 12494 30466
rect 12546 30414 12560 30466
rect 12480 30400 12560 30414
rect 12640 30466 12720 30480
rect 12640 30414 12654 30466
rect 12706 30414 12720 30466
rect 12640 30400 12720 30414
rect 12800 30466 12880 30480
rect 12800 30414 12814 30466
rect 12866 30414 12880 30466
rect 12800 30400 12880 30414
rect 12960 30466 13040 30480
rect 12960 30414 12974 30466
rect 13026 30414 13040 30466
rect 12960 30400 13040 30414
rect 13120 30466 13200 30480
rect 13120 30414 13134 30466
rect 13186 30414 13200 30466
rect 13120 30400 13200 30414
rect 13280 30466 13360 30480
rect 13280 30414 13294 30466
rect 13346 30414 13360 30466
rect 13280 30400 13360 30414
rect 13440 30466 13520 30480
rect 13440 30414 13454 30466
rect 13506 30414 13520 30466
rect 13440 30400 13520 30414
rect 13600 30466 13680 30480
rect 13600 30414 13614 30466
rect 13666 30414 13680 30466
rect 13600 30400 13680 30414
rect 13760 30466 13840 30480
rect 13760 30414 13774 30466
rect 13826 30414 13840 30466
rect 13760 30400 13840 30414
rect 13920 30466 14000 30480
rect 13920 30414 13934 30466
rect 13986 30414 14000 30466
rect 13920 30400 14000 30414
rect 14080 30466 14160 30480
rect 14080 30414 14094 30466
rect 14146 30414 14160 30466
rect 14080 30400 14160 30414
rect 14240 30466 14320 30480
rect 14240 30414 14254 30466
rect 14306 30414 14320 30466
rect 14240 30400 14320 30414
rect 14400 30466 14480 30480
rect 14400 30414 14414 30466
rect 14466 30414 14480 30466
rect 14400 30400 14480 30414
rect 14560 30466 14640 30480
rect 14560 30414 14574 30466
rect 14626 30414 14640 30466
rect 14560 30400 14640 30414
rect 14720 30466 14800 30480
rect 14720 30414 14734 30466
rect 14786 30414 14800 30466
rect 14720 30400 14800 30414
rect 14880 30466 14960 30480
rect 14880 30414 14894 30466
rect 14946 30414 14960 30466
rect 14880 30400 14960 30414
rect 15040 30466 15120 30480
rect 15040 30414 15054 30466
rect 15106 30414 15120 30466
rect 15040 30400 15120 30414
rect 15200 30466 15280 30480
rect 15200 30414 15214 30466
rect 15266 30414 15280 30466
rect 15200 30400 15280 30414
rect 15360 30466 15440 30480
rect 15360 30414 15374 30466
rect 15426 30414 15440 30466
rect 15360 30400 15440 30414
rect 15520 30466 15600 30480
rect 15520 30414 15534 30466
rect 15586 30414 15600 30466
rect 15520 30400 15600 30414
rect 15680 30466 15760 30480
rect 15680 30414 15694 30466
rect 15746 30414 15760 30466
rect 15680 30400 15760 30414
rect 15840 30466 15920 30480
rect 15840 30414 15854 30466
rect 15906 30414 15920 30466
rect 15840 30400 15920 30414
rect 16000 30466 16080 30480
rect 16000 30414 16014 30466
rect 16066 30414 16080 30466
rect 16000 30400 16080 30414
rect 16160 30466 16240 30480
rect 16160 30414 16174 30466
rect 16226 30414 16240 30466
rect 16160 30400 16240 30414
rect 16320 30466 16400 30480
rect 16320 30414 16334 30466
rect 16386 30414 16400 30466
rect 16320 30400 16400 30414
rect 16480 30466 16560 30480
rect 16480 30414 16494 30466
rect 16546 30414 16560 30466
rect 16480 30400 16560 30414
rect 16640 30466 16720 30480
rect 16640 30414 16654 30466
rect 16706 30414 16720 30466
rect 16640 30400 16720 30414
rect 16800 30466 16880 30480
rect 16800 30414 16814 30466
rect 16866 30414 16880 30466
rect 16800 30400 16880 30414
rect 16960 30466 17040 30480
rect 16960 30414 16974 30466
rect 17026 30414 17040 30466
rect 16960 30400 17040 30414
rect 17120 30466 17200 30480
rect 17120 30414 17134 30466
rect 17186 30414 17200 30466
rect 17120 30400 17200 30414
rect 17280 30466 17360 30480
rect 17280 30414 17294 30466
rect 17346 30414 17360 30466
rect 17280 30400 17360 30414
rect 17440 30466 17520 30480
rect 17440 30414 17454 30466
rect 17506 30414 17520 30466
rect 17440 30400 17520 30414
rect 17600 30466 17680 30480
rect 17600 30414 17614 30466
rect 17666 30414 17680 30466
rect 17600 30400 17680 30414
rect 17760 30466 17840 30480
rect 17760 30414 17774 30466
rect 17826 30414 17840 30466
rect 17760 30400 17840 30414
rect 17920 30466 18000 30480
rect 17920 30414 17934 30466
rect 17986 30414 18000 30466
rect 17920 30400 18000 30414
rect 18080 30466 18160 30480
rect 18080 30414 18094 30466
rect 18146 30414 18160 30466
rect 18080 30400 18160 30414
rect 18240 30466 18320 30480
rect 18240 30414 18254 30466
rect 18306 30414 18320 30466
rect 18240 30400 18320 30414
rect 18400 30466 18480 30480
rect 18400 30414 18414 30466
rect 18466 30414 18480 30466
rect 18400 30400 18480 30414
rect 18560 30466 18640 30480
rect 18560 30414 18574 30466
rect 18626 30414 18640 30466
rect 18560 30400 18640 30414
rect 18720 30466 18800 30480
rect 18720 30414 18734 30466
rect 18786 30414 18800 30466
rect 18720 30400 18800 30414
rect 18880 30466 18960 30480
rect 18880 30414 18894 30466
rect 18946 30414 18960 30466
rect 18880 30400 18960 30414
rect 23120 30466 23200 30480
rect 23120 30414 23134 30466
rect 23186 30414 23200 30466
rect 23120 30400 23200 30414
rect 23280 30466 23360 30480
rect 23280 30414 23294 30466
rect 23346 30414 23360 30466
rect 23280 30400 23360 30414
rect 23440 30466 23520 30480
rect 23440 30414 23454 30466
rect 23506 30414 23520 30466
rect 23440 30400 23520 30414
rect 23600 30466 23680 30480
rect 23600 30414 23614 30466
rect 23666 30414 23680 30466
rect 23600 30400 23680 30414
rect 23760 30466 23840 30480
rect 23760 30414 23774 30466
rect 23826 30414 23840 30466
rect 23760 30400 23840 30414
rect 23920 30466 24000 30480
rect 23920 30414 23934 30466
rect 23986 30414 24000 30466
rect 23920 30400 24000 30414
rect 24080 30466 24160 30480
rect 24080 30414 24094 30466
rect 24146 30414 24160 30466
rect 24080 30400 24160 30414
rect 24240 30466 24320 30480
rect 24240 30414 24254 30466
rect 24306 30414 24320 30466
rect 24240 30400 24320 30414
rect 24400 30466 24480 30480
rect 24400 30414 24414 30466
rect 24466 30414 24480 30466
rect 24400 30400 24480 30414
rect 24560 30466 24640 30480
rect 24560 30414 24574 30466
rect 24626 30414 24640 30466
rect 24560 30400 24640 30414
rect 24720 30466 24800 30480
rect 24720 30414 24734 30466
rect 24786 30414 24800 30466
rect 24720 30400 24800 30414
rect 24880 30466 24960 30480
rect 24880 30414 24894 30466
rect 24946 30414 24960 30466
rect 24880 30400 24960 30414
rect 25040 30466 25120 30480
rect 25040 30414 25054 30466
rect 25106 30414 25120 30466
rect 25040 30400 25120 30414
rect 25200 30466 25280 30480
rect 25200 30414 25214 30466
rect 25266 30414 25280 30466
rect 25200 30400 25280 30414
rect 25360 30466 25440 30480
rect 25360 30414 25374 30466
rect 25426 30414 25440 30466
rect 25360 30400 25440 30414
rect 25520 30466 25600 30480
rect 25520 30414 25534 30466
rect 25586 30414 25600 30466
rect 25520 30400 25600 30414
rect 25680 30466 25760 30480
rect 25680 30414 25694 30466
rect 25746 30414 25760 30466
rect 25680 30400 25760 30414
rect 25840 30466 25920 30480
rect 25840 30414 25854 30466
rect 25906 30414 25920 30466
rect 25840 30400 25920 30414
rect 26000 30466 26080 30480
rect 26000 30414 26014 30466
rect 26066 30414 26080 30466
rect 26000 30400 26080 30414
rect 26160 30466 26240 30480
rect 26160 30414 26174 30466
rect 26226 30414 26240 30466
rect 26160 30400 26240 30414
rect 26320 30466 26400 30480
rect 26320 30414 26334 30466
rect 26386 30414 26400 30466
rect 26320 30400 26400 30414
rect 26480 30466 26560 30480
rect 26480 30414 26494 30466
rect 26546 30414 26560 30466
rect 26480 30400 26560 30414
rect 26640 30466 26720 30480
rect 26640 30414 26654 30466
rect 26706 30414 26720 30466
rect 26640 30400 26720 30414
rect 26800 30466 26880 30480
rect 26800 30414 26814 30466
rect 26866 30414 26880 30466
rect 26800 30400 26880 30414
rect 26960 30466 27040 30480
rect 26960 30414 26974 30466
rect 27026 30414 27040 30466
rect 26960 30400 27040 30414
rect 27120 30466 27200 30480
rect 27120 30414 27134 30466
rect 27186 30414 27200 30466
rect 27120 30400 27200 30414
rect 27280 30466 27360 30480
rect 27280 30414 27294 30466
rect 27346 30414 27360 30466
rect 27280 30400 27360 30414
rect 27440 30466 27520 30480
rect 27440 30414 27454 30466
rect 27506 30414 27520 30466
rect 27440 30400 27520 30414
rect 27600 30466 27680 30480
rect 27600 30414 27614 30466
rect 27666 30414 27680 30466
rect 27600 30400 27680 30414
rect 27760 30466 27840 30480
rect 27760 30414 27774 30466
rect 27826 30414 27840 30466
rect 27760 30400 27840 30414
rect 27920 30466 28000 30480
rect 27920 30414 27934 30466
rect 27986 30414 28000 30466
rect 27920 30400 28000 30414
rect 28080 30466 28160 30480
rect 28080 30414 28094 30466
rect 28146 30414 28160 30466
rect 28080 30400 28160 30414
rect 28240 30466 28320 30480
rect 28240 30414 28254 30466
rect 28306 30414 28320 30466
rect 28240 30400 28320 30414
rect 28400 30466 28480 30480
rect 28400 30414 28414 30466
rect 28466 30414 28480 30466
rect 28400 30400 28480 30414
rect 28560 30466 28640 30480
rect 28560 30414 28574 30466
rect 28626 30414 28640 30466
rect 28560 30400 28640 30414
rect 28720 30466 28800 30480
rect 28720 30414 28734 30466
rect 28786 30414 28800 30466
rect 28720 30400 28800 30414
rect 28880 30466 28960 30480
rect 28880 30414 28894 30466
rect 28946 30414 28960 30466
rect 28880 30400 28960 30414
rect 29040 30466 29120 30480
rect 29040 30414 29054 30466
rect 29106 30414 29120 30466
rect 29040 30400 29120 30414
rect 29200 30466 29280 30480
rect 29200 30414 29214 30466
rect 29266 30414 29280 30466
rect 29200 30400 29280 30414
rect 29360 30466 29440 30480
rect 29360 30414 29374 30466
rect 29426 30414 29440 30466
rect 29360 30400 29440 30414
rect 33520 30466 33600 30480
rect 33520 30414 33534 30466
rect 33586 30414 33600 30466
rect 33520 30400 33600 30414
rect 33680 30466 33760 30480
rect 33680 30414 33694 30466
rect 33746 30414 33760 30466
rect 33680 30400 33760 30414
rect 33840 30466 33920 30480
rect 33840 30414 33854 30466
rect 33906 30414 33920 30466
rect 33840 30400 33920 30414
rect 34000 30466 34080 30480
rect 34000 30414 34014 30466
rect 34066 30414 34080 30466
rect 34000 30400 34080 30414
rect 34160 30466 34240 30480
rect 34160 30414 34174 30466
rect 34226 30414 34240 30466
rect 34160 30400 34240 30414
rect 34320 30466 34400 30480
rect 34320 30414 34334 30466
rect 34386 30414 34400 30466
rect 34320 30400 34400 30414
rect 34480 30466 34560 30480
rect 34480 30414 34494 30466
rect 34546 30414 34560 30466
rect 34480 30400 34560 30414
rect 34640 30466 34720 30480
rect 34640 30414 34654 30466
rect 34706 30414 34720 30466
rect 34640 30400 34720 30414
rect 34800 30466 34880 30480
rect 34800 30414 34814 30466
rect 34866 30414 34880 30466
rect 34800 30400 34880 30414
rect 34960 30466 35040 30480
rect 34960 30414 34974 30466
rect 35026 30414 35040 30466
rect 34960 30400 35040 30414
rect 35120 30466 35200 30480
rect 35120 30414 35134 30466
rect 35186 30414 35200 30466
rect 35120 30400 35200 30414
rect 35280 30466 35360 30480
rect 35280 30414 35294 30466
rect 35346 30414 35360 30466
rect 35280 30400 35360 30414
rect 35440 30466 35520 30480
rect 35440 30414 35454 30466
rect 35506 30414 35520 30466
rect 35440 30400 35520 30414
rect 35600 30466 35680 30480
rect 35600 30414 35614 30466
rect 35666 30414 35680 30466
rect 35600 30400 35680 30414
rect 35760 30466 35840 30480
rect 35760 30414 35774 30466
rect 35826 30414 35840 30466
rect 35760 30400 35840 30414
rect 35920 30466 36000 30480
rect 35920 30414 35934 30466
rect 35986 30414 36000 30466
rect 35920 30400 36000 30414
rect 36080 30466 36160 30480
rect 36080 30414 36094 30466
rect 36146 30414 36160 30466
rect 36080 30400 36160 30414
rect 36240 30466 36320 30480
rect 36240 30414 36254 30466
rect 36306 30414 36320 30466
rect 36240 30400 36320 30414
rect 36400 30466 36480 30480
rect 36400 30414 36414 30466
rect 36466 30414 36480 30466
rect 36400 30400 36480 30414
rect 36560 30466 36640 30480
rect 36560 30414 36574 30466
rect 36626 30414 36640 30466
rect 36560 30400 36640 30414
rect 36720 30466 36800 30480
rect 36720 30414 36734 30466
rect 36786 30414 36800 30466
rect 36720 30400 36800 30414
rect 36880 30466 36960 30480
rect 36880 30414 36894 30466
rect 36946 30414 36960 30466
rect 36880 30400 36960 30414
rect 37040 30466 37120 30480
rect 37040 30414 37054 30466
rect 37106 30414 37120 30466
rect 37040 30400 37120 30414
rect 37200 30466 37280 30480
rect 37200 30414 37214 30466
rect 37266 30414 37280 30466
rect 37200 30400 37280 30414
rect 37360 30466 37440 30480
rect 37360 30414 37374 30466
rect 37426 30414 37440 30466
rect 37360 30400 37440 30414
rect 37520 30466 37600 30480
rect 37520 30414 37534 30466
rect 37586 30414 37600 30466
rect 37520 30400 37600 30414
rect 37680 30466 37760 30480
rect 37680 30414 37694 30466
rect 37746 30414 37760 30466
rect 37680 30400 37760 30414
rect 37840 30466 37920 30480
rect 37840 30414 37854 30466
rect 37906 30414 37920 30466
rect 37840 30400 37920 30414
rect 38000 30466 38080 30480
rect 38000 30414 38014 30466
rect 38066 30414 38080 30466
rect 38000 30400 38080 30414
rect 38160 30466 38240 30480
rect 38160 30414 38174 30466
rect 38226 30414 38240 30466
rect 38160 30400 38240 30414
rect 38320 30466 38400 30480
rect 38320 30414 38334 30466
rect 38386 30414 38400 30466
rect 38320 30400 38400 30414
rect 38480 30466 38560 30480
rect 38480 30414 38494 30466
rect 38546 30414 38560 30466
rect 38480 30400 38560 30414
rect 38640 30466 38720 30480
rect 38640 30414 38654 30466
rect 38706 30414 38720 30466
rect 38640 30400 38720 30414
rect 38800 30466 38880 30480
rect 38800 30414 38814 30466
rect 38866 30414 38880 30466
rect 38800 30400 38880 30414
rect 38960 30466 39040 30480
rect 38960 30414 38974 30466
rect 39026 30414 39040 30466
rect 38960 30400 39040 30414
rect 39120 30466 39200 30480
rect 39120 30414 39134 30466
rect 39186 30414 39200 30466
rect 39120 30400 39200 30414
rect 39280 30466 39360 30480
rect 39280 30414 39294 30466
rect 39346 30414 39360 30466
rect 39280 30400 39360 30414
rect 39440 30466 39520 30480
rect 39440 30414 39454 30466
rect 39506 30414 39520 30466
rect 39440 30400 39520 30414
rect 39600 30466 39680 30480
rect 39600 30414 39614 30466
rect 39666 30414 39680 30466
rect 39600 30400 39680 30414
rect 39760 30466 39840 30480
rect 39760 30414 39774 30466
rect 39826 30414 39840 30466
rect 39760 30400 39840 30414
rect 39920 30466 40000 30480
rect 39920 30414 39934 30466
rect 39986 30414 40000 30466
rect 39920 30400 40000 30414
rect 40080 30466 40160 30480
rect 40080 30414 40094 30466
rect 40146 30414 40160 30466
rect 40080 30400 40160 30414
rect 40240 30466 40320 30480
rect 40240 30414 40254 30466
rect 40306 30414 40320 30466
rect 40240 30400 40320 30414
rect 40400 30466 40480 30480
rect 40400 30414 40414 30466
rect 40466 30414 40480 30466
rect 40400 30400 40480 30414
rect 40560 30466 40640 30480
rect 40560 30414 40574 30466
rect 40626 30414 40640 30466
rect 40560 30400 40640 30414
rect 40720 30466 40800 30480
rect 40720 30414 40734 30466
rect 40786 30414 40800 30466
rect 40720 30400 40800 30414
rect 40880 30466 40960 30480
rect 40880 30414 40894 30466
rect 40946 30414 40960 30466
rect 40880 30400 40960 30414
rect 41040 30466 41120 30480
rect 41040 30414 41054 30466
rect 41106 30414 41120 30466
rect 41040 30400 41120 30414
rect 41200 30466 41280 30480
rect 41200 30414 41214 30466
rect 41266 30414 41280 30466
rect 41200 30400 41280 30414
rect 41360 30466 41440 30480
rect 41360 30414 41374 30466
rect 41426 30414 41440 30466
rect 41360 30400 41440 30414
rect 41520 30466 41600 30480
rect 41520 30414 41534 30466
rect 41586 30414 41600 30466
rect 41520 30400 41600 30414
rect 41680 30466 41760 30480
rect 41680 30414 41694 30466
rect 41746 30414 41760 30466
rect 41680 30400 41760 30414
rect 41840 30466 41920 30480
rect 41840 30414 41854 30466
rect 41906 30414 41920 30466
rect 41840 30400 41920 30414
rect 0 30306 80 30320
rect 0 30254 14 30306
rect 66 30254 80 30306
rect 0 30240 80 30254
rect 160 30306 240 30320
rect 160 30254 174 30306
rect 226 30254 240 30306
rect 160 30240 240 30254
rect 320 30306 400 30320
rect 320 30254 334 30306
rect 386 30254 400 30306
rect 320 30240 400 30254
rect 480 30306 560 30320
rect 480 30254 494 30306
rect 546 30254 560 30306
rect 480 30240 560 30254
rect 640 30306 720 30320
rect 640 30254 654 30306
rect 706 30254 720 30306
rect 640 30240 720 30254
rect 800 30306 880 30320
rect 800 30254 814 30306
rect 866 30254 880 30306
rect 800 30240 880 30254
rect 960 30306 1040 30320
rect 960 30254 974 30306
rect 1026 30254 1040 30306
rect 960 30240 1040 30254
rect 1120 30306 1200 30320
rect 1120 30254 1134 30306
rect 1186 30254 1200 30306
rect 1120 30240 1200 30254
rect 1280 30306 1360 30320
rect 1280 30254 1294 30306
rect 1346 30254 1360 30306
rect 1280 30240 1360 30254
rect 1440 30306 1520 30320
rect 1440 30254 1454 30306
rect 1506 30254 1520 30306
rect 1440 30240 1520 30254
rect 1600 30306 1680 30320
rect 1600 30254 1614 30306
rect 1666 30254 1680 30306
rect 1600 30240 1680 30254
rect 1760 30306 1840 30320
rect 1760 30254 1774 30306
rect 1826 30254 1840 30306
rect 1760 30240 1840 30254
rect 1920 30306 2000 30320
rect 1920 30254 1934 30306
rect 1986 30254 2000 30306
rect 1920 30240 2000 30254
rect 2080 30306 2160 30320
rect 2080 30254 2094 30306
rect 2146 30254 2160 30306
rect 2080 30240 2160 30254
rect 2240 30306 2320 30320
rect 2240 30254 2254 30306
rect 2306 30254 2320 30306
rect 2240 30240 2320 30254
rect 2400 30306 2480 30320
rect 2400 30254 2414 30306
rect 2466 30254 2480 30306
rect 2400 30240 2480 30254
rect 2560 30306 2640 30320
rect 2560 30254 2574 30306
rect 2626 30254 2640 30306
rect 2560 30240 2640 30254
rect 2720 30306 2800 30320
rect 2720 30254 2734 30306
rect 2786 30254 2800 30306
rect 2720 30240 2800 30254
rect 2880 30306 2960 30320
rect 2880 30254 2894 30306
rect 2946 30254 2960 30306
rect 2880 30240 2960 30254
rect 3040 30306 3120 30320
rect 3040 30254 3054 30306
rect 3106 30254 3120 30306
rect 3040 30240 3120 30254
rect 3200 30306 3280 30320
rect 3200 30254 3214 30306
rect 3266 30254 3280 30306
rect 3200 30240 3280 30254
rect 3360 30306 3440 30320
rect 3360 30254 3374 30306
rect 3426 30254 3440 30306
rect 3360 30240 3440 30254
rect 3520 30306 3600 30320
rect 3520 30254 3534 30306
rect 3586 30254 3600 30306
rect 3520 30240 3600 30254
rect 3680 30306 3760 30320
rect 3680 30254 3694 30306
rect 3746 30254 3760 30306
rect 3680 30240 3760 30254
rect 3840 30306 3920 30320
rect 3840 30254 3854 30306
rect 3906 30254 3920 30306
rect 3840 30240 3920 30254
rect 4000 30306 4080 30320
rect 4000 30254 4014 30306
rect 4066 30254 4080 30306
rect 4000 30240 4080 30254
rect 4160 30306 4240 30320
rect 4160 30254 4174 30306
rect 4226 30254 4240 30306
rect 4160 30240 4240 30254
rect 4320 30306 4400 30320
rect 4320 30254 4334 30306
rect 4386 30254 4400 30306
rect 4320 30240 4400 30254
rect 4480 30306 4560 30320
rect 4480 30254 4494 30306
rect 4546 30254 4560 30306
rect 4480 30240 4560 30254
rect 4640 30306 4720 30320
rect 4640 30254 4654 30306
rect 4706 30254 4720 30306
rect 4640 30240 4720 30254
rect 4800 30306 4880 30320
rect 4800 30254 4814 30306
rect 4866 30254 4880 30306
rect 4800 30240 4880 30254
rect 4960 30306 5040 30320
rect 4960 30254 4974 30306
rect 5026 30254 5040 30306
rect 4960 30240 5040 30254
rect 5120 30306 5200 30320
rect 5120 30254 5134 30306
rect 5186 30254 5200 30306
rect 5120 30240 5200 30254
rect 5280 30306 5360 30320
rect 5280 30254 5294 30306
rect 5346 30254 5360 30306
rect 5280 30240 5360 30254
rect 5440 30306 5520 30320
rect 5440 30254 5454 30306
rect 5506 30254 5520 30306
rect 5440 30240 5520 30254
rect 5600 30306 5680 30320
rect 5600 30254 5614 30306
rect 5666 30254 5680 30306
rect 5600 30240 5680 30254
rect 5760 30306 5840 30320
rect 5760 30254 5774 30306
rect 5826 30254 5840 30306
rect 5760 30240 5840 30254
rect 5920 30306 6000 30320
rect 5920 30254 5934 30306
rect 5986 30254 6000 30306
rect 5920 30240 6000 30254
rect 6080 30306 6160 30320
rect 6080 30254 6094 30306
rect 6146 30254 6160 30306
rect 6080 30240 6160 30254
rect 6240 30306 6320 30320
rect 6240 30254 6254 30306
rect 6306 30254 6320 30306
rect 6240 30240 6320 30254
rect 6400 30306 6480 30320
rect 6400 30254 6414 30306
rect 6466 30254 6480 30306
rect 6400 30240 6480 30254
rect 6560 30306 6640 30320
rect 6560 30254 6574 30306
rect 6626 30254 6640 30306
rect 6560 30240 6640 30254
rect 6720 30306 6800 30320
rect 6720 30254 6734 30306
rect 6786 30254 6800 30306
rect 6720 30240 6800 30254
rect 6880 30306 6960 30320
rect 6880 30254 6894 30306
rect 6946 30254 6960 30306
rect 6880 30240 6960 30254
rect 7040 30306 7120 30320
rect 7040 30254 7054 30306
rect 7106 30254 7120 30306
rect 7040 30240 7120 30254
rect 7200 30306 7280 30320
rect 7200 30254 7214 30306
rect 7266 30254 7280 30306
rect 7200 30240 7280 30254
rect 7360 30306 7440 30320
rect 7360 30254 7374 30306
rect 7426 30254 7440 30306
rect 7360 30240 7440 30254
rect 7520 30306 7600 30320
rect 7520 30254 7534 30306
rect 7586 30254 7600 30306
rect 7520 30240 7600 30254
rect 7680 30306 7760 30320
rect 7680 30254 7694 30306
rect 7746 30254 7760 30306
rect 7680 30240 7760 30254
rect 7840 30306 7920 30320
rect 7840 30254 7854 30306
rect 7906 30254 7920 30306
rect 7840 30240 7920 30254
rect 8000 30306 8080 30320
rect 8000 30254 8014 30306
rect 8066 30254 8080 30306
rect 8000 30240 8080 30254
rect 8160 30306 8240 30320
rect 8160 30254 8174 30306
rect 8226 30254 8240 30306
rect 8160 30240 8240 30254
rect 8320 30306 8400 30320
rect 8320 30254 8334 30306
rect 8386 30254 8400 30306
rect 8320 30240 8400 30254
rect 12480 30306 12560 30320
rect 12480 30254 12494 30306
rect 12546 30254 12560 30306
rect 12480 30240 12560 30254
rect 12640 30306 12720 30320
rect 12640 30254 12654 30306
rect 12706 30254 12720 30306
rect 12640 30240 12720 30254
rect 12800 30306 12880 30320
rect 12800 30254 12814 30306
rect 12866 30254 12880 30306
rect 12800 30240 12880 30254
rect 12960 30306 13040 30320
rect 12960 30254 12974 30306
rect 13026 30254 13040 30306
rect 12960 30240 13040 30254
rect 13120 30306 13200 30320
rect 13120 30254 13134 30306
rect 13186 30254 13200 30306
rect 13120 30240 13200 30254
rect 13280 30306 13360 30320
rect 13280 30254 13294 30306
rect 13346 30254 13360 30306
rect 13280 30240 13360 30254
rect 13440 30306 13520 30320
rect 13440 30254 13454 30306
rect 13506 30254 13520 30306
rect 13440 30240 13520 30254
rect 13600 30306 13680 30320
rect 13600 30254 13614 30306
rect 13666 30254 13680 30306
rect 13600 30240 13680 30254
rect 13760 30306 13840 30320
rect 13760 30254 13774 30306
rect 13826 30254 13840 30306
rect 13760 30240 13840 30254
rect 13920 30306 14000 30320
rect 13920 30254 13934 30306
rect 13986 30254 14000 30306
rect 13920 30240 14000 30254
rect 14080 30306 14160 30320
rect 14080 30254 14094 30306
rect 14146 30254 14160 30306
rect 14080 30240 14160 30254
rect 14240 30306 14320 30320
rect 14240 30254 14254 30306
rect 14306 30254 14320 30306
rect 14240 30240 14320 30254
rect 14400 30306 14480 30320
rect 14400 30254 14414 30306
rect 14466 30254 14480 30306
rect 14400 30240 14480 30254
rect 14560 30306 14640 30320
rect 14560 30254 14574 30306
rect 14626 30254 14640 30306
rect 14560 30240 14640 30254
rect 14720 30306 14800 30320
rect 14720 30254 14734 30306
rect 14786 30254 14800 30306
rect 14720 30240 14800 30254
rect 14880 30306 14960 30320
rect 14880 30254 14894 30306
rect 14946 30254 14960 30306
rect 14880 30240 14960 30254
rect 15040 30306 15120 30320
rect 15040 30254 15054 30306
rect 15106 30254 15120 30306
rect 15040 30240 15120 30254
rect 15200 30306 15280 30320
rect 15200 30254 15214 30306
rect 15266 30254 15280 30306
rect 15200 30240 15280 30254
rect 15360 30306 15440 30320
rect 15360 30254 15374 30306
rect 15426 30254 15440 30306
rect 15360 30240 15440 30254
rect 15520 30306 15600 30320
rect 15520 30254 15534 30306
rect 15586 30254 15600 30306
rect 15520 30240 15600 30254
rect 15680 30306 15760 30320
rect 15680 30254 15694 30306
rect 15746 30254 15760 30306
rect 15680 30240 15760 30254
rect 15840 30306 15920 30320
rect 15840 30254 15854 30306
rect 15906 30254 15920 30306
rect 15840 30240 15920 30254
rect 16000 30306 16080 30320
rect 16000 30254 16014 30306
rect 16066 30254 16080 30306
rect 16000 30240 16080 30254
rect 16160 30306 16240 30320
rect 16160 30254 16174 30306
rect 16226 30254 16240 30306
rect 16160 30240 16240 30254
rect 16320 30306 16400 30320
rect 16320 30254 16334 30306
rect 16386 30254 16400 30306
rect 16320 30240 16400 30254
rect 16480 30306 16560 30320
rect 16480 30254 16494 30306
rect 16546 30254 16560 30306
rect 16480 30240 16560 30254
rect 16640 30306 16720 30320
rect 16640 30254 16654 30306
rect 16706 30254 16720 30306
rect 16640 30240 16720 30254
rect 16800 30306 16880 30320
rect 16800 30254 16814 30306
rect 16866 30254 16880 30306
rect 16800 30240 16880 30254
rect 16960 30306 17040 30320
rect 16960 30254 16974 30306
rect 17026 30254 17040 30306
rect 16960 30240 17040 30254
rect 17120 30306 17200 30320
rect 17120 30254 17134 30306
rect 17186 30254 17200 30306
rect 17120 30240 17200 30254
rect 17280 30306 17360 30320
rect 17280 30254 17294 30306
rect 17346 30254 17360 30306
rect 17280 30240 17360 30254
rect 17440 30306 17520 30320
rect 17440 30254 17454 30306
rect 17506 30254 17520 30306
rect 17440 30240 17520 30254
rect 17600 30306 17680 30320
rect 17600 30254 17614 30306
rect 17666 30254 17680 30306
rect 17600 30240 17680 30254
rect 17760 30306 17840 30320
rect 17760 30254 17774 30306
rect 17826 30254 17840 30306
rect 17760 30240 17840 30254
rect 17920 30306 18000 30320
rect 17920 30254 17934 30306
rect 17986 30254 18000 30306
rect 17920 30240 18000 30254
rect 18080 30306 18160 30320
rect 18080 30254 18094 30306
rect 18146 30254 18160 30306
rect 18080 30240 18160 30254
rect 18240 30306 18320 30320
rect 18240 30254 18254 30306
rect 18306 30254 18320 30306
rect 18240 30240 18320 30254
rect 18400 30306 18480 30320
rect 18400 30254 18414 30306
rect 18466 30254 18480 30306
rect 18400 30240 18480 30254
rect 18560 30306 18640 30320
rect 18560 30254 18574 30306
rect 18626 30254 18640 30306
rect 18560 30240 18640 30254
rect 18720 30306 18800 30320
rect 18720 30254 18734 30306
rect 18786 30254 18800 30306
rect 18720 30240 18800 30254
rect 18880 30306 18960 30320
rect 18880 30254 18894 30306
rect 18946 30254 18960 30306
rect 18880 30240 18960 30254
rect 23120 30306 23200 30320
rect 23120 30254 23134 30306
rect 23186 30254 23200 30306
rect 23120 30240 23200 30254
rect 23280 30306 23360 30320
rect 23280 30254 23294 30306
rect 23346 30254 23360 30306
rect 23280 30240 23360 30254
rect 23440 30306 23520 30320
rect 23440 30254 23454 30306
rect 23506 30254 23520 30306
rect 23440 30240 23520 30254
rect 23600 30306 23680 30320
rect 23600 30254 23614 30306
rect 23666 30254 23680 30306
rect 23600 30240 23680 30254
rect 23760 30306 23840 30320
rect 23760 30254 23774 30306
rect 23826 30254 23840 30306
rect 23760 30240 23840 30254
rect 23920 30306 24000 30320
rect 23920 30254 23934 30306
rect 23986 30254 24000 30306
rect 23920 30240 24000 30254
rect 24080 30306 24160 30320
rect 24080 30254 24094 30306
rect 24146 30254 24160 30306
rect 24080 30240 24160 30254
rect 24240 30306 24320 30320
rect 24240 30254 24254 30306
rect 24306 30254 24320 30306
rect 24240 30240 24320 30254
rect 24400 30306 24480 30320
rect 24400 30254 24414 30306
rect 24466 30254 24480 30306
rect 24400 30240 24480 30254
rect 24560 30306 24640 30320
rect 24560 30254 24574 30306
rect 24626 30254 24640 30306
rect 24560 30240 24640 30254
rect 24720 30306 24800 30320
rect 24720 30254 24734 30306
rect 24786 30254 24800 30306
rect 24720 30240 24800 30254
rect 24880 30306 24960 30320
rect 24880 30254 24894 30306
rect 24946 30254 24960 30306
rect 24880 30240 24960 30254
rect 25040 30306 25120 30320
rect 25040 30254 25054 30306
rect 25106 30254 25120 30306
rect 25040 30240 25120 30254
rect 25200 30306 25280 30320
rect 25200 30254 25214 30306
rect 25266 30254 25280 30306
rect 25200 30240 25280 30254
rect 25360 30306 25440 30320
rect 25360 30254 25374 30306
rect 25426 30254 25440 30306
rect 25360 30240 25440 30254
rect 25520 30306 25600 30320
rect 25520 30254 25534 30306
rect 25586 30254 25600 30306
rect 25520 30240 25600 30254
rect 25680 30306 25760 30320
rect 25680 30254 25694 30306
rect 25746 30254 25760 30306
rect 25680 30240 25760 30254
rect 25840 30306 25920 30320
rect 25840 30254 25854 30306
rect 25906 30254 25920 30306
rect 25840 30240 25920 30254
rect 26000 30306 26080 30320
rect 26000 30254 26014 30306
rect 26066 30254 26080 30306
rect 26000 30240 26080 30254
rect 26160 30306 26240 30320
rect 26160 30254 26174 30306
rect 26226 30254 26240 30306
rect 26160 30240 26240 30254
rect 26320 30306 26400 30320
rect 26320 30254 26334 30306
rect 26386 30254 26400 30306
rect 26320 30240 26400 30254
rect 26480 30306 26560 30320
rect 26480 30254 26494 30306
rect 26546 30254 26560 30306
rect 26480 30240 26560 30254
rect 26640 30306 26720 30320
rect 26640 30254 26654 30306
rect 26706 30254 26720 30306
rect 26640 30240 26720 30254
rect 26800 30306 26880 30320
rect 26800 30254 26814 30306
rect 26866 30254 26880 30306
rect 26800 30240 26880 30254
rect 26960 30306 27040 30320
rect 26960 30254 26974 30306
rect 27026 30254 27040 30306
rect 26960 30240 27040 30254
rect 27120 30306 27200 30320
rect 27120 30254 27134 30306
rect 27186 30254 27200 30306
rect 27120 30240 27200 30254
rect 27280 30306 27360 30320
rect 27280 30254 27294 30306
rect 27346 30254 27360 30306
rect 27280 30240 27360 30254
rect 27440 30306 27520 30320
rect 27440 30254 27454 30306
rect 27506 30254 27520 30306
rect 27440 30240 27520 30254
rect 27600 30306 27680 30320
rect 27600 30254 27614 30306
rect 27666 30254 27680 30306
rect 27600 30240 27680 30254
rect 27760 30306 27840 30320
rect 27760 30254 27774 30306
rect 27826 30254 27840 30306
rect 27760 30240 27840 30254
rect 27920 30306 28000 30320
rect 27920 30254 27934 30306
rect 27986 30254 28000 30306
rect 27920 30240 28000 30254
rect 28080 30306 28160 30320
rect 28080 30254 28094 30306
rect 28146 30254 28160 30306
rect 28080 30240 28160 30254
rect 28240 30306 28320 30320
rect 28240 30254 28254 30306
rect 28306 30254 28320 30306
rect 28240 30240 28320 30254
rect 28400 30306 28480 30320
rect 28400 30254 28414 30306
rect 28466 30254 28480 30306
rect 28400 30240 28480 30254
rect 28560 30306 28640 30320
rect 28560 30254 28574 30306
rect 28626 30254 28640 30306
rect 28560 30240 28640 30254
rect 28720 30306 28800 30320
rect 28720 30254 28734 30306
rect 28786 30254 28800 30306
rect 28720 30240 28800 30254
rect 28880 30306 28960 30320
rect 28880 30254 28894 30306
rect 28946 30254 28960 30306
rect 28880 30240 28960 30254
rect 29040 30306 29120 30320
rect 29040 30254 29054 30306
rect 29106 30254 29120 30306
rect 29040 30240 29120 30254
rect 29200 30306 29280 30320
rect 29200 30254 29214 30306
rect 29266 30254 29280 30306
rect 29200 30240 29280 30254
rect 29360 30306 29440 30320
rect 29360 30254 29374 30306
rect 29426 30254 29440 30306
rect 29360 30240 29440 30254
rect 33520 30306 33600 30320
rect 33520 30254 33534 30306
rect 33586 30254 33600 30306
rect 33520 30240 33600 30254
rect 33680 30306 33760 30320
rect 33680 30254 33694 30306
rect 33746 30254 33760 30306
rect 33680 30240 33760 30254
rect 33840 30306 33920 30320
rect 33840 30254 33854 30306
rect 33906 30254 33920 30306
rect 33840 30240 33920 30254
rect 34000 30306 34080 30320
rect 34000 30254 34014 30306
rect 34066 30254 34080 30306
rect 34000 30240 34080 30254
rect 34160 30306 34240 30320
rect 34160 30254 34174 30306
rect 34226 30254 34240 30306
rect 34160 30240 34240 30254
rect 34320 30306 34400 30320
rect 34320 30254 34334 30306
rect 34386 30254 34400 30306
rect 34320 30240 34400 30254
rect 34480 30306 34560 30320
rect 34480 30254 34494 30306
rect 34546 30254 34560 30306
rect 34480 30240 34560 30254
rect 34640 30306 34720 30320
rect 34640 30254 34654 30306
rect 34706 30254 34720 30306
rect 34640 30240 34720 30254
rect 34800 30306 34880 30320
rect 34800 30254 34814 30306
rect 34866 30254 34880 30306
rect 34800 30240 34880 30254
rect 34960 30306 35040 30320
rect 34960 30254 34974 30306
rect 35026 30254 35040 30306
rect 34960 30240 35040 30254
rect 35120 30306 35200 30320
rect 35120 30254 35134 30306
rect 35186 30254 35200 30306
rect 35120 30240 35200 30254
rect 35280 30306 35360 30320
rect 35280 30254 35294 30306
rect 35346 30254 35360 30306
rect 35280 30240 35360 30254
rect 35440 30306 35520 30320
rect 35440 30254 35454 30306
rect 35506 30254 35520 30306
rect 35440 30240 35520 30254
rect 35600 30306 35680 30320
rect 35600 30254 35614 30306
rect 35666 30254 35680 30306
rect 35600 30240 35680 30254
rect 35760 30306 35840 30320
rect 35760 30254 35774 30306
rect 35826 30254 35840 30306
rect 35760 30240 35840 30254
rect 35920 30306 36000 30320
rect 35920 30254 35934 30306
rect 35986 30254 36000 30306
rect 35920 30240 36000 30254
rect 36080 30306 36160 30320
rect 36080 30254 36094 30306
rect 36146 30254 36160 30306
rect 36080 30240 36160 30254
rect 36240 30306 36320 30320
rect 36240 30254 36254 30306
rect 36306 30254 36320 30306
rect 36240 30240 36320 30254
rect 36400 30306 36480 30320
rect 36400 30254 36414 30306
rect 36466 30254 36480 30306
rect 36400 30240 36480 30254
rect 36560 30306 36640 30320
rect 36560 30254 36574 30306
rect 36626 30254 36640 30306
rect 36560 30240 36640 30254
rect 36720 30306 36800 30320
rect 36720 30254 36734 30306
rect 36786 30254 36800 30306
rect 36720 30240 36800 30254
rect 36880 30306 36960 30320
rect 36880 30254 36894 30306
rect 36946 30254 36960 30306
rect 36880 30240 36960 30254
rect 37040 30306 37120 30320
rect 37040 30254 37054 30306
rect 37106 30254 37120 30306
rect 37040 30240 37120 30254
rect 37200 30306 37280 30320
rect 37200 30254 37214 30306
rect 37266 30254 37280 30306
rect 37200 30240 37280 30254
rect 37360 30306 37440 30320
rect 37360 30254 37374 30306
rect 37426 30254 37440 30306
rect 37360 30240 37440 30254
rect 37520 30306 37600 30320
rect 37520 30254 37534 30306
rect 37586 30254 37600 30306
rect 37520 30240 37600 30254
rect 37680 30306 37760 30320
rect 37680 30254 37694 30306
rect 37746 30254 37760 30306
rect 37680 30240 37760 30254
rect 37840 30306 37920 30320
rect 37840 30254 37854 30306
rect 37906 30254 37920 30306
rect 37840 30240 37920 30254
rect 38000 30306 38080 30320
rect 38000 30254 38014 30306
rect 38066 30254 38080 30306
rect 38000 30240 38080 30254
rect 38160 30306 38240 30320
rect 38160 30254 38174 30306
rect 38226 30254 38240 30306
rect 38160 30240 38240 30254
rect 38320 30306 38400 30320
rect 38320 30254 38334 30306
rect 38386 30254 38400 30306
rect 38320 30240 38400 30254
rect 38480 30306 38560 30320
rect 38480 30254 38494 30306
rect 38546 30254 38560 30306
rect 38480 30240 38560 30254
rect 38640 30306 38720 30320
rect 38640 30254 38654 30306
rect 38706 30254 38720 30306
rect 38640 30240 38720 30254
rect 38800 30306 38880 30320
rect 38800 30254 38814 30306
rect 38866 30254 38880 30306
rect 38800 30240 38880 30254
rect 38960 30306 39040 30320
rect 38960 30254 38974 30306
rect 39026 30254 39040 30306
rect 38960 30240 39040 30254
rect 39120 30306 39200 30320
rect 39120 30254 39134 30306
rect 39186 30254 39200 30306
rect 39120 30240 39200 30254
rect 39280 30306 39360 30320
rect 39280 30254 39294 30306
rect 39346 30254 39360 30306
rect 39280 30240 39360 30254
rect 39440 30306 39520 30320
rect 39440 30254 39454 30306
rect 39506 30254 39520 30306
rect 39440 30240 39520 30254
rect 39600 30306 39680 30320
rect 39600 30254 39614 30306
rect 39666 30254 39680 30306
rect 39600 30240 39680 30254
rect 39760 30306 39840 30320
rect 39760 30254 39774 30306
rect 39826 30254 39840 30306
rect 39760 30240 39840 30254
rect 39920 30306 40000 30320
rect 39920 30254 39934 30306
rect 39986 30254 40000 30306
rect 39920 30240 40000 30254
rect 40080 30306 40160 30320
rect 40080 30254 40094 30306
rect 40146 30254 40160 30306
rect 40080 30240 40160 30254
rect 40240 30306 40320 30320
rect 40240 30254 40254 30306
rect 40306 30254 40320 30306
rect 40240 30240 40320 30254
rect 40400 30306 40480 30320
rect 40400 30254 40414 30306
rect 40466 30254 40480 30306
rect 40400 30240 40480 30254
rect 40560 30306 40640 30320
rect 40560 30254 40574 30306
rect 40626 30254 40640 30306
rect 40560 30240 40640 30254
rect 40720 30306 40800 30320
rect 40720 30254 40734 30306
rect 40786 30254 40800 30306
rect 40720 30240 40800 30254
rect 40880 30306 40960 30320
rect 40880 30254 40894 30306
rect 40946 30254 40960 30306
rect 40880 30240 40960 30254
rect 41040 30306 41120 30320
rect 41040 30254 41054 30306
rect 41106 30254 41120 30306
rect 41040 30240 41120 30254
rect 41200 30306 41280 30320
rect 41200 30254 41214 30306
rect 41266 30254 41280 30306
rect 41200 30240 41280 30254
rect 41360 30306 41440 30320
rect 41360 30254 41374 30306
rect 41426 30254 41440 30306
rect 41360 30240 41440 30254
rect 41520 30306 41600 30320
rect 41520 30254 41534 30306
rect 41586 30254 41600 30306
rect 41520 30240 41600 30254
rect 41680 30306 41760 30320
rect 41680 30254 41694 30306
rect 41746 30254 41760 30306
rect 41680 30240 41760 30254
rect 41840 30306 41920 30320
rect 41840 30254 41854 30306
rect 41906 30254 41920 30306
rect 41840 30240 41920 30254
rect 0 29986 80 30000
rect 0 29934 14 29986
rect 66 29934 80 29986
rect 0 29920 80 29934
rect 160 29986 240 30000
rect 160 29934 174 29986
rect 226 29934 240 29986
rect 160 29920 240 29934
rect 320 29986 400 30000
rect 320 29934 334 29986
rect 386 29934 400 29986
rect 320 29920 400 29934
rect 480 29986 560 30000
rect 480 29934 494 29986
rect 546 29934 560 29986
rect 480 29920 560 29934
rect 640 29986 720 30000
rect 640 29934 654 29986
rect 706 29934 720 29986
rect 640 29920 720 29934
rect 800 29986 880 30000
rect 800 29934 814 29986
rect 866 29934 880 29986
rect 800 29920 880 29934
rect 960 29986 1040 30000
rect 960 29934 974 29986
rect 1026 29934 1040 29986
rect 960 29920 1040 29934
rect 1120 29986 1200 30000
rect 1120 29934 1134 29986
rect 1186 29934 1200 29986
rect 1120 29920 1200 29934
rect 1280 29986 1360 30000
rect 1280 29934 1294 29986
rect 1346 29934 1360 29986
rect 1280 29920 1360 29934
rect 1440 29986 1520 30000
rect 1440 29934 1454 29986
rect 1506 29934 1520 29986
rect 1440 29920 1520 29934
rect 1600 29986 1680 30000
rect 1600 29934 1614 29986
rect 1666 29934 1680 29986
rect 1600 29920 1680 29934
rect 1760 29986 1840 30000
rect 1760 29934 1774 29986
rect 1826 29934 1840 29986
rect 1760 29920 1840 29934
rect 1920 29986 2000 30000
rect 1920 29934 1934 29986
rect 1986 29934 2000 29986
rect 1920 29920 2000 29934
rect 2080 29986 2160 30000
rect 2080 29934 2094 29986
rect 2146 29934 2160 29986
rect 2080 29920 2160 29934
rect 2240 29986 2320 30000
rect 2240 29934 2254 29986
rect 2306 29934 2320 29986
rect 2240 29920 2320 29934
rect 2400 29986 2480 30000
rect 2400 29934 2414 29986
rect 2466 29934 2480 29986
rect 2400 29920 2480 29934
rect 2560 29986 2640 30000
rect 2560 29934 2574 29986
rect 2626 29934 2640 29986
rect 2560 29920 2640 29934
rect 2720 29986 2800 30000
rect 2720 29934 2734 29986
rect 2786 29934 2800 29986
rect 2720 29920 2800 29934
rect 2880 29986 2960 30000
rect 2880 29934 2894 29986
rect 2946 29934 2960 29986
rect 2880 29920 2960 29934
rect 3040 29986 3120 30000
rect 3040 29934 3054 29986
rect 3106 29934 3120 29986
rect 3040 29920 3120 29934
rect 3200 29986 3280 30000
rect 3200 29934 3214 29986
rect 3266 29934 3280 29986
rect 3200 29920 3280 29934
rect 3360 29986 3440 30000
rect 3360 29934 3374 29986
rect 3426 29934 3440 29986
rect 3360 29920 3440 29934
rect 3520 29986 3600 30000
rect 3520 29934 3534 29986
rect 3586 29934 3600 29986
rect 3520 29920 3600 29934
rect 3680 29986 3760 30000
rect 3680 29934 3694 29986
rect 3746 29934 3760 29986
rect 3680 29920 3760 29934
rect 3840 29986 3920 30000
rect 3840 29934 3854 29986
rect 3906 29934 3920 29986
rect 3840 29920 3920 29934
rect 4000 29986 4080 30000
rect 4000 29934 4014 29986
rect 4066 29934 4080 29986
rect 4000 29920 4080 29934
rect 4160 29986 4240 30000
rect 4160 29934 4174 29986
rect 4226 29934 4240 29986
rect 4160 29920 4240 29934
rect 4320 29986 4400 30000
rect 4320 29934 4334 29986
rect 4386 29934 4400 29986
rect 4320 29920 4400 29934
rect 4480 29986 4560 30000
rect 4480 29934 4494 29986
rect 4546 29934 4560 29986
rect 4480 29920 4560 29934
rect 4640 29986 4720 30000
rect 4640 29934 4654 29986
rect 4706 29934 4720 29986
rect 4640 29920 4720 29934
rect 4800 29986 4880 30000
rect 4800 29934 4814 29986
rect 4866 29934 4880 29986
rect 4800 29920 4880 29934
rect 4960 29986 5040 30000
rect 4960 29934 4974 29986
rect 5026 29934 5040 29986
rect 4960 29920 5040 29934
rect 5120 29986 5200 30000
rect 5120 29934 5134 29986
rect 5186 29934 5200 29986
rect 5120 29920 5200 29934
rect 5280 29986 5360 30000
rect 5280 29934 5294 29986
rect 5346 29934 5360 29986
rect 5280 29920 5360 29934
rect 5440 29986 5520 30000
rect 5440 29934 5454 29986
rect 5506 29934 5520 29986
rect 5440 29920 5520 29934
rect 5600 29986 5680 30000
rect 5600 29934 5614 29986
rect 5666 29934 5680 29986
rect 5600 29920 5680 29934
rect 5760 29986 5840 30000
rect 5760 29934 5774 29986
rect 5826 29934 5840 29986
rect 5760 29920 5840 29934
rect 5920 29986 6000 30000
rect 5920 29934 5934 29986
rect 5986 29934 6000 29986
rect 5920 29920 6000 29934
rect 6080 29986 6160 30000
rect 6080 29934 6094 29986
rect 6146 29934 6160 29986
rect 6080 29920 6160 29934
rect 6240 29986 6320 30000
rect 6240 29934 6254 29986
rect 6306 29934 6320 29986
rect 6240 29920 6320 29934
rect 6400 29986 6480 30000
rect 6400 29934 6414 29986
rect 6466 29934 6480 29986
rect 6400 29920 6480 29934
rect 6560 29986 6640 30000
rect 6560 29934 6574 29986
rect 6626 29934 6640 29986
rect 6560 29920 6640 29934
rect 6720 29986 6800 30000
rect 6720 29934 6734 29986
rect 6786 29934 6800 29986
rect 6720 29920 6800 29934
rect 6880 29986 6960 30000
rect 6880 29934 6894 29986
rect 6946 29934 6960 29986
rect 6880 29920 6960 29934
rect 7040 29986 7120 30000
rect 7040 29934 7054 29986
rect 7106 29934 7120 29986
rect 7040 29920 7120 29934
rect 7200 29986 7280 30000
rect 7200 29934 7214 29986
rect 7266 29934 7280 29986
rect 7200 29920 7280 29934
rect 7360 29986 7440 30000
rect 7360 29934 7374 29986
rect 7426 29934 7440 29986
rect 7360 29920 7440 29934
rect 7520 29986 7600 30000
rect 7520 29934 7534 29986
rect 7586 29934 7600 29986
rect 7520 29920 7600 29934
rect 7680 29986 7760 30000
rect 7680 29934 7694 29986
rect 7746 29934 7760 29986
rect 7680 29920 7760 29934
rect 7840 29986 7920 30000
rect 7840 29934 7854 29986
rect 7906 29934 7920 29986
rect 7840 29920 7920 29934
rect 8000 29986 8080 30000
rect 8000 29934 8014 29986
rect 8066 29934 8080 29986
rect 8000 29920 8080 29934
rect 8160 29986 8240 30000
rect 8160 29934 8174 29986
rect 8226 29934 8240 29986
rect 8160 29920 8240 29934
rect 8320 29986 8400 30000
rect 8320 29934 8334 29986
rect 8386 29934 8400 29986
rect 8320 29920 8400 29934
rect 12480 29986 12560 30000
rect 12480 29934 12494 29986
rect 12546 29934 12560 29986
rect 12480 29920 12560 29934
rect 12640 29986 12720 30000
rect 12640 29934 12654 29986
rect 12706 29934 12720 29986
rect 12640 29920 12720 29934
rect 12800 29986 12880 30000
rect 12800 29934 12814 29986
rect 12866 29934 12880 29986
rect 12800 29920 12880 29934
rect 12960 29986 13040 30000
rect 12960 29934 12974 29986
rect 13026 29934 13040 29986
rect 12960 29920 13040 29934
rect 13120 29986 13200 30000
rect 13120 29934 13134 29986
rect 13186 29934 13200 29986
rect 13120 29920 13200 29934
rect 13280 29986 13360 30000
rect 13280 29934 13294 29986
rect 13346 29934 13360 29986
rect 13280 29920 13360 29934
rect 13440 29986 13520 30000
rect 13440 29934 13454 29986
rect 13506 29934 13520 29986
rect 13440 29920 13520 29934
rect 13600 29986 13680 30000
rect 13600 29934 13614 29986
rect 13666 29934 13680 29986
rect 13600 29920 13680 29934
rect 13760 29986 13840 30000
rect 13760 29934 13774 29986
rect 13826 29934 13840 29986
rect 13760 29920 13840 29934
rect 13920 29986 14000 30000
rect 13920 29934 13934 29986
rect 13986 29934 14000 29986
rect 13920 29920 14000 29934
rect 14080 29986 14160 30000
rect 14080 29934 14094 29986
rect 14146 29934 14160 29986
rect 14080 29920 14160 29934
rect 14240 29986 14320 30000
rect 14240 29934 14254 29986
rect 14306 29934 14320 29986
rect 14240 29920 14320 29934
rect 14400 29986 14480 30000
rect 14400 29934 14414 29986
rect 14466 29934 14480 29986
rect 14400 29920 14480 29934
rect 14560 29986 14640 30000
rect 14560 29934 14574 29986
rect 14626 29934 14640 29986
rect 14560 29920 14640 29934
rect 14720 29986 14800 30000
rect 14720 29934 14734 29986
rect 14786 29934 14800 29986
rect 14720 29920 14800 29934
rect 14880 29986 14960 30000
rect 14880 29934 14894 29986
rect 14946 29934 14960 29986
rect 14880 29920 14960 29934
rect 15040 29986 15120 30000
rect 15040 29934 15054 29986
rect 15106 29934 15120 29986
rect 15040 29920 15120 29934
rect 15200 29986 15280 30000
rect 15200 29934 15214 29986
rect 15266 29934 15280 29986
rect 15200 29920 15280 29934
rect 15360 29986 15440 30000
rect 15360 29934 15374 29986
rect 15426 29934 15440 29986
rect 15360 29920 15440 29934
rect 15520 29986 15600 30000
rect 15520 29934 15534 29986
rect 15586 29934 15600 29986
rect 15520 29920 15600 29934
rect 15680 29986 15760 30000
rect 15680 29934 15694 29986
rect 15746 29934 15760 29986
rect 15680 29920 15760 29934
rect 15840 29986 15920 30000
rect 15840 29934 15854 29986
rect 15906 29934 15920 29986
rect 15840 29920 15920 29934
rect 16000 29986 16080 30000
rect 16000 29934 16014 29986
rect 16066 29934 16080 29986
rect 16000 29920 16080 29934
rect 16160 29986 16240 30000
rect 16160 29934 16174 29986
rect 16226 29934 16240 29986
rect 16160 29920 16240 29934
rect 16320 29986 16400 30000
rect 16320 29934 16334 29986
rect 16386 29934 16400 29986
rect 16320 29920 16400 29934
rect 16480 29986 16560 30000
rect 16480 29934 16494 29986
rect 16546 29934 16560 29986
rect 16480 29920 16560 29934
rect 16640 29986 16720 30000
rect 16640 29934 16654 29986
rect 16706 29934 16720 29986
rect 16640 29920 16720 29934
rect 16800 29986 16880 30000
rect 16800 29934 16814 29986
rect 16866 29934 16880 29986
rect 16800 29920 16880 29934
rect 16960 29986 17040 30000
rect 16960 29934 16974 29986
rect 17026 29934 17040 29986
rect 16960 29920 17040 29934
rect 17120 29986 17200 30000
rect 17120 29934 17134 29986
rect 17186 29934 17200 29986
rect 17120 29920 17200 29934
rect 17280 29986 17360 30000
rect 17280 29934 17294 29986
rect 17346 29934 17360 29986
rect 17280 29920 17360 29934
rect 17440 29986 17520 30000
rect 17440 29934 17454 29986
rect 17506 29934 17520 29986
rect 17440 29920 17520 29934
rect 17600 29986 17680 30000
rect 17600 29934 17614 29986
rect 17666 29934 17680 29986
rect 17600 29920 17680 29934
rect 17760 29986 17840 30000
rect 17760 29934 17774 29986
rect 17826 29934 17840 29986
rect 17760 29920 17840 29934
rect 17920 29986 18000 30000
rect 17920 29934 17934 29986
rect 17986 29934 18000 29986
rect 17920 29920 18000 29934
rect 18080 29986 18160 30000
rect 18080 29934 18094 29986
rect 18146 29934 18160 29986
rect 18080 29920 18160 29934
rect 18240 29986 18320 30000
rect 18240 29934 18254 29986
rect 18306 29934 18320 29986
rect 18240 29920 18320 29934
rect 18400 29986 18480 30000
rect 18400 29934 18414 29986
rect 18466 29934 18480 29986
rect 18400 29920 18480 29934
rect 18560 29986 18640 30000
rect 18560 29934 18574 29986
rect 18626 29934 18640 29986
rect 18560 29920 18640 29934
rect 18720 29986 18800 30000
rect 18720 29934 18734 29986
rect 18786 29934 18800 29986
rect 18720 29920 18800 29934
rect 18880 29986 18960 30000
rect 18880 29934 18894 29986
rect 18946 29934 18960 29986
rect 18880 29920 18960 29934
rect 23120 29986 23200 30000
rect 23120 29934 23134 29986
rect 23186 29934 23200 29986
rect 23120 29920 23200 29934
rect 23280 29986 23360 30000
rect 23280 29934 23294 29986
rect 23346 29934 23360 29986
rect 23280 29920 23360 29934
rect 23440 29986 23520 30000
rect 23440 29934 23454 29986
rect 23506 29934 23520 29986
rect 23440 29920 23520 29934
rect 23600 29986 23680 30000
rect 23600 29934 23614 29986
rect 23666 29934 23680 29986
rect 23600 29920 23680 29934
rect 23760 29986 23840 30000
rect 23760 29934 23774 29986
rect 23826 29934 23840 29986
rect 23760 29920 23840 29934
rect 23920 29986 24000 30000
rect 23920 29934 23934 29986
rect 23986 29934 24000 29986
rect 23920 29920 24000 29934
rect 24080 29986 24160 30000
rect 24080 29934 24094 29986
rect 24146 29934 24160 29986
rect 24080 29920 24160 29934
rect 24240 29986 24320 30000
rect 24240 29934 24254 29986
rect 24306 29934 24320 29986
rect 24240 29920 24320 29934
rect 24400 29986 24480 30000
rect 24400 29934 24414 29986
rect 24466 29934 24480 29986
rect 24400 29920 24480 29934
rect 24560 29986 24640 30000
rect 24560 29934 24574 29986
rect 24626 29934 24640 29986
rect 24560 29920 24640 29934
rect 24720 29986 24800 30000
rect 24720 29934 24734 29986
rect 24786 29934 24800 29986
rect 24720 29920 24800 29934
rect 24880 29986 24960 30000
rect 24880 29934 24894 29986
rect 24946 29934 24960 29986
rect 24880 29920 24960 29934
rect 25040 29986 25120 30000
rect 25040 29934 25054 29986
rect 25106 29934 25120 29986
rect 25040 29920 25120 29934
rect 25200 29986 25280 30000
rect 25200 29934 25214 29986
rect 25266 29934 25280 29986
rect 25200 29920 25280 29934
rect 25360 29986 25440 30000
rect 25360 29934 25374 29986
rect 25426 29934 25440 29986
rect 25360 29920 25440 29934
rect 25520 29986 25600 30000
rect 25520 29934 25534 29986
rect 25586 29934 25600 29986
rect 25520 29920 25600 29934
rect 25680 29986 25760 30000
rect 25680 29934 25694 29986
rect 25746 29934 25760 29986
rect 25680 29920 25760 29934
rect 25840 29986 25920 30000
rect 25840 29934 25854 29986
rect 25906 29934 25920 29986
rect 25840 29920 25920 29934
rect 26000 29986 26080 30000
rect 26000 29934 26014 29986
rect 26066 29934 26080 29986
rect 26000 29920 26080 29934
rect 26160 29986 26240 30000
rect 26160 29934 26174 29986
rect 26226 29934 26240 29986
rect 26160 29920 26240 29934
rect 26320 29986 26400 30000
rect 26320 29934 26334 29986
rect 26386 29934 26400 29986
rect 26320 29920 26400 29934
rect 26480 29986 26560 30000
rect 26480 29934 26494 29986
rect 26546 29934 26560 29986
rect 26480 29920 26560 29934
rect 26640 29986 26720 30000
rect 26640 29934 26654 29986
rect 26706 29934 26720 29986
rect 26640 29920 26720 29934
rect 26800 29986 26880 30000
rect 26800 29934 26814 29986
rect 26866 29934 26880 29986
rect 26800 29920 26880 29934
rect 26960 29986 27040 30000
rect 26960 29934 26974 29986
rect 27026 29934 27040 29986
rect 26960 29920 27040 29934
rect 27120 29986 27200 30000
rect 27120 29934 27134 29986
rect 27186 29934 27200 29986
rect 27120 29920 27200 29934
rect 27280 29986 27360 30000
rect 27280 29934 27294 29986
rect 27346 29934 27360 29986
rect 27280 29920 27360 29934
rect 27440 29986 27520 30000
rect 27440 29934 27454 29986
rect 27506 29934 27520 29986
rect 27440 29920 27520 29934
rect 27600 29986 27680 30000
rect 27600 29934 27614 29986
rect 27666 29934 27680 29986
rect 27600 29920 27680 29934
rect 27760 29986 27840 30000
rect 27760 29934 27774 29986
rect 27826 29934 27840 29986
rect 27760 29920 27840 29934
rect 27920 29986 28000 30000
rect 27920 29934 27934 29986
rect 27986 29934 28000 29986
rect 27920 29920 28000 29934
rect 28080 29986 28160 30000
rect 28080 29934 28094 29986
rect 28146 29934 28160 29986
rect 28080 29920 28160 29934
rect 28240 29986 28320 30000
rect 28240 29934 28254 29986
rect 28306 29934 28320 29986
rect 28240 29920 28320 29934
rect 28400 29986 28480 30000
rect 28400 29934 28414 29986
rect 28466 29934 28480 29986
rect 28400 29920 28480 29934
rect 28560 29986 28640 30000
rect 28560 29934 28574 29986
rect 28626 29934 28640 29986
rect 28560 29920 28640 29934
rect 28720 29986 28800 30000
rect 28720 29934 28734 29986
rect 28786 29934 28800 29986
rect 28720 29920 28800 29934
rect 28880 29986 28960 30000
rect 28880 29934 28894 29986
rect 28946 29934 28960 29986
rect 28880 29920 28960 29934
rect 29040 29986 29120 30000
rect 29040 29934 29054 29986
rect 29106 29934 29120 29986
rect 29040 29920 29120 29934
rect 29200 29986 29280 30000
rect 29200 29934 29214 29986
rect 29266 29934 29280 29986
rect 29200 29920 29280 29934
rect 29360 29986 29440 30000
rect 29360 29934 29374 29986
rect 29426 29934 29440 29986
rect 29360 29920 29440 29934
rect 33520 29986 33600 30000
rect 33520 29934 33534 29986
rect 33586 29934 33600 29986
rect 33520 29920 33600 29934
rect 33680 29986 33760 30000
rect 33680 29934 33694 29986
rect 33746 29934 33760 29986
rect 33680 29920 33760 29934
rect 33840 29986 33920 30000
rect 33840 29934 33854 29986
rect 33906 29934 33920 29986
rect 33840 29920 33920 29934
rect 34000 29986 34080 30000
rect 34000 29934 34014 29986
rect 34066 29934 34080 29986
rect 34000 29920 34080 29934
rect 34160 29986 34240 30000
rect 34160 29934 34174 29986
rect 34226 29934 34240 29986
rect 34160 29920 34240 29934
rect 34320 29986 34400 30000
rect 34320 29934 34334 29986
rect 34386 29934 34400 29986
rect 34320 29920 34400 29934
rect 34480 29986 34560 30000
rect 34480 29934 34494 29986
rect 34546 29934 34560 29986
rect 34480 29920 34560 29934
rect 34640 29986 34720 30000
rect 34640 29934 34654 29986
rect 34706 29934 34720 29986
rect 34640 29920 34720 29934
rect 34800 29986 34880 30000
rect 34800 29934 34814 29986
rect 34866 29934 34880 29986
rect 34800 29920 34880 29934
rect 34960 29986 35040 30000
rect 34960 29934 34974 29986
rect 35026 29934 35040 29986
rect 34960 29920 35040 29934
rect 35120 29986 35200 30000
rect 35120 29934 35134 29986
rect 35186 29934 35200 29986
rect 35120 29920 35200 29934
rect 35280 29986 35360 30000
rect 35280 29934 35294 29986
rect 35346 29934 35360 29986
rect 35280 29920 35360 29934
rect 35440 29986 35520 30000
rect 35440 29934 35454 29986
rect 35506 29934 35520 29986
rect 35440 29920 35520 29934
rect 35600 29986 35680 30000
rect 35600 29934 35614 29986
rect 35666 29934 35680 29986
rect 35600 29920 35680 29934
rect 35760 29986 35840 30000
rect 35760 29934 35774 29986
rect 35826 29934 35840 29986
rect 35760 29920 35840 29934
rect 35920 29986 36000 30000
rect 35920 29934 35934 29986
rect 35986 29934 36000 29986
rect 35920 29920 36000 29934
rect 36080 29986 36160 30000
rect 36080 29934 36094 29986
rect 36146 29934 36160 29986
rect 36080 29920 36160 29934
rect 36240 29986 36320 30000
rect 36240 29934 36254 29986
rect 36306 29934 36320 29986
rect 36240 29920 36320 29934
rect 36400 29986 36480 30000
rect 36400 29934 36414 29986
rect 36466 29934 36480 29986
rect 36400 29920 36480 29934
rect 36560 29986 36640 30000
rect 36560 29934 36574 29986
rect 36626 29934 36640 29986
rect 36560 29920 36640 29934
rect 36720 29986 36800 30000
rect 36720 29934 36734 29986
rect 36786 29934 36800 29986
rect 36720 29920 36800 29934
rect 36880 29986 36960 30000
rect 36880 29934 36894 29986
rect 36946 29934 36960 29986
rect 36880 29920 36960 29934
rect 37040 29986 37120 30000
rect 37040 29934 37054 29986
rect 37106 29934 37120 29986
rect 37040 29920 37120 29934
rect 37200 29986 37280 30000
rect 37200 29934 37214 29986
rect 37266 29934 37280 29986
rect 37200 29920 37280 29934
rect 37360 29986 37440 30000
rect 37360 29934 37374 29986
rect 37426 29934 37440 29986
rect 37360 29920 37440 29934
rect 37520 29986 37600 30000
rect 37520 29934 37534 29986
rect 37586 29934 37600 29986
rect 37520 29920 37600 29934
rect 37680 29986 37760 30000
rect 37680 29934 37694 29986
rect 37746 29934 37760 29986
rect 37680 29920 37760 29934
rect 37840 29986 37920 30000
rect 37840 29934 37854 29986
rect 37906 29934 37920 29986
rect 37840 29920 37920 29934
rect 38000 29986 38080 30000
rect 38000 29934 38014 29986
rect 38066 29934 38080 29986
rect 38000 29920 38080 29934
rect 38160 29986 38240 30000
rect 38160 29934 38174 29986
rect 38226 29934 38240 29986
rect 38160 29920 38240 29934
rect 38320 29986 38400 30000
rect 38320 29934 38334 29986
rect 38386 29934 38400 29986
rect 38320 29920 38400 29934
rect 38480 29986 38560 30000
rect 38480 29934 38494 29986
rect 38546 29934 38560 29986
rect 38480 29920 38560 29934
rect 38640 29986 38720 30000
rect 38640 29934 38654 29986
rect 38706 29934 38720 29986
rect 38640 29920 38720 29934
rect 38800 29986 38880 30000
rect 38800 29934 38814 29986
rect 38866 29934 38880 29986
rect 38800 29920 38880 29934
rect 38960 29986 39040 30000
rect 38960 29934 38974 29986
rect 39026 29934 39040 29986
rect 38960 29920 39040 29934
rect 39120 29986 39200 30000
rect 39120 29934 39134 29986
rect 39186 29934 39200 29986
rect 39120 29920 39200 29934
rect 39280 29986 39360 30000
rect 39280 29934 39294 29986
rect 39346 29934 39360 29986
rect 39280 29920 39360 29934
rect 39440 29986 39520 30000
rect 39440 29934 39454 29986
rect 39506 29934 39520 29986
rect 39440 29920 39520 29934
rect 39600 29986 39680 30000
rect 39600 29934 39614 29986
rect 39666 29934 39680 29986
rect 39600 29920 39680 29934
rect 39760 29986 39840 30000
rect 39760 29934 39774 29986
rect 39826 29934 39840 29986
rect 39760 29920 39840 29934
rect 39920 29986 40000 30000
rect 39920 29934 39934 29986
rect 39986 29934 40000 29986
rect 39920 29920 40000 29934
rect 40080 29986 40160 30000
rect 40080 29934 40094 29986
rect 40146 29934 40160 29986
rect 40080 29920 40160 29934
rect 40240 29986 40320 30000
rect 40240 29934 40254 29986
rect 40306 29934 40320 29986
rect 40240 29920 40320 29934
rect 40400 29986 40480 30000
rect 40400 29934 40414 29986
rect 40466 29934 40480 29986
rect 40400 29920 40480 29934
rect 40560 29986 40640 30000
rect 40560 29934 40574 29986
rect 40626 29934 40640 29986
rect 40560 29920 40640 29934
rect 40720 29986 40800 30000
rect 40720 29934 40734 29986
rect 40786 29934 40800 29986
rect 40720 29920 40800 29934
rect 40880 29986 40960 30000
rect 40880 29934 40894 29986
rect 40946 29934 40960 29986
rect 40880 29920 40960 29934
rect 41040 29986 41120 30000
rect 41040 29934 41054 29986
rect 41106 29934 41120 29986
rect 41040 29920 41120 29934
rect 41200 29986 41280 30000
rect 41200 29934 41214 29986
rect 41266 29934 41280 29986
rect 41200 29920 41280 29934
rect 41360 29986 41440 30000
rect 41360 29934 41374 29986
rect 41426 29934 41440 29986
rect 41360 29920 41440 29934
rect 41520 29986 41600 30000
rect 41520 29934 41534 29986
rect 41586 29934 41600 29986
rect 41520 29920 41600 29934
rect 41680 29986 41760 30000
rect 41680 29934 41694 29986
rect 41746 29934 41760 29986
rect 41680 29920 41760 29934
rect 41840 29986 41920 30000
rect 41840 29934 41854 29986
rect 41906 29934 41920 29986
rect 41840 29920 41920 29934
rect 0 29826 80 29840
rect 0 29774 14 29826
rect 66 29774 80 29826
rect 0 29760 80 29774
rect 160 29826 240 29840
rect 160 29774 174 29826
rect 226 29774 240 29826
rect 160 29760 240 29774
rect 320 29826 400 29840
rect 320 29774 334 29826
rect 386 29774 400 29826
rect 320 29760 400 29774
rect 480 29826 560 29840
rect 480 29774 494 29826
rect 546 29774 560 29826
rect 480 29760 560 29774
rect 640 29826 720 29840
rect 640 29774 654 29826
rect 706 29774 720 29826
rect 640 29760 720 29774
rect 800 29826 880 29840
rect 800 29774 814 29826
rect 866 29774 880 29826
rect 800 29760 880 29774
rect 960 29826 1040 29840
rect 960 29774 974 29826
rect 1026 29774 1040 29826
rect 960 29760 1040 29774
rect 1120 29826 1200 29840
rect 1120 29774 1134 29826
rect 1186 29774 1200 29826
rect 1120 29760 1200 29774
rect 1280 29826 1360 29840
rect 1280 29774 1294 29826
rect 1346 29774 1360 29826
rect 1280 29760 1360 29774
rect 1440 29826 1520 29840
rect 1440 29774 1454 29826
rect 1506 29774 1520 29826
rect 1440 29760 1520 29774
rect 1600 29826 1680 29840
rect 1600 29774 1614 29826
rect 1666 29774 1680 29826
rect 1600 29760 1680 29774
rect 1760 29826 1840 29840
rect 1760 29774 1774 29826
rect 1826 29774 1840 29826
rect 1760 29760 1840 29774
rect 1920 29826 2000 29840
rect 1920 29774 1934 29826
rect 1986 29774 2000 29826
rect 1920 29760 2000 29774
rect 2080 29826 2160 29840
rect 2080 29774 2094 29826
rect 2146 29774 2160 29826
rect 2080 29760 2160 29774
rect 2240 29826 2320 29840
rect 2240 29774 2254 29826
rect 2306 29774 2320 29826
rect 2240 29760 2320 29774
rect 2400 29826 2480 29840
rect 2400 29774 2414 29826
rect 2466 29774 2480 29826
rect 2400 29760 2480 29774
rect 2560 29826 2640 29840
rect 2560 29774 2574 29826
rect 2626 29774 2640 29826
rect 2560 29760 2640 29774
rect 2720 29826 2800 29840
rect 2720 29774 2734 29826
rect 2786 29774 2800 29826
rect 2720 29760 2800 29774
rect 2880 29826 2960 29840
rect 2880 29774 2894 29826
rect 2946 29774 2960 29826
rect 2880 29760 2960 29774
rect 3040 29826 3120 29840
rect 3040 29774 3054 29826
rect 3106 29774 3120 29826
rect 3040 29760 3120 29774
rect 3200 29826 3280 29840
rect 3200 29774 3214 29826
rect 3266 29774 3280 29826
rect 3200 29760 3280 29774
rect 3360 29826 3440 29840
rect 3360 29774 3374 29826
rect 3426 29774 3440 29826
rect 3360 29760 3440 29774
rect 3520 29826 3600 29840
rect 3520 29774 3534 29826
rect 3586 29774 3600 29826
rect 3520 29760 3600 29774
rect 3680 29826 3760 29840
rect 3680 29774 3694 29826
rect 3746 29774 3760 29826
rect 3680 29760 3760 29774
rect 3840 29826 3920 29840
rect 3840 29774 3854 29826
rect 3906 29774 3920 29826
rect 3840 29760 3920 29774
rect 4000 29826 4080 29840
rect 4000 29774 4014 29826
rect 4066 29774 4080 29826
rect 4000 29760 4080 29774
rect 4160 29826 4240 29840
rect 4160 29774 4174 29826
rect 4226 29774 4240 29826
rect 4160 29760 4240 29774
rect 4320 29826 4400 29840
rect 4320 29774 4334 29826
rect 4386 29774 4400 29826
rect 4320 29760 4400 29774
rect 4480 29826 4560 29840
rect 4480 29774 4494 29826
rect 4546 29774 4560 29826
rect 4480 29760 4560 29774
rect 4640 29826 4720 29840
rect 4640 29774 4654 29826
rect 4706 29774 4720 29826
rect 4640 29760 4720 29774
rect 4800 29826 4880 29840
rect 4800 29774 4814 29826
rect 4866 29774 4880 29826
rect 4800 29760 4880 29774
rect 4960 29826 5040 29840
rect 4960 29774 4974 29826
rect 5026 29774 5040 29826
rect 4960 29760 5040 29774
rect 5120 29826 5200 29840
rect 5120 29774 5134 29826
rect 5186 29774 5200 29826
rect 5120 29760 5200 29774
rect 5280 29826 5360 29840
rect 5280 29774 5294 29826
rect 5346 29774 5360 29826
rect 5280 29760 5360 29774
rect 5440 29826 5520 29840
rect 5440 29774 5454 29826
rect 5506 29774 5520 29826
rect 5440 29760 5520 29774
rect 5600 29826 5680 29840
rect 5600 29774 5614 29826
rect 5666 29774 5680 29826
rect 5600 29760 5680 29774
rect 5760 29826 5840 29840
rect 5760 29774 5774 29826
rect 5826 29774 5840 29826
rect 5760 29760 5840 29774
rect 5920 29826 6000 29840
rect 5920 29774 5934 29826
rect 5986 29774 6000 29826
rect 5920 29760 6000 29774
rect 6080 29826 6160 29840
rect 6080 29774 6094 29826
rect 6146 29774 6160 29826
rect 6080 29760 6160 29774
rect 6240 29826 6320 29840
rect 6240 29774 6254 29826
rect 6306 29774 6320 29826
rect 6240 29760 6320 29774
rect 6400 29826 6480 29840
rect 6400 29774 6414 29826
rect 6466 29774 6480 29826
rect 6400 29760 6480 29774
rect 6560 29826 6640 29840
rect 6560 29774 6574 29826
rect 6626 29774 6640 29826
rect 6560 29760 6640 29774
rect 6720 29826 6800 29840
rect 6720 29774 6734 29826
rect 6786 29774 6800 29826
rect 6720 29760 6800 29774
rect 6880 29826 6960 29840
rect 6880 29774 6894 29826
rect 6946 29774 6960 29826
rect 6880 29760 6960 29774
rect 7040 29826 7120 29840
rect 7040 29774 7054 29826
rect 7106 29774 7120 29826
rect 7040 29760 7120 29774
rect 7200 29826 7280 29840
rect 7200 29774 7214 29826
rect 7266 29774 7280 29826
rect 7200 29760 7280 29774
rect 7360 29826 7440 29840
rect 7360 29774 7374 29826
rect 7426 29774 7440 29826
rect 7360 29760 7440 29774
rect 7520 29826 7600 29840
rect 7520 29774 7534 29826
rect 7586 29774 7600 29826
rect 7520 29760 7600 29774
rect 7680 29826 7760 29840
rect 7680 29774 7694 29826
rect 7746 29774 7760 29826
rect 7680 29760 7760 29774
rect 7840 29826 7920 29840
rect 7840 29774 7854 29826
rect 7906 29774 7920 29826
rect 7840 29760 7920 29774
rect 8000 29826 8080 29840
rect 8000 29774 8014 29826
rect 8066 29774 8080 29826
rect 8000 29760 8080 29774
rect 8160 29826 8240 29840
rect 8160 29774 8174 29826
rect 8226 29774 8240 29826
rect 8160 29760 8240 29774
rect 8320 29826 8400 29840
rect 8320 29774 8334 29826
rect 8386 29774 8400 29826
rect 8320 29760 8400 29774
rect 12480 29826 12560 29840
rect 12480 29774 12494 29826
rect 12546 29774 12560 29826
rect 12480 29760 12560 29774
rect 12640 29826 12720 29840
rect 12640 29774 12654 29826
rect 12706 29774 12720 29826
rect 12640 29760 12720 29774
rect 12800 29826 12880 29840
rect 12800 29774 12814 29826
rect 12866 29774 12880 29826
rect 12800 29760 12880 29774
rect 12960 29826 13040 29840
rect 12960 29774 12974 29826
rect 13026 29774 13040 29826
rect 12960 29760 13040 29774
rect 13120 29826 13200 29840
rect 13120 29774 13134 29826
rect 13186 29774 13200 29826
rect 13120 29760 13200 29774
rect 13280 29826 13360 29840
rect 13280 29774 13294 29826
rect 13346 29774 13360 29826
rect 13280 29760 13360 29774
rect 13440 29826 13520 29840
rect 13440 29774 13454 29826
rect 13506 29774 13520 29826
rect 13440 29760 13520 29774
rect 13600 29826 13680 29840
rect 13600 29774 13614 29826
rect 13666 29774 13680 29826
rect 13600 29760 13680 29774
rect 13760 29826 13840 29840
rect 13760 29774 13774 29826
rect 13826 29774 13840 29826
rect 13760 29760 13840 29774
rect 13920 29826 14000 29840
rect 13920 29774 13934 29826
rect 13986 29774 14000 29826
rect 13920 29760 14000 29774
rect 14080 29826 14160 29840
rect 14080 29774 14094 29826
rect 14146 29774 14160 29826
rect 14080 29760 14160 29774
rect 14240 29826 14320 29840
rect 14240 29774 14254 29826
rect 14306 29774 14320 29826
rect 14240 29760 14320 29774
rect 14400 29826 14480 29840
rect 14400 29774 14414 29826
rect 14466 29774 14480 29826
rect 14400 29760 14480 29774
rect 14560 29826 14640 29840
rect 14560 29774 14574 29826
rect 14626 29774 14640 29826
rect 14560 29760 14640 29774
rect 14720 29826 14800 29840
rect 14720 29774 14734 29826
rect 14786 29774 14800 29826
rect 14720 29760 14800 29774
rect 14880 29826 14960 29840
rect 14880 29774 14894 29826
rect 14946 29774 14960 29826
rect 14880 29760 14960 29774
rect 15040 29826 15120 29840
rect 15040 29774 15054 29826
rect 15106 29774 15120 29826
rect 15040 29760 15120 29774
rect 15200 29826 15280 29840
rect 15200 29774 15214 29826
rect 15266 29774 15280 29826
rect 15200 29760 15280 29774
rect 15360 29826 15440 29840
rect 15360 29774 15374 29826
rect 15426 29774 15440 29826
rect 15360 29760 15440 29774
rect 15520 29826 15600 29840
rect 15520 29774 15534 29826
rect 15586 29774 15600 29826
rect 15520 29760 15600 29774
rect 15680 29826 15760 29840
rect 15680 29774 15694 29826
rect 15746 29774 15760 29826
rect 15680 29760 15760 29774
rect 15840 29826 15920 29840
rect 15840 29774 15854 29826
rect 15906 29774 15920 29826
rect 15840 29760 15920 29774
rect 16000 29826 16080 29840
rect 16000 29774 16014 29826
rect 16066 29774 16080 29826
rect 16000 29760 16080 29774
rect 16160 29826 16240 29840
rect 16160 29774 16174 29826
rect 16226 29774 16240 29826
rect 16160 29760 16240 29774
rect 16320 29826 16400 29840
rect 16320 29774 16334 29826
rect 16386 29774 16400 29826
rect 16320 29760 16400 29774
rect 16480 29826 16560 29840
rect 16480 29774 16494 29826
rect 16546 29774 16560 29826
rect 16480 29760 16560 29774
rect 16640 29826 16720 29840
rect 16640 29774 16654 29826
rect 16706 29774 16720 29826
rect 16640 29760 16720 29774
rect 16800 29826 16880 29840
rect 16800 29774 16814 29826
rect 16866 29774 16880 29826
rect 16800 29760 16880 29774
rect 16960 29826 17040 29840
rect 16960 29774 16974 29826
rect 17026 29774 17040 29826
rect 16960 29760 17040 29774
rect 17120 29826 17200 29840
rect 17120 29774 17134 29826
rect 17186 29774 17200 29826
rect 17120 29760 17200 29774
rect 17280 29826 17360 29840
rect 17280 29774 17294 29826
rect 17346 29774 17360 29826
rect 17280 29760 17360 29774
rect 17440 29826 17520 29840
rect 17440 29774 17454 29826
rect 17506 29774 17520 29826
rect 17440 29760 17520 29774
rect 17600 29826 17680 29840
rect 17600 29774 17614 29826
rect 17666 29774 17680 29826
rect 17600 29760 17680 29774
rect 17760 29826 17840 29840
rect 17760 29774 17774 29826
rect 17826 29774 17840 29826
rect 17760 29760 17840 29774
rect 17920 29826 18000 29840
rect 17920 29774 17934 29826
rect 17986 29774 18000 29826
rect 17920 29760 18000 29774
rect 18080 29826 18160 29840
rect 18080 29774 18094 29826
rect 18146 29774 18160 29826
rect 18080 29760 18160 29774
rect 18240 29826 18320 29840
rect 18240 29774 18254 29826
rect 18306 29774 18320 29826
rect 18240 29760 18320 29774
rect 18400 29826 18480 29840
rect 18400 29774 18414 29826
rect 18466 29774 18480 29826
rect 18400 29760 18480 29774
rect 18560 29826 18640 29840
rect 18560 29774 18574 29826
rect 18626 29774 18640 29826
rect 18560 29760 18640 29774
rect 18720 29826 18800 29840
rect 18720 29774 18734 29826
rect 18786 29774 18800 29826
rect 18720 29760 18800 29774
rect 18880 29826 18960 29840
rect 18880 29774 18894 29826
rect 18946 29774 18960 29826
rect 18880 29760 18960 29774
rect 23120 29826 23200 29840
rect 23120 29774 23134 29826
rect 23186 29774 23200 29826
rect 23120 29760 23200 29774
rect 23280 29826 23360 29840
rect 23280 29774 23294 29826
rect 23346 29774 23360 29826
rect 23280 29760 23360 29774
rect 23440 29826 23520 29840
rect 23440 29774 23454 29826
rect 23506 29774 23520 29826
rect 23440 29760 23520 29774
rect 23600 29826 23680 29840
rect 23600 29774 23614 29826
rect 23666 29774 23680 29826
rect 23600 29760 23680 29774
rect 23760 29826 23840 29840
rect 23760 29774 23774 29826
rect 23826 29774 23840 29826
rect 23760 29760 23840 29774
rect 23920 29826 24000 29840
rect 23920 29774 23934 29826
rect 23986 29774 24000 29826
rect 23920 29760 24000 29774
rect 24080 29826 24160 29840
rect 24080 29774 24094 29826
rect 24146 29774 24160 29826
rect 24080 29760 24160 29774
rect 24240 29826 24320 29840
rect 24240 29774 24254 29826
rect 24306 29774 24320 29826
rect 24240 29760 24320 29774
rect 24400 29826 24480 29840
rect 24400 29774 24414 29826
rect 24466 29774 24480 29826
rect 24400 29760 24480 29774
rect 24560 29826 24640 29840
rect 24560 29774 24574 29826
rect 24626 29774 24640 29826
rect 24560 29760 24640 29774
rect 24720 29826 24800 29840
rect 24720 29774 24734 29826
rect 24786 29774 24800 29826
rect 24720 29760 24800 29774
rect 24880 29826 24960 29840
rect 24880 29774 24894 29826
rect 24946 29774 24960 29826
rect 24880 29760 24960 29774
rect 25040 29826 25120 29840
rect 25040 29774 25054 29826
rect 25106 29774 25120 29826
rect 25040 29760 25120 29774
rect 25200 29826 25280 29840
rect 25200 29774 25214 29826
rect 25266 29774 25280 29826
rect 25200 29760 25280 29774
rect 25360 29826 25440 29840
rect 25360 29774 25374 29826
rect 25426 29774 25440 29826
rect 25360 29760 25440 29774
rect 25520 29826 25600 29840
rect 25520 29774 25534 29826
rect 25586 29774 25600 29826
rect 25520 29760 25600 29774
rect 25680 29826 25760 29840
rect 25680 29774 25694 29826
rect 25746 29774 25760 29826
rect 25680 29760 25760 29774
rect 25840 29826 25920 29840
rect 25840 29774 25854 29826
rect 25906 29774 25920 29826
rect 25840 29760 25920 29774
rect 26000 29826 26080 29840
rect 26000 29774 26014 29826
rect 26066 29774 26080 29826
rect 26000 29760 26080 29774
rect 26160 29826 26240 29840
rect 26160 29774 26174 29826
rect 26226 29774 26240 29826
rect 26160 29760 26240 29774
rect 26320 29826 26400 29840
rect 26320 29774 26334 29826
rect 26386 29774 26400 29826
rect 26320 29760 26400 29774
rect 26480 29826 26560 29840
rect 26480 29774 26494 29826
rect 26546 29774 26560 29826
rect 26480 29760 26560 29774
rect 26640 29826 26720 29840
rect 26640 29774 26654 29826
rect 26706 29774 26720 29826
rect 26640 29760 26720 29774
rect 26800 29826 26880 29840
rect 26800 29774 26814 29826
rect 26866 29774 26880 29826
rect 26800 29760 26880 29774
rect 26960 29826 27040 29840
rect 26960 29774 26974 29826
rect 27026 29774 27040 29826
rect 26960 29760 27040 29774
rect 27120 29826 27200 29840
rect 27120 29774 27134 29826
rect 27186 29774 27200 29826
rect 27120 29760 27200 29774
rect 27280 29826 27360 29840
rect 27280 29774 27294 29826
rect 27346 29774 27360 29826
rect 27280 29760 27360 29774
rect 27440 29826 27520 29840
rect 27440 29774 27454 29826
rect 27506 29774 27520 29826
rect 27440 29760 27520 29774
rect 27600 29826 27680 29840
rect 27600 29774 27614 29826
rect 27666 29774 27680 29826
rect 27600 29760 27680 29774
rect 27760 29826 27840 29840
rect 27760 29774 27774 29826
rect 27826 29774 27840 29826
rect 27760 29760 27840 29774
rect 27920 29826 28000 29840
rect 27920 29774 27934 29826
rect 27986 29774 28000 29826
rect 27920 29760 28000 29774
rect 28080 29826 28160 29840
rect 28080 29774 28094 29826
rect 28146 29774 28160 29826
rect 28080 29760 28160 29774
rect 28240 29826 28320 29840
rect 28240 29774 28254 29826
rect 28306 29774 28320 29826
rect 28240 29760 28320 29774
rect 28400 29826 28480 29840
rect 28400 29774 28414 29826
rect 28466 29774 28480 29826
rect 28400 29760 28480 29774
rect 28560 29826 28640 29840
rect 28560 29774 28574 29826
rect 28626 29774 28640 29826
rect 28560 29760 28640 29774
rect 28720 29826 28800 29840
rect 28720 29774 28734 29826
rect 28786 29774 28800 29826
rect 28720 29760 28800 29774
rect 28880 29826 28960 29840
rect 28880 29774 28894 29826
rect 28946 29774 28960 29826
rect 28880 29760 28960 29774
rect 29040 29826 29120 29840
rect 29040 29774 29054 29826
rect 29106 29774 29120 29826
rect 29040 29760 29120 29774
rect 29200 29826 29280 29840
rect 29200 29774 29214 29826
rect 29266 29774 29280 29826
rect 29200 29760 29280 29774
rect 29360 29826 29440 29840
rect 29360 29774 29374 29826
rect 29426 29774 29440 29826
rect 29360 29760 29440 29774
rect 33520 29826 33600 29840
rect 33520 29774 33534 29826
rect 33586 29774 33600 29826
rect 33520 29760 33600 29774
rect 33680 29826 33760 29840
rect 33680 29774 33694 29826
rect 33746 29774 33760 29826
rect 33680 29760 33760 29774
rect 33840 29826 33920 29840
rect 33840 29774 33854 29826
rect 33906 29774 33920 29826
rect 33840 29760 33920 29774
rect 34000 29826 34080 29840
rect 34000 29774 34014 29826
rect 34066 29774 34080 29826
rect 34000 29760 34080 29774
rect 34160 29826 34240 29840
rect 34160 29774 34174 29826
rect 34226 29774 34240 29826
rect 34160 29760 34240 29774
rect 34320 29826 34400 29840
rect 34320 29774 34334 29826
rect 34386 29774 34400 29826
rect 34320 29760 34400 29774
rect 34480 29826 34560 29840
rect 34480 29774 34494 29826
rect 34546 29774 34560 29826
rect 34480 29760 34560 29774
rect 34640 29826 34720 29840
rect 34640 29774 34654 29826
rect 34706 29774 34720 29826
rect 34640 29760 34720 29774
rect 34800 29826 34880 29840
rect 34800 29774 34814 29826
rect 34866 29774 34880 29826
rect 34800 29760 34880 29774
rect 34960 29826 35040 29840
rect 34960 29774 34974 29826
rect 35026 29774 35040 29826
rect 34960 29760 35040 29774
rect 35120 29826 35200 29840
rect 35120 29774 35134 29826
rect 35186 29774 35200 29826
rect 35120 29760 35200 29774
rect 35280 29826 35360 29840
rect 35280 29774 35294 29826
rect 35346 29774 35360 29826
rect 35280 29760 35360 29774
rect 35440 29826 35520 29840
rect 35440 29774 35454 29826
rect 35506 29774 35520 29826
rect 35440 29760 35520 29774
rect 35600 29826 35680 29840
rect 35600 29774 35614 29826
rect 35666 29774 35680 29826
rect 35600 29760 35680 29774
rect 35760 29826 35840 29840
rect 35760 29774 35774 29826
rect 35826 29774 35840 29826
rect 35760 29760 35840 29774
rect 35920 29826 36000 29840
rect 35920 29774 35934 29826
rect 35986 29774 36000 29826
rect 35920 29760 36000 29774
rect 36080 29826 36160 29840
rect 36080 29774 36094 29826
rect 36146 29774 36160 29826
rect 36080 29760 36160 29774
rect 36240 29826 36320 29840
rect 36240 29774 36254 29826
rect 36306 29774 36320 29826
rect 36240 29760 36320 29774
rect 36400 29826 36480 29840
rect 36400 29774 36414 29826
rect 36466 29774 36480 29826
rect 36400 29760 36480 29774
rect 36560 29826 36640 29840
rect 36560 29774 36574 29826
rect 36626 29774 36640 29826
rect 36560 29760 36640 29774
rect 36720 29826 36800 29840
rect 36720 29774 36734 29826
rect 36786 29774 36800 29826
rect 36720 29760 36800 29774
rect 36880 29826 36960 29840
rect 36880 29774 36894 29826
rect 36946 29774 36960 29826
rect 36880 29760 36960 29774
rect 37040 29826 37120 29840
rect 37040 29774 37054 29826
rect 37106 29774 37120 29826
rect 37040 29760 37120 29774
rect 37200 29826 37280 29840
rect 37200 29774 37214 29826
rect 37266 29774 37280 29826
rect 37200 29760 37280 29774
rect 37360 29826 37440 29840
rect 37360 29774 37374 29826
rect 37426 29774 37440 29826
rect 37360 29760 37440 29774
rect 37520 29826 37600 29840
rect 37520 29774 37534 29826
rect 37586 29774 37600 29826
rect 37520 29760 37600 29774
rect 37680 29826 37760 29840
rect 37680 29774 37694 29826
rect 37746 29774 37760 29826
rect 37680 29760 37760 29774
rect 37840 29826 37920 29840
rect 37840 29774 37854 29826
rect 37906 29774 37920 29826
rect 37840 29760 37920 29774
rect 38000 29826 38080 29840
rect 38000 29774 38014 29826
rect 38066 29774 38080 29826
rect 38000 29760 38080 29774
rect 38160 29826 38240 29840
rect 38160 29774 38174 29826
rect 38226 29774 38240 29826
rect 38160 29760 38240 29774
rect 38320 29826 38400 29840
rect 38320 29774 38334 29826
rect 38386 29774 38400 29826
rect 38320 29760 38400 29774
rect 38480 29826 38560 29840
rect 38480 29774 38494 29826
rect 38546 29774 38560 29826
rect 38480 29760 38560 29774
rect 38640 29826 38720 29840
rect 38640 29774 38654 29826
rect 38706 29774 38720 29826
rect 38640 29760 38720 29774
rect 38800 29826 38880 29840
rect 38800 29774 38814 29826
rect 38866 29774 38880 29826
rect 38800 29760 38880 29774
rect 38960 29826 39040 29840
rect 38960 29774 38974 29826
rect 39026 29774 39040 29826
rect 38960 29760 39040 29774
rect 39120 29826 39200 29840
rect 39120 29774 39134 29826
rect 39186 29774 39200 29826
rect 39120 29760 39200 29774
rect 39280 29826 39360 29840
rect 39280 29774 39294 29826
rect 39346 29774 39360 29826
rect 39280 29760 39360 29774
rect 39440 29826 39520 29840
rect 39440 29774 39454 29826
rect 39506 29774 39520 29826
rect 39440 29760 39520 29774
rect 39600 29826 39680 29840
rect 39600 29774 39614 29826
rect 39666 29774 39680 29826
rect 39600 29760 39680 29774
rect 39760 29826 39840 29840
rect 39760 29774 39774 29826
rect 39826 29774 39840 29826
rect 39760 29760 39840 29774
rect 39920 29826 40000 29840
rect 39920 29774 39934 29826
rect 39986 29774 40000 29826
rect 39920 29760 40000 29774
rect 40080 29826 40160 29840
rect 40080 29774 40094 29826
rect 40146 29774 40160 29826
rect 40080 29760 40160 29774
rect 40240 29826 40320 29840
rect 40240 29774 40254 29826
rect 40306 29774 40320 29826
rect 40240 29760 40320 29774
rect 40400 29826 40480 29840
rect 40400 29774 40414 29826
rect 40466 29774 40480 29826
rect 40400 29760 40480 29774
rect 40560 29826 40640 29840
rect 40560 29774 40574 29826
rect 40626 29774 40640 29826
rect 40560 29760 40640 29774
rect 40720 29826 40800 29840
rect 40720 29774 40734 29826
rect 40786 29774 40800 29826
rect 40720 29760 40800 29774
rect 40880 29826 40960 29840
rect 40880 29774 40894 29826
rect 40946 29774 40960 29826
rect 40880 29760 40960 29774
rect 41040 29826 41120 29840
rect 41040 29774 41054 29826
rect 41106 29774 41120 29826
rect 41040 29760 41120 29774
rect 41200 29826 41280 29840
rect 41200 29774 41214 29826
rect 41266 29774 41280 29826
rect 41200 29760 41280 29774
rect 41360 29826 41440 29840
rect 41360 29774 41374 29826
rect 41426 29774 41440 29826
rect 41360 29760 41440 29774
rect 41520 29826 41600 29840
rect 41520 29774 41534 29826
rect 41586 29774 41600 29826
rect 41520 29760 41600 29774
rect 41680 29826 41760 29840
rect 41680 29774 41694 29826
rect 41746 29774 41760 29826
rect 41680 29760 41760 29774
rect 41840 29826 41920 29840
rect 41840 29774 41854 29826
rect 41906 29774 41920 29826
rect 41840 29760 41920 29774
rect 0 29506 80 29520
rect 0 29454 14 29506
rect 66 29454 80 29506
rect 0 29440 80 29454
rect 160 29506 240 29520
rect 160 29454 174 29506
rect 226 29454 240 29506
rect 160 29440 240 29454
rect 320 29506 400 29520
rect 320 29454 334 29506
rect 386 29454 400 29506
rect 320 29440 400 29454
rect 480 29506 560 29520
rect 480 29454 494 29506
rect 546 29454 560 29506
rect 480 29440 560 29454
rect 640 29506 720 29520
rect 640 29454 654 29506
rect 706 29454 720 29506
rect 640 29440 720 29454
rect 800 29506 880 29520
rect 800 29454 814 29506
rect 866 29454 880 29506
rect 800 29440 880 29454
rect 960 29506 1040 29520
rect 960 29454 974 29506
rect 1026 29454 1040 29506
rect 960 29440 1040 29454
rect 1120 29506 1200 29520
rect 1120 29454 1134 29506
rect 1186 29454 1200 29506
rect 1120 29440 1200 29454
rect 1280 29506 1360 29520
rect 1280 29454 1294 29506
rect 1346 29454 1360 29506
rect 1280 29440 1360 29454
rect 1440 29506 1520 29520
rect 1440 29454 1454 29506
rect 1506 29454 1520 29506
rect 1440 29440 1520 29454
rect 1600 29506 1680 29520
rect 1600 29454 1614 29506
rect 1666 29454 1680 29506
rect 1600 29440 1680 29454
rect 1760 29506 1840 29520
rect 1760 29454 1774 29506
rect 1826 29454 1840 29506
rect 1760 29440 1840 29454
rect 1920 29506 2000 29520
rect 1920 29454 1934 29506
rect 1986 29454 2000 29506
rect 1920 29440 2000 29454
rect 2080 29506 2160 29520
rect 2080 29454 2094 29506
rect 2146 29454 2160 29506
rect 2080 29440 2160 29454
rect 2240 29506 2320 29520
rect 2240 29454 2254 29506
rect 2306 29454 2320 29506
rect 2240 29440 2320 29454
rect 2400 29506 2480 29520
rect 2400 29454 2414 29506
rect 2466 29454 2480 29506
rect 2400 29440 2480 29454
rect 2560 29506 2640 29520
rect 2560 29454 2574 29506
rect 2626 29454 2640 29506
rect 2560 29440 2640 29454
rect 2720 29506 2800 29520
rect 2720 29454 2734 29506
rect 2786 29454 2800 29506
rect 2720 29440 2800 29454
rect 2880 29506 2960 29520
rect 2880 29454 2894 29506
rect 2946 29454 2960 29506
rect 2880 29440 2960 29454
rect 3040 29506 3120 29520
rect 3040 29454 3054 29506
rect 3106 29454 3120 29506
rect 3040 29440 3120 29454
rect 3200 29506 3280 29520
rect 3200 29454 3214 29506
rect 3266 29454 3280 29506
rect 3200 29440 3280 29454
rect 3360 29506 3440 29520
rect 3360 29454 3374 29506
rect 3426 29454 3440 29506
rect 3360 29440 3440 29454
rect 3520 29506 3600 29520
rect 3520 29454 3534 29506
rect 3586 29454 3600 29506
rect 3520 29440 3600 29454
rect 3680 29506 3760 29520
rect 3680 29454 3694 29506
rect 3746 29454 3760 29506
rect 3680 29440 3760 29454
rect 3840 29506 3920 29520
rect 3840 29454 3854 29506
rect 3906 29454 3920 29506
rect 3840 29440 3920 29454
rect 4000 29506 4080 29520
rect 4000 29454 4014 29506
rect 4066 29454 4080 29506
rect 4000 29440 4080 29454
rect 4160 29506 4240 29520
rect 4160 29454 4174 29506
rect 4226 29454 4240 29506
rect 4160 29440 4240 29454
rect 4320 29506 4400 29520
rect 4320 29454 4334 29506
rect 4386 29454 4400 29506
rect 4320 29440 4400 29454
rect 4480 29506 4560 29520
rect 4480 29454 4494 29506
rect 4546 29454 4560 29506
rect 4480 29440 4560 29454
rect 4640 29506 4720 29520
rect 4640 29454 4654 29506
rect 4706 29454 4720 29506
rect 4640 29440 4720 29454
rect 4800 29506 4880 29520
rect 4800 29454 4814 29506
rect 4866 29454 4880 29506
rect 4800 29440 4880 29454
rect 4960 29506 5040 29520
rect 4960 29454 4974 29506
rect 5026 29454 5040 29506
rect 4960 29440 5040 29454
rect 5120 29506 5200 29520
rect 5120 29454 5134 29506
rect 5186 29454 5200 29506
rect 5120 29440 5200 29454
rect 5280 29506 5360 29520
rect 5280 29454 5294 29506
rect 5346 29454 5360 29506
rect 5280 29440 5360 29454
rect 5440 29506 5520 29520
rect 5440 29454 5454 29506
rect 5506 29454 5520 29506
rect 5440 29440 5520 29454
rect 5600 29506 5680 29520
rect 5600 29454 5614 29506
rect 5666 29454 5680 29506
rect 5600 29440 5680 29454
rect 5760 29506 5840 29520
rect 5760 29454 5774 29506
rect 5826 29454 5840 29506
rect 5760 29440 5840 29454
rect 5920 29506 6000 29520
rect 5920 29454 5934 29506
rect 5986 29454 6000 29506
rect 5920 29440 6000 29454
rect 6080 29506 6160 29520
rect 6080 29454 6094 29506
rect 6146 29454 6160 29506
rect 6080 29440 6160 29454
rect 6240 29506 6320 29520
rect 6240 29454 6254 29506
rect 6306 29454 6320 29506
rect 6240 29440 6320 29454
rect 6400 29506 6480 29520
rect 6400 29454 6414 29506
rect 6466 29454 6480 29506
rect 6400 29440 6480 29454
rect 6560 29506 6640 29520
rect 6560 29454 6574 29506
rect 6626 29454 6640 29506
rect 6560 29440 6640 29454
rect 6720 29506 6800 29520
rect 6720 29454 6734 29506
rect 6786 29454 6800 29506
rect 6720 29440 6800 29454
rect 6880 29506 6960 29520
rect 6880 29454 6894 29506
rect 6946 29454 6960 29506
rect 6880 29440 6960 29454
rect 7040 29506 7120 29520
rect 7040 29454 7054 29506
rect 7106 29454 7120 29506
rect 7040 29440 7120 29454
rect 7200 29506 7280 29520
rect 7200 29454 7214 29506
rect 7266 29454 7280 29506
rect 7200 29440 7280 29454
rect 7360 29506 7440 29520
rect 7360 29454 7374 29506
rect 7426 29454 7440 29506
rect 7360 29440 7440 29454
rect 7520 29506 7600 29520
rect 7520 29454 7534 29506
rect 7586 29454 7600 29506
rect 7520 29440 7600 29454
rect 7680 29506 7760 29520
rect 7680 29454 7694 29506
rect 7746 29454 7760 29506
rect 7680 29440 7760 29454
rect 7840 29506 7920 29520
rect 7840 29454 7854 29506
rect 7906 29454 7920 29506
rect 7840 29440 7920 29454
rect 8000 29506 8080 29520
rect 8000 29454 8014 29506
rect 8066 29454 8080 29506
rect 8000 29440 8080 29454
rect 8160 29506 8240 29520
rect 8160 29454 8174 29506
rect 8226 29454 8240 29506
rect 8160 29440 8240 29454
rect 8320 29506 8400 29520
rect 8320 29454 8334 29506
rect 8386 29454 8400 29506
rect 8320 29440 8400 29454
rect 12480 29506 12560 29520
rect 12480 29454 12494 29506
rect 12546 29454 12560 29506
rect 12480 29440 12560 29454
rect 12640 29506 12720 29520
rect 12640 29454 12654 29506
rect 12706 29454 12720 29506
rect 12640 29440 12720 29454
rect 12800 29506 12880 29520
rect 12800 29454 12814 29506
rect 12866 29454 12880 29506
rect 12800 29440 12880 29454
rect 12960 29506 13040 29520
rect 12960 29454 12974 29506
rect 13026 29454 13040 29506
rect 12960 29440 13040 29454
rect 13120 29506 13200 29520
rect 13120 29454 13134 29506
rect 13186 29454 13200 29506
rect 13120 29440 13200 29454
rect 13280 29506 13360 29520
rect 13280 29454 13294 29506
rect 13346 29454 13360 29506
rect 13280 29440 13360 29454
rect 13440 29506 13520 29520
rect 13440 29454 13454 29506
rect 13506 29454 13520 29506
rect 13440 29440 13520 29454
rect 13600 29506 13680 29520
rect 13600 29454 13614 29506
rect 13666 29454 13680 29506
rect 13600 29440 13680 29454
rect 13760 29506 13840 29520
rect 13760 29454 13774 29506
rect 13826 29454 13840 29506
rect 13760 29440 13840 29454
rect 13920 29506 14000 29520
rect 13920 29454 13934 29506
rect 13986 29454 14000 29506
rect 13920 29440 14000 29454
rect 14080 29506 14160 29520
rect 14080 29454 14094 29506
rect 14146 29454 14160 29506
rect 14080 29440 14160 29454
rect 14240 29506 14320 29520
rect 14240 29454 14254 29506
rect 14306 29454 14320 29506
rect 14240 29440 14320 29454
rect 14400 29506 14480 29520
rect 14400 29454 14414 29506
rect 14466 29454 14480 29506
rect 14400 29440 14480 29454
rect 14560 29506 14640 29520
rect 14560 29454 14574 29506
rect 14626 29454 14640 29506
rect 14560 29440 14640 29454
rect 14720 29506 14800 29520
rect 14720 29454 14734 29506
rect 14786 29454 14800 29506
rect 14720 29440 14800 29454
rect 14880 29506 14960 29520
rect 14880 29454 14894 29506
rect 14946 29454 14960 29506
rect 14880 29440 14960 29454
rect 15040 29506 15120 29520
rect 15040 29454 15054 29506
rect 15106 29454 15120 29506
rect 15040 29440 15120 29454
rect 15200 29506 15280 29520
rect 15200 29454 15214 29506
rect 15266 29454 15280 29506
rect 15200 29440 15280 29454
rect 15360 29506 15440 29520
rect 15360 29454 15374 29506
rect 15426 29454 15440 29506
rect 15360 29440 15440 29454
rect 15520 29506 15600 29520
rect 15520 29454 15534 29506
rect 15586 29454 15600 29506
rect 15520 29440 15600 29454
rect 15680 29506 15760 29520
rect 15680 29454 15694 29506
rect 15746 29454 15760 29506
rect 15680 29440 15760 29454
rect 15840 29506 15920 29520
rect 15840 29454 15854 29506
rect 15906 29454 15920 29506
rect 15840 29440 15920 29454
rect 16000 29506 16080 29520
rect 16000 29454 16014 29506
rect 16066 29454 16080 29506
rect 16000 29440 16080 29454
rect 16160 29506 16240 29520
rect 16160 29454 16174 29506
rect 16226 29454 16240 29506
rect 16160 29440 16240 29454
rect 16320 29506 16400 29520
rect 16320 29454 16334 29506
rect 16386 29454 16400 29506
rect 16320 29440 16400 29454
rect 16480 29506 16560 29520
rect 16480 29454 16494 29506
rect 16546 29454 16560 29506
rect 16480 29440 16560 29454
rect 16640 29506 16720 29520
rect 16640 29454 16654 29506
rect 16706 29454 16720 29506
rect 16640 29440 16720 29454
rect 16800 29506 16880 29520
rect 16800 29454 16814 29506
rect 16866 29454 16880 29506
rect 16800 29440 16880 29454
rect 16960 29506 17040 29520
rect 16960 29454 16974 29506
rect 17026 29454 17040 29506
rect 16960 29440 17040 29454
rect 17120 29506 17200 29520
rect 17120 29454 17134 29506
rect 17186 29454 17200 29506
rect 17120 29440 17200 29454
rect 17280 29506 17360 29520
rect 17280 29454 17294 29506
rect 17346 29454 17360 29506
rect 17280 29440 17360 29454
rect 17440 29506 17520 29520
rect 17440 29454 17454 29506
rect 17506 29454 17520 29506
rect 17440 29440 17520 29454
rect 17600 29506 17680 29520
rect 17600 29454 17614 29506
rect 17666 29454 17680 29506
rect 17600 29440 17680 29454
rect 17760 29506 17840 29520
rect 17760 29454 17774 29506
rect 17826 29454 17840 29506
rect 17760 29440 17840 29454
rect 17920 29506 18000 29520
rect 17920 29454 17934 29506
rect 17986 29454 18000 29506
rect 17920 29440 18000 29454
rect 18080 29506 18160 29520
rect 18080 29454 18094 29506
rect 18146 29454 18160 29506
rect 18080 29440 18160 29454
rect 18240 29506 18320 29520
rect 18240 29454 18254 29506
rect 18306 29454 18320 29506
rect 18240 29440 18320 29454
rect 18400 29506 18480 29520
rect 18400 29454 18414 29506
rect 18466 29454 18480 29506
rect 18400 29440 18480 29454
rect 18560 29506 18640 29520
rect 18560 29454 18574 29506
rect 18626 29454 18640 29506
rect 18560 29440 18640 29454
rect 18720 29506 18800 29520
rect 18720 29454 18734 29506
rect 18786 29454 18800 29506
rect 18720 29440 18800 29454
rect 18880 29506 18960 29520
rect 18880 29454 18894 29506
rect 18946 29454 18960 29506
rect 18880 29440 18960 29454
rect 23120 29506 23200 29520
rect 23120 29454 23134 29506
rect 23186 29454 23200 29506
rect 23120 29440 23200 29454
rect 23280 29506 23360 29520
rect 23280 29454 23294 29506
rect 23346 29454 23360 29506
rect 23280 29440 23360 29454
rect 23440 29506 23520 29520
rect 23440 29454 23454 29506
rect 23506 29454 23520 29506
rect 23440 29440 23520 29454
rect 23600 29506 23680 29520
rect 23600 29454 23614 29506
rect 23666 29454 23680 29506
rect 23600 29440 23680 29454
rect 23760 29506 23840 29520
rect 23760 29454 23774 29506
rect 23826 29454 23840 29506
rect 23760 29440 23840 29454
rect 23920 29506 24000 29520
rect 23920 29454 23934 29506
rect 23986 29454 24000 29506
rect 23920 29440 24000 29454
rect 24080 29506 24160 29520
rect 24080 29454 24094 29506
rect 24146 29454 24160 29506
rect 24080 29440 24160 29454
rect 24240 29506 24320 29520
rect 24240 29454 24254 29506
rect 24306 29454 24320 29506
rect 24240 29440 24320 29454
rect 24400 29506 24480 29520
rect 24400 29454 24414 29506
rect 24466 29454 24480 29506
rect 24400 29440 24480 29454
rect 24560 29506 24640 29520
rect 24560 29454 24574 29506
rect 24626 29454 24640 29506
rect 24560 29440 24640 29454
rect 24720 29506 24800 29520
rect 24720 29454 24734 29506
rect 24786 29454 24800 29506
rect 24720 29440 24800 29454
rect 24880 29506 24960 29520
rect 24880 29454 24894 29506
rect 24946 29454 24960 29506
rect 24880 29440 24960 29454
rect 25040 29506 25120 29520
rect 25040 29454 25054 29506
rect 25106 29454 25120 29506
rect 25040 29440 25120 29454
rect 25200 29506 25280 29520
rect 25200 29454 25214 29506
rect 25266 29454 25280 29506
rect 25200 29440 25280 29454
rect 25360 29506 25440 29520
rect 25360 29454 25374 29506
rect 25426 29454 25440 29506
rect 25360 29440 25440 29454
rect 25520 29506 25600 29520
rect 25520 29454 25534 29506
rect 25586 29454 25600 29506
rect 25520 29440 25600 29454
rect 25680 29506 25760 29520
rect 25680 29454 25694 29506
rect 25746 29454 25760 29506
rect 25680 29440 25760 29454
rect 25840 29506 25920 29520
rect 25840 29454 25854 29506
rect 25906 29454 25920 29506
rect 25840 29440 25920 29454
rect 26000 29506 26080 29520
rect 26000 29454 26014 29506
rect 26066 29454 26080 29506
rect 26000 29440 26080 29454
rect 26160 29506 26240 29520
rect 26160 29454 26174 29506
rect 26226 29454 26240 29506
rect 26160 29440 26240 29454
rect 26320 29506 26400 29520
rect 26320 29454 26334 29506
rect 26386 29454 26400 29506
rect 26320 29440 26400 29454
rect 26480 29506 26560 29520
rect 26480 29454 26494 29506
rect 26546 29454 26560 29506
rect 26480 29440 26560 29454
rect 26640 29506 26720 29520
rect 26640 29454 26654 29506
rect 26706 29454 26720 29506
rect 26640 29440 26720 29454
rect 26800 29506 26880 29520
rect 26800 29454 26814 29506
rect 26866 29454 26880 29506
rect 26800 29440 26880 29454
rect 26960 29506 27040 29520
rect 26960 29454 26974 29506
rect 27026 29454 27040 29506
rect 26960 29440 27040 29454
rect 27120 29506 27200 29520
rect 27120 29454 27134 29506
rect 27186 29454 27200 29506
rect 27120 29440 27200 29454
rect 27280 29506 27360 29520
rect 27280 29454 27294 29506
rect 27346 29454 27360 29506
rect 27280 29440 27360 29454
rect 27440 29506 27520 29520
rect 27440 29454 27454 29506
rect 27506 29454 27520 29506
rect 27440 29440 27520 29454
rect 27600 29506 27680 29520
rect 27600 29454 27614 29506
rect 27666 29454 27680 29506
rect 27600 29440 27680 29454
rect 27760 29506 27840 29520
rect 27760 29454 27774 29506
rect 27826 29454 27840 29506
rect 27760 29440 27840 29454
rect 27920 29506 28000 29520
rect 27920 29454 27934 29506
rect 27986 29454 28000 29506
rect 27920 29440 28000 29454
rect 28080 29506 28160 29520
rect 28080 29454 28094 29506
rect 28146 29454 28160 29506
rect 28080 29440 28160 29454
rect 28240 29506 28320 29520
rect 28240 29454 28254 29506
rect 28306 29454 28320 29506
rect 28240 29440 28320 29454
rect 28400 29506 28480 29520
rect 28400 29454 28414 29506
rect 28466 29454 28480 29506
rect 28400 29440 28480 29454
rect 28560 29506 28640 29520
rect 28560 29454 28574 29506
rect 28626 29454 28640 29506
rect 28560 29440 28640 29454
rect 28720 29506 28800 29520
rect 28720 29454 28734 29506
rect 28786 29454 28800 29506
rect 28720 29440 28800 29454
rect 28880 29506 28960 29520
rect 28880 29454 28894 29506
rect 28946 29454 28960 29506
rect 28880 29440 28960 29454
rect 29040 29506 29120 29520
rect 29040 29454 29054 29506
rect 29106 29454 29120 29506
rect 29040 29440 29120 29454
rect 29200 29506 29280 29520
rect 29200 29454 29214 29506
rect 29266 29454 29280 29506
rect 29200 29440 29280 29454
rect 29360 29506 29440 29520
rect 29360 29454 29374 29506
rect 29426 29454 29440 29506
rect 29360 29440 29440 29454
rect 33520 29506 33600 29520
rect 33520 29454 33534 29506
rect 33586 29454 33600 29506
rect 33520 29440 33600 29454
rect 33680 29506 33760 29520
rect 33680 29454 33694 29506
rect 33746 29454 33760 29506
rect 33680 29440 33760 29454
rect 33840 29506 33920 29520
rect 33840 29454 33854 29506
rect 33906 29454 33920 29506
rect 33840 29440 33920 29454
rect 34000 29506 34080 29520
rect 34000 29454 34014 29506
rect 34066 29454 34080 29506
rect 34000 29440 34080 29454
rect 34160 29506 34240 29520
rect 34160 29454 34174 29506
rect 34226 29454 34240 29506
rect 34160 29440 34240 29454
rect 34320 29506 34400 29520
rect 34320 29454 34334 29506
rect 34386 29454 34400 29506
rect 34320 29440 34400 29454
rect 34480 29506 34560 29520
rect 34480 29454 34494 29506
rect 34546 29454 34560 29506
rect 34480 29440 34560 29454
rect 34640 29506 34720 29520
rect 34640 29454 34654 29506
rect 34706 29454 34720 29506
rect 34640 29440 34720 29454
rect 34800 29506 34880 29520
rect 34800 29454 34814 29506
rect 34866 29454 34880 29506
rect 34800 29440 34880 29454
rect 34960 29506 35040 29520
rect 34960 29454 34974 29506
rect 35026 29454 35040 29506
rect 34960 29440 35040 29454
rect 35120 29506 35200 29520
rect 35120 29454 35134 29506
rect 35186 29454 35200 29506
rect 35120 29440 35200 29454
rect 35280 29506 35360 29520
rect 35280 29454 35294 29506
rect 35346 29454 35360 29506
rect 35280 29440 35360 29454
rect 35440 29506 35520 29520
rect 35440 29454 35454 29506
rect 35506 29454 35520 29506
rect 35440 29440 35520 29454
rect 35600 29506 35680 29520
rect 35600 29454 35614 29506
rect 35666 29454 35680 29506
rect 35600 29440 35680 29454
rect 35760 29506 35840 29520
rect 35760 29454 35774 29506
rect 35826 29454 35840 29506
rect 35760 29440 35840 29454
rect 35920 29506 36000 29520
rect 35920 29454 35934 29506
rect 35986 29454 36000 29506
rect 35920 29440 36000 29454
rect 36080 29506 36160 29520
rect 36080 29454 36094 29506
rect 36146 29454 36160 29506
rect 36080 29440 36160 29454
rect 36240 29506 36320 29520
rect 36240 29454 36254 29506
rect 36306 29454 36320 29506
rect 36240 29440 36320 29454
rect 36400 29506 36480 29520
rect 36400 29454 36414 29506
rect 36466 29454 36480 29506
rect 36400 29440 36480 29454
rect 36560 29506 36640 29520
rect 36560 29454 36574 29506
rect 36626 29454 36640 29506
rect 36560 29440 36640 29454
rect 36720 29506 36800 29520
rect 36720 29454 36734 29506
rect 36786 29454 36800 29506
rect 36720 29440 36800 29454
rect 36880 29506 36960 29520
rect 36880 29454 36894 29506
rect 36946 29454 36960 29506
rect 36880 29440 36960 29454
rect 37040 29506 37120 29520
rect 37040 29454 37054 29506
rect 37106 29454 37120 29506
rect 37040 29440 37120 29454
rect 37200 29506 37280 29520
rect 37200 29454 37214 29506
rect 37266 29454 37280 29506
rect 37200 29440 37280 29454
rect 37360 29506 37440 29520
rect 37360 29454 37374 29506
rect 37426 29454 37440 29506
rect 37360 29440 37440 29454
rect 37520 29506 37600 29520
rect 37520 29454 37534 29506
rect 37586 29454 37600 29506
rect 37520 29440 37600 29454
rect 37680 29506 37760 29520
rect 37680 29454 37694 29506
rect 37746 29454 37760 29506
rect 37680 29440 37760 29454
rect 37840 29506 37920 29520
rect 37840 29454 37854 29506
rect 37906 29454 37920 29506
rect 37840 29440 37920 29454
rect 38000 29506 38080 29520
rect 38000 29454 38014 29506
rect 38066 29454 38080 29506
rect 38000 29440 38080 29454
rect 38160 29506 38240 29520
rect 38160 29454 38174 29506
rect 38226 29454 38240 29506
rect 38160 29440 38240 29454
rect 38320 29506 38400 29520
rect 38320 29454 38334 29506
rect 38386 29454 38400 29506
rect 38320 29440 38400 29454
rect 38480 29506 38560 29520
rect 38480 29454 38494 29506
rect 38546 29454 38560 29506
rect 38480 29440 38560 29454
rect 38640 29506 38720 29520
rect 38640 29454 38654 29506
rect 38706 29454 38720 29506
rect 38640 29440 38720 29454
rect 38800 29506 38880 29520
rect 38800 29454 38814 29506
rect 38866 29454 38880 29506
rect 38800 29440 38880 29454
rect 38960 29506 39040 29520
rect 38960 29454 38974 29506
rect 39026 29454 39040 29506
rect 38960 29440 39040 29454
rect 39120 29506 39200 29520
rect 39120 29454 39134 29506
rect 39186 29454 39200 29506
rect 39120 29440 39200 29454
rect 39280 29506 39360 29520
rect 39280 29454 39294 29506
rect 39346 29454 39360 29506
rect 39280 29440 39360 29454
rect 39440 29506 39520 29520
rect 39440 29454 39454 29506
rect 39506 29454 39520 29506
rect 39440 29440 39520 29454
rect 39600 29506 39680 29520
rect 39600 29454 39614 29506
rect 39666 29454 39680 29506
rect 39600 29440 39680 29454
rect 39760 29506 39840 29520
rect 39760 29454 39774 29506
rect 39826 29454 39840 29506
rect 39760 29440 39840 29454
rect 39920 29506 40000 29520
rect 39920 29454 39934 29506
rect 39986 29454 40000 29506
rect 39920 29440 40000 29454
rect 40080 29506 40160 29520
rect 40080 29454 40094 29506
rect 40146 29454 40160 29506
rect 40080 29440 40160 29454
rect 40240 29506 40320 29520
rect 40240 29454 40254 29506
rect 40306 29454 40320 29506
rect 40240 29440 40320 29454
rect 40400 29506 40480 29520
rect 40400 29454 40414 29506
rect 40466 29454 40480 29506
rect 40400 29440 40480 29454
rect 40560 29506 40640 29520
rect 40560 29454 40574 29506
rect 40626 29454 40640 29506
rect 40560 29440 40640 29454
rect 40720 29506 40800 29520
rect 40720 29454 40734 29506
rect 40786 29454 40800 29506
rect 40720 29440 40800 29454
rect 40880 29506 40960 29520
rect 40880 29454 40894 29506
rect 40946 29454 40960 29506
rect 40880 29440 40960 29454
rect 41040 29506 41120 29520
rect 41040 29454 41054 29506
rect 41106 29454 41120 29506
rect 41040 29440 41120 29454
rect 41200 29506 41280 29520
rect 41200 29454 41214 29506
rect 41266 29454 41280 29506
rect 41200 29440 41280 29454
rect 41360 29506 41440 29520
rect 41360 29454 41374 29506
rect 41426 29454 41440 29506
rect 41360 29440 41440 29454
rect 41520 29506 41600 29520
rect 41520 29454 41534 29506
rect 41586 29454 41600 29506
rect 41520 29440 41600 29454
rect 41680 29506 41760 29520
rect 41680 29454 41694 29506
rect 41746 29454 41760 29506
rect 41680 29440 41760 29454
rect 41840 29506 41920 29520
rect 41840 29454 41854 29506
rect 41906 29454 41920 29506
rect 41840 29440 41920 29454
<< via1 >>
rect 14 37337 66 37346
rect 14 37303 23 37337
rect 23 37303 57 37337
rect 57 37303 66 37337
rect 14 37294 66 37303
rect 174 37337 226 37346
rect 174 37303 183 37337
rect 183 37303 217 37337
rect 217 37303 226 37337
rect 174 37294 226 37303
rect 334 37337 386 37346
rect 334 37303 343 37337
rect 343 37303 377 37337
rect 377 37303 386 37337
rect 334 37294 386 37303
rect 494 37337 546 37346
rect 494 37303 503 37337
rect 503 37303 537 37337
rect 537 37303 546 37337
rect 494 37294 546 37303
rect 654 37337 706 37346
rect 654 37303 663 37337
rect 663 37303 697 37337
rect 697 37303 706 37337
rect 654 37294 706 37303
rect 814 37337 866 37346
rect 814 37303 823 37337
rect 823 37303 857 37337
rect 857 37303 866 37337
rect 814 37294 866 37303
rect 974 37337 1026 37346
rect 974 37303 983 37337
rect 983 37303 1017 37337
rect 1017 37303 1026 37337
rect 974 37294 1026 37303
rect 1134 37337 1186 37346
rect 1134 37303 1143 37337
rect 1143 37303 1177 37337
rect 1177 37303 1186 37337
rect 1134 37294 1186 37303
rect 1294 37337 1346 37346
rect 1294 37303 1303 37337
rect 1303 37303 1337 37337
rect 1337 37303 1346 37337
rect 1294 37294 1346 37303
rect 1454 37337 1506 37346
rect 1454 37303 1463 37337
rect 1463 37303 1497 37337
rect 1497 37303 1506 37337
rect 1454 37294 1506 37303
rect 1614 37337 1666 37346
rect 1614 37303 1623 37337
rect 1623 37303 1657 37337
rect 1657 37303 1666 37337
rect 1614 37294 1666 37303
rect 1774 37337 1826 37346
rect 1774 37303 1783 37337
rect 1783 37303 1817 37337
rect 1817 37303 1826 37337
rect 1774 37294 1826 37303
rect 1934 37337 1986 37346
rect 1934 37303 1943 37337
rect 1943 37303 1977 37337
rect 1977 37303 1986 37337
rect 1934 37294 1986 37303
rect 2094 37337 2146 37346
rect 2094 37303 2103 37337
rect 2103 37303 2137 37337
rect 2137 37303 2146 37337
rect 2094 37294 2146 37303
rect 2254 37337 2306 37346
rect 2254 37303 2263 37337
rect 2263 37303 2297 37337
rect 2297 37303 2306 37337
rect 2254 37294 2306 37303
rect 2414 37337 2466 37346
rect 2414 37303 2423 37337
rect 2423 37303 2457 37337
rect 2457 37303 2466 37337
rect 2414 37294 2466 37303
rect 2574 37337 2626 37346
rect 2574 37303 2583 37337
rect 2583 37303 2617 37337
rect 2617 37303 2626 37337
rect 2574 37294 2626 37303
rect 2734 37337 2786 37346
rect 2734 37303 2743 37337
rect 2743 37303 2777 37337
rect 2777 37303 2786 37337
rect 2734 37294 2786 37303
rect 2894 37337 2946 37346
rect 2894 37303 2903 37337
rect 2903 37303 2937 37337
rect 2937 37303 2946 37337
rect 2894 37294 2946 37303
rect 3054 37337 3106 37346
rect 3054 37303 3063 37337
rect 3063 37303 3097 37337
rect 3097 37303 3106 37337
rect 3054 37294 3106 37303
rect 3214 37337 3266 37346
rect 3214 37303 3223 37337
rect 3223 37303 3257 37337
rect 3257 37303 3266 37337
rect 3214 37294 3266 37303
rect 3374 37337 3426 37346
rect 3374 37303 3383 37337
rect 3383 37303 3417 37337
rect 3417 37303 3426 37337
rect 3374 37294 3426 37303
rect 3534 37337 3586 37346
rect 3534 37303 3543 37337
rect 3543 37303 3577 37337
rect 3577 37303 3586 37337
rect 3534 37294 3586 37303
rect 3694 37337 3746 37346
rect 3694 37303 3703 37337
rect 3703 37303 3737 37337
rect 3737 37303 3746 37337
rect 3694 37294 3746 37303
rect 3854 37337 3906 37346
rect 3854 37303 3863 37337
rect 3863 37303 3897 37337
rect 3897 37303 3906 37337
rect 3854 37294 3906 37303
rect 4014 37337 4066 37346
rect 4014 37303 4023 37337
rect 4023 37303 4057 37337
rect 4057 37303 4066 37337
rect 4014 37294 4066 37303
rect 4174 37337 4226 37346
rect 4174 37303 4183 37337
rect 4183 37303 4217 37337
rect 4217 37303 4226 37337
rect 4174 37294 4226 37303
rect 4334 37337 4386 37346
rect 4334 37303 4343 37337
rect 4343 37303 4377 37337
rect 4377 37303 4386 37337
rect 4334 37294 4386 37303
rect 4494 37337 4546 37346
rect 4494 37303 4503 37337
rect 4503 37303 4537 37337
rect 4537 37303 4546 37337
rect 4494 37294 4546 37303
rect 4654 37337 4706 37346
rect 4654 37303 4663 37337
rect 4663 37303 4697 37337
rect 4697 37303 4706 37337
rect 4654 37294 4706 37303
rect 4814 37337 4866 37346
rect 4814 37303 4823 37337
rect 4823 37303 4857 37337
rect 4857 37303 4866 37337
rect 4814 37294 4866 37303
rect 4974 37337 5026 37346
rect 4974 37303 4983 37337
rect 4983 37303 5017 37337
rect 5017 37303 5026 37337
rect 4974 37294 5026 37303
rect 5134 37337 5186 37346
rect 5134 37303 5143 37337
rect 5143 37303 5177 37337
rect 5177 37303 5186 37337
rect 5134 37294 5186 37303
rect 5294 37337 5346 37346
rect 5294 37303 5303 37337
rect 5303 37303 5337 37337
rect 5337 37303 5346 37337
rect 5294 37294 5346 37303
rect 5454 37337 5506 37346
rect 5454 37303 5463 37337
rect 5463 37303 5497 37337
rect 5497 37303 5506 37337
rect 5454 37294 5506 37303
rect 5614 37337 5666 37346
rect 5614 37303 5623 37337
rect 5623 37303 5657 37337
rect 5657 37303 5666 37337
rect 5614 37294 5666 37303
rect 5774 37337 5826 37346
rect 5774 37303 5783 37337
rect 5783 37303 5817 37337
rect 5817 37303 5826 37337
rect 5774 37294 5826 37303
rect 5934 37337 5986 37346
rect 5934 37303 5943 37337
rect 5943 37303 5977 37337
rect 5977 37303 5986 37337
rect 5934 37294 5986 37303
rect 6094 37337 6146 37346
rect 6094 37303 6103 37337
rect 6103 37303 6137 37337
rect 6137 37303 6146 37337
rect 6094 37294 6146 37303
rect 6254 37337 6306 37346
rect 6254 37303 6263 37337
rect 6263 37303 6297 37337
rect 6297 37303 6306 37337
rect 6254 37294 6306 37303
rect 6414 37337 6466 37346
rect 6414 37303 6423 37337
rect 6423 37303 6457 37337
rect 6457 37303 6466 37337
rect 6414 37294 6466 37303
rect 6574 37337 6626 37346
rect 6574 37303 6583 37337
rect 6583 37303 6617 37337
rect 6617 37303 6626 37337
rect 6574 37294 6626 37303
rect 6734 37337 6786 37346
rect 6734 37303 6743 37337
rect 6743 37303 6777 37337
rect 6777 37303 6786 37337
rect 6734 37294 6786 37303
rect 6894 37337 6946 37346
rect 6894 37303 6903 37337
rect 6903 37303 6937 37337
rect 6937 37303 6946 37337
rect 6894 37294 6946 37303
rect 7054 37337 7106 37346
rect 7054 37303 7063 37337
rect 7063 37303 7097 37337
rect 7097 37303 7106 37337
rect 7054 37294 7106 37303
rect 7214 37337 7266 37346
rect 7214 37303 7223 37337
rect 7223 37303 7257 37337
rect 7257 37303 7266 37337
rect 7214 37294 7266 37303
rect 7374 37337 7426 37346
rect 7374 37303 7383 37337
rect 7383 37303 7417 37337
rect 7417 37303 7426 37337
rect 7374 37294 7426 37303
rect 7534 37337 7586 37346
rect 7534 37303 7543 37337
rect 7543 37303 7577 37337
rect 7577 37303 7586 37337
rect 7534 37294 7586 37303
rect 7694 37337 7746 37346
rect 7694 37303 7703 37337
rect 7703 37303 7737 37337
rect 7737 37303 7746 37337
rect 7694 37294 7746 37303
rect 7854 37337 7906 37346
rect 7854 37303 7863 37337
rect 7863 37303 7897 37337
rect 7897 37303 7906 37337
rect 7854 37294 7906 37303
rect 8014 37337 8066 37346
rect 8014 37303 8023 37337
rect 8023 37303 8057 37337
rect 8057 37303 8066 37337
rect 8014 37294 8066 37303
rect 8174 37337 8226 37346
rect 8174 37303 8183 37337
rect 8183 37303 8217 37337
rect 8217 37303 8226 37337
rect 8174 37294 8226 37303
rect 8334 37337 8386 37346
rect 8334 37303 8343 37337
rect 8343 37303 8377 37337
rect 8377 37303 8386 37337
rect 8334 37294 8386 37303
rect 12494 37337 12546 37346
rect 12494 37303 12503 37337
rect 12503 37303 12537 37337
rect 12537 37303 12546 37337
rect 12494 37294 12546 37303
rect 12654 37337 12706 37346
rect 12654 37303 12663 37337
rect 12663 37303 12697 37337
rect 12697 37303 12706 37337
rect 12654 37294 12706 37303
rect 12814 37337 12866 37346
rect 12814 37303 12823 37337
rect 12823 37303 12857 37337
rect 12857 37303 12866 37337
rect 12814 37294 12866 37303
rect 12974 37337 13026 37346
rect 12974 37303 12983 37337
rect 12983 37303 13017 37337
rect 13017 37303 13026 37337
rect 12974 37294 13026 37303
rect 13134 37337 13186 37346
rect 13134 37303 13143 37337
rect 13143 37303 13177 37337
rect 13177 37303 13186 37337
rect 13134 37294 13186 37303
rect 13294 37337 13346 37346
rect 13294 37303 13303 37337
rect 13303 37303 13337 37337
rect 13337 37303 13346 37337
rect 13294 37294 13346 37303
rect 13454 37337 13506 37346
rect 13454 37303 13463 37337
rect 13463 37303 13497 37337
rect 13497 37303 13506 37337
rect 13454 37294 13506 37303
rect 13614 37337 13666 37346
rect 13614 37303 13623 37337
rect 13623 37303 13657 37337
rect 13657 37303 13666 37337
rect 13614 37294 13666 37303
rect 13774 37337 13826 37346
rect 13774 37303 13783 37337
rect 13783 37303 13817 37337
rect 13817 37303 13826 37337
rect 13774 37294 13826 37303
rect 13934 37337 13986 37346
rect 13934 37303 13943 37337
rect 13943 37303 13977 37337
rect 13977 37303 13986 37337
rect 13934 37294 13986 37303
rect 14094 37337 14146 37346
rect 14094 37303 14103 37337
rect 14103 37303 14137 37337
rect 14137 37303 14146 37337
rect 14094 37294 14146 37303
rect 14254 37337 14306 37346
rect 14254 37303 14263 37337
rect 14263 37303 14297 37337
rect 14297 37303 14306 37337
rect 14254 37294 14306 37303
rect 14414 37337 14466 37346
rect 14414 37303 14423 37337
rect 14423 37303 14457 37337
rect 14457 37303 14466 37337
rect 14414 37294 14466 37303
rect 14574 37337 14626 37346
rect 14574 37303 14583 37337
rect 14583 37303 14617 37337
rect 14617 37303 14626 37337
rect 14574 37294 14626 37303
rect 14734 37337 14786 37346
rect 14734 37303 14743 37337
rect 14743 37303 14777 37337
rect 14777 37303 14786 37337
rect 14734 37294 14786 37303
rect 14894 37337 14946 37346
rect 14894 37303 14903 37337
rect 14903 37303 14937 37337
rect 14937 37303 14946 37337
rect 14894 37294 14946 37303
rect 15054 37337 15106 37346
rect 15054 37303 15063 37337
rect 15063 37303 15097 37337
rect 15097 37303 15106 37337
rect 15054 37294 15106 37303
rect 15214 37337 15266 37346
rect 15214 37303 15223 37337
rect 15223 37303 15257 37337
rect 15257 37303 15266 37337
rect 15214 37294 15266 37303
rect 15374 37337 15426 37346
rect 15374 37303 15383 37337
rect 15383 37303 15417 37337
rect 15417 37303 15426 37337
rect 15374 37294 15426 37303
rect 15534 37337 15586 37346
rect 15534 37303 15543 37337
rect 15543 37303 15577 37337
rect 15577 37303 15586 37337
rect 15534 37294 15586 37303
rect 15694 37337 15746 37346
rect 15694 37303 15703 37337
rect 15703 37303 15737 37337
rect 15737 37303 15746 37337
rect 15694 37294 15746 37303
rect 15854 37337 15906 37346
rect 15854 37303 15863 37337
rect 15863 37303 15897 37337
rect 15897 37303 15906 37337
rect 15854 37294 15906 37303
rect 16014 37337 16066 37346
rect 16014 37303 16023 37337
rect 16023 37303 16057 37337
rect 16057 37303 16066 37337
rect 16014 37294 16066 37303
rect 16174 37337 16226 37346
rect 16174 37303 16183 37337
rect 16183 37303 16217 37337
rect 16217 37303 16226 37337
rect 16174 37294 16226 37303
rect 16334 37337 16386 37346
rect 16334 37303 16343 37337
rect 16343 37303 16377 37337
rect 16377 37303 16386 37337
rect 16334 37294 16386 37303
rect 16494 37337 16546 37346
rect 16494 37303 16503 37337
rect 16503 37303 16537 37337
rect 16537 37303 16546 37337
rect 16494 37294 16546 37303
rect 16654 37337 16706 37346
rect 16654 37303 16663 37337
rect 16663 37303 16697 37337
rect 16697 37303 16706 37337
rect 16654 37294 16706 37303
rect 16814 37337 16866 37346
rect 16814 37303 16823 37337
rect 16823 37303 16857 37337
rect 16857 37303 16866 37337
rect 16814 37294 16866 37303
rect 16974 37337 17026 37346
rect 16974 37303 16983 37337
rect 16983 37303 17017 37337
rect 17017 37303 17026 37337
rect 16974 37294 17026 37303
rect 17134 37337 17186 37346
rect 17134 37303 17143 37337
rect 17143 37303 17177 37337
rect 17177 37303 17186 37337
rect 17134 37294 17186 37303
rect 17294 37337 17346 37346
rect 17294 37303 17303 37337
rect 17303 37303 17337 37337
rect 17337 37303 17346 37337
rect 17294 37294 17346 37303
rect 17454 37337 17506 37346
rect 17454 37303 17463 37337
rect 17463 37303 17497 37337
rect 17497 37303 17506 37337
rect 17454 37294 17506 37303
rect 17614 37337 17666 37346
rect 17614 37303 17623 37337
rect 17623 37303 17657 37337
rect 17657 37303 17666 37337
rect 17614 37294 17666 37303
rect 17774 37337 17826 37346
rect 17774 37303 17783 37337
rect 17783 37303 17817 37337
rect 17817 37303 17826 37337
rect 17774 37294 17826 37303
rect 17934 37337 17986 37346
rect 17934 37303 17943 37337
rect 17943 37303 17977 37337
rect 17977 37303 17986 37337
rect 17934 37294 17986 37303
rect 18094 37337 18146 37346
rect 18094 37303 18103 37337
rect 18103 37303 18137 37337
rect 18137 37303 18146 37337
rect 18094 37294 18146 37303
rect 18254 37337 18306 37346
rect 18254 37303 18263 37337
rect 18263 37303 18297 37337
rect 18297 37303 18306 37337
rect 18254 37294 18306 37303
rect 18414 37337 18466 37346
rect 18414 37303 18423 37337
rect 18423 37303 18457 37337
rect 18457 37303 18466 37337
rect 18414 37294 18466 37303
rect 18574 37337 18626 37346
rect 18574 37303 18583 37337
rect 18583 37303 18617 37337
rect 18617 37303 18626 37337
rect 18574 37294 18626 37303
rect 18734 37337 18786 37346
rect 18734 37303 18743 37337
rect 18743 37303 18777 37337
rect 18777 37303 18786 37337
rect 18734 37294 18786 37303
rect 18894 37337 18946 37346
rect 18894 37303 18903 37337
rect 18903 37303 18937 37337
rect 18937 37303 18946 37337
rect 18894 37294 18946 37303
rect 23134 37337 23186 37346
rect 23134 37303 23143 37337
rect 23143 37303 23177 37337
rect 23177 37303 23186 37337
rect 23134 37294 23186 37303
rect 23294 37337 23346 37346
rect 23294 37303 23303 37337
rect 23303 37303 23337 37337
rect 23337 37303 23346 37337
rect 23294 37294 23346 37303
rect 23454 37337 23506 37346
rect 23454 37303 23463 37337
rect 23463 37303 23497 37337
rect 23497 37303 23506 37337
rect 23454 37294 23506 37303
rect 23614 37337 23666 37346
rect 23614 37303 23623 37337
rect 23623 37303 23657 37337
rect 23657 37303 23666 37337
rect 23614 37294 23666 37303
rect 23774 37337 23826 37346
rect 23774 37303 23783 37337
rect 23783 37303 23817 37337
rect 23817 37303 23826 37337
rect 23774 37294 23826 37303
rect 23934 37337 23986 37346
rect 23934 37303 23943 37337
rect 23943 37303 23977 37337
rect 23977 37303 23986 37337
rect 23934 37294 23986 37303
rect 24094 37337 24146 37346
rect 24094 37303 24103 37337
rect 24103 37303 24137 37337
rect 24137 37303 24146 37337
rect 24094 37294 24146 37303
rect 24254 37337 24306 37346
rect 24254 37303 24263 37337
rect 24263 37303 24297 37337
rect 24297 37303 24306 37337
rect 24254 37294 24306 37303
rect 24414 37337 24466 37346
rect 24414 37303 24423 37337
rect 24423 37303 24457 37337
rect 24457 37303 24466 37337
rect 24414 37294 24466 37303
rect 24574 37337 24626 37346
rect 24574 37303 24583 37337
rect 24583 37303 24617 37337
rect 24617 37303 24626 37337
rect 24574 37294 24626 37303
rect 24734 37337 24786 37346
rect 24734 37303 24743 37337
rect 24743 37303 24777 37337
rect 24777 37303 24786 37337
rect 24734 37294 24786 37303
rect 24894 37337 24946 37346
rect 24894 37303 24903 37337
rect 24903 37303 24937 37337
rect 24937 37303 24946 37337
rect 24894 37294 24946 37303
rect 25054 37337 25106 37346
rect 25054 37303 25063 37337
rect 25063 37303 25097 37337
rect 25097 37303 25106 37337
rect 25054 37294 25106 37303
rect 25214 37337 25266 37346
rect 25214 37303 25223 37337
rect 25223 37303 25257 37337
rect 25257 37303 25266 37337
rect 25214 37294 25266 37303
rect 25374 37337 25426 37346
rect 25374 37303 25383 37337
rect 25383 37303 25417 37337
rect 25417 37303 25426 37337
rect 25374 37294 25426 37303
rect 25534 37337 25586 37346
rect 25534 37303 25543 37337
rect 25543 37303 25577 37337
rect 25577 37303 25586 37337
rect 25534 37294 25586 37303
rect 25694 37337 25746 37346
rect 25694 37303 25703 37337
rect 25703 37303 25737 37337
rect 25737 37303 25746 37337
rect 25694 37294 25746 37303
rect 25854 37337 25906 37346
rect 25854 37303 25863 37337
rect 25863 37303 25897 37337
rect 25897 37303 25906 37337
rect 25854 37294 25906 37303
rect 26014 37337 26066 37346
rect 26014 37303 26023 37337
rect 26023 37303 26057 37337
rect 26057 37303 26066 37337
rect 26014 37294 26066 37303
rect 26174 37337 26226 37346
rect 26174 37303 26183 37337
rect 26183 37303 26217 37337
rect 26217 37303 26226 37337
rect 26174 37294 26226 37303
rect 26334 37337 26386 37346
rect 26334 37303 26343 37337
rect 26343 37303 26377 37337
rect 26377 37303 26386 37337
rect 26334 37294 26386 37303
rect 26494 37337 26546 37346
rect 26494 37303 26503 37337
rect 26503 37303 26537 37337
rect 26537 37303 26546 37337
rect 26494 37294 26546 37303
rect 26654 37337 26706 37346
rect 26654 37303 26663 37337
rect 26663 37303 26697 37337
rect 26697 37303 26706 37337
rect 26654 37294 26706 37303
rect 26814 37337 26866 37346
rect 26814 37303 26823 37337
rect 26823 37303 26857 37337
rect 26857 37303 26866 37337
rect 26814 37294 26866 37303
rect 26974 37337 27026 37346
rect 26974 37303 26983 37337
rect 26983 37303 27017 37337
rect 27017 37303 27026 37337
rect 26974 37294 27026 37303
rect 27134 37337 27186 37346
rect 27134 37303 27143 37337
rect 27143 37303 27177 37337
rect 27177 37303 27186 37337
rect 27134 37294 27186 37303
rect 27294 37337 27346 37346
rect 27294 37303 27303 37337
rect 27303 37303 27337 37337
rect 27337 37303 27346 37337
rect 27294 37294 27346 37303
rect 27454 37337 27506 37346
rect 27454 37303 27463 37337
rect 27463 37303 27497 37337
rect 27497 37303 27506 37337
rect 27454 37294 27506 37303
rect 27614 37337 27666 37346
rect 27614 37303 27623 37337
rect 27623 37303 27657 37337
rect 27657 37303 27666 37337
rect 27614 37294 27666 37303
rect 27774 37337 27826 37346
rect 27774 37303 27783 37337
rect 27783 37303 27817 37337
rect 27817 37303 27826 37337
rect 27774 37294 27826 37303
rect 27934 37337 27986 37346
rect 27934 37303 27943 37337
rect 27943 37303 27977 37337
rect 27977 37303 27986 37337
rect 27934 37294 27986 37303
rect 28094 37337 28146 37346
rect 28094 37303 28103 37337
rect 28103 37303 28137 37337
rect 28137 37303 28146 37337
rect 28094 37294 28146 37303
rect 28254 37337 28306 37346
rect 28254 37303 28263 37337
rect 28263 37303 28297 37337
rect 28297 37303 28306 37337
rect 28254 37294 28306 37303
rect 28414 37337 28466 37346
rect 28414 37303 28423 37337
rect 28423 37303 28457 37337
rect 28457 37303 28466 37337
rect 28414 37294 28466 37303
rect 28574 37337 28626 37346
rect 28574 37303 28583 37337
rect 28583 37303 28617 37337
rect 28617 37303 28626 37337
rect 28574 37294 28626 37303
rect 28734 37337 28786 37346
rect 28734 37303 28743 37337
rect 28743 37303 28777 37337
rect 28777 37303 28786 37337
rect 28734 37294 28786 37303
rect 28894 37337 28946 37346
rect 28894 37303 28903 37337
rect 28903 37303 28937 37337
rect 28937 37303 28946 37337
rect 28894 37294 28946 37303
rect 29054 37337 29106 37346
rect 29054 37303 29063 37337
rect 29063 37303 29097 37337
rect 29097 37303 29106 37337
rect 29054 37294 29106 37303
rect 29214 37337 29266 37346
rect 29214 37303 29223 37337
rect 29223 37303 29257 37337
rect 29257 37303 29266 37337
rect 29214 37294 29266 37303
rect 29374 37337 29426 37346
rect 29374 37303 29383 37337
rect 29383 37303 29417 37337
rect 29417 37303 29426 37337
rect 29374 37294 29426 37303
rect 33534 37337 33586 37346
rect 33534 37303 33543 37337
rect 33543 37303 33577 37337
rect 33577 37303 33586 37337
rect 33534 37294 33586 37303
rect 33694 37337 33746 37346
rect 33694 37303 33703 37337
rect 33703 37303 33737 37337
rect 33737 37303 33746 37337
rect 33694 37294 33746 37303
rect 33854 37337 33906 37346
rect 33854 37303 33863 37337
rect 33863 37303 33897 37337
rect 33897 37303 33906 37337
rect 33854 37294 33906 37303
rect 34014 37337 34066 37346
rect 34014 37303 34023 37337
rect 34023 37303 34057 37337
rect 34057 37303 34066 37337
rect 34014 37294 34066 37303
rect 34174 37337 34226 37346
rect 34174 37303 34183 37337
rect 34183 37303 34217 37337
rect 34217 37303 34226 37337
rect 34174 37294 34226 37303
rect 34334 37337 34386 37346
rect 34334 37303 34343 37337
rect 34343 37303 34377 37337
rect 34377 37303 34386 37337
rect 34334 37294 34386 37303
rect 34494 37337 34546 37346
rect 34494 37303 34503 37337
rect 34503 37303 34537 37337
rect 34537 37303 34546 37337
rect 34494 37294 34546 37303
rect 34654 37337 34706 37346
rect 34654 37303 34663 37337
rect 34663 37303 34697 37337
rect 34697 37303 34706 37337
rect 34654 37294 34706 37303
rect 34814 37337 34866 37346
rect 34814 37303 34823 37337
rect 34823 37303 34857 37337
rect 34857 37303 34866 37337
rect 34814 37294 34866 37303
rect 34974 37337 35026 37346
rect 34974 37303 34983 37337
rect 34983 37303 35017 37337
rect 35017 37303 35026 37337
rect 34974 37294 35026 37303
rect 35134 37337 35186 37346
rect 35134 37303 35143 37337
rect 35143 37303 35177 37337
rect 35177 37303 35186 37337
rect 35134 37294 35186 37303
rect 35294 37337 35346 37346
rect 35294 37303 35303 37337
rect 35303 37303 35337 37337
rect 35337 37303 35346 37337
rect 35294 37294 35346 37303
rect 35454 37337 35506 37346
rect 35454 37303 35463 37337
rect 35463 37303 35497 37337
rect 35497 37303 35506 37337
rect 35454 37294 35506 37303
rect 35614 37337 35666 37346
rect 35614 37303 35623 37337
rect 35623 37303 35657 37337
rect 35657 37303 35666 37337
rect 35614 37294 35666 37303
rect 35774 37337 35826 37346
rect 35774 37303 35783 37337
rect 35783 37303 35817 37337
rect 35817 37303 35826 37337
rect 35774 37294 35826 37303
rect 35934 37337 35986 37346
rect 35934 37303 35943 37337
rect 35943 37303 35977 37337
rect 35977 37303 35986 37337
rect 35934 37294 35986 37303
rect 36094 37337 36146 37346
rect 36094 37303 36103 37337
rect 36103 37303 36137 37337
rect 36137 37303 36146 37337
rect 36094 37294 36146 37303
rect 36254 37337 36306 37346
rect 36254 37303 36263 37337
rect 36263 37303 36297 37337
rect 36297 37303 36306 37337
rect 36254 37294 36306 37303
rect 36414 37337 36466 37346
rect 36414 37303 36423 37337
rect 36423 37303 36457 37337
rect 36457 37303 36466 37337
rect 36414 37294 36466 37303
rect 36574 37337 36626 37346
rect 36574 37303 36583 37337
rect 36583 37303 36617 37337
rect 36617 37303 36626 37337
rect 36574 37294 36626 37303
rect 36734 37337 36786 37346
rect 36734 37303 36743 37337
rect 36743 37303 36777 37337
rect 36777 37303 36786 37337
rect 36734 37294 36786 37303
rect 36894 37337 36946 37346
rect 36894 37303 36903 37337
rect 36903 37303 36937 37337
rect 36937 37303 36946 37337
rect 36894 37294 36946 37303
rect 37054 37337 37106 37346
rect 37054 37303 37063 37337
rect 37063 37303 37097 37337
rect 37097 37303 37106 37337
rect 37054 37294 37106 37303
rect 37214 37337 37266 37346
rect 37214 37303 37223 37337
rect 37223 37303 37257 37337
rect 37257 37303 37266 37337
rect 37214 37294 37266 37303
rect 37374 37337 37426 37346
rect 37374 37303 37383 37337
rect 37383 37303 37417 37337
rect 37417 37303 37426 37337
rect 37374 37294 37426 37303
rect 37534 37337 37586 37346
rect 37534 37303 37543 37337
rect 37543 37303 37577 37337
rect 37577 37303 37586 37337
rect 37534 37294 37586 37303
rect 37694 37337 37746 37346
rect 37694 37303 37703 37337
rect 37703 37303 37737 37337
rect 37737 37303 37746 37337
rect 37694 37294 37746 37303
rect 37854 37337 37906 37346
rect 37854 37303 37863 37337
rect 37863 37303 37897 37337
rect 37897 37303 37906 37337
rect 37854 37294 37906 37303
rect 38014 37337 38066 37346
rect 38014 37303 38023 37337
rect 38023 37303 38057 37337
rect 38057 37303 38066 37337
rect 38014 37294 38066 37303
rect 38174 37337 38226 37346
rect 38174 37303 38183 37337
rect 38183 37303 38217 37337
rect 38217 37303 38226 37337
rect 38174 37294 38226 37303
rect 38334 37337 38386 37346
rect 38334 37303 38343 37337
rect 38343 37303 38377 37337
rect 38377 37303 38386 37337
rect 38334 37294 38386 37303
rect 38494 37337 38546 37346
rect 38494 37303 38503 37337
rect 38503 37303 38537 37337
rect 38537 37303 38546 37337
rect 38494 37294 38546 37303
rect 38654 37337 38706 37346
rect 38654 37303 38663 37337
rect 38663 37303 38697 37337
rect 38697 37303 38706 37337
rect 38654 37294 38706 37303
rect 38814 37337 38866 37346
rect 38814 37303 38823 37337
rect 38823 37303 38857 37337
rect 38857 37303 38866 37337
rect 38814 37294 38866 37303
rect 38974 37337 39026 37346
rect 38974 37303 38983 37337
rect 38983 37303 39017 37337
rect 39017 37303 39026 37337
rect 38974 37294 39026 37303
rect 39134 37337 39186 37346
rect 39134 37303 39143 37337
rect 39143 37303 39177 37337
rect 39177 37303 39186 37337
rect 39134 37294 39186 37303
rect 39294 37337 39346 37346
rect 39294 37303 39303 37337
rect 39303 37303 39337 37337
rect 39337 37303 39346 37337
rect 39294 37294 39346 37303
rect 39454 37337 39506 37346
rect 39454 37303 39463 37337
rect 39463 37303 39497 37337
rect 39497 37303 39506 37337
rect 39454 37294 39506 37303
rect 39614 37337 39666 37346
rect 39614 37303 39623 37337
rect 39623 37303 39657 37337
rect 39657 37303 39666 37337
rect 39614 37294 39666 37303
rect 39774 37337 39826 37346
rect 39774 37303 39783 37337
rect 39783 37303 39817 37337
rect 39817 37303 39826 37337
rect 39774 37294 39826 37303
rect 39934 37337 39986 37346
rect 39934 37303 39943 37337
rect 39943 37303 39977 37337
rect 39977 37303 39986 37337
rect 39934 37294 39986 37303
rect 40094 37337 40146 37346
rect 40094 37303 40103 37337
rect 40103 37303 40137 37337
rect 40137 37303 40146 37337
rect 40094 37294 40146 37303
rect 40254 37337 40306 37346
rect 40254 37303 40263 37337
rect 40263 37303 40297 37337
rect 40297 37303 40306 37337
rect 40254 37294 40306 37303
rect 40414 37337 40466 37346
rect 40414 37303 40423 37337
rect 40423 37303 40457 37337
rect 40457 37303 40466 37337
rect 40414 37294 40466 37303
rect 40574 37337 40626 37346
rect 40574 37303 40583 37337
rect 40583 37303 40617 37337
rect 40617 37303 40626 37337
rect 40574 37294 40626 37303
rect 40734 37337 40786 37346
rect 40734 37303 40743 37337
rect 40743 37303 40777 37337
rect 40777 37303 40786 37337
rect 40734 37294 40786 37303
rect 40894 37337 40946 37346
rect 40894 37303 40903 37337
rect 40903 37303 40937 37337
rect 40937 37303 40946 37337
rect 40894 37294 40946 37303
rect 41054 37337 41106 37346
rect 41054 37303 41063 37337
rect 41063 37303 41097 37337
rect 41097 37303 41106 37337
rect 41054 37294 41106 37303
rect 41214 37337 41266 37346
rect 41214 37303 41223 37337
rect 41223 37303 41257 37337
rect 41257 37303 41266 37337
rect 41214 37294 41266 37303
rect 41374 37337 41426 37346
rect 41374 37303 41383 37337
rect 41383 37303 41417 37337
rect 41417 37303 41426 37337
rect 41374 37294 41426 37303
rect 41534 37337 41586 37346
rect 41534 37303 41543 37337
rect 41543 37303 41577 37337
rect 41577 37303 41586 37337
rect 41534 37294 41586 37303
rect 41694 37337 41746 37346
rect 41694 37303 41703 37337
rect 41703 37303 41737 37337
rect 41737 37303 41746 37337
rect 41694 37294 41746 37303
rect 41854 37337 41906 37346
rect 41854 37303 41863 37337
rect 41863 37303 41897 37337
rect 41897 37303 41906 37337
rect 41854 37294 41906 37303
rect 14 37017 66 37026
rect 14 36983 23 37017
rect 23 36983 57 37017
rect 57 36983 66 37017
rect 14 36974 66 36983
rect 174 37017 226 37026
rect 174 36983 183 37017
rect 183 36983 217 37017
rect 217 36983 226 37017
rect 174 36974 226 36983
rect 334 37017 386 37026
rect 334 36983 343 37017
rect 343 36983 377 37017
rect 377 36983 386 37017
rect 334 36974 386 36983
rect 494 37017 546 37026
rect 494 36983 503 37017
rect 503 36983 537 37017
rect 537 36983 546 37017
rect 494 36974 546 36983
rect 654 37017 706 37026
rect 654 36983 663 37017
rect 663 36983 697 37017
rect 697 36983 706 37017
rect 654 36974 706 36983
rect 814 37017 866 37026
rect 814 36983 823 37017
rect 823 36983 857 37017
rect 857 36983 866 37017
rect 814 36974 866 36983
rect 974 37017 1026 37026
rect 974 36983 983 37017
rect 983 36983 1017 37017
rect 1017 36983 1026 37017
rect 974 36974 1026 36983
rect 1134 37017 1186 37026
rect 1134 36983 1143 37017
rect 1143 36983 1177 37017
rect 1177 36983 1186 37017
rect 1134 36974 1186 36983
rect 1294 37017 1346 37026
rect 1294 36983 1303 37017
rect 1303 36983 1337 37017
rect 1337 36983 1346 37017
rect 1294 36974 1346 36983
rect 1454 37017 1506 37026
rect 1454 36983 1463 37017
rect 1463 36983 1497 37017
rect 1497 36983 1506 37017
rect 1454 36974 1506 36983
rect 1614 37017 1666 37026
rect 1614 36983 1623 37017
rect 1623 36983 1657 37017
rect 1657 36983 1666 37017
rect 1614 36974 1666 36983
rect 1774 37017 1826 37026
rect 1774 36983 1783 37017
rect 1783 36983 1817 37017
rect 1817 36983 1826 37017
rect 1774 36974 1826 36983
rect 1934 37017 1986 37026
rect 1934 36983 1943 37017
rect 1943 36983 1977 37017
rect 1977 36983 1986 37017
rect 1934 36974 1986 36983
rect 2094 37017 2146 37026
rect 2094 36983 2103 37017
rect 2103 36983 2137 37017
rect 2137 36983 2146 37017
rect 2094 36974 2146 36983
rect 2254 37017 2306 37026
rect 2254 36983 2263 37017
rect 2263 36983 2297 37017
rect 2297 36983 2306 37017
rect 2254 36974 2306 36983
rect 2414 37017 2466 37026
rect 2414 36983 2423 37017
rect 2423 36983 2457 37017
rect 2457 36983 2466 37017
rect 2414 36974 2466 36983
rect 2574 37017 2626 37026
rect 2574 36983 2583 37017
rect 2583 36983 2617 37017
rect 2617 36983 2626 37017
rect 2574 36974 2626 36983
rect 2734 37017 2786 37026
rect 2734 36983 2743 37017
rect 2743 36983 2777 37017
rect 2777 36983 2786 37017
rect 2734 36974 2786 36983
rect 2894 37017 2946 37026
rect 2894 36983 2903 37017
rect 2903 36983 2937 37017
rect 2937 36983 2946 37017
rect 2894 36974 2946 36983
rect 3054 37017 3106 37026
rect 3054 36983 3063 37017
rect 3063 36983 3097 37017
rect 3097 36983 3106 37017
rect 3054 36974 3106 36983
rect 3214 37017 3266 37026
rect 3214 36983 3223 37017
rect 3223 36983 3257 37017
rect 3257 36983 3266 37017
rect 3214 36974 3266 36983
rect 3374 37017 3426 37026
rect 3374 36983 3383 37017
rect 3383 36983 3417 37017
rect 3417 36983 3426 37017
rect 3374 36974 3426 36983
rect 3534 37017 3586 37026
rect 3534 36983 3543 37017
rect 3543 36983 3577 37017
rect 3577 36983 3586 37017
rect 3534 36974 3586 36983
rect 3694 37017 3746 37026
rect 3694 36983 3703 37017
rect 3703 36983 3737 37017
rect 3737 36983 3746 37017
rect 3694 36974 3746 36983
rect 3854 37017 3906 37026
rect 3854 36983 3863 37017
rect 3863 36983 3897 37017
rect 3897 36983 3906 37017
rect 3854 36974 3906 36983
rect 4014 37017 4066 37026
rect 4014 36983 4023 37017
rect 4023 36983 4057 37017
rect 4057 36983 4066 37017
rect 4014 36974 4066 36983
rect 4174 37017 4226 37026
rect 4174 36983 4183 37017
rect 4183 36983 4217 37017
rect 4217 36983 4226 37017
rect 4174 36974 4226 36983
rect 4334 37017 4386 37026
rect 4334 36983 4343 37017
rect 4343 36983 4377 37017
rect 4377 36983 4386 37017
rect 4334 36974 4386 36983
rect 4494 37017 4546 37026
rect 4494 36983 4503 37017
rect 4503 36983 4537 37017
rect 4537 36983 4546 37017
rect 4494 36974 4546 36983
rect 4654 37017 4706 37026
rect 4654 36983 4663 37017
rect 4663 36983 4697 37017
rect 4697 36983 4706 37017
rect 4654 36974 4706 36983
rect 4814 37017 4866 37026
rect 4814 36983 4823 37017
rect 4823 36983 4857 37017
rect 4857 36983 4866 37017
rect 4814 36974 4866 36983
rect 4974 37017 5026 37026
rect 4974 36983 4983 37017
rect 4983 36983 5017 37017
rect 5017 36983 5026 37017
rect 4974 36974 5026 36983
rect 5134 37017 5186 37026
rect 5134 36983 5143 37017
rect 5143 36983 5177 37017
rect 5177 36983 5186 37017
rect 5134 36974 5186 36983
rect 5294 37017 5346 37026
rect 5294 36983 5303 37017
rect 5303 36983 5337 37017
rect 5337 36983 5346 37017
rect 5294 36974 5346 36983
rect 5454 37017 5506 37026
rect 5454 36983 5463 37017
rect 5463 36983 5497 37017
rect 5497 36983 5506 37017
rect 5454 36974 5506 36983
rect 5614 37017 5666 37026
rect 5614 36983 5623 37017
rect 5623 36983 5657 37017
rect 5657 36983 5666 37017
rect 5614 36974 5666 36983
rect 5774 37017 5826 37026
rect 5774 36983 5783 37017
rect 5783 36983 5817 37017
rect 5817 36983 5826 37017
rect 5774 36974 5826 36983
rect 5934 37017 5986 37026
rect 5934 36983 5943 37017
rect 5943 36983 5977 37017
rect 5977 36983 5986 37017
rect 5934 36974 5986 36983
rect 6094 37017 6146 37026
rect 6094 36983 6103 37017
rect 6103 36983 6137 37017
rect 6137 36983 6146 37017
rect 6094 36974 6146 36983
rect 6254 37017 6306 37026
rect 6254 36983 6263 37017
rect 6263 36983 6297 37017
rect 6297 36983 6306 37017
rect 6254 36974 6306 36983
rect 6414 37017 6466 37026
rect 6414 36983 6423 37017
rect 6423 36983 6457 37017
rect 6457 36983 6466 37017
rect 6414 36974 6466 36983
rect 6574 37017 6626 37026
rect 6574 36983 6583 37017
rect 6583 36983 6617 37017
rect 6617 36983 6626 37017
rect 6574 36974 6626 36983
rect 6734 37017 6786 37026
rect 6734 36983 6743 37017
rect 6743 36983 6777 37017
rect 6777 36983 6786 37017
rect 6734 36974 6786 36983
rect 6894 37017 6946 37026
rect 6894 36983 6903 37017
rect 6903 36983 6937 37017
rect 6937 36983 6946 37017
rect 6894 36974 6946 36983
rect 7054 37017 7106 37026
rect 7054 36983 7063 37017
rect 7063 36983 7097 37017
rect 7097 36983 7106 37017
rect 7054 36974 7106 36983
rect 7214 37017 7266 37026
rect 7214 36983 7223 37017
rect 7223 36983 7257 37017
rect 7257 36983 7266 37017
rect 7214 36974 7266 36983
rect 7374 37017 7426 37026
rect 7374 36983 7383 37017
rect 7383 36983 7417 37017
rect 7417 36983 7426 37017
rect 7374 36974 7426 36983
rect 7534 37017 7586 37026
rect 7534 36983 7543 37017
rect 7543 36983 7577 37017
rect 7577 36983 7586 37017
rect 7534 36974 7586 36983
rect 7694 37017 7746 37026
rect 7694 36983 7703 37017
rect 7703 36983 7737 37017
rect 7737 36983 7746 37017
rect 7694 36974 7746 36983
rect 7854 37017 7906 37026
rect 7854 36983 7863 37017
rect 7863 36983 7897 37017
rect 7897 36983 7906 37017
rect 7854 36974 7906 36983
rect 8014 37017 8066 37026
rect 8014 36983 8023 37017
rect 8023 36983 8057 37017
rect 8057 36983 8066 37017
rect 8014 36974 8066 36983
rect 8174 37017 8226 37026
rect 8174 36983 8183 37017
rect 8183 36983 8217 37017
rect 8217 36983 8226 37017
rect 8174 36974 8226 36983
rect 8334 37017 8386 37026
rect 8334 36983 8343 37017
rect 8343 36983 8377 37017
rect 8377 36983 8386 37017
rect 8334 36974 8386 36983
rect 12494 37017 12546 37026
rect 12494 36983 12503 37017
rect 12503 36983 12537 37017
rect 12537 36983 12546 37017
rect 12494 36974 12546 36983
rect 12654 37017 12706 37026
rect 12654 36983 12663 37017
rect 12663 36983 12697 37017
rect 12697 36983 12706 37017
rect 12654 36974 12706 36983
rect 12814 37017 12866 37026
rect 12814 36983 12823 37017
rect 12823 36983 12857 37017
rect 12857 36983 12866 37017
rect 12814 36974 12866 36983
rect 12974 37017 13026 37026
rect 12974 36983 12983 37017
rect 12983 36983 13017 37017
rect 13017 36983 13026 37017
rect 12974 36974 13026 36983
rect 13134 37017 13186 37026
rect 13134 36983 13143 37017
rect 13143 36983 13177 37017
rect 13177 36983 13186 37017
rect 13134 36974 13186 36983
rect 13294 37017 13346 37026
rect 13294 36983 13303 37017
rect 13303 36983 13337 37017
rect 13337 36983 13346 37017
rect 13294 36974 13346 36983
rect 13454 37017 13506 37026
rect 13454 36983 13463 37017
rect 13463 36983 13497 37017
rect 13497 36983 13506 37017
rect 13454 36974 13506 36983
rect 13614 37017 13666 37026
rect 13614 36983 13623 37017
rect 13623 36983 13657 37017
rect 13657 36983 13666 37017
rect 13614 36974 13666 36983
rect 13774 37017 13826 37026
rect 13774 36983 13783 37017
rect 13783 36983 13817 37017
rect 13817 36983 13826 37017
rect 13774 36974 13826 36983
rect 13934 37017 13986 37026
rect 13934 36983 13943 37017
rect 13943 36983 13977 37017
rect 13977 36983 13986 37017
rect 13934 36974 13986 36983
rect 14094 37017 14146 37026
rect 14094 36983 14103 37017
rect 14103 36983 14137 37017
rect 14137 36983 14146 37017
rect 14094 36974 14146 36983
rect 14254 37017 14306 37026
rect 14254 36983 14263 37017
rect 14263 36983 14297 37017
rect 14297 36983 14306 37017
rect 14254 36974 14306 36983
rect 14414 37017 14466 37026
rect 14414 36983 14423 37017
rect 14423 36983 14457 37017
rect 14457 36983 14466 37017
rect 14414 36974 14466 36983
rect 14574 37017 14626 37026
rect 14574 36983 14583 37017
rect 14583 36983 14617 37017
rect 14617 36983 14626 37017
rect 14574 36974 14626 36983
rect 14734 37017 14786 37026
rect 14734 36983 14743 37017
rect 14743 36983 14777 37017
rect 14777 36983 14786 37017
rect 14734 36974 14786 36983
rect 14894 37017 14946 37026
rect 14894 36983 14903 37017
rect 14903 36983 14937 37017
rect 14937 36983 14946 37017
rect 14894 36974 14946 36983
rect 15054 37017 15106 37026
rect 15054 36983 15063 37017
rect 15063 36983 15097 37017
rect 15097 36983 15106 37017
rect 15054 36974 15106 36983
rect 15214 37017 15266 37026
rect 15214 36983 15223 37017
rect 15223 36983 15257 37017
rect 15257 36983 15266 37017
rect 15214 36974 15266 36983
rect 15374 37017 15426 37026
rect 15374 36983 15383 37017
rect 15383 36983 15417 37017
rect 15417 36983 15426 37017
rect 15374 36974 15426 36983
rect 15534 37017 15586 37026
rect 15534 36983 15543 37017
rect 15543 36983 15577 37017
rect 15577 36983 15586 37017
rect 15534 36974 15586 36983
rect 15694 37017 15746 37026
rect 15694 36983 15703 37017
rect 15703 36983 15737 37017
rect 15737 36983 15746 37017
rect 15694 36974 15746 36983
rect 15854 37017 15906 37026
rect 15854 36983 15863 37017
rect 15863 36983 15897 37017
rect 15897 36983 15906 37017
rect 15854 36974 15906 36983
rect 16014 37017 16066 37026
rect 16014 36983 16023 37017
rect 16023 36983 16057 37017
rect 16057 36983 16066 37017
rect 16014 36974 16066 36983
rect 16174 37017 16226 37026
rect 16174 36983 16183 37017
rect 16183 36983 16217 37017
rect 16217 36983 16226 37017
rect 16174 36974 16226 36983
rect 16334 37017 16386 37026
rect 16334 36983 16343 37017
rect 16343 36983 16377 37017
rect 16377 36983 16386 37017
rect 16334 36974 16386 36983
rect 16494 37017 16546 37026
rect 16494 36983 16503 37017
rect 16503 36983 16537 37017
rect 16537 36983 16546 37017
rect 16494 36974 16546 36983
rect 16654 37017 16706 37026
rect 16654 36983 16663 37017
rect 16663 36983 16697 37017
rect 16697 36983 16706 37017
rect 16654 36974 16706 36983
rect 16814 37017 16866 37026
rect 16814 36983 16823 37017
rect 16823 36983 16857 37017
rect 16857 36983 16866 37017
rect 16814 36974 16866 36983
rect 16974 37017 17026 37026
rect 16974 36983 16983 37017
rect 16983 36983 17017 37017
rect 17017 36983 17026 37017
rect 16974 36974 17026 36983
rect 17134 37017 17186 37026
rect 17134 36983 17143 37017
rect 17143 36983 17177 37017
rect 17177 36983 17186 37017
rect 17134 36974 17186 36983
rect 17294 37017 17346 37026
rect 17294 36983 17303 37017
rect 17303 36983 17337 37017
rect 17337 36983 17346 37017
rect 17294 36974 17346 36983
rect 17454 37017 17506 37026
rect 17454 36983 17463 37017
rect 17463 36983 17497 37017
rect 17497 36983 17506 37017
rect 17454 36974 17506 36983
rect 17614 37017 17666 37026
rect 17614 36983 17623 37017
rect 17623 36983 17657 37017
rect 17657 36983 17666 37017
rect 17614 36974 17666 36983
rect 17774 37017 17826 37026
rect 17774 36983 17783 37017
rect 17783 36983 17817 37017
rect 17817 36983 17826 37017
rect 17774 36974 17826 36983
rect 17934 37017 17986 37026
rect 17934 36983 17943 37017
rect 17943 36983 17977 37017
rect 17977 36983 17986 37017
rect 17934 36974 17986 36983
rect 18094 37017 18146 37026
rect 18094 36983 18103 37017
rect 18103 36983 18137 37017
rect 18137 36983 18146 37017
rect 18094 36974 18146 36983
rect 18254 37017 18306 37026
rect 18254 36983 18263 37017
rect 18263 36983 18297 37017
rect 18297 36983 18306 37017
rect 18254 36974 18306 36983
rect 18414 37017 18466 37026
rect 18414 36983 18423 37017
rect 18423 36983 18457 37017
rect 18457 36983 18466 37017
rect 18414 36974 18466 36983
rect 18574 37017 18626 37026
rect 18574 36983 18583 37017
rect 18583 36983 18617 37017
rect 18617 36983 18626 37017
rect 18574 36974 18626 36983
rect 18734 37017 18786 37026
rect 18734 36983 18743 37017
rect 18743 36983 18777 37017
rect 18777 36983 18786 37017
rect 18734 36974 18786 36983
rect 18894 37017 18946 37026
rect 18894 36983 18903 37017
rect 18903 36983 18937 37017
rect 18937 36983 18946 37017
rect 18894 36974 18946 36983
rect 23134 37017 23186 37026
rect 23134 36983 23143 37017
rect 23143 36983 23177 37017
rect 23177 36983 23186 37017
rect 23134 36974 23186 36983
rect 23294 37017 23346 37026
rect 23294 36983 23303 37017
rect 23303 36983 23337 37017
rect 23337 36983 23346 37017
rect 23294 36974 23346 36983
rect 23454 37017 23506 37026
rect 23454 36983 23463 37017
rect 23463 36983 23497 37017
rect 23497 36983 23506 37017
rect 23454 36974 23506 36983
rect 23614 37017 23666 37026
rect 23614 36983 23623 37017
rect 23623 36983 23657 37017
rect 23657 36983 23666 37017
rect 23614 36974 23666 36983
rect 23774 37017 23826 37026
rect 23774 36983 23783 37017
rect 23783 36983 23817 37017
rect 23817 36983 23826 37017
rect 23774 36974 23826 36983
rect 23934 37017 23986 37026
rect 23934 36983 23943 37017
rect 23943 36983 23977 37017
rect 23977 36983 23986 37017
rect 23934 36974 23986 36983
rect 24094 37017 24146 37026
rect 24094 36983 24103 37017
rect 24103 36983 24137 37017
rect 24137 36983 24146 37017
rect 24094 36974 24146 36983
rect 24254 37017 24306 37026
rect 24254 36983 24263 37017
rect 24263 36983 24297 37017
rect 24297 36983 24306 37017
rect 24254 36974 24306 36983
rect 24414 37017 24466 37026
rect 24414 36983 24423 37017
rect 24423 36983 24457 37017
rect 24457 36983 24466 37017
rect 24414 36974 24466 36983
rect 24574 37017 24626 37026
rect 24574 36983 24583 37017
rect 24583 36983 24617 37017
rect 24617 36983 24626 37017
rect 24574 36974 24626 36983
rect 24734 37017 24786 37026
rect 24734 36983 24743 37017
rect 24743 36983 24777 37017
rect 24777 36983 24786 37017
rect 24734 36974 24786 36983
rect 24894 37017 24946 37026
rect 24894 36983 24903 37017
rect 24903 36983 24937 37017
rect 24937 36983 24946 37017
rect 24894 36974 24946 36983
rect 25054 37017 25106 37026
rect 25054 36983 25063 37017
rect 25063 36983 25097 37017
rect 25097 36983 25106 37017
rect 25054 36974 25106 36983
rect 25214 37017 25266 37026
rect 25214 36983 25223 37017
rect 25223 36983 25257 37017
rect 25257 36983 25266 37017
rect 25214 36974 25266 36983
rect 25374 37017 25426 37026
rect 25374 36983 25383 37017
rect 25383 36983 25417 37017
rect 25417 36983 25426 37017
rect 25374 36974 25426 36983
rect 25534 37017 25586 37026
rect 25534 36983 25543 37017
rect 25543 36983 25577 37017
rect 25577 36983 25586 37017
rect 25534 36974 25586 36983
rect 25694 37017 25746 37026
rect 25694 36983 25703 37017
rect 25703 36983 25737 37017
rect 25737 36983 25746 37017
rect 25694 36974 25746 36983
rect 25854 37017 25906 37026
rect 25854 36983 25863 37017
rect 25863 36983 25897 37017
rect 25897 36983 25906 37017
rect 25854 36974 25906 36983
rect 26014 37017 26066 37026
rect 26014 36983 26023 37017
rect 26023 36983 26057 37017
rect 26057 36983 26066 37017
rect 26014 36974 26066 36983
rect 26174 37017 26226 37026
rect 26174 36983 26183 37017
rect 26183 36983 26217 37017
rect 26217 36983 26226 37017
rect 26174 36974 26226 36983
rect 26334 37017 26386 37026
rect 26334 36983 26343 37017
rect 26343 36983 26377 37017
rect 26377 36983 26386 37017
rect 26334 36974 26386 36983
rect 26494 37017 26546 37026
rect 26494 36983 26503 37017
rect 26503 36983 26537 37017
rect 26537 36983 26546 37017
rect 26494 36974 26546 36983
rect 26654 37017 26706 37026
rect 26654 36983 26663 37017
rect 26663 36983 26697 37017
rect 26697 36983 26706 37017
rect 26654 36974 26706 36983
rect 26814 37017 26866 37026
rect 26814 36983 26823 37017
rect 26823 36983 26857 37017
rect 26857 36983 26866 37017
rect 26814 36974 26866 36983
rect 26974 37017 27026 37026
rect 26974 36983 26983 37017
rect 26983 36983 27017 37017
rect 27017 36983 27026 37017
rect 26974 36974 27026 36983
rect 27134 37017 27186 37026
rect 27134 36983 27143 37017
rect 27143 36983 27177 37017
rect 27177 36983 27186 37017
rect 27134 36974 27186 36983
rect 27294 37017 27346 37026
rect 27294 36983 27303 37017
rect 27303 36983 27337 37017
rect 27337 36983 27346 37017
rect 27294 36974 27346 36983
rect 27454 37017 27506 37026
rect 27454 36983 27463 37017
rect 27463 36983 27497 37017
rect 27497 36983 27506 37017
rect 27454 36974 27506 36983
rect 27614 37017 27666 37026
rect 27614 36983 27623 37017
rect 27623 36983 27657 37017
rect 27657 36983 27666 37017
rect 27614 36974 27666 36983
rect 27774 37017 27826 37026
rect 27774 36983 27783 37017
rect 27783 36983 27817 37017
rect 27817 36983 27826 37017
rect 27774 36974 27826 36983
rect 27934 37017 27986 37026
rect 27934 36983 27943 37017
rect 27943 36983 27977 37017
rect 27977 36983 27986 37017
rect 27934 36974 27986 36983
rect 28094 37017 28146 37026
rect 28094 36983 28103 37017
rect 28103 36983 28137 37017
rect 28137 36983 28146 37017
rect 28094 36974 28146 36983
rect 28254 37017 28306 37026
rect 28254 36983 28263 37017
rect 28263 36983 28297 37017
rect 28297 36983 28306 37017
rect 28254 36974 28306 36983
rect 28414 37017 28466 37026
rect 28414 36983 28423 37017
rect 28423 36983 28457 37017
rect 28457 36983 28466 37017
rect 28414 36974 28466 36983
rect 28574 37017 28626 37026
rect 28574 36983 28583 37017
rect 28583 36983 28617 37017
rect 28617 36983 28626 37017
rect 28574 36974 28626 36983
rect 28734 37017 28786 37026
rect 28734 36983 28743 37017
rect 28743 36983 28777 37017
rect 28777 36983 28786 37017
rect 28734 36974 28786 36983
rect 28894 37017 28946 37026
rect 28894 36983 28903 37017
rect 28903 36983 28937 37017
rect 28937 36983 28946 37017
rect 28894 36974 28946 36983
rect 29054 37017 29106 37026
rect 29054 36983 29063 37017
rect 29063 36983 29097 37017
rect 29097 36983 29106 37017
rect 29054 36974 29106 36983
rect 29214 37017 29266 37026
rect 29214 36983 29223 37017
rect 29223 36983 29257 37017
rect 29257 36983 29266 37017
rect 29214 36974 29266 36983
rect 29374 37017 29426 37026
rect 29374 36983 29383 37017
rect 29383 36983 29417 37017
rect 29417 36983 29426 37017
rect 29374 36974 29426 36983
rect 33534 37017 33586 37026
rect 33534 36983 33543 37017
rect 33543 36983 33577 37017
rect 33577 36983 33586 37017
rect 33534 36974 33586 36983
rect 33694 37017 33746 37026
rect 33694 36983 33703 37017
rect 33703 36983 33737 37017
rect 33737 36983 33746 37017
rect 33694 36974 33746 36983
rect 33854 37017 33906 37026
rect 33854 36983 33863 37017
rect 33863 36983 33897 37017
rect 33897 36983 33906 37017
rect 33854 36974 33906 36983
rect 34014 37017 34066 37026
rect 34014 36983 34023 37017
rect 34023 36983 34057 37017
rect 34057 36983 34066 37017
rect 34014 36974 34066 36983
rect 34174 37017 34226 37026
rect 34174 36983 34183 37017
rect 34183 36983 34217 37017
rect 34217 36983 34226 37017
rect 34174 36974 34226 36983
rect 34334 37017 34386 37026
rect 34334 36983 34343 37017
rect 34343 36983 34377 37017
rect 34377 36983 34386 37017
rect 34334 36974 34386 36983
rect 34494 37017 34546 37026
rect 34494 36983 34503 37017
rect 34503 36983 34537 37017
rect 34537 36983 34546 37017
rect 34494 36974 34546 36983
rect 34654 37017 34706 37026
rect 34654 36983 34663 37017
rect 34663 36983 34697 37017
rect 34697 36983 34706 37017
rect 34654 36974 34706 36983
rect 34814 37017 34866 37026
rect 34814 36983 34823 37017
rect 34823 36983 34857 37017
rect 34857 36983 34866 37017
rect 34814 36974 34866 36983
rect 34974 37017 35026 37026
rect 34974 36983 34983 37017
rect 34983 36983 35017 37017
rect 35017 36983 35026 37017
rect 34974 36974 35026 36983
rect 35134 37017 35186 37026
rect 35134 36983 35143 37017
rect 35143 36983 35177 37017
rect 35177 36983 35186 37017
rect 35134 36974 35186 36983
rect 35294 37017 35346 37026
rect 35294 36983 35303 37017
rect 35303 36983 35337 37017
rect 35337 36983 35346 37017
rect 35294 36974 35346 36983
rect 35454 37017 35506 37026
rect 35454 36983 35463 37017
rect 35463 36983 35497 37017
rect 35497 36983 35506 37017
rect 35454 36974 35506 36983
rect 35614 37017 35666 37026
rect 35614 36983 35623 37017
rect 35623 36983 35657 37017
rect 35657 36983 35666 37017
rect 35614 36974 35666 36983
rect 35774 37017 35826 37026
rect 35774 36983 35783 37017
rect 35783 36983 35817 37017
rect 35817 36983 35826 37017
rect 35774 36974 35826 36983
rect 35934 37017 35986 37026
rect 35934 36983 35943 37017
rect 35943 36983 35977 37017
rect 35977 36983 35986 37017
rect 35934 36974 35986 36983
rect 36094 37017 36146 37026
rect 36094 36983 36103 37017
rect 36103 36983 36137 37017
rect 36137 36983 36146 37017
rect 36094 36974 36146 36983
rect 36254 37017 36306 37026
rect 36254 36983 36263 37017
rect 36263 36983 36297 37017
rect 36297 36983 36306 37017
rect 36254 36974 36306 36983
rect 36414 37017 36466 37026
rect 36414 36983 36423 37017
rect 36423 36983 36457 37017
rect 36457 36983 36466 37017
rect 36414 36974 36466 36983
rect 36574 37017 36626 37026
rect 36574 36983 36583 37017
rect 36583 36983 36617 37017
rect 36617 36983 36626 37017
rect 36574 36974 36626 36983
rect 36734 37017 36786 37026
rect 36734 36983 36743 37017
rect 36743 36983 36777 37017
rect 36777 36983 36786 37017
rect 36734 36974 36786 36983
rect 36894 37017 36946 37026
rect 36894 36983 36903 37017
rect 36903 36983 36937 37017
rect 36937 36983 36946 37017
rect 36894 36974 36946 36983
rect 37054 37017 37106 37026
rect 37054 36983 37063 37017
rect 37063 36983 37097 37017
rect 37097 36983 37106 37017
rect 37054 36974 37106 36983
rect 37214 37017 37266 37026
rect 37214 36983 37223 37017
rect 37223 36983 37257 37017
rect 37257 36983 37266 37017
rect 37214 36974 37266 36983
rect 37374 37017 37426 37026
rect 37374 36983 37383 37017
rect 37383 36983 37417 37017
rect 37417 36983 37426 37017
rect 37374 36974 37426 36983
rect 37534 37017 37586 37026
rect 37534 36983 37543 37017
rect 37543 36983 37577 37017
rect 37577 36983 37586 37017
rect 37534 36974 37586 36983
rect 37694 37017 37746 37026
rect 37694 36983 37703 37017
rect 37703 36983 37737 37017
rect 37737 36983 37746 37017
rect 37694 36974 37746 36983
rect 37854 37017 37906 37026
rect 37854 36983 37863 37017
rect 37863 36983 37897 37017
rect 37897 36983 37906 37017
rect 37854 36974 37906 36983
rect 38014 37017 38066 37026
rect 38014 36983 38023 37017
rect 38023 36983 38057 37017
rect 38057 36983 38066 37017
rect 38014 36974 38066 36983
rect 38174 37017 38226 37026
rect 38174 36983 38183 37017
rect 38183 36983 38217 37017
rect 38217 36983 38226 37017
rect 38174 36974 38226 36983
rect 38334 37017 38386 37026
rect 38334 36983 38343 37017
rect 38343 36983 38377 37017
rect 38377 36983 38386 37017
rect 38334 36974 38386 36983
rect 38494 37017 38546 37026
rect 38494 36983 38503 37017
rect 38503 36983 38537 37017
rect 38537 36983 38546 37017
rect 38494 36974 38546 36983
rect 38654 37017 38706 37026
rect 38654 36983 38663 37017
rect 38663 36983 38697 37017
rect 38697 36983 38706 37017
rect 38654 36974 38706 36983
rect 38814 37017 38866 37026
rect 38814 36983 38823 37017
rect 38823 36983 38857 37017
rect 38857 36983 38866 37017
rect 38814 36974 38866 36983
rect 38974 37017 39026 37026
rect 38974 36983 38983 37017
rect 38983 36983 39017 37017
rect 39017 36983 39026 37017
rect 38974 36974 39026 36983
rect 39134 37017 39186 37026
rect 39134 36983 39143 37017
rect 39143 36983 39177 37017
rect 39177 36983 39186 37017
rect 39134 36974 39186 36983
rect 39294 37017 39346 37026
rect 39294 36983 39303 37017
rect 39303 36983 39337 37017
rect 39337 36983 39346 37017
rect 39294 36974 39346 36983
rect 39454 37017 39506 37026
rect 39454 36983 39463 37017
rect 39463 36983 39497 37017
rect 39497 36983 39506 37017
rect 39454 36974 39506 36983
rect 39614 37017 39666 37026
rect 39614 36983 39623 37017
rect 39623 36983 39657 37017
rect 39657 36983 39666 37017
rect 39614 36974 39666 36983
rect 39774 37017 39826 37026
rect 39774 36983 39783 37017
rect 39783 36983 39817 37017
rect 39817 36983 39826 37017
rect 39774 36974 39826 36983
rect 39934 37017 39986 37026
rect 39934 36983 39943 37017
rect 39943 36983 39977 37017
rect 39977 36983 39986 37017
rect 39934 36974 39986 36983
rect 40094 37017 40146 37026
rect 40094 36983 40103 37017
rect 40103 36983 40137 37017
rect 40137 36983 40146 37017
rect 40094 36974 40146 36983
rect 40254 37017 40306 37026
rect 40254 36983 40263 37017
rect 40263 36983 40297 37017
rect 40297 36983 40306 37017
rect 40254 36974 40306 36983
rect 40414 37017 40466 37026
rect 40414 36983 40423 37017
rect 40423 36983 40457 37017
rect 40457 36983 40466 37017
rect 40414 36974 40466 36983
rect 40574 37017 40626 37026
rect 40574 36983 40583 37017
rect 40583 36983 40617 37017
rect 40617 36983 40626 37017
rect 40574 36974 40626 36983
rect 40734 37017 40786 37026
rect 40734 36983 40743 37017
rect 40743 36983 40777 37017
rect 40777 36983 40786 37017
rect 40734 36974 40786 36983
rect 40894 37017 40946 37026
rect 40894 36983 40903 37017
rect 40903 36983 40937 37017
rect 40937 36983 40946 37017
rect 40894 36974 40946 36983
rect 41054 37017 41106 37026
rect 41054 36983 41063 37017
rect 41063 36983 41097 37017
rect 41097 36983 41106 37017
rect 41054 36974 41106 36983
rect 41214 37017 41266 37026
rect 41214 36983 41223 37017
rect 41223 36983 41257 37017
rect 41257 36983 41266 37017
rect 41214 36974 41266 36983
rect 41374 37017 41426 37026
rect 41374 36983 41383 37017
rect 41383 36983 41417 37017
rect 41417 36983 41426 37017
rect 41374 36974 41426 36983
rect 41534 37017 41586 37026
rect 41534 36983 41543 37017
rect 41543 36983 41577 37017
rect 41577 36983 41586 37017
rect 41534 36974 41586 36983
rect 41694 37017 41746 37026
rect 41694 36983 41703 37017
rect 41703 36983 41737 37017
rect 41737 36983 41746 37017
rect 41694 36974 41746 36983
rect 41854 37017 41906 37026
rect 41854 36983 41863 37017
rect 41863 36983 41897 37017
rect 41897 36983 41906 37017
rect 41854 36974 41906 36983
rect 14 36857 66 36866
rect 14 36823 23 36857
rect 23 36823 57 36857
rect 57 36823 66 36857
rect 14 36814 66 36823
rect 174 36857 226 36866
rect 174 36823 183 36857
rect 183 36823 217 36857
rect 217 36823 226 36857
rect 174 36814 226 36823
rect 334 36857 386 36866
rect 334 36823 343 36857
rect 343 36823 377 36857
rect 377 36823 386 36857
rect 334 36814 386 36823
rect 494 36857 546 36866
rect 494 36823 503 36857
rect 503 36823 537 36857
rect 537 36823 546 36857
rect 494 36814 546 36823
rect 654 36857 706 36866
rect 654 36823 663 36857
rect 663 36823 697 36857
rect 697 36823 706 36857
rect 654 36814 706 36823
rect 814 36857 866 36866
rect 814 36823 823 36857
rect 823 36823 857 36857
rect 857 36823 866 36857
rect 814 36814 866 36823
rect 974 36857 1026 36866
rect 974 36823 983 36857
rect 983 36823 1017 36857
rect 1017 36823 1026 36857
rect 974 36814 1026 36823
rect 1134 36857 1186 36866
rect 1134 36823 1143 36857
rect 1143 36823 1177 36857
rect 1177 36823 1186 36857
rect 1134 36814 1186 36823
rect 1294 36857 1346 36866
rect 1294 36823 1303 36857
rect 1303 36823 1337 36857
rect 1337 36823 1346 36857
rect 1294 36814 1346 36823
rect 1454 36857 1506 36866
rect 1454 36823 1463 36857
rect 1463 36823 1497 36857
rect 1497 36823 1506 36857
rect 1454 36814 1506 36823
rect 1614 36857 1666 36866
rect 1614 36823 1623 36857
rect 1623 36823 1657 36857
rect 1657 36823 1666 36857
rect 1614 36814 1666 36823
rect 1774 36857 1826 36866
rect 1774 36823 1783 36857
rect 1783 36823 1817 36857
rect 1817 36823 1826 36857
rect 1774 36814 1826 36823
rect 1934 36857 1986 36866
rect 1934 36823 1943 36857
rect 1943 36823 1977 36857
rect 1977 36823 1986 36857
rect 1934 36814 1986 36823
rect 2094 36857 2146 36866
rect 2094 36823 2103 36857
rect 2103 36823 2137 36857
rect 2137 36823 2146 36857
rect 2094 36814 2146 36823
rect 2254 36857 2306 36866
rect 2254 36823 2263 36857
rect 2263 36823 2297 36857
rect 2297 36823 2306 36857
rect 2254 36814 2306 36823
rect 2414 36857 2466 36866
rect 2414 36823 2423 36857
rect 2423 36823 2457 36857
rect 2457 36823 2466 36857
rect 2414 36814 2466 36823
rect 2574 36857 2626 36866
rect 2574 36823 2583 36857
rect 2583 36823 2617 36857
rect 2617 36823 2626 36857
rect 2574 36814 2626 36823
rect 2734 36857 2786 36866
rect 2734 36823 2743 36857
rect 2743 36823 2777 36857
rect 2777 36823 2786 36857
rect 2734 36814 2786 36823
rect 2894 36857 2946 36866
rect 2894 36823 2903 36857
rect 2903 36823 2937 36857
rect 2937 36823 2946 36857
rect 2894 36814 2946 36823
rect 3054 36857 3106 36866
rect 3054 36823 3063 36857
rect 3063 36823 3097 36857
rect 3097 36823 3106 36857
rect 3054 36814 3106 36823
rect 3214 36857 3266 36866
rect 3214 36823 3223 36857
rect 3223 36823 3257 36857
rect 3257 36823 3266 36857
rect 3214 36814 3266 36823
rect 3374 36857 3426 36866
rect 3374 36823 3383 36857
rect 3383 36823 3417 36857
rect 3417 36823 3426 36857
rect 3374 36814 3426 36823
rect 3534 36857 3586 36866
rect 3534 36823 3543 36857
rect 3543 36823 3577 36857
rect 3577 36823 3586 36857
rect 3534 36814 3586 36823
rect 3694 36857 3746 36866
rect 3694 36823 3703 36857
rect 3703 36823 3737 36857
rect 3737 36823 3746 36857
rect 3694 36814 3746 36823
rect 3854 36857 3906 36866
rect 3854 36823 3863 36857
rect 3863 36823 3897 36857
rect 3897 36823 3906 36857
rect 3854 36814 3906 36823
rect 4014 36857 4066 36866
rect 4014 36823 4023 36857
rect 4023 36823 4057 36857
rect 4057 36823 4066 36857
rect 4014 36814 4066 36823
rect 4174 36857 4226 36866
rect 4174 36823 4183 36857
rect 4183 36823 4217 36857
rect 4217 36823 4226 36857
rect 4174 36814 4226 36823
rect 4334 36857 4386 36866
rect 4334 36823 4343 36857
rect 4343 36823 4377 36857
rect 4377 36823 4386 36857
rect 4334 36814 4386 36823
rect 4494 36857 4546 36866
rect 4494 36823 4503 36857
rect 4503 36823 4537 36857
rect 4537 36823 4546 36857
rect 4494 36814 4546 36823
rect 4654 36857 4706 36866
rect 4654 36823 4663 36857
rect 4663 36823 4697 36857
rect 4697 36823 4706 36857
rect 4654 36814 4706 36823
rect 4814 36857 4866 36866
rect 4814 36823 4823 36857
rect 4823 36823 4857 36857
rect 4857 36823 4866 36857
rect 4814 36814 4866 36823
rect 4974 36857 5026 36866
rect 4974 36823 4983 36857
rect 4983 36823 5017 36857
rect 5017 36823 5026 36857
rect 4974 36814 5026 36823
rect 5134 36857 5186 36866
rect 5134 36823 5143 36857
rect 5143 36823 5177 36857
rect 5177 36823 5186 36857
rect 5134 36814 5186 36823
rect 5294 36857 5346 36866
rect 5294 36823 5303 36857
rect 5303 36823 5337 36857
rect 5337 36823 5346 36857
rect 5294 36814 5346 36823
rect 5454 36857 5506 36866
rect 5454 36823 5463 36857
rect 5463 36823 5497 36857
rect 5497 36823 5506 36857
rect 5454 36814 5506 36823
rect 5614 36857 5666 36866
rect 5614 36823 5623 36857
rect 5623 36823 5657 36857
rect 5657 36823 5666 36857
rect 5614 36814 5666 36823
rect 5774 36857 5826 36866
rect 5774 36823 5783 36857
rect 5783 36823 5817 36857
rect 5817 36823 5826 36857
rect 5774 36814 5826 36823
rect 5934 36857 5986 36866
rect 5934 36823 5943 36857
rect 5943 36823 5977 36857
rect 5977 36823 5986 36857
rect 5934 36814 5986 36823
rect 6094 36857 6146 36866
rect 6094 36823 6103 36857
rect 6103 36823 6137 36857
rect 6137 36823 6146 36857
rect 6094 36814 6146 36823
rect 6254 36857 6306 36866
rect 6254 36823 6263 36857
rect 6263 36823 6297 36857
rect 6297 36823 6306 36857
rect 6254 36814 6306 36823
rect 6414 36857 6466 36866
rect 6414 36823 6423 36857
rect 6423 36823 6457 36857
rect 6457 36823 6466 36857
rect 6414 36814 6466 36823
rect 6574 36857 6626 36866
rect 6574 36823 6583 36857
rect 6583 36823 6617 36857
rect 6617 36823 6626 36857
rect 6574 36814 6626 36823
rect 6734 36857 6786 36866
rect 6734 36823 6743 36857
rect 6743 36823 6777 36857
rect 6777 36823 6786 36857
rect 6734 36814 6786 36823
rect 6894 36857 6946 36866
rect 6894 36823 6903 36857
rect 6903 36823 6937 36857
rect 6937 36823 6946 36857
rect 6894 36814 6946 36823
rect 7054 36857 7106 36866
rect 7054 36823 7063 36857
rect 7063 36823 7097 36857
rect 7097 36823 7106 36857
rect 7054 36814 7106 36823
rect 7214 36857 7266 36866
rect 7214 36823 7223 36857
rect 7223 36823 7257 36857
rect 7257 36823 7266 36857
rect 7214 36814 7266 36823
rect 7374 36857 7426 36866
rect 7374 36823 7383 36857
rect 7383 36823 7417 36857
rect 7417 36823 7426 36857
rect 7374 36814 7426 36823
rect 7534 36857 7586 36866
rect 7534 36823 7543 36857
rect 7543 36823 7577 36857
rect 7577 36823 7586 36857
rect 7534 36814 7586 36823
rect 7694 36857 7746 36866
rect 7694 36823 7703 36857
rect 7703 36823 7737 36857
rect 7737 36823 7746 36857
rect 7694 36814 7746 36823
rect 7854 36857 7906 36866
rect 7854 36823 7863 36857
rect 7863 36823 7897 36857
rect 7897 36823 7906 36857
rect 7854 36814 7906 36823
rect 8014 36857 8066 36866
rect 8014 36823 8023 36857
rect 8023 36823 8057 36857
rect 8057 36823 8066 36857
rect 8014 36814 8066 36823
rect 8174 36857 8226 36866
rect 8174 36823 8183 36857
rect 8183 36823 8217 36857
rect 8217 36823 8226 36857
rect 8174 36814 8226 36823
rect 8334 36857 8386 36866
rect 8334 36823 8343 36857
rect 8343 36823 8377 36857
rect 8377 36823 8386 36857
rect 8334 36814 8386 36823
rect 12494 36857 12546 36866
rect 12494 36823 12503 36857
rect 12503 36823 12537 36857
rect 12537 36823 12546 36857
rect 12494 36814 12546 36823
rect 12654 36857 12706 36866
rect 12654 36823 12663 36857
rect 12663 36823 12697 36857
rect 12697 36823 12706 36857
rect 12654 36814 12706 36823
rect 12814 36857 12866 36866
rect 12814 36823 12823 36857
rect 12823 36823 12857 36857
rect 12857 36823 12866 36857
rect 12814 36814 12866 36823
rect 12974 36857 13026 36866
rect 12974 36823 12983 36857
rect 12983 36823 13017 36857
rect 13017 36823 13026 36857
rect 12974 36814 13026 36823
rect 13134 36857 13186 36866
rect 13134 36823 13143 36857
rect 13143 36823 13177 36857
rect 13177 36823 13186 36857
rect 13134 36814 13186 36823
rect 13294 36857 13346 36866
rect 13294 36823 13303 36857
rect 13303 36823 13337 36857
rect 13337 36823 13346 36857
rect 13294 36814 13346 36823
rect 13454 36857 13506 36866
rect 13454 36823 13463 36857
rect 13463 36823 13497 36857
rect 13497 36823 13506 36857
rect 13454 36814 13506 36823
rect 13614 36857 13666 36866
rect 13614 36823 13623 36857
rect 13623 36823 13657 36857
rect 13657 36823 13666 36857
rect 13614 36814 13666 36823
rect 13774 36857 13826 36866
rect 13774 36823 13783 36857
rect 13783 36823 13817 36857
rect 13817 36823 13826 36857
rect 13774 36814 13826 36823
rect 13934 36857 13986 36866
rect 13934 36823 13943 36857
rect 13943 36823 13977 36857
rect 13977 36823 13986 36857
rect 13934 36814 13986 36823
rect 14094 36857 14146 36866
rect 14094 36823 14103 36857
rect 14103 36823 14137 36857
rect 14137 36823 14146 36857
rect 14094 36814 14146 36823
rect 14254 36857 14306 36866
rect 14254 36823 14263 36857
rect 14263 36823 14297 36857
rect 14297 36823 14306 36857
rect 14254 36814 14306 36823
rect 14414 36857 14466 36866
rect 14414 36823 14423 36857
rect 14423 36823 14457 36857
rect 14457 36823 14466 36857
rect 14414 36814 14466 36823
rect 14574 36857 14626 36866
rect 14574 36823 14583 36857
rect 14583 36823 14617 36857
rect 14617 36823 14626 36857
rect 14574 36814 14626 36823
rect 14734 36857 14786 36866
rect 14734 36823 14743 36857
rect 14743 36823 14777 36857
rect 14777 36823 14786 36857
rect 14734 36814 14786 36823
rect 14894 36857 14946 36866
rect 14894 36823 14903 36857
rect 14903 36823 14937 36857
rect 14937 36823 14946 36857
rect 14894 36814 14946 36823
rect 15054 36857 15106 36866
rect 15054 36823 15063 36857
rect 15063 36823 15097 36857
rect 15097 36823 15106 36857
rect 15054 36814 15106 36823
rect 15214 36857 15266 36866
rect 15214 36823 15223 36857
rect 15223 36823 15257 36857
rect 15257 36823 15266 36857
rect 15214 36814 15266 36823
rect 15374 36857 15426 36866
rect 15374 36823 15383 36857
rect 15383 36823 15417 36857
rect 15417 36823 15426 36857
rect 15374 36814 15426 36823
rect 15534 36857 15586 36866
rect 15534 36823 15543 36857
rect 15543 36823 15577 36857
rect 15577 36823 15586 36857
rect 15534 36814 15586 36823
rect 15694 36857 15746 36866
rect 15694 36823 15703 36857
rect 15703 36823 15737 36857
rect 15737 36823 15746 36857
rect 15694 36814 15746 36823
rect 15854 36857 15906 36866
rect 15854 36823 15863 36857
rect 15863 36823 15897 36857
rect 15897 36823 15906 36857
rect 15854 36814 15906 36823
rect 16014 36857 16066 36866
rect 16014 36823 16023 36857
rect 16023 36823 16057 36857
rect 16057 36823 16066 36857
rect 16014 36814 16066 36823
rect 16174 36857 16226 36866
rect 16174 36823 16183 36857
rect 16183 36823 16217 36857
rect 16217 36823 16226 36857
rect 16174 36814 16226 36823
rect 16334 36857 16386 36866
rect 16334 36823 16343 36857
rect 16343 36823 16377 36857
rect 16377 36823 16386 36857
rect 16334 36814 16386 36823
rect 16494 36857 16546 36866
rect 16494 36823 16503 36857
rect 16503 36823 16537 36857
rect 16537 36823 16546 36857
rect 16494 36814 16546 36823
rect 16654 36857 16706 36866
rect 16654 36823 16663 36857
rect 16663 36823 16697 36857
rect 16697 36823 16706 36857
rect 16654 36814 16706 36823
rect 16814 36857 16866 36866
rect 16814 36823 16823 36857
rect 16823 36823 16857 36857
rect 16857 36823 16866 36857
rect 16814 36814 16866 36823
rect 16974 36857 17026 36866
rect 16974 36823 16983 36857
rect 16983 36823 17017 36857
rect 17017 36823 17026 36857
rect 16974 36814 17026 36823
rect 17134 36857 17186 36866
rect 17134 36823 17143 36857
rect 17143 36823 17177 36857
rect 17177 36823 17186 36857
rect 17134 36814 17186 36823
rect 17294 36857 17346 36866
rect 17294 36823 17303 36857
rect 17303 36823 17337 36857
rect 17337 36823 17346 36857
rect 17294 36814 17346 36823
rect 17454 36857 17506 36866
rect 17454 36823 17463 36857
rect 17463 36823 17497 36857
rect 17497 36823 17506 36857
rect 17454 36814 17506 36823
rect 17614 36857 17666 36866
rect 17614 36823 17623 36857
rect 17623 36823 17657 36857
rect 17657 36823 17666 36857
rect 17614 36814 17666 36823
rect 17774 36857 17826 36866
rect 17774 36823 17783 36857
rect 17783 36823 17817 36857
rect 17817 36823 17826 36857
rect 17774 36814 17826 36823
rect 17934 36857 17986 36866
rect 17934 36823 17943 36857
rect 17943 36823 17977 36857
rect 17977 36823 17986 36857
rect 17934 36814 17986 36823
rect 18094 36857 18146 36866
rect 18094 36823 18103 36857
rect 18103 36823 18137 36857
rect 18137 36823 18146 36857
rect 18094 36814 18146 36823
rect 18254 36857 18306 36866
rect 18254 36823 18263 36857
rect 18263 36823 18297 36857
rect 18297 36823 18306 36857
rect 18254 36814 18306 36823
rect 18414 36857 18466 36866
rect 18414 36823 18423 36857
rect 18423 36823 18457 36857
rect 18457 36823 18466 36857
rect 18414 36814 18466 36823
rect 18574 36857 18626 36866
rect 18574 36823 18583 36857
rect 18583 36823 18617 36857
rect 18617 36823 18626 36857
rect 18574 36814 18626 36823
rect 18734 36857 18786 36866
rect 18734 36823 18743 36857
rect 18743 36823 18777 36857
rect 18777 36823 18786 36857
rect 18734 36814 18786 36823
rect 18894 36857 18946 36866
rect 18894 36823 18903 36857
rect 18903 36823 18937 36857
rect 18937 36823 18946 36857
rect 18894 36814 18946 36823
rect 23134 36857 23186 36866
rect 23134 36823 23143 36857
rect 23143 36823 23177 36857
rect 23177 36823 23186 36857
rect 23134 36814 23186 36823
rect 23294 36857 23346 36866
rect 23294 36823 23303 36857
rect 23303 36823 23337 36857
rect 23337 36823 23346 36857
rect 23294 36814 23346 36823
rect 23454 36857 23506 36866
rect 23454 36823 23463 36857
rect 23463 36823 23497 36857
rect 23497 36823 23506 36857
rect 23454 36814 23506 36823
rect 23614 36857 23666 36866
rect 23614 36823 23623 36857
rect 23623 36823 23657 36857
rect 23657 36823 23666 36857
rect 23614 36814 23666 36823
rect 23774 36857 23826 36866
rect 23774 36823 23783 36857
rect 23783 36823 23817 36857
rect 23817 36823 23826 36857
rect 23774 36814 23826 36823
rect 23934 36857 23986 36866
rect 23934 36823 23943 36857
rect 23943 36823 23977 36857
rect 23977 36823 23986 36857
rect 23934 36814 23986 36823
rect 24094 36857 24146 36866
rect 24094 36823 24103 36857
rect 24103 36823 24137 36857
rect 24137 36823 24146 36857
rect 24094 36814 24146 36823
rect 24254 36857 24306 36866
rect 24254 36823 24263 36857
rect 24263 36823 24297 36857
rect 24297 36823 24306 36857
rect 24254 36814 24306 36823
rect 24414 36857 24466 36866
rect 24414 36823 24423 36857
rect 24423 36823 24457 36857
rect 24457 36823 24466 36857
rect 24414 36814 24466 36823
rect 24574 36857 24626 36866
rect 24574 36823 24583 36857
rect 24583 36823 24617 36857
rect 24617 36823 24626 36857
rect 24574 36814 24626 36823
rect 24734 36857 24786 36866
rect 24734 36823 24743 36857
rect 24743 36823 24777 36857
rect 24777 36823 24786 36857
rect 24734 36814 24786 36823
rect 24894 36857 24946 36866
rect 24894 36823 24903 36857
rect 24903 36823 24937 36857
rect 24937 36823 24946 36857
rect 24894 36814 24946 36823
rect 25054 36857 25106 36866
rect 25054 36823 25063 36857
rect 25063 36823 25097 36857
rect 25097 36823 25106 36857
rect 25054 36814 25106 36823
rect 25214 36857 25266 36866
rect 25214 36823 25223 36857
rect 25223 36823 25257 36857
rect 25257 36823 25266 36857
rect 25214 36814 25266 36823
rect 25374 36857 25426 36866
rect 25374 36823 25383 36857
rect 25383 36823 25417 36857
rect 25417 36823 25426 36857
rect 25374 36814 25426 36823
rect 25534 36857 25586 36866
rect 25534 36823 25543 36857
rect 25543 36823 25577 36857
rect 25577 36823 25586 36857
rect 25534 36814 25586 36823
rect 25694 36857 25746 36866
rect 25694 36823 25703 36857
rect 25703 36823 25737 36857
rect 25737 36823 25746 36857
rect 25694 36814 25746 36823
rect 25854 36857 25906 36866
rect 25854 36823 25863 36857
rect 25863 36823 25897 36857
rect 25897 36823 25906 36857
rect 25854 36814 25906 36823
rect 26014 36857 26066 36866
rect 26014 36823 26023 36857
rect 26023 36823 26057 36857
rect 26057 36823 26066 36857
rect 26014 36814 26066 36823
rect 26174 36857 26226 36866
rect 26174 36823 26183 36857
rect 26183 36823 26217 36857
rect 26217 36823 26226 36857
rect 26174 36814 26226 36823
rect 26334 36857 26386 36866
rect 26334 36823 26343 36857
rect 26343 36823 26377 36857
rect 26377 36823 26386 36857
rect 26334 36814 26386 36823
rect 26494 36857 26546 36866
rect 26494 36823 26503 36857
rect 26503 36823 26537 36857
rect 26537 36823 26546 36857
rect 26494 36814 26546 36823
rect 26654 36857 26706 36866
rect 26654 36823 26663 36857
rect 26663 36823 26697 36857
rect 26697 36823 26706 36857
rect 26654 36814 26706 36823
rect 26814 36857 26866 36866
rect 26814 36823 26823 36857
rect 26823 36823 26857 36857
rect 26857 36823 26866 36857
rect 26814 36814 26866 36823
rect 26974 36857 27026 36866
rect 26974 36823 26983 36857
rect 26983 36823 27017 36857
rect 27017 36823 27026 36857
rect 26974 36814 27026 36823
rect 27134 36857 27186 36866
rect 27134 36823 27143 36857
rect 27143 36823 27177 36857
rect 27177 36823 27186 36857
rect 27134 36814 27186 36823
rect 27294 36857 27346 36866
rect 27294 36823 27303 36857
rect 27303 36823 27337 36857
rect 27337 36823 27346 36857
rect 27294 36814 27346 36823
rect 27454 36857 27506 36866
rect 27454 36823 27463 36857
rect 27463 36823 27497 36857
rect 27497 36823 27506 36857
rect 27454 36814 27506 36823
rect 27614 36857 27666 36866
rect 27614 36823 27623 36857
rect 27623 36823 27657 36857
rect 27657 36823 27666 36857
rect 27614 36814 27666 36823
rect 27774 36857 27826 36866
rect 27774 36823 27783 36857
rect 27783 36823 27817 36857
rect 27817 36823 27826 36857
rect 27774 36814 27826 36823
rect 27934 36857 27986 36866
rect 27934 36823 27943 36857
rect 27943 36823 27977 36857
rect 27977 36823 27986 36857
rect 27934 36814 27986 36823
rect 28094 36857 28146 36866
rect 28094 36823 28103 36857
rect 28103 36823 28137 36857
rect 28137 36823 28146 36857
rect 28094 36814 28146 36823
rect 28254 36857 28306 36866
rect 28254 36823 28263 36857
rect 28263 36823 28297 36857
rect 28297 36823 28306 36857
rect 28254 36814 28306 36823
rect 28414 36857 28466 36866
rect 28414 36823 28423 36857
rect 28423 36823 28457 36857
rect 28457 36823 28466 36857
rect 28414 36814 28466 36823
rect 28574 36857 28626 36866
rect 28574 36823 28583 36857
rect 28583 36823 28617 36857
rect 28617 36823 28626 36857
rect 28574 36814 28626 36823
rect 28734 36857 28786 36866
rect 28734 36823 28743 36857
rect 28743 36823 28777 36857
rect 28777 36823 28786 36857
rect 28734 36814 28786 36823
rect 28894 36857 28946 36866
rect 28894 36823 28903 36857
rect 28903 36823 28937 36857
rect 28937 36823 28946 36857
rect 28894 36814 28946 36823
rect 29054 36857 29106 36866
rect 29054 36823 29063 36857
rect 29063 36823 29097 36857
rect 29097 36823 29106 36857
rect 29054 36814 29106 36823
rect 29214 36857 29266 36866
rect 29214 36823 29223 36857
rect 29223 36823 29257 36857
rect 29257 36823 29266 36857
rect 29214 36814 29266 36823
rect 29374 36857 29426 36866
rect 29374 36823 29383 36857
rect 29383 36823 29417 36857
rect 29417 36823 29426 36857
rect 29374 36814 29426 36823
rect 33534 36857 33586 36866
rect 33534 36823 33543 36857
rect 33543 36823 33577 36857
rect 33577 36823 33586 36857
rect 33534 36814 33586 36823
rect 33694 36857 33746 36866
rect 33694 36823 33703 36857
rect 33703 36823 33737 36857
rect 33737 36823 33746 36857
rect 33694 36814 33746 36823
rect 33854 36857 33906 36866
rect 33854 36823 33863 36857
rect 33863 36823 33897 36857
rect 33897 36823 33906 36857
rect 33854 36814 33906 36823
rect 34014 36857 34066 36866
rect 34014 36823 34023 36857
rect 34023 36823 34057 36857
rect 34057 36823 34066 36857
rect 34014 36814 34066 36823
rect 34174 36857 34226 36866
rect 34174 36823 34183 36857
rect 34183 36823 34217 36857
rect 34217 36823 34226 36857
rect 34174 36814 34226 36823
rect 34334 36857 34386 36866
rect 34334 36823 34343 36857
rect 34343 36823 34377 36857
rect 34377 36823 34386 36857
rect 34334 36814 34386 36823
rect 34494 36857 34546 36866
rect 34494 36823 34503 36857
rect 34503 36823 34537 36857
rect 34537 36823 34546 36857
rect 34494 36814 34546 36823
rect 34654 36857 34706 36866
rect 34654 36823 34663 36857
rect 34663 36823 34697 36857
rect 34697 36823 34706 36857
rect 34654 36814 34706 36823
rect 34814 36857 34866 36866
rect 34814 36823 34823 36857
rect 34823 36823 34857 36857
rect 34857 36823 34866 36857
rect 34814 36814 34866 36823
rect 34974 36857 35026 36866
rect 34974 36823 34983 36857
rect 34983 36823 35017 36857
rect 35017 36823 35026 36857
rect 34974 36814 35026 36823
rect 35134 36857 35186 36866
rect 35134 36823 35143 36857
rect 35143 36823 35177 36857
rect 35177 36823 35186 36857
rect 35134 36814 35186 36823
rect 35294 36857 35346 36866
rect 35294 36823 35303 36857
rect 35303 36823 35337 36857
rect 35337 36823 35346 36857
rect 35294 36814 35346 36823
rect 35454 36857 35506 36866
rect 35454 36823 35463 36857
rect 35463 36823 35497 36857
rect 35497 36823 35506 36857
rect 35454 36814 35506 36823
rect 35614 36857 35666 36866
rect 35614 36823 35623 36857
rect 35623 36823 35657 36857
rect 35657 36823 35666 36857
rect 35614 36814 35666 36823
rect 35774 36857 35826 36866
rect 35774 36823 35783 36857
rect 35783 36823 35817 36857
rect 35817 36823 35826 36857
rect 35774 36814 35826 36823
rect 35934 36857 35986 36866
rect 35934 36823 35943 36857
rect 35943 36823 35977 36857
rect 35977 36823 35986 36857
rect 35934 36814 35986 36823
rect 36094 36857 36146 36866
rect 36094 36823 36103 36857
rect 36103 36823 36137 36857
rect 36137 36823 36146 36857
rect 36094 36814 36146 36823
rect 36254 36857 36306 36866
rect 36254 36823 36263 36857
rect 36263 36823 36297 36857
rect 36297 36823 36306 36857
rect 36254 36814 36306 36823
rect 36414 36857 36466 36866
rect 36414 36823 36423 36857
rect 36423 36823 36457 36857
rect 36457 36823 36466 36857
rect 36414 36814 36466 36823
rect 36574 36857 36626 36866
rect 36574 36823 36583 36857
rect 36583 36823 36617 36857
rect 36617 36823 36626 36857
rect 36574 36814 36626 36823
rect 36734 36857 36786 36866
rect 36734 36823 36743 36857
rect 36743 36823 36777 36857
rect 36777 36823 36786 36857
rect 36734 36814 36786 36823
rect 36894 36857 36946 36866
rect 36894 36823 36903 36857
rect 36903 36823 36937 36857
rect 36937 36823 36946 36857
rect 36894 36814 36946 36823
rect 37054 36857 37106 36866
rect 37054 36823 37063 36857
rect 37063 36823 37097 36857
rect 37097 36823 37106 36857
rect 37054 36814 37106 36823
rect 37214 36857 37266 36866
rect 37214 36823 37223 36857
rect 37223 36823 37257 36857
rect 37257 36823 37266 36857
rect 37214 36814 37266 36823
rect 37374 36857 37426 36866
rect 37374 36823 37383 36857
rect 37383 36823 37417 36857
rect 37417 36823 37426 36857
rect 37374 36814 37426 36823
rect 37534 36857 37586 36866
rect 37534 36823 37543 36857
rect 37543 36823 37577 36857
rect 37577 36823 37586 36857
rect 37534 36814 37586 36823
rect 37694 36857 37746 36866
rect 37694 36823 37703 36857
rect 37703 36823 37737 36857
rect 37737 36823 37746 36857
rect 37694 36814 37746 36823
rect 37854 36857 37906 36866
rect 37854 36823 37863 36857
rect 37863 36823 37897 36857
rect 37897 36823 37906 36857
rect 37854 36814 37906 36823
rect 38014 36857 38066 36866
rect 38014 36823 38023 36857
rect 38023 36823 38057 36857
rect 38057 36823 38066 36857
rect 38014 36814 38066 36823
rect 38174 36857 38226 36866
rect 38174 36823 38183 36857
rect 38183 36823 38217 36857
rect 38217 36823 38226 36857
rect 38174 36814 38226 36823
rect 38334 36857 38386 36866
rect 38334 36823 38343 36857
rect 38343 36823 38377 36857
rect 38377 36823 38386 36857
rect 38334 36814 38386 36823
rect 38494 36857 38546 36866
rect 38494 36823 38503 36857
rect 38503 36823 38537 36857
rect 38537 36823 38546 36857
rect 38494 36814 38546 36823
rect 38654 36857 38706 36866
rect 38654 36823 38663 36857
rect 38663 36823 38697 36857
rect 38697 36823 38706 36857
rect 38654 36814 38706 36823
rect 38814 36857 38866 36866
rect 38814 36823 38823 36857
rect 38823 36823 38857 36857
rect 38857 36823 38866 36857
rect 38814 36814 38866 36823
rect 38974 36857 39026 36866
rect 38974 36823 38983 36857
rect 38983 36823 39017 36857
rect 39017 36823 39026 36857
rect 38974 36814 39026 36823
rect 39134 36857 39186 36866
rect 39134 36823 39143 36857
rect 39143 36823 39177 36857
rect 39177 36823 39186 36857
rect 39134 36814 39186 36823
rect 39294 36857 39346 36866
rect 39294 36823 39303 36857
rect 39303 36823 39337 36857
rect 39337 36823 39346 36857
rect 39294 36814 39346 36823
rect 39454 36857 39506 36866
rect 39454 36823 39463 36857
rect 39463 36823 39497 36857
rect 39497 36823 39506 36857
rect 39454 36814 39506 36823
rect 39614 36857 39666 36866
rect 39614 36823 39623 36857
rect 39623 36823 39657 36857
rect 39657 36823 39666 36857
rect 39614 36814 39666 36823
rect 39774 36857 39826 36866
rect 39774 36823 39783 36857
rect 39783 36823 39817 36857
rect 39817 36823 39826 36857
rect 39774 36814 39826 36823
rect 39934 36857 39986 36866
rect 39934 36823 39943 36857
rect 39943 36823 39977 36857
rect 39977 36823 39986 36857
rect 39934 36814 39986 36823
rect 40094 36857 40146 36866
rect 40094 36823 40103 36857
rect 40103 36823 40137 36857
rect 40137 36823 40146 36857
rect 40094 36814 40146 36823
rect 40254 36857 40306 36866
rect 40254 36823 40263 36857
rect 40263 36823 40297 36857
rect 40297 36823 40306 36857
rect 40254 36814 40306 36823
rect 40414 36857 40466 36866
rect 40414 36823 40423 36857
rect 40423 36823 40457 36857
rect 40457 36823 40466 36857
rect 40414 36814 40466 36823
rect 40574 36857 40626 36866
rect 40574 36823 40583 36857
rect 40583 36823 40617 36857
rect 40617 36823 40626 36857
rect 40574 36814 40626 36823
rect 40734 36857 40786 36866
rect 40734 36823 40743 36857
rect 40743 36823 40777 36857
rect 40777 36823 40786 36857
rect 40734 36814 40786 36823
rect 40894 36857 40946 36866
rect 40894 36823 40903 36857
rect 40903 36823 40937 36857
rect 40937 36823 40946 36857
rect 40894 36814 40946 36823
rect 41054 36857 41106 36866
rect 41054 36823 41063 36857
rect 41063 36823 41097 36857
rect 41097 36823 41106 36857
rect 41054 36814 41106 36823
rect 41214 36857 41266 36866
rect 41214 36823 41223 36857
rect 41223 36823 41257 36857
rect 41257 36823 41266 36857
rect 41214 36814 41266 36823
rect 41374 36857 41426 36866
rect 41374 36823 41383 36857
rect 41383 36823 41417 36857
rect 41417 36823 41426 36857
rect 41374 36814 41426 36823
rect 41534 36857 41586 36866
rect 41534 36823 41543 36857
rect 41543 36823 41577 36857
rect 41577 36823 41586 36857
rect 41534 36814 41586 36823
rect 41694 36857 41746 36866
rect 41694 36823 41703 36857
rect 41703 36823 41737 36857
rect 41737 36823 41746 36857
rect 41694 36814 41746 36823
rect 41854 36857 41906 36866
rect 41854 36823 41863 36857
rect 41863 36823 41897 36857
rect 41897 36823 41906 36857
rect 41854 36814 41906 36823
rect 14 36537 66 36546
rect 14 36503 23 36537
rect 23 36503 57 36537
rect 57 36503 66 36537
rect 14 36494 66 36503
rect 174 36537 226 36546
rect 174 36503 183 36537
rect 183 36503 217 36537
rect 217 36503 226 36537
rect 174 36494 226 36503
rect 334 36537 386 36546
rect 334 36503 343 36537
rect 343 36503 377 36537
rect 377 36503 386 36537
rect 334 36494 386 36503
rect 494 36537 546 36546
rect 494 36503 503 36537
rect 503 36503 537 36537
rect 537 36503 546 36537
rect 494 36494 546 36503
rect 654 36537 706 36546
rect 654 36503 663 36537
rect 663 36503 697 36537
rect 697 36503 706 36537
rect 654 36494 706 36503
rect 814 36537 866 36546
rect 814 36503 823 36537
rect 823 36503 857 36537
rect 857 36503 866 36537
rect 814 36494 866 36503
rect 974 36537 1026 36546
rect 974 36503 983 36537
rect 983 36503 1017 36537
rect 1017 36503 1026 36537
rect 974 36494 1026 36503
rect 1134 36537 1186 36546
rect 1134 36503 1143 36537
rect 1143 36503 1177 36537
rect 1177 36503 1186 36537
rect 1134 36494 1186 36503
rect 1294 36537 1346 36546
rect 1294 36503 1303 36537
rect 1303 36503 1337 36537
rect 1337 36503 1346 36537
rect 1294 36494 1346 36503
rect 1454 36537 1506 36546
rect 1454 36503 1463 36537
rect 1463 36503 1497 36537
rect 1497 36503 1506 36537
rect 1454 36494 1506 36503
rect 1614 36537 1666 36546
rect 1614 36503 1623 36537
rect 1623 36503 1657 36537
rect 1657 36503 1666 36537
rect 1614 36494 1666 36503
rect 1774 36537 1826 36546
rect 1774 36503 1783 36537
rect 1783 36503 1817 36537
rect 1817 36503 1826 36537
rect 1774 36494 1826 36503
rect 1934 36537 1986 36546
rect 1934 36503 1943 36537
rect 1943 36503 1977 36537
rect 1977 36503 1986 36537
rect 1934 36494 1986 36503
rect 2094 36537 2146 36546
rect 2094 36503 2103 36537
rect 2103 36503 2137 36537
rect 2137 36503 2146 36537
rect 2094 36494 2146 36503
rect 2254 36537 2306 36546
rect 2254 36503 2263 36537
rect 2263 36503 2297 36537
rect 2297 36503 2306 36537
rect 2254 36494 2306 36503
rect 2414 36537 2466 36546
rect 2414 36503 2423 36537
rect 2423 36503 2457 36537
rect 2457 36503 2466 36537
rect 2414 36494 2466 36503
rect 2574 36537 2626 36546
rect 2574 36503 2583 36537
rect 2583 36503 2617 36537
rect 2617 36503 2626 36537
rect 2574 36494 2626 36503
rect 2734 36537 2786 36546
rect 2734 36503 2743 36537
rect 2743 36503 2777 36537
rect 2777 36503 2786 36537
rect 2734 36494 2786 36503
rect 2894 36537 2946 36546
rect 2894 36503 2903 36537
rect 2903 36503 2937 36537
rect 2937 36503 2946 36537
rect 2894 36494 2946 36503
rect 3054 36537 3106 36546
rect 3054 36503 3063 36537
rect 3063 36503 3097 36537
rect 3097 36503 3106 36537
rect 3054 36494 3106 36503
rect 3214 36537 3266 36546
rect 3214 36503 3223 36537
rect 3223 36503 3257 36537
rect 3257 36503 3266 36537
rect 3214 36494 3266 36503
rect 3374 36537 3426 36546
rect 3374 36503 3383 36537
rect 3383 36503 3417 36537
rect 3417 36503 3426 36537
rect 3374 36494 3426 36503
rect 3534 36537 3586 36546
rect 3534 36503 3543 36537
rect 3543 36503 3577 36537
rect 3577 36503 3586 36537
rect 3534 36494 3586 36503
rect 3694 36537 3746 36546
rect 3694 36503 3703 36537
rect 3703 36503 3737 36537
rect 3737 36503 3746 36537
rect 3694 36494 3746 36503
rect 3854 36537 3906 36546
rect 3854 36503 3863 36537
rect 3863 36503 3897 36537
rect 3897 36503 3906 36537
rect 3854 36494 3906 36503
rect 4014 36537 4066 36546
rect 4014 36503 4023 36537
rect 4023 36503 4057 36537
rect 4057 36503 4066 36537
rect 4014 36494 4066 36503
rect 4174 36537 4226 36546
rect 4174 36503 4183 36537
rect 4183 36503 4217 36537
rect 4217 36503 4226 36537
rect 4174 36494 4226 36503
rect 4334 36537 4386 36546
rect 4334 36503 4343 36537
rect 4343 36503 4377 36537
rect 4377 36503 4386 36537
rect 4334 36494 4386 36503
rect 4494 36537 4546 36546
rect 4494 36503 4503 36537
rect 4503 36503 4537 36537
rect 4537 36503 4546 36537
rect 4494 36494 4546 36503
rect 4654 36537 4706 36546
rect 4654 36503 4663 36537
rect 4663 36503 4697 36537
rect 4697 36503 4706 36537
rect 4654 36494 4706 36503
rect 4814 36537 4866 36546
rect 4814 36503 4823 36537
rect 4823 36503 4857 36537
rect 4857 36503 4866 36537
rect 4814 36494 4866 36503
rect 4974 36537 5026 36546
rect 4974 36503 4983 36537
rect 4983 36503 5017 36537
rect 5017 36503 5026 36537
rect 4974 36494 5026 36503
rect 5134 36537 5186 36546
rect 5134 36503 5143 36537
rect 5143 36503 5177 36537
rect 5177 36503 5186 36537
rect 5134 36494 5186 36503
rect 5294 36537 5346 36546
rect 5294 36503 5303 36537
rect 5303 36503 5337 36537
rect 5337 36503 5346 36537
rect 5294 36494 5346 36503
rect 5454 36537 5506 36546
rect 5454 36503 5463 36537
rect 5463 36503 5497 36537
rect 5497 36503 5506 36537
rect 5454 36494 5506 36503
rect 5614 36537 5666 36546
rect 5614 36503 5623 36537
rect 5623 36503 5657 36537
rect 5657 36503 5666 36537
rect 5614 36494 5666 36503
rect 5774 36537 5826 36546
rect 5774 36503 5783 36537
rect 5783 36503 5817 36537
rect 5817 36503 5826 36537
rect 5774 36494 5826 36503
rect 5934 36537 5986 36546
rect 5934 36503 5943 36537
rect 5943 36503 5977 36537
rect 5977 36503 5986 36537
rect 5934 36494 5986 36503
rect 6094 36537 6146 36546
rect 6094 36503 6103 36537
rect 6103 36503 6137 36537
rect 6137 36503 6146 36537
rect 6094 36494 6146 36503
rect 6254 36537 6306 36546
rect 6254 36503 6263 36537
rect 6263 36503 6297 36537
rect 6297 36503 6306 36537
rect 6254 36494 6306 36503
rect 6414 36537 6466 36546
rect 6414 36503 6423 36537
rect 6423 36503 6457 36537
rect 6457 36503 6466 36537
rect 6414 36494 6466 36503
rect 6574 36537 6626 36546
rect 6574 36503 6583 36537
rect 6583 36503 6617 36537
rect 6617 36503 6626 36537
rect 6574 36494 6626 36503
rect 6734 36537 6786 36546
rect 6734 36503 6743 36537
rect 6743 36503 6777 36537
rect 6777 36503 6786 36537
rect 6734 36494 6786 36503
rect 6894 36537 6946 36546
rect 6894 36503 6903 36537
rect 6903 36503 6937 36537
rect 6937 36503 6946 36537
rect 6894 36494 6946 36503
rect 7054 36537 7106 36546
rect 7054 36503 7063 36537
rect 7063 36503 7097 36537
rect 7097 36503 7106 36537
rect 7054 36494 7106 36503
rect 7214 36537 7266 36546
rect 7214 36503 7223 36537
rect 7223 36503 7257 36537
rect 7257 36503 7266 36537
rect 7214 36494 7266 36503
rect 7374 36537 7426 36546
rect 7374 36503 7383 36537
rect 7383 36503 7417 36537
rect 7417 36503 7426 36537
rect 7374 36494 7426 36503
rect 7534 36537 7586 36546
rect 7534 36503 7543 36537
rect 7543 36503 7577 36537
rect 7577 36503 7586 36537
rect 7534 36494 7586 36503
rect 7694 36537 7746 36546
rect 7694 36503 7703 36537
rect 7703 36503 7737 36537
rect 7737 36503 7746 36537
rect 7694 36494 7746 36503
rect 7854 36537 7906 36546
rect 7854 36503 7863 36537
rect 7863 36503 7897 36537
rect 7897 36503 7906 36537
rect 7854 36494 7906 36503
rect 8014 36537 8066 36546
rect 8014 36503 8023 36537
rect 8023 36503 8057 36537
rect 8057 36503 8066 36537
rect 8014 36494 8066 36503
rect 8174 36537 8226 36546
rect 8174 36503 8183 36537
rect 8183 36503 8217 36537
rect 8217 36503 8226 36537
rect 8174 36494 8226 36503
rect 8334 36537 8386 36546
rect 8334 36503 8343 36537
rect 8343 36503 8377 36537
rect 8377 36503 8386 36537
rect 8334 36494 8386 36503
rect 12494 36537 12546 36546
rect 12494 36503 12503 36537
rect 12503 36503 12537 36537
rect 12537 36503 12546 36537
rect 12494 36494 12546 36503
rect 12654 36537 12706 36546
rect 12654 36503 12663 36537
rect 12663 36503 12697 36537
rect 12697 36503 12706 36537
rect 12654 36494 12706 36503
rect 12814 36537 12866 36546
rect 12814 36503 12823 36537
rect 12823 36503 12857 36537
rect 12857 36503 12866 36537
rect 12814 36494 12866 36503
rect 12974 36537 13026 36546
rect 12974 36503 12983 36537
rect 12983 36503 13017 36537
rect 13017 36503 13026 36537
rect 12974 36494 13026 36503
rect 13134 36537 13186 36546
rect 13134 36503 13143 36537
rect 13143 36503 13177 36537
rect 13177 36503 13186 36537
rect 13134 36494 13186 36503
rect 13294 36537 13346 36546
rect 13294 36503 13303 36537
rect 13303 36503 13337 36537
rect 13337 36503 13346 36537
rect 13294 36494 13346 36503
rect 13454 36537 13506 36546
rect 13454 36503 13463 36537
rect 13463 36503 13497 36537
rect 13497 36503 13506 36537
rect 13454 36494 13506 36503
rect 13614 36537 13666 36546
rect 13614 36503 13623 36537
rect 13623 36503 13657 36537
rect 13657 36503 13666 36537
rect 13614 36494 13666 36503
rect 13774 36537 13826 36546
rect 13774 36503 13783 36537
rect 13783 36503 13817 36537
rect 13817 36503 13826 36537
rect 13774 36494 13826 36503
rect 13934 36537 13986 36546
rect 13934 36503 13943 36537
rect 13943 36503 13977 36537
rect 13977 36503 13986 36537
rect 13934 36494 13986 36503
rect 14094 36537 14146 36546
rect 14094 36503 14103 36537
rect 14103 36503 14137 36537
rect 14137 36503 14146 36537
rect 14094 36494 14146 36503
rect 14254 36537 14306 36546
rect 14254 36503 14263 36537
rect 14263 36503 14297 36537
rect 14297 36503 14306 36537
rect 14254 36494 14306 36503
rect 14414 36537 14466 36546
rect 14414 36503 14423 36537
rect 14423 36503 14457 36537
rect 14457 36503 14466 36537
rect 14414 36494 14466 36503
rect 14574 36537 14626 36546
rect 14574 36503 14583 36537
rect 14583 36503 14617 36537
rect 14617 36503 14626 36537
rect 14574 36494 14626 36503
rect 14734 36537 14786 36546
rect 14734 36503 14743 36537
rect 14743 36503 14777 36537
rect 14777 36503 14786 36537
rect 14734 36494 14786 36503
rect 14894 36537 14946 36546
rect 14894 36503 14903 36537
rect 14903 36503 14937 36537
rect 14937 36503 14946 36537
rect 14894 36494 14946 36503
rect 15054 36537 15106 36546
rect 15054 36503 15063 36537
rect 15063 36503 15097 36537
rect 15097 36503 15106 36537
rect 15054 36494 15106 36503
rect 15214 36537 15266 36546
rect 15214 36503 15223 36537
rect 15223 36503 15257 36537
rect 15257 36503 15266 36537
rect 15214 36494 15266 36503
rect 15374 36537 15426 36546
rect 15374 36503 15383 36537
rect 15383 36503 15417 36537
rect 15417 36503 15426 36537
rect 15374 36494 15426 36503
rect 15534 36537 15586 36546
rect 15534 36503 15543 36537
rect 15543 36503 15577 36537
rect 15577 36503 15586 36537
rect 15534 36494 15586 36503
rect 15694 36537 15746 36546
rect 15694 36503 15703 36537
rect 15703 36503 15737 36537
rect 15737 36503 15746 36537
rect 15694 36494 15746 36503
rect 15854 36537 15906 36546
rect 15854 36503 15863 36537
rect 15863 36503 15897 36537
rect 15897 36503 15906 36537
rect 15854 36494 15906 36503
rect 16014 36537 16066 36546
rect 16014 36503 16023 36537
rect 16023 36503 16057 36537
rect 16057 36503 16066 36537
rect 16014 36494 16066 36503
rect 16174 36537 16226 36546
rect 16174 36503 16183 36537
rect 16183 36503 16217 36537
rect 16217 36503 16226 36537
rect 16174 36494 16226 36503
rect 16334 36537 16386 36546
rect 16334 36503 16343 36537
rect 16343 36503 16377 36537
rect 16377 36503 16386 36537
rect 16334 36494 16386 36503
rect 16494 36537 16546 36546
rect 16494 36503 16503 36537
rect 16503 36503 16537 36537
rect 16537 36503 16546 36537
rect 16494 36494 16546 36503
rect 16654 36537 16706 36546
rect 16654 36503 16663 36537
rect 16663 36503 16697 36537
rect 16697 36503 16706 36537
rect 16654 36494 16706 36503
rect 16814 36537 16866 36546
rect 16814 36503 16823 36537
rect 16823 36503 16857 36537
rect 16857 36503 16866 36537
rect 16814 36494 16866 36503
rect 16974 36537 17026 36546
rect 16974 36503 16983 36537
rect 16983 36503 17017 36537
rect 17017 36503 17026 36537
rect 16974 36494 17026 36503
rect 17134 36537 17186 36546
rect 17134 36503 17143 36537
rect 17143 36503 17177 36537
rect 17177 36503 17186 36537
rect 17134 36494 17186 36503
rect 17294 36537 17346 36546
rect 17294 36503 17303 36537
rect 17303 36503 17337 36537
rect 17337 36503 17346 36537
rect 17294 36494 17346 36503
rect 17454 36537 17506 36546
rect 17454 36503 17463 36537
rect 17463 36503 17497 36537
rect 17497 36503 17506 36537
rect 17454 36494 17506 36503
rect 17614 36537 17666 36546
rect 17614 36503 17623 36537
rect 17623 36503 17657 36537
rect 17657 36503 17666 36537
rect 17614 36494 17666 36503
rect 17774 36537 17826 36546
rect 17774 36503 17783 36537
rect 17783 36503 17817 36537
rect 17817 36503 17826 36537
rect 17774 36494 17826 36503
rect 17934 36537 17986 36546
rect 17934 36503 17943 36537
rect 17943 36503 17977 36537
rect 17977 36503 17986 36537
rect 17934 36494 17986 36503
rect 18094 36537 18146 36546
rect 18094 36503 18103 36537
rect 18103 36503 18137 36537
rect 18137 36503 18146 36537
rect 18094 36494 18146 36503
rect 18254 36537 18306 36546
rect 18254 36503 18263 36537
rect 18263 36503 18297 36537
rect 18297 36503 18306 36537
rect 18254 36494 18306 36503
rect 18414 36537 18466 36546
rect 18414 36503 18423 36537
rect 18423 36503 18457 36537
rect 18457 36503 18466 36537
rect 18414 36494 18466 36503
rect 18574 36537 18626 36546
rect 18574 36503 18583 36537
rect 18583 36503 18617 36537
rect 18617 36503 18626 36537
rect 18574 36494 18626 36503
rect 18734 36537 18786 36546
rect 18734 36503 18743 36537
rect 18743 36503 18777 36537
rect 18777 36503 18786 36537
rect 18734 36494 18786 36503
rect 18894 36537 18946 36546
rect 18894 36503 18903 36537
rect 18903 36503 18937 36537
rect 18937 36503 18946 36537
rect 18894 36494 18946 36503
rect 23134 36537 23186 36546
rect 23134 36503 23143 36537
rect 23143 36503 23177 36537
rect 23177 36503 23186 36537
rect 23134 36494 23186 36503
rect 23294 36537 23346 36546
rect 23294 36503 23303 36537
rect 23303 36503 23337 36537
rect 23337 36503 23346 36537
rect 23294 36494 23346 36503
rect 23454 36537 23506 36546
rect 23454 36503 23463 36537
rect 23463 36503 23497 36537
rect 23497 36503 23506 36537
rect 23454 36494 23506 36503
rect 23614 36537 23666 36546
rect 23614 36503 23623 36537
rect 23623 36503 23657 36537
rect 23657 36503 23666 36537
rect 23614 36494 23666 36503
rect 23774 36537 23826 36546
rect 23774 36503 23783 36537
rect 23783 36503 23817 36537
rect 23817 36503 23826 36537
rect 23774 36494 23826 36503
rect 23934 36537 23986 36546
rect 23934 36503 23943 36537
rect 23943 36503 23977 36537
rect 23977 36503 23986 36537
rect 23934 36494 23986 36503
rect 24094 36537 24146 36546
rect 24094 36503 24103 36537
rect 24103 36503 24137 36537
rect 24137 36503 24146 36537
rect 24094 36494 24146 36503
rect 24254 36537 24306 36546
rect 24254 36503 24263 36537
rect 24263 36503 24297 36537
rect 24297 36503 24306 36537
rect 24254 36494 24306 36503
rect 24414 36537 24466 36546
rect 24414 36503 24423 36537
rect 24423 36503 24457 36537
rect 24457 36503 24466 36537
rect 24414 36494 24466 36503
rect 24574 36537 24626 36546
rect 24574 36503 24583 36537
rect 24583 36503 24617 36537
rect 24617 36503 24626 36537
rect 24574 36494 24626 36503
rect 24734 36537 24786 36546
rect 24734 36503 24743 36537
rect 24743 36503 24777 36537
rect 24777 36503 24786 36537
rect 24734 36494 24786 36503
rect 24894 36537 24946 36546
rect 24894 36503 24903 36537
rect 24903 36503 24937 36537
rect 24937 36503 24946 36537
rect 24894 36494 24946 36503
rect 25054 36537 25106 36546
rect 25054 36503 25063 36537
rect 25063 36503 25097 36537
rect 25097 36503 25106 36537
rect 25054 36494 25106 36503
rect 25214 36537 25266 36546
rect 25214 36503 25223 36537
rect 25223 36503 25257 36537
rect 25257 36503 25266 36537
rect 25214 36494 25266 36503
rect 25374 36537 25426 36546
rect 25374 36503 25383 36537
rect 25383 36503 25417 36537
rect 25417 36503 25426 36537
rect 25374 36494 25426 36503
rect 25534 36537 25586 36546
rect 25534 36503 25543 36537
rect 25543 36503 25577 36537
rect 25577 36503 25586 36537
rect 25534 36494 25586 36503
rect 25694 36537 25746 36546
rect 25694 36503 25703 36537
rect 25703 36503 25737 36537
rect 25737 36503 25746 36537
rect 25694 36494 25746 36503
rect 25854 36537 25906 36546
rect 25854 36503 25863 36537
rect 25863 36503 25897 36537
rect 25897 36503 25906 36537
rect 25854 36494 25906 36503
rect 26014 36537 26066 36546
rect 26014 36503 26023 36537
rect 26023 36503 26057 36537
rect 26057 36503 26066 36537
rect 26014 36494 26066 36503
rect 26174 36537 26226 36546
rect 26174 36503 26183 36537
rect 26183 36503 26217 36537
rect 26217 36503 26226 36537
rect 26174 36494 26226 36503
rect 26334 36537 26386 36546
rect 26334 36503 26343 36537
rect 26343 36503 26377 36537
rect 26377 36503 26386 36537
rect 26334 36494 26386 36503
rect 26494 36537 26546 36546
rect 26494 36503 26503 36537
rect 26503 36503 26537 36537
rect 26537 36503 26546 36537
rect 26494 36494 26546 36503
rect 26654 36537 26706 36546
rect 26654 36503 26663 36537
rect 26663 36503 26697 36537
rect 26697 36503 26706 36537
rect 26654 36494 26706 36503
rect 26814 36537 26866 36546
rect 26814 36503 26823 36537
rect 26823 36503 26857 36537
rect 26857 36503 26866 36537
rect 26814 36494 26866 36503
rect 26974 36537 27026 36546
rect 26974 36503 26983 36537
rect 26983 36503 27017 36537
rect 27017 36503 27026 36537
rect 26974 36494 27026 36503
rect 27134 36537 27186 36546
rect 27134 36503 27143 36537
rect 27143 36503 27177 36537
rect 27177 36503 27186 36537
rect 27134 36494 27186 36503
rect 27294 36537 27346 36546
rect 27294 36503 27303 36537
rect 27303 36503 27337 36537
rect 27337 36503 27346 36537
rect 27294 36494 27346 36503
rect 27454 36537 27506 36546
rect 27454 36503 27463 36537
rect 27463 36503 27497 36537
rect 27497 36503 27506 36537
rect 27454 36494 27506 36503
rect 27614 36537 27666 36546
rect 27614 36503 27623 36537
rect 27623 36503 27657 36537
rect 27657 36503 27666 36537
rect 27614 36494 27666 36503
rect 27774 36537 27826 36546
rect 27774 36503 27783 36537
rect 27783 36503 27817 36537
rect 27817 36503 27826 36537
rect 27774 36494 27826 36503
rect 27934 36537 27986 36546
rect 27934 36503 27943 36537
rect 27943 36503 27977 36537
rect 27977 36503 27986 36537
rect 27934 36494 27986 36503
rect 28094 36537 28146 36546
rect 28094 36503 28103 36537
rect 28103 36503 28137 36537
rect 28137 36503 28146 36537
rect 28094 36494 28146 36503
rect 28254 36537 28306 36546
rect 28254 36503 28263 36537
rect 28263 36503 28297 36537
rect 28297 36503 28306 36537
rect 28254 36494 28306 36503
rect 28414 36537 28466 36546
rect 28414 36503 28423 36537
rect 28423 36503 28457 36537
rect 28457 36503 28466 36537
rect 28414 36494 28466 36503
rect 28574 36537 28626 36546
rect 28574 36503 28583 36537
rect 28583 36503 28617 36537
rect 28617 36503 28626 36537
rect 28574 36494 28626 36503
rect 28734 36537 28786 36546
rect 28734 36503 28743 36537
rect 28743 36503 28777 36537
rect 28777 36503 28786 36537
rect 28734 36494 28786 36503
rect 28894 36537 28946 36546
rect 28894 36503 28903 36537
rect 28903 36503 28937 36537
rect 28937 36503 28946 36537
rect 28894 36494 28946 36503
rect 29054 36537 29106 36546
rect 29054 36503 29063 36537
rect 29063 36503 29097 36537
rect 29097 36503 29106 36537
rect 29054 36494 29106 36503
rect 29214 36537 29266 36546
rect 29214 36503 29223 36537
rect 29223 36503 29257 36537
rect 29257 36503 29266 36537
rect 29214 36494 29266 36503
rect 29374 36537 29426 36546
rect 29374 36503 29383 36537
rect 29383 36503 29417 36537
rect 29417 36503 29426 36537
rect 29374 36494 29426 36503
rect 33534 36537 33586 36546
rect 33534 36503 33543 36537
rect 33543 36503 33577 36537
rect 33577 36503 33586 36537
rect 33534 36494 33586 36503
rect 33694 36537 33746 36546
rect 33694 36503 33703 36537
rect 33703 36503 33737 36537
rect 33737 36503 33746 36537
rect 33694 36494 33746 36503
rect 33854 36537 33906 36546
rect 33854 36503 33863 36537
rect 33863 36503 33897 36537
rect 33897 36503 33906 36537
rect 33854 36494 33906 36503
rect 34014 36537 34066 36546
rect 34014 36503 34023 36537
rect 34023 36503 34057 36537
rect 34057 36503 34066 36537
rect 34014 36494 34066 36503
rect 34174 36537 34226 36546
rect 34174 36503 34183 36537
rect 34183 36503 34217 36537
rect 34217 36503 34226 36537
rect 34174 36494 34226 36503
rect 34334 36537 34386 36546
rect 34334 36503 34343 36537
rect 34343 36503 34377 36537
rect 34377 36503 34386 36537
rect 34334 36494 34386 36503
rect 34494 36537 34546 36546
rect 34494 36503 34503 36537
rect 34503 36503 34537 36537
rect 34537 36503 34546 36537
rect 34494 36494 34546 36503
rect 34654 36537 34706 36546
rect 34654 36503 34663 36537
rect 34663 36503 34697 36537
rect 34697 36503 34706 36537
rect 34654 36494 34706 36503
rect 34814 36537 34866 36546
rect 34814 36503 34823 36537
rect 34823 36503 34857 36537
rect 34857 36503 34866 36537
rect 34814 36494 34866 36503
rect 34974 36537 35026 36546
rect 34974 36503 34983 36537
rect 34983 36503 35017 36537
rect 35017 36503 35026 36537
rect 34974 36494 35026 36503
rect 35134 36537 35186 36546
rect 35134 36503 35143 36537
rect 35143 36503 35177 36537
rect 35177 36503 35186 36537
rect 35134 36494 35186 36503
rect 35294 36537 35346 36546
rect 35294 36503 35303 36537
rect 35303 36503 35337 36537
rect 35337 36503 35346 36537
rect 35294 36494 35346 36503
rect 35454 36537 35506 36546
rect 35454 36503 35463 36537
rect 35463 36503 35497 36537
rect 35497 36503 35506 36537
rect 35454 36494 35506 36503
rect 35614 36537 35666 36546
rect 35614 36503 35623 36537
rect 35623 36503 35657 36537
rect 35657 36503 35666 36537
rect 35614 36494 35666 36503
rect 35774 36537 35826 36546
rect 35774 36503 35783 36537
rect 35783 36503 35817 36537
rect 35817 36503 35826 36537
rect 35774 36494 35826 36503
rect 35934 36537 35986 36546
rect 35934 36503 35943 36537
rect 35943 36503 35977 36537
rect 35977 36503 35986 36537
rect 35934 36494 35986 36503
rect 36094 36537 36146 36546
rect 36094 36503 36103 36537
rect 36103 36503 36137 36537
rect 36137 36503 36146 36537
rect 36094 36494 36146 36503
rect 36254 36537 36306 36546
rect 36254 36503 36263 36537
rect 36263 36503 36297 36537
rect 36297 36503 36306 36537
rect 36254 36494 36306 36503
rect 36414 36537 36466 36546
rect 36414 36503 36423 36537
rect 36423 36503 36457 36537
rect 36457 36503 36466 36537
rect 36414 36494 36466 36503
rect 36574 36537 36626 36546
rect 36574 36503 36583 36537
rect 36583 36503 36617 36537
rect 36617 36503 36626 36537
rect 36574 36494 36626 36503
rect 36734 36537 36786 36546
rect 36734 36503 36743 36537
rect 36743 36503 36777 36537
rect 36777 36503 36786 36537
rect 36734 36494 36786 36503
rect 36894 36537 36946 36546
rect 36894 36503 36903 36537
rect 36903 36503 36937 36537
rect 36937 36503 36946 36537
rect 36894 36494 36946 36503
rect 37054 36537 37106 36546
rect 37054 36503 37063 36537
rect 37063 36503 37097 36537
rect 37097 36503 37106 36537
rect 37054 36494 37106 36503
rect 37214 36537 37266 36546
rect 37214 36503 37223 36537
rect 37223 36503 37257 36537
rect 37257 36503 37266 36537
rect 37214 36494 37266 36503
rect 37374 36537 37426 36546
rect 37374 36503 37383 36537
rect 37383 36503 37417 36537
rect 37417 36503 37426 36537
rect 37374 36494 37426 36503
rect 37534 36537 37586 36546
rect 37534 36503 37543 36537
rect 37543 36503 37577 36537
rect 37577 36503 37586 36537
rect 37534 36494 37586 36503
rect 37694 36537 37746 36546
rect 37694 36503 37703 36537
rect 37703 36503 37737 36537
rect 37737 36503 37746 36537
rect 37694 36494 37746 36503
rect 37854 36537 37906 36546
rect 37854 36503 37863 36537
rect 37863 36503 37897 36537
rect 37897 36503 37906 36537
rect 37854 36494 37906 36503
rect 38014 36537 38066 36546
rect 38014 36503 38023 36537
rect 38023 36503 38057 36537
rect 38057 36503 38066 36537
rect 38014 36494 38066 36503
rect 38174 36537 38226 36546
rect 38174 36503 38183 36537
rect 38183 36503 38217 36537
rect 38217 36503 38226 36537
rect 38174 36494 38226 36503
rect 38334 36537 38386 36546
rect 38334 36503 38343 36537
rect 38343 36503 38377 36537
rect 38377 36503 38386 36537
rect 38334 36494 38386 36503
rect 38494 36537 38546 36546
rect 38494 36503 38503 36537
rect 38503 36503 38537 36537
rect 38537 36503 38546 36537
rect 38494 36494 38546 36503
rect 38654 36537 38706 36546
rect 38654 36503 38663 36537
rect 38663 36503 38697 36537
rect 38697 36503 38706 36537
rect 38654 36494 38706 36503
rect 38814 36537 38866 36546
rect 38814 36503 38823 36537
rect 38823 36503 38857 36537
rect 38857 36503 38866 36537
rect 38814 36494 38866 36503
rect 38974 36537 39026 36546
rect 38974 36503 38983 36537
rect 38983 36503 39017 36537
rect 39017 36503 39026 36537
rect 38974 36494 39026 36503
rect 39134 36537 39186 36546
rect 39134 36503 39143 36537
rect 39143 36503 39177 36537
rect 39177 36503 39186 36537
rect 39134 36494 39186 36503
rect 39294 36537 39346 36546
rect 39294 36503 39303 36537
rect 39303 36503 39337 36537
rect 39337 36503 39346 36537
rect 39294 36494 39346 36503
rect 39454 36537 39506 36546
rect 39454 36503 39463 36537
rect 39463 36503 39497 36537
rect 39497 36503 39506 36537
rect 39454 36494 39506 36503
rect 39614 36537 39666 36546
rect 39614 36503 39623 36537
rect 39623 36503 39657 36537
rect 39657 36503 39666 36537
rect 39614 36494 39666 36503
rect 39774 36537 39826 36546
rect 39774 36503 39783 36537
rect 39783 36503 39817 36537
rect 39817 36503 39826 36537
rect 39774 36494 39826 36503
rect 39934 36537 39986 36546
rect 39934 36503 39943 36537
rect 39943 36503 39977 36537
rect 39977 36503 39986 36537
rect 39934 36494 39986 36503
rect 40094 36537 40146 36546
rect 40094 36503 40103 36537
rect 40103 36503 40137 36537
rect 40137 36503 40146 36537
rect 40094 36494 40146 36503
rect 40254 36537 40306 36546
rect 40254 36503 40263 36537
rect 40263 36503 40297 36537
rect 40297 36503 40306 36537
rect 40254 36494 40306 36503
rect 40414 36537 40466 36546
rect 40414 36503 40423 36537
rect 40423 36503 40457 36537
rect 40457 36503 40466 36537
rect 40414 36494 40466 36503
rect 40574 36537 40626 36546
rect 40574 36503 40583 36537
rect 40583 36503 40617 36537
rect 40617 36503 40626 36537
rect 40574 36494 40626 36503
rect 40734 36537 40786 36546
rect 40734 36503 40743 36537
rect 40743 36503 40777 36537
rect 40777 36503 40786 36537
rect 40734 36494 40786 36503
rect 40894 36537 40946 36546
rect 40894 36503 40903 36537
rect 40903 36503 40937 36537
rect 40937 36503 40946 36537
rect 40894 36494 40946 36503
rect 41054 36537 41106 36546
rect 41054 36503 41063 36537
rect 41063 36503 41097 36537
rect 41097 36503 41106 36537
rect 41054 36494 41106 36503
rect 41214 36537 41266 36546
rect 41214 36503 41223 36537
rect 41223 36503 41257 36537
rect 41257 36503 41266 36537
rect 41214 36494 41266 36503
rect 41374 36537 41426 36546
rect 41374 36503 41383 36537
rect 41383 36503 41417 36537
rect 41417 36503 41426 36537
rect 41374 36494 41426 36503
rect 41534 36537 41586 36546
rect 41534 36503 41543 36537
rect 41543 36503 41577 36537
rect 41577 36503 41586 36537
rect 41534 36494 41586 36503
rect 41694 36537 41746 36546
rect 41694 36503 41703 36537
rect 41703 36503 41737 36537
rect 41737 36503 41746 36537
rect 41694 36494 41746 36503
rect 41854 36537 41906 36546
rect 41854 36503 41863 36537
rect 41863 36503 41897 36537
rect 41897 36503 41906 36537
rect 41854 36494 41906 36503
rect 14 36377 66 36386
rect 14 36343 23 36377
rect 23 36343 57 36377
rect 57 36343 66 36377
rect 14 36334 66 36343
rect 174 36377 226 36386
rect 174 36343 183 36377
rect 183 36343 217 36377
rect 217 36343 226 36377
rect 174 36334 226 36343
rect 334 36377 386 36386
rect 334 36343 343 36377
rect 343 36343 377 36377
rect 377 36343 386 36377
rect 334 36334 386 36343
rect 494 36377 546 36386
rect 494 36343 503 36377
rect 503 36343 537 36377
rect 537 36343 546 36377
rect 494 36334 546 36343
rect 654 36377 706 36386
rect 654 36343 663 36377
rect 663 36343 697 36377
rect 697 36343 706 36377
rect 654 36334 706 36343
rect 814 36377 866 36386
rect 814 36343 823 36377
rect 823 36343 857 36377
rect 857 36343 866 36377
rect 814 36334 866 36343
rect 974 36377 1026 36386
rect 974 36343 983 36377
rect 983 36343 1017 36377
rect 1017 36343 1026 36377
rect 974 36334 1026 36343
rect 1134 36377 1186 36386
rect 1134 36343 1143 36377
rect 1143 36343 1177 36377
rect 1177 36343 1186 36377
rect 1134 36334 1186 36343
rect 1294 36377 1346 36386
rect 1294 36343 1303 36377
rect 1303 36343 1337 36377
rect 1337 36343 1346 36377
rect 1294 36334 1346 36343
rect 1454 36377 1506 36386
rect 1454 36343 1463 36377
rect 1463 36343 1497 36377
rect 1497 36343 1506 36377
rect 1454 36334 1506 36343
rect 1614 36377 1666 36386
rect 1614 36343 1623 36377
rect 1623 36343 1657 36377
rect 1657 36343 1666 36377
rect 1614 36334 1666 36343
rect 1774 36377 1826 36386
rect 1774 36343 1783 36377
rect 1783 36343 1817 36377
rect 1817 36343 1826 36377
rect 1774 36334 1826 36343
rect 1934 36377 1986 36386
rect 1934 36343 1943 36377
rect 1943 36343 1977 36377
rect 1977 36343 1986 36377
rect 1934 36334 1986 36343
rect 2094 36377 2146 36386
rect 2094 36343 2103 36377
rect 2103 36343 2137 36377
rect 2137 36343 2146 36377
rect 2094 36334 2146 36343
rect 2254 36377 2306 36386
rect 2254 36343 2263 36377
rect 2263 36343 2297 36377
rect 2297 36343 2306 36377
rect 2254 36334 2306 36343
rect 2414 36377 2466 36386
rect 2414 36343 2423 36377
rect 2423 36343 2457 36377
rect 2457 36343 2466 36377
rect 2414 36334 2466 36343
rect 2574 36377 2626 36386
rect 2574 36343 2583 36377
rect 2583 36343 2617 36377
rect 2617 36343 2626 36377
rect 2574 36334 2626 36343
rect 2734 36377 2786 36386
rect 2734 36343 2743 36377
rect 2743 36343 2777 36377
rect 2777 36343 2786 36377
rect 2734 36334 2786 36343
rect 2894 36377 2946 36386
rect 2894 36343 2903 36377
rect 2903 36343 2937 36377
rect 2937 36343 2946 36377
rect 2894 36334 2946 36343
rect 3054 36377 3106 36386
rect 3054 36343 3063 36377
rect 3063 36343 3097 36377
rect 3097 36343 3106 36377
rect 3054 36334 3106 36343
rect 3214 36377 3266 36386
rect 3214 36343 3223 36377
rect 3223 36343 3257 36377
rect 3257 36343 3266 36377
rect 3214 36334 3266 36343
rect 3374 36377 3426 36386
rect 3374 36343 3383 36377
rect 3383 36343 3417 36377
rect 3417 36343 3426 36377
rect 3374 36334 3426 36343
rect 3534 36377 3586 36386
rect 3534 36343 3543 36377
rect 3543 36343 3577 36377
rect 3577 36343 3586 36377
rect 3534 36334 3586 36343
rect 3694 36377 3746 36386
rect 3694 36343 3703 36377
rect 3703 36343 3737 36377
rect 3737 36343 3746 36377
rect 3694 36334 3746 36343
rect 3854 36377 3906 36386
rect 3854 36343 3863 36377
rect 3863 36343 3897 36377
rect 3897 36343 3906 36377
rect 3854 36334 3906 36343
rect 4014 36377 4066 36386
rect 4014 36343 4023 36377
rect 4023 36343 4057 36377
rect 4057 36343 4066 36377
rect 4014 36334 4066 36343
rect 4174 36377 4226 36386
rect 4174 36343 4183 36377
rect 4183 36343 4217 36377
rect 4217 36343 4226 36377
rect 4174 36334 4226 36343
rect 4334 36377 4386 36386
rect 4334 36343 4343 36377
rect 4343 36343 4377 36377
rect 4377 36343 4386 36377
rect 4334 36334 4386 36343
rect 4494 36377 4546 36386
rect 4494 36343 4503 36377
rect 4503 36343 4537 36377
rect 4537 36343 4546 36377
rect 4494 36334 4546 36343
rect 4654 36377 4706 36386
rect 4654 36343 4663 36377
rect 4663 36343 4697 36377
rect 4697 36343 4706 36377
rect 4654 36334 4706 36343
rect 4814 36377 4866 36386
rect 4814 36343 4823 36377
rect 4823 36343 4857 36377
rect 4857 36343 4866 36377
rect 4814 36334 4866 36343
rect 4974 36377 5026 36386
rect 4974 36343 4983 36377
rect 4983 36343 5017 36377
rect 5017 36343 5026 36377
rect 4974 36334 5026 36343
rect 5134 36377 5186 36386
rect 5134 36343 5143 36377
rect 5143 36343 5177 36377
rect 5177 36343 5186 36377
rect 5134 36334 5186 36343
rect 5294 36377 5346 36386
rect 5294 36343 5303 36377
rect 5303 36343 5337 36377
rect 5337 36343 5346 36377
rect 5294 36334 5346 36343
rect 5454 36377 5506 36386
rect 5454 36343 5463 36377
rect 5463 36343 5497 36377
rect 5497 36343 5506 36377
rect 5454 36334 5506 36343
rect 5614 36377 5666 36386
rect 5614 36343 5623 36377
rect 5623 36343 5657 36377
rect 5657 36343 5666 36377
rect 5614 36334 5666 36343
rect 5774 36377 5826 36386
rect 5774 36343 5783 36377
rect 5783 36343 5817 36377
rect 5817 36343 5826 36377
rect 5774 36334 5826 36343
rect 5934 36377 5986 36386
rect 5934 36343 5943 36377
rect 5943 36343 5977 36377
rect 5977 36343 5986 36377
rect 5934 36334 5986 36343
rect 6094 36377 6146 36386
rect 6094 36343 6103 36377
rect 6103 36343 6137 36377
rect 6137 36343 6146 36377
rect 6094 36334 6146 36343
rect 6254 36377 6306 36386
rect 6254 36343 6263 36377
rect 6263 36343 6297 36377
rect 6297 36343 6306 36377
rect 6254 36334 6306 36343
rect 6414 36377 6466 36386
rect 6414 36343 6423 36377
rect 6423 36343 6457 36377
rect 6457 36343 6466 36377
rect 6414 36334 6466 36343
rect 6574 36377 6626 36386
rect 6574 36343 6583 36377
rect 6583 36343 6617 36377
rect 6617 36343 6626 36377
rect 6574 36334 6626 36343
rect 6734 36377 6786 36386
rect 6734 36343 6743 36377
rect 6743 36343 6777 36377
rect 6777 36343 6786 36377
rect 6734 36334 6786 36343
rect 6894 36377 6946 36386
rect 6894 36343 6903 36377
rect 6903 36343 6937 36377
rect 6937 36343 6946 36377
rect 6894 36334 6946 36343
rect 7054 36377 7106 36386
rect 7054 36343 7063 36377
rect 7063 36343 7097 36377
rect 7097 36343 7106 36377
rect 7054 36334 7106 36343
rect 7214 36377 7266 36386
rect 7214 36343 7223 36377
rect 7223 36343 7257 36377
rect 7257 36343 7266 36377
rect 7214 36334 7266 36343
rect 7374 36377 7426 36386
rect 7374 36343 7383 36377
rect 7383 36343 7417 36377
rect 7417 36343 7426 36377
rect 7374 36334 7426 36343
rect 7534 36377 7586 36386
rect 7534 36343 7543 36377
rect 7543 36343 7577 36377
rect 7577 36343 7586 36377
rect 7534 36334 7586 36343
rect 7694 36377 7746 36386
rect 7694 36343 7703 36377
rect 7703 36343 7737 36377
rect 7737 36343 7746 36377
rect 7694 36334 7746 36343
rect 7854 36377 7906 36386
rect 7854 36343 7863 36377
rect 7863 36343 7897 36377
rect 7897 36343 7906 36377
rect 7854 36334 7906 36343
rect 8014 36377 8066 36386
rect 8014 36343 8023 36377
rect 8023 36343 8057 36377
rect 8057 36343 8066 36377
rect 8014 36334 8066 36343
rect 8174 36377 8226 36386
rect 8174 36343 8183 36377
rect 8183 36343 8217 36377
rect 8217 36343 8226 36377
rect 8174 36334 8226 36343
rect 8334 36377 8386 36386
rect 8334 36343 8343 36377
rect 8343 36343 8377 36377
rect 8377 36343 8386 36377
rect 8334 36334 8386 36343
rect 12494 36377 12546 36386
rect 12494 36343 12503 36377
rect 12503 36343 12537 36377
rect 12537 36343 12546 36377
rect 12494 36334 12546 36343
rect 12654 36377 12706 36386
rect 12654 36343 12663 36377
rect 12663 36343 12697 36377
rect 12697 36343 12706 36377
rect 12654 36334 12706 36343
rect 12814 36377 12866 36386
rect 12814 36343 12823 36377
rect 12823 36343 12857 36377
rect 12857 36343 12866 36377
rect 12814 36334 12866 36343
rect 12974 36377 13026 36386
rect 12974 36343 12983 36377
rect 12983 36343 13017 36377
rect 13017 36343 13026 36377
rect 12974 36334 13026 36343
rect 13134 36377 13186 36386
rect 13134 36343 13143 36377
rect 13143 36343 13177 36377
rect 13177 36343 13186 36377
rect 13134 36334 13186 36343
rect 13294 36377 13346 36386
rect 13294 36343 13303 36377
rect 13303 36343 13337 36377
rect 13337 36343 13346 36377
rect 13294 36334 13346 36343
rect 13454 36377 13506 36386
rect 13454 36343 13463 36377
rect 13463 36343 13497 36377
rect 13497 36343 13506 36377
rect 13454 36334 13506 36343
rect 13614 36377 13666 36386
rect 13614 36343 13623 36377
rect 13623 36343 13657 36377
rect 13657 36343 13666 36377
rect 13614 36334 13666 36343
rect 13774 36377 13826 36386
rect 13774 36343 13783 36377
rect 13783 36343 13817 36377
rect 13817 36343 13826 36377
rect 13774 36334 13826 36343
rect 13934 36377 13986 36386
rect 13934 36343 13943 36377
rect 13943 36343 13977 36377
rect 13977 36343 13986 36377
rect 13934 36334 13986 36343
rect 14094 36377 14146 36386
rect 14094 36343 14103 36377
rect 14103 36343 14137 36377
rect 14137 36343 14146 36377
rect 14094 36334 14146 36343
rect 14254 36377 14306 36386
rect 14254 36343 14263 36377
rect 14263 36343 14297 36377
rect 14297 36343 14306 36377
rect 14254 36334 14306 36343
rect 14414 36377 14466 36386
rect 14414 36343 14423 36377
rect 14423 36343 14457 36377
rect 14457 36343 14466 36377
rect 14414 36334 14466 36343
rect 14574 36377 14626 36386
rect 14574 36343 14583 36377
rect 14583 36343 14617 36377
rect 14617 36343 14626 36377
rect 14574 36334 14626 36343
rect 14734 36377 14786 36386
rect 14734 36343 14743 36377
rect 14743 36343 14777 36377
rect 14777 36343 14786 36377
rect 14734 36334 14786 36343
rect 14894 36377 14946 36386
rect 14894 36343 14903 36377
rect 14903 36343 14937 36377
rect 14937 36343 14946 36377
rect 14894 36334 14946 36343
rect 15054 36377 15106 36386
rect 15054 36343 15063 36377
rect 15063 36343 15097 36377
rect 15097 36343 15106 36377
rect 15054 36334 15106 36343
rect 15214 36377 15266 36386
rect 15214 36343 15223 36377
rect 15223 36343 15257 36377
rect 15257 36343 15266 36377
rect 15214 36334 15266 36343
rect 15374 36377 15426 36386
rect 15374 36343 15383 36377
rect 15383 36343 15417 36377
rect 15417 36343 15426 36377
rect 15374 36334 15426 36343
rect 15534 36377 15586 36386
rect 15534 36343 15543 36377
rect 15543 36343 15577 36377
rect 15577 36343 15586 36377
rect 15534 36334 15586 36343
rect 15694 36377 15746 36386
rect 15694 36343 15703 36377
rect 15703 36343 15737 36377
rect 15737 36343 15746 36377
rect 15694 36334 15746 36343
rect 15854 36377 15906 36386
rect 15854 36343 15863 36377
rect 15863 36343 15897 36377
rect 15897 36343 15906 36377
rect 15854 36334 15906 36343
rect 16014 36377 16066 36386
rect 16014 36343 16023 36377
rect 16023 36343 16057 36377
rect 16057 36343 16066 36377
rect 16014 36334 16066 36343
rect 16174 36377 16226 36386
rect 16174 36343 16183 36377
rect 16183 36343 16217 36377
rect 16217 36343 16226 36377
rect 16174 36334 16226 36343
rect 16334 36377 16386 36386
rect 16334 36343 16343 36377
rect 16343 36343 16377 36377
rect 16377 36343 16386 36377
rect 16334 36334 16386 36343
rect 16494 36377 16546 36386
rect 16494 36343 16503 36377
rect 16503 36343 16537 36377
rect 16537 36343 16546 36377
rect 16494 36334 16546 36343
rect 16654 36377 16706 36386
rect 16654 36343 16663 36377
rect 16663 36343 16697 36377
rect 16697 36343 16706 36377
rect 16654 36334 16706 36343
rect 16814 36377 16866 36386
rect 16814 36343 16823 36377
rect 16823 36343 16857 36377
rect 16857 36343 16866 36377
rect 16814 36334 16866 36343
rect 16974 36377 17026 36386
rect 16974 36343 16983 36377
rect 16983 36343 17017 36377
rect 17017 36343 17026 36377
rect 16974 36334 17026 36343
rect 17134 36377 17186 36386
rect 17134 36343 17143 36377
rect 17143 36343 17177 36377
rect 17177 36343 17186 36377
rect 17134 36334 17186 36343
rect 17294 36377 17346 36386
rect 17294 36343 17303 36377
rect 17303 36343 17337 36377
rect 17337 36343 17346 36377
rect 17294 36334 17346 36343
rect 17454 36377 17506 36386
rect 17454 36343 17463 36377
rect 17463 36343 17497 36377
rect 17497 36343 17506 36377
rect 17454 36334 17506 36343
rect 17614 36377 17666 36386
rect 17614 36343 17623 36377
rect 17623 36343 17657 36377
rect 17657 36343 17666 36377
rect 17614 36334 17666 36343
rect 17774 36377 17826 36386
rect 17774 36343 17783 36377
rect 17783 36343 17817 36377
rect 17817 36343 17826 36377
rect 17774 36334 17826 36343
rect 17934 36377 17986 36386
rect 17934 36343 17943 36377
rect 17943 36343 17977 36377
rect 17977 36343 17986 36377
rect 17934 36334 17986 36343
rect 18094 36377 18146 36386
rect 18094 36343 18103 36377
rect 18103 36343 18137 36377
rect 18137 36343 18146 36377
rect 18094 36334 18146 36343
rect 18254 36377 18306 36386
rect 18254 36343 18263 36377
rect 18263 36343 18297 36377
rect 18297 36343 18306 36377
rect 18254 36334 18306 36343
rect 18414 36377 18466 36386
rect 18414 36343 18423 36377
rect 18423 36343 18457 36377
rect 18457 36343 18466 36377
rect 18414 36334 18466 36343
rect 18574 36377 18626 36386
rect 18574 36343 18583 36377
rect 18583 36343 18617 36377
rect 18617 36343 18626 36377
rect 18574 36334 18626 36343
rect 18734 36377 18786 36386
rect 18734 36343 18743 36377
rect 18743 36343 18777 36377
rect 18777 36343 18786 36377
rect 18734 36334 18786 36343
rect 18894 36377 18946 36386
rect 18894 36343 18903 36377
rect 18903 36343 18937 36377
rect 18937 36343 18946 36377
rect 18894 36334 18946 36343
rect 23134 36377 23186 36386
rect 23134 36343 23143 36377
rect 23143 36343 23177 36377
rect 23177 36343 23186 36377
rect 23134 36334 23186 36343
rect 23294 36377 23346 36386
rect 23294 36343 23303 36377
rect 23303 36343 23337 36377
rect 23337 36343 23346 36377
rect 23294 36334 23346 36343
rect 23454 36377 23506 36386
rect 23454 36343 23463 36377
rect 23463 36343 23497 36377
rect 23497 36343 23506 36377
rect 23454 36334 23506 36343
rect 23614 36377 23666 36386
rect 23614 36343 23623 36377
rect 23623 36343 23657 36377
rect 23657 36343 23666 36377
rect 23614 36334 23666 36343
rect 23774 36377 23826 36386
rect 23774 36343 23783 36377
rect 23783 36343 23817 36377
rect 23817 36343 23826 36377
rect 23774 36334 23826 36343
rect 23934 36377 23986 36386
rect 23934 36343 23943 36377
rect 23943 36343 23977 36377
rect 23977 36343 23986 36377
rect 23934 36334 23986 36343
rect 24094 36377 24146 36386
rect 24094 36343 24103 36377
rect 24103 36343 24137 36377
rect 24137 36343 24146 36377
rect 24094 36334 24146 36343
rect 24254 36377 24306 36386
rect 24254 36343 24263 36377
rect 24263 36343 24297 36377
rect 24297 36343 24306 36377
rect 24254 36334 24306 36343
rect 24414 36377 24466 36386
rect 24414 36343 24423 36377
rect 24423 36343 24457 36377
rect 24457 36343 24466 36377
rect 24414 36334 24466 36343
rect 24574 36377 24626 36386
rect 24574 36343 24583 36377
rect 24583 36343 24617 36377
rect 24617 36343 24626 36377
rect 24574 36334 24626 36343
rect 24734 36377 24786 36386
rect 24734 36343 24743 36377
rect 24743 36343 24777 36377
rect 24777 36343 24786 36377
rect 24734 36334 24786 36343
rect 24894 36377 24946 36386
rect 24894 36343 24903 36377
rect 24903 36343 24937 36377
rect 24937 36343 24946 36377
rect 24894 36334 24946 36343
rect 25054 36377 25106 36386
rect 25054 36343 25063 36377
rect 25063 36343 25097 36377
rect 25097 36343 25106 36377
rect 25054 36334 25106 36343
rect 25214 36377 25266 36386
rect 25214 36343 25223 36377
rect 25223 36343 25257 36377
rect 25257 36343 25266 36377
rect 25214 36334 25266 36343
rect 25374 36377 25426 36386
rect 25374 36343 25383 36377
rect 25383 36343 25417 36377
rect 25417 36343 25426 36377
rect 25374 36334 25426 36343
rect 25534 36377 25586 36386
rect 25534 36343 25543 36377
rect 25543 36343 25577 36377
rect 25577 36343 25586 36377
rect 25534 36334 25586 36343
rect 25694 36377 25746 36386
rect 25694 36343 25703 36377
rect 25703 36343 25737 36377
rect 25737 36343 25746 36377
rect 25694 36334 25746 36343
rect 25854 36377 25906 36386
rect 25854 36343 25863 36377
rect 25863 36343 25897 36377
rect 25897 36343 25906 36377
rect 25854 36334 25906 36343
rect 26014 36377 26066 36386
rect 26014 36343 26023 36377
rect 26023 36343 26057 36377
rect 26057 36343 26066 36377
rect 26014 36334 26066 36343
rect 26174 36377 26226 36386
rect 26174 36343 26183 36377
rect 26183 36343 26217 36377
rect 26217 36343 26226 36377
rect 26174 36334 26226 36343
rect 26334 36377 26386 36386
rect 26334 36343 26343 36377
rect 26343 36343 26377 36377
rect 26377 36343 26386 36377
rect 26334 36334 26386 36343
rect 26494 36377 26546 36386
rect 26494 36343 26503 36377
rect 26503 36343 26537 36377
rect 26537 36343 26546 36377
rect 26494 36334 26546 36343
rect 26654 36377 26706 36386
rect 26654 36343 26663 36377
rect 26663 36343 26697 36377
rect 26697 36343 26706 36377
rect 26654 36334 26706 36343
rect 26814 36377 26866 36386
rect 26814 36343 26823 36377
rect 26823 36343 26857 36377
rect 26857 36343 26866 36377
rect 26814 36334 26866 36343
rect 26974 36377 27026 36386
rect 26974 36343 26983 36377
rect 26983 36343 27017 36377
rect 27017 36343 27026 36377
rect 26974 36334 27026 36343
rect 27134 36377 27186 36386
rect 27134 36343 27143 36377
rect 27143 36343 27177 36377
rect 27177 36343 27186 36377
rect 27134 36334 27186 36343
rect 27294 36377 27346 36386
rect 27294 36343 27303 36377
rect 27303 36343 27337 36377
rect 27337 36343 27346 36377
rect 27294 36334 27346 36343
rect 27454 36377 27506 36386
rect 27454 36343 27463 36377
rect 27463 36343 27497 36377
rect 27497 36343 27506 36377
rect 27454 36334 27506 36343
rect 27614 36377 27666 36386
rect 27614 36343 27623 36377
rect 27623 36343 27657 36377
rect 27657 36343 27666 36377
rect 27614 36334 27666 36343
rect 27774 36377 27826 36386
rect 27774 36343 27783 36377
rect 27783 36343 27817 36377
rect 27817 36343 27826 36377
rect 27774 36334 27826 36343
rect 27934 36377 27986 36386
rect 27934 36343 27943 36377
rect 27943 36343 27977 36377
rect 27977 36343 27986 36377
rect 27934 36334 27986 36343
rect 28094 36377 28146 36386
rect 28094 36343 28103 36377
rect 28103 36343 28137 36377
rect 28137 36343 28146 36377
rect 28094 36334 28146 36343
rect 28254 36377 28306 36386
rect 28254 36343 28263 36377
rect 28263 36343 28297 36377
rect 28297 36343 28306 36377
rect 28254 36334 28306 36343
rect 28414 36377 28466 36386
rect 28414 36343 28423 36377
rect 28423 36343 28457 36377
rect 28457 36343 28466 36377
rect 28414 36334 28466 36343
rect 28574 36377 28626 36386
rect 28574 36343 28583 36377
rect 28583 36343 28617 36377
rect 28617 36343 28626 36377
rect 28574 36334 28626 36343
rect 28734 36377 28786 36386
rect 28734 36343 28743 36377
rect 28743 36343 28777 36377
rect 28777 36343 28786 36377
rect 28734 36334 28786 36343
rect 28894 36377 28946 36386
rect 28894 36343 28903 36377
rect 28903 36343 28937 36377
rect 28937 36343 28946 36377
rect 28894 36334 28946 36343
rect 29054 36377 29106 36386
rect 29054 36343 29063 36377
rect 29063 36343 29097 36377
rect 29097 36343 29106 36377
rect 29054 36334 29106 36343
rect 29214 36377 29266 36386
rect 29214 36343 29223 36377
rect 29223 36343 29257 36377
rect 29257 36343 29266 36377
rect 29214 36334 29266 36343
rect 29374 36377 29426 36386
rect 29374 36343 29383 36377
rect 29383 36343 29417 36377
rect 29417 36343 29426 36377
rect 29374 36334 29426 36343
rect 33534 36377 33586 36386
rect 33534 36343 33543 36377
rect 33543 36343 33577 36377
rect 33577 36343 33586 36377
rect 33534 36334 33586 36343
rect 33694 36377 33746 36386
rect 33694 36343 33703 36377
rect 33703 36343 33737 36377
rect 33737 36343 33746 36377
rect 33694 36334 33746 36343
rect 33854 36377 33906 36386
rect 33854 36343 33863 36377
rect 33863 36343 33897 36377
rect 33897 36343 33906 36377
rect 33854 36334 33906 36343
rect 34014 36377 34066 36386
rect 34014 36343 34023 36377
rect 34023 36343 34057 36377
rect 34057 36343 34066 36377
rect 34014 36334 34066 36343
rect 34174 36377 34226 36386
rect 34174 36343 34183 36377
rect 34183 36343 34217 36377
rect 34217 36343 34226 36377
rect 34174 36334 34226 36343
rect 34334 36377 34386 36386
rect 34334 36343 34343 36377
rect 34343 36343 34377 36377
rect 34377 36343 34386 36377
rect 34334 36334 34386 36343
rect 34494 36377 34546 36386
rect 34494 36343 34503 36377
rect 34503 36343 34537 36377
rect 34537 36343 34546 36377
rect 34494 36334 34546 36343
rect 34654 36377 34706 36386
rect 34654 36343 34663 36377
rect 34663 36343 34697 36377
rect 34697 36343 34706 36377
rect 34654 36334 34706 36343
rect 34814 36377 34866 36386
rect 34814 36343 34823 36377
rect 34823 36343 34857 36377
rect 34857 36343 34866 36377
rect 34814 36334 34866 36343
rect 34974 36377 35026 36386
rect 34974 36343 34983 36377
rect 34983 36343 35017 36377
rect 35017 36343 35026 36377
rect 34974 36334 35026 36343
rect 35134 36377 35186 36386
rect 35134 36343 35143 36377
rect 35143 36343 35177 36377
rect 35177 36343 35186 36377
rect 35134 36334 35186 36343
rect 35294 36377 35346 36386
rect 35294 36343 35303 36377
rect 35303 36343 35337 36377
rect 35337 36343 35346 36377
rect 35294 36334 35346 36343
rect 35454 36377 35506 36386
rect 35454 36343 35463 36377
rect 35463 36343 35497 36377
rect 35497 36343 35506 36377
rect 35454 36334 35506 36343
rect 35614 36377 35666 36386
rect 35614 36343 35623 36377
rect 35623 36343 35657 36377
rect 35657 36343 35666 36377
rect 35614 36334 35666 36343
rect 35774 36377 35826 36386
rect 35774 36343 35783 36377
rect 35783 36343 35817 36377
rect 35817 36343 35826 36377
rect 35774 36334 35826 36343
rect 35934 36377 35986 36386
rect 35934 36343 35943 36377
rect 35943 36343 35977 36377
rect 35977 36343 35986 36377
rect 35934 36334 35986 36343
rect 36094 36377 36146 36386
rect 36094 36343 36103 36377
rect 36103 36343 36137 36377
rect 36137 36343 36146 36377
rect 36094 36334 36146 36343
rect 36254 36377 36306 36386
rect 36254 36343 36263 36377
rect 36263 36343 36297 36377
rect 36297 36343 36306 36377
rect 36254 36334 36306 36343
rect 36414 36377 36466 36386
rect 36414 36343 36423 36377
rect 36423 36343 36457 36377
rect 36457 36343 36466 36377
rect 36414 36334 36466 36343
rect 36574 36377 36626 36386
rect 36574 36343 36583 36377
rect 36583 36343 36617 36377
rect 36617 36343 36626 36377
rect 36574 36334 36626 36343
rect 36734 36377 36786 36386
rect 36734 36343 36743 36377
rect 36743 36343 36777 36377
rect 36777 36343 36786 36377
rect 36734 36334 36786 36343
rect 36894 36377 36946 36386
rect 36894 36343 36903 36377
rect 36903 36343 36937 36377
rect 36937 36343 36946 36377
rect 36894 36334 36946 36343
rect 37054 36377 37106 36386
rect 37054 36343 37063 36377
rect 37063 36343 37097 36377
rect 37097 36343 37106 36377
rect 37054 36334 37106 36343
rect 37214 36377 37266 36386
rect 37214 36343 37223 36377
rect 37223 36343 37257 36377
rect 37257 36343 37266 36377
rect 37214 36334 37266 36343
rect 37374 36377 37426 36386
rect 37374 36343 37383 36377
rect 37383 36343 37417 36377
rect 37417 36343 37426 36377
rect 37374 36334 37426 36343
rect 37534 36377 37586 36386
rect 37534 36343 37543 36377
rect 37543 36343 37577 36377
rect 37577 36343 37586 36377
rect 37534 36334 37586 36343
rect 37694 36377 37746 36386
rect 37694 36343 37703 36377
rect 37703 36343 37737 36377
rect 37737 36343 37746 36377
rect 37694 36334 37746 36343
rect 37854 36377 37906 36386
rect 37854 36343 37863 36377
rect 37863 36343 37897 36377
rect 37897 36343 37906 36377
rect 37854 36334 37906 36343
rect 38014 36377 38066 36386
rect 38014 36343 38023 36377
rect 38023 36343 38057 36377
rect 38057 36343 38066 36377
rect 38014 36334 38066 36343
rect 38174 36377 38226 36386
rect 38174 36343 38183 36377
rect 38183 36343 38217 36377
rect 38217 36343 38226 36377
rect 38174 36334 38226 36343
rect 38334 36377 38386 36386
rect 38334 36343 38343 36377
rect 38343 36343 38377 36377
rect 38377 36343 38386 36377
rect 38334 36334 38386 36343
rect 38494 36377 38546 36386
rect 38494 36343 38503 36377
rect 38503 36343 38537 36377
rect 38537 36343 38546 36377
rect 38494 36334 38546 36343
rect 38654 36377 38706 36386
rect 38654 36343 38663 36377
rect 38663 36343 38697 36377
rect 38697 36343 38706 36377
rect 38654 36334 38706 36343
rect 38814 36377 38866 36386
rect 38814 36343 38823 36377
rect 38823 36343 38857 36377
rect 38857 36343 38866 36377
rect 38814 36334 38866 36343
rect 38974 36377 39026 36386
rect 38974 36343 38983 36377
rect 38983 36343 39017 36377
rect 39017 36343 39026 36377
rect 38974 36334 39026 36343
rect 39134 36377 39186 36386
rect 39134 36343 39143 36377
rect 39143 36343 39177 36377
rect 39177 36343 39186 36377
rect 39134 36334 39186 36343
rect 39294 36377 39346 36386
rect 39294 36343 39303 36377
rect 39303 36343 39337 36377
rect 39337 36343 39346 36377
rect 39294 36334 39346 36343
rect 39454 36377 39506 36386
rect 39454 36343 39463 36377
rect 39463 36343 39497 36377
rect 39497 36343 39506 36377
rect 39454 36334 39506 36343
rect 39614 36377 39666 36386
rect 39614 36343 39623 36377
rect 39623 36343 39657 36377
rect 39657 36343 39666 36377
rect 39614 36334 39666 36343
rect 39774 36377 39826 36386
rect 39774 36343 39783 36377
rect 39783 36343 39817 36377
rect 39817 36343 39826 36377
rect 39774 36334 39826 36343
rect 39934 36377 39986 36386
rect 39934 36343 39943 36377
rect 39943 36343 39977 36377
rect 39977 36343 39986 36377
rect 39934 36334 39986 36343
rect 40094 36377 40146 36386
rect 40094 36343 40103 36377
rect 40103 36343 40137 36377
rect 40137 36343 40146 36377
rect 40094 36334 40146 36343
rect 40254 36377 40306 36386
rect 40254 36343 40263 36377
rect 40263 36343 40297 36377
rect 40297 36343 40306 36377
rect 40254 36334 40306 36343
rect 40414 36377 40466 36386
rect 40414 36343 40423 36377
rect 40423 36343 40457 36377
rect 40457 36343 40466 36377
rect 40414 36334 40466 36343
rect 40574 36377 40626 36386
rect 40574 36343 40583 36377
rect 40583 36343 40617 36377
rect 40617 36343 40626 36377
rect 40574 36334 40626 36343
rect 40734 36377 40786 36386
rect 40734 36343 40743 36377
rect 40743 36343 40777 36377
rect 40777 36343 40786 36377
rect 40734 36334 40786 36343
rect 40894 36377 40946 36386
rect 40894 36343 40903 36377
rect 40903 36343 40937 36377
rect 40937 36343 40946 36377
rect 40894 36334 40946 36343
rect 41054 36377 41106 36386
rect 41054 36343 41063 36377
rect 41063 36343 41097 36377
rect 41097 36343 41106 36377
rect 41054 36334 41106 36343
rect 41214 36377 41266 36386
rect 41214 36343 41223 36377
rect 41223 36343 41257 36377
rect 41257 36343 41266 36377
rect 41214 36334 41266 36343
rect 41374 36377 41426 36386
rect 41374 36343 41383 36377
rect 41383 36343 41417 36377
rect 41417 36343 41426 36377
rect 41374 36334 41426 36343
rect 41534 36377 41586 36386
rect 41534 36343 41543 36377
rect 41543 36343 41577 36377
rect 41577 36343 41586 36377
rect 41534 36334 41586 36343
rect 41694 36377 41746 36386
rect 41694 36343 41703 36377
rect 41703 36343 41737 36377
rect 41737 36343 41746 36377
rect 41694 36334 41746 36343
rect 41854 36377 41906 36386
rect 41854 36343 41863 36377
rect 41863 36343 41897 36377
rect 41897 36343 41906 36377
rect 41854 36334 41906 36343
rect 14 36057 66 36066
rect 14 36023 23 36057
rect 23 36023 57 36057
rect 57 36023 66 36057
rect 14 36014 66 36023
rect 174 36057 226 36066
rect 174 36023 183 36057
rect 183 36023 217 36057
rect 217 36023 226 36057
rect 174 36014 226 36023
rect 334 36057 386 36066
rect 334 36023 343 36057
rect 343 36023 377 36057
rect 377 36023 386 36057
rect 334 36014 386 36023
rect 494 36057 546 36066
rect 494 36023 503 36057
rect 503 36023 537 36057
rect 537 36023 546 36057
rect 494 36014 546 36023
rect 654 36057 706 36066
rect 654 36023 663 36057
rect 663 36023 697 36057
rect 697 36023 706 36057
rect 654 36014 706 36023
rect 814 36057 866 36066
rect 814 36023 823 36057
rect 823 36023 857 36057
rect 857 36023 866 36057
rect 814 36014 866 36023
rect 974 36057 1026 36066
rect 974 36023 983 36057
rect 983 36023 1017 36057
rect 1017 36023 1026 36057
rect 974 36014 1026 36023
rect 1134 36057 1186 36066
rect 1134 36023 1143 36057
rect 1143 36023 1177 36057
rect 1177 36023 1186 36057
rect 1134 36014 1186 36023
rect 1294 36057 1346 36066
rect 1294 36023 1303 36057
rect 1303 36023 1337 36057
rect 1337 36023 1346 36057
rect 1294 36014 1346 36023
rect 1454 36057 1506 36066
rect 1454 36023 1463 36057
rect 1463 36023 1497 36057
rect 1497 36023 1506 36057
rect 1454 36014 1506 36023
rect 1614 36057 1666 36066
rect 1614 36023 1623 36057
rect 1623 36023 1657 36057
rect 1657 36023 1666 36057
rect 1614 36014 1666 36023
rect 1774 36057 1826 36066
rect 1774 36023 1783 36057
rect 1783 36023 1817 36057
rect 1817 36023 1826 36057
rect 1774 36014 1826 36023
rect 1934 36057 1986 36066
rect 1934 36023 1943 36057
rect 1943 36023 1977 36057
rect 1977 36023 1986 36057
rect 1934 36014 1986 36023
rect 2094 36057 2146 36066
rect 2094 36023 2103 36057
rect 2103 36023 2137 36057
rect 2137 36023 2146 36057
rect 2094 36014 2146 36023
rect 2254 36057 2306 36066
rect 2254 36023 2263 36057
rect 2263 36023 2297 36057
rect 2297 36023 2306 36057
rect 2254 36014 2306 36023
rect 2414 36057 2466 36066
rect 2414 36023 2423 36057
rect 2423 36023 2457 36057
rect 2457 36023 2466 36057
rect 2414 36014 2466 36023
rect 2574 36057 2626 36066
rect 2574 36023 2583 36057
rect 2583 36023 2617 36057
rect 2617 36023 2626 36057
rect 2574 36014 2626 36023
rect 2734 36057 2786 36066
rect 2734 36023 2743 36057
rect 2743 36023 2777 36057
rect 2777 36023 2786 36057
rect 2734 36014 2786 36023
rect 2894 36057 2946 36066
rect 2894 36023 2903 36057
rect 2903 36023 2937 36057
rect 2937 36023 2946 36057
rect 2894 36014 2946 36023
rect 3054 36057 3106 36066
rect 3054 36023 3063 36057
rect 3063 36023 3097 36057
rect 3097 36023 3106 36057
rect 3054 36014 3106 36023
rect 3214 36057 3266 36066
rect 3214 36023 3223 36057
rect 3223 36023 3257 36057
rect 3257 36023 3266 36057
rect 3214 36014 3266 36023
rect 3374 36057 3426 36066
rect 3374 36023 3383 36057
rect 3383 36023 3417 36057
rect 3417 36023 3426 36057
rect 3374 36014 3426 36023
rect 3534 36057 3586 36066
rect 3534 36023 3543 36057
rect 3543 36023 3577 36057
rect 3577 36023 3586 36057
rect 3534 36014 3586 36023
rect 3694 36057 3746 36066
rect 3694 36023 3703 36057
rect 3703 36023 3737 36057
rect 3737 36023 3746 36057
rect 3694 36014 3746 36023
rect 3854 36057 3906 36066
rect 3854 36023 3863 36057
rect 3863 36023 3897 36057
rect 3897 36023 3906 36057
rect 3854 36014 3906 36023
rect 4014 36057 4066 36066
rect 4014 36023 4023 36057
rect 4023 36023 4057 36057
rect 4057 36023 4066 36057
rect 4014 36014 4066 36023
rect 4174 36057 4226 36066
rect 4174 36023 4183 36057
rect 4183 36023 4217 36057
rect 4217 36023 4226 36057
rect 4174 36014 4226 36023
rect 4334 36057 4386 36066
rect 4334 36023 4343 36057
rect 4343 36023 4377 36057
rect 4377 36023 4386 36057
rect 4334 36014 4386 36023
rect 4494 36057 4546 36066
rect 4494 36023 4503 36057
rect 4503 36023 4537 36057
rect 4537 36023 4546 36057
rect 4494 36014 4546 36023
rect 4654 36057 4706 36066
rect 4654 36023 4663 36057
rect 4663 36023 4697 36057
rect 4697 36023 4706 36057
rect 4654 36014 4706 36023
rect 4814 36057 4866 36066
rect 4814 36023 4823 36057
rect 4823 36023 4857 36057
rect 4857 36023 4866 36057
rect 4814 36014 4866 36023
rect 4974 36057 5026 36066
rect 4974 36023 4983 36057
rect 4983 36023 5017 36057
rect 5017 36023 5026 36057
rect 4974 36014 5026 36023
rect 5134 36057 5186 36066
rect 5134 36023 5143 36057
rect 5143 36023 5177 36057
rect 5177 36023 5186 36057
rect 5134 36014 5186 36023
rect 5294 36057 5346 36066
rect 5294 36023 5303 36057
rect 5303 36023 5337 36057
rect 5337 36023 5346 36057
rect 5294 36014 5346 36023
rect 5454 36057 5506 36066
rect 5454 36023 5463 36057
rect 5463 36023 5497 36057
rect 5497 36023 5506 36057
rect 5454 36014 5506 36023
rect 5614 36057 5666 36066
rect 5614 36023 5623 36057
rect 5623 36023 5657 36057
rect 5657 36023 5666 36057
rect 5614 36014 5666 36023
rect 5774 36057 5826 36066
rect 5774 36023 5783 36057
rect 5783 36023 5817 36057
rect 5817 36023 5826 36057
rect 5774 36014 5826 36023
rect 5934 36057 5986 36066
rect 5934 36023 5943 36057
rect 5943 36023 5977 36057
rect 5977 36023 5986 36057
rect 5934 36014 5986 36023
rect 6094 36057 6146 36066
rect 6094 36023 6103 36057
rect 6103 36023 6137 36057
rect 6137 36023 6146 36057
rect 6094 36014 6146 36023
rect 6254 36057 6306 36066
rect 6254 36023 6263 36057
rect 6263 36023 6297 36057
rect 6297 36023 6306 36057
rect 6254 36014 6306 36023
rect 6414 36057 6466 36066
rect 6414 36023 6423 36057
rect 6423 36023 6457 36057
rect 6457 36023 6466 36057
rect 6414 36014 6466 36023
rect 6574 36057 6626 36066
rect 6574 36023 6583 36057
rect 6583 36023 6617 36057
rect 6617 36023 6626 36057
rect 6574 36014 6626 36023
rect 6734 36057 6786 36066
rect 6734 36023 6743 36057
rect 6743 36023 6777 36057
rect 6777 36023 6786 36057
rect 6734 36014 6786 36023
rect 6894 36057 6946 36066
rect 6894 36023 6903 36057
rect 6903 36023 6937 36057
rect 6937 36023 6946 36057
rect 6894 36014 6946 36023
rect 7054 36057 7106 36066
rect 7054 36023 7063 36057
rect 7063 36023 7097 36057
rect 7097 36023 7106 36057
rect 7054 36014 7106 36023
rect 7214 36057 7266 36066
rect 7214 36023 7223 36057
rect 7223 36023 7257 36057
rect 7257 36023 7266 36057
rect 7214 36014 7266 36023
rect 7374 36057 7426 36066
rect 7374 36023 7383 36057
rect 7383 36023 7417 36057
rect 7417 36023 7426 36057
rect 7374 36014 7426 36023
rect 7534 36057 7586 36066
rect 7534 36023 7543 36057
rect 7543 36023 7577 36057
rect 7577 36023 7586 36057
rect 7534 36014 7586 36023
rect 7694 36057 7746 36066
rect 7694 36023 7703 36057
rect 7703 36023 7737 36057
rect 7737 36023 7746 36057
rect 7694 36014 7746 36023
rect 7854 36057 7906 36066
rect 7854 36023 7863 36057
rect 7863 36023 7897 36057
rect 7897 36023 7906 36057
rect 7854 36014 7906 36023
rect 8014 36057 8066 36066
rect 8014 36023 8023 36057
rect 8023 36023 8057 36057
rect 8057 36023 8066 36057
rect 8014 36014 8066 36023
rect 8174 36057 8226 36066
rect 8174 36023 8183 36057
rect 8183 36023 8217 36057
rect 8217 36023 8226 36057
rect 8174 36014 8226 36023
rect 8334 36057 8386 36066
rect 8334 36023 8343 36057
rect 8343 36023 8377 36057
rect 8377 36023 8386 36057
rect 8334 36014 8386 36023
rect 12494 36057 12546 36066
rect 12494 36023 12503 36057
rect 12503 36023 12537 36057
rect 12537 36023 12546 36057
rect 12494 36014 12546 36023
rect 12654 36057 12706 36066
rect 12654 36023 12663 36057
rect 12663 36023 12697 36057
rect 12697 36023 12706 36057
rect 12654 36014 12706 36023
rect 12814 36057 12866 36066
rect 12814 36023 12823 36057
rect 12823 36023 12857 36057
rect 12857 36023 12866 36057
rect 12814 36014 12866 36023
rect 12974 36057 13026 36066
rect 12974 36023 12983 36057
rect 12983 36023 13017 36057
rect 13017 36023 13026 36057
rect 12974 36014 13026 36023
rect 13134 36057 13186 36066
rect 13134 36023 13143 36057
rect 13143 36023 13177 36057
rect 13177 36023 13186 36057
rect 13134 36014 13186 36023
rect 13294 36057 13346 36066
rect 13294 36023 13303 36057
rect 13303 36023 13337 36057
rect 13337 36023 13346 36057
rect 13294 36014 13346 36023
rect 13454 36057 13506 36066
rect 13454 36023 13463 36057
rect 13463 36023 13497 36057
rect 13497 36023 13506 36057
rect 13454 36014 13506 36023
rect 13614 36057 13666 36066
rect 13614 36023 13623 36057
rect 13623 36023 13657 36057
rect 13657 36023 13666 36057
rect 13614 36014 13666 36023
rect 13774 36057 13826 36066
rect 13774 36023 13783 36057
rect 13783 36023 13817 36057
rect 13817 36023 13826 36057
rect 13774 36014 13826 36023
rect 13934 36057 13986 36066
rect 13934 36023 13943 36057
rect 13943 36023 13977 36057
rect 13977 36023 13986 36057
rect 13934 36014 13986 36023
rect 14094 36057 14146 36066
rect 14094 36023 14103 36057
rect 14103 36023 14137 36057
rect 14137 36023 14146 36057
rect 14094 36014 14146 36023
rect 14254 36057 14306 36066
rect 14254 36023 14263 36057
rect 14263 36023 14297 36057
rect 14297 36023 14306 36057
rect 14254 36014 14306 36023
rect 14414 36057 14466 36066
rect 14414 36023 14423 36057
rect 14423 36023 14457 36057
rect 14457 36023 14466 36057
rect 14414 36014 14466 36023
rect 14574 36057 14626 36066
rect 14574 36023 14583 36057
rect 14583 36023 14617 36057
rect 14617 36023 14626 36057
rect 14574 36014 14626 36023
rect 14734 36057 14786 36066
rect 14734 36023 14743 36057
rect 14743 36023 14777 36057
rect 14777 36023 14786 36057
rect 14734 36014 14786 36023
rect 14894 36057 14946 36066
rect 14894 36023 14903 36057
rect 14903 36023 14937 36057
rect 14937 36023 14946 36057
rect 14894 36014 14946 36023
rect 15054 36057 15106 36066
rect 15054 36023 15063 36057
rect 15063 36023 15097 36057
rect 15097 36023 15106 36057
rect 15054 36014 15106 36023
rect 15214 36057 15266 36066
rect 15214 36023 15223 36057
rect 15223 36023 15257 36057
rect 15257 36023 15266 36057
rect 15214 36014 15266 36023
rect 15374 36057 15426 36066
rect 15374 36023 15383 36057
rect 15383 36023 15417 36057
rect 15417 36023 15426 36057
rect 15374 36014 15426 36023
rect 15534 36057 15586 36066
rect 15534 36023 15543 36057
rect 15543 36023 15577 36057
rect 15577 36023 15586 36057
rect 15534 36014 15586 36023
rect 15694 36057 15746 36066
rect 15694 36023 15703 36057
rect 15703 36023 15737 36057
rect 15737 36023 15746 36057
rect 15694 36014 15746 36023
rect 15854 36057 15906 36066
rect 15854 36023 15863 36057
rect 15863 36023 15897 36057
rect 15897 36023 15906 36057
rect 15854 36014 15906 36023
rect 16014 36057 16066 36066
rect 16014 36023 16023 36057
rect 16023 36023 16057 36057
rect 16057 36023 16066 36057
rect 16014 36014 16066 36023
rect 16174 36057 16226 36066
rect 16174 36023 16183 36057
rect 16183 36023 16217 36057
rect 16217 36023 16226 36057
rect 16174 36014 16226 36023
rect 16334 36057 16386 36066
rect 16334 36023 16343 36057
rect 16343 36023 16377 36057
rect 16377 36023 16386 36057
rect 16334 36014 16386 36023
rect 16494 36057 16546 36066
rect 16494 36023 16503 36057
rect 16503 36023 16537 36057
rect 16537 36023 16546 36057
rect 16494 36014 16546 36023
rect 16654 36057 16706 36066
rect 16654 36023 16663 36057
rect 16663 36023 16697 36057
rect 16697 36023 16706 36057
rect 16654 36014 16706 36023
rect 16814 36057 16866 36066
rect 16814 36023 16823 36057
rect 16823 36023 16857 36057
rect 16857 36023 16866 36057
rect 16814 36014 16866 36023
rect 16974 36057 17026 36066
rect 16974 36023 16983 36057
rect 16983 36023 17017 36057
rect 17017 36023 17026 36057
rect 16974 36014 17026 36023
rect 17134 36057 17186 36066
rect 17134 36023 17143 36057
rect 17143 36023 17177 36057
rect 17177 36023 17186 36057
rect 17134 36014 17186 36023
rect 17294 36057 17346 36066
rect 17294 36023 17303 36057
rect 17303 36023 17337 36057
rect 17337 36023 17346 36057
rect 17294 36014 17346 36023
rect 17454 36057 17506 36066
rect 17454 36023 17463 36057
rect 17463 36023 17497 36057
rect 17497 36023 17506 36057
rect 17454 36014 17506 36023
rect 17614 36057 17666 36066
rect 17614 36023 17623 36057
rect 17623 36023 17657 36057
rect 17657 36023 17666 36057
rect 17614 36014 17666 36023
rect 17774 36057 17826 36066
rect 17774 36023 17783 36057
rect 17783 36023 17817 36057
rect 17817 36023 17826 36057
rect 17774 36014 17826 36023
rect 17934 36057 17986 36066
rect 17934 36023 17943 36057
rect 17943 36023 17977 36057
rect 17977 36023 17986 36057
rect 17934 36014 17986 36023
rect 18094 36057 18146 36066
rect 18094 36023 18103 36057
rect 18103 36023 18137 36057
rect 18137 36023 18146 36057
rect 18094 36014 18146 36023
rect 18254 36057 18306 36066
rect 18254 36023 18263 36057
rect 18263 36023 18297 36057
rect 18297 36023 18306 36057
rect 18254 36014 18306 36023
rect 18414 36057 18466 36066
rect 18414 36023 18423 36057
rect 18423 36023 18457 36057
rect 18457 36023 18466 36057
rect 18414 36014 18466 36023
rect 18574 36057 18626 36066
rect 18574 36023 18583 36057
rect 18583 36023 18617 36057
rect 18617 36023 18626 36057
rect 18574 36014 18626 36023
rect 18734 36057 18786 36066
rect 18734 36023 18743 36057
rect 18743 36023 18777 36057
rect 18777 36023 18786 36057
rect 18734 36014 18786 36023
rect 18894 36057 18946 36066
rect 18894 36023 18903 36057
rect 18903 36023 18937 36057
rect 18937 36023 18946 36057
rect 18894 36014 18946 36023
rect 23134 36057 23186 36066
rect 23134 36023 23143 36057
rect 23143 36023 23177 36057
rect 23177 36023 23186 36057
rect 23134 36014 23186 36023
rect 23294 36057 23346 36066
rect 23294 36023 23303 36057
rect 23303 36023 23337 36057
rect 23337 36023 23346 36057
rect 23294 36014 23346 36023
rect 23454 36057 23506 36066
rect 23454 36023 23463 36057
rect 23463 36023 23497 36057
rect 23497 36023 23506 36057
rect 23454 36014 23506 36023
rect 23614 36057 23666 36066
rect 23614 36023 23623 36057
rect 23623 36023 23657 36057
rect 23657 36023 23666 36057
rect 23614 36014 23666 36023
rect 23774 36057 23826 36066
rect 23774 36023 23783 36057
rect 23783 36023 23817 36057
rect 23817 36023 23826 36057
rect 23774 36014 23826 36023
rect 23934 36057 23986 36066
rect 23934 36023 23943 36057
rect 23943 36023 23977 36057
rect 23977 36023 23986 36057
rect 23934 36014 23986 36023
rect 24094 36057 24146 36066
rect 24094 36023 24103 36057
rect 24103 36023 24137 36057
rect 24137 36023 24146 36057
rect 24094 36014 24146 36023
rect 24254 36057 24306 36066
rect 24254 36023 24263 36057
rect 24263 36023 24297 36057
rect 24297 36023 24306 36057
rect 24254 36014 24306 36023
rect 24414 36057 24466 36066
rect 24414 36023 24423 36057
rect 24423 36023 24457 36057
rect 24457 36023 24466 36057
rect 24414 36014 24466 36023
rect 24574 36057 24626 36066
rect 24574 36023 24583 36057
rect 24583 36023 24617 36057
rect 24617 36023 24626 36057
rect 24574 36014 24626 36023
rect 24734 36057 24786 36066
rect 24734 36023 24743 36057
rect 24743 36023 24777 36057
rect 24777 36023 24786 36057
rect 24734 36014 24786 36023
rect 24894 36057 24946 36066
rect 24894 36023 24903 36057
rect 24903 36023 24937 36057
rect 24937 36023 24946 36057
rect 24894 36014 24946 36023
rect 25054 36057 25106 36066
rect 25054 36023 25063 36057
rect 25063 36023 25097 36057
rect 25097 36023 25106 36057
rect 25054 36014 25106 36023
rect 25214 36057 25266 36066
rect 25214 36023 25223 36057
rect 25223 36023 25257 36057
rect 25257 36023 25266 36057
rect 25214 36014 25266 36023
rect 25374 36057 25426 36066
rect 25374 36023 25383 36057
rect 25383 36023 25417 36057
rect 25417 36023 25426 36057
rect 25374 36014 25426 36023
rect 25534 36057 25586 36066
rect 25534 36023 25543 36057
rect 25543 36023 25577 36057
rect 25577 36023 25586 36057
rect 25534 36014 25586 36023
rect 25694 36057 25746 36066
rect 25694 36023 25703 36057
rect 25703 36023 25737 36057
rect 25737 36023 25746 36057
rect 25694 36014 25746 36023
rect 25854 36057 25906 36066
rect 25854 36023 25863 36057
rect 25863 36023 25897 36057
rect 25897 36023 25906 36057
rect 25854 36014 25906 36023
rect 26014 36057 26066 36066
rect 26014 36023 26023 36057
rect 26023 36023 26057 36057
rect 26057 36023 26066 36057
rect 26014 36014 26066 36023
rect 26174 36057 26226 36066
rect 26174 36023 26183 36057
rect 26183 36023 26217 36057
rect 26217 36023 26226 36057
rect 26174 36014 26226 36023
rect 26334 36057 26386 36066
rect 26334 36023 26343 36057
rect 26343 36023 26377 36057
rect 26377 36023 26386 36057
rect 26334 36014 26386 36023
rect 26494 36057 26546 36066
rect 26494 36023 26503 36057
rect 26503 36023 26537 36057
rect 26537 36023 26546 36057
rect 26494 36014 26546 36023
rect 26654 36057 26706 36066
rect 26654 36023 26663 36057
rect 26663 36023 26697 36057
rect 26697 36023 26706 36057
rect 26654 36014 26706 36023
rect 26814 36057 26866 36066
rect 26814 36023 26823 36057
rect 26823 36023 26857 36057
rect 26857 36023 26866 36057
rect 26814 36014 26866 36023
rect 26974 36057 27026 36066
rect 26974 36023 26983 36057
rect 26983 36023 27017 36057
rect 27017 36023 27026 36057
rect 26974 36014 27026 36023
rect 27134 36057 27186 36066
rect 27134 36023 27143 36057
rect 27143 36023 27177 36057
rect 27177 36023 27186 36057
rect 27134 36014 27186 36023
rect 27294 36057 27346 36066
rect 27294 36023 27303 36057
rect 27303 36023 27337 36057
rect 27337 36023 27346 36057
rect 27294 36014 27346 36023
rect 27454 36057 27506 36066
rect 27454 36023 27463 36057
rect 27463 36023 27497 36057
rect 27497 36023 27506 36057
rect 27454 36014 27506 36023
rect 27614 36057 27666 36066
rect 27614 36023 27623 36057
rect 27623 36023 27657 36057
rect 27657 36023 27666 36057
rect 27614 36014 27666 36023
rect 27774 36057 27826 36066
rect 27774 36023 27783 36057
rect 27783 36023 27817 36057
rect 27817 36023 27826 36057
rect 27774 36014 27826 36023
rect 27934 36057 27986 36066
rect 27934 36023 27943 36057
rect 27943 36023 27977 36057
rect 27977 36023 27986 36057
rect 27934 36014 27986 36023
rect 28094 36057 28146 36066
rect 28094 36023 28103 36057
rect 28103 36023 28137 36057
rect 28137 36023 28146 36057
rect 28094 36014 28146 36023
rect 28254 36057 28306 36066
rect 28254 36023 28263 36057
rect 28263 36023 28297 36057
rect 28297 36023 28306 36057
rect 28254 36014 28306 36023
rect 28414 36057 28466 36066
rect 28414 36023 28423 36057
rect 28423 36023 28457 36057
rect 28457 36023 28466 36057
rect 28414 36014 28466 36023
rect 28574 36057 28626 36066
rect 28574 36023 28583 36057
rect 28583 36023 28617 36057
rect 28617 36023 28626 36057
rect 28574 36014 28626 36023
rect 28734 36057 28786 36066
rect 28734 36023 28743 36057
rect 28743 36023 28777 36057
rect 28777 36023 28786 36057
rect 28734 36014 28786 36023
rect 28894 36057 28946 36066
rect 28894 36023 28903 36057
rect 28903 36023 28937 36057
rect 28937 36023 28946 36057
rect 28894 36014 28946 36023
rect 29054 36057 29106 36066
rect 29054 36023 29063 36057
rect 29063 36023 29097 36057
rect 29097 36023 29106 36057
rect 29054 36014 29106 36023
rect 29214 36057 29266 36066
rect 29214 36023 29223 36057
rect 29223 36023 29257 36057
rect 29257 36023 29266 36057
rect 29214 36014 29266 36023
rect 29374 36057 29426 36066
rect 29374 36023 29383 36057
rect 29383 36023 29417 36057
rect 29417 36023 29426 36057
rect 29374 36014 29426 36023
rect 33534 36057 33586 36066
rect 33534 36023 33543 36057
rect 33543 36023 33577 36057
rect 33577 36023 33586 36057
rect 33534 36014 33586 36023
rect 33694 36057 33746 36066
rect 33694 36023 33703 36057
rect 33703 36023 33737 36057
rect 33737 36023 33746 36057
rect 33694 36014 33746 36023
rect 33854 36057 33906 36066
rect 33854 36023 33863 36057
rect 33863 36023 33897 36057
rect 33897 36023 33906 36057
rect 33854 36014 33906 36023
rect 34014 36057 34066 36066
rect 34014 36023 34023 36057
rect 34023 36023 34057 36057
rect 34057 36023 34066 36057
rect 34014 36014 34066 36023
rect 34174 36057 34226 36066
rect 34174 36023 34183 36057
rect 34183 36023 34217 36057
rect 34217 36023 34226 36057
rect 34174 36014 34226 36023
rect 34334 36057 34386 36066
rect 34334 36023 34343 36057
rect 34343 36023 34377 36057
rect 34377 36023 34386 36057
rect 34334 36014 34386 36023
rect 34494 36057 34546 36066
rect 34494 36023 34503 36057
rect 34503 36023 34537 36057
rect 34537 36023 34546 36057
rect 34494 36014 34546 36023
rect 34654 36057 34706 36066
rect 34654 36023 34663 36057
rect 34663 36023 34697 36057
rect 34697 36023 34706 36057
rect 34654 36014 34706 36023
rect 34814 36057 34866 36066
rect 34814 36023 34823 36057
rect 34823 36023 34857 36057
rect 34857 36023 34866 36057
rect 34814 36014 34866 36023
rect 34974 36057 35026 36066
rect 34974 36023 34983 36057
rect 34983 36023 35017 36057
rect 35017 36023 35026 36057
rect 34974 36014 35026 36023
rect 35134 36057 35186 36066
rect 35134 36023 35143 36057
rect 35143 36023 35177 36057
rect 35177 36023 35186 36057
rect 35134 36014 35186 36023
rect 35294 36057 35346 36066
rect 35294 36023 35303 36057
rect 35303 36023 35337 36057
rect 35337 36023 35346 36057
rect 35294 36014 35346 36023
rect 35454 36057 35506 36066
rect 35454 36023 35463 36057
rect 35463 36023 35497 36057
rect 35497 36023 35506 36057
rect 35454 36014 35506 36023
rect 35614 36057 35666 36066
rect 35614 36023 35623 36057
rect 35623 36023 35657 36057
rect 35657 36023 35666 36057
rect 35614 36014 35666 36023
rect 35774 36057 35826 36066
rect 35774 36023 35783 36057
rect 35783 36023 35817 36057
rect 35817 36023 35826 36057
rect 35774 36014 35826 36023
rect 35934 36057 35986 36066
rect 35934 36023 35943 36057
rect 35943 36023 35977 36057
rect 35977 36023 35986 36057
rect 35934 36014 35986 36023
rect 36094 36057 36146 36066
rect 36094 36023 36103 36057
rect 36103 36023 36137 36057
rect 36137 36023 36146 36057
rect 36094 36014 36146 36023
rect 36254 36057 36306 36066
rect 36254 36023 36263 36057
rect 36263 36023 36297 36057
rect 36297 36023 36306 36057
rect 36254 36014 36306 36023
rect 36414 36057 36466 36066
rect 36414 36023 36423 36057
rect 36423 36023 36457 36057
rect 36457 36023 36466 36057
rect 36414 36014 36466 36023
rect 36574 36057 36626 36066
rect 36574 36023 36583 36057
rect 36583 36023 36617 36057
rect 36617 36023 36626 36057
rect 36574 36014 36626 36023
rect 36734 36057 36786 36066
rect 36734 36023 36743 36057
rect 36743 36023 36777 36057
rect 36777 36023 36786 36057
rect 36734 36014 36786 36023
rect 36894 36057 36946 36066
rect 36894 36023 36903 36057
rect 36903 36023 36937 36057
rect 36937 36023 36946 36057
rect 36894 36014 36946 36023
rect 37054 36057 37106 36066
rect 37054 36023 37063 36057
rect 37063 36023 37097 36057
rect 37097 36023 37106 36057
rect 37054 36014 37106 36023
rect 37214 36057 37266 36066
rect 37214 36023 37223 36057
rect 37223 36023 37257 36057
rect 37257 36023 37266 36057
rect 37214 36014 37266 36023
rect 37374 36057 37426 36066
rect 37374 36023 37383 36057
rect 37383 36023 37417 36057
rect 37417 36023 37426 36057
rect 37374 36014 37426 36023
rect 37534 36057 37586 36066
rect 37534 36023 37543 36057
rect 37543 36023 37577 36057
rect 37577 36023 37586 36057
rect 37534 36014 37586 36023
rect 37694 36057 37746 36066
rect 37694 36023 37703 36057
rect 37703 36023 37737 36057
rect 37737 36023 37746 36057
rect 37694 36014 37746 36023
rect 37854 36057 37906 36066
rect 37854 36023 37863 36057
rect 37863 36023 37897 36057
rect 37897 36023 37906 36057
rect 37854 36014 37906 36023
rect 38014 36057 38066 36066
rect 38014 36023 38023 36057
rect 38023 36023 38057 36057
rect 38057 36023 38066 36057
rect 38014 36014 38066 36023
rect 38174 36057 38226 36066
rect 38174 36023 38183 36057
rect 38183 36023 38217 36057
rect 38217 36023 38226 36057
rect 38174 36014 38226 36023
rect 38334 36057 38386 36066
rect 38334 36023 38343 36057
rect 38343 36023 38377 36057
rect 38377 36023 38386 36057
rect 38334 36014 38386 36023
rect 38494 36057 38546 36066
rect 38494 36023 38503 36057
rect 38503 36023 38537 36057
rect 38537 36023 38546 36057
rect 38494 36014 38546 36023
rect 38654 36057 38706 36066
rect 38654 36023 38663 36057
rect 38663 36023 38697 36057
rect 38697 36023 38706 36057
rect 38654 36014 38706 36023
rect 38814 36057 38866 36066
rect 38814 36023 38823 36057
rect 38823 36023 38857 36057
rect 38857 36023 38866 36057
rect 38814 36014 38866 36023
rect 38974 36057 39026 36066
rect 38974 36023 38983 36057
rect 38983 36023 39017 36057
rect 39017 36023 39026 36057
rect 38974 36014 39026 36023
rect 39134 36057 39186 36066
rect 39134 36023 39143 36057
rect 39143 36023 39177 36057
rect 39177 36023 39186 36057
rect 39134 36014 39186 36023
rect 39294 36057 39346 36066
rect 39294 36023 39303 36057
rect 39303 36023 39337 36057
rect 39337 36023 39346 36057
rect 39294 36014 39346 36023
rect 39454 36057 39506 36066
rect 39454 36023 39463 36057
rect 39463 36023 39497 36057
rect 39497 36023 39506 36057
rect 39454 36014 39506 36023
rect 39614 36057 39666 36066
rect 39614 36023 39623 36057
rect 39623 36023 39657 36057
rect 39657 36023 39666 36057
rect 39614 36014 39666 36023
rect 39774 36057 39826 36066
rect 39774 36023 39783 36057
rect 39783 36023 39817 36057
rect 39817 36023 39826 36057
rect 39774 36014 39826 36023
rect 39934 36057 39986 36066
rect 39934 36023 39943 36057
rect 39943 36023 39977 36057
rect 39977 36023 39986 36057
rect 39934 36014 39986 36023
rect 40094 36057 40146 36066
rect 40094 36023 40103 36057
rect 40103 36023 40137 36057
rect 40137 36023 40146 36057
rect 40094 36014 40146 36023
rect 40254 36057 40306 36066
rect 40254 36023 40263 36057
rect 40263 36023 40297 36057
rect 40297 36023 40306 36057
rect 40254 36014 40306 36023
rect 40414 36057 40466 36066
rect 40414 36023 40423 36057
rect 40423 36023 40457 36057
rect 40457 36023 40466 36057
rect 40414 36014 40466 36023
rect 40574 36057 40626 36066
rect 40574 36023 40583 36057
rect 40583 36023 40617 36057
rect 40617 36023 40626 36057
rect 40574 36014 40626 36023
rect 40734 36057 40786 36066
rect 40734 36023 40743 36057
rect 40743 36023 40777 36057
rect 40777 36023 40786 36057
rect 40734 36014 40786 36023
rect 40894 36057 40946 36066
rect 40894 36023 40903 36057
rect 40903 36023 40937 36057
rect 40937 36023 40946 36057
rect 40894 36014 40946 36023
rect 41054 36057 41106 36066
rect 41054 36023 41063 36057
rect 41063 36023 41097 36057
rect 41097 36023 41106 36057
rect 41054 36014 41106 36023
rect 41214 36057 41266 36066
rect 41214 36023 41223 36057
rect 41223 36023 41257 36057
rect 41257 36023 41266 36057
rect 41214 36014 41266 36023
rect 41374 36057 41426 36066
rect 41374 36023 41383 36057
rect 41383 36023 41417 36057
rect 41417 36023 41426 36057
rect 41374 36014 41426 36023
rect 41534 36057 41586 36066
rect 41534 36023 41543 36057
rect 41543 36023 41577 36057
rect 41577 36023 41586 36057
rect 41534 36014 41586 36023
rect 41694 36057 41746 36066
rect 41694 36023 41703 36057
rect 41703 36023 41737 36057
rect 41737 36023 41746 36057
rect 41694 36014 41746 36023
rect 41854 36057 41906 36066
rect 41854 36023 41863 36057
rect 41863 36023 41897 36057
rect 41897 36023 41906 36057
rect 41854 36014 41906 36023
rect 14 35737 66 35746
rect 14 35703 23 35737
rect 23 35703 57 35737
rect 57 35703 66 35737
rect 14 35694 66 35703
rect 174 35737 226 35746
rect 174 35703 183 35737
rect 183 35703 217 35737
rect 217 35703 226 35737
rect 174 35694 226 35703
rect 334 35737 386 35746
rect 334 35703 343 35737
rect 343 35703 377 35737
rect 377 35703 386 35737
rect 334 35694 386 35703
rect 494 35737 546 35746
rect 494 35703 503 35737
rect 503 35703 537 35737
rect 537 35703 546 35737
rect 494 35694 546 35703
rect 654 35737 706 35746
rect 654 35703 663 35737
rect 663 35703 697 35737
rect 697 35703 706 35737
rect 654 35694 706 35703
rect 814 35737 866 35746
rect 814 35703 823 35737
rect 823 35703 857 35737
rect 857 35703 866 35737
rect 814 35694 866 35703
rect 974 35737 1026 35746
rect 974 35703 983 35737
rect 983 35703 1017 35737
rect 1017 35703 1026 35737
rect 974 35694 1026 35703
rect 1134 35737 1186 35746
rect 1134 35703 1143 35737
rect 1143 35703 1177 35737
rect 1177 35703 1186 35737
rect 1134 35694 1186 35703
rect 1294 35737 1346 35746
rect 1294 35703 1303 35737
rect 1303 35703 1337 35737
rect 1337 35703 1346 35737
rect 1294 35694 1346 35703
rect 1454 35737 1506 35746
rect 1454 35703 1463 35737
rect 1463 35703 1497 35737
rect 1497 35703 1506 35737
rect 1454 35694 1506 35703
rect 1614 35737 1666 35746
rect 1614 35703 1623 35737
rect 1623 35703 1657 35737
rect 1657 35703 1666 35737
rect 1614 35694 1666 35703
rect 1774 35737 1826 35746
rect 1774 35703 1783 35737
rect 1783 35703 1817 35737
rect 1817 35703 1826 35737
rect 1774 35694 1826 35703
rect 1934 35737 1986 35746
rect 1934 35703 1943 35737
rect 1943 35703 1977 35737
rect 1977 35703 1986 35737
rect 1934 35694 1986 35703
rect 2094 35737 2146 35746
rect 2094 35703 2103 35737
rect 2103 35703 2137 35737
rect 2137 35703 2146 35737
rect 2094 35694 2146 35703
rect 2254 35737 2306 35746
rect 2254 35703 2263 35737
rect 2263 35703 2297 35737
rect 2297 35703 2306 35737
rect 2254 35694 2306 35703
rect 2414 35737 2466 35746
rect 2414 35703 2423 35737
rect 2423 35703 2457 35737
rect 2457 35703 2466 35737
rect 2414 35694 2466 35703
rect 2574 35737 2626 35746
rect 2574 35703 2583 35737
rect 2583 35703 2617 35737
rect 2617 35703 2626 35737
rect 2574 35694 2626 35703
rect 2734 35737 2786 35746
rect 2734 35703 2743 35737
rect 2743 35703 2777 35737
rect 2777 35703 2786 35737
rect 2734 35694 2786 35703
rect 2894 35737 2946 35746
rect 2894 35703 2903 35737
rect 2903 35703 2937 35737
rect 2937 35703 2946 35737
rect 2894 35694 2946 35703
rect 3054 35737 3106 35746
rect 3054 35703 3063 35737
rect 3063 35703 3097 35737
rect 3097 35703 3106 35737
rect 3054 35694 3106 35703
rect 3214 35737 3266 35746
rect 3214 35703 3223 35737
rect 3223 35703 3257 35737
rect 3257 35703 3266 35737
rect 3214 35694 3266 35703
rect 3374 35737 3426 35746
rect 3374 35703 3383 35737
rect 3383 35703 3417 35737
rect 3417 35703 3426 35737
rect 3374 35694 3426 35703
rect 3534 35737 3586 35746
rect 3534 35703 3543 35737
rect 3543 35703 3577 35737
rect 3577 35703 3586 35737
rect 3534 35694 3586 35703
rect 3694 35737 3746 35746
rect 3694 35703 3703 35737
rect 3703 35703 3737 35737
rect 3737 35703 3746 35737
rect 3694 35694 3746 35703
rect 3854 35737 3906 35746
rect 3854 35703 3863 35737
rect 3863 35703 3897 35737
rect 3897 35703 3906 35737
rect 3854 35694 3906 35703
rect 4014 35737 4066 35746
rect 4014 35703 4023 35737
rect 4023 35703 4057 35737
rect 4057 35703 4066 35737
rect 4014 35694 4066 35703
rect 4174 35737 4226 35746
rect 4174 35703 4183 35737
rect 4183 35703 4217 35737
rect 4217 35703 4226 35737
rect 4174 35694 4226 35703
rect 4334 35737 4386 35746
rect 4334 35703 4343 35737
rect 4343 35703 4377 35737
rect 4377 35703 4386 35737
rect 4334 35694 4386 35703
rect 4494 35737 4546 35746
rect 4494 35703 4503 35737
rect 4503 35703 4537 35737
rect 4537 35703 4546 35737
rect 4494 35694 4546 35703
rect 4654 35737 4706 35746
rect 4654 35703 4663 35737
rect 4663 35703 4697 35737
rect 4697 35703 4706 35737
rect 4654 35694 4706 35703
rect 4814 35737 4866 35746
rect 4814 35703 4823 35737
rect 4823 35703 4857 35737
rect 4857 35703 4866 35737
rect 4814 35694 4866 35703
rect 4974 35737 5026 35746
rect 4974 35703 4983 35737
rect 4983 35703 5017 35737
rect 5017 35703 5026 35737
rect 4974 35694 5026 35703
rect 5134 35737 5186 35746
rect 5134 35703 5143 35737
rect 5143 35703 5177 35737
rect 5177 35703 5186 35737
rect 5134 35694 5186 35703
rect 5294 35737 5346 35746
rect 5294 35703 5303 35737
rect 5303 35703 5337 35737
rect 5337 35703 5346 35737
rect 5294 35694 5346 35703
rect 5454 35737 5506 35746
rect 5454 35703 5463 35737
rect 5463 35703 5497 35737
rect 5497 35703 5506 35737
rect 5454 35694 5506 35703
rect 5614 35737 5666 35746
rect 5614 35703 5623 35737
rect 5623 35703 5657 35737
rect 5657 35703 5666 35737
rect 5614 35694 5666 35703
rect 5774 35737 5826 35746
rect 5774 35703 5783 35737
rect 5783 35703 5817 35737
rect 5817 35703 5826 35737
rect 5774 35694 5826 35703
rect 5934 35737 5986 35746
rect 5934 35703 5943 35737
rect 5943 35703 5977 35737
rect 5977 35703 5986 35737
rect 5934 35694 5986 35703
rect 6094 35737 6146 35746
rect 6094 35703 6103 35737
rect 6103 35703 6137 35737
rect 6137 35703 6146 35737
rect 6094 35694 6146 35703
rect 6254 35737 6306 35746
rect 6254 35703 6263 35737
rect 6263 35703 6297 35737
rect 6297 35703 6306 35737
rect 6254 35694 6306 35703
rect 6414 35737 6466 35746
rect 6414 35703 6423 35737
rect 6423 35703 6457 35737
rect 6457 35703 6466 35737
rect 6414 35694 6466 35703
rect 6574 35737 6626 35746
rect 6574 35703 6583 35737
rect 6583 35703 6617 35737
rect 6617 35703 6626 35737
rect 6574 35694 6626 35703
rect 6734 35737 6786 35746
rect 6734 35703 6743 35737
rect 6743 35703 6777 35737
rect 6777 35703 6786 35737
rect 6734 35694 6786 35703
rect 6894 35737 6946 35746
rect 6894 35703 6903 35737
rect 6903 35703 6937 35737
rect 6937 35703 6946 35737
rect 6894 35694 6946 35703
rect 7054 35737 7106 35746
rect 7054 35703 7063 35737
rect 7063 35703 7097 35737
rect 7097 35703 7106 35737
rect 7054 35694 7106 35703
rect 7214 35737 7266 35746
rect 7214 35703 7223 35737
rect 7223 35703 7257 35737
rect 7257 35703 7266 35737
rect 7214 35694 7266 35703
rect 7374 35737 7426 35746
rect 7374 35703 7383 35737
rect 7383 35703 7417 35737
rect 7417 35703 7426 35737
rect 7374 35694 7426 35703
rect 7534 35737 7586 35746
rect 7534 35703 7543 35737
rect 7543 35703 7577 35737
rect 7577 35703 7586 35737
rect 7534 35694 7586 35703
rect 7694 35737 7746 35746
rect 7694 35703 7703 35737
rect 7703 35703 7737 35737
rect 7737 35703 7746 35737
rect 7694 35694 7746 35703
rect 7854 35737 7906 35746
rect 7854 35703 7863 35737
rect 7863 35703 7897 35737
rect 7897 35703 7906 35737
rect 7854 35694 7906 35703
rect 8014 35737 8066 35746
rect 8014 35703 8023 35737
rect 8023 35703 8057 35737
rect 8057 35703 8066 35737
rect 8014 35694 8066 35703
rect 8174 35737 8226 35746
rect 8174 35703 8183 35737
rect 8183 35703 8217 35737
rect 8217 35703 8226 35737
rect 8174 35694 8226 35703
rect 8334 35737 8386 35746
rect 8334 35703 8343 35737
rect 8343 35703 8377 35737
rect 8377 35703 8386 35737
rect 8334 35694 8386 35703
rect 12494 35737 12546 35746
rect 12494 35703 12503 35737
rect 12503 35703 12537 35737
rect 12537 35703 12546 35737
rect 12494 35694 12546 35703
rect 12654 35737 12706 35746
rect 12654 35703 12663 35737
rect 12663 35703 12697 35737
rect 12697 35703 12706 35737
rect 12654 35694 12706 35703
rect 12814 35737 12866 35746
rect 12814 35703 12823 35737
rect 12823 35703 12857 35737
rect 12857 35703 12866 35737
rect 12814 35694 12866 35703
rect 12974 35737 13026 35746
rect 12974 35703 12983 35737
rect 12983 35703 13017 35737
rect 13017 35703 13026 35737
rect 12974 35694 13026 35703
rect 13134 35737 13186 35746
rect 13134 35703 13143 35737
rect 13143 35703 13177 35737
rect 13177 35703 13186 35737
rect 13134 35694 13186 35703
rect 13294 35737 13346 35746
rect 13294 35703 13303 35737
rect 13303 35703 13337 35737
rect 13337 35703 13346 35737
rect 13294 35694 13346 35703
rect 13454 35737 13506 35746
rect 13454 35703 13463 35737
rect 13463 35703 13497 35737
rect 13497 35703 13506 35737
rect 13454 35694 13506 35703
rect 13614 35737 13666 35746
rect 13614 35703 13623 35737
rect 13623 35703 13657 35737
rect 13657 35703 13666 35737
rect 13614 35694 13666 35703
rect 13774 35737 13826 35746
rect 13774 35703 13783 35737
rect 13783 35703 13817 35737
rect 13817 35703 13826 35737
rect 13774 35694 13826 35703
rect 13934 35737 13986 35746
rect 13934 35703 13943 35737
rect 13943 35703 13977 35737
rect 13977 35703 13986 35737
rect 13934 35694 13986 35703
rect 14094 35737 14146 35746
rect 14094 35703 14103 35737
rect 14103 35703 14137 35737
rect 14137 35703 14146 35737
rect 14094 35694 14146 35703
rect 14254 35737 14306 35746
rect 14254 35703 14263 35737
rect 14263 35703 14297 35737
rect 14297 35703 14306 35737
rect 14254 35694 14306 35703
rect 14414 35737 14466 35746
rect 14414 35703 14423 35737
rect 14423 35703 14457 35737
rect 14457 35703 14466 35737
rect 14414 35694 14466 35703
rect 14574 35737 14626 35746
rect 14574 35703 14583 35737
rect 14583 35703 14617 35737
rect 14617 35703 14626 35737
rect 14574 35694 14626 35703
rect 14734 35737 14786 35746
rect 14734 35703 14743 35737
rect 14743 35703 14777 35737
rect 14777 35703 14786 35737
rect 14734 35694 14786 35703
rect 14894 35737 14946 35746
rect 14894 35703 14903 35737
rect 14903 35703 14937 35737
rect 14937 35703 14946 35737
rect 14894 35694 14946 35703
rect 15054 35737 15106 35746
rect 15054 35703 15063 35737
rect 15063 35703 15097 35737
rect 15097 35703 15106 35737
rect 15054 35694 15106 35703
rect 15214 35737 15266 35746
rect 15214 35703 15223 35737
rect 15223 35703 15257 35737
rect 15257 35703 15266 35737
rect 15214 35694 15266 35703
rect 15374 35737 15426 35746
rect 15374 35703 15383 35737
rect 15383 35703 15417 35737
rect 15417 35703 15426 35737
rect 15374 35694 15426 35703
rect 15534 35737 15586 35746
rect 15534 35703 15543 35737
rect 15543 35703 15577 35737
rect 15577 35703 15586 35737
rect 15534 35694 15586 35703
rect 15694 35737 15746 35746
rect 15694 35703 15703 35737
rect 15703 35703 15737 35737
rect 15737 35703 15746 35737
rect 15694 35694 15746 35703
rect 15854 35737 15906 35746
rect 15854 35703 15863 35737
rect 15863 35703 15897 35737
rect 15897 35703 15906 35737
rect 15854 35694 15906 35703
rect 16014 35737 16066 35746
rect 16014 35703 16023 35737
rect 16023 35703 16057 35737
rect 16057 35703 16066 35737
rect 16014 35694 16066 35703
rect 16174 35737 16226 35746
rect 16174 35703 16183 35737
rect 16183 35703 16217 35737
rect 16217 35703 16226 35737
rect 16174 35694 16226 35703
rect 16334 35737 16386 35746
rect 16334 35703 16343 35737
rect 16343 35703 16377 35737
rect 16377 35703 16386 35737
rect 16334 35694 16386 35703
rect 16494 35737 16546 35746
rect 16494 35703 16503 35737
rect 16503 35703 16537 35737
rect 16537 35703 16546 35737
rect 16494 35694 16546 35703
rect 16654 35737 16706 35746
rect 16654 35703 16663 35737
rect 16663 35703 16697 35737
rect 16697 35703 16706 35737
rect 16654 35694 16706 35703
rect 16814 35737 16866 35746
rect 16814 35703 16823 35737
rect 16823 35703 16857 35737
rect 16857 35703 16866 35737
rect 16814 35694 16866 35703
rect 16974 35737 17026 35746
rect 16974 35703 16983 35737
rect 16983 35703 17017 35737
rect 17017 35703 17026 35737
rect 16974 35694 17026 35703
rect 17134 35737 17186 35746
rect 17134 35703 17143 35737
rect 17143 35703 17177 35737
rect 17177 35703 17186 35737
rect 17134 35694 17186 35703
rect 17294 35737 17346 35746
rect 17294 35703 17303 35737
rect 17303 35703 17337 35737
rect 17337 35703 17346 35737
rect 17294 35694 17346 35703
rect 17454 35737 17506 35746
rect 17454 35703 17463 35737
rect 17463 35703 17497 35737
rect 17497 35703 17506 35737
rect 17454 35694 17506 35703
rect 17614 35737 17666 35746
rect 17614 35703 17623 35737
rect 17623 35703 17657 35737
rect 17657 35703 17666 35737
rect 17614 35694 17666 35703
rect 17774 35737 17826 35746
rect 17774 35703 17783 35737
rect 17783 35703 17817 35737
rect 17817 35703 17826 35737
rect 17774 35694 17826 35703
rect 17934 35737 17986 35746
rect 17934 35703 17943 35737
rect 17943 35703 17977 35737
rect 17977 35703 17986 35737
rect 17934 35694 17986 35703
rect 18094 35737 18146 35746
rect 18094 35703 18103 35737
rect 18103 35703 18137 35737
rect 18137 35703 18146 35737
rect 18094 35694 18146 35703
rect 18254 35737 18306 35746
rect 18254 35703 18263 35737
rect 18263 35703 18297 35737
rect 18297 35703 18306 35737
rect 18254 35694 18306 35703
rect 18414 35737 18466 35746
rect 18414 35703 18423 35737
rect 18423 35703 18457 35737
rect 18457 35703 18466 35737
rect 18414 35694 18466 35703
rect 18574 35737 18626 35746
rect 18574 35703 18583 35737
rect 18583 35703 18617 35737
rect 18617 35703 18626 35737
rect 18574 35694 18626 35703
rect 18734 35737 18786 35746
rect 18734 35703 18743 35737
rect 18743 35703 18777 35737
rect 18777 35703 18786 35737
rect 18734 35694 18786 35703
rect 18894 35737 18946 35746
rect 18894 35703 18903 35737
rect 18903 35703 18937 35737
rect 18937 35703 18946 35737
rect 18894 35694 18946 35703
rect 23134 35737 23186 35746
rect 23134 35703 23143 35737
rect 23143 35703 23177 35737
rect 23177 35703 23186 35737
rect 23134 35694 23186 35703
rect 23294 35737 23346 35746
rect 23294 35703 23303 35737
rect 23303 35703 23337 35737
rect 23337 35703 23346 35737
rect 23294 35694 23346 35703
rect 23454 35737 23506 35746
rect 23454 35703 23463 35737
rect 23463 35703 23497 35737
rect 23497 35703 23506 35737
rect 23454 35694 23506 35703
rect 23614 35737 23666 35746
rect 23614 35703 23623 35737
rect 23623 35703 23657 35737
rect 23657 35703 23666 35737
rect 23614 35694 23666 35703
rect 23774 35737 23826 35746
rect 23774 35703 23783 35737
rect 23783 35703 23817 35737
rect 23817 35703 23826 35737
rect 23774 35694 23826 35703
rect 23934 35737 23986 35746
rect 23934 35703 23943 35737
rect 23943 35703 23977 35737
rect 23977 35703 23986 35737
rect 23934 35694 23986 35703
rect 24094 35737 24146 35746
rect 24094 35703 24103 35737
rect 24103 35703 24137 35737
rect 24137 35703 24146 35737
rect 24094 35694 24146 35703
rect 24254 35737 24306 35746
rect 24254 35703 24263 35737
rect 24263 35703 24297 35737
rect 24297 35703 24306 35737
rect 24254 35694 24306 35703
rect 24414 35737 24466 35746
rect 24414 35703 24423 35737
rect 24423 35703 24457 35737
rect 24457 35703 24466 35737
rect 24414 35694 24466 35703
rect 24574 35737 24626 35746
rect 24574 35703 24583 35737
rect 24583 35703 24617 35737
rect 24617 35703 24626 35737
rect 24574 35694 24626 35703
rect 24734 35737 24786 35746
rect 24734 35703 24743 35737
rect 24743 35703 24777 35737
rect 24777 35703 24786 35737
rect 24734 35694 24786 35703
rect 24894 35737 24946 35746
rect 24894 35703 24903 35737
rect 24903 35703 24937 35737
rect 24937 35703 24946 35737
rect 24894 35694 24946 35703
rect 25054 35737 25106 35746
rect 25054 35703 25063 35737
rect 25063 35703 25097 35737
rect 25097 35703 25106 35737
rect 25054 35694 25106 35703
rect 25214 35737 25266 35746
rect 25214 35703 25223 35737
rect 25223 35703 25257 35737
rect 25257 35703 25266 35737
rect 25214 35694 25266 35703
rect 25374 35737 25426 35746
rect 25374 35703 25383 35737
rect 25383 35703 25417 35737
rect 25417 35703 25426 35737
rect 25374 35694 25426 35703
rect 25534 35737 25586 35746
rect 25534 35703 25543 35737
rect 25543 35703 25577 35737
rect 25577 35703 25586 35737
rect 25534 35694 25586 35703
rect 25694 35737 25746 35746
rect 25694 35703 25703 35737
rect 25703 35703 25737 35737
rect 25737 35703 25746 35737
rect 25694 35694 25746 35703
rect 25854 35737 25906 35746
rect 25854 35703 25863 35737
rect 25863 35703 25897 35737
rect 25897 35703 25906 35737
rect 25854 35694 25906 35703
rect 26014 35737 26066 35746
rect 26014 35703 26023 35737
rect 26023 35703 26057 35737
rect 26057 35703 26066 35737
rect 26014 35694 26066 35703
rect 26174 35737 26226 35746
rect 26174 35703 26183 35737
rect 26183 35703 26217 35737
rect 26217 35703 26226 35737
rect 26174 35694 26226 35703
rect 26334 35737 26386 35746
rect 26334 35703 26343 35737
rect 26343 35703 26377 35737
rect 26377 35703 26386 35737
rect 26334 35694 26386 35703
rect 26494 35737 26546 35746
rect 26494 35703 26503 35737
rect 26503 35703 26537 35737
rect 26537 35703 26546 35737
rect 26494 35694 26546 35703
rect 26654 35737 26706 35746
rect 26654 35703 26663 35737
rect 26663 35703 26697 35737
rect 26697 35703 26706 35737
rect 26654 35694 26706 35703
rect 26814 35737 26866 35746
rect 26814 35703 26823 35737
rect 26823 35703 26857 35737
rect 26857 35703 26866 35737
rect 26814 35694 26866 35703
rect 26974 35737 27026 35746
rect 26974 35703 26983 35737
rect 26983 35703 27017 35737
rect 27017 35703 27026 35737
rect 26974 35694 27026 35703
rect 27134 35737 27186 35746
rect 27134 35703 27143 35737
rect 27143 35703 27177 35737
rect 27177 35703 27186 35737
rect 27134 35694 27186 35703
rect 27294 35737 27346 35746
rect 27294 35703 27303 35737
rect 27303 35703 27337 35737
rect 27337 35703 27346 35737
rect 27294 35694 27346 35703
rect 27454 35737 27506 35746
rect 27454 35703 27463 35737
rect 27463 35703 27497 35737
rect 27497 35703 27506 35737
rect 27454 35694 27506 35703
rect 27614 35737 27666 35746
rect 27614 35703 27623 35737
rect 27623 35703 27657 35737
rect 27657 35703 27666 35737
rect 27614 35694 27666 35703
rect 27774 35737 27826 35746
rect 27774 35703 27783 35737
rect 27783 35703 27817 35737
rect 27817 35703 27826 35737
rect 27774 35694 27826 35703
rect 27934 35737 27986 35746
rect 27934 35703 27943 35737
rect 27943 35703 27977 35737
rect 27977 35703 27986 35737
rect 27934 35694 27986 35703
rect 28094 35737 28146 35746
rect 28094 35703 28103 35737
rect 28103 35703 28137 35737
rect 28137 35703 28146 35737
rect 28094 35694 28146 35703
rect 28254 35737 28306 35746
rect 28254 35703 28263 35737
rect 28263 35703 28297 35737
rect 28297 35703 28306 35737
rect 28254 35694 28306 35703
rect 28414 35737 28466 35746
rect 28414 35703 28423 35737
rect 28423 35703 28457 35737
rect 28457 35703 28466 35737
rect 28414 35694 28466 35703
rect 28574 35737 28626 35746
rect 28574 35703 28583 35737
rect 28583 35703 28617 35737
rect 28617 35703 28626 35737
rect 28574 35694 28626 35703
rect 28734 35737 28786 35746
rect 28734 35703 28743 35737
rect 28743 35703 28777 35737
rect 28777 35703 28786 35737
rect 28734 35694 28786 35703
rect 28894 35737 28946 35746
rect 28894 35703 28903 35737
rect 28903 35703 28937 35737
rect 28937 35703 28946 35737
rect 28894 35694 28946 35703
rect 29054 35737 29106 35746
rect 29054 35703 29063 35737
rect 29063 35703 29097 35737
rect 29097 35703 29106 35737
rect 29054 35694 29106 35703
rect 29214 35737 29266 35746
rect 29214 35703 29223 35737
rect 29223 35703 29257 35737
rect 29257 35703 29266 35737
rect 29214 35694 29266 35703
rect 29374 35737 29426 35746
rect 29374 35703 29383 35737
rect 29383 35703 29417 35737
rect 29417 35703 29426 35737
rect 29374 35694 29426 35703
rect 33534 35737 33586 35746
rect 33534 35703 33543 35737
rect 33543 35703 33577 35737
rect 33577 35703 33586 35737
rect 33534 35694 33586 35703
rect 33694 35737 33746 35746
rect 33694 35703 33703 35737
rect 33703 35703 33737 35737
rect 33737 35703 33746 35737
rect 33694 35694 33746 35703
rect 33854 35737 33906 35746
rect 33854 35703 33863 35737
rect 33863 35703 33897 35737
rect 33897 35703 33906 35737
rect 33854 35694 33906 35703
rect 34014 35737 34066 35746
rect 34014 35703 34023 35737
rect 34023 35703 34057 35737
rect 34057 35703 34066 35737
rect 34014 35694 34066 35703
rect 34174 35737 34226 35746
rect 34174 35703 34183 35737
rect 34183 35703 34217 35737
rect 34217 35703 34226 35737
rect 34174 35694 34226 35703
rect 34334 35737 34386 35746
rect 34334 35703 34343 35737
rect 34343 35703 34377 35737
rect 34377 35703 34386 35737
rect 34334 35694 34386 35703
rect 34494 35737 34546 35746
rect 34494 35703 34503 35737
rect 34503 35703 34537 35737
rect 34537 35703 34546 35737
rect 34494 35694 34546 35703
rect 34654 35737 34706 35746
rect 34654 35703 34663 35737
rect 34663 35703 34697 35737
rect 34697 35703 34706 35737
rect 34654 35694 34706 35703
rect 34814 35737 34866 35746
rect 34814 35703 34823 35737
rect 34823 35703 34857 35737
rect 34857 35703 34866 35737
rect 34814 35694 34866 35703
rect 34974 35737 35026 35746
rect 34974 35703 34983 35737
rect 34983 35703 35017 35737
rect 35017 35703 35026 35737
rect 34974 35694 35026 35703
rect 35134 35737 35186 35746
rect 35134 35703 35143 35737
rect 35143 35703 35177 35737
rect 35177 35703 35186 35737
rect 35134 35694 35186 35703
rect 35294 35737 35346 35746
rect 35294 35703 35303 35737
rect 35303 35703 35337 35737
rect 35337 35703 35346 35737
rect 35294 35694 35346 35703
rect 35454 35737 35506 35746
rect 35454 35703 35463 35737
rect 35463 35703 35497 35737
rect 35497 35703 35506 35737
rect 35454 35694 35506 35703
rect 35614 35737 35666 35746
rect 35614 35703 35623 35737
rect 35623 35703 35657 35737
rect 35657 35703 35666 35737
rect 35614 35694 35666 35703
rect 35774 35737 35826 35746
rect 35774 35703 35783 35737
rect 35783 35703 35817 35737
rect 35817 35703 35826 35737
rect 35774 35694 35826 35703
rect 35934 35737 35986 35746
rect 35934 35703 35943 35737
rect 35943 35703 35977 35737
rect 35977 35703 35986 35737
rect 35934 35694 35986 35703
rect 36094 35737 36146 35746
rect 36094 35703 36103 35737
rect 36103 35703 36137 35737
rect 36137 35703 36146 35737
rect 36094 35694 36146 35703
rect 36254 35737 36306 35746
rect 36254 35703 36263 35737
rect 36263 35703 36297 35737
rect 36297 35703 36306 35737
rect 36254 35694 36306 35703
rect 36414 35737 36466 35746
rect 36414 35703 36423 35737
rect 36423 35703 36457 35737
rect 36457 35703 36466 35737
rect 36414 35694 36466 35703
rect 36574 35737 36626 35746
rect 36574 35703 36583 35737
rect 36583 35703 36617 35737
rect 36617 35703 36626 35737
rect 36574 35694 36626 35703
rect 36734 35737 36786 35746
rect 36734 35703 36743 35737
rect 36743 35703 36777 35737
rect 36777 35703 36786 35737
rect 36734 35694 36786 35703
rect 36894 35737 36946 35746
rect 36894 35703 36903 35737
rect 36903 35703 36937 35737
rect 36937 35703 36946 35737
rect 36894 35694 36946 35703
rect 37054 35737 37106 35746
rect 37054 35703 37063 35737
rect 37063 35703 37097 35737
rect 37097 35703 37106 35737
rect 37054 35694 37106 35703
rect 37214 35737 37266 35746
rect 37214 35703 37223 35737
rect 37223 35703 37257 35737
rect 37257 35703 37266 35737
rect 37214 35694 37266 35703
rect 37374 35737 37426 35746
rect 37374 35703 37383 35737
rect 37383 35703 37417 35737
rect 37417 35703 37426 35737
rect 37374 35694 37426 35703
rect 37534 35737 37586 35746
rect 37534 35703 37543 35737
rect 37543 35703 37577 35737
rect 37577 35703 37586 35737
rect 37534 35694 37586 35703
rect 37694 35737 37746 35746
rect 37694 35703 37703 35737
rect 37703 35703 37737 35737
rect 37737 35703 37746 35737
rect 37694 35694 37746 35703
rect 37854 35737 37906 35746
rect 37854 35703 37863 35737
rect 37863 35703 37897 35737
rect 37897 35703 37906 35737
rect 37854 35694 37906 35703
rect 38014 35737 38066 35746
rect 38014 35703 38023 35737
rect 38023 35703 38057 35737
rect 38057 35703 38066 35737
rect 38014 35694 38066 35703
rect 38174 35737 38226 35746
rect 38174 35703 38183 35737
rect 38183 35703 38217 35737
rect 38217 35703 38226 35737
rect 38174 35694 38226 35703
rect 38334 35737 38386 35746
rect 38334 35703 38343 35737
rect 38343 35703 38377 35737
rect 38377 35703 38386 35737
rect 38334 35694 38386 35703
rect 38494 35737 38546 35746
rect 38494 35703 38503 35737
rect 38503 35703 38537 35737
rect 38537 35703 38546 35737
rect 38494 35694 38546 35703
rect 38654 35737 38706 35746
rect 38654 35703 38663 35737
rect 38663 35703 38697 35737
rect 38697 35703 38706 35737
rect 38654 35694 38706 35703
rect 38814 35737 38866 35746
rect 38814 35703 38823 35737
rect 38823 35703 38857 35737
rect 38857 35703 38866 35737
rect 38814 35694 38866 35703
rect 38974 35737 39026 35746
rect 38974 35703 38983 35737
rect 38983 35703 39017 35737
rect 39017 35703 39026 35737
rect 38974 35694 39026 35703
rect 39134 35737 39186 35746
rect 39134 35703 39143 35737
rect 39143 35703 39177 35737
rect 39177 35703 39186 35737
rect 39134 35694 39186 35703
rect 39294 35737 39346 35746
rect 39294 35703 39303 35737
rect 39303 35703 39337 35737
rect 39337 35703 39346 35737
rect 39294 35694 39346 35703
rect 39454 35737 39506 35746
rect 39454 35703 39463 35737
rect 39463 35703 39497 35737
rect 39497 35703 39506 35737
rect 39454 35694 39506 35703
rect 39614 35737 39666 35746
rect 39614 35703 39623 35737
rect 39623 35703 39657 35737
rect 39657 35703 39666 35737
rect 39614 35694 39666 35703
rect 39774 35737 39826 35746
rect 39774 35703 39783 35737
rect 39783 35703 39817 35737
rect 39817 35703 39826 35737
rect 39774 35694 39826 35703
rect 39934 35737 39986 35746
rect 39934 35703 39943 35737
rect 39943 35703 39977 35737
rect 39977 35703 39986 35737
rect 39934 35694 39986 35703
rect 40094 35737 40146 35746
rect 40094 35703 40103 35737
rect 40103 35703 40137 35737
rect 40137 35703 40146 35737
rect 40094 35694 40146 35703
rect 40254 35737 40306 35746
rect 40254 35703 40263 35737
rect 40263 35703 40297 35737
rect 40297 35703 40306 35737
rect 40254 35694 40306 35703
rect 40414 35737 40466 35746
rect 40414 35703 40423 35737
rect 40423 35703 40457 35737
rect 40457 35703 40466 35737
rect 40414 35694 40466 35703
rect 40574 35737 40626 35746
rect 40574 35703 40583 35737
rect 40583 35703 40617 35737
rect 40617 35703 40626 35737
rect 40574 35694 40626 35703
rect 40734 35737 40786 35746
rect 40734 35703 40743 35737
rect 40743 35703 40777 35737
rect 40777 35703 40786 35737
rect 40734 35694 40786 35703
rect 40894 35737 40946 35746
rect 40894 35703 40903 35737
rect 40903 35703 40937 35737
rect 40937 35703 40946 35737
rect 40894 35694 40946 35703
rect 41054 35737 41106 35746
rect 41054 35703 41063 35737
rect 41063 35703 41097 35737
rect 41097 35703 41106 35737
rect 41054 35694 41106 35703
rect 41214 35737 41266 35746
rect 41214 35703 41223 35737
rect 41223 35703 41257 35737
rect 41257 35703 41266 35737
rect 41214 35694 41266 35703
rect 41374 35737 41426 35746
rect 41374 35703 41383 35737
rect 41383 35703 41417 35737
rect 41417 35703 41426 35737
rect 41374 35694 41426 35703
rect 41534 35737 41586 35746
rect 41534 35703 41543 35737
rect 41543 35703 41577 35737
rect 41577 35703 41586 35737
rect 41534 35694 41586 35703
rect 41694 35737 41746 35746
rect 41694 35703 41703 35737
rect 41703 35703 41737 35737
rect 41737 35703 41746 35737
rect 41694 35694 41746 35703
rect 41854 35737 41906 35746
rect 41854 35703 41863 35737
rect 41863 35703 41897 35737
rect 41897 35703 41906 35737
rect 41854 35694 41906 35703
rect 14 35417 66 35426
rect 14 35383 23 35417
rect 23 35383 57 35417
rect 57 35383 66 35417
rect 14 35374 66 35383
rect 174 35417 226 35426
rect 174 35383 183 35417
rect 183 35383 217 35417
rect 217 35383 226 35417
rect 174 35374 226 35383
rect 334 35417 386 35426
rect 334 35383 343 35417
rect 343 35383 377 35417
rect 377 35383 386 35417
rect 334 35374 386 35383
rect 494 35417 546 35426
rect 494 35383 503 35417
rect 503 35383 537 35417
rect 537 35383 546 35417
rect 494 35374 546 35383
rect 654 35417 706 35426
rect 654 35383 663 35417
rect 663 35383 697 35417
rect 697 35383 706 35417
rect 654 35374 706 35383
rect 814 35417 866 35426
rect 814 35383 823 35417
rect 823 35383 857 35417
rect 857 35383 866 35417
rect 814 35374 866 35383
rect 974 35417 1026 35426
rect 974 35383 983 35417
rect 983 35383 1017 35417
rect 1017 35383 1026 35417
rect 974 35374 1026 35383
rect 1134 35417 1186 35426
rect 1134 35383 1143 35417
rect 1143 35383 1177 35417
rect 1177 35383 1186 35417
rect 1134 35374 1186 35383
rect 1294 35417 1346 35426
rect 1294 35383 1303 35417
rect 1303 35383 1337 35417
rect 1337 35383 1346 35417
rect 1294 35374 1346 35383
rect 1454 35417 1506 35426
rect 1454 35383 1463 35417
rect 1463 35383 1497 35417
rect 1497 35383 1506 35417
rect 1454 35374 1506 35383
rect 1614 35417 1666 35426
rect 1614 35383 1623 35417
rect 1623 35383 1657 35417
rect 1657 35383 1666 35417
rect 1614 35374 1666 35383
rect 1774 35417 1826 35426
rect 1774 35383 1783 35417
rect 1783 35383 1817 35417
rect 1817 35383 1826 35417
rect 1774 35374 1826 35383
rect 1934 35417 1986 35426
rect 1934 35383 1943 35417
rect 1943 35383 1977 35417
rect 1977 35383 1986 35417
rect 1934 35374 1986 35383
rect 2094 35417 2146 35426
rect 2094 35383 2103 35417
rect 2103 35383 2137 35417
rect 2137 35383 2146 35417
rect 2094 35374 2146 35383
rect 2254 35417 2306 35426
rect 2254 35383 2263 35417
rect 2263 35383 2297 35417
rect 2297 35383 2306 35417
rect 2254 35374 2306 35383
rect 2414 35417 2466 35426
rect 2414 35383 2423 35417
rect 2423 35383 2457 35417
rect 2457 35383 2466 35417
rect 2414 35374 2466 35383
rect 2574 35417 2626 35426
rect 2574 35383 2583 35417
rect 2583 35383 2617 35417
rect 2617 35383 2626 35417
rect 2574 35374 2626 35383
rect 2734 35417 2786 35426
rect 2734 35383 2743 35417
rect 2743 35383 2777 35417
rect 2777 35383 2786 35417
rect 2734 35374 2786 35383
rect 2894 35417 2946 35426
rect 2894 35383 2903 35417
rect 2903 35383 2937 35417
rect 2937 35383 2946 35417
rect 2894 35374 2946 35383
rect 3054 35417 3106 35426
rect 3054 35383 3063 35417
rect 3063 35383 3097 35417
rect 3097 35383 3106 35417
rect 3054 35374 3106 35383
rect 3214 35417 3266 35426
rect 3214 35383 3223 35417
rect 3223 35383 3257 35417
rect 3257 35383 3266 35417
rect 3214 35374 3266 35383
rect 3374 35417 3426 35426
rect 3374 35383 3383 35417
rect 3383 35383 3417 35417
rect 3417 35383 3426 35417
rect 3374 35374 3426 35383
rect 3534 35417 3586 35426
rect 3534 35383 3543 35417
rect 3543 35383 3577 35417
rect 3577 35383 3586 35417
rect 3534 35374 3586 35383
rect 3694 35417 3746 35426
rect 3694 35383 3703 35417
rect 3703 35383 3737 35417
rect 3737 35383 3746 35417
rect 3694 35374 3746 35383
rect 3854 35417 3906 35426
rect 3854 35383 3863 35417
rect 3863 35383 3897 35417
rect 3897 35383 3906 35417
rect 3854 35374 3906 35383
rect 4014 35417 4066 35426
rect 4014 35383 4023 35417
rect 4023 35383 4057 35417
rect 4057 35383 4066 35417
rect 4014 35374 4066 35383
rect 4174 35417 4226 35426
rect 4174 35383 4183 35417
rect 4183 35383 4217 35417
rect 4217 35383 4226 35417
rect 4174 35374 4226 35383
rect 4334 35417 4386 35426
rect 4334 35383 4343 35417
rect 4343 35383 4377 35417
rect 4377 35383 4386 35417
rect 4334 35374 4386 35383
rect 4494 35417 4546 35426
rect 4494 35383 4503 35417
rect 4503 35383 4537 35417
rect 4537 35383 4546 35417
rect 4494 35374 4546 35383
rect 4654 35417 4706 35426
rect 4654 35383 4663 35417
rect 4663 35383 4697 35417
rect 4697 35383 4706 35417
rect 4654 35374 4706 35383
rect 4814 35417 4866 35426
rect 4814 35383 4823 35417
rect 4823 35383 4857 35417
rect 4857 35383 4866 35417
rect 4814 35374 4866 35383
rect 4974 35417 5026 35426
rect 4974 35383 4983 35417
rect 4983 35383 5017 35417
rect 5017 35383 5026 35417
rect 4974 35374 5026 35383
rect 5134 35417 5186 35426
rect 5134 35383 5143 35417
rect 5143 35383 5177 35417
rect 5177 35383 5186 35417
rect 5134 35374 5186 35383
rect 5294 35417 5346 35426
rect 5294 35383 5303 35417
rect 5303 35383 5337 35417
rect 5337 35383 5346 35417
rect 5294 35374 5346 35383
rect 5454 35417 5506 35426
rect 5454 35383 5463 35417
rect 5463 35383 5497 35417
rect 5497 35383 5506 35417
rect 5454 35374 5506 35383
rect 5614 35417 5666 35426
rect 5614 35383 5623 35417
rect 5623 35383 5657 35417
rect 5657 35383 5666 35417
rect 5614 35374 5666 35383
rect 5774 35417 5826 35426
rect 5774 35383 5783 35417
rect 5783 35383 5817 35417
rect 5817 35383 5826 35417
rect 5774 35374 5826 35383
rect 5934 35417 5986 35426
rect 5934 35383 5943 35417
rect 5943 35383 5977 35417
rect 5977 35383 5986 35417
rect 5934 35374 5986 35383
rect 6094 35417 6146 35426
rect 6094 35383 6103 35417
rect 6103 35383 6137 35417
rect 6137 35383 6146 35417
rect 6094 35374 6146 35383
rect 6254 35417 6306 35426
rect 6254 35383 6263 35417
rect 6263 35383 6297 35417
rect 6297 35383 6306 35417
rect 6254 35374 6306 35383
rect 6414 35417 6466 35426
rect 6414 35383 6423 35417
rect 6423 35383 6457 35417
rect 6457 35383 6466 35417
rect 6414 35374 6466 35383
rect 6574 35417 6626 35426
rect 6574 35383 6583 35417
rect 6583 35383 6617 35417
rect 6617 35383 6626 35417
rect 6574 35374 6626 35383
rect 6734 35417 6786 35426
rect 6734 35383 6743 35417
rect 6743 35383 6777 35417
rect 6777 35383 6786 35417
rect 6734 35374 6786 35383
rect 6894 35417 6946 35426
rect 6894 35383 6903 35417
rect 6903 35383 6937 35417
rect 6937 35383 6946 35417
rect 6894 35374 6946 35383
rect 7054 35417 7106 35426
rect 7054 35383 7063 35417
rect 7063 35383 7097 35417
rect 7097 35383 7106 35417
rect 7054 35374 7106 35383
rect 7214 35417 7266 35426
rect 7214 35383 7223 35417
rect 7223 35383 7257 35417
rect 7257 35383 7266 35417
rect 7214 35374 7266 35383
rect 7374 35417 7426 35426
rect 7374 35383 7383 35417
rect 7383 35383 7417 35417
rect 7417 35383 7426 35417
rect 7374 35374 7426 35383
rect 7534 35417 7586 35426
rect 7534 35383 7543 35417
rect 7543 35383 7577 35417
rect 7577 35383 7586 35417
rect 7534 35374 7586 35383
rect 7694 35417 7746 35426
rect 7694 35383 7703 35417
rect 7703 35383 7737 35417
rect 7737 35383 7746 35417
rect 7694 35374 7746 35383
rect 7854 35417 7906 35426
rect 7854 35383 7863 35417
rect 7863 35383 7897 35417
rect 7897 35383 7906 35417
rect 7854 35374 7906 35383
rect 8014 35417 8066 35426
rect 8014 35383 8023 35417
rect 8023 35383 8057 35417
rect 8057 35383 8066 35417
rect 8014 35374 8066 35383
rect 8174 35417 8226 35426
rect 8174 35383 8183 35417
rect 8183 35383 8217 35417
rect 8217 35383 8226 35417
rect 8174 35374 8226 35383
rect 8334 35417 8386 35426
rect 8334 35383 8343 35417
rect 8343 35383 8377 35417
rect 8377 35383 8386 35417
rect 8334 35374 8386 35383
rect 12494 35417 12546 35426
rect 12494 35383 12503 35417
rect 12503 35383 12537 35417
rect 12537 35383 12546 35417
rect 12494 35374 12546 35383
rect 12654 35417 12706 35426
rect 12654 35383 12663 35417
rect 12663 35383 12697 35417
rect 12697 35383 12706 35417
rect 12654 35374 12706 35383
rect 12814 35417 12866 35426
rect 12814 35383 12823 35417
rect 12823 35383 12857 35417
rect 12857 35383 12866 35417
rect 12814 35374 12866 35383
rect 12974 35417 13026 35426
rect 12974 35383 12983 35417
rect 12983 35383 13017 35417
rect 13017 35383 13026 35417
rect 12974 35374 13026 35383
rect 13134 35417 13186 35426
rect 13134 35383 13143 35417
rect 13143 35383 13177 35417
rect 13177 35383 13186 35417
rect 13134 35374 13186 35383
rect 13294 35417 13346 35426
rect 13294 35383 13303 35417
rect 13303 35383 13337 35417
rect 13337 35383 13346 35417
rect 13294 35374 13346 35383
rect 13454 35417 13506 35426
rect 13454 35383 13463 35417
rect 13463 35383 13497 35417
rect 13497 35383 13506 35417
rect 13454 35374 13506 35383
rect 13614 35417 13666 35426
rect 13614 35383 13623 35417
rect 13623 35383 13657 35417
rect 13657 35383 13666 35417
rect 13614 35374 13666 35383
rect 13774 35417 13826 35426
rect 13774 35383 13783 35417
rect 13783 35383 13817 35417
rect 13817 35383 13826 35417
rect 13774 35374 13826 35383
rect 13934 35417 13986 35426
rect 13934 35383 13943 35417
rect 13943 35383 13977 35417
rect 13977 35383 13986 35417
rect 13934 35374 13986 35383
rect 14094 35417 14146 35426
rect 14094 35383 14103 35417
rect 14103 35383 14137 35417
rect 14137 35383 14146 35417
rect 14094 35374 14146 35383
rect 14254 35417 14306 35426
rect 14254 35383 14263 35417
rect 14263 35383 14297 35417
rect 14297 35383 14306 35417
rect 14254 35374 14306 35383
rect 14414 35417 14466 35426
rect 14414 35383 14423 35417
rect 14423 35383 14457 35417
rect 14457 35383 14466 35417
rect 14414 35374 14466 35383
rect 14574 35417 14626 35426
rect 14574 35383 14583 35417
rect 14583 35383 14617 35417
rect 14617 35383 14626 35417
rect 14574 35374 14626 35383
rect 14734 35417 14786 35426
rect 14734 35383 14743 35417
rect 14743 35383 14777 35417
rect 14777 35383 14786 35417
rect 14734 35374 14786 35383
rect 14894 35417 14946 35426
rect 14894 35383 14903 35417
rect 14903 35383 14937 35417
rect 14937 35383 14946 35417
rect 14894 35374 14946 35383
rect 15054 35417 15106 35426
rect 15054 35383 15063 35417
rect 15063 35383 15097 35417
rect 15097 35383 15106 35417
rect 15054 35374 15106 35383
rect 15214 35417 15266 35426
rect 15214 35383 15223 35417
rect 15223 35383 15257 35417
rect 15257 35383 15266 35417
rect 15214 35374 15266 35383
rect 15374 35417 15426 35426
rect 15374 35383 15383 35417
rect 15383 35383 15417 35417
rect 15417 35383 15426 35417
rect 15374 35374 15426 35383
rect 15534 35417 15586 35426
rect 15534 35383 15543 35417
rect 15543 35383 15577 35417
rect 15577 35383 15586 35417
rect 15534 35374 15586 35383
rect 15694 35417 15746 35426
rect 15694 35383 15703 35417
rect 15703 35383 15737 35417
rect 15737 35383 15746 35417
rect 15694 35374 15746 35383
rect 15854 35417 15906 35426
rect 15854 35383 15863 35417
rect 15863 35383 15897 35417
rect 15897 35383 15906 35417
rect 15854 35374 15906 35383
rect 16014 35417 16066 35426
rect 16014 35383 16023 35417
rect 16023 35383 16057 35417
rect 16057 35383 16066 35417
rect 16014 35374 16066 35383
rect 16174 35417 16226 35426
rect 16174 35383 16183 35417
rect 16183 35383 16217 35417
rect 16217 35383 16226 35417
rect 16174 35374 16226 35383
rect 16334 35417 16386 35426
rect 16334 35383 16343 35417
rect 16343 35383 16377 35417
rect 16377 35383 16386 35417
rect 16334 35374 16386 35383
rect 16494 35417 16546 35426
rect 16494 35383 16503 35417
rect 16503 35383 16537 35417
rect 16537 35383 16546 35417
rect 16494 35374 16546 35383
rect 16654 35417 16706 35426
rect 16654 35383 16663 35417
rect 16663 35383 16697 35417
rect 16697 35383 16706 35417
rect 16654 35374 16706 35383
rect 16814 35417 16866 35426
rect 16814 35383 16823 35417
rect 16823 35383 16857 35417
rect 16857 35383 16866 35417
rect 16814 35374 16866 35383
rect 16974 35417 17026 35426
rect 16974 35383 16983 35417
rect 16983 35383 17017 35417
rect 17017 35383 17026 35417
rect 16974 35374 17026 35383
rect 17134 35417 17186 35426
rect 17134 35383 17143 35417
rect 17143 35383 17177 35417
rect 17177 35383 17186 35417
rect 17134 35374 17186 35383
rect 17294 35417 17346 35426
rect 17294 35383 17303 35417
rect 17303 35383 17337 35417
rect 17337 35383 17346 35417
rect 17294 35374 17346 35383
rect 17454 35417 17506 35426
rect 17454 35383 17463 35417
rect 17463 35383 17497 35417
rect 17497 35383 17506 35417
rect 17454 35374 17506 35383
rect 17614 35417 17666 35426
rect 17614 35383 17623 35417
rect 17623 35383 17657 35417
rect 17657 35383 17666 35417
rect 17614 35374 17666 35383
rect 17774 35417 17826 35426
rect 17774 35383 17783 35417
rect 17783 35383 17817 35417
rect 17817 35383 17826 35417
rect 17774 35374 17826 35383
rect 17934 35417 17986 35426
rect 17934 35383 17943 35417
rect 17943 35383 17977 35417
rect 17977 35383 17986 35417
rect 17934 35374 17986 35383
rect 18094 35417 18146 35426
rect 18094 35383 18103 35417
rect 18103 35383 18137 35417
rect 18137 35383 18146 35417
rect 18094 35374 18146 35383
rect 18254 35417 18306 35426
rect 18254 35383 18263 35417
rect 18263 35383 18297 35417
rect 18297 35383 18306 35417
rect 18254 35374 18306 35383
rect 18414 35417 18466 35426
rect 18414 35383 18423 35417
rect 18423 35383 18457 35417
rect 18457 35383 18466 35417
rect 18414 35374 18466 35383
rect 18574 35417 18626 35426
rect 18574 35383 18583 35417
rect 18583 35383 18617 35417
rect 18617 35383 18626 35417
rect 18574 35374 18626 35383
rect 18734 35417 18786 35426
rect 18734 35383 18743 35417
rect 18743 35383 18777 35417
rect 18777 35383 18786 35417
rect 18734 35374 18786 35383
rect 18894 35417 18946 35426
rect 18894 35383 18903 35417
rect 18903 35383 18937 35417
rect 18937 35383 18946 35417
rect 18894 35374 18946 35383
rect 23134 35417 23186 35426
rect 23134 35383 23143 35417
rect 23143 35383 23177 35417
rect 23177 35383 23186 35417
rect 23134 35374 23186 35383
rect 23294 35417 23346 35426
rect 23294 35383 23303 35417
rect 23303 35383 23337 35417
rect 23337 35383 23346 35417
rect 23294 35374 23346 35383
rect 23454 35417 23506 35426
rect 23454 35383 23463 35417
rect 23463 35383 23497 35417
rect 23497 35383 23506 35417
rect 23454 35374 23506 35383
rect 23614 35417 23666 35426
rect 23614 35383 23623 35417
rect 23623 35383 23657 35417
rect 23657 35383 23666 35417
rect 23614 35374 23666 35383
rect 23774 35417 23826 35426
rect 23774 35383 23783 35417
rect 23783 35383 23817 35417
rect 23817 35383 23826 35417
rect 23774 35374 23826 35383
rect 23934 35417 23986 35426
rect 23934 35383 23943 35417
rect 23943 35383 23977 35417
rect 23977 35383 23986 35417
rect 23934 35374 23986 35383
rect 24094 35417 24146 35426
rect 24094 35383 24103 35417
rect 24103 35383 24137 35417
rect 24137 35383 24146 35417
rect 24094 35374 24146 35383
rect 24254 35417 24306 35426
rect 24254 35383 24263 35417
rect 24263 35383 24297 35417
rect 24297 35383 24306 35417
rect 24254 35374 24306 35383
rect 24414 35417 24466 35426
rect 24414 35383 24423 35417
rect 24423 35383 24457 35417
rect 24457 35383 24466 35417
rect 24414 35374 24466 35383
rect 24574 35417 24626 35426
rect 24574 35383 24583 35417
rect 24583 35383 24617 35417
rect 24617 35383 24626 35417
rect 24574 35374 24626 35383
rect 24734 35417 24786 35426
rect 24734 35383 24743 35417
rect 24743 35383 24777 35417
rect 24777 35383 24786 35417
rect 24734 35374 24786 35383
rect 24894 35417 24946 35426
rect 24894 35383 24903 35417
rect 24903 35383 24937 35417
rect 24937 35383 24946 35417
rect 24894 35374 24946 35383
rect 25054 35417 25106 35426
rect 25054 35383 25063 35417
rect 25063 35383 25097 35417
rect 25097 35383 25106 35417
rect 25054 35374 25106 35383
rect 25214 35417 25266 35426
rect 25214 35383 25223 35417
rect 25223 35383 25257 35417
rect 25257 35383 25266 35417
rect 25214 35374 25266 35383
rect 25374 35417 25426 35426
rect 25374 35383 25383 35417
rect 25383 35383 25417 35417
rect 25417 35383 25426 35417
rect 25374 35374 25426 35383
rect 25534 35417 25586 35426
rect 25534 35383 25543 35417
rect 25543 35383 25577 35417
rect 25577 35383 25586 35417
rect 25534 35374 25586 35383
rect 25694 35417 25746 35426
rect 25694 35383 25703 35417
rect 25703 35383 25737 35417
rect 25737 35383 25746 35417
rect 25694 35374 25746 35383
rect 25854 35417 25906 35426
rect 25854 35383 25863 35417
rect 25863 35383 25897 35417
rect 25897 35383 25906 35417
rect 25854 35374 25906 35383
rect 26014 35417 26066 35426
rect 26014 35383 26023 35417
rect 26023 35383 26057 35417
rect 26057 35383 26066 35417
rect 26014 35374 26066 35383
rect 26174 35417 26226 35426
rect 26174 35383 26183 35417
rect 26183 35383 26217 35417
rect 26217 35383 26226 35417
rect 26174 35374 26226 35383
rect 26334 35417 26386 35426
rect 26334 35383 26343 35417
rect 26343 35383 26377 35417
rect 26377 35383 26386 35417
rect 26334 35374 26386 35383
rect 26494 35417 26546 35426
rect 26494 35383 26503 35417
rect 26503 35383 26537 35417
rect 26537 35383 26546 35417
rect 26494 35374 26546 35383
rect 26654 35417 26706 35426
rect 26654 35383 26663 35417
rect 26663 35383 26697 35417
rect 26697 35383 26706 35417
rect 26654 35374 26706 35383
rect 26814 35417 26866 35426
rect 26814 35383 26823 35417
rect 26823 35383 26857 35417
rect 26857 35383 26866 35417
rect 26814 35374 26866 35383
rect 26974 35417 27026 35426
rect 26974 35383 26983 35417
rect 26983 35383 27017 35417
rect 27017 35383 27026 35417
rect 26974 35374 27026 35383
rect 27134 35417 27186 35426
rect 27134 35383 27143 35417
rect 27143 35383 27177 35417
rect 27177 35383 27186 35417
rect 27134 35374 27186 35383
rect 27294 35417 27346 35426
rect 27294 35383 27303 35417
rect 27303 35383 27337 35417
rect 27337 35383 27346 35417
rect 27294 35374 27346 35383
rect 27454 35417 27506 35426
rect 27454 35383 27463 35417
rect 27463 35383 27497 35417
rect 27497 35383 27506 35417
rect 27454 35374 27506 35383
rect 27614 35417 27666 35426
rect 27614 35383 27623 35417
rect 27623 35383 27657 35417
rect 27657 35383 27666 35417
rect 27614 35374 27666 35383
rect 27774 35417 27826 35426
rect 27774 35383 27783 35417
rect 27783 35383 27817 35417
rect 27817 35383 27826 35417
rect 27774 35374 27826 35383
rect 27934 35417 27986 35426
rect 27934 35383 27943 35417
rect 27943 35383 27977 35417
rect 27977 35383 27986 35417
rect 27934 35374 27986 35383
rect 28094 35417 28146 35426
rect 28094 35383 28103 35417
rect 28103 35383 28137 35417
rect 28137 35383 28146 35417
rect 28094 35374 28146 35383
rect 28254 35417 28306 35426
rect 28254 35383 28263 35417
rect 28263 35383 28297 35417
rect 28297 35383 28306 35417
rect 28254 35374 28306 35383
rect 28414 35417 28466 35426
rect 28414 35383 28423 35417
rect 28423 35383 28457 35417
rect 28457 35383 28466 35417
rect 28414 35374 28466 35383
rect 28574 35417 28626 35426
rect 28574 35383 28583 35417
rect 28583 35383 28617 35417
rect 28617 35383 28626 35417
rect 28574 35374 28626 35383
rect 28734 35417 28786 35426
rect 28734 35383 28743 35417
rect 28743 35383 28777 35417
rect 28777 35383 28786 35417
rect 28734 35374 28786 35383
rect 28894 35417 28946 35426
rect 28894 35383 28903 35417
rect 28903 35383 28937 35417
rect 28937 35383 28946 35417
rect 28894 35374 28946 35383
rect 29054 35417 29106 35426
rect 29054 35383 29063 35417
rect 29063 35383 29097 35417
rect 29097 35383 29106 35417
rect 29054 35374 29106 35383
rect 29214 35417 29266 35426
rect 29214 35383 29223 35417
rect 29223 35383 29257 35417
rect 29257 35383 29266 35417
rect 29214 35374 29266 35383
rect 29374 35417 29426 35426
rect 29374 35383 29383 35417
rect 29383 35383 29417 35417
rect 29417 35383 29426 35417
rect 29374 35374 29426 35383
rect 33534 35417 33586 35426
rect 33534 35383 33543 35417
rect 33543 35383 33577 35417
rect 33577 35383 33586 35417
rect 33534 35374 33586 35383
rect 33694 35417 33746 35426
rect 33694 35383 33703 35417
rect 33703 35383 33737 35417
rect 33737 35383 33746 35417
rect 33694 35374 33746 35383
rect 33854 35417 33906 35426
rect 33854 35383 33863 35417
rect 33863 35383 33897 35417
rect 33897 35383 33906 35417
rect 33854 35374 33906 35383
rect 34014 35417 34066 35426
rect 34014 35383 34023 35417
rect 34023 35383 34057 35417
rect 34057 35383 34066 35417
rect 34014 35374 34066 35383
rect 34174 35417 34226 35426
rect 34174 35383 34183 35417
rect 34183 35383 34217 35417
rect 34217 35383 34226 35417
rect 34174 35374 34226 35383
rect 34334 35417 34386 35426
rect 34334 35383 34343 35417
rect 34343 35383 34377 35417
rect 34377 35383 34386 35417
rect 34334 35374 34386 35383
rect 34494 35417 34546 35426
rect 34494 35383 34503 35417
rect 34503 35383 34537 35417
rect 34537 35383 34546 35417
rect 34494 35374 34546 35383
rect 34654 35417 34706 35426
rect 34654 35383 34663 35417
rect 34663 35383 34697 35417
rect 34697 35383 34706 35417
rect 34654 35374 34706 35383
rect 34814 35417 34866 35426
rect 34814 35383 34823 35417
rect 34823 35383 34857 35417
rect 34857 35383 34866 35417
rect 34814 35374 34866 35383
rect 34974 35417 35026 35426
rect 34974 35383 34983 35417
rect 34983 35383 35017 35417
rect 35017 35383 35026 35417
rect 34974 35374 35026 35383
rect 35134 35417 35186 35426
rect 35134 35383 35143 35417
rect 35143 35383 35177 35417
rect 35177 35383 35186 35417
rect 35134 35374 35186 35383
rect 35294 35417 35346 35426
rect 35294 35383 35303 35417
rect 35303 35383 35337 35417
rect 35337 35383 35346 35417
rect 35294 35374 35346 35383
rect 35454 35417 35506 35426
rect 35454 35383 35463 35417
rect 35463 35383 35497 35417
rect 35497 35383 35506 35417
rect 35454 35374 35506 35383
rect 35614 35417 35666 35426
rect 35614 35383 35623 35417
rect 35623 35383 35657 35417
rect 35657 35383 35666 35417
rect 35614 35374 35666 35383
rect 35774 35417 35826 35426
rect 35774 35383 35783 35417
rect 35783 35383 35817 35417
rect 35817 35383 35826 35417
rect 35774 35374 35826 35383
rect 35934 35417 35986 35426
rect 35934 35383 35943 35417
rect 35943 35383 35977 35417
rect 35977 35383 35986 35417
rect 35934 35374 35986 35383
rect 36094 35417 36146 35426
rect 36094 35383 36103 35417
rect 36103 35383 36137 35417
rect 36137 35383 36146 35417
rect 36094 35374 36146 35383
rect 36254 35417 36306 35426
rect 36254 35383 36263 35417
rect 36263 35383 36297 35417
rect 36297 35383 36306 35417
rect 36254 35374 36306 35383
rect 36414 35417 36466 35426
rect 36414 35383 36423 35417
rect 36423 35383 36457 35417
rect 36457 35383 36466 35417
rect 36414 35374 36466 35383
rect 36574 35417 36626 35426
rect 36574 35383 36583 35417
rect 36583 35383 36617 35417
rect 36617 35383 36626 35417
rect 36574 35374 36626 35383
rect 36734 35417 36786 35426
rect 36734 35383 36743 35417
rect 36743 35383 36777 35417
rect 36777 35383 36786 35417
rect 36734 35374 36786 35383
rect 36894 35417 36946 35426
rect 36894 35383 36903 35417
rect 36903 35383 36937 35417
rect 36937 35383 36946 35417
rect 36894 35374 36946 35383
rect 37054 35417 37106 35426
rect 37054 35383 37063 35417
rect 37063 35383 37097 35417
rect 37097 35383 37106 35417
rect 37054 35374 37106 35383
rect 37214 35417 37266 35426
rect 37214 35383 37223 35417
rect 37223 35383 37257 35417
rect 37257 35383 37266 35417
rect 37214 35374 37266 35383
rect 37374 35417 37426 35426
rect 37374 35383 37383 35417
rect 37383 35383 37417 35417
rect 37417 35383 37426 35417
rect 37374 35374 37426 35383
rect 37534 35417 37586 35426
rect 37534 35383 37543 35417
rect 37543 35383 37577 35417
rect 37577 35383 37586 35417
rect 37534 35374 37586 35383
rect 37694 35417 37746 35426
rect 37694 35383 37703 35417
rect 37703 35383 37737 35417
rect 37737 35383 37746 35417
rect 37694 35374 37746 35383
rect 37854 35417 37906 35426
rect 37854 35383 37863 35417
rect 37863 35383 37897 35417
rect 37897 35383 37906 35417
rect 37854 35374 37906 35383
rect 38014 35417 38066 35426
rect 38014 35383 38023 35417
rect 38023 35383 38057 35417
rect 38057 35383 38066 35417
rect 38014 35374 38066 35383
rect 38174 35417 38226 35426
rect 38174 35383 38183 35417
rect 38183 35383 38217 35417
rect 38217 35383 38226 35417
rect 38174 35374 38226 35383
rect 38334 35417 38386 35426
rect 38334 35383 38343 35417
rect 38343 35383 38377 35417
rect 38377 35383 38386 35417
rect 38334 35374 38386 35383
rect 38494 35417 38546 35426
rect 38494 35383 38503 35417
rect 38503 35383 38537 35417
rect 38537 35383 38546 35417
rect 38494 35374 38546 35383
rect 38654 35417 38706 35426
rect 38654 35383 38663 35417
rect 38663 35383 38697 35417
rect 38697 35383 38706 35417
rect 38654 35374 38706 35383
rect 38814 35417 38866 35426
rect 38814 35383 38823 35417
rect 38823 35383 38857 35417
rect 38857 35383 38866 35417
rect 38814 35374 38866 35383
rect 38974 35417 39026 35426
rect 38974 35383 38983 35417
rect 38983 35383 39017 35417
rect 39017 35383 39026 35417
rect 38974 35374 39026 35383
rect 39134 35417 39186 35426
rect 39134 35383 39143 35417
rect 39143 35383 39177 35417
rect 39177 35383 39186 35417
rect 39134 35374 39186 35383
rect 39294 35417 39346 35426
rect 39294 35383 39303 35417
rect 39303 35383 39337 35417
rect 39337 35383 39346 35417
rect 39294 35374 39346 35383
rect 39454 35417 39506 35426
rect 39454 35383 39463 35417
rect 39463 35383 39497 35417
rect 39497 35383 39506 35417
rect 39454 35374 39506 35383
rect 39614 35417 39666 35426
rect 39614 35383 39623 35417
rect 39623 35383 39657 35417
rect 39657 35383 39666 35417
rect 39614 35374 39666 35383
rect 39774 35417 39826 35426
rect 39774 35383 39783 35417
rect 39783 35383 39817 35417
rect 39817 35383 39826 35417
rect 39774 35374 39826 35383
rect 39934 35417 39986 35426
rect 39934 35383 39943 35417
rect 39943 35383 39977 35417
rect 39977 35383 39986 35417
rect 39934 35374 39986 35383
rect 40094 35417 40146 35426
rect 40094 35383 40103 35417
rect 40103 35383 40137 35417
rect 40137 35383 40146 35417
rect 40094 35374 40146 35383
rect 40254 35417 40306 35426
rect 40254 35383 40263 35417
rect 40263 35383 40297 35417
rect 40297 35383 40306 35417
rect 40254 35374 40306 35383
rect 40414 35417 40466 35426
rect 40414 35383 40423 35417
rect 40423 35383 40457 35417
rect 40457 35383 40466 35417
rect 40414 35374 40466 35383
rect 40574 35417 40626 35426
rect 40574 35383 40583 35417
rect 40583 35383 40617 35417
rect 40617 35383 40626 35417
rect 40574 35374 40626 35383
rect 40734 35417 40786 35426
rect 40734 35383 40743 35417
rect 40743 35383 40777 35417
rect 40777 35383 40786 35417
rect 40734 35374 40786 35383
rect 40894 35417 40946 35426
rect 40894 35383 40903 35417
rect 40903 35383 40937 35417
rect 40937 35383 40946 35417
rect 40894 35374 40946 35383
rect 41054 35417 41106 35426
rect 41054 35383 41063 35417
rect 41063 35383 41097 35417
rect 41097 35383 41106 35417
rect 41054 35374 41106 35383
rect 41214 35417 41266 35426
rect 41214 35383 41223 35417
rect 41223 35383 41257 35417
rect 41257 35383 41266 35417
rect 41214 35374 41266 35383
rect 41374 35417 41426 35426
rect 41374 35383 41383 35417
rect 41383 35383 41417 35417
rect 41417 35383 41426 35417
rect 41374 35374 41426 35383
rect 41534 35417 41586 35426
rect 41534 35383 41543 35417
rect 41543 35383 41577 35417
rect 41577 35383 41586 35417
rect 41534 35374 41586 35383
rect 41694 35417 41746 35426
rect 41694 35383 41703 35417
rect 41703 35383 41737 35417
rect 41737 35383 41746 35417
rect 41694 35374 41746 35383
rect 41854 35417 41906 35426
rect 41854 35383 41863 35417
rect 41863 35383 41897 35417
rect 41897 35383 41906 35417
rect 41854 35374 41906 35383
rect 14 35097 66 35106
rect 14 35063 23 35097
rect 23 35063 57 35097
rect 57 35063 66 35097
rect 14 35054 66 35063
rect 174 35097 226 35106
rect 174 35063 183 35097
rect 183 35063 217 35097
rect 217 35063 226 35097
rect 174 35054 226 35063
rect 334 35097 386 35106
rect 334 35063 343 35097
rect 343 35063 377 35097
rect 377 35063 386 35097
rect 334 35054 386 35063
rect 494 35097 546 35106
rect 494 35063 503 35097
rect 503 35063 537 35097
rect 537 35063 546 35097
rect 494 35054 546 35063
rect 654 35097 706 35106
rect 654 35063 663 35097
rect 663 35063 697 35097
rect 697 35063 706 35097
rect 654 35054 706 35063
rect 814 35097 866 35106
rect 814 35063 823 35097
rect 823 35063 857 35097
rect 857 35063 866 35097
rect 814 35054 866 35063
rect 974 35097 1026 35106
rect 974 35063 983 35097
rect 983 35063 1017 35097
rect 1017 35063 1026 35097
rect 974 35054 1026 35063
rect 1134 35097 1186 35106
rect 1134 35063 1143 35097
rect 1143 35063 1177 35097
rect 1177 35063 1186 35097
rect 1134 35054 1186 35063
rect 1294 35097 1346 35106
rect 1294 35063 1303 35097
rect 1303 35063 1337 35097
rect 1337 35063 1346 35097
rect 1294 35054 1346 35063
rect 1454 35097 1506 35106
rect 1454 35063 1463 35097
rect 1463 35063 1497 35097
rect 1497 35063 1506 35097
rect 1454 35054 1506 35063
rect 1614 35097 1666 35106
rect 1614 35063 1623 35097
rect 1623 35063 1657 35097
rect 1657 35063 1666 35097
rect 1614 35054 1666 35063
rect 1774 35097 1826 35106
rect 1774 35063 1783 35097
rect 1783 35063 1817 35097
rect 1817 35063 1826 35097
rect 1774 35054 1826 35063
rect 1934 35097 1986 35106
rect 1934 35063 1943 35097
rect 1943 35063 1977 35097
rect 1977 35063 1986 35097
rect 1934 35054 1986 35063
rect 2094 35097 2146 35106
rect 2094 35063 2103 35097
rect 2103 35063 2137 35097
rect 2137 35063 2146 35097
rect 2094 35054 2146 35063
rect 2254 35097 2306 35106
rect 2254 35063 2263 35097
rect 2263 35063 2297 35097
rect 2297 35063 2306 35097
rect 2254 35054 2306 35063
rect 2414 35097 2466 35106
rect 2414 35063 2423 35097
rect 2423 35063 2457 35097
rect 2457 35063 2466 35097
rect 2414 35054 2466 35063
rect 2574 35097 2626 35106
rect 2574 35063 2583 35097
rect 2583 35063 2617 35097
rect 2617 35063 2626 35097
rect 2574 35054 2626 35063
rect 2734 35097 2786 35106
rect 2734 35063 2743 35097
rect 2743 35063 2777 35097
rect 2777 35063 2786 35097
rect 2734 35054 2786 35063
rect 2894 35097 2946 35106
rect 2894 35063 2903 35097
rect 2903 35063 2937 35097
rect 2937 35063 2946 35097
rect 2894 35054 2946 35063
rect 3054 35097 3106 35106
rect 3054 35063 3063 35097
rect 3063 35063 3097 35097
rect 3097 35063 3106 35097
rect 3054 35054 3106 35063
rect 3214 35097 3266 35106
rect 3214 35063 3223 35097
rect 3223 35063 3257 35097
rect 3257 35063 3266 35097
rect 3214 35054 3266 35063
rect 3374 35097 3426 35106
rect 3374 35063 3383 35097
rect 3383 35063 3417 35097
rect 3417 35063 3426 35097
rect 3374 35054 3426 35063
rect 3534 35097 3586 35106
rect 3534 35063 3543 35097
rect 3543 35063 3577 35097
rect 3577 35063 3586 35097
rect 3534 35054 3586 35063
rect 3694 35097 3746 35106
rect 3694 35063 3703 35097
rect 3703 35063 3737 35097
rect 3737 35063 3746 35097
rect 3694 35054 3746 35063
rect 3854 35097 3906 35106
rect 3854 35063 3863 35097
rect 3863 35063 3897 35097
rect 3897 35063 3906 35097
rect 3854 35054 3906 35063
rect 4014 35097 4066 35106
rect 4014 35063 4023 35097
rect 4023 35063 4057 35097
rect 4057 35063 4066 35097
rect 4014 35054 4066 35063
rect 4174 35097 4226 35106
rect 4174 35063 4183 35097
rect 4183 35063 4217 35097
rect 4217 35063 4226 35097
rect 4174 35054 4226 35063
rect 4334 35097 4386 35106
rect 4334 35063 4343 35097
rect 4343 35063 4377 35097
rect 4377 35063 4386 35097
rect 4334 35054 4386 35063
rect 4494 35097 4546 35106
rect 4494 35063 4503 35097
rect 4503 35063 4537 35097
rect 4537 35063 4546 35097
rect 4494 35054 4546 35063
rect 4654 35097 4706 35106
rect 4654 35063 4663 35097
rect 4663 35063 4697 35097
rect 4697 35063 4706 35097
rect 4654 35054 4706 35063
rect 4814 35097 4866 35106
rect 4814 35063 4823 35097
rect 4823 35063 4857 35097
rect 4857 35063 4866 35097
rect 4814 35054 4866 35063
rect 4974 35097 5026 35106
rect 4974 35063 4983 35097
rect 4983 35063 5017 35097
rect 5017 35063 5026 35097
rect 4974 35054 5026 35063
rect 5134 35097 5186 35106
rect 5134 35063 5143 35097
rect 5143 35063 5177 35097
rect 5177 35063 5186 35097
rect 5134 35054 5186 35063
rect 5294 35097 5346 35106
rect 5294 35063 5303 35097
rect 5303 35063 5337 35097
rect 5337 35063 5346 35097
rect 5294 35054 5346 35063
rect 5454 35097 5506 35106
rect 5454 35063 5463 35097
rect 5463 35063 5497 35097
rect 5497 35063 5506 35097
rect 5454 35054 5506 35063
rect 5614 35097 5666 35106
rect 5614 35063 5623 35097
rect 5623 35063 5657 35097
rect 5657 35063 5666 35097
rect 5614 35054 5666 35063
rect 5774 35097 5826 35106
rect 5774 35063 5783 35097
rect 5783 35063 5817 35097
rect 5817 35063 5826 35097
rect 5774 35054 5826 35063
rect 5934 35097 5986 35106
rect 5934 35063 5943 35097
rect 5943 35063 5977 35097
rect 5977 35063 5986 35097
rect 5934 35054 5986 35063
rect 6094 35097 6146 35106
rect 6094 35063 6103 35097
rect 6103 35063 6137 35097
rect 6137 35063 6146 35097
rect 6094 35054 6146 35063
rect 6254 35097 6306 35106
rect 6254 35063 6263 35097
rect 6263 35063 6297 35097
rect 6297 35063 6306 35097
rect 6254 35054 6306 35063
rect 6414 35097 6466 35106
rect 6414 35063 6423 35097
rect 6423 35063 6457 35097
rect 6457 35063 6466 35097
rect 6414 35054 6466 35063
rect 6574 35097 6626 35106
rect 6574 35063 6583 35097
rect 6583 35063 6617 35097
rect 6617 35063 6626 35097
rect 6574 35054 6626 35063
rect 6734 35097 6786 35106
rect 6734 35063 6743 35097
rect 6743 35063 6777 35097
rect 6777 35063 6786 35097
rect 6734 35054 6786 35063
rect 6894 35097 6946 35106
rect 6894 35063 6903 35097
rect 6903 35063 6937 35097
rect 6937 35063 6946 35097
rect 6894 35054 6946 35063
rect 7054 35097 7106 35106
rect 7054 35063 7063 35097
rect 7063 35063 7097 35097
rect 7097 35063 7106 35097
rect 7054 35054 7106 35063
rect 7214 35097 7266 35106
rect 7214 35063 7223 35097
rect 7223 35063 7257 35097
rect 7257 35063 7266 35097
rect 7214 35054 7266 35063
rect 7374 35097 7426 35106
rect 7374 35063 7383 35097
rect 7383 35063 7417 35097
rect 7417 35063 7426 35097
rect 7374 35054 7426 35063
rect 7534 35097 7586 35106
rect 7534 35063 7543 35097
rect 7543 35063 7577 35097
rect 7577 35063 7586 35097
rect 7534 35054 7586 35063
rect 7694 35097 7746 35106
rect 7694 35063 7703 35097
rect 7703 35063 7737 35097
rect 7737 35063 7746 35097
rect 7694 35054 7746 35063
rect 7854 35097 7906 35106
rect 7854 35063 7863 35097
rect 7863 35063 7897 35097
rect 7897 35063 7906 35097
rect 7854 35054 7906 35063
rect 8014 35097 8066 35106
rect 8014 35063 8023 35097
rect 8023 35063 8057 35097
rect 8057 35063 8066 35097
rect 8014 35054 8066 35063
rect 8174 35097 8226 35106
rect 8174 35063 8183 35097
rect 8183 35063 8217 35097
rect 8217 35063 8226 35097
rect 8174 35054 8226 35063
rect 8334 35097 8386 35106
rect 8334 35063 8343 35097
rect 8343 35063 8377 35097
rect 8377 35063 8386 35097
rect 8334 35054 8386 35063
rect 12494 35097 12546 35106
rect 12494 35063 12503 35097
rect 12503 35063 12537 35097
rect 12537 35063 12546 35097
rect 12494 35054 12546 35063
rect 12654 35097 12706 35106
rect 12654 35063 12663 35097
rect 12663 35063 12697 35097
rect 12697 35063 12706 35097
rect 12654 35054 12706 35063
rect 12814 35097 12866 35106
rect 12814 35063 12823 35097
rect 12823 35063 12857 35097
rect 12857 35063 12866 35097
rect 12814 35054 12866 35063
rect 12974 35097 13026 35106
rect 12974 35063 12983 35097
rect 12983 35063 13017 35097
rect 13017 35063 13026 35097
rect 12974 35054 13026 35063
rect 13134 35097 13186 35106
rect 13134 35063 13143 35097
rect 13143 35063 13177 35097
rect 13177 35063 13186 35097
rect 13134 35054 13186 35063
rect 13294 35097 13346 35106
rect 13294 35063 13303 35097
rect 13303 35063 13337 35097
rect 13337 35063 13346 35097
rect 13294 35054 13346 35063
rect 13454 35097 13506 35106
rect 13454 35063 13463 35097
rect 13463 35063 13497 35097
rect 13497 35063 13506 35097
rect 13454 35054 13506 35063
rect 13614 35097 13666 35106
rect 13614 35063 13623 35097
rect 13623 35063 13657 35097
rect 13657 35063 13666 35097
rect 13614 35054 13666 35063
rect 13774 35097 13826 35106
rect 13774 35063 13783 35097
rect 13783 35063 13817 35097
rect 13817 35063 13826 35097
rect 13774 35054 13826 35063
rect 13934 35097 13986 35106
rect 13934 35063 13943 35097
rect 13943 35063 13977 35097
rect 13977 35063 13986 35097
rect 13934 35054 13986 35063
rect 14094 35097 14146 35106
rect 14094 35063 14103 35097
rect 14103 35063 14137 35097
rect 14137 35063 14146 35097
rect 14094 35054 14146 35063
rect 14254 35097 14306 35106
rect 14254 35063 14263 35097
rect 14263 35063 14297 35097
rect 14297 35063 14306 35097
rect 14254 35054 14306 35063
rect 14414 35097 14466 35106
rect 14414 35063 14423 35097
rect 14423 35063 14457 35097
rect 14457 35063 14466 35097
rect 14414 35054 14466 35063
rect 14574 35097 14626 35106
rect 14574 35063 14583 35097
rect 14583 35063 14617 35097
rect 14617 35063 14626 35097
rect 14574 35054 14626 35063
rect 14734 35097 14786 35106
rect 14734 35063 14743 35097
rect 14743 35063 14777 35097
rect 14777 35063 14786 35097
rect 14734 35054 14786 35063
rect 14894 35097 14946 35106
rect 14894 35063 14903 35097
rect 14903 35063 14937 35097
rect 14937 35063 14946 35097
rect 14894 35054 14946 35063
rect 15054 35097 15106 35106
rect 15054 35063 15063 35097
rect 15063 35063 15097 35097
rect 15097 35063 15106 35097
rect 15054 35054 15106 35063
rect 15214 35097 15266 35106
rect 15214 35063 15223 35097
rect 15223 35063 15257 35097
rect 15257 35063 15266 35097
rect 15214 35054 15266 35063
rect 15374 35097 15426 35106
rect 15374 35063 15383 35097
rect 15383 35063 15417 35097
rect 15417 35063 15426 35097
rect 15374 35054 15426 35063
rect 15534 35097 15586 35106
rect 15534 35063 15543 35097
rect 15543 35063 15577 35097
rect 15577 35063 15586 35097
rect 15534 35054 15586 35063
rect 15694 35097 15746 35106
rect 15694 35063 15703 35097
rect 15703 35063 15737 35097
rect 15737 35063 15746 35097
rect 15694 35054 15746 35063
rect 15854 35097 15906 35106
rect 15854 35063 15863 35097
rect 15863 35063 15897 35097
rect 15897 35063 15906 35097
rect 15854 35054 15906 35063
rect 16014 35097 16066 35106
rect 16014 35063 16023 35097
rect 16023 35063 16057 35097
rect 16057 35063 16066 35097
rect 16014 35054 16066 35063
rect 16174 35097 16226 35106
rect 16174 35063 16183 35097
rect 16183 35063 16217 35097
rect 16217 35063 16226 35097
rect 16174 35054 16226 35063
rect 16334 35097 16386 35106
rect 16334 35063 16343 35097
rect 16343 35063 16377 35097
rect 16377 35063 16386 35097
rect 16334 35054 16386 35063
rect 16494 35097 16546 35106
rect 16494 35063 16503 35097
rect 16503 35063 16537 35097
rect 16537 35063 16546 35097
rect 16494 35054 16546 35063
rect 16654 35097 16706 35106
rect 16654 35063 16663 35097
rect 16663 35063 16697 35097
rect 16697 35063 16706 35097
rect 16654 35054 16706 35063
rect 16814 35097 16866 35106
rect 16814 35063 16823 35097
rect 16823 35063 16857 35097
rect 16857 35063 16866 35097
rect 16814 35054 16866 35063
rect 16974 35097 17026 35106
rect 16974 35063 16983 35097
rect 16983 35063 17017 35097
rect 17017 35063 17026 35097
rect 16974 35054 17026 35063
rect 17134 35097 17186 35106
rect 17134 35063 17143 35097
rect 17143 35063 17177 35097
rect 17177 35063 17186 35097
rect 17134 35054 17186 35063
rect 17294 35097 17346 35106
rect 17294 35063 17303 35097
rect 17303 35063 17337 35097
rect 17337 35063 17346 35097
rect 17294 35054 17346 35063
rect 17454 35097 17506 35106
rect 17454 35063 17463 35097
rect 17463 35063 17497 35097
rect 17497 35063 17506 35097
rect 17454 35054 17506 35063
rect 17614 35097 17666 35106
rect 17614 35063 17623 35097
rect 17623 35063 17657 35097
rect 17657 35063 17666 35097
rect 17614 35054 17666 35063
rect 17774 35097 17826 35106
rect 17774 35063 17783 35097
rect 17783 35063 17817 35097
rect 17817 35063 17826 35097
rect 17774 35054 17826 35063
rect 17934 35097 17986 35106
rect 17934 35063 17943 35097
rect 17943 35063 17977 35097
rect 17977 35063 17986 35097
rect 17934 35054 17986 35063
rect 18094 35097 18146 35106
rect 18094 35063 18103 35097
rect 18103 35063 18137 35097
rect 18137 35063 18146 35097
rect 18094 35054 18146 35063
rect 18254 35097 18306 35106
rect 18254 35063 18263 35097
rect 18263 35063 18297 35097
rect 18297 35063 18306 35097
rect 18254 35054 18306 35063
rect 18414 35097 18466 35106
rect 18414 35063 18423 35097
rect 18423 35063 18457 35097
rect 18457 35063 18466 35097
rect 18414 35054 18466 35063
rect 18574 35097 18626 35106
rect 18574 35063 18583 35097
rect 18583 35063 18617 35097
rect 18617 35063 18626 35097
rect 18574 35054 18626 35063
rect 18734 35097 18786 35106
rect 18734 35063 18743 35097
rect 18743 35063 18777 35097
rect 18777 35063 18786 35097
rect 18734 35054 18786 35063
rect 18894 35097 18946 35106
rect 18894 35063 18903 35097
rect 18903 35063 18937 35097
rect 18937 35063 18946 35097
rect 18894 35054 18946 35063
rect 23134 35097 23186 35106
rect 23134 35063 23143 35097
rect 23143 35063 23177 35097
rect 23177 35063 23186 35097
rect 23134 35054 23186 35063
rect 23294 35097 23346 35106
rect 23294 35063 23303 35097
rect 23303 35063 23337 35097
rect 23337 35063 23346 35097
rect 23294 35054 23346 35063
rect 23454 35097 23506 35106
rect 23454 35063 23463 35097
rect 23463 35063 23497 35097
rect 23497 35063 23506 35097
rect 23454 35054 23506 35063
rect 23614 35097 23666 35106
rect 23614 35063 23623 35097
rect 23623 35063 23657 35097
rect 23657 35063 23666 35097
rect 23614 35054 23666 35063
rect 23774 35097 23826 35106
rect 23774 35063 23783 35097
rect 23783 35063 23817 35097
rect 23817 35063 23826 35097
rect 23774 35054 23826 35063
rect 23934 35097 23986 35106
rect 23934 35063 23943 35097
rect 23943 35063 23977 35097
rect 23977 35063 23986 35097
rect 23934 35054 23986 35063
rect 24094 35097 24146 35106
rect 24094 35063 24103 35097
rect 24103 35063 24137 35097
rect 24137 35063 24146 35097
rect 24094 35054 24146 35063
rect 24254 35097 24306 35106
rect 24254 35063 24263 35097
rect 24263 35063 24297 35097
rect 24297 35063 24306 35097
rect 24254 35054 24306 35063
rect 24414 35097 24466 35106
rect 24414 35063 24423 35097
rect 24423 35063 24457 35097
rect 24457 35063 24466 35097
rect 24414 35054 24466 35063
rect 24574 35097 24626 35106
rect 24574 35063 24583 35097
rect 24583 35063 24617 35097
rect 24617 35063 24626 35097
rect 24574 35054 24626 35063
rect 24734 35097 24786 35106
rect 24734 35063 24743 35097
rect 24743 35063 24777 35097
rect 24777 35063 24786 35097
rect 24734 35054 24786 35063
rect 24894 35097 24946 35106
rect 24894 35063 24903 35097
rect 24903 35063 24937 35097
rect 24937 35063 24946 35097
rect 24894 35054 24946 35063
rect 25054 35097 25106 35106
rect 25054 35063 25063 35097
rect 25063 35063 25097 35097
rect 25097 35063 25106 35097
rect 25054 35054 25106 35063
rect 25214 35097 25266 35106
rect 25214 35063 25223 35097
rect 25223 35063 25257 35097
rect 25257 35063 25266 35097
rect 25214 35054 25266 35063
rect 25374 35097 25426 35106
rect 25374 35063 25383 35097
rect 25383 35063 25417 35097
rect 25417 35063 25426 35097
rect 25374 35054 25426 35063
rect 25534 35097 25586 35106
rect 25534 35063 25543 35097
rect 25543 35063 25577 35097
rect 25577 35063 25586 35097
rect 25534 35054 25586 35063
rect 25694 35097 25746 35106
rect 25694 35063 25703 35097
rect 25703 35063 25737 35097
rect 25737 35063 25746 35097
rect 25694 35054 25746 35063
rect 25854 35097 25906 35106
rect 25854 35063 25863 35097
rect 25863 35063 25897 35097
rect 25897 35063 25906 35097
rect 25854 35054 25906 35063
rect 26014 35097 26066 35106
rect 26014 35063 26023 35097
rect 26023 35063 26057 35097
rect 26057 35063 26066 35097
rect 26014 35054 26066 35063
rect 26174 35097 26226 35106
rect 26174 35063 26183 35097
rect 26183 35063 26217 35097
rect 26217 35063 26226 35097
rect 26174 35054 26226 35063
rect 26334 35097 26386 35106
rect 26334 35063 26343 35097
rect 26343 35063 26377 35097
rect 26377 35063 26386 35097
rect 26334 35054 26386 35063
rect 26494 35097 26546 35106
rect 26494 35063 26503 35097
rect 26503 35063 26537 35097
rect 26537 35063 26546 35097
rect 26494 35054 26546 35063
rect 26654 35097 26706 35106
rect 26654 35063 26663 35097
rect 26663 35063 26697 35097
rect 26697 35063 26706 35097
rect 26654 35054 26706 35063
rect 26814 35097 26866 35106
rect 26814 35063 26823 35097
rect 26823 35063 26857 35097
rect 26857 35063 26866 35097
rect 26814 35054 26866 35063
rect 26974 35097 27026 35106
rect 26974 35063 26983 35097
rect 26983 35063 27017 35097
rect 27017 35063 27026 35097
rect 26974 35054 27026 35063
rect 27134 35097 27186 35106
rect 27134 35063 27143 35097
rect 27143 35063 27177 35097
rect 27177 35063 27186 35097
rect 27134 35054 27186 35063
rect 27294 35097 27346 35106
rect 27294 35063 27303 35097
rect 27303 35063 27337 35097
rect 27337 35063 27346 35097
rect 27294 35054 27346 35063
rect 27454 35097 27506 35106
rect 27454 35063 27463 35097
rect 27463 35063 27497 35097
rect 27497 35063 27506 35097
rect 27454 35054 27506 35063
rect 27614 35097 27666 35106
rect 27614 35063 27623 35097
rect 27623 35063 27657 35097
rect 27657 35063 27666 35097
rect 27614 35054 27666 35063
rect 27774 35097 27826 35106
rect 27774 35063 27783 35097
rect 27783 35063 27817 35097
rect 27817 35063 27826 35097
rect 27774 35054 27826 35063
rect 27934 35097 27986 35106
rect 27934 35063 27943 35097
rect 27943 35063 27977 35097
rect 27977 35063 27986 35097
rect 27934 35054 27986 35063
rect 28094 35097 28146 35106
rect 28094 35063 28103 35097
rect 28103 35063 28137 35097
rect 28137 35063 28146 35097
rect 28094 35054 28146 35063
rect 28254 35097 28306 35106
rect 28254 35063 28263 35097
rect 28263 35063 28297 35097
rect 28297 35063 28306 35097
rect 28254 35054 28306 35063
rect 28414 35097 28466 35106
rect 28414 35063 28423 35097
rect 28423 35063 28457 35097
rect 28457 35063 28466 35097
rect 28414 35054 28466 35063
rect 28574 35097 28626 35106
rect 28574 35063 28583 35097
rect 28583 35063 28617 35097
rect 28617 35063 28626 35097
rect 28574 35054 28626 35063
rect 28734 35097 28786 35106
rect 28734 35063 28743 35097
rect 28743 35063 28777 35097
rect 28777 35063 28786 35097
rect 28734 35054 28786 35063
rect 28894 35097 28946 35106
rect 28894 35063 28903 35097
rect 28903 35063 28937 35097
rect 28937 35063 28946 35097
rect 28894 35054 28946 35063
rect 29054 35097 29106 35106
rect 29054 35063 29063 35097
rect 29063 35063 29097 35097
rect 29097 35063 29106 35097
rect 29054 35054 29106 35063
rect 29214 35097 29266 35106
rect 29214 35063 29223 35097
rect 29223 35063 29257 35097
rect 29257 35063 29266 35097
rect 29214 35054 29266 35063
rect 29374 35097 29426 35106
rect 29374 35063 29383 35097
rect 29383 35063 29417 35097
rect 29417 35063 29426 35097
rect 29374 35054 29426 35063
rect 33534 35097 33586 35106
rect 33534 35063 33543 35097
rect 33543 35063 33577 35097
rect 33577 35063 33586 35097
rect 33534 35054 33586 35063
rect 33694 35097 33746 35106
rect 33694 35063 33703 35097
rect 33703 35063 33737 35097
rect 33737 35063 33746 35097
rect 33694 35054 33746 35063
rect 33854 35097 33906 35106
rect 33854 35063 33863 35097
rect 33863 35063 33897 35097
rect 33897 35063 33906 35097
rect 33854 35054 33906 35063
rect 34014 35097 34066 35106
rect 34014 35063 34023 35097
rect 34023 35063 34057 35097
rect 34057 35063 34066 35097
rect 34014 35054 34066 35063
rect 34174 35097 34226 35106
rect 34174 35063 34183 35097
rect 34183 35063 34217 35097
rect 34217 35063 34226 35097
rect 34174 35054 34226 35063
rect 34334 35097 34386 35106
rect 34334 35063 34343 35097
rect 34343 35063 34377 35097
rect 34377 35063 34386 35097
rect 34334 35054 34386 35063
rect 34494 35097 34546 35106
rect 34494 35063 34503 35097
rect 34503 35063 34537 35097
rect 34537 35063 34546 35097
rect 34494 35054 34546 35063
rect 34654 35097 34706 35106
rect 34654 35063 34663 35097
rect 34663 35063 34697 35097
rect 34697 35063 34706 35097
rect 34654 35054 34706 35063
rect 34814 35097 34866 35106
rect 34814 35063 34823 35097
rect 34823 35063 34857 35097
rect 34857 35063 34866 35097
rect 34814 35054 34866 35063
rect 34974 35097 35026 35106
rect 34974 35063 34983 35097
rect 34983 35063 35017 35097
rect 35017 35063 35026 35097
rect 34974 35054 35026 35063
rect 35134 35097 35186 35106
rect 35134 35063 35143 35097
rect 35143 35063 35177 35097
rect 35177 35063 35186 35097
rect 35134 35054 35186 35063
rect 35294 35097 35346 35106
rect 35294 35063 35303 35097
rect 35303 35063 35337 35097
rect 35337 35063 35346 35097
rect 35294 35054 35346 35063
rect 35454 35097 35506 35106
rect 35454 35063 35463 35097
rect 35463 35063 35497 35097
rect 35497 35063 35506 35097
rect 35454 35054 35506 35063
rect 35614 35097 35666 35106
rect 35614 35063 35623 35097
rect 35623 35063 35657 35097
rect 35657 35063 35666 35097
rect 35614 35054 35666 35063
rect 35774 35097 35826 35106
rect 35774 35063 35783 35097
rect 35783 35063 35817 35097
rect 35817 35063 35826 35097
rect 35774 35054 35826 35063
rect 35934 35097 35986 35106
rect 35934 35063 35943 35097
rect 35943 35063 35977 35097
rect 35977 35063 35986 35097
rect 35934 35054 35986 35063
rect 36094 35097 36146 35106
rect 36094 35063 36103 35097
rect 36103 35063 36137 35097
rect 36137 35063 36146 35097
rect 36094 35054 36146 35063
rect 36254 35097 36306 35106
rect 36254 35063 36263 35097
rect 36263 35063 36297 35097
rect 36297 35063 36306 35097
rect 36254 35054 36306 35063
rect 36414 35097 36466 35106
rect 36414 35063 36423 35097
rect 36423 35063 36457 35097
rect 36457 35063 36466 35097
rect 36414 35054 36466 35063
rect 36574 35097 36626 35106
rect 36574 35063 36583 35097
rect 36583 35063 36617 35097
rect 36617 35063 36626 35097
rect 36574 35054 36626 35063
rect 36734 35097 36786 35106
rect 36734 35063 36743 35097
rect 36743 35063 36777 35097
rect 36777 35063 36786 35097
rect 36734 35054 36786 35063
rect 36894 35097 36946 35106
rect 36894 35063 36903 35097
rect 36903 35063 36937 35097
rect 36937 35063 36946 35097
rect 36894 35054 36946 35063
rect 37054 35097 37106 35106
rect 37054 35063 37063 35097
rect 37063 35063 37097 35097
rect 37097 35063 37106 35097
rect 37054 35054 37106 35063
rect 37214 35097 37266 35106
rect 37214 35063 37223 35097
rect 37223 35063 37257 35097
rect 37257 35063 37266 35097
rect 37214 35054 37266 35063
rect 37374 35097 37426 35106
rect 37374 35063 37383 35097
rect 37383 35063 37417 35097
rect 37417 35063 37426 35097
rect 37374 35054 37426 35063
rect 37534 35097 37586 35106
rect 37534 35063 37543 35097
rect 37543 35063 37577 35097
rect 37577 35063 37586 35097
rect 37534 35054 37586 35063
rect 37694 35097 37746 35106
rect 37694 35063 37703 35097
rect 37703 35063 37737 35097
rect 37737 35063 37746 35097
rect 37694 35054 37746 35063
rect 37854 35097 37906 35106
rect 37854 35063 37863 35097
rect 37863 35063 37897 35097
rect 37897 35063 37906 35097
rect 37854 35054 37906 35063
rect 38014 35097 38066 35106
rect 38014 35063 38023 35097
rect 38023 35063 38057 35097
rect 38057 35063 38066 35097
rect 38014 35054 38066 35063
rect 38174 35097 38226 35106
rect 38174 35063 38183 35097
rect 38183 35063 38217 35097
rect 38217 35063 38226 35097
rect 38174 35054 38226 35063
rect 38334 35097 38386 35106
rect 38334 35063 38343 35097
rect 38343 35063 38377 35097
rect 38377 35063 38386 35097
rect 38334 35054 38386 35063
rect 38494 35097 38546 35106
rect 38494 35063 38503 35097
rect 38503 35063 38537 35097
rect 38537 35063 38546 35097
rect 38494 35054 38546 35063
rect 38654 35097 38706 35106
rect 38654 35063 38663 35097
rect 38663 35063 38697 35097
rect 38697 35063 38706 35097
rect 38654 35054 38706 35063
rect 38814 35097 38866 35106
rect 38814 35063 38823 35097
rect 38823 35063 38857 35097
rect 38857 35063 38866 35097
rect 38814 35054 38866 35063
rect 38974 35097 39026 35106
rect 38974 35063 38983 35097
rect 38983 35063 39017 35097
rect 39017 35063 39026 35097
rect 38974 35054 39026 35063
rect 39134 35097 39186 35106
rect 39134 35063 39143 35097
rect 39143 35063 39177 35097
rect 39177 35063 39186 35097
rect 39134 35054 39186 35063
rect 39294 35097 39346 35106
rect 39294 35063 39303 35097
rect 39303 35063 39337 35097
rect 39337 35063 39346 35097
rect 39294 35054 39346 35063
rect 39454 35097 39506 35106
rect 39454 35063 39463 35097
rect 39463 35063 39497 35097
rect 39497 35063 39506 35097
rect 39454 35054 39506 35063
rect 39614 35097 39666 35106
rect 39614 35063 39623 35097
rect 39623 35063 39657 35097
rect 39657 35063 39666 35097
rect 39614 35054 39666 35063
rect 39774 35097 39826 35106
rect 39774 35063 39783 35097
rect 39783 35063 39817 35097
rect 39817 35063 39826 35097
rect 39774 35054 39826 35063
rect 39934 35097 39986 35106
rect 39934 35063 39943 35097
rect 39943 35063 39977 35097
rect 39977 35063 39986 35097
rect 39934 35054 39986 35063
rect 40094 35097 40146 35106
rect 40094 35063 40103 35097
rect 40103 35063 40137 35097
rect 40137 35063 40146 35097
rect 40094 35054 40146 35063
rect 40254 35097 40306 35106
rect 40254 35063 40263 35097
rect 40263 35063 40297 35097
rect 40297 35063 40306 35097
rect 40254 35054 40306 35063
rect 40414 35097 40466 35106
rect 40414 35063 40423 35097
rect 40423 35063 40457 35097
rect 40457 35063 40466 35097
rect 40414 35054 40466 35063
rect 40574 35097 40626 35106
rect 40574 35063 40583 35097
rect 40583 35063 40617 35097
rect 40617 35063 40626 35097
rect 40574 35054 40626 35063
rect 40734 35097 40786 35106
rect 40734 35063 40743 35097
rect 40743 35063 40777 35097
rect 40777 35063 40786 35097
rect 40734 35054 40786 35063
rect 40894 35097 40946 35106
rect 40894 35063 40903 35097
rect 40903 35063 40937 35097
rect 40937 35063 40946 35097
rect 40894 35054 40946 35063
rect 41054 35097 41106 35106
rect 41054 35063 41063 35097
rect 41063 35063 41097 35097
rect 41097 35063 41106 35097
rect 41054 35054 41106 35063
rect 41214 35097 41266 35106
rect 41214 35063 41223 35097
rect 41223 35063 41257 35097
rect 41257 35063 41266 35097
rect 41214 35054 41266 35063
rect 41374 35097 41426 35106
rect 41374 35063 41383 35097
rect 41383 35063 41417 35097
rect 41417 35063 41426 35097
rect 41374 35054 41426 35063
rect 41534 35097 41586 35106
rect 41534 35063 41543 35097
rect 41543 35063 41577 35097
rect 41577 35063 41586 35097
rect 41534 35054 41586 35063
rect 41694 35097 41746 35106
rect 41694 35063 41703 35097
rect 41703 35063 41737 35097
rect 41737 35063 41746 35097
rect 41694 35054 41746 35063
rect 41854 35097 41906 35106
rect 41854 35063 41863 35097
rect 41863 35063 41897 35097
rect 41897 35063 41906 35097
rect 41854 35054 41906 35063
rect 14 34777 66 34786
rect 14 34743 23 34777
rect 23 34743 57 34777
rect 57 34743 66 34777
rect 14 34734 66 34743
rect 174 34777 226 34786
rect 174 34743 183 34777
rect 183 34743 217 34777
rect 217 34743 226 34777
rect 174 34734 226 34743
rect 334 34777 386 34786
rect 334 34743 343 34777
rect 343 34743 377 34777
rect 377 34743 386 34777
rect 334 34734 386 34743
rect 494 34777 546 34786
rect 494 34743 503 34777
rect 503 34743 537 34777
rect 537 34743 546 34777
rect 494 34734 546 34743
rect 654 34777 706 34786
rect 654 34743 663 34777
rect 663 34743 697 34777
rect 697 34743 706 34777
rect 654 34734 706 34743
rect 814 34777 866 34786
rect 814 34743 823 34777
rect 823 34743 857 34777
rect 857 34743 866 34777
rect 814 34734 866 34743
rect 974 34777 1026 34786
rect 974 34743 983 34777
rect 983 34743 1017 34777
rect 1017 34743 1026 34777
rect 974 34734 1026 34743
rect 1134 34777 1186 34786
rect 1134 34743 1143 34777
rect 1143 34743 1177 34777
rect 1177 34743 1186 34777
rect 1134 34734 1186 34743
rect 1294 34777 1346 34786
rect 1294 34743 1303 34777
rect 1303 34743 1337 34777
rect 1337 34743 1346 34777
rect 1294 34734 1346 34743
rect 1454 34777 1506 34786
rect 1454 34743 1463 34777
rect 1463 34743 1497 34777
rect 1497 34743 1506 34777
rect 1454 34734 1506 34743
rect 1614 34777 1666 34786
rect 1614 34743 1623 34777
rect 1623 34743 1657 34777
rect 1657 34743 1666 34777
rect 1614 34734 1666 34743
rect 1774 34777 1826 34786
rect 1774 34743 1783 34777
rect 1783 34743 1817 34777
rect 1817 34743 1826 34777
rect 1774 34734 1826 34743
rect 1934 34777 1986 34786
rect 1934 34743 1943 34777
rect 1943 34743 1977 34777
rect 1977 34743 1986 34777
rect 1934 34734 1986 34743
rect 2094 34777 2146 34786
rect 2094 34743 2103 34777
rect 2103 34743 2137 34777
rect 2137 34743 2146 34777
rect 2094 34734 2146 34743
rect 2254 34777 2306 34786
rect 2254 34743 2263 34777
rect 2263 34743 2297 34777
rect 2297 34743 2306 34777
rect 2254 34734 2306 34743
rect 2414 34777 2466 34786
rect 2414 34743 2423 34777
rect 2423 34743 2457 34777
rect 2457 34743 2466 34777
rect 2414 34734 2466 34743
rect 2574 34777 2626 34786
rect 2574 34743 2583 34777
rect 2583 34743 2617 34777
rect 2617 34743 2626 34777
rect 2574 34734 2626 34743
rect 2734 34777 2786 34786
rect 2734 34743 2743 34777
rect 2743 34743 2777 34777
rect 2777 34743 2786 34777
rect 2734 34734 2786 34743
rect 2894 34777 2946 34786
rect 2894 34743 2903 34777
rect 2903 34743 2937 34777
rect 2937 34743 2946 34777
rect 2894 34734 2946 34743
rect 3054 34777 3106 34786
rect 3054 34743 3063 34777
rect 3063 34743 3097 34777
rect 3097 34743 3106 34777
rect 3054 34734 3106 34743
rect 3214 34777 3266 34786
rect 3214 34743 3223 34777
rect 3223 34743 3257 34777
rect 3257 34743 3266 34777
rect 3214 34734 3266 34743
rect 3374 34777 3426 34786
rect 3374 34743 3383 34777
rect 3383 34743 3417 34777
rect 3417 34743 3426 34777
rect 3374 34734 3426 34743
rect 3534 34777 3586 34786
rect 3534 34743 3543 34777
rect 3543 34743 3577 34777
rect 3577 34743 3586 34777
rect 3534 34734 3586 34743
rect 3694 34777 3746 34786
rect 3694 34743 3703 34777
rect 3703 34743 3737 34777
rect 3737 34743 3746 34777
rect 3694 34734 3746 34743
rect 3854 34777 3906 34786
rect 3854 34743 3863 34777
rect 3863 34743 3897 34777
rect 3897 34743 3906 34777
rect 3854 34734 3906 34743
rect 4014 34777 4066 34786
rect 4014 34743 4023 34777
rect 4023 34743 4057 34777
rect 4057 34743 4066 34777
rect 4014 34734 4066 34743
rect 4174 34777 4226 34786
rect 4174 34743 4183 34777
rect 4183 34743 4217 34777
rect 4217 34743 4226 34777
rect 4174 34734 4226 34743
rect 4334 34777 4386 34786
rect 4334 34743 4343 34777
rect 4343 34743 4377 34777
rect 4377 34743 4386 34777
rect 4334 34734 4386 34743
rect 4494 34777 4546 34786
rect 4494 34743 4503 34777
rect 4503 34743 4537 34777
rect 4537 34743 4546 34777
rect 4494 34734 4546 34743
rect 4654 34777 4706 34786
rect 4654 34743 4663 34777
rect 4663 34743 4697 34777
rect 4697 34743 4706 34777
rect 4654 34734 4706 34743
rect 4814 34777 4866 34786
rect 4814 34743 4823 34777
rect 4823 34743 4857 34777
rect 4857 34743 4866 34777
rect 4814 34734 4866 34743
rect 4974 34777 5026 34786
rect 4974 34743 4983 34777
rect 4983 34743 5017 34777
rect 5017 34743 5026 34777
rect 4974 34734 5026 34743
rect 5134 34777 5186 34786
rect 5134 34743 5143 34777
rect 5143 34743 5177 34777
rect 5177 34743 5186 34777
rect 5134 34734 5186 34743
rect 5294 34777 5346 34786
rect 5294 34743 5303 34777
rect 5303 34743 5337 34777
rect 5337 34743 5346 34777
rect 5294 34734 5346 34743
rect 5454 34777 5506 34786
rect 5454 34743 5463 34777
rect 5463 34743 5497 34777
rect 5497 34743 5506 34777
rect 5454 34734 5506 34743
rect 5614 34777 5666 34786
rect 5614 34743 5623 34777
rect 5623 34743 5657 34777
rect 5657 34743 5666 34777
rect 5614 34734 5666 34743
rect 5774 34777 5826 34786
rect 5774 34743 5783 34777
rect 5783 34743 5817 34777
rect 5817 34743 5826 34777
rect 5774 34734 5826 34743
rect 5934 34777 5986 34786
rect 5934 34743 5943 34777
rect 5943 34743 5977 34777
rect 5977 34743 5986 34777
rect 5934 34734 5986 34743
rect 6094 34777 6146 34786
rect 6094 34743 6103 34777
rect 6103 34743 6137 34777
rect 6137 34743 6146 34777
rect 6094 34734 6146 34743
rect 6254 34777 6306 34786
rect 6254 34743 6263 34777
rect 6263 34743 6297 34777
rect 6297 34743 6306 34777
rect 6254 34734 6306 34743
rect 6414 34777 6466 34786
rect 6414 34743 6423 34777
rect 6423 34743 6457 34777
rect 6457 34743 6466 34777
rect 6414 34734 6466 34743
rect 6574 34777 6626 34786
rect 6574 34743 6583 34777
rect 6583 34743 6617 34777
rect 6617 34743 6626 34777
rect 6574 34734 6626 34743
rect 6734 34777 6786 34786
rect 6734 34743 6743 34777
rect 6743 34743 6777 34777
rect 6777 34743 6786 34777
rect 6734 34734 6786 34743
rect 6894 34777 6946 34786
rect 6894 34743 6903 34777
rect 6903 34743 6937 34777
rect 6937 34743 6946 34777
rect 6894 34734 6946 34743
rect 7054 34777 7106 34786
rect 7054 34743 7063 34777
rect 7063 34743 7097 34777
rect 7097 34743 7106 34777
rect 7054 34734 7106 34743
rect 7214 34777 7266 34786
rect 7214 34743 7223 34777
rect 7223 34743 7257 34777
rect 7257 34743 7266 34777
rect 7214 34734 7266 34743
rect 7374 34777 7426 34786
rect 7374 34743 7383 34777
rect 7383 34743 7417 34777
rect 7417 34743 7426 34777
rect 7374 34734 7426 34743
rect 7534 34777 7586 34786
rect 7534 34743 7543 34777
rect 7543 34743 7577 34777
rect 7577 34743 7586 34777
rect 7534 34734 7586 34743
rect 7694 34777 7746 34786
rect 7694 34743 7703 34777
rect 7703 34743 7737 34777
rect 7737 34743 7746 34777
rect 7694 34734 7746 34743
rect 7854 34777 7906 34786
rect 7854 34743 7863 34777
rect 7863 34743 7897 34777
rect 7897 34743 7906 34777
rect 7854 34734 7906 34743
rect 8014 34777 8066 34786
rect 8014 34743 8023 34777
rect 8023 34743 8057 34777
rect 8057 34743 8066 34777
rect 8014 34734 8066 34743
rect 8174 34777 8226 34786
rect 8174 34743 8183 34777
rect 8183 34743 8217 34777
rect 8217 34743 8226 34777
rect 8174 34734 8226 34743
rect 8334 34777 8386 34786
rect 8334 34743 8343 34777
rect 8343 34743 8377 34777
rect 8377 34743 8386 34777
rect 8334 34734 8386 34743
rect 12494 34777 12546 34786
rect 12494 34743 12503 34777
rect 12503 34743 12537 34777
rect 12537 34743 12546 34777
rect 12494 34734 12546 34743
rect 12654 34777 12706 34786
rect 12654 34743 12663 34777
rect 12663 34743 12697 34777
rect 12697 34743 12706 34777
rect 12654 34734 12706 34743
rect 12814 34777 12866 34786
rect 12814 34743 12823 34777
rect 12823 34743 12857 34777
rect 12857 34743 12866 34777
rect 12814 34734 12866 34743
rect 12974 34777 13026 34786
rect 12974 34743 12983 34777
rect 12983 34743 13017 34777
rect 13017 34743 13026 34777
rect 12974 34734 13026 34743
rect 13134 34777 13186 34786
rect 13134 34743 13143 34777
rect 13143 34743 13177 34777
rect 13177 34743 13186 34777
rect 13134 34734 13186 34743
rect 13294 34777 13346 34786
rect 13294 34743 13303 34777
rect 13303 34743 13337 34777
rect 13337 34743 13346 34777
rect 13294 34734 13346 34743
rect 13454 34777 13506 34786
rect 13454 34743 13463 34777
rect 13463 34743 13497 34777
rect 13497 34743 13506 34777
rect 13454 34734 13506 34743
rect 13614 34777 13666 34786
rect 13614 34743 13623 34777
rect 13623 34743 13657 34777
rect 13657 34743 13666 34777
rect 13614 34734 13666 34743
rect 13774 34777 13826 34786
rect 13774 34743 13783 34777
rect 13783 34743 13817 34777
rect 13817 34743 13826 34777
rect 13774 34734 13826 34743
rect 13934 34777 13986 34786
rect 13934 34743 13943 34777
rect 13943 34743 13977 34777
rect 13977 34743 13986 34777
rect 13934 34734 13986 34743
rect 14094 34777 14146 34786
rect 14094 34743 14103 34777
rect 14103 34743 14137 34777
rect 14137 34743 14146 34777
rect 14094 34734 14146 34743
rect 14254 34777 14306 34786
rect 14254 34743 14263 34777
rect 14263 34743 14297 34777
rect 14297 34743 14306 34777
rect 14254 34734 14306 34743
rect 14414 34777 14466 34786
rect 14414 34743 14423 34777
rect 14423 34743 14457 34777
rect 14457 34743 14466 34777
rect 14414 34734 14466 34743
rect 14574 34777 14626 34786
rect 14574 34743 14583 34777
rect 14583 34743 14617 34777
rect 14617 34743 14626 34777
rect 14574 34734 14626 34743
rect 14734 34777 14786 34786
rect 14734 34743 14743 34777
rect 14743 34743 14777 34777
rect 14777 34743 14786 34777
rect 14734 34734 14786 34743
rect 14894 34777 14946 34786
rect 14894 34743 14903 34777
rect 14903 34743 14937 34777
rect 14937 34743 14946 34777
rect 14894 34734 14946 34743
rect 15054 34777 15106 34786
rect 15054 34743 15063 34777
rect 15063 34743 15097 34777
rect 15097 34743 15106 34777
rect 15054 34734 15106 34743
rect 15214 34777 15266 34786
rect 15214 34743 15223 34777
rect 15223 34743 15257 34777
rect 15257 34743 15266 34777
rect 15214 34734 15266 34743
rect 15374 34777 15426 34786
rect 15374 34743 15383 34777
rect 15383 34743 15417 34777
rect 15417 34743 15426 34777
rect 15374 34734 15426 34743
rect 15534 34777 15586 34786
rect 15534 34743 15543 34777
rect 15543 34743 15577 34777
rect 15577 34743 15586 34777
rect 15534 34734 15586 34743
rect 15694 34777 15746 34786
rect 15694 34743 15703 34777
rect 15703 34743 15737 34777
rect 15737 34743 15746 34777
rect 15694 34734 15746 34743
rect 15854 34777 15906 34786
rect 15854 34743 15863 34777
rect 15863 34743 15897 34777
rect 15897 34743 15906 34777
rect 15854 34734 15906 34743
rect 16014 34777 16066 34786
rect 16014 34743 16023 34777
rect 16023 34743 16057 34777
rect 16057 34743 16066 34777
rect 16014 34734 16066 34743
rect 16174 34777 16226 34786
rect 16174 34743 16183 34777
rect 16183 34743 16217 34777
rect 16217 34743 16226 34777
rect 16174 34734 16226 34743
rect 16334 34777 16386 34786
rect 16334 34743 16343 34777
rect 16343 34743 16377 34777
rect 16377 34743 16386 34777
rect 16334 34734 16386 34743
rect 16494 34777 16546 34786
rect 16494 34743 16503 34777
rect 16503 34743 16537 34777
rect 16537 34743 16546 34777
rect 16494 34734 16546 34743
rect 16654 34777 16706 34786
rect 16654 34743 16663 34777
rect 16663 34743 16697 34777
rect 16697 34743 16706 34777
rect 16654 34734 16706 34743
rect 16814 34777 16866 34786
rect 16814 34743 16823 34777
rect 16823 34743 16857 34777
rect 16857 34743 16866 34777
rect 16814 34734 16866 34743
rect 16974 34777 17026 34786
rect 16974 34743 16983 34777
rect 16983 34743 17017 34777
rect 17017 34743 17026 34777
rect 16974 34734 17026 34743
rect 17134 34777 17186 34786
rect 17134 34743 17143 34777
rect 17143 34743 17177 34777
rect 17177 34743 17186 34777
rect 17134 34734 17186 34743
rect 17294 34777 17346 34786
rect 17294 34743 17303 34777
rect 17303 34743 17337 34777
rect 17337 34743 17346 34777
rect 17294 34734 17346 34743
rect 17454 34777 17506 34786
rect 17454 34743 17463 34777
rect 17463 34743 17497 34777
rect 17497 34743 17506 34777
rect 17454 34734 17506 34743
rect 17614 34777 17666 34786
rect 17614 34743 17623 34777
rect 17623 34743 17657 34777
rect 17657 34743 17666 34777
rect 17614 34734 17666 34743
rect 17774 34777 17826 34786
rect 17774 34743 17783 34777
rect 17783 34743 17817 34777
rect 17817 34743 17826 34777
rect 17774 34734 17826 34743
rect 17934 34777 17986 34786
rect 17934 34743 17943 34777
rect 17943 34743 17977 34777
rect 17977 34743 17986 34777
rect 17934 34734 17986 34743
rect 18094 34777 18146 34786
rect 18094 34743 18103 34777
rect 18103 34743 18137 34777
rect 18137 34743 18146 34777
rect 18094 34734 18146 34743
rect 18254 34777 18306 34786
rect 18254 34743 18263 34777
rect 18263 34743 18297 34777
rect 18297 34743 18306 34777
rect 18254 34734 18306 34743
rect 18414 34777 18466 34786
rect 18414 34743 18423 34777
rect 18423 34743 18457 34777
rect 18457 34743 18466 34777
rect 18414 34734 18466 34743
rect 18574 34777 18626 34786
rect 18574 34743 18583 34777
rect 18583 34743 18617 34777
rect 18617 34743 18626 34777
rect 18574 34734 18626 34743
rect 18734 34777 18786 34786
rect 18734 34743 18743 34777
rect 18743 34743 18777 34777
rect 18777 34743 18786 34777
rect 18734 34734 18786 34743
rect 18894 34777 18946 34786
rect 18894 34743 18903 34777
rect 18903 34743 18937 34777
rect 18937 34743 18946 34777
rect 18894 34734 18946 34743
rect 23134 34777 23186 34786
rect 23134 34743 23143 34777
rect 23143 34743 23177 34777
rect 23177 34743 23186 34777
rect 23134 34734 23186 34743
rect 23294 34777 23346 34786
rect 23294 34743 23303 34777
rect 23303 34743 23337 34777
rect 23337 34743 23346 34777
rect 23294 34734 23346 34743
rect 23454 34777 23506 34786
rect 23454 34743 23463 34777
rect 23463 34743 23497 34777
rect 23497 34743 23506 34777
rect 23454 34734 23506 34743
rect 23614 34777 23666 34786
rect 23614 34743 23623 34777
rect 23623 34743 23657 34777
rect 23657 34743 23666 34777
rect 23614 34734 23666 34743
rect 23774 34777 23826 34786
rect 23774 34743 23783 34777
rect 23783 34743 23817 34777
rect 23817 34743 23826 34777
rect 23774 34734 23826 34743
rect 23934 34777 23986 34786
rect 23934 34743 23943 34777
rect 23943 34743 23977 34777
rect 23977 34743 23986 34777
rect 23934 34734 23986 34743
rect 24094 34777 24146 34786
rect 24094 34743 24103 34777
rect 24103 34743 24137 34777
rect 24137 34743 24146 34777
rect 24094 34734 24146 34743
rect 24254 34777 24306 34786
rect 24254 34743 24263 34777
rect 24263 34743 24297 34777
rect 24297 34743 24306 34777
rect 24254 34734 24306 34743
rect 24414 34777 24466 34786
rect 24414 34743 24423 34777
rect 24423 34743 24457 34777
rect 24457 34743 24466 34777
rect 24414 34734 24466 34743
rect 24574 34777 24626 34786
rect 24574 34743 24583 34777
rect 24583 34743 24617 34777
rect 24617 34743 24626 34777
rect 24574 34734 24626 34743
rect 24734 34777 24786 34786
rect 24734 34743 24743 34777
rect 24743 34743 24777 34777
rect 24777 34743 24786 34777
rect 24734 34734 24786 34743
rect 24894 34777 24946 34786
rect 24894 34743 24903 34777
rect 24903 34743 24937 34777
rect 24937 34743 24946 34777
rect 24894 34734 24946 34743
rect 25054 34777 25106 34786
rect 25054 34743 25063 34777
rect 25063 34743 25097 34777
rect 25097 34743 25106 34777
rect 25054 34734 25106 34743
rect 25214 34777 25266 34786
rect 25214 34743 25223 34777
rect 25223 34743 25257 34777
rect 25257 34743 25266 34777
rect 25214 34734 25266 34743
rect 25374 34777 25426 34786
rect 25374 34743 25383 34777
rect 25383 34743 25417 34777
rect 25417 34743 25426 34777
rect 25374 34734 25426 34743
rect 25534 34777 25586 34786
rect 25534 34743 25543 34777
rect 25543 34743 25577 34777
rect 25577 34743 25586 34777
rect 25534 34734 25586 34743
rect 25694 34777 25746 34786
rect 25694 34743 25703 34777
rect 25703 34743 25737 34777
rect 25737 34743 25746 34777
rect 25694 34734 25746 34743
rect 25854 34777 25906 34786
rect 25854 34743 25863 34777
rect 25863 34743 25897 34777
rect 25897 34743 25906 34777
rect 25854 34734 25906 34743
rect 26014 34777 26066 34786
rect 26014 34743 26023 34777
rect 26023 34743 26057 34777
rect 26057 34743 26066 34777
rect 26014 34734 26066 34743
rect 26174 34777 26226 34786
rect 26174 34743 26183 34777
rect 26183 34743 26217 34777
rect 26217 34743 26226 34777
rect 26174 34734 26226 34743
rect 26334 34777 26386 34786
rect 26334 34743 26343 34777
rect 26343 34743 26377 34777
rect 26377 34743 26386 34777
rect 26334 34734 26386 34743
rect 26494 34777 26546 34786
rect 26494 34743 26503 34777
rect 26503 34743 26537 34777
rect 26537 34743 26546 34777
rect 26494 34734 26546 34743
rect 26654 34777 26706 34786
rect 26654 34743 26663 34777
rect 26663 34743 26697 34777
rect 26697 34743 26706 34777
rect 26654 34734 26706 34743
rect 26814 34777 26866 34786
rect 26814 34743 26823 34777
rect 26823 34743 26857 34777
rect 26857 34743 26866 34777
rect 26814 34734 26866 34743
rect 26974 34777 27026 34786
rect 26974 34743 26983 34777
rect 26983 34743 27017 34777
rect 27017 34743 27026 34777
rect 26974 34734 27026 34743
rect 27134 34777 27186 34786
rect 27134 34743 27143 34777
rect 27143 34743 27177 34777
rect 27177 34743 27186 34777
rect 27134 34734 27186 34743
rect 27294 34777 27346 34786
rect 27294 34743 27303 34777
rect 27303 34743 27337 34777
rect 27337 34743 27346 34777
rect 27294 34734 27346 34743
rect 27454 34777 27506 34786
rect 27454 34743 27463 34777
rect 27463 34743 27497 34777
rect 27497 34743 27506 34777
rect 27454 34734 27506 34743
rect 27614 34777 27666 34786
rect 27614 34743 27623 34777
rect 27623 34743 27657 34777
rect 27657 34743 27666 34777
rect 27614 34734 27666 34743
rect 27774 34777 27826 34786
rect 27774 34743 27783 34777
rect 27783 34743 27817 34777
rect 27817 34743 27826 34777
rect 27774 34734 27826 34743
rect 27934 34777 27986 34786
rect 27934 34743 27943 34777
rect 27943 34743 27977 34777
rect 27977 34743 27986 34777
rect 27934 34734 27986 34743
rect 28094 34777 28146 34786
rect 28094 34743 28103 34777
rect 28103 34743 28137 34777
rect 28137 34743 28146 34777
rect 28094 34734 28146 34743
rect 28254 34777 28306 34786
rect 28254 34743 28263 34777
rect 28263 34743 28297 34777
rect 28297 34743 28306 34777
rect 28254 34734 28306 34743
rect 28414 34777 28466 34786
rect 28414 34743 28423 34777
rect 28423 34743 28457 34777
rect 28457 34743 28466 34777
rect 28414 34734 28466 34743
rect 28574 34777 28626 34786
rect 28574 34743 28583 34777
rect 28583 34743 28617 34777
rect 28617 34743 28626 34777
rect 28574 34734 28626 34743
rect 28734 34777 28786 34786
rect 28734 34743 28743 34777
rect 28743 34743 28777 34777
rect 28777 34743 28786 34777
rect 28734 34734 28786 34743
rect 28894 34777 28946 34786
rect 28894 34743 28903 34777
rect 28903 34743 28937 34777
rect 28937 34743 28946 34777
rect 28894 34734 28946 34743
rect 29054 34777 29106 34786
rect 29054 34743 29063 34777
rect 29063 34743 29097 34777
rect 29097 34743 29106 34777
rect 29054 34734 29106 34743
rect 29214 34777 29266 34786
rect 29214 34743 29223 34777
rect 29223 34743 29257 34777
rect 29257 34743 29266 34777
rect 29214 34734 29266 34743
rect 29374 34777 29426 34786
rect 29374 34743 29383 34777
rect 29383 34743 29417 34777
rect 29417 34743 29426 34777
rect 29374 34734 29426 34743
rect 33534 34777 33586 34786
rect 33534 34743 33543 34777
rect 33543 34743 33577 34777
rect 33577 34743 33586 34777
rect 33534 34734 33586 34743
rect 33694 34777 33746 34786
rect 33694 34743 33703 34777
rect 33703 34743 33737 34777
rect 33737 34743 33746 34777
rect 33694 34734 33746 34743
rect 33854 34777 33906 34786
rect 33854 34743 33863 34777
rect 33863 34743 33897 34777
rect 33897 34743 33906 34777
rect 33854 34734 33906 34743
rect 34014 34777 34066 34786
rect 34014 34743 34023 34777
rect 34023 34743 34057 34777
rect 34057 34743 34066 34777
rect 34014 34734 34066 34743
rect 34174 34777 34226 34786
rect 34174 34743 34183 34777
rect 34183 34743 34217 34777
rect 34217 34743 34226 34777
rect 34174 34734 34226 34743
rect 34334 34777 34386 34786
rect 34334 34743 34343 34777
rect 34343 34743 34377 34777
rect 34377 34743 34386 34777
rect 34334 34734 34386 34743
rect 34494 34777 34546 34786
rect 34494 34743 34503 34777
rect 34503 34743 34537 34777
rect 34537 34743 34546 34777
rect 34494 34734 34546 34743
rect 34654 34777 34706 34786
rect 34654 34743 34663 34777
rect 34663 34743 34697 34777
rect 34697 34743 34706 34777
rect 34654 34734 34706 34743
rect 34814 34777 34866 34786
rect 34814 34743 34823 34777
rect 34823 34743 34857 34777
rect 34857 34743 34866 34777
rect 34814 34734 34866 34743
rect 34974 34777 35026 34786
rect 34974 34743 34983 34777
rect 34983 34743 35017 34777
rect 35017 34743 35026 34777
rect 34974 34734 35026 34743
rect 35134 34777 35186 34786
rect 35134 34743 35143 34777
rect 35143 34743 35177 34777
rect 35177 34743 35186 34777
rect 35134 34734 35186 34743
rect 35294 34777 35346 34786
rect 35294 34743 35303 34777
rect 35303 34743 35337 34777
rect 35337 34743 35346 34777
rect 35294 34734 35346 34743
rect 35454 34777 35506 34786
rect 35454 34743 35463 34777
rect 35463 34743 35497 34777
rect 35497 34743 35506 34777
rect 35454 34734 35506 34743
rect 35614 34777 35666 34786
rect 35614 34743 35623 34777
rect 35623 34743 35657 34777
rect 35657 34743 35666 34777
rect 35614 34734 35666 34743
rect 35774 34777 35826 34786
rect 35774 34743 35783 34777
rect 35783 34743 35817 34777
rect 35817 34743 35826 34777
rect 35774 34734 35826 34743
rect 35934 34777 35986 34786
rect 35934 34743 35943 34777
rect 35943 34743 35977 34777
rect 35977 34743 35986 34777
rect 35934 34734 35986 34743
rect 36094 34777 36146 34786
rect 36094 34743 36103 34777
rect 36103 34743 36137 34777
rect 36137 34743 36146 34777
rect 36094 34734 36146 34743
rect 36254 34777 36306 34786
rect 36254 34743 36263 34777
rect 36263 34743 36297 34777
rect 36297 34743 36306 34777
rect 36254 34734 36306 34743
rect 36414 34777 36466 34786
rect 36414 34743 36423 34777
rect 36423 34743 36457 34777
rect 36457 34743 36466 34777
rect 36414 34734 36466 34743
rect 36574 34777 36626 34786
rect 36574 34743 36583 34777
rect 36583 34743 36617 34777
rect 36617 34743 36626 34777
rect 36574 34734 36626 34743
rect 36734 34777 36786 34786
rect 36734 34743 36743 34777
rect 36743 34743 36777 34777
rect 36777 34743 36786 34777
rect 36734 34734 36786 34743
rect 36894 34777 36946 34786
rect 36894 34743 36903 34777
rect 36903 34743 36937 34777
rect 36937 34743 36946 34777
rect 36894 34734 36946 34743
rect 37054 34777 37106 34786
rect 37054 34743 37063 34777
rect 37063 34743 37097 34777
rect 37097 34743 37106 34777
rect 37054 34734 37106 34743
rect 37214 34777 37266 34786
rect 37214 34743 37223 34777
rect 37223 34743 37257 34777
rect 37257 34743 37266 34777
rect 37214 34734 37266 34743
rect 37374 34777 37426 34786
rect 37374 34743 37383 34777
rect 37383 34743 37417 34777
rect 37417 34743 37426 34777
rect 37374 34734 37426 34743
rect 37534 34777 37586 34786
rect 37534 34743 37543 34777
rect 37543 34743 37577 34777
rect 37577 34743 37586 34777
rect 37534 34734 37586 34743
rect 37694 34777 37746 34786
rect 37694 34743 37703 34777
rect 37703 34743 37737 34777
rect 37737 34743 37746 34777
rect 37694 34734 37746 34743
rect 37854 34777 37906 34786
rect 37854 34743 37863 34777
rect 37863 34743 37897 34777
rect 37897 34743 37906 34777
rect 37854 34734 37906 34743
rect 38014 34777 38066 34786
rect 38014 34743 38023 34777
rect 38023 34743 38057 34777
rect 38057 34743 38066 34777
rect 38014 34734 38066 34743
rect 38174 34777 38226 34786
rect 38174 34743 38183 34777
rect 38183 34743 38217 34777
rect 38217 34743 38226 34777
rect 38174 34734 38226 34743
rect 38334 34777 38386 34786
rect 38334 34743 38343 34777
rect 38343 34743 38377 34777
rect 38377 34743 38386 34777
rect 38334 34734 38386 34743
rect 38494 34777 38546 34786
rect 38494 34743 38503 34777
rect 38503 34743 38537 34777
rect 38537 34743 38546 34777
rect 38494 34734 38546 34743
rect 38654 34777 38706 34786
rect 38654 34743 38663 34777
rect 38663 34743 38697 34777
rect 38697 34743 38706 34777
rect 38654 34734 38706 34743
rect 38814 34777 38866 34786
rect 38814 34743 38823 34777
rect 38823 34743 38857 34777
rect 38857 34743 38866 34777
rect 38814 34734 38866 34743
rect 38974 34777 39026 34786
rect 38974 34743 38983 34777
rect 38983 34743 39017 34777
rect 39017 34743 39026 34777
rect 38974 34734 39026 34743
rect 39134 34777 39186 34786
rect 39134 34743 39143 34777
rect 39143 34743 39177 34777
rect 39177 34743 39186 34777
rect 39134 34734 39186 34743
rect 39294 34777 39346 34786
rect 39294 34743 39303 34777
rect 39303 34743 39337 34777
rect 39337 34743 39346 34777
rect 39294 34734 39346 34743
rect 39454 34777 39506 34786
rect 39454 34743 39463 34777
rect 39463 34743 39497 34777
rect 39497 34743 39506 34777
rect 39454 34734 39506 34743
rect 39614 34777 39666 34786
rect 39614 34743 39623 34777
rect 39623 34743 39657 34777
rect 39657 34743 39666 34777
rect 39614 34734 39666 34743
rect 39774 34777 39826 34786
rect 39774 34743 39783 34777
rect 39783 34743 39817 34777
rect 39817 34743 39826 34777
rect 39774 34734 39826 34743
rect 39934 34777 39986 34786
rect 39934 34743 39943 34777
rect 39943 34743 39977 34777
rect 39977 34743 39986 34777
rect 39934 34734 39986 34743
rect 40094 34777 40146 34786
rect 40094 34743 40103 34777
rect 40103 34743 40137 34777
rect 40137 34743 40146 34777
rect 40094 34734 40146 34743
rect 40254 34777 40306 34786
rect 40254 34743 40263 34777
rect 40263 34743 40297 34777
rect 40297 34743 40306 34777
rect 40254 34734 40306 34743
rect 40414 34777 40466 34786
rect 40414 34743 40423 34777
rect 40423 34743 40457 34777
rect 40457 34743 40466 34777
rect 40414 34734 40466 34743
rect 40574 34777 40626 34786
rect 40574 34743 40583 34777
rect 40583 34743 40617 34777
rect 40617 34743 40626 34777
rect 40574 34734 40626 34743
rect 40734 34777 40786 34786
rect 40734 34743 40743 34777
rect 40743 34743 40777 34777
rect 40777 34743 40786 34777
rect 40734 34734 40786 34743
rect 40894 34777 40946 34786
rect 40894 34743 40903 34777
rect 40903 34743 40937 34777
rect 40937 34743 40946 34777
rect 40894 34734 40946 34743
rect 41054 34777 41106 34786
rect 41054 34743 41063 34777
rect 41063 34743 41097 34777
rect 41097 34743 41106 34777
rect 41054 34734 41106 34743
rect 41214 34777 41266 34786
rect 41214 34743 41223 34777
rect 41223 34743 41257 34777
rect 41257 34743 41266 34777
rect 41214 34734 41266 34743
rect 41374 34777 41426 34786
rect 41374 34743 41383 34777
rect 41383 34743 41417 34777
rect 41417 34743 41426 34777
rect 41374 34734 41426 34743
rect 41534 34777 41586 34786
rect 41534 34743 41543 34777
rect 41543 34743 41577 34777
rect 41577 34743 41586 34777
rect 41534 34734 41586 34743
rect 41694 34777 41746 34786
rect 41694 34743 41703 34777
rect 41703 34743 41737 34777
rect 41737 34743 41746 34777
rect 41694 34734 41746 34743
rect 41854 34777 41906 34786
rect 41854 34743 41863 34777
rect 41863 34743 41897 34777
rect 41897 34743 41906 34777
rect 41854 34734 41906 34743
rect 14 34457 66 34466
rect 14 34423 23 34457
rect 23 34423 57 34457
rect 57 34423 66 34457
rect 14 34414 66 34423
rect 174 34457 226 34466
rect 174 34423 183 34457
rect 183 34423 217 34457
rect 217 34423 226 34457
rect 174 34414 226 34423
rect 334 34457 386 34466
rect 334 34423 343 34457
rect 343 34423 377 34457
rect 377 34423 386 34457
rect 334 34414 386 34423
rect 494 34457 546 34466
rect 494 34423 503 34457
rect 503 34423 537 34457
rect 537 34423 546 34457
rect 494 34414 546 34423
rect 654 34457 706 34466
rect 654 34423 663 34457
rect 663 34423 697 34457
rect 697 34423 706 34457
rect 654 34414 706 34423
rect 814 34457 866 34466
rect 814 34423 823 34457
rect 823 34423 857 34457
rect 857 34423 866 34457
rect 814 34414 866 34423
rect 974 34457 1026 34466
rect 974 34423 983 34457
rect 983 34423 1017 34457
rect 1017 34423 1026 34457
rect 974 34414 1026 34423
rect 1134 34457 1186 34466
rect 1134 34423 1143 34457
rect 1143 34423 1177 34457
rect 1177 34423 1186 34457
rect 1134 34414 1186 34423
rect 1294 34457 1346 34466
rect 1294 34423 1303 34457
rect 1303 34423 1337 34457
rect 1337 34423 1346 34457
rect 1294 34414 1346 34423
rect 1454 34457 1506 34466
rect 1454 34423 1463 34457
rect 1463 34423 1497 34457
rect 1497 34423 1506 34457
rect 1454 34414 1506 34423
rect 1614 34457 1666 34466
rect 1614 34423 1623 34457
rect 1623 34423 1657 34457
rect 1657 34423 1666 34457
rect 1614 34414 1666 34423
rect 1774 34457 1826 34466
rect 1774 34423 1783 34457
rect 1783 34423 1817 34457
rect 1817 34423 1826 34457
rect 1774 34414 1826 34423
rect 1934 34457 1986 34466
rect 1934 34423 1943 34457
rect 1943 34423 1977 34457
rect 1977 34423 1986 34457
rect 1934 34414 1986 34423
rect 2094 34457 2146 34466
rect 2094 34423 2103 34457
rect 2103 34423 2137 34457
rect 2137 34423 2146 34457
rect 2094 34414 2146 34423
rect 2254 34457 2306 34466
rect 2254 34423 2263 34457
rect 2263 34423 2297 34457
rect 2297 34423 2306 34457
rect 2254 34414 2306 34423
rect 2414 34457 2466 34466
rect 2414 34423 2423 34457
rect 2423 34423 2457 34457
rect 2457 34423 2466 34457
rect 2414 34414 2466 34423
rect 2574 34457 2626 34466
rect 2574 34423 2583 34457
rect 2583 34423 2617 34457
rect 2617 34423 2626 34457
rect 2574 34414 2626 34423
rect 2734 34457 2786 34466
rect 2734 34423 2743 34457
rect 2743 34423 2777 34457
rect 2777 34423 2786 34457
rect 2734 34414 2786 34423
rect 2894 34457 2946 34466
rect 2894 34423 2903 34457
rect 2903 34423 2937 34457
rect 2937 34423 2946 34457
rect 2894 34414 2946 34423
rect 3054 34457 3106 34466
rect 3054 34423 3063 34457
rect 3063 34423 3097 34457
rect 3097 34423 3106 34457
rect 3054 34414 3106 34423
rect 3214 34457 3266 34466
rect 3214 34423 3223 34457
rect 3223 34423 3257 34457
rect 3257 34423 3266 34457
rect 3214 34414 3266 34423
rect 3374 34457 3426 34466
rect 3374 34423 3383 34457
rect 3383 34423 3417 34457
rect 3417 34423 3426 34457
rect 3374 34414 3426 34423
rect 3534 34457 3586 34466
rect 3534 34423 3543 34457
rect 3543 34423 3577 34457
rect 3577 34423 3586 34457
rect 3534 34414 3586 34423
rect 3694 34457 3746 34466
rect 3694 34423 3703 34457
rect 3703 34423 3737 34457
rect 3737 34423 3746 34457
rect 3694 34414 3746 34423
rect 3854 34457 3906 34466
rect 3854 34423 3863 34457
rect 3863 34423 3897 34457
rect 3897 34423 3906 34457
rect 3854 34414 3906 34423
rect 4014 34457 4066 34466
rect 4014 34423 4023 34457
rect 4023 34423 4057 34457
rect 4057 34423 4066 34457
rect 4014 34414 4066 34423
rect 4174 34457 4226 34466
rect 4174 34423 4183 34457
rect 4183 34423 4217 34457
rect 4217 34423 4226 34457
rect 4174 34414 4226 34423
rect 4334 34457 4386 34466
rect 4334 34423 4343 34457
rect 4343 34423 4377 34457
rect 4377 34423 4386 34457
rect 4334 34414 4386 34423
rect 4494 34457 4546 34466
rect 4494 34423 4503 34457
rect 4503 34423 4537 34457
rect 4537 34423 4546 34457
rect 4494 34414 4546 34423
rect 4654 34457 4706 34466
rect 4654 34423 4663 34457
rect 4663 34423 4697 34457
rect 4697 34423 4706 34457
rect 4654 34414 4706 34423
rect 4814 34457 4866 34466
rect 4814 34423 4823 34457
rect 4823 34423 4857 34457
rect 4857 34423 4866 34457
rect 4814 34414 4866 34423
rect 4974 34457 5026 34466
rect 4974 34423 4983 34457
rect 4983 34423 5017 34457
rect 5017 34423 5026 34457
rect 4974 34414 5026 34423
rect 5134 34457 5186 34466
rect 5134 34423 5143 34457
rect 5143 34423 5177 34457
rect 5177 34423 5186 34457
rect 5134 34414 5186 34423
rect 5294 34457 5346 34466
rect 5294 34423 5303 34457
rect 5303 34423 5337 34457
rect 5337 34423 5346 34457
rect 5294 34414 5346 34423
rect 5454 34457 5506 34466
rect 5454 34423 5463 34457
rect 5463 34423 5497 34457
rect 5497 34423 5506 34457
rect 5454 34414 5506 34423
rect 5614 34457 5666 34466
rect 5614 34423 5623 34457
rect 5623 34423 5657 34457
rect 5657 34423 5666 34457
rect 5614 34414 5666 34423
rect 5774 34457 5826 34466
rect 5774 34423 5783 34457
rect 5783 34423 5817 34457
rect 5817 34423 5826 34457
rect 5774 34414 5826 34423
rect 5934 34457 5986 34466
rect 5934 34423 5943 34457
rect 5943 34423 5977 34457
rect 5977 34423 5986 34457
rect 5934 34414 5986 34423
rect 6094 34457 6146 34466
rect 6094 34423 6103 34457
rect 6103 34423 6137 34457
rect 6137 34423 6146 34457
rect 6094 34414 6146 34423
rect 6254 34457 6306 34466
rect 6254 34423 6263 34457
rect 6263 34423 6297 34457
rect 6297 34423 6306 34457
rect 6254 34414 6306 34423
rect 6414 34457 6466 34466
rect 6414 34423 6423 34457
rect 6423 34423 6457 34457
rect 6457 34423 6466 34457
rect 6414 34414 6466 34423
rect 6574 34457 6626 34466
rect 6574 34423 6583 34457
rect 6583 34423 6617 34457
rect 6617 34423 6626 34457
rect 6574 34414 6626 34423
rect 6734 34457 6786 34466
rect 6734 34423 6743 34457
rect 6743 34423 6777 34457
rect 6777 34423 6786 34457
rect 6734 34414 6786 34423
rect 6894 34457 6946 34466
rect 6894 34423 6903 34457
rect 6903 34423 6937 34457
rect 6937 34423 6946 34457
rect 6894 34414 6946 34423
rect 7054 34457 7106 34466
rect 7054 34423 7063 34457
rect 7063 34423 7097 34457
rect 7097 34423 7106 34457
rect 7054 34414 7106 34423
rect 7214 34457 7266 34466
rect 7214 34423 7223 34457
rect 7223 34423 7257 34457
rect 7257 34423 7266 34457
rect 7214 34414 7266 34423
rect 7374 34457 7426 34466
rect 7374 34423 7383 34457
rect 7383 34423 7417 34457
rect 7417 34423 7426 34457
rect 7374 34414 7426 34423
rect 7534 34457 7586 34466
rect 7534 34423 7543 34457
rect 7543 34423 7577 34457
rect 7577 34423 7586 34457
rect 7534 34414 7586 34423
rect 7694 34457 7746 34466
rect 7694 34423 7703 34457
rect 7703 34423 7737 34457
rect 7737 34423 7746 34457
rect 7694 34414 7746 34423
rect 7854 34457 7906 34466
rect 7854 34423 7863 34457
rect 7863 34423 7897 34457
rect 7897 34423 7906 34457
rect 7854 34414 7906 34423
rect 8014 34457 8066 34466
rect 8014 34423 8023 34457
rect 8023 34423 8057 34457
rect 8057 34423 8066 34457
rect 8014 34414 8066 34423
rect 8174 34457 8226 34466
rect 8174 34423 8183 34457
rect 8183 34423 8217 34457
rect 8217 34423 8226 34457
rect 8174 34414 8226 34423
rect 8334 34457 8386 34466
rect 8334 34423 8343 34457
rect 8343 34423 8377 34457
rect 8377 34423 8386 34457
rect 8334 34414 8386 34423
rect 12494 34457 12546 34466
rect 12494 34423 12503 34457
rect 12503 34423 12537 34457
rect 12537 34423 12546 34457
rect 12494 34414 12546 34423
rect 12654 34457 12706 34466
rect 12654 34423 12663 34457
rect 12663 34423 12697 34457
rect 12697 34423 12706 34457
rect 12654 34414 12706 34423
rect 12814 34457 12866 34466
rect 12814 34423 12823 34457
rect 12823 34423 12857 34457
rect 12857 34423 12866 34457
rect 12814 34414 12866 34423
rect 12974 34457 13026 34466
rect 12974 34423 12983 34457
rect 12983 34423 13017 34457
rect 13017 34423 13026 34457
rect 12974 34414 13026 34423
rect 13134 34457 13186 34466
rect 13134 34423 13143 34457
rect 13143 34423 13177 34457
rect 13177 34423 13186 34457
rect 13134 34414 13186 34423
rect 13294 34457 13346 34466
rect 13294 34423 13303 34457
rect 13303 34423 13337 34457
rect 13337 34423 13346 34457
rect 13294 34414 13346 34423
rect 13454 34457 13506 34466
rect 13454 34423 13463 34457
rect 13463 34423 13497 34457
rect 13497 34423 13506 34457
rect 13454 34414 13506 34423
rect 13614 34457 13666 34466
rect 13614 34423 13623 34457
rect 13623 34423 13657 34457
rect 13657 34423 13666 34457
rect 13614 34414 13666 34423
rect 13774 34457 13826 34466
rect 13774 34423 13783 34457
rect 13783 34423 13817 34457
rect 13817 34423 13826 34457
rect 13774 34414 13826 34423
rect 13934 34457 13986 34466
rect 13934 34423 13943 34457
rect 13943 34423 13977 34457
rect 13977 34423 13986 34457
rect 13934 34414 13986 34423
rect 14094 34457 14146 34466
rect 14094 34423 14103 34457
rect 14103 34423 14137 34457
rect 14137 34423 14146 34457
rect 14094 34414 14146 34423
rect 14254 34457 14306 34466
rect 14254 34423 14263 34457
rect 14263 34423 14297 34457
rect 14297 34423 14306 34457
rect 14254 34414 14306 34423
rect 14414 34457 14466 34466
rect 14414 34423 14423 34457
rect 14423 34423 14457 34457
rect 14457 34423 14466 34457
rect 14414 34414 14466 34423
rect 14574 34457 14626 34466
rect 14574 34423 14583 34457
rect 14583 34423 14617 34457
rect 14617 34423 14626 34457
rect 14574 34414 14626 34423
rect 14734 34457 14786 34466
rect 14734 34423 14743 34457
rect 14743 34423 14777 34457
rect 14777 34423 14786 34457
rect 14734 34414 14786 34423
rect 14894 34457 14946 34466
rect 14894 34423 14903 34457
rect 14903 34423 14937 34457
rect 14937 34423 14946 34457
rect 14894 34414 14946 34423
rect 15054 34457 15106 34466
rect 15054 34423 15063 34457
rect 15063 34423 15097 34457
rect 15097 34423 15106 34457
rect 15054 34414 15106 34423
rect 15214 34457 15266 34466
rect 15214 34423 15223 34457
rect 15223 34423 15257 34457
rect 15257 34423 15266 34457
rect 15214 34414 15266 34423
rect 15374 34457 15426 34466
rect 15374 34423 15383 34457
rect 15383 34423 15417 34457
rect 15417 34423 15426 34457
rect 15374 34414 15426 34423
rect 15534 34457 15586 34466
rect 15534 34423 15543 34457
rect 15543 34423 15577 34457
rect 15577 34423 15586 34457
rect 15534 34414 15586 34423
rect 15694 34457 15746 34466
rect 15694 34423 15703 34457
rect 15703 34423 15737 34457
rect 15737 34423 15746 34457
rect 15694 34414 15746 34423
rect 15854 34457 15906 34466
rect 15854 34423 15863 34457
rect 15863 34423 15897 34457
rect 15897 34423 15906 34457
rect 15854 34414 15906 34423
rect 16014 34457 16066 34466
rect 16014 34423 16023 34457
rect 16023 34423 16057 34457
rect 16057 34423 16066 34457
rect 16014 34414 16066 34423
rect 16174 34457 16226 34466
rect 16174 34423 16183 34457
rect 16183 34423 16217 34457
rect 16217 34423 16226 34457
rect 16174 34414 16226 34423
rect 16334 34457 16386 34466
rect 16334 34423 16343 34457
rect 16343 34423 16377 34457
rect 16377 34423 16386 34457
rect 16334 34414 16386 34423
rect 16494 34457 16546 34466
rect 16494 34423 16503 34457
rect 16503 34423 16537 34457
rect 16537 34423 16546 34457
rect 16494 34414 16546 34423
rect 16654 34457 16706 34466
rect 16654 34423 16663 34457
rect 16663 34423 16697 34457
rect 16697 34423 16706 34457
rect 16654 34414 16706 34423
rect 16814 34457 16866 34466
rect 16814 34423 16823 34457
rect 16823 34423 16857 34457
rect 16857 34423 16866 34457
rect 16814 34414 16866 34423
rect 16974 34457 17026 34466
rect 16974 34423 16983 34457
rect 16983 34423 17017 34457
rect 17017 34423 17026 34457
rect 16974 34414 17026 34423
rect 17134 34457 17186 34466
rect 17134 34423 17143 34457
rect 17143 34423 17177 34457
rect 17177 34423 17186 34457
rect 17134 34414 17186 34423
rect 17294 34457 17346 34466
rect 17294 34423 17303 34457
rect 17303 34423 17337 34457
rect 17337 34423 17346 34457
rect 17294 34414 17346 34423
rect 17454 34457 17506 34466
rect 17454 34423 17463 34457
rect 17463 34423 17497 34457
rect 17497 34423 17506 34457
rect 17454 34414 17506 34423
rect 17614 34457 17666 34466
rect 17614 34423 17623 34457
rect 17623 34423 17657 34457
rect 17657 34423 17666 34457
rect 17614 34414 17666 34423
rect 17774 34457 17826 34466
rect 17774 34423 17783 34457
rect 17783 34423 17817 34457
rect 17817 34423 17826 34457
rect 17774 34414 17826 34423
rect 17934 34457 17986 34466
rect 17934 34423 17943 34457
rect 17943 34423 17977 34457
rect 17977 34423 17986 34457
rect 17934 34414 17986 34423
rect 18094 34457 18146 34466
rect 18094 34423 18103 34457
rect 18103 34423 18137 34457
rect 18137 34423 18146 34457
rect 18094 34414 18146 34423
rect 18254 34457 18306 34466
rect 18254 34423 18263 34457
rect 18263 34423 18297 34457
rect 18297 34423 18306 34457
rect 18254 34414 18306 34423
rect 18414 34457 18466 34466
rect 18414 34423 18423 34457
rect 18423 34423 18457 34457
rect 18457 34423 18466 34457
rect 18414 34414 18466 34423
rect 18574 34457 18626 34466
rect 18574 34423 18583 34457
rect 18583 34423 18617 34457
rect 18617 34423 18626 34457
rect 18574 34414 18626 34423
rect 18734 34457 18786 34466
rect 18734 34423 18743 34457
rect 18743 34423 18777 34457
rect 18777 34423 18786 34457
rect 18734 34414 18786 34423
rect 18894 34457 18946 34466
rect 18894 34423 18903 34457
rect 18903 34423 18937 34457
rect 18937 34423 18946 34457
rect 18894 34414 18946 34423
rect 23134 34457 23186 34466
rect 23134 34423 23143 34457
rect 23143 34423 23177 34457
rect 23177 34423 23186 34457
rect 23134 34414 23186 34423
rect 23294 34457 23346 34466
rect 23294 34423 23303 34457
rect 23303 34423 23337 34457
rect 23337 34423 23346 34457
rect 23294 34414 23346 34423
rect 23454 34457 23506 34466
rect 23454 34423 23463 34457
rect 23463 34423 23497 34457
rect 23497 34423 23506 34457
rect 23454 34414 23506 34423
rect 23614 34457 23666 34466
rect 23614 34423 23623 34457
rect 23623 34423 23657 34457
rect 23657 34423 23666 34457
rect 23614 34414 23666 34423
rect 23774 34457 23826 34466
rect 23774 34423 23783 34457
rect 23783 34423 23817 34457
rect 23817 34423 23826 34457
rect 23774 34414 23826 34423
rect 23934 34457 23986 34466
rect 23934 34423 23943 34457
rect 23943 34423 23977 34457
rect 23977 34423 23986 34457
rect 23934 34414 23986 34423
rect 24094 34457 24146 34466
rect 24094 34423 24103 34457
rect 24103 34423 24137 34457
rect 24137 34423 24146 34457
rect 24094 34414 24146 34423
rect 24254 34457 24306 34466
rect 24254 34423 24263 34457
rect 24263 34423 24297 34457
rect 24297 34423 24306 34457
rect 24254 34414 24306 34423
rect 24414 34457 24466 34466
rect 24414 34423 24423 34457
rect 24423 34423 24457 34457
rect 24457 34423 24466 34457
rect 24414 34414 24466 34423
rect 24574 34457 24626 34466
rect 24574 34423 24583 34457
rect 24583 34423 24617 34457
rect 24617 34423 24626 34457
rect 24574 34414 24626 34423
rect 24734 34457 24786 34466
rect 24734 34423 24743 34457
rect 24743 34423 24777 34457
rect 24777 34423 24786 34457
rect 24734 34414 24786 34423
rect 24894 34457 24946 34466
rect 24894 34423 24903 34457
rect 24903 34423 24937 34457
rect 24937 34423 24946 34457
rect 24894 34414 24946 34423
rect 25054 34457 25106 34466
rect 25054 34423 25063 34457
rect 25063 34423 25097 34457
rect 25097 34423 25106 34457
rect 25054 34414 25106 34423
rect 25214 34457 25266 34466
rect 25214 34423 25223 34457
rect 25223 34423 25257 34457
rect 25257 34423 25266 34457
rect 25214 34414 25266 34423
rect 25374 34457 25426 34466
rect 25374 34423 25383 34457
rect 25383 34423 25417 34457
rect 25417 34423 25426 34457
rect 25374 34414 25426 34423
rect 25534 34457 25586 34466
rect 25534 34423 25543 34457
rect 25543 34423 25577 34457
rect 25577 34423 25586 34457
rect 25534 34414 25586 34423
rect 25694 34457 25746 34466
rect 25694 34423 25703 34457
rect 25703 34423 25737 34457
rect 25737 34423 25746 34457
rect 25694 34414 25746 34423
rect 25854 34457 25906 34466
rect 25854 34423 25863 34457
rect 25863 34423 25897 34457
rect 25897 34423 25906 34457
rect 25854 34414 25906 34423
rect 26014 34457 26066 34466
rect 26014 34423 26023 34457
rect 26023 34423 26057 34457
rect 26057 34423 26066 34457
rect 26014 34414 26066 34423
rect 26174 34457 26226 34466
rect 26174 34423 26183 34457
rect 26183 34423 26217 34457
rect 26217 34423 26226 34457
rect 26174 34414 26226 34423
rect 26334 34457 26386 34466
rect 26334 34423 26343 34457
rect 26343 34423 26377 34457
rect 26377 34423 26386 34457
rect 26334 34414 26386 34423
rect 26494 34457 26546 34466
rect 26494 34423 26503 34457
rect 26503 34423 26537 34457
rect 26537 34423 26546 34457
rect 26494 34414 26546 34423
rect 26654 34457 26706 34466
rect 26654 34423 26663 34457
rect 26663 34423 26697 34457
rect 26697 34423 26706 34457
rect 26654 34414 26706 34423
rect 26814 34457 26866 34466
rect 26814 34423 26823 34457
rect 26823 34423 26857 34457
rect 26857 34423 26866 34457
rect 26814 34414 26866 34423
rect 26974 34457 27026 34466
rect 26974 34423 26983 34457
rect 26983 34423 27017 34457
rect 27017 34423 27026 34457
rect 26974 34414 27026 34423
rect 27134 34457 27186 34466
rect 27134 34423 27143 34457
rect 27143 34423 27177 34457
rect 27177 34423 27186 34457
rect 27134 34414 27186 34423
rect 27294 34457 27346 34466
rect 27294 34423 27303 34457
rect 27303 34423 27337 34457
rect 27337 34423 27346 34457
rect 27294 34414 27346 34423
rect 27454 34457 27506 34466
rect 27454 34423 27463 34457
rect 27463 34423 27497 34457
rect 27497 34423 27506 34457
rect 27454 34414 27506 34423
rect 27614 34457 27666 34466
rect 27614 34423 27623 34457
rect 27623 34423 27657 34457
rect 27657 34423 27666 34457
rect 27614 34414 27666 34423
rect 27774 34457 27826 34466
rect 27774 34423 27783 34457
rect 27783 34423 27817 34457
rect 27817 34423 27826 34457
rect 27774 34414 27826 34423
rect 27934 34457 27986 34466
rect 27934 34423 27943 34457
rect 27943 34423 27977 34457
rect 27977 34423 27986 34457
rect 27934 34414 27986 34423
rect 28094 34457 28146 34466
rect 28094 34423 28103 34457
rect 28103 34423 28137 34457
rect 28137 34423 28146 34457
rect 28094 34414 28146 34423
rect 28254 34457 28306 34466
rect 28254 34423 28263 34457
rect 28263 34423 28297 34457
rect 28297 34423 28306 34457
rect 28254 34414 28306 34423
rect 28414 34457 28466 34466
rect 28414 34423 28423 34457
rect 28423 34423 28457 34457
rect 28457 34423 28466 34457
rect 28414 34414 28466 34423
rect 28574 34457 28626 34466
rect 28574 34423 28583 34457
rect 28583 34423 28617 34457
rect 28617 34423 28626 34457
rect 28574 34414 28626 34423
rect 28734 34457 28786 34466
rect 28734 34423 28743 34457
rect 28743 34423 28777 34457
rect 28777 34423 28786 34457
rect 28734 34414 28786 34423
rect 28894 34457 28946 34466
rect 28894 34423 28903 34457
rect 28903 34423 28937 34457
rect 28937 34423 28946 34457
rect 28894 34414 28946 34423
rect 29054 34457 29106 34466
rect 29054 34423 29063 34457
rect 29063 34423 29097 34457
rect 29097 34423 29106 34457
rect 29054 34414 29106 34423
rect 29214 34457 29266 34466
rect 29214 34423 29223 34457
rect 29223 34423 29257 34457
rect 29257 34423 29266 34457
rect 29214 34414 29266 34423
rect 29374 34457 29426 34466
rect 29374 34423 29383 34457
rect 29383 34423 29417 34457
rect 29417 34423 29426 34457
rect 29374 34414 29426 34423
rect 33534 34457 33586 34466
rect 33534 34423 33543 34457
rect 33543 34423 33577 34457
rect 33577 34423 33586 34457
rect 33534 34414 33586 34423
rect 33694 34457 33746 34466
rect 33694 34423 33703 34457
rect 33703 34423 33737 34457
rect 33737 34423 33746 34457
rect 33694 34414 33746 34423
rect 33854 34457 33906 34466
rect 33854 34423 33863 34457
rect 33863 34423 33897 34457
rect 33897 34423 33906 34457
rect 33854 34414 33906 34423
rect 34014 34457 34066 34466
rect 34014 34423 34023 34457
rect 34023 34423 34057 34457
rect 34057 34423 34066 34457
rect 34014 34414 34066 34423
rect 34174 34457 34226 34466
rect 34174 34423 34183 34457
rect 34183 34423 34217 34457
rect 34217 34423 34226 34457
rect 34174 34414 34226 34423
rect 34334 34457 34386 34466
rect 34334 34423 34343 34457
rect 34343 34423 34377 34457
rect 34377 34423 34386 34457
rect 34334 34414 34386 34423
rect 34494 34457 34546 34466
rect 34494 34423 34503 34457
rect 34503 34423 34537 34457
rect 34537 34423 34546 34457
rect 34494 34414 34546 34423
rect 34654 34457 34706 34466
rect 34654 34423 34663 34457
rect 34663 34423 34697 34457
rect 34697 34423 34706 34457
rect 34654 34414 34706 34423
rect 34814 34457 34866 34466
rect 34814 34423 34823 34457
rect 34823 34423 34857 34457
rect 34857 34423 34866 34457
rect 34814 34414 34866 34423
rect 34974 34457 35026 34466
rect 34974 34423 34983 34457
rect 34983 34423 35017 34457
rect 35017 34423 35026 34457
rect 34974 34414 35026 34423
rect 35134 34457 35186 34466
rect 35134 34423 35143 34457
rect 35143 34423 35177 34457
rect 35177 34423 35186 34457
rect 35134 34414 35186 34423
rect 35294 34457 35346 34466
rect 35294 34423 35303 34457
rect 35303 34423 35337 34457
rect 35337 34423 35346 34457
rect 35294 34414 35346 34423
rect 35454 34457 35506 34466
rect 35454 34423 35463 34457
rect 35463 34423 35497 34457
rect 35497 34423 35506 34457
rect 35454 34414 35506 34423
rect 35614 34457 35666 34466
rect 35614 34423 35623 34457
rect 35623 34423 35657 34457
rect 35657 34423 35666 34457
rect 35614 34414 35666 34423
rect 35774 34457 35826 34466
rect 35774 34423 35783 34457
rect 35783 34423 35817 34457
rect 35817 34423 35826 34457
rect 35774 34414 35826 34423
rect 35934 34457 35986 34466
rect 35934 34423 35943 34457
rect 35943 34423 35977 34457
rect 35977 34423 35986 34457
rect 35934 34414 35986 34423
rect 36094 34457 36146 34466
rect 36094 34423 36103 34457
rect 36103 34423 36137 34457
rect 36137 34423 36146 34457
rect 36094 34414 36146 34423
rect 36254 34457 36306 34466
rect 36254 34423 36263 34457
rect 36263 34423 36297 34457
rect 36297 34423 36306 34457
rect 36254 34414 36306 34423
rect 36414 34457 36466 34466
rect 36414 34423 36423 34457
rect 36423 34423 36457 34457
rect 36457 34423 36466 34457
rect 36414 34414 36466 34423
rect 36574 34457 36626 34466
rect 36574 34423 36583 34457
rect 36583 34423 36617 34457
rect 36617 34423 36626 34457
rect 36574 34414 36626 34423
rect 36734 34457 36786 34466
rect 36734 34423 36743 34457
rect 36743 34423 36777 34457
rect 36777 34423 36786 34457
rect 36734 34414 36786 34423
rect 36894 34457 36946 34466
rect 36894 34423 36903 34457
rect 36903 34423 36937 34457
rect 36937 34423 36946 34457
rect 36894 34414 36946 34423
rect 37054 34457 37106 34466
rect 37054 34423 37063 34457
rect 37063 34423 37097 34457
rect 37097 34423 37106 34457
rect 37054 34414 37106 34423
rect 37214 34457 37266 34466
rect 37214 34423 37223 34457
rect 37223 34423 37257 34457
rect 37257 34423 37266 34457
rect 37214 34414 37266 34423
rect 37374 34457 37426 34466
rect 37374 34423 37383 34457
rect 37383 34423 37417 34457
rect 37417 34423 37426 34457
rect 37374 34414 37426 34423
rect 37534 34457 37586 34466
rect 37534 34423 37543 34457
rect 37543 34423 37577 34457
rect 37577 34423 37586 34457
rect 37534 34414 37586 34423
rect 37694 34457 37746 34466
rect 37694 34423 37703 34457
rect 37703 34423 37737 34457
rect 37737 34423 37746 34457
rect 37694 34414 37746 34423
rect 37854 34457 37906 34466
rect 37854 34423 37863 34457
rect 37863 34423 37897 34457
rect 37897 34423 37906 34457
rect 37854 34414 37906 34423
rect 38014 34457 38066 34466
rect 38014 34423 38023 34457
rect 38023 34423 38057 34457
rect 38057 34423 38066 34457
rect 38014 34414 38066 34423
rect 38174 34457 38226 34466
rect 38174 34423 38183 34457
rect 38183 34423 38217 34457
rect 38217 34423 38226 34457
rect 38174 34414 38226 34423
rect 38334 34457 38386 34466
rect 38334 34423 38343 34457
rect 38343 34423 38377 34457
rect 38377 34423 38386 34457
rect 38334 34414 38386 34423
rect 38494 34457 38546 34466
rect 38494 34423 38503 34457
rect 38503 34423 38537 34457
rect 38537 34423 38546 34457
rect 38494 34414 38546 34423
rect 38654 34457 38706 34466
rect 38654 34423 38663 34457
rect 38663 34423 38697 34457
rect 38697 34423 38706 34457
rect 38654 34414 38706 34423
rect 38814 34457 38866 34466
rect 38814 34423 38823 34457
rect 38823 34423 38857 34457
rect 38857 34423 38866 34457
rect 38814 34414 38866 34423
rect 38974 34457 39026 34466
rect 38974 34423 38983 34457
rect 38983 34423 39017 34457
rect 39017 34423 39026 34457
rect 38974 34414 39026 34423
rect 39134 34457 39186 34466
rect 39134 34423 39143 34457
rect 39143 34423 39177 34457
rect 39177 34423 39186 34457
rect 39134 34414 39186 34423
rect 39294 34457 39346 34466
rect 39294 34423 39303 34457
rect 39303 34423 39337 34457
rect 39337 34423 39346 34457
rect 39294 34414 39346 34423
rect 39454 34457 39506 34466
rect 39454 34423 39463 34457
rect 39463 34423 39497 34457
rect 39497 34423 39506 34457
rect 39454 34414 39506 34423
rect 39614 34457 39666 34466
rect 39614 34423 39623 34457
rect 39623 34423 39657 34457
rect 39657 34423 39666 34457
rect 39614 34414 39666 34423
rect 39774 34457 39826 34466
rect 39774 34423 39783 34457
rect 39783 34423 39817 34457
rect 39817 34423 39826 34457
rect 39774 34414 39826 34423
rect 39934 34457 39986 34466
rect 39934 34423 39943 34457
rect 39943 34423 39977 34457
rect 39977 34423 39986 34457
rect 39934 34414 39986 34423
rect 40094 34457 40146 34466
rect 40094 34423 40103 34457
rect 40103 34423 40137 34457
rect 40137 34423 40146 34457
rect 40094 34414 40146 34423
rect 40254 34457 40306 34466
rect 40254 34423 40263 34457
rect 40263 34423 40297 34457
rect 40297 34423 40306 34457
rect 40254 34414 40306 34423
rect 40414 34457 40466 34466
rect 40414 34423 40423 34457
rect 40423 34423 40457 34457
rect 40457 34423 40466 34457
rect 40414 34414 40466 34423
rect 40574 34457 40626 34466
rect 40574 34423 40583 34457
rect 40583 34423 40617 34457
rect 40617 34423 40626 34457
rect 40574 34414 40626 34423
rect 40734 34457 40786 34466
rect 40734 34423 40743 34457
rect 40743 34423 40777 34457
rect 40777 34423 40786 34457
rect 40734 34414 40786 34423
rect 40894 34457 40946 34466
rect 40894 34423 40903 34457
rect 40903 34423 40937 34457
rect 40937 34423 40946 34457
rect 40894 34414 40946 34423
rect 41054 34457 41106 34466
rect 41054 34423 41063 34457
rect 41063 34423 41097 34457
rect 41097 34423 41106 34457
rect 41054 34414 41106 34423
rect 41214 34457 41266 34466
rect 41214 34423 41223 34457
rect 41223 34423 41257 34457
rect 41257 34423 41266 34457
rect 41214 34414 41266 34423
rect 41374 34457 41426 34466
rect 41374 34423 41383 34457
rect 41383 34423 41417 34457
rect 41417 34423 41426 34457
rect 41374 34414 41426 34423
rect 41534 34457 41586 34466
rect 41534 34423 41543 34457
rect 41543 34423 41577 34457
rect 41577 34423 41586 34457
rect 41534 34414 41586 34423
rect 41694 34457 41746 34466
rect 41694 34423 41703 34457
rect 41703 34423 41737 34457
rect 41737 34423 41746 34457
rect 41694 34414 41746 34423
rect 41854 34457 41906 34466
rect 41854 34423 41863 34457
rect 41863 34423 41897 34457
rect 41897 34423 41906 34457
rect 41854 34414 41906 34423
rect 14 34297 66 34306
rect 14 34263 23 34297
rect 23 34263 57 34297
rect 57 34263 66 34297
rect 14 34254 66 34263
rect 174 34297 226 34306
rect 174 34263 183 34297
rect 183 34263 217 34297
rect 217 34263 226 34297
rect 174 34254 226 34263
rect 334 34297 386 34306
rect 334 34263 343 34297
rect 343 34263 377 34297
rect 377 34263 386 34297
rect 334 34254 386 34263
rect 494 34297 546 34306
rect 494 34263 503 34297
rect 503 34263 537 34297
rect 537 34263 546 34297
rect 494 34254 546 34263
rect 654 34297 706 34306
rect 654 34263 663 34297
rect 663 34263 697 34297
rect 697 34263 706 34297
rect 654 34254 706 34263
rect 814 34297 866 34306
rect 814 34263 823 34297
rect 823 34263 857 34297
rect 857 34263 866 34297
rect 814 34254 866 34263
rect 974 34297 1026 34306
rect 974 34263 983 34297
rect 983 34263 1017 34297
rect 1017 34263 1026 34297
rect 974 34254 1026 34263
rect 1134 34297 1186 34306
rect 1134 34263 1143 34297
rect 1143 34263 1177 34297
rect 1177 34263 1186 34297
rect 1134 34254 1186 34263
rect 1294 34297 1346 34306
rect 1294 34263 1303 34297
rect 1303 34263 1337 34297
rect 1337 34263 1346 34297
rect 1294 34254 1346 34263
rect 1454 34297 1506 34306
rect 1454 34263 1463 34297
rect 1463 34263 1497 34297
rect 1497 34263 1506 34297
rect 1454 34254 1506 34263
rect 1614 34297 1666 34306
rect 1614 34263 1623 34297
rect 1623 34263 1657 34297
rect 1657 34263 1666 34297
rect 1614 34254 1666 34263
rect 1774 34297 1826 34306
rect 1774 34263 1783 34297
rect 1783 34263 1817 34297
rect 1817 34263 1826 34297
rect 1774 34254 1826 34263
rect 1934 34297 1986 34306
rect 1934 34263 1943 34297
rect 1943 34263 1977 34297
rect 1977 34263 1986 34297
rect 1934 34254 1986 34263
rect 2094 34297 2146 34306
rect 2094 34263 2103 34297
rect 2103 34263 2137 34297
rect 2137 34263 2146 34297
rect 2094 34254 2146 34263
rect 2254 34297 2306 34306
rect 2254 34263 2263 34297
rect 2263 34263 2297 34297
rect 2297 34263 2306 34297
rect 2254 34254 2306 34263
rect 2414 34297 2466 34306
rect 2414 34263 2423 34297
rect 2423 34263 2457 34297
rect 2457 34263 2466 34297
rect 2414 34254 2466 34263
rect 2574 34297 2626 34306
rect 2574 34263 2583 34297
rect 2583 34263 2617 34297
rect 2617 34263 2626 34297
rect 2574 34254 2626 34263
rect 2734 34297 2786 34306
rect 2734 34263 2743 34297
rect 2743 34263 2777 34297
rect 2777 34263 2786 34297
rect 2734 34254 2786 34263
rect 2894 34297 2946 34306
rect 2894 34263 2903 34297
rect 2903 34263 2937 34297
rect 2937 34263 2946 34297
rect 2894 34254 2946 34263
rect 3054 34297 3106 34306
rect 3054 34263 3063 34297
rect 3063 34263 3097 34297
rect 3097 34263 3106 34297
rect 3054 34254 3106 34263
rect 3214 34297 3266 34306
rect 3214 34263 3223 34297
rect 3223 34263 3257 34297
rect 3257 34263 3266 34297
rect 3214 34254 3266 34263
rect 3374 34297 3426 34306
rect 3374 34263 3383 34297
rect 3383 34263 3417 34297
rect 3417 34263 3426 34297
rect 3374 34254 3426 34263
rect 3534 34297 3586 34306
rect 3534 34263 3543 34297
rect 3543 34263 3577 34297
rect 3577 34263 3586 34297
rect 3534 34254 3586 34263
rect 3694 34297 3746 34306
rect 3694 34263 3703 34297
rect 3703 34263 3737 34297
rect 3737 34263 3746 34297
rect 3694 34254 3746 34263
rect 3854 34297 3906 34306
rect 3854 34263 3863 34297
rect 3863 34263 3897 34297
rect 3897 34263 3906 34297
rect 3854 34254 3906 34263
rect 4014 34297 4066 34306
rect 4014 34263 4023 34297
rect 4023 34263 4057 34297
rect 4057 34263 4066 34297
rect 4014 34254 4066 34263
rect 4174 34297 4226 34306
rect 4174 34263 4183 34297
rect 4183 34263 4217 34297
rect 4217 34263 4226 34297
rect 4174 34254 4226 34263
rect 4334 34297 4386 34306
rect 4334 34263 4343 34297
rect 4343 34263 4377 34297
rect 4377 34263 4386 34297
rect 4334 34254 4386 34263
rect 4494 34297 4546 34306
rect 4494 34263 4503 34297
rect 4503 34263 4537 34297
rect 4537 34263 4546 34297
rect 4494 34254 4546 34263
rect 4654 34297 4706 34306
rect 4654 34263 4663 34297
rect 4663 34263 4697 34297
rect 4697 34263 4706 34297
rect 4654 34254 4706 34263
rect 4814 34297 4866 34306
rect 4814 34263 4823 34297
rect 4823 34263 4857 34297
rect 4857 34263 4866 34297
rect 4814 34254 4866 34263
rect 4974 34297 5026 34306
rect 4974 34263 4983 34297
rect 4983 34263 5017 34297
rect 5017 34263 5026 34297
rect 4974 34254 5026 34263
rect 5134 34297 5186 34306
rect 5134 34263 5143 34297
rect 5143 34263 5177 34297
rect 5177 34263 5186 34297
rect 5134 34254 5186 34263
rect 5294 34297 5346 34306
rect 5294 34263 5303 34297
rect 5303 34263 5337 34297
rect 5337 34263 5346 34297
rect 5294 34254 5346 34263
rect 5454 34297 5506 34306
rect 5454 34263 5463 34297
rect 5463 34263 5497 34297
rect 5497 34263 5506 34297
rect 5454 34254 5506 34263
rect 5614 34297 5666 34306
rect 5614 34263 5623 34297
rect 5623 34263 5657 34297
rect 5657 34263 5666 34297
rect 5614 34254 5666 34263
rect 5774 34297 5826 34306
rect 5774 34263 5783 34297
rect 5783 34263 5817 34297
rect 5817 34263 5826 34297
rect 5774 34254 5826 34263
rect 5934 34297 5986 34306
rect 5934 34263 5943 34297
rect 5943 34263 5977 34297
rect 5977 34263 5986 34297
rect 5934 34254 5986 34263
rect 6094 34297 6146 34306
rect 6094 34263 6103 34297
rect 6103 34263 6137 34297
rect 6137 34263 6146 34297
rect 6094 34254 6146 34263
rect 6254 34297 6306 34306
rect 6254 34263 6263 34297
rect 6263 34263 6297 34297
rect 6297 34263 6306 34297
rect 6254 34254 6306 34263
rect 6414 34297 6466 34306
rect 6414 34263 6423 34297
rect 6423 34263 6457 34297
rect 6457 34263 6466 34297
rect 6414 34254 6466 34263
rect 6574 34297 6626 34306
rect 6574 34263 6583 34297
rect 6583 34263 6617 34297
rect 6617 34263 6626 34297
rect 6574 34254 6626 34263
rect 6734 34297 6786 34306
rect 6734 34263 6743 34297
rect 6743 34263 6777 34297
rect 6777 34263 6786 34297
rect 6734 34254 6786 34263
rect 6894 34297 6946 34306
rect 6894 34263 6903 34297
rect 6903 34263 6937 34297
rect 6937 34263 6946 34297
rect 6894 34254 6946 34263
rect 7054 34297 7106 34306
rect 7054 34263 7063 34297
rect 7063 34263 7097 34297
rect 7097 34263 7106 34297
rect 7054 34254 7106 34263
rect 7214 34297 7266 34306
rect 7214 34263 7223 34297
rect 7223 34263 7257 34297
rect 7257 34263 7266 34297
rect 7214 34254 7266 34263
rect 7374 34297 7426 34306
rect 7374 34263 7383 34297
rect 7383 34263 7417 34297
rect 7417 34263 7426 34297
rect 7374 34254 7426 34263
rect 7534 34297 7586 34306
rect 7534 34263 7543 34297
rect 7543 34263 7577 34297
rect 7577 34263 7586 34297
rect 7534 34254 7586 34263
rect 7694 34297 7746 34306
rect 7694 34263 7703 34297
rect 7703 34263 7737 34297
rect 7737 34263 7746 34297
rect 7694 34254 7746 34263
rect 7854 34297 7906 34306
rect 7854 34263 7863 34297
rect 7863 34263 7897 34297
rect 7897 34263 7906 34297
rect 7854 34254 7906 34263
rect 8014 34297 8066 34306
rect 8014 34263 8023 34297
rect 8023 34263 8057 34297
rect 8057 34263 8066 34297
rect 8014 34254 8066 34263
rect 8174 34297 8226 34306
rect 8174 34263 8183 34297
rect 8183 34263 8217 34297
rect 8217 34263 8226 34297
rect 8174 34254 8226 34263
rect 8334 34297 8386 34306
rect 8334 34263 8343 34297
rect 8343 34263 8377 34297
rect 8377 34263 8386 34297
rect 8334 34254 8386 34263
rect 12494 34297 12546 34306
rect 12494 34263 12503 34297
rect 12503 34263 12537 34297
rect 12537 34263 12546 34297
rect 12494 34254 12546 34263
rect 12654 34297 12706 34306
rect 12654 34263 12663 34297
rect 12663 34263 12697 34297
rect 12697 34263 12706 34297
rect 12654 34254 12706 34263
rect 12814 34297 12866 34306
rect 12814 34263 12823 34297
rect 12823 34263 12857 34297
rect 12857 34263 12866 34297
rect 12814 34254 12866 34263
rect 12974 34297 13026 34306
rect 12974 34263 12983 34297
rect 12983 34263 13017 34297
rect 13017 34263 13026 34297
rect 12974 34254 13026 34263
rect 13134 34297 13186 34306
rect 13134 34263 13143 34297
rect 13143 34263 13177 34297
rect 13177 34263 13186 34297
rect 13134 34254 13186 34263
rect 13294 34297 13346 34306
rect 13294 34263 13303 34297
rect 13303 34263 13337 34297
rect 13337 34263 13346 34297
rect 13294 34254 13346 34263
rect 13454 34297 13506 34306
rect 13454 34263 13463 34297
rect 13463 34263 13497 34297
rect 13497 34263 13506 34297
rect 13454 34254 13506 34263
rect 13614 34297 13666 34306
rect 13614 34263 13623 34297
rect 13623 34263 13657 34297
rect 13657 34263 13666 34297
rect 13614 34254 13666 34263
rect 13774 34297 13826 34306
rect 13774 34263 13783 34297
rect 13783 34263 13817 34297
rect 13817 34263 13826 34297
rect 13774 34254 13826 34263
rect 13934 34297 13986 34306
rect 13934 34263 13943 34297
rect 13943 34263 13977 34297
rect 13977 34263 13986 34297
rect 13934 34254 13986 34263
rect 14094 34297 14146 34306
rect 14094 34263 14103 34297
rect 14103 34263 14137 34297
rect 14137 34263 14146 34297
rect 14094 34254 14146 34263
rect 14254 34297 14306 34306
rect 14254 34263 14263 34297
rect 14263 34263 14297 34297
rect 14297 34263 14306 34297
rect 14254 34254 14306 34263
rect 14414 34297 14466 34306
rect 14414 34263 14423 34297
rect 14423 34263 14457 34297
rect 14457 34263 14466 34297
rect 14414 34254 14466 34263
rect 14574 34297 14626 34306
rect 14574 34263 14583 34297
rect 14583 34263 14617 34297
rect 14617 34263 14626 34297
rect 14574 34254 14626 34263
rect 14734 34297 14786 34306
rect 14734 34263 14743 34297
rect 14743 34263 14777 34297
rect 14777 34263 14786 34297
rect 14734 34254 14786 34263
rect 14894 34297 14946 34306
rect 14894 34263 14903 34297
rect 14903 34263 14937 34297
rect 14937 34263 14946 34297
rect 14894 34254 14946 34263
rect 15054 34297 15106 34306
rect 15054 34263 15063 34297
rect 15063 34263 15097 34297
rect 15097 34263 15106 34297
rect 15054 34254 15106 34263
rect 15214 34297 15266 34306
rect 15214 34263 15223 34297
rect 15223 34263 15257 34297
rect 15257 34263 15266 34297
rect 15214 34254 15266 34263
rect 15374 34297 15426 34306
rect 15374 34263 15383 34297
rect 15383 34263 15417 34297
rect 15417 34263 15426 34297
rect 15374 34254 15426 34263
rect 15534 34297 15586 34306
rect 15534 34263 15543 34297
rect 15543 34263 15577 34297
rect 15577 34263 15586 34297
rect 15534 34254 15586 34263
rect 15694 34297 15746 34306
rect 15694 34263 15703 34297
rect 15703 34263 15737 34297
rect 15737 34263 15746 34297
rect 15694 34254 15746 34263
rect 15854 34297 15906 34306
rect 15854 34263 15863 34297
rect 15863 34263 15897 34297
rect 15897 34263 15906 34297
rect 15854 34254 15906 34263
rect 16014 34297 16066 34306
rect 16014 34263 16023 34297
rect 16023 34263 16057 34297
rect 16057 34263 16066 34297
rect 16014 34254 16066 34263
rect 16174 34297 16226 34306
rect 16174 34263 16183 34297
rect 16183 34263 16217 34297
rect 16217 34263 16226 34297
rect 16174 34254 16226 34263
rect 16334 34297 16386 34306
rect 16334 34263 16343 34297
rect 16343 34263 16377 34297
rect 16377 34263 16386 34297
rect 16334 34254 16386 34263
rect 16494 34297 16546 34306
rect 16494 34263 16503 34297
rect 16503 34263 16537 34297
rect 16537 34263 16546 34297
rect 16494 34254 16546 34263
rect 16654 34297 16706 34306
rect 16654 34263 16663 34297
rect 16663 34263 16697 34297
rect 16697 34263 16706 34297
rect 16654 34254 16706 34263
rect 16814 34297 16866 34306
rect 16814 34263 16823 34297
rect 16823 34263 16857 34297
rect 16857 34263 16866 34297
rect 16814 34254 16866 34263
rect 16974 34297 17026 34306
rect 16974 34263 16983 34297
rect 16983 34263 17017 34297
rect 17017 34263 17026 34297
rect 16974 34254 17026 34263
rect 17134 34297 17186 34306
rect 17134 34263 17143 34297
rect 17143 34263 17177 34297
rect 17177 34263 17186 34297
rect 17134 34254 17186 34263
rect 17294 34297 17346 34306
rect 17294 34263 17303 34297
rect 17303 34263 17337 34297
rect 17337 34263 17346 34297
rect 17294 34254 17346 34263
rect 17454 34297 17506 34306
rect 17454 34263 17463 34297
rect 17463 34263 17497 34297
rect 17497 34263 17506 34297
rect 17454 34254 17506 34263
rect 17614 34297 17666 34306
rect 17614 34263 17623 34297
rect 17623 34263 17657 34297
rect 17657 34263 17666 34297
rect 17614 34254 17666 34263
rect 17774 34297 17826 34306
rect 17774 34263 17783 34297
rect 17783 34263 17817 34297
rect 17817 34263 17826 34297
rect 17774 34254 17826 34263
rect 17934 34297 17986 34306
rect 17934 34263 17943 34297
rect 17943 34263 17977 34297
rect 17977 34263 17986 34297
rect 17934 34254 17986 34263
rect 18094 34297 18146 34306
rect 18094 34263 18103 34297
rect 18103 34263 18137 34297
rect 18137 34263 18146 34297
rect 18094 34254 18146 34263
rect 18254 34297 18306 34306
rect 18254 34263 18263 34297
rect 18263 34263 18297 34297
rect 18297 34263 18306 34297
rect 18254 34254 18306 34263
rect 18414 34297 18466 34306
rect 18414 34263 18423 34297
rect 18423 34263 18457 34297
rect 18457 34263 18466 34297
rect 18414 34254 18466 34263
rect 18574 34297 18626 34306
rect 18574 34263 18583 34297
rect 18583 34263 18617 34297
rect 18617 34263 18626 34297
rect 18574 34254 18626 34263
rect 18734 34297 18786 34306
rect 18734 34263 18743 34297
rect 18743 34263 18777 34297
rect 18777 34263 18786 34297
rect 18734 34254 18786 34263
rect 18894 34297 18946 34306
rect 18894 34263 18903 34297
rect 18903 34263 18937 34297
rect 18937 34263 18946 34297
rect 18894 34254 18946 34263
rect 23134 34297 23186 34306
rect 23134 34263 23143 34297
rect 23143 34263 23177 34297
rect 23177 34263 23186 34297
rect 23134 34254 23186 34263
rect 23294 34297 23346 34306
rect 23294 34263 23303 34297
rect 23303 34263 23337 34297
rect 23337 34263 23346 34297
rect 23294 34254 23346 34263
rect 23454 34297 23506 34306
rect 23454 34263 23463 34297
rect 23463 34263 23497 34297
rect 23497 34263 23506 34297
rect 23454 34254 23506 34263
rect 23614 34297 23666 34306
rect 23614 34263 23623 34297
rect 23623 34263 23657 34297
rect 23657 34263 23666 34297
rect 23614 34254 23666 34263
rect 23774 34297 23826 34306
rect 23774 34263 23783 34297
rect 23783 34263 23817 34297
rect 23817 34263 23826 34297
rect 23774 34254 23826 34263
rect 23934 34297 23986 34306
rect 23934 34263 23943 34297
rect 23943 34263 23977 34297
rect 23977 34263 23986 34297
rect 23934 34254 23986 34263
rect 24094 34297 24146 34306
rect 24094 34263 24103 34297
rect 24103 34263 24137 34297
rect 24137 34263 24146 34297
rect 24094 34254 24146 34263
rect 24254 34297 24306 34306
rect 24254 34263 24263 34297
rect 24263 34263 24297 34297
rect 24297 34263 24306 34297
rect 24254 34254 24306 34263
rect 24414 34297 24466 34306
rect 24414 34263 24423 34297
rect 24423 34263 24457 34297
rect 24457 34263 24466 34297
rect 24414 34254 24466 34263
rect 24574 34297 24626 34306
rect 24574 34263 24583 34297
rect 24583 34263 24617 34297
rect 24617 34263 24626 34297
rect 24574 34254 24626 34263
rect 24734 34297 24786 34306
rect 24734 34263 24743 34297
rect 24743 34263 24777 34297
rect 24777 34263 24786 34297
rect 24734 34254 24786 34263
rect 24894 34297 24946 34306
rect 24894 34263 24903 34297
rect 24903 34263 24937 34297
rect 24937 34263 24946 34297
rect 24894 34254 24946 34263
rect 25054 34297 25106 34306
rect 25054 34263 25063 34297
rect 25063 34263 25097 34297
rect 25097 34263 25106 34297
rect 25054 34254 25106 34263
rect 25214 34297 25266 34306
rect 25214 34263 25223 34297
rect 25223 34263 25257 34297
rect 25257 34263 25266 34297
rect 25214 34254 25266 34263
rect 25374 34297 25426 34306
rect 25374 34263 25383 34297
rect 25383 34263 25417 34297
rect 25417 34263 25426 34297
rect 25374 34254 25426 34263
rect 25534 34297 25586 34306
rect 25534 34263 25543 34297
rect 25543 34263 25577 34297
rect 25577 34263 25586 34297
rect 25534 34254 25586 34263
rect 25694 34297 25746 34306
rect 25694 34263 25703 34297
rect 25703 34263 25737 34297
rect 25737 34263 25746 34297
rect 25694 34254 25746 34263
rect 25854 34297 25906 34306
rect 25854 34263 25863 34297
rect 25863 34263 25897 34297
rect 25897 34263 25906 34297
rect 25854 34254 25906 34263
rect 26014 34297 26066 34306
rect 26014 34263 26023 34297
rect 26023 34263 26057 34297
rect 26057 34263 26066 34297
rect 26014 34254 26066 34263
rect 26174 34297 26226 34306
rect 26174 34263 26183 34297
rect 26183 34263 26217 34297
rect 26217 34263 26226 34297
rect 26174 34254 26226 34263
rect 26334 34297 26386 34306
rect 26334 34263 26343 34297
rect 26343 34263 26377 34297
rect 26377 34263 26386 34297
rect 26334 34254 26386 34263
rect 26494 34297 26546 34306
rect 26494 34263 26503 34297
rect 26503 34263 26537 34297
rect 26537 34263 26546 34297
rect 26494 34254 26546 34263
rect 26654 34297 26706 34306
rect 26654 34263 26663 34297
rect 26663 34263 26697 34297
rect 26697 34263 26706 34297
rect 26654 34254 26706 34263
rect 26814 34297 26866 34306
rect 26814 34263 26823 34297
rect 26823 34263 26857 34297
rect 26857 34263 26866 34297
rect 26814 34254 26866 34263
rect 26974 34297 27026 34306
rect 26974 34263 26983 34297
rect 26983 34263 27017 34297
rect 27017 34263 27026 34297
rect 26974 34254 27026 34263
rect 27134 34297 27186 34306
rect 27134 34263 27143 34297
rect 27143 34263 27177 34297
rect 27177 34263 27186 34297
rect 27134 34254 27186 34263
rect 27294 34297 27346 34306
rect 27294 34263 27303 34297
rect 27303 34263 27337 34297
rect 27337 34263 27346 34297
rect 27294 34254 27346 34263
rect 27454 34297 27506 34306
rect 27454 34263 27463 34297
rect 27463 34263 27497 34297
rect 27497 34263 27506 34297
rect 27454 34254 27506 34263
rect 27614 34297 27666 34306
rect 27614 34263 27623 34297
rect 27623 34263 27657 34297
rect 27657 34263 27666 34297
rect 27614 34254 27666 34263
rect 27774 34297 27826 34306
rect 27774 34263 27783 34297
rect 27783 34263 27817 34297
rect 27817 34263 27826 34297
rect 27774 34254 27826 34263
rect 27934 34297 27986 34306
rect 27934 34263 27943 34297
rect 27943 34263 27977 34297
rect 27977 34263 27986 34297
rect 27934 34254 27986 34263
rect 28094 34297 28146 34306
rect 28094 34263 28103 34297
rect 28103 34263 28137 34297
rect 28137 34263 28146 34297
rect 28094 34254 28146 34263
rect 28254 34297 28306 34306
rect 28254 34263 28263 34297
rect 28263 34263 28297 34297
rect 28297 34263 28306 34297
rect 28254 34254 28306 34263
rect 28414 34297 28466 34306
rect 28414 34263 28423 34297
rect 28423 34263 28457 34297
rect 28457 34263 28466 34297
rect 28414 34254 28466 34263
rect 28574 34297 28626 34306
rect 28574 34263 28583 34297
rect 28583 34263 28617 34297
rect 28617 34263 28626 34297
rect 28574 34254 28626 34263
rect 28734 34297 28786 34306
rect 28734 34263 28743 34297
rect 28743 34263 28777 34297
rect 28777 34263 28786 34297
rect 28734 34254 28786 34263
rect 28894 34297 28946 34306
rect 28894 34263 28903 34297
rect 28903 34263 28937 34297
rect 28937 34263 28946 34297
rect 28894 34254 28946 34263
rect 29054 34297 29106 34306
rect 29054 34263 29063 34297
rect 29063 34263 29097 34297
rect 29097 34263 29106 34297
rect 29054 34254 29106 34263
rect 29214 34297 29266 34306
rect 29214 34263 29223 34297
rect 29223 34263 29257 34297
rect 29257 34263 29266 34297
rect 29214 34254 29266 34263
rect 29374 34297 29426 34306
rect 29374 34263 29383 34297
rect 29383 34263 29417 34297
rect 29417 34263 29426 34297
rect 29374 34254 29426 34263
rect 33534 34297 33586 34306
rect 33534 34263 33543 34297
rect 33543 34263 33577 34297
rect 33577 34263 33586 34297
rect 33534 34254 33586 34263
rect 33694 34297 33746 34306
rect 33694 34263 33703 34297
rect 33703 34263 33737 34297
rect 33737 34263 33746 34297
rect 33694 34254 33746 34263
rect 33854 34297 33906 34306
rect 33854 34263 33863 34297
rect 33863 34263 33897 34297
rect 33897 34263 33906 34297
rect 33854 34254 33906 34263
rect 34014 34297 34066 34306
rect 34014 34263 34023 34297
rect 34023 34263 34057 34297
rect 34057 34263 34066 34297
rect 34014 34254 34066 34263
rect 34174 34297 34226 34306
rect 34174 34263 34183 34297
rect 34183 34263 34217 34297
rect 34217 34263 34226 34297
rect 34174 34254 34226 34263
rect 34334 34297 34386 34306
rect 34334 34263 34343 34297
rect 34343 34263 34377 34297
rect 34377 34263 34386 34297
rect 34334 34254 34386 34263
rect 34494 34297 34546 34306
rect 34494 34263 34503 34297
rect 34503 34263 34537 34297
rect 34537 34263 34546 34297
rect 34494 34254 34546 34263
rect 34654 34297 34706 34306
rect 34654 34263 34663 34297
rect 34663 34263 34697 34297
rect 34697 34263 34706 34297
rect 34654 34254 34706 34263
rect 34814 34297 34866 34306
rect 34814 34263 34823 34297
rect 34823 34263 34857 34297
rect 34857 34263 34866 34297
rect 34814 34254 34866 34263
rect 34974 34297 35026 34306
rect 34974 34263 34983 34297
rect 34983 34263 35017 34297
rect 35017 34263 35026 34297
rect 34974 34254 35026 34263
rect 35134 34297 35186 34306
rect 35134 34263 35143 34297
rect 35143 34263 35177 34297
rect 35177 34263 35186 34297
rect 35134 34254 35186 34263
rect 35294 34297 35346 34306
rect 35294 34263 35303 34297
rect 35303 34263 35337 34297
rect 35337 34263 35346 34297
rect 35294 34254 35346 34263
rect 35454 34297 35506 34306
rect 35454 34263 35463 34297
rect 35463 34263 35497 34297
rect 35497 34263 35506 34297
rect 35454 34254 35506 34263
rect 35614 34297 35666 34306
rect 35614 34263 35623 34297
rect 35623 34263 35657 34297
rect 35657 34263 35666 34297
rect 35614 34254 35666 34263
rect 35774 34297 35826 34306
rect 35774 34263 35783 34297
rect 35783 34263 35817 34297
rect 35817 34263 35826 34297
rect 35774 34254 35826 34263
rect 35934 34297 35986 34306
rect 35934 34263 35943 34297
rect 35943 34263 35977 34297
rect 35977 34263 35986 34297
rect 35934 34254 35986 34263
rect 36094 34297 36146 34306
rect 36094 34263 36103 34297
rect 36103 34263 36137 34297
rect 36137 34263 36146 34297
rect 36094 34254 36146 34263
rect 36254 34297 36306 34306
rect 36254 34263 36263 34297
rect 36263 34263 36297 34297
rect 36297 34263 36306 34297
rect 36254 34254 36306 34263
rect 36414 34297 36466 34306
rect 36414 34263 36423 34297
rect 36423 34263 36457 34297
rect 36457 34263 36466 34297
rect 36414 34254 36466 34263
rect 36574 34297 36626 34306
rect 36574 34263 36583 34297
rect 36583 34263 36617 34297
rect 36617 34263 36626 34297
rect 36574 34254 36626 34263
rect 36734 34297 36786 34306
rect 36734 34263 36743 34297
rect 36743 34263 36777 34297
rect 36777 34263 36786 34297
rect 36734 34254 36786 34263
rect 36894 34297 36946 34306
rect 36894 34263 36903 34297
rect 36903 34263 36937 34297
rect 36937 34263 36946 34297
rect 36894 34254 36946 34263
rect 37054 34297 37106 34306
rect 37054 34263 37063 34297
rect 37063 34263 37097 34297
rect 37097 34263 37106 34297
rect 37054 34254 37106 34263
rect 37214 34297 37266 34306
rect 37214 34263 37223 34297
rect 37223 34263 37257 34297
rect 37257 34263 37266 34297
rect 37214 34254 37266 34263
rect 37374 34297 37426 34306
rect 37374 34263 37383 34297
rect 37383 34263 37417 34297
rect 37417 34263 37426 34297
rect 37374 34254 37426 34263
rect 37534 34297 37586 34306
rect 37534 34263 37543 34297
rect 37543 34263 37577 34297
rect 37577 34263 37586 34297
rect 37534 34254 37586 34263
rect 37694 34297 37746 34306
rect 37694 34263 37703 34297
rect 37703 34263 37737 34297
rect 37737 34263 37746 34297
rect 37694 34254 37746 34263
rect 37854 34297 37906 34306
rect 37854 34263 37863 34297
rect 37863 34263 37897 34297
rect 37897 34263 37906 34297
rect 37854 34254 37906 34263
rect 38014 34297 38066 34306
rect 38014 34263 38023 34297
rect 38023 34263 38057 34297
rect 38057 34263 38066 34297
rect 38014 34254 38066 34263
rect 38174 34297 38226 34306
rect 38174 34263 38183 34297
rect 38183 34263 38217 34297
rect 38217 34263 38226 34297
rect 38174 34254 38226 34263
rect 38334 34297 38386 34306
rect 38334 34263 38343 34297
rect 38343 34263 38377 34297
rect 38377 34263 38386 34297
rect 38334 34254 38386 34263
rect 38494 34297 38546 34306
rect 38494 34263 38503 34297
rect 38503 34263 38537 34297
rect 38537 34263 38546 34297
rect 38494 34254 38546 34263
rect 38654 34297 38706 34306
rect 38654 34263 38663 34297
rect 38663 34263 38697 34297
rect 38697 34263 38706 34297
rect 38654 34254 38706 34263
rect 38814 34297 38866 34306
rect 38814 34263 38823 34297
rect 38823 34263 38857 34297
rect 38857 34263 38866 34297
rect 38814 34254 38866 34263
rect 38974 34297 39026 34306
rect 38974 34263 38983 34297
rect 38983 34263 39017 34297
rect 39017 34263 39026 34297
rect 38974 34254 39026 34263
rect 39134 34297 39186 34306
rect 39134 34263 39143 34297
rect 39143 34263 39177 34297
rect 39177 34263 39186 34297
rect 39134 34254 39186 34263
rect 39294 34297 39346 34306
rect 39294 34263 39303 34297
rect 39303 34263 39337 34297
rect 39337 34263 39346 34297
rect 39294 34254 39346 34263
rect 39454 34297 39506 34306
rect 39454 34263 39463 34297
rect 39463 34263 39497 34297
rect 39497 34263 39506 34297
rect 39454 34254 39506 34263
rect 39614 34297 39666 34306
rect 39614 34263 39623 34297
rect 39623 34263 39657 34297
rect 39657 34263 39666 34297
rect 39614 34254 39666 34263
rect 39774 34297 39826 34306
rect 39774 34263 39783 34297
rect 39783 34263 39817 34297
rect 39817 34263 39826 34297
rect 39774 34254 39826 34263
rect 39934 34297 39986 34306
rect 39934 34263 39943 34297
rect 39943 34263 39977 34297
rect 39977 34263 39986 34297
rect 39934 34254 39986 34263
rect 40094 34297 40146 34306
rect 40094 34263 40103 34297
rect 40103 34263 40137 34297
rect 40137 34263 40146 34297
rect 40094 34254 40146 34263
rect 40254 34297 40306 34306
rect 40254 34263 40263 34297
rect 40263 34263 40297 34297
rect 40297 34263 40306 34297
rect 40254 34254 40306 34263
rect 40414 34297 40466 34306
rect 40414 34263 40423 34297
rect 40423 34263 40457 34297
rect 40457 34263 40466 34297
rect 40414 34254 40466 34263
rect 40574 34297 40626 34306
rect 40574 34263 40583 34297
rect 40583 34263 40617 34297
rect 40617 34263 40626 34297
rect 40574 34254 40626 34263
rect 40734 34297 40786 34306
rect 40734 34263 40743 34297
rect 40743 34263 40777 34297
rect 40777 34263 40786 34297
rect 40734 34254 40786 34263
rect 40894 34297 40946 34306
rect 40894 34263 40903 34297
rect 40903 34263 40937 34297
rect 40937 34263 40946 34297
rect 40894 34254 40946 34263
rect 41054 34297 41106 34306
rect 41054 34263 41063 34297
rect 41063 34263 41097 34297
rect 41097 34263 41106 34297
rect 41054 34254 41106 34263
rect 41214 34297 41266 34306
rect 41214 34263 41223 34297
rect 41223 34263 41257 34297
rect 41257 34263 41266 34297
rect 41214 34254 41266 34263
rect 41374 34297 41426 34306
rect 41374 34263 41383 34297
rect 41383 34263 41417 34297
rect 41417 34263 41426 34297
rect 41374 34254 41426 34263
rect 41534 34297 41586 34306
rect 41534 34263 41543 34297
rect 41543 34263 41577 34297
rect 41577 34263 41586 34297
rect 41534 34254 41586 34263
rect 41694 34297 41746 34306
rect 41694 34263 41703 34297
rect 41703 34263 41737 34297
rect 41737 34263 41746 34297
rect 41694 34254 41746 34263
rect 41854 34297 41906 34306
rect 41854 34263 41863 34297
rect 41863 34263 41897 34297
rect 41897 34263 41906 34297
rect 41854 34254 41906 34263
rect 14 33977 66 33986
rect 14 33943 23 33977
rect 23 33943 57 33977
rect 57 33943 66 33977
rect 14 33934 66 33943
rect 174 33977 226 33986
rect 174 33943 183 33977
rect 183 33943 217 33977
rect 217 33943 226 33977
rect 174 33934 226 33943
rect 334 33977 386 33986
rect 334 33943 343 33977
rect 343 33943 377 33977
rect 377 33943 386 33977
rect 334 33934 386 33943
rect 494 33977 546 33986
rect 494 33943 503 33977
rect 503 33943 537 33977
rect 537 33943 546 33977
rect 494 33934 546 33943
rect 654 33977 706 33986
rect 654 33943 663 33977
rect 663 33943 697 33977
rect 697 33943 706 33977
rect 654 33934 706 33943
rect 814 33977 866 33986
rect 814 33943 823 33977
rect 823 33943 857 33977
rect 857 33943 866 33977
rect 814 33934 866 33943
rect 974 33977 1026 33986
rect 974 33943 983 33977
rect 983 33943 1017 33977
rect 1017 33943 1026 33977
rect 974 33934 1026 33943
rect 1134 33977 1186 33986
rect 1134 33943 1143 33977
rect 1143 33943 1177 33977
rect 1177 33943 1186 33977
rect 1134 33934 1186 33943
rect 1294 33977 1346 33986
rect 1294 33943 1303 33977
rect 1303 33943 1337 33977
rect 1337 33943 1346 33977
rect 1294 33934 1346 33943
rect 1454 33977 1506 33986
rect 1454 33943 1463 33977
rect 1463 33943 1497 33977
rect 1497 33943 1506 33977
rect 1454 33934 1506 33943
rect 1614 33977 1666 33986
rect 1614 33943 1623 33977
rect 1623 33943 1657 33977
rect 1657 33943 1666 33977
rect 1614 33934 1666 33943
rect 1774 33977 1826 33986
rect 1774 33943 1783 33977
rect 1783 33943 1817 33977
rect 1817 33943 1826 33977
rect 1774 33934 1826 33943
rect 1934 33977 1986 33986
rect 1934 33943 1943 33977
rect 1943 33943 1977 33977
rect 1977 33943 1986 33977
rect 1934 33934 1986 33943
rect 2094 33977 2146 33986
rect 2094 33943 2103 33977
rect 2103 33943 2137 33977
rect 2137 33943 2146 33977
rect 2094 33934 2146 33943
rect 2254 33977 2306 33986
rect 2254 33943 2263 33977
rect 2263 33943 2297 33977
rect 2297 33943 2306 33977
rect 2254 33934 2306 33943
rect 2414 33977 2466 33986
rect 2414 33943 2423 33977
rect 2423 33943 2457 33977
rect 2457 33943 2466 33977
rect 2414 33934 2466 33943
rect 2574 33977 2626 33986
rect 2574 33943 2583 33977
rect 2583 33943 2617 33977
rect 2617 33943 2626 33977
rect 2574 33934 2626 33943
rect 2734 33977 2786 33986
rect 2734 33943 2743 33977
rect 2743 33943 2777 33977
rect 2777 33943 2786 33977
rect 2734 33934 2786 33943
rect 2894 33977 2946 33986
rect 2894 33943 2903 33977
rect 2903 33943 2937 33977
rect 2937 33943 2946 33977
rect 2894 33934 2946 33943
rect 3054 33977 3106 33986
rect 3054 33943 3063 33977
rect 3063 33943 3097 33977
rect 3097 33943 3106 33977
rect 3054 33934 3106 33943
rect 3214 33977 3266 33986
rect 3214 33943 3223 33977
rect 3223 33943 3257 33977
rect 3257 33943 3266 33977
rect 3214 33934 3266 33943
rect 3374 33977 3426 33986
rect 3374 33943 3383 33977
rect 3383 33943 3417 33977
rect 3417 33943 3426 33977
rect 3374 33934 3426 33943
rect 3534 33977 3586 33986
rect 3534 33943 3543 33977
rect 3543 33943 3577 33977
rect 3577 33943 3586 33977
rect 3534 33934 3586 33943
rect 3694 33977 3746 33986
rect 3694 33943 3703 33977
rect 3703 33943 3737 33977
rect 3737 33943 3746 33977
rect 3694 33934 3746 33943
rect 3854 33977 3906 33986
rect 3854 33943 3863 33977
rect 3863 33943 3897 33977
rect 3897 33943 3906 33977
rect 3854 33934 3906 33943
rect 4014 33977 4066 33986
rect 4014 33943 4023 33977
rect 4023 33943 4057 33977
rect 4057 33943 4066 33977
rect 4014 33934 4066 33943
rect 4174 33977 4226 33986
rect 4174 33943 4183 33977
rect 4183 33943 4217 33977
rect 4217 33943 4226 33977
rect 4174 33934 4226 33943
rect 4334 33977 4386 33986
rect 4334 33943 4343 33977
rect 4343 33943 4377 33977
rect 4377 33943 4386 33977
rect 4334 33934 4386 33943
rect 4494 33977 4546 33986
rect 4494 33943 4503 33977
rect 4503 33943 4537 33977
rect 4537 33943 4546 33977
rect 4494 33934 4546 33943
rect 4654 33977 4706 33986
rect 4654 33943 4663 33977
rect 4663 33943 4697 33977
rect 4697 33943 4706 33977
rect 4654 33934 4706 33943
rect 4814 33977 4866 33986
rect 4814 33943 4823 33977
rect 4823 33943 4857 33977
rect 4857 33943 4866 33977
rect 4814 33934 4866 33943
rect 4974 33977 5026 33986
rect 4974 33943 4983 33977
rect 4983 33943 5017 33977
rect 5017 33943 5026 33977
rect 4974 33934 5026 33943
rect 5134 33977 5186 33986
rect 5134 33943 5143 33977
rect 5143 33943 5177 33977
rect 5177 33943 5186 33977
rect 5134 33934 5186 33943
rect 5294 33977 5346 33986
rect 5294 33943 5303 33977
rect 5303 33943 5337 33977
rect 5337 33943 5346 33977
rect 5294 33934 5346 33943
rect 5454 33977 5506 33986
rect 5454 33943 5463 33977
rect 5463 33943 5497 33977
rect 5497 33943 5506 33977
rect 5454 33934 5506 33943
rect 5614 33977 5666 33986
rect 5614 33943 5623 33977
rect 5623 33943 5657 33977
rect 5657 33943 5666 33977
rect 5614 33934 5666 33943
rect 5774 33977 5826 33986
rect 5774 33943 5783 33977
rect 5783 33943 5817 33977
rect 5817 33943 5826 33977
rect 5774 33934 5826 33943
rect 5934 33977 5986 33986
rect 5934 33943 5943 33977
rect 5943 33943 5977 33977
rect 5977 33943 5986 33977
rect 5934 33934 5986 33943
rect 6094 33977 6146 33986
rect 6094 33943 6103 33977
rect 6103 33943 6137 33977
rect 6137 33943 6146 33977
rect 6094 33934 6146 33943
rect 6254 33977 6306 33986
rect 6254 33943 6263 33977
rect 6263 33943 6297 33977
rect 6297 33943 6306 33977
rect 6254 33934 6306 33943
rect 6414 33977 6466 33986
rect 6414 33943 6423 33977
rect 6423 33943 6457 33977
rect 6457 33943 6466 33977
rect 6414 33934 6466 33943
rect 6574 33977 6626 33986
rect 6574 33943 6583 33977
rect 6583 33943 6617 33977
rect 6617 33943 6626 33977
rect 6574 33934 6626 33943
rect 6734 33977 6786 33986
rect 6734 33943 6743 33977
rect 6743 33943 6777 33977
rect 6777 33943 6786 33977
rect 6734 33934 6786 33943
rect 6894 33977 6946 33986
rect 6894 33943 6903 33977
rect 6903 33943 6937 33977
rect 6937 33943 6946 33977
rect 6894 33934 6946 33943
rect 7054 33977 7106 33986
rect 7054 33943 7063 33977
rect 7063 33943 7097 33977
rect 7097 33943 7106 33977
rect 7054 33934 7106 33943
rect 7214 33977 7266 33986
rect 7214 33943 7223 33977
rect 7223 33943 7257 33977
rect 7257 33943 7266 33977
rect 7214 33934 7266 33943
rect 7374 33977 7426 33986
rect 7374 33943 7383 33977
rect 7383 33943 7417 33977
rect 7417 33943 7426 33977
rect 7374 33934 7426 33943
rect 7534 33977 7586 33986
rect 7534 33943 7543 33977
rect 7543 33943 7577 33977
rect 7577 33943 7586 33977
rect 7534 33934 7586 33943
rect 7694 33977 7746 33986
rect 7694 33943 7703 33977
rect 7703 33943 7737 33977
rect 7737 33943 7746 33977
rect 7694 33934 7746 33943
rect 7854 33977 7906 33986
rect 7854 33943 7863 33977
rect 7863 33943 7897 33977
rect 7897 33943 7906 33977
rect 7854 33934 7906 33943
rect 8014 33977 8066 33986
rect 8014 33943 8023 33977
rect 8023 33943 8057 33977
rect 8057 33943 8066 33977
rect 8014 33934 8066 33943
rect 8174 33977 8226 33986
rect 8174 33943 8183 33977
rect 8183 33943 8217 33977
rect 8217 33943 8226 33977
rect 8174 33934 8226 33943
rect 8334 33977 8386 33986
rect 8334 33943 8343 33977
rect 8343 33943 8377 33977
rect 8377 33943 8386 33977
rect 8334 33934 8386 33943
rect 12494 33977 12546 33986
rect 12494 33943 12503 33977
rect 12503 33943 12537 33977
rect 12537 33943 12546 33977
rect 12494 33934 12546 33943
rect 12654 33977 12706 33986
rect 12654 33943 12663 33977
rect 12663 33943 12697 33977
rect 12697 33943 12706 33977
rect 12654 33934 12706 33943
rect 12814 33977 12866 33986
rect 12814 33943 12823 33977
rect 12823 33943 12857 33977
rect 12857 33943 12866 33977
rect 12814 33934 12866 33943
rect 12974 33977 13026 33986
rect 12974 33943 12983 33977
rect 12983 33943 13017 33977
rect 13017 33943 13026 33977
rect 12974 33934 13026 33943
rect 13134 33977 13186 33986
rect 13134 33943 13143 33977
rect 13143 33943 13177 33977
rect 13177 33943 13186 33977
rect 13134 33934 13186 33943
rect 13294 33977 13346 33986
rect 13294 33943 13303 33977
rect 13303 33943 13337 33977
rect 13337 33943 13346 33977
rect 13294 33934 13346 33943
rect 13454 33977 13506 33986
rect 13454 33943 13463 33977
rect 13463 33943 13497 33977
rect 13497 33943 13506 33977
rect 13454 33934 13506 33943
rect 13614 33977 13666 33986
rect 13614 33943 13623 33977
rect 13623 33943 13657 33977
rect 13657 33943 13666 33977
rect 13614 33934 13666 33943
rect 13774 33977 13826 33986
rect 13774 33943 13783 33977
rect 13783 33943 13817 33977
rect 13817 33943 13826 33977
rect 13774 33934 13826 33943
rect 13934 33977 13986 33986
rect 13934 33943 13943 33977
rect 13943 33943 13977 33977
rect 13977 33943 13986 33977
rect 13934 33934 13986 33943
rect 14094 33977 14146 33986
rect 14094 33943 14103 33977
rect 14103 33943 14137 33977
rect 14137 33943 14146 33977
rect 14094 33934 14146 33943
rect 14254 33977 14306 33986
rect 14254 33943 14263 33977
rect 14263 33943 14297 33977
rect 14297 33943 14306 33977
rect 14254 33934 14306 33943
rect 14414 33977 14466 33986
rect 14414 33943 14423 33977
rect 14423 33943 14457 33977
rect 14457 33943 14466 33977
rect 14414 33934 14466 33943
rect 14574 33977 14626 33986
rect 14574 33943 14583 33977
rect 14583 33943 14617 33977
rect 14617 33943 14626 33977
rect 14574 33934 14626 33943
rect 14734 33977 14786 33986
rect 14734 33943 14743 33977
rect 14743 33943 14777 33977
rect 14777 33943 14786 33977
rect 14734 33934 14786 33943
rect 14894 33977 14946 33986
rect 14894 33943 14903 33977
rect 14903 33943 14937 33977
rect 14937 33943 14946 33977
rect 14894 33934 14946 33943
rect 15054 33977 15106 33986
rect 15054 33943 15063 33977
rect 15063 33943 15097 33977
rect 15097 33943 15106 33977
rect 15054 33934 15106 33943
rect 15214 33977 15266 33986
rect 15214 33943 15223 33977
rect 15223 33943 15257 33977
rect 15257 33943 15266 33977
rect 15214 33934 15266 33943
rect 15374 33977 15426 33986
rect 15374 33943 15383 33977
rect 15383 33943 15417 33977
rect 15417 33943 15426 33977
rect 15374 33934 15426 33943
rect 15534 33977 15586 33986
rect 15534 33943 15543 33977
rect 15543 33943 15577 33977
rect 15577 33943 15586 33977
rect 15534 33934 15586 33943
rect 15694 33977 15746 33986
rect 15694 33943 15703 33977
rect 15703 33943 15737 33977
rect 15737 33943 15746 33977
rect 15694 33934 15746 33943
rect 15854 33977 15906 33986
rect 15854 33943 15863 33977
rect 15863 33943 15897 33977
rect 15897 33943 15906 33977
rect 15854 33934 15906 33943
rect 16014 33977 16066 33986
rect 16014 33943 16023 33977
rect 16023 33943 16057 33977
rect 16057 33943 16066 33977
rect 16014 33934 16066 33943
rect 16174 33977 16226 33986
rect 16174 33943 16183 33977
rect 16183 33943 16217 33977
rect 16217 33943 16226 33977
rect 16174 33934 16226 33943
rect 16334 33977 16386 33986
rect 16334 33943 16343 33977
rect 16343 33943 16377 33977
rect 16377 33943 16386 33977
rect 16334 33934 16386 33943
rect 16494 33977 16546 33986
rect 16494 33943 16503 33977
rect 16503 33943 16537 33977
rect 16537 33943 16546 33977
rect 16494 33934 16546 33943
rect 16654 33977 16706 33986
rect 16654 33943 16663 33977
rect 16663 33943 16697 33977
rect 16697 33943 16706 33977
rect 16654 33934 16706 33943
rect 16814 33977 16866 33986
rect 16814 33943 16823 33977
rect 16823 33943 16857 33977
rect 16857 33943 16866 33977
rect 16814 33934 16866 33943
rect 16974 33977 17026 33986
rect 16974 33943 16983 33977
rect 16983 33943 17017 33977
rect 17017 33943 17026 33977
rect 16974 33934 17026 33943
rect 17134 33977 17186 33986
rect 17134 33943 17143 33977
rect 17143 33943 17177 33977
rect 17177 33943 17186 33977
rect 17134 33934 17186 33943
rect 17294 33977 17346 33986
rect 17294 33943 17303 33977
rect 17303 33943 17337 33977
rect 17337 33943 17346 33977
rect 17294 33934 17346 33943
rect 17454 33977 17506 33986
rect 17454 33943 17463 33977
rect 17463 33943 17497 33977
rect 17497 33943 17506 33977
rect 17454 33934 17506 33943
rect 17614 33977 17666 33986
rect 17614 33943 17623 33977
rect 17623 33943 17657 33977
rect 17657 33943 17666 33977
rect 17614 33934 17666 33943
rect 17774 33977 17826 33986
rect 17774 33943 17783 33977
rect 17783 33943 17817 33977
rect 17817 33943 17826 33977
rect 17774 33934 17826 33943
rect 17934 33977 17986 33986
rect 17934 33943 17943 33977
rect 17943 33943 17977 33977
rect 17977 33943 17986 33977
rect 17934 33934 17986 33943
rect 18094 33977 18146 33986
rect 18094 33943 18103 33977
rect 18103 33943 18137 33977
rect 18137 33943 18146 33977
rect 18094 33934 18146 33943
rect 18254 33977 18306 33986
rect 18254 33943 18263 33977
rect 18263 33943 18297 33977
rect 18297 33943 18306 33977
rect 18254 33934 18306 33943
rect 18414 33977 18466 33986
rect 18414 33943 18423 33977
rect 18423 33943 18457 33977
rect 18457 33943 18466 33977
rect 18414 33934 18466 33943
rect 18574 33977 18626 33986
rect 18574 33943 18583 33977
rect 18583 33943 18617 33977
rect 18617 33943 18626 33977
rect 18574 33934 18626 33943
rect 18734 33977 18786 33986
rect 18734 33943 18743 33977
rect 18743 33943 18777 33977
rect 18777 33943 18786 33977
rect 18734 33934 18786 33943
rect 18894 33977 18946 33986
rect 18894 33943 18903 33977
rect 18903 33943 18937 33977
rect 18937 33943 18946 33977
rect 18894 33934 18946 33943
rect 23134 33977 23186 33986
rect 23134 33943 23143 33977
rect 23143 33943 23177 33977
rect 23177 33943 23186 33977
rect 23134 33934 23186 33943
rect 23294 33977 23346 33986
rect 23294 33943 23303 33977
rect 23303 33943 23337 33977
rect 23337 33943 23346 33977
rect 23294 33934 23346 33943
rect 23454 33977 23506 33986
rect 23454 33943 23463 33977
rect 23463 33943 23497 33977
rect 23497 33943 23506 33977
rect 23454 33934 23506 33943
rect 23614 33977 23666 33986
rect 23614 33943 23623 33977
rect 23623 33943 23657 33977
rect 23657 33943 23666 33977
rect 23614 33934 23666 33943
rect 23774 33977 23826 33986
rect 23774 33943 23783 33977
rect 23783 33943 23817 33977
rect 23817 33943 23826 33977
rect 23774 33934 23826 33943
rect 23934 33977 23986 33986
rect 23934 33943 23943 33977
rect 23943 33943 23977 33977
rect 23977 33943 23986 33977
rect 23934 33934 23986 33943
rect 24094 33977 24146 33986
rect 24094 33943 24103 33977
rect 24103 33943 24137 33977
rect 24137 33943 24146 33977
rect 24094 33934 24146 33943
rect 24254 33977 24306 33986
rect 24254 33943 24263 33977
rect 24263 33943 24297 33977
rect 24297 33943 24306 33977
rect 24254 33934 24306 33943
rect 24414 33977 24466 33986
rect 24414 33943 24423 33977
rect 24423 33943 24457 33977
rect 24457 33943 24466 33977
rect 24414 33934 24466 33943
rect 24574 33977 24626 33986
rect 24574 33943 24583 33977
rect 24583 33943 24617 33977
rect 24617 33943 24626 33977
rect 24574 33934 24626 33943
rect 24734 33977 24786 33986
rect 24734 33943 24743 33977
rect 24743 33943 24777 33977
rect 24777 33943 24786 33977
rect 24734 33934 24786 33943
rect 24894 33977 24946 33986
rect 24894 33943 24903 33977
rect 24903 33943 24937 33977
rect 24937 33943 24946 33977
rect 24894 33934 24946 33943
rect 25054 33977 25106 33986
rect 25054 33943 25063 33977
rect 25063 33943 25097 33977
rect 25097 33943 25106 33977
rect 25054 33934 25106 33943
rect 25214 33977 25266 33986
rect 25214 33943 25223 33977
rect 25223 33943 25257 33977
rect 25257 33943 25266 33977
rect 25214 33934 25266 33943
rect 25374 33977 25426 33986
rect 25374 33943 25383 33977
rect 25383 33943 25417 33977
rect 25417 33943 25426 33977
rect 25374 33934 25426 33943
rect 25534 33977 25586 33986
rect 25534 33943 25543 33977
rect 25543 33943 25577 33977
rect 25577 33943 25586 33977
rect 25534 33934 25586 33943
rect 25694 33977 25746 33986
rect 25694 33943 25703 33977
rect 25703 33943 25737 33977
rect 25737 33943 25746 33977
rect 25694 33934 25746 33943
rect 25854 33977 25906 33986
rect 25854 33943 25863 33977
rect 25863 33943 25897 33977
rect 25897 33943 25906 33977
rect 25854 33934 25906 33943
rect 26014 33977 26066 33986
rect 26014 33943 26023 33977
rect 26023 33943 26057 33977
rect 26057 33943 26066 33977
rect 26014 33934 26066 33943
rect 26174 33977 26226 33986
rect 26174 33943 26183 33977
rect 26183 33943 26217 33977
rect 26217 33943 26226 33977
rect 26174 33934 26226 33943
rect 26334 33977 26386 33986
rect 26334 33943 26343 33977
rect 26343 33943 26377 33977
rect 26377 33943 26386 33977
rect 26334 33934 26386 33943
rect 26494 33977 26546 33986
rect 26494 33943 26503 33977
rect 26503 33943 26537 33977
rect 26537 33943 26546 33977
rect 26494 33934 26546 33943
rect 26654 33977 26706 33986
rect 26654 33943 26663 33977
rect 26663 33943 26697 33977
rect 26697 33943 26706 33977
rect 26654 33934 26706 33943
rect 26814 33977 26866 33986
rect 26814 33943 26823 33977
rect 26823 33943 26857 33977
rect 26857 33943 26866 33977
rect 26814 33934 26866 33943
rect 26974 33977 27026 33986
rect 26974 33943 26983 33977
rect 26983 33943 27017 33977
rect 27017 33943 27026 33977
rect 26974 33934 27026 33943
rect 27134 33977 27186 33986
rect 27134 33943 27143 33977
rect 27143 33943 27177 33977
rect 27177 33943 27186 33977
rect 27134 33934 27186 33943
rect 27294 33977 27346 33986
rect 27294 33943 27303 33977
rect 27303 33943 27337 33977
rect 27337 33943 27346 33977
rect 27294 33934 27346 33943
rect 27454 33977 27506 33986
rect 27454 33943 27463 33977
rect 27463 33943 27497 33977
rect 27497 33943 27506 33977
rect 27454 33934 27506 33943
rect 27614 33977 27666 33986
rect 27614 33943 27623 33977
rect 27623 33943 27657 33977
rect 27657 33943 27666 33977
rect 27614 33934 27666 33943
rect 27774 33977 27826 33986
rect 27774 33943 27783 33977
rect 27783 33943 27817 33977
rect 27817 33943 27826 33977
rect 27774 33934 27826 33943
rect 27934 33977 27986 33986
rect 27934 33943 27943 33977
rect 27943 33943 27977 33977
rect 27977 33943 27986 33977
rect 27934 33934 27986 33943
rect 28094 33977 28146 33986
rect 28094 33943 28103 33977
rect 28103 33943 28137 33977
rect 28137 33943 28146 33977
rect 28094 33934 28146 33943
rect 28254 33977 28306 33986
rect 28254 33943 28263 33977
rect 28263 33943 28297 33977
rect 28297 33943 28306 33977
rect 28254 33934 28306 33943
rect 28414 33977 28466 33986
rect 28414 33943 28423 33977
rect 28423 33943 28457 33977
rect 28457 33943 28466 33977
rect 28414 33934 28466 33943
rect 28574 33977 28626 33986
rect 28574 33943 28583 33977
rect 28583 33943 28617 33977
rect 28617 33943 28626 33977
rect 28574 33934 28626 33943
rect 28734 33977 28786 33986
rect 28734 33943 28743 33977
rect 28743 33943 28777 33977
rect 28777 33943 28786 33977
rect 28734 33934 28786 33943
rect 28894 33977 28946 33986
rect 28894 33943 28903 33977
rect 28903 33943 28937 33977
rect 28937 33943 28946 33977
rect 28894 33934 28946 33943
rect 29054 33977 29106 33986
rect 29054 33943 29063 33977
rect 29063 33943 29097 33977
rect 29097 33943 29106 33977
rect 29054 33934 29106 33943
rect 29214 33977 29266 33986
rect 29214 33943 29223 33977
rect 29223 33943 29257 33977
rect 29257 33943 29266 33977
rect 29214 33934 29266 33943
rect 29374 33977 29426 33986
rect 29374 33943 29383 33977
rect 29383 33943 29417 33977
rect 29417 33943 29426 33977
rect 29374 33934 29426 33943
rect 33534 33977 33586 33986
rect 33534 33943 33543 33977
rect 33543 33943 33577 33977
rect 33577 33943 33586 33977
rect 33534 33934 33586 33943
rect 33694 33977 33746 33986
rect 33694 33943 33703 33977
rect 33703 33943 33737 33977
rect 33737 33943 33746 33977
rect 33694 33934 33746 33943
rect 33854 33977 33906 33986
rect 33854 33943 33863 33977
rect 33863 33943 33897 33977
rect 33897 33943 33906 33977
rect 33854 33934 33906 33943
rect 34014 33977 34066 33986
rect 34014 33943 34023 33977
rect 34023 33943 34057 33977
rect 34057 33943 34066 33977
rect 34014 33934 34066 33943
rect 34174 33977 34226 33986
rect 34174 33943 34183 33977
rect 34183 33943 34217 33977
rect 34217 33943 34226 33977
rect 34174 33934 34226 33943
rect 34334 33977 34386 33986
rect 34334 33943 34343 33977
rect 34343 33943 34377 33977
rect 34377 33943 34386 33977
rect 34334 33934 34386 33943
rect 34494 33977 34546 33986
rect 34494 33943 34503 33977
rect 34503 33943 34537 33977
rect 34537 33943 34546 33977
rect 34494 33934 34546 33943
rect 34654 33977 34706 33986
rect 34654 33943 34663 33977
rect 34663 33943 34697 33977
rect 34697 33943 34706 33977
rect 34654 33934 34706 33943
rect 34814 33977 34866 33986
rect 34814 33943 34823 33977
rect 34823 33943 34857 33977
rect 34857 33943 34866 33977
rect 34814 33934 34866 33943
rect 34974 33977 35026 33986
rect 34974 33943 34983 33977
rect 34983 33943 35017 33977
rect 35017 33943 35026 33977
rect 34974 33934 35026 33943
rect 35134 33977 35186 33986
rect 35134 33943 35143 33977
rect 35143 33943 35177 33977
rect 35177 33943 35186 33977
rect 35134 33934 35186 33943
rect 35294 33977 35346 33986
rect 35294 33943 35303 33977
rect 35303 33943 35337 33977
rect 35337 33943 35346 33977
rect 35294 33934 35346 33943
rect 35454 33977 35506 33986
rect 35454 33943 35463 33977
rect 35463 33943 35497 33977
rect 35497 33943 35506 33977
rect 35454 33934 35506 33943
rect 35614 33977 35666 33986
rect 35614 33943 35623 33977
rect 35623 33943 35657 33977
rect 35657 33943 35666 33977
rect 35614 33934 35666 33943
rect 35774 33977 35826 33986
rect 35774 33943 35783 33977
rect 35783 33943 35817 33977
rect 35817 33943 35826 33977
rect 35774 33934 35826 33943
rect 35934 33977 35986 33986
rect 35934 33943 35943 33977
rect 35943 33943 35977 33977
rect 35977 33943 35986 33977
rect 35934 33934 35986 33943
rect 36094 33977 36146 33986
rect 36094 33943 36103 33977
rect 36103 33943 36137 33977
rect 36137 33943 36146 33977
rect 36094 33934 36146 33943
rect 36254 33977 36306 33986
rect 36254 33943 36263 33977
rect 36263 33943 36297 33977
rect 36297 33943 36306 33977
rect 36254 33934 36306 33943
rect 36414 33977 36466 33986
rect 36414 33943 36423 33977
rect 36423 33943 36457 33977
rect 36457 33943 36466 33977
rect 36414 33934 36466 33943
rect 36574 33977 36626 33986
rect 36574 33943 36583 33977
rect 36583 33943 36617 33977
rect 36617 33943 36626 33977
rect 36574 33934 36626 33943
rect 36734 33977 36786 33986
rect 36734 33943 36743 33977
rect 36743 33943 36777 33977
rect 36777 33943 36786 33977
rect 36734 33934 36786 33943
rect 36894 33977 36946 33986
rect 36894 33943 36903 33977
rect 36903 33943 36937 33977
rect 36937 33943 36946 33977
rect 36894 33934 36946 33943
rect 37054 33977 37106 33986
rect 37054 33943 37063 33977
rect 37063 33943 37097 33977
rect 37097 33943 37106 33977
rect 37054 33934 37106 33943
rect 37214 33977 37266 33986
rect 37214 33943 37223 33977
rect 37223 33943 37257 33977
rect 37257 33943 37266 33977
rect 37214 33934 37266 33943
rect 37374 33977 37426 33986
rect 37374 33943 37383 33977
rect 37383 33943 37417 33977
rect 37417 33943 37426 33977
rect 37374 33934 37426 33943
rect 37534 33977 37586 33986
rect 37534 33943 37543 33977
rect 37543 33943 37577 33977
rect 37577 33943 37586 33977
rect 37534 33934 37586 33943
rect 37694 33977 37746 33986
rect 37694 33943 37703 33977
rect 37703 33943 37737 33977
rect 37737 33943 37746 33977
rect 37694 33934 37746 33943
rect 37854 33977 37906 33986
rect 37854 33943 37863 33977
rect 37863 33943 37897 33977
rect 37897 33943 37906 33977
rect 37854 33934 37906 33943
rect 38014 33977 38066 33986
rect 38014 33943 38023 33977
rect 38023 33943 38057 33977
rect 38057 33943 38066 33977
rect 38014 33934 38066 33943
rect 38174 33977 38226 33986
rect 38174 33943 38183 33977
rect 38183 33943 38217 33977
rect 38217 33943 38226 33977
rect 38174 33934 38226 33943
rect 38334 33977 38386 33986
rect 38334 33943 38343 33977
rect 38343 33943 38377 33977
rect 38377 33943 38386 33977
rect 38334 33934 38386 33943
rect 38494 33977 38546 33986
rect 38494 33943 38503 33977
rect 38503 33943 38537 33977
rect 38537 33943 38546 33977
rect 38494 33934 38546 33943
rect 38654 33977 38706 33986
rect 38654 33943 38663 33977
rect 38663 33943 38697 33977
rect 38697 33943 38706 33977
rect 38654 33934 38706 33943
rect 38814 33977 38866 33986
rect 38814 33943 38823 33977
rect 38823 33943 38857 33977
rect 38857 33943 38866 33977
rect 38814 33934 38866 33943
rect 38974 33977 39026 33986
rect 38974 33943 38983 33977
rect 38983 33943 39017 33977
rect 39017 33943 39026 33977
rect 38974 33934 39026 33943
rect 39134 33977 39186 33986
rect 39134 33943 39143 33977
rect 39143 33943 39177 33977
rect 39177 33943 39186 33977
rect 39134 33934 39186 33943
rect 39294 33977 39346 33986
rect 39294 33943 39303 33977
rect 39303 33943 39337 33977
rect 39337 33943 39346 33977
rect 39294 33934 39346 33943
rect 39454 33977 39506 33986
rect 39454 33943 39463 33977
rect 39463 33943 39497 33977
rect 39497 33943 39506 33977
rect 39454 33934 39506 33943
rect 39614 33977 39666 33986
rect 39614 33943 39623 33977
rect 39623 33943 39657 33977
rect 39657 33943 39666 33977
rect 39614 33934 39666 33943
rect 39774 33977 39826 33986
rect 39774 33943 39783 33977
rect 39783 33943 39817 33977
rect 39817 33943 39826 33977
rect 39774 33934 39826 33943
rect 39934 33977 39986 33986
rect 39934 33943 39943 33977
rect 39943 33943 39977 33977
rect 39977 33943 39986 33977
rect 39934 33934 39986 33943
rect 40094 33977 40146 33986
rect 40094 33943 40103 33977
rect 40103 33943 40137 33977
rect 40137 33943 40146 33977
rect 40094 33934 40146 33943
rect 40254 33977 40306 33986
rect 40254 33943 40263 33977
rect 40263 33943 40297 33977
rect 40297 33943 40306 33977
rect 40254 33934 40306 33943
rect 40414 33977 40466 33986
rect 40414 33943 40423 33977
rect 40423 33943 40457 33977
rect 40457 33943 40466 33977
rect 40414 33934 40466 33943
rect 40574 33977 40626 33986
rect 40574 33943 40583 33977
rect 40583 33943 40617 33977
rect 40617 33943 40626 33977
rect 40574 33934 40626 33943
rect 40734 33977 40786 33986
rect 40734 33943 40743 33977
rect 40743 33943 40777 33977
rect 40777 33943 40786 33977
rect 40734 33934 40786 33943
rect 40894 33977 40946 33986
rect 40894 33943 40903 33977
rect 40903 33943 40937 33977
rect 40937 33943 40946 33977
rect 40894 33934 40946 33943
rect 41054 33977 41106 33986
rect 41054 33943 41063 33977
rect 41063 33943 41097 33977
rect 41097 33943 41106 33977
rect 41054 33934 41106 33943
rect 41214 33977 41266 33986
rect 41214 33943 41223 33977
rect 41223 33943 41257 33977
rect 41257 33943 41266 33977
rect 41214 33934 41266 33943
rect 41374 33977 41426 33986
rect 41374 33943 41383 33977
rect 41383 33943 41417 33977
rect 41417 33943 41426 33977
rect 41374 33934 41426 33943
rect 41534 33977 41586 33986
rect 41534 33943 41543 33977
rect 41543 33943 41577 33977
rect 41577 33943 41586 33977
rect 41534 33934 41586 33943
rect 41694 33977 41746 33986
rect 41694 33943 41703 33977
rect 41703 33943 41737 33977
rect 41737 33943 41746 33977
rect 41694 33934 41746 33943
rect 41854 33977 41906 33986
rect 41854 33943 41863 33977
rect 41863 33943 41897 33977
rect 41897 33943 41906 33977
rect 41854 33934 41906 33943
rect 14 33817 66 33826
rect 14 33783 23 33817
rect 23 33783 57 33817
rect 57 33783 66 33817
rect 14 33774 66 33783
rect 174 33817 226 33826
rect 174 33783 183 33817
rect 183 33783 217 33817
rect 217 33783 226 33817
rect 174 33774 226 33783
rect 334 33817 386 33826
rect 334 33783 343 33817
rect 343 33783 377 33817
rect 377 33783 386 33817
rect 334 33774 386 33783
rect 494 33817 546 33826
rect 494 33783 503 33817
rect 503 33783 537 33817
rect 537 33783 546 33817
rect 494 33774 546 33783
rect 654 33817 706 33826
rect 654 33783 663 33817
rect 663 33783 697 33817
rect 697 33783 706 33817
rect 654 33774 706 33783
rect 814 33817 866 33826
rect 814 33783 823 33817
rect 823 33783 857 33817
rect 857 33783 866 33817
rect 814 33774 866 33783
rect 974 33817 1026 33826
rect 974 33783 983 33817
rect 983 33783 1017 33817
rect 1017 33783 1026 33817
rect 974 33774 1026 33783
rect 1134 33817 1186 33826
rect 1134 33783 1143 33817
rect 1143 33783 1177 33817
rect 1177 33783 1186 33817
rect 1134 33774 1186 33783
rect 1294 33817 1346 33826
rect 1294 33783 1303 33817
rect 1303 33783 1337 33817
rect 1337 33783 1346 33817
rect 1294 33774 1346 33783
rect 1454 33817 1506 33826
rect 1454 33783 1463 33817
rect 1463 33783 1497 33817
rect 1497 33783 1506 33817
rect 1454 33774 1506 33783
rect 1614 33817 1666 33826
rect 1614 33783 1623 33817
rect 1623 33783 1657 33817
rect 1657 33783 1666 33817
rect 1614 33774 1666 33783
rect 1774 33817 1826 33826
rect 1774 33783 1783 33817
rect 1783 33783 1817 33817
rect 1817 33783 1826 33817
rect 1774 33774 1826 33783
rect 1934 33817 1986 33826
rect 1934 33783 1943 33817
rect 1943 33783 1977 33817
rect 1977 33783 1986 33817
rect 1934 33774 1986 33783
rect 2094 33817 2146 33826
rect 2094 33783 2103 33817
rect 2103 33783 2137 33817
rect 2137 33783 2146 33817
rect 2094 33774 2146 33783
rect 2254 33817 2306 33826
rect 2254 33783 2263 33817
rect 2263 33783 2297 33817
rect 2297 33783 2306 33817
rect 2254 33774 2306 33783
rect 2414 33817 2466 33826
rect 2414 33783 2423 33817
rect 2423 33783 2457 33817
rect 2457 33783 2466 33817
rect 2414 33774 2466 33783
rect 2574 33817 2626 33826
rect 2574 33783 2583 33817
rect 2583 33783 2617 33817
rect 2617 33783 2626 33817
rect 2574 33774 2626 33783
rect 2734 33817 2786 33826
rect 2734 33783 2743 33817
rect 2743 33783 2777 33817
rect 2777 33783 2786 33817
rect 2734 33774 2786 33783
rect 2894 33817 2946 33826
rect 2894 33783 2903 33817
rect 2903 33783 2937 33817
rect 2937 33783 2946 33817
rect 2894 33774 2946 33783
rect 3054 33817 3106 33826
rect 3054 33783 3063 33817
rect 3063 33783 3097 33817
rect 3097 33783 3106 33817
rect 3054 33774 3106 33783
rect 3214 33817 3266 33826
rect 3214 33783 3223 33817
rect 3223 33783 3257 33817
rect 3257 33783 3266 33817
rect 3214 33774 3266 33783
rect 3374 33817 3426 33826
rect 3374 33783 3383 33817
rect 3383 33783 3417 33817
rect 3417 33783 3426 33817
rect 3374 33774 3426 33783
rect 3534 33817 3586 33826
rect 3534 33783 3543 33817
rect 3543 33783 3577 33817
rect 3577 33783 3586 33817
rect 3534 33774 3586 33783
rect 3694 33817 3746 33826
rect 3694 33783 3703 33817
rect 3703 33783 3737 33817
rect 3737 33783 3746 33817
rect 3694 33774 3746 33783
rect 3854 33817 3906 33826
rect 3854 33783 3863 33817
rect 3863 33783 3897 33817
rect 3897 33783 3906 33817
rect 3854 33774 3906 33783
rect 4014 33817 4066 33826
rect 4014 33783 4023 33817
rect 4023 33783 4057 33817
rect 4057 33783 4066 33817
rect 4014 33774 4066 33783
rect 4174 33817 4226 33826
rect 4174 33783 4183 33817
rect 4183 33783 4217 33817
rect 4217 33783 4226 33817
rect 4174 33774 4226 33783
rect 4334 33817 4386 33826
rect 4334 33783 4343 33817
rect 4343 33783 4377 33817
rect 4377 33783 4386 33817
rect 4334 33774 4386 33783
rect 4494 33817 4546 33826
rect 4494 33783 4503 33817
rect 4503 33783 4537 33817
rect 4537 33783 4546 33817
rect 4494 33774 4546 33783
rect 4654 33817 4706 33826
rect 4654 33783 4663 33817
rect 4663 33783 4697 33817
rect 4697 33783 4706 33817
rect 4654 33774 4706 33783
rect 4814 33817 4866 33826
rect 4814 33783 4823 33817
rect 4823 33783 4857 33817
rect 4857 33783 4866 33817
rect 4814 33774 4866 33783
rect 4974 33817 5026 33826
rect 4974 33783 4983 33817
rect 4983 33783 5017 33817
rect 5017 33783 5026 33817
rect 4974 33774 5026 33783
rect 5134 33817 5186 33826
rect 5134 33783 5143 33817
rect 5143 33783 5177 33817
rect 5177 33783 5186 33817
rect 5134 33774 5186 33783
rect 5294 33817 5346 33826
rect 5294 33783 5303 33817
rect 5303 33783 5337 33817
rect 5337 33783 5346 33817
rect 5294 33774 5346 33783
rect 5454 33817 5506 33826
rect 5454 33783 5463 33817
rect 5463 33783 5497 33817
rect 5497 33783 5506 33817
rect 5454 33774 5506 33783
rect 5614 33817 5666 33826
rect 5614 33783 5623 33817
rect 5623 33783 5657 33817
rect 5657 33783 5666 33817
rect 5614 33774 5666 33783
rect 5774 33817 5826 33826
rect 5774 33783 5783 33817
rect 5783 33783 5817 33817
rect 5817 33783 5826 33817
rect 5774 33774 5826 33783
rect 5934 33817 5986 33826
rect 5934 33783 5943 33817
rect 5943 33783 5977 33817
rect 5977 33783 5986 33817
rect 5934 33774 5986 33783
rect 6094 33817 6146 33826
rect 6094 33783 6103 33817
rect 6103 33783 6137 33817
rect 6137 33783 6146 33817
rect 6094 33774 6146 33783
rect 6254 33817 6306 33826
rect 6254 33783 6263 33817
rect 6263 33783 6297 33817
rect 6297 33783 6306 33817
rect 6254 33774 6306 33783
rect 6414 33817 6466 33826
rect 6414 33783 6423 33817
rect 6423 33783 6457 33817
rect 6457 33783 6466 33817
rect 6414 33774 6466 33783
rect 6574 33817 6626 33826
rect 6574 33783 6583 33817
rect 6583 33783 6617 33817
rect 6617 33783 6626 33817
rect 6574 33774 6626 33783
rect 6734 33817 6786 33826
rect 6734 33783 6743 33817
rect 6743 33783 6777 33817
rect 6777 33783 6786 33817
rect 6734 33774 6786 33783
rect 6894 33817 6946 33826
rect 6894 33783 6903 33817
rect 6903 33783 6937 33817
rect 6937 33783 6946 33817
rect 6894 33774 6946 33783
rect 7054 33817 7106 33826
rect 7054 33783 7063 33817
rect 7063 33783 7097 33817
rect 7097 33783 7106 33817
rect 7054 33774 7106 33783
rect 7214 33817 7266 33826
rect 7214 33783 7223 33817
rect 7223 33783 7257 33817
rect 7257 33783 7266 33817
rect 7214 33774 7266 33783
rect 7374 33817 7426 33826
rect 7374 33783 7383 33817
rect 7383 33783 7417 33817
rect 7417 33783 7426 33817
rect 7374 33774 7426 33783
rect 7534 33817 7586 33826
rect 7534 33783 7543 33817
rect 7543 33783 7577 33817
rect 7577 33783 7586 33817
rect 7534 33774 7586 33783
rect 7694 33817 7746 33826
rect 7694 33783 7703 33817
rect 7703 33783 7737 33817
rect 7737 33783 7746 33817
rect 7694 33774 7746 33783
rect 7854 33817 7906 33826
rect 7854 33783 7863 33817
rect 7863 33783 7897 33817
rect 7897 33783 7906 33817
rect 7854 33774 7906 33783
rect 8014 33817 8066 33826
rect 8014 33783 8023 33817
rect 8023 33783 8057 33817
rect 8057 33783 8066 33817
rect 8014 33774 8066 33783
rect 8174 33817 8226 33826
rect 8174 33783 8183 33817
rect 8183 33783 8217 33817
rect 8217 33783 8226 33817
rect 8174 33774 8226 33783
rect 8334 33817 8386 33826
rect 8334 33783 8343 33817
rect 8343 33783 8377 33817
rect 8377 33783 8386 33817
rect 8334 33774 8386 33783
rect 12494 33817 12546 33826
rect 12494 33783 12503 33817
rect 12503 33783 12537 33817
rect 12537 33783 12546 33817
rect 12494 33774 12546 33783
rect 12654 33817 12706 33826
rect 12654 33783 12663 33817
rect 12663 33783 12697 33817
rect 12697 33783 12706 33817
rect 12654 33774 12706 33783
rect 12814 33817 12866 33826
rect 12814 33783 12823 33817
rect 12823 33783 12857 33817
rect 12857 33783 12866 33817
rect 12814 33774 12866 33783
rect 12974 33817 13026 33826
rect 12974 33783 12983 33817
rect 12983 33783 13017 33817
rect 13017 33783 13026 33817
rect 12974 33774 13026 33783
rect 13134 33817 13186 33826
rect 13134 33783 13143 33817
rect 13143 33783 13177 33817
rect 13177 33783 13186 33817
rect 13134 33774 13186 33783
rect 13294 33817 13346 33826
rect 13294 33783 13303 33817
rect 13303 33783 13337 33817
rect 13337 33783 13346 33817
rect 13294 33774 13346 33783
rect 13454 33817 13506 33826
rect 13454 33783 13463 33817
rect 13463 33783 13497 33817
rect 13497 33783 13506 33817
rect 13454 33774 13506 33783
rect 13614 33817 13666 33826
rect 13614 33783 13623 33817
rect 13623 33783 13657 33817
rect 13657 33783 13666 33817
rect 13614 33774 13666 33783
rect 13774 33817 13826 33826
rect 13774 33783 13783 33817
rect 13783 33783 13817 33817
rect 13817 33783 13826 33817
rect 13774 33774 13826 33783
rect 13934 33817 13986 33826
rect 13934 33783 13943 33817
rect 13943 33783 13977 33817
rect 13977 33783 13986 33817
rect 13934 33774 13986 33783
rect 14094 33817 14146 33826
rect 14094 33783 14103 33817
rect 14103 33783 14137 33817
rect 14137 33783 14146 33817
rect 14094 33774 14146 33783
rect 14254 33817 14306 33826
rect 14254 33783 14263 33817
rect 14263 33783 14297 33817
rect 14297 33783 14306 33817
rect 14254 33774 14306 33783
rect 14414 33817 14466 33826
rect 14414 33783 14423 33817
rect 14423 33783 14457 33817
rect 14457 33783 14466 33817
rect 14414 33774 14466 33783
rect 14574 33817 14626 33826
rect 14574 33783 14583 33817
rect 14583 33783 14617 33817
rect 14617 33783 14626 33817
rect 14574 33774 14626 33783
rect 14734 33817 14786 33826
rect 14734 33783 14743 33817
rect 14743 33783 14777 33817
rect 14777 33783 14786 33817
rect 14734 33774 14786 33783
rect 14894 33817 14946 33826
rect 14894 33783 14903 33817
rect 14903 33783 14937 33817
rect 14937 33783 14946 33817
rect 14894 33774 14946 33783
rect 15054 33817 15106 33826
rect 15054 33783 15063 33817
rect 15063 33783 15097 33817
rect 15097 33783 15106 33817
rect 15054 33774 15106 33783
rect 15214 33817 15266 33826
rect 15214 33783 15223 33817
rect 15223 33783 15257 33817
rect 15257 33783 15266 33817
rect 15214 33774 15266 33783
rect 15374 33817 15426 33826
rect 15374 33783 15383 33817
rect 15383 33783 15417 33817
rect 15417 33783 15426 33817
rect 15374 33774 15426 33783
rect 15534 33817 15586 33826
rect 15534 33783 15543 33817
rect 15543 33783 15577 33817
rect 15577 33783 15586 33817
rect 15534 33774 15586 33783
rect 15694 33817 15746 33826
rect 15694 33783 15703 33817
rect 15703 33783 15737 33817
rect 15737 33783 15746 33817
rect 15694 33774 15746 33783
rect 15854 33817 15906 33826
rect 15854 33783 15863 33817
rect 15863 33783 15897 33817
rect 15897 33783 15906 33817
rect 15854 33774 15906 33783
rect 16014 33817 16066 33826
rect 16014 33783 16023 33817
rect 16023 33783 16057 33817
rect 16057 33783 16066 33817
rect 16014 33774 16066 33783
rect 16174 33817 16226 33826
rect 16174 33783 16183 33817
rect 16183 33783 16217 33817
rect 16217 33783 16226 33817
rect 16174 33774 16226 33783
rect 16334 33817 16386 33826
rect 16334 33783 16343 33817
rect 16343 33783 16377 33817
rect 16377 33783 16386 33817
rect 16334 33774 16386 33783
rect 16494 33817 16546 33826
rect 16494 33783 16503 33817
rect 16503 33783 16537 33817
rect 16537 33783 16546 33817
rect 16494 33774 16546 33783
rect 16654 33817 16706 33826
rect 16654 33783 16663 33817
rect 16663 33783 16697 33817
rect 16697 33783 16706 33817
rect 16654 33774 16706 33783
rect 16814 33817 16866 33826
rect 16814 33783 16823 33817
rect 16823 33783 16857 33817
rect 16857 33783 16866 33817
rect 16814 33774 16866 33783
rect 16974 33817 17026 33826
rect 16974 33783 16983 33817
rect 16983 33783 17017 33817
rect 17017 33783 17026 33817
rect 16974 33774 17026 33783
rect 17134 33817 17186 33826
rect 17134 33783 17143 33817
rect 17143 33783 17177 33817
rect 17177 33783 17186 33817
rect 17134 33774 17186 33783
rect 17294 33817 17346 33826
rect 17294 33783 17303 33817
rect 17303 33783 17337 33817
rect 17337 33783 17346 33817
rect 17294 33774 17346 33783
rect 17454 33817 17506 33826
rect 17454 33783 17463 33817
rect 17463 33783 17497 33817
rect 17497 33783 17506 33817
rect 17454 33774 17506 33783
rect 17614 33817 17666 33826
rect 17614 33783 17623 33817
rect 17623 33783 17657 33817
rect 17657 33783 17666 33817
rect 17614 33774 17666 33783
rect 17774 33817 17826 33826
rect 17774 33783 17783 33817
rect 17783 33783 17817 33817
rect 17817 33783 17826 33817
rect 17774 33774 17826 33783
rect 17934 33817 17986 33826
rect 17934 33783 17943 33817
rect 17943 33783 17977 33817
rect 17977 33783 17986 33817
rect 17934 33774 17986 33783
rect 18094 33817 18146 33826
rect 18094 33783 18103 33817
rect 18103 33783 18137 33817
rect 18137 33783 18146 33817
rect 18094 33774 18146 33783
rect 18254 33817 18306 33826
rect 18254 33783 18263 33817
rect 18263 33783 18297 33817
rect 18297 33783 18306 33817
rect 18254 33774 18306 33783
rect 18414 33817 18466 33826
rect 18414 33783 18423 33817
rect 18423 33783 18457 33817
rect 18457 33783 18466 33817
rect 18414 33774 18466 33783
rect 18574 33817 18626 33826
rect 18574 33783 18583 33817
rect 18583 33783 18617 33817
rect 18617 33783 18626 33817
rect 18574 33774 18626 33783
rect 18734 33817 18786 33826
rect 18734 33783 18743 33817
rect 18743 33783 18777 33817
rect 18777 33783 18786 33817
rect 18734 33774 18786 33783
rect 18894 33817 18946 33826
rect 18894 33783 18903 33817
rect 18903 33783 18937 33817
rect 18937 33783 18946 33817
rect 18894 33774 18946 33783
rect 23134 33817 23186 33826
rect 23134 33783 23143 33817
rect 23143 33783 23177 33817
rect 23177 33783 23186 33817
rect 23134 33774 23186 33783
rect 23294 33817 23346 33826
rect 23294 33783 23303 33817
rect 23303 33783 23337 33817
rect 23337 33783 23346 33817
rect 23294 33774 23346 33783
rect 23454 33817 23506 33826
rect 23454 33783 23463 33817
rect 23463 33783 23497 33817
rect 23497 33783 23506 33817
rect 23454 33774 23506 33783
rect 23614 33817 23666 33826
rect 23614 33783 23623 33817
rect 23623 33783 23657 33817
rect 23657 33783 23666 33817
rect 23614 33774 23666 33783
rect 23774 33817 23826 33826
rect 23774 33783 23783 33817
rect 23783 33783 23817 33817
rect 23817 33783 23826 33817
rect 23774 33774 23826 33783
rect 23934 33817 23986 33826
rect 23934 33783 23943 33817
rect 23943 33783 23977 33817
rect 23977 33783 23986 33817
rect 23934 33774 23986 33783
rect 24094 33817 24146 33826
rect 24094 33783 24103 33817
rect 24103 33783 24137 33817
rect 24137 33783 24146 33817
rect 24094 33774 24146 33783
rect 24254 33817 24306 33826
rect 24254 33783 24263 33817
rect 24263 33783 24297 33817
rect 24297 33783 24306 33817
rect 24254 33774 24306 33783
rect 24414 33817 24466 33826
rect 24414 33783 24423 33817
rect 24423 33783 24457 33817
rect 24457 33783 24466 33817
rect 24414 33774 24466 33783
rect 24574 33817 24626 33826
rect 24574 33783 24583 33817
rect 24583 33783 24617 33817
rect 24617 33783 24626 33817
rect 24574 33774 24626 33783
rect 24734 33817 24786 33826
rect 24734 33783 24743 33817
rect 24743 33783 24777 33817
rect 24777 33783 24786 33817
rect 24734 33774 24786 33783
rect 24894 33817 24946 33826
rect 24894 33783 24903 33817
rect 24903 33783 24937 33817
rect 24937 33783 24946 33817
rect 24894 33774 24946 33783
rect 25054 33817 25106 33826
rect 25054 33783 25063 33817
rect 25063 33783 25097 33817
rect 25097 33783 25106 33817
rect 25054 33774 25106 33783
rect 25214 33817 25266 33826
rect 25214 33783 25223 33817
rect 25223 33783 25257 33817
rect 25257 33783 25266 33817
rect 25214 33774 25266 33783
rect 25374 33817 25426 33826
rect 25374 33783 25383 33817
rect 25383 33783 25417 33817
rect 25417 33783 25426 33817
rect 25374 33774 25426 33783
rect 25534 33817 25586 33826
rect 25534 33783 25543 33817
rect 25543 33783 25577 33817
rect 25577 33783 25586 33817
rect 25534 33774 25586 33783
rect 25694 33817 25746 33826
rect 25694 33783 25703 33817
rect 25703 33783 25737 33817
rect 25737 33783 25746 33817
rect 25694 33774 25746 33783
rect 25854 33817 25906 33826
rect 25854 33783 25863 33817
rect 25863 33783 25897 33817
rect 25897 33783 25906 33817
rect 25854 33774 25906 33783
rect 26014 33817 26066 33826
rect 26014 33783 26023 33817
rect 26023 33783 26057 33817
rect 26057 33783 26066 33817
rect 26014 33774 26066 33783
rect 26174 33817 26226 33826
rect 26174 33783 26183 33817
rect 26183 33783 26217 33817
rect 26217 33783 26226 33817
rect 26174 33774 26226 33783
rect 26334 33817 26386 33826
rect 26334 33783 26343 33817
rect 26343 33783 26377 33817
rect 26377 33783 26386 33817
rect 26334 33774 26386 33783
rect 26494 33817 26546 33826
rect 26494 33783 26503 33817
rect 26503 33783 26537 33817
rect 26537 33783 26546 33817
rect 26494 33774 26546 33783
rect 26654 33817 26706 33826
rect 26654 33783 26663 33817
rect 26663 33783 26697 33817
rect 26697 33783 26706 33817
rect 26654 33774 26706 33783
rect 26814 33817 26866 33826
rect 26814 33783 26823 33817
rect 26823 33783 26857 33817
rect 26857 33783 26866 33817
rect 26814 33774 26866 33783
rect 26974 33817 27026 33826
rect 26974 33783 26983 33817
rect 26983 33783 27017 33817
rect 27017 33783 27026 33817
rect 26974 33774 27026 33783
rect 27134 33817 27186 33826
rect 27134 33783 27143 33817
rect 27143 33783 27177 33817
rect 27177 33783 27186 33817
rect 27134 33774 27186 33783
rect 27294 33817 27346 33826
rect 27294 33783 27303 33817
rect 27303 33783 27337 33817
rect 27337 33783 27346 33817
rect 27294 33774 27346 33783
rect 27454 33817 27506 33826
rect 27454 33783 27463 33817
rect 27463 33783 27497 33817
rect 27497 33783 27506 33817
rect 27454 33774 27506 33783
rect 27614 33817 27666 33826
rect 27614 33783 27623 33817
rect 27623 33783 27657 33817
rect 27657 33783 27666 33817
rect 27614 33774 27666 33783
rect 27774 33817 27826 33826
rect 27774 33783 27783 33817
rect 27783 33783 27817 33817
rect 27817 33783 27826 33817
rect 27774 33774 27826 33783
rect 27934 33817 27986 33826
rect 27934 33783 27943 33817
rect 27943 33783 27977 33817
rect 27977 33783 27986 33817
rect 27934 33774 27986 33783
rect 28094 33817 28146 33826
rect 28094 33783 28103 33817
rect 28103 33783 28137 33817
rect 28137 33783 28146 33817
rect 28094 33774 28146 33783
rect 28254 33817 28306 33826
rect 28254 33783 28263 33817
rect 28263 33783 28297 33817
rect 28297 33783 28306 33817
rect 28254 33774 28306 33783
rect 28414 33817 28466 33826
rect 28414 33783 28423 33817
rect 28423 33783 28457 33817
rect 28457 33783 28466 33817
rect 28414 33774 28466 33783
rect 28574 33817 28626 33826
rect 28574 33783 28583 33817
rect 28583 33783 28617 33817
rect 28617 33783 28626 33817
rect 28574 33774 28626 33783
rect 28734 33817 28786 33826
rect 28734 33783 28743 33817
rect 28743 33783 28777 33817
rect 28777 33783 28786 33817
rect 28734 33774 28786 33783
rect 28894 33817 28946 33826
rect 28894 33783 28903 33817
rect 28903 33783 28937 33817
rect 28937 33783 28946 33817
rect 28894 33774 28946 33783
rect 29054 33817 29106 33826
rect 29054 33783 29063 33817
rect 29063 33783 29097 33817
rect 29097 33783 29106 33817
rect 29054 33774 29106 33783
rect 29214 33817 29266 33826
rect 29214 33783 29223 33817
rect 29223 33783 29257 33817
rect 29257 33783 29266 33817
rect 29214 33774 29266 33783
rect 29374 33817 29426 33826
rect 29374 33783 29383 33817
rect 29383 33783 29417 33817
rect 29417 33783 29426 33817
rect 29374 33774 29426 33783
rect 33534 33817 33586 33826
rect 33534 33783 33543 33817
rect 33543 33783 33577 33817
rect 33577 33783 33586 33817
rect 33534 33774 33586 33783
rect 33694 33817 33746 33826
rect 33694 33783 33703 33817
rect 33703 33783 33737 33817
rect 33737 33783 33746 33817
rect 33694 33774 33746 33783
rect 33854 33817 33906 33826
rect 33854 33783 33863 33817
rect 33863 33783 33897 33817
rect 33897 33783 33906 33817
rect 33854 33774 33906 33783
rect 34014 33817 34066 33826
rect 34014 33783 34023 33817
rect 34023 33783 34057 33817
rect 34057 33783 34066 33817
rect 34014 33774 34066 33783
rect 34174 33817 34226 33826
rect 34174 33783 34183 33817
rect 34183 33783 34217 33817
rect 34217 33783 34226 33817
rect 34174 33774 34226 33783
rect 34334 33817 34386 33826
rect 34334 33783 34343 33817
rect 34343 33783 34377 33817
rect 34377 33783 34386 33817
rect 34334 33774 34386 33783
rect 34494 33817 34546 33826
rect 34494 33783 34503 33817
rect 34503 33783 34537 33817
rect 34537 33783 34546 33817
rect 34494 33774 34546 33783
rect 34654 33817 34706 33826
rect 34654 33783 34663 33817
rect 34663 33783 34697 33817
rect 34697 33783 34706 33817
rect 34654 33774 34706 33783
rect 34814 33817 34866 33826
rect 34814 33783 34823 33817
rect 34823 33783 34857 33817
rect 34857 33783 34866 33817
rect 34814 33774 34866 33783
rect 34974 33817 35026 33826
rect 34974 33783 34983 33817
rect 34983 33783 35017 33817
rect 35017 33783 35026 33817
rect 34974 33774 35026 33783
rect 35134 33817 35186 33826
rect 35134 33783 35143 33817
rect 35143 33783 35177 33817
rect 35177 33783 35186 33817
rect 35134 33774 35186 33783
rect 35294 33817 35346 33826
rect 35294 33783 35303 33817
rect 35303 33783 35337 33817
rect 35337 33783 35346 33817
rect 35294 33774 35346 33783
rect 35454 33817 35506 33826
rect 35454 33783 35463 33817
rect 35463 33783 35497 33817
rect 35497 33783 35506 33817
rect 35454 33774 35506 33783
rect 35614 33817 35666 33826
rect 35614 33783 35623 33817
rect 35623 33783 35657 33817
rect 35657 33783 35666 33817
rect 35614 33774 35666 33783
rect 35774 33817 35826 33826
rect 35774 33783 35783 33817
rect 35783 33783 35817 33817
rect 35817 33783 35826 33817
rect 35774 33774 35826 33783
rect 35934 33817 35986 33826
rect 35934 33783 35943 33817
rect 35943 33783 35977 33817
rect 35977 33783 35986 33817
rect 35934 33774 35986 33783
rect 36094 33817 36146 33826
rect 36094 33783 36103 33817
rect 36103 33783 36137 33817
rect 36137 33783 36146 33817
rect 36094 33774 36146 33783
rect 36254 33817 36306 33826
rect 36254 33783 36263 33817
rect 36263 33783 36297 33817
rect 36297 33783 36306 33817
rect 36254 33774 36306 33783
rect 36414 33817 36466 33826
rect 36414 33783 36423 33817
rect 36423 33783 36457 33817
rect 36457 33783 36466 33817
rect 36414 33774 36466 33783
rect 36574 33817 36626 33826
rect 36574 33783 36583 33817
rect 36583 33783 36617 33817
rect 36617 33783 36626 33817
rect 36574 33774 36626 33783
rect 36734 33817 36786 33826
rect 36734 33783 36743 33817
rect 36743 33783 36777 33817
rect 36777 33783 36786 33817
rect 36734 33774 36786 33783
rect 36894 33817 36946 33826
rect 36894 33783 36903 33817
rect 36903 33783 36937 33817
rect 36937 33783 36946 33817
rect 36894 33774 36946 33783
rect 37054 33817 37106 33826
rect 37054 33783 37063 33817
rect 37063 33783 37097 33817
rect 37097 33783 37106 33817
rect 37054 33774 37106 33783
rect 37214 33817 37266 33826
rect 37214 33783 37223 33817
rect 37223 33783 37257 33817
rect 37257 33783 37266 33817
rect 37214 33774 37266 33783
rect 37374 33817 37426 33826
rect 37374 33783 37383 33817
rect 37383 33783 37417 33817
rect 37417 33783 37426 33817
rect 37374 33774 37426 33783
rect 37534 33817 37586 33826
rect 37534 33783 37543 33817
rect 37543 33783 37577 33817
rect 37577 33783 37586 33817
rect 37534 33774 37586 33783
rect 37694 33817 37746 33826
rect 37694 33783 37703 33817
rect 37703 33783 37737 33817
rect 37737 33783 37746 33817
rect 37694 33774 37746 33783
rect 37854 33817 37906 33826
rect 37854 33783 37863 33817
rect 37863 33783 37897 33817
rect 37897 33783 37906 33817
rect 37854 33774 37906 33783
rect 38014 33817 38066 33826
rect 38014 33783 38023 33817
rect 38023 33783 38057 33817
rect 38057 33783 38066 33817
rect 38014 33774 38066 33783
rect 38174 33817 38226 33826
rect 38174 33783 38183 33817
rect 38183 33783 38217 33817
rect 38217 33783 38226 33817
rect 38174 33774 38226 33783
rect 38334 33817 38386 33826
rect 38334 33783 38343 33817
rect 38343 33783 38377 33817
rect 38377 33783 38386 33817
rect 38334 33774 38386 33783
rect 38494 33817 38546 33826
rect 38494 33783 38503 33817
rect 38503 33783 38537 33817
rect 38537 33783 38546 33817
rect 38494 33774 38546 33783
rect 38654 33817 38706 33826
rect 38654 33783 38663 33817
rect 38663 33783 38697 33817
rect 38697 33783 38706 33817
rect 38654 33774 38706 33783
rect 38814 33817 38866 33826
rect 38814 33783 38823 33817
rect 38823 33783 38857 33817
rect 38857 33783 38866 33817
rect 38814 33774 38866 33783
rect 38974 33817 39026 33826
rect 38974 33783 38983 33817
rect 38983 33783 39017 33817
rect 39017 33783 39026 33817
rect 38974 33774 39026 33783
rect 39134 33817 39186 33826
rect 39134 33783 39143 33817
rect 39143 33783 39177 33817
rect 39177 33783 39186 33817
rect 39134 33774 39186 33783
rect 39294 33817 39346 33826
rect 39294 33783 39303 33817
rect 39303 33783 39337 33817
rect 39337 33783 39346 33817
rect 39294 33774 39346 33783
rect 39454 33817 39506 33826
rect 39454 33783 39463 33817
rect 39463 33783 39497 33817
rect 39497 33783 39506 33817
rect 39454 33774 39506 33783
rect 39614 33817 39666 33826
rect 39614 33783 39623 33817
rect 39623 33783 39657 33817
rect 39657 33783 39666 33817
rect 39614 33774 39666 33783
rect 39774 33817 39826 33826
rect 39774 33783 39783 33817
rect 39783 33783 39817 33817
rect 39817 33783 39826 33817
rect 39774 33774 39826 33783
rect 39934 33817 39986 33826
rect 39934 33783 39943 33817
rect 39943 33783 39977 33817
rect 39977 33783 39986 33817
rect 39934 33774 39986 33783
rect 40094 33817 40146 33826
rect 40094 33783 40103 33817
rect 40103 33783 40137 33817
rect 40137 33783 40146 33817
rect 40094 33774 40146 33783
rect 40254 33817 40306 33826
rect 40254 33783 40263 33817
rect 40263 33783 40297 33817
rect 40297 33783 40306 33817
rect 40254 33774 40306 33783
rect 40414 33817 40466 33826
rect 40414 33783 40423 33817
rect 40423 33783 40457 33817
rect 40457 33783 40466 33817
rect 40414 33774 40466 33783
rect 40574 33817 40626 33826
rect 40574 33783 40583 33817
rect 40583 33783 40617 33817
rect 40617 33783 40626 33817
rect 40574 33774 40626 33783
rect 40734 33817 40786 33826
rect 40734 33783 40743 33817
rect 40743 33783 40777 33817
rect 40777 33783 40786 33817
rect 40734 33774 40786 33783
rect 40894 33817 40946 33826
rect 40894 33783 40903 33817
rect 40903 33783 40937 33817
rect 40937 33783 40946 33817
rect 40894 33774 40946 33783
rect 41054 33817 41106 33826
rect 41054 33783 41063 33817
rect 41063 33783 41097 33817
rect 41097 33783 41106 33817
rect 41054 33774 41106 33783
rect 41214 33817 41266 33826
rect 41214 33783 41223 33817
rect 41223 33783 41257 33817
rect 41257 33783 41266 33817
rect 41214 33774 41266 33783
rect 41374 33817 41426 33826
rect 41374 33783 41383 33817
rect 41383 33783 41417 33817
rect 41417 33783 41426 33817
rect 41374 33774 41426 33783
rect 41534 33817 41586 33826
rect 41534 33783 41543 33817
rect 41543 33783 41577 33817
rect 41577 33783 41586 33817
rect 41534 33774 41586 33783
rect 41694 33817 41746 33826
rect 41694 33783 41703 33817
rect 41703 33783 41737 33817
rect 41737 33783 41746 33817
rect 41694 33774 41746 33783
rect 41854 33817 41906 33826
rect 41854 33783 41863 33817
rect 41863 33783 41897 33817
rect 41897 33783 41906 33817
rect 41854 33774 41906 33783
rect 14 33497 66 33506
rect 14 33463 23 33497
rect 23 33463 57 33497
rect 57 33463 66 33497
rect 14 33454 66 33463
rect 174 33497 226 33506
rect 174 33463 183 33497
rect 183 33463 217 33497
rect 217 33463 226 33497
rect 174 33454 226 33463
rect 334 33497 386 33506
rect 334 33463 343 33497
rect 343 33463 377 33497
rect 377 33463 386 33497
rect 334 33454 386 33463
rect 494 33497 546 33506
rect 494 33463 503 33497
rect 503 33463 537 33497
rect 537 33463 546 33497
rect 494 33454 546 33463
rect 654 33497 706 33506
rect 654 33463 663 33497
rect 663 33463 697 33497
rect 697 33463 706 33497
rect 654 33454 706 33463
rect 814 33497 866 33506
rect 814 33463 823 33497
rect 823 33463 857 33497
rect 857 33463 866 33497
rect 814 33454 866 33463
rect 974 33497 1026 33506
rect 974 33463 983 33497
rect 983 33463 1017 33497
rect 1017 33463 1026 33497
rect 974 33454 1026 33463
rect 1134 33497 1186 33506
rect 1134 33463 1143 33497
rect 1143 33463 1177 33497
rect 1177 33463 1186 33497
rect 1134 33454 1186 33463
rect 1294 33497 1346 33506
rect 1294 33463 1303 33497
rect 1303 33463 1337 33497
rect 1337 33463 1346 33497
rect 1294 33454 1346 33463
rect 1454 33497 1506 33506
rect 1454 33463 1463 33497
rect 1463 33463 1497 33497
rect 1497 33463 1506 33497
rect 1454 33454 1506 33463
rect 1614 33497 1666 33506
rect 1614 33463 1623 33497
rect 1623 33463 1657 33497
rect 1657 33463 1666 33497
rect 1614 33454 1666 33463
rect 1774 33497 1826 33506
rect 1774 33463 1783 33497
rect 1783 33463 1817 33497
rect 1817 33463 1826 33497
rect 1774 33454 1826 33463
rect 1934 33497 1986 33506
rect 1934 33463 1943 33497
rect 1943 33463 1977 33497
rect 1977 33463 1986 33497
rect 1934 33454 1986 33463
rect 2094 33497 2146 33506
rect 2094 33463 2103 33497
rect 2103 33463 2137 33497
rect 2137 33463 2146 33497
rect 2094 33454 2146 33463
rect 2254 33497 2306 33506
rect 2254 33463 2263 33497
rect 2263 33463 2297 33497
rect 2297 33463 2306 33497
rect 2254 33454 2306 33463
rect 2414 33497 2466 33506
rect 2414 33463 2423 33497
rect 2423 33463 2457 33497
rect 2457 33463 2466 33497
rect 2414 33454 2466 33463
rect 2574 33497 2626 33506
rect 2574 33463 2583 33497
rect 2583 33463 2617 33497
rect 2617 33463 2626 33497
rect 2574 33454 2626 33463
rect 2734 33497 2786 33506
rect 2734 33463 2743 33497
rect 2743 33463 2777 33497
rect 2777 33463 2786 33497
rect 2734 33454 2786 33463
rect 2894 33497 2946 33506
rect 2894 33463 2903 33497
rect 2903 33463 2937 33497
rect 2937 33463 2946 33497
rect 2894 33454 2946 33463
rect 3054 33497 3106 33506
rect 3054 33463 3063 33497
rect 3063 33463 3097 33497
rect 3097 33463 3106 33497
rect 3054 33454 3106 33463
rect 3214 33497 3266 33506
rect 3214 33463 3223 33497
rect 3223 33463 3257 33497
rect 3257 33463 3266 33497
rect 3214 33454 3266 33463
rect 3374 33497 3426 33506
rect 3374 33463 3383 33497
rect 3383 33463 3417 33497
rect 3417 33463 3426 33497
rect 3374 33454 3426 33463
rect 3534 33497 3586 33506
rect 3534 33463 3543 33497
rect 3543 33463 3577 33497
rect 3577 33463 3586 33497
rect 3534 33454 3586 33463
rect 3694 33497 3746 33506
rect 3694 33463 3703 33497
rect 3703 33463 3737 33497
rect 3737 33463 3746 33497
rect 3694 33454 3746 33463
rect 3854 33497 3906 33506
rect 3854 33463 3863 33497
rect 3863 33463 3897 33497
rect 3897 33463 3906 33497
rect 3854 33454 3906 33463
rect 4014 33497 4066 33506
rect 4014 33463 4023 33497
rect 4023 33463 4057 33497
rect 4057 33463 4066 33497
rect 4014 33454 4066 33463
rect 4174 33497 4226 33506
rect 4174 33463 4183 33497
rect 4183 33463 4217 33497
rect 4217 33463 4226 33497
rect 4174 33454 4226 33463
rect 4334 33497 4386 33506
rect 4334 33463 4343 33497
rect 4343 33463 4377 33497
rect 4377 33463 4386 33497
rect 4334 33454 4386 33463
rect 4494 33497 4546 33506
rect 4494 33463 4503 33497
rect 4503 33463 4537 33497
rect 4537 33463 4546 33497
rect 4494 33454 4546 33463
rect 4654 33497 4706 33506
rect 4654 33463 4663 33497
rect 4663 33463 4697 33497
rect 4697 33463 4706 33497
rect 4654 33454 4706 33463
rect 4814 33497 4866 33506
rect 4814 33463 4823 33497
rect 4823 33463 4857 33497
rect 4857 33463 4866 33497
rect 4814 33454 4866 33463
rect 4974 33497 5026 33506
rect 4974 33463 4983 33497
rect 4983 33463 5017 33497
rect 5017 33463 5026 33497
rect 4974 33454 5026 33463
rect 5134 33497 5186 33506
rect 5134 33463 5143 33497
rect 5143 33463 5177 33497
rect 5177 33463 5186 33497
rect 5134 33454 5186 33463
rect 5294 33497 5346 33506
rect 5294 33463 5303 33497
rect 5303 33463 5337 33497
rect 5337 33463 5346 33497
rect 5294 33454 5346 33463
rect 5454 33497 5506 33506
rect 5454 33463 5463 33497
rect 5463 33463 5497 33497
rect 5497 33463 5506 33497
rect 5454 33454 5506 33463
rect 5614 33497 5666 33506
rect 5614 33463 5623 33497
rect 5623 33463 5657 33497
rect 5657 33463 5666 33497
rect 5614 33454 5666 33463
rect 5774 33497 5826 33506
rect 5774 33463 5783 33497
rect 5783 33463 5817 33497
rect 5817 33463 5826 33497
rect 5774 33454 5826 33463
rect 5934 33497 5986 33506
rect 5934 33463 5943 33497
rect 5943 33463 5977 33497
rect 5977 33463 5986 33497
rect 5934 33454 5986 33463
rect 6094 33497 6146 33506
rect 6094 33463 6103 33497
rect 6103 33463 6137 33497
rect 6137 33463 6146 33497
rect 6094 33454 6146 33463
rect 6254 33497 6306 33506
rect 6254 33463 6263 33497
rect 6263 33463 6297 33497
rect 6297 33463 6306 33497
rect 6254 33454 6306 33463
rect 6414 33497 6466 33506
rect 6414 33463 6423 33497
rect 6423 33463 6457 33497
rect 6457 33463 6466 33497
rect 6414 33454 6466 33463
rect 6574 33497 6626 33506
rect 6574 33463 6583 33497
rect 6583 33463 6617 33497
rect 6617 33463 6626 33497
rect 6574 33454 6626 33463
rect 6734 33497 6786 33506
rect 6734 33463 6743 33497
rect 6743 33463 6777 33497
rect 6777 33463 6786 33497
rect 6734 33454 6786 33463
rect 6894 33497 6946 33506
rect 6894 33463 6903 33497
rect 6903 33463 6937 33497
rect 6937 33463 6946 33497
rect 6894 33454 6946 33463
rect 7054 33497 7106 33506
rect 7054 33463 7063 33497
rect 7063 33463 7097 33497
rect 7097 33463 7106 33497
rect 7054 33454 7106 33463
rect 7214 33497 7266 33506
rect 7214 33463 7223 33497
rect 7223 33463 7257 33497
rect 7257 33463 7266 33497
rect 7214 33454 7266 33463
rect 7374 33497 7426 33506
rect 7374 33463 7383 33497
rect 7383 33463 7417 33497
rect 7417 33463 7426 33497
rect 7374 33454 7426 33463
rect 7534 33497 7586 33506
rect 7534 33463 7543 33497
rect 7543 33463 7577 33497
rect 7577 33463 7586 33497
rect 7534 33454 7586 33463
rect 7694 33497 7746 33506
rect 7694 33463 7703 33497
rect 7703 33463 7737 33497
rect 7737 33463 7746 33497
rect 7694 33454 7746 33463
rect 7854 33497 7906 33506
rect 7854 33463 7863 33497
rect 7863 33463 7897 33497
rect 7897 33463 7906 33497
rect 7854 33454 7906 33463
rect 8014 33497 8066 33506
rect 8014 33463 8023 33497
rect 8023 33463 8057 33497
rect 8057 33463 8066 33497
rect 8014 33454 8066 33463
rect 8174 33497 8226 33506
rect 8174 33463 8183 33497
rect 8183 33463 8217 33497
rect 8217 33463 8226 33497
rect 8174 33454 8226 33463
rect 8334 33497 8386 33506
rect 8334 33463 8343 33497
rect 8343 33463 8377 33497
rect 8377 33463 8386 33497
rect 8334 33454 8386 33463
rect 12494 33497 12546 33506
rect 12494 33463 12503 33497
rect 12503 33463 12537 33497
rect 12537 33463 12546 33497
rect 12494 33454 12546 33463
rect 12654 33497 12706 33506
rect 12654 33463 12663 33497
rect 12663 33463 12697 33497
rect 12697 33463 12706 33497
rect 12654 33454 12706 33463
rect 12814 33497 12866 33506
rect 12814 33463 12823 33497
rect 12823 33463 12857 33497
rect 12857 33463 12866 33497
rect 12814 33454 12866 33463
rect 12974 33497 13026 33506
rect 12974 33463 12983 33497
rect 12983 33463 13017 33497
rect 13017 33463 13026 33497
rect 12974 33454 13026 33463
rect 13134 33497 13186 33506
rect 13134 33463 13143 33497
rect 13143 33463 13177 33497
rect 13177 33463 13186 33497
rect 13134 33454 13186 33463
rect 13294 33497 13346 33506
rect 13294 33463 13303 33497
rect 13303 33463 13337 33497
rect 13337 33463 13346 33497
rect 13294 33454 13346 33463
rect 13454 33497 13506 33506
rect 13454 33463 13463 33497
rect 13463 33463 13497 33497
rect 13497 33463 13506 33497
rect 13454 33454 13506 33463
rect 13614 33497 13666 33506
rect 13614 33463 13623 33497
rect 13623 33463 13657 33497
rect 13657 33463 13666 33497
rect 13614 33454 13666 33463
rect 13774 33497 13826 33506
rect 13774 33463 13783 33497
rect 13783 33463 13817 33497
rect 13817 33463 13826 33497
rect 13774 33454 13826 33463
rect 13934 33497 13986 33506
rect 13934 33463 13943 33497
rect 13943 33463 13977 33497
rect 13977 33463 13986 33497
rect 13934 33454 13986 33463
rect 14094 33497 14146 33506
rect 14094 33463 14103 33497
rect 14103 33463 14137 33497
rect 14137 33463 14146 33497
rect 14094 33454 14146 33463
rect 14254 33497 14306 33506
rect 14254 33463 14263 33497
rect 14263 33463 14297 33497
rect 14297 33463 14306 33497
rect 14254 33454 14306 33463
rect 14414 33497 14466 33506
rect 14414 33463 14423 33497
rect 14423 33463 14457 33497
rect 14457 33463 14466 33497
rect 14414 33454 14466 33463
rect 14574 33497 14626 33506
rect 14574 33463 14583 33497
rect 14583 33463 14617 33497
rect 14617 33463 14626 33497
rect 14574 33454 14626 33463
rect 14734 33497 14786 33506
rect 14734 33463 14743 33497
rect 14743 33463 14777 33497
rect 14777 33463 14786 33497
rect 14734 33454 14786 33463
rect 14894 33497 14946 33506
rect 14894 33463 14903 33497
rect 14903 33463 14937 33497
rect 14937 33463 14946 33497
rect 14894 33454 14946 33463
rect 15054 33497 15106 33506
rect 15054 33463 15063 33497
rect 15063 33463 15097 33497
rect 15097 33463 15106 33497
rect 15054 33454 15106 33463
rect 15214 33497 15266 33506
rect 15214 33463 15223 33497
rect 15223 33463 15257 33497
rect 15257 33463 15266 33497
rect 15214 33454 15266 33463
rect 15374 33497 15426 33506
rect 15374 33463 15383 33497
rect 15383 33463 15417 33497
rect 15417 33463 15426 33497
rect 15374 33454 15426 33463
rect 15534 33497 15586 33506
rect 15534 33463 15543 33497
rect 15543 33463 15577 33497
rect 15577 33463 15586 33497
rect 15534 33454 15586 33463
rect 15694 33497 15746 33506
rect 15694 33463 15703 33497
rect 15703 33463 15737 33497
rect 15737 33463 15746 33497
rect 15694 33454 15746 33463
rect 15854 33497 15906 33506
rect 15854 33463 15863 33497
rect 15863 33463 15897 33497
rect 15897 33463 15906 33497
rect 15854 33454 15906 33463
rect 16014 33497 16066 33506
rect 16014 33463 16023 33497
rect 16023 33463 16057 33497
rect 16057 33463 16066 33497
rect 16014 33454 16066 33463
rect 16174 33497 16226 33506
rect 16174 33463 16183 33497
rect 16183 33463 16217 33497
rect 16217 33463 16226 33497
rect 16174 33454 16226 33463
rect 16334 33497 16386 33506
rect 16334 33463 16343 33497
rect 16343 33463 16377 33497
rect 16377 33463 16386 33497
rect 16334 33454 16386 33463
rect 16494 33497 16546 33506
rect 16494 33463 16503 33497
rect 16503 33463 16537 33497
rect 16537 33463 16546 33497
rect 16494 33454 16546 33463
rect 16654 33497 16706 33506
rect 16654 33463 16663 33497
rect 16663 33463 16697 33497
rect 16697 33463 16706 33497
rect 16654 33454 16706 33463
rect 16814 33497 16866 33506
rect 16814 33463 16823 33497
rect 16823 33463 16857 33497
rect 16857 33463 16866 33497
rect 16814 33454 16866 33463
rect 16974 33497 17026 33506
rect 16974 33463 16983 33497
rect 16983 33463 17017 33497
rect 17017 33463 17026 33497
rect 16974 33454 17026 33463
rect 17134 33497 17186 33506
rect 17134 33463 17143 33497
rect 17143 33463 17177 33497
rect 17177 33463 17186 33497
rect 17134 33454 17186 33463
rect 17294 33497 17346 33506
rect 17294 33463 17303 33497
rect 17303 33463 17337 33497
rect 17337 33463 17346 33497
rect 17294 33454 17346 33463
rect 17454 33497 17506 33506
rect 17454 33463 17463 33497
rect 17463 33463 17497 33497
rect 17497 33463 17506 33497
rect 17454 33454 17506 33463
rect 17614 33497 17666 33506
rect 17614 33463 17623 33497
rect 17623 33463 17657 33497
rect 17657 33463 17666 33497
rect 17614 33454 17666 33463
rect 17774 33497 17826 33506
rect 17774 33463 17783 33497
rect 17783 33463 17817 33497
rect 17817 33463 17826 33497
rect 17774 33454 17826 33463
rect 17934 33497 17986 33506
rect 17934 33463 17943 33497
rect 17943 33463 17977 33497
rect 17977 33463 17986 33497
rect 17934 33454 17986 33463
rect 18094 33497 18146 33506
rect 18094 33463 18103 33497
rect 18103 33463 18137 33497
rect 18137 33463 18146 33497
rect 18094 33454 18146 33463
rect 18254 33497 18306 33506
rect 18254 33463 18263 33497
rect 18263 33463 18297 33497
rect 18297 33463 18306 33497
rect 18254 33454 18306 33463
rect 18414 33497 18466 33506
rect 18414 33463 18423 33497
rect 18423 33463 18457 33497
rect 18457 33463 18466 33497
rect 18414 33454 18466 33463
rect 18574 33497 18626 33506
rect 18574 33463 18583 33497
rect 18583 33463 18617 33497
rect 18617 33463 18626 33497
rect 18574 33454 18626 33463
rect 18734 33497 18786 33506
rect 18734 33463 18743 33497
rect 18743 33463 18777 33497
rect 18777 33463 18786 33497
rect 18734 33454 18786 33463
rect 18894 33497 18946 33506
rect 18894 33463 18903 33497
rect 18903 33463 18937 33497
rect 18937 33463 18946 33497
rect 18894 33454 18946 33463
rect 23134 33497 23186 33506
rect 23134 33463 23143 33497
rect 23143 33463 23177 33497
rect 23177 33463 23186 33497
rect 23134 33454 23186 33463
rect 23294 33497 23346 33506
rect 23294 33463 23303 33497
rect 23303 33463 23337 33497
rect 23337 33463 23346 33497
rect 23294 33454 23346 33463
rect 23454 33497 23506 33506
rect 23454 33463 23463 33497
rect 23463 33463 23497 33497
rect 23497 33463 23506 33497
rect 23454 33454 23506 33463
rect 23614 33497 23666 33506
rect 23614 33463 23623 33497
rect 23623 33463 23657 33497
rect 23657 33463 23666 33497
rect 23614 33454 23666 33463
rect 23774 33497 23826 33506
rect 23774 33463 23783 33497
rect 23783 33463 23817 33497
rect 23817 33463 23826 33497
rect 23774 33454 23826 33463
rect 23934 33497 23986 33506
rect 23934 33463 23943 33497
rect 23943 33463 23977 33497
rect 23977 33463 23986 33497
rect 23934 33454 23986 33463
rect 24094 33497 24146 33506
rect 24094 33463 24103 33497
rect 24103 33463 24137 33497
rect 24137 33463 24146 33497
rect 24094 33454 24146 33463
rect 24254 33497 24306 33506
rect 24254 33463 24263 33497
rect 24263 33463 24297 33497
rect 24297 33463 24306 33497
rect 24254 33454 24306 33463
rect 24414 33497 24466 33506
rect 24414 33463 24423 33497
rect 24423 33463 24457 33497
rect 24457 33463 24466 33497
rect 24414 33454 24466 33463
rect 24574 33497 24626 33506
rect 24574 33463 24583 33497
rect 24583 33463 24617 33497
rect 24617 33463 24626 33497
rect 24574 33454 24626 33463
rect 24734 33497 24786 33506
rect 24734 33463 24743 33497
rect 24743 33463 24777 33497
rect 24777 33463 24786 33497
rect 24734 33454 24786 33463
rect 24894 33497 24946 33506
rect 24894 33463 24903 33497
rect 24903 33463 24937 33497
rect 24937 33463 24946 33497
rect 24894 33454 24946 33463
rect 25054 33497 25106 33506
rect 25054 33463 25063 33497
rect 25063 33463 25097 33497
rect 25097 33463 25106 33497
rect 25054 33454 25106 33463
rect 25214 33497 25266 33506
rect 25214 33463 25223 33497
rect 25223 33463 25257 33497
rect 25257 33463 25266 33497
rect 25214 33454 25266 33463
rect 25374 33497 25426 33506
rect 25374 33463 25383 33497
rect 25383 33463 25417 33497
rect 25417 33463 25426 33497
rect 25374 33454 25426 33463
rect 25534 33497 25586 33506
rect 25534 33463 25543 33497
rect 25543 33463 25577 33497
rect 25577 33463 25586 33497
rect 25534 33454 25586 33463
rect 25694 33497 25746 33506
rect 25694 33463 25703 33497
rect 25703 33463 25737 33497
rect 25737 33463 25746 33497
rect 25694 33454 25746 33463
rect 25854 33497 25906 33506
rect 25854 33463 25863 33497
rect 25863 33463 25897 33497
rect 25897 33463 25906 33497
rect 25854 33454 25906 33463
rect 26014 33497 26066 33506
rect 26014 33463 26023 33497
rect 26023 33463 26057 33497
rect 26057 33463 26066 33497
rect 26014 33454 26066 33463
rect 26174 33497 26226 33506
rect 26174 33463 26183 33497
rect 26183 33463 26217 33497
rect 26217 33463 26226 33497
rect 26174 33454 26226 33463
rect 26334 33497 26386 33506
rect 26334 33463 26343 33497
rect 26343 33463 26377 33497
rect 26377 33463 26386 33497
rect 26334 33454 26386 33463
rect 26494 33497 26546 33506
rect 26494 33463 26503 33497
rect 26503 33463 26537 33497
rect 26537 33463 26546 33497
rect 26494 33454 26546 33463
rect 26654 33497 26706 33506
rect 26654 33463 26663 33497
rect 26663 33463 26697 33497
rect 26697 33463 26706 33497
rect 26654 33454 26706 33463
rect 26814 33497 26866 33506
rect 26814 33463 26823 33497
rect 26823 33463 26857 33497
rect 26857 33463 26866 33497
rect 26814 33454 26866 33463
rect 26974 33497 27026 33506
rect 26974 33463 26983 33497
rect 26983 33463 27017 33497
rect 27017 33463 27026 33497
rect 26974 33454 27026 33463
rect 27134 33497 27186 33506
rect 27134 33463 27143 33497
rect 27143 33463 27177 33497
rect 27177 33463 27186 33497
rect 27134 33454 27186 33463
rect 27294 33497 27346 33506
rect 27294 33463 27303 33497
rect 27303 33463 27337 33497
rect 27337 33463 27346 33497
rect 27294 33454 27346 33463
rect 27454 33497 27506 33506
rect 27454 33463 27463 33497
rect 27463 33463 27497 33497
rect 27497 33463 27506 33497
rect 27454 33454 27506 33463
rect 27614 33497 27666 33506
rect 27614 33463 27623 33497
rect 27623 33463 27657 33497
rect 27657 33463 27666 33497
rect 27614 33454 27666 33463
rect 27774 33497 27826 33506
rect 27774 33463 27783 33497
rect 27783 33463 27817 33497
rect 27817 33463 27826 33497
rect 27774 33454 27826 33463
rect 27934 33497 27986 33506
rect 27934 33463 27943 33497
rect 27943 33463 27977 33497
rect 27977 33463 27986 33497
rect 27934 33454 27986 33463
rect 28094 33497 28146 33506
rect 28094 33463 28103 33497
rect 28103 33463 28137 33497
rect 28137 33463 28146 33497
rect 28094 33454 28146 33463
rect 28254 33497 28306 33506
rect 28254 33463 28263 33497
rect 28263 33463 28297 33497
rect 28297 33463 28306 33497
rect 28254 33454 28306 33463
rect 28414 33497 28466 33506
rect 28414 33463 28423 33497
rect 28423 33463 28457 33497
rect 28457 33463 28466 33497
rect 28414 33454 28466 33463
rect 28574 33497 28626 33506
rect 28574 33463 28583 33497
rect 28583 33463 28617 33497
rect 28617 33463 28626 33497
rect 28574 33454 28626 33463
rect 28734 33497 28786 33506
rect 28734 33463 28743 33497
rect 28743 33463 28777 33497
rect 28777 33463 28786 33497
rect 28734 33454 28786 33463
rect 28894 33497 28946 33506
rect 28894 33463 28903 33497
rect 28903 33463 28937 33497
rect 28937 33463 28946 33497
rect 28894 33454 28946 33463
rect 29054 33497 29106 33506
rect 29054 33463 29063 33497
rect 29063 33463 29097 33497
rect 29097 33463 29106 33497
rect 29054 33454 29106 33463
rect 29214 33497 29266 33506
rect 29214 33463 29223 33497
rect 29223 33463 29257 33497
rect 29257 33463 29266 33497
rect 29214 33454 29266 33463
rect 29374 33497 29426 33506
rect 29374 33463 29383 33497
rect 29383 33463 29417 33497
rect 29417 33463 29426 33497
rect 29374 33454 29426 33463
rect 33534 33497 33586 33506
rect 33534 33463 33543 33497
rect 33543 33463 33577 33497
rect 33577 33463 33586 33497
rect 33534 33454 33586 33463
rect 33694 33497 33746 33506
rect 33694 33463 33703 33497
rect 33703 33463 33737 33497
rect 33737 33463 33746 33497
rect 33694 33454 33746 33463
rect 33854 33497 33906 33506
rect 33854 33463 33863 33497
rect 33863 33463 33897 33497
rect 33897 33463 33906 33497
rect 33854 33454 33906 33463
rect 34014 33497 34066 33506
rect 34014 33463 34023 33497
rect 34023 33463 34057 33497
rect 34057 33463 34066 33497
rect 34014 33454 34066 33463
rect 34174 33497 34226 33506
rect 34174 33463 34183 33497
rect 34183 33463 34217 33497
rect 34217 33463 34226 33497
rect 34174 33454 34226 33463
rect 34334 33497 34386 33506
rect 34334 33463 34343 33497
rect 34343 33463 34377 33497
rect 34377 33463 34386 33497
rect 34334 33454 34386 33463
rect 34494 33497 34546 33506
rect 34494 33463 34503 33497
rect 34503 33463 34537 33497
rect 34537 33463 34546 33497
rect 34494 33454 34546 33463
rect 34654 33497 34706 33506
rect 34654 33463 34663 33497
rect 34663 33463 34697 33497
rect 34697 33463 34706 33497
rect 34654 33454 34706 33463
rect 34814 33497 34866 33506
rect 34814 33463 34823 33497
rect 34823 33463 34857 33497
rect 34857 33463 34866 33497
rect 34814 33454 34866 33463
rect 34974 33497 35026 33506
rect 34974 33463 34983 33497
rect 34983 33463 35017 33497
rect 35017 33463 35026 33497
rect 34974 33454 35026 33463
rect 35134 33497 35186 33506
rect 35134 33463 35143 33497
rect 35143 33463 35177 33497
rect 35177 33463 35186 33497
rect 35134 33454 35186 33463
rect 35294 33497 35346 33506
rect 35294 33463 35303 33497
rect 35303 33463 35337 33497
rect 35337 33463 35346 33497
rect 35294 33454 35346 33463
rect 35454 33497 35506 33506
rect 35454 33463 35463 33497
rect 35463 33463 35497 33497
rect 35497 33463 35506 33497
rect 35454 33454 35506 33463
rect 35614 33497 35666 33506
rect 35614 33463 35623 33497
rect 35623 33463 35657 33497
rect 35657 33463 35666 33497
rect 35614 33454 35666 33463
rect 35774 33497 35826 33506
rect 35774 33463 35783 33497
rect 35783 33463 35817 33497
rect 35817 33463 35826 33497
rect 35774 33454 35826 33463
rect 35934 33497 35986 33506
rect 35934 33463 35943 33497
rect 35943 33463 35977 33497
rect 35977 33463 35986 33497
rect 35934 33454 35986 33463
rect 36094 33497 36146 33506
rect 36094 33463 36103 33497
rect 36103 33463 36137 33497
rect 36137 33463 36146 33497
rect 36094 33454 36146 33463
rect 36254 33497 36306 33506
rect 36254 33463 36263 33497
rect 36263 33463 36297 33497
rect 36297 33463 36306 33497
rect 36254 33454 36306 33463
rect 36414 33497 36466 33506
rect 36414 33463 36423 33497
rect 36423 33463 36457 33497
rect 36457 33463 36466 33497
rect 36414 33454 36466 33463
rect 36574 33497 36626 33506
rect 36574 33463 36583 33497
rect 36583 33463 36617 33497
rect 36617 33463 36626 33497
rect 36574 33454 36626 33463
rect 36734 33497 36786 33506
rect 36734 33463 36743 33497
rect 36743 33463 36777 33497
rect 36777 33463 36786 33497
rect 36734 33454 36786 33463
rect 36894 33497 36946 33506
rect 36894 33463 36903 33497
rect 36903 33463 36937 33497
rect 36937 33463 36946 33497
rect 36894 33454 36946 33463
rect 37054 33497 37106 33506
rect 37054 33463 37063 33497
rect 37063 33463 37097 33497
rect 37097 33463 37106 33497
rect 37054 33454 37106 33463
rect 37214 33497 37266 33506
rect 37214 33463 37223 33497
rect 37223 33463 37257 33497
rect 37257 33463 37266 33497
rect 37214 33454 37266 33463
rect 37374 33497 37426 33506
rect 37374 33463 37383 33497
rect 37383 33463 37417 33497
rect 37417 33463 37426 33497
rect 37374 33454 37426 33463
rect 37534 33497 37586 33506
rect 37534 33463 37543 33497
rect 37543 33463 37577 33497
rect 37577 33463 37586 33497
rect 37534 33454 37586 33463
rect 37694 33497 37746 33506
rect 37694 33463 37703 33497
rect 37703 33463 37737 33497
rect 37737 33463 37746 33497
rect 37694 33454 37746 33463
rect 37854 33497 37906 33506
rect 37854 33463 37863 33497
rect 37863 33463 37897 33497
rect 37897 33463 37906 33497
rect 37854 33454 37906 33463
rect 38014 33497 38066 33506
rect 38014 33463 38023 33497
rect 38023 33463 38057 33497
rect 38057 33463 38066 33497
rect 38014 33454 38066 33463
rect 38174 33497 38226 33506
rect 38174 33463 38183 33497
rect 38183 33463 38217 33497
rect 38217 33463 38226 33497
rect 38174 33454 38226 33463
rect 38334 33497 38386 33506
rect 38334 33463 38343 33497
rect 38343 33463 38377 33497
rect 38377 33463 38386 33497
rect 38334 33454 38386 33463
rect 38494 33497 38546 33506
rect 38494 33463 38503 33497
rect 38503 33463 38537 33497
rect 38537 33463 38546 33497
rect 38494 33454 38546 33463
rect 38654 33497 38706 33506
rect 38654 33463 38663 33497
rect 38663 33463 38697 33497
rect 38697 33463 38706 33497
rect 38654 33454 38706 33463
rect 38814 33497 38866 33506
rect 38814 33463 38823 33497
rect 38823 33463 38857 33497
rect 38857 33463 38866 33497
rect 38814 33454 38866 33463
rect 38974 33497 39026 33506
rect 38974 33463 38983 33497
rect 38983 33463 39017 33497
rect 39017 33463 39026 33497
rect 38974 33454 39026 33463
rect 39134 33497 39186 33506
rect 39134 33463 39143 33497
rect 39143 33463 39177 33497
rect 39177 33463 39186 33497
rect 39134 33454 39186 33463
rect 39294 33497 39346 33506
rect 39294 33463 39303 33497
rect 39303 33463 39337 33497
rect 39337 33463 39346 33497
rect 39294 33454 39346 33463
rect 39454 33497 39506 33506
rect 39454 33463 39463 33497
rect 39463 33463 39497 33497
rect 39497 33463 39506 33497
rect 39454 33454 39506 33463
rect 39614 33497 39666 33506
rect 39614 33463 39623 33497
rect 39623 33463 39657 33497
rect 39657 33463 39666 33497
rect 39614 33454 39666 33463
rect 39774 33497 39826 33506
rect 39774 33463 39783 33497
rect 39783 33463 39817 33497
rect 39817 33463 39826 33497
rect 39774 33454 39826 33463
rect 39934 33497 39986 33506
rect 39934 33463 39943 33497
rect 39943 33463 39977 33497
rect 39977 33463 39986 33497
rect 39934 33454 39986 33463
rect 40094 33497 40146 33506
rect 40094 33463 40103 33497
rect 40103 33463 40137 33497
rect 40137 33463 40146 33497
rect 40094 33454 40146 33463
rect 40254 33497 40306 33506
rect 40254 33463 40263 33497
rect 40263 33463 40297 33497
rect 40297 33463 40306 33497
rect 40254 33454 40306 33463
rect 40414 33497 40466 33506
rect 40414 33463 40423 33497
rect 40423 33463 40457 33497
rect 40457 33463 40466 33497
rect 40414 33454 40466 33463
rect 40574 33497 40626 33506
rect 40574 33463 40583 33497
rect 40583 33463 40617 33497
rect 40617 33463 40626 33497
rect 40574 33454 40626 33463
rect 40734 33497 40786 33506
rect 40734 33463 40743 33497
rect 40743 33463 40777 33497
rect 40777 33463 40786 33497
rect 40734 33454 40786 33463
rect 40894 33497 40946 33506
rect 40894 33463 40903 33497
rect 40903 33463 40937 33497
rect 40937 33463 40946 33497
rect 40894 33454 40946 33463
rect 41054 33497 41106 33506
rect 41054 33463 41063 33497
rect 41063 33463 41097 33497
rect 41097 33463 41106 33497
rect 41054 33454 41106 33463
rect 41214 33497 41266 33506
rect 41214 33463 41223 33497
rect 41223 33463 41257 33497
rect 41257 33463 41266 33497
rect 41214 33454 41266 33463
rect 41374 33497 41426 33506
rect 41374 33463 41383 33497
rect 41383 33463 41417 33497
rect 41417 33463 41426 33497
rect 41374 33454 41426 33463
rect 41534 33497 41586 33506
rect 41534 33463 41543 33497
rect 41543 33463 41577 33497
rect 41577 33463 41586 33497
rect 41534 33454 41586 33463
rect 41694 33497 41746 33506
rect 41694 33463 41703 33497
rect 41703 33463 41737 33497
rect 41737 33463 41746 33497
rect 41694 33454 41746 33463
rect 41854 33497 41906 33506
rect 41854 33463 41863 33497
rect 41863 33463 41897 33497
rect 41897 33463 41906 33497
rect 41854 33454 41906 33463
rect 14 33337 66 33346
rect 14 33303 23 33337
rect 23 33303 57 33337
rect 57 33303 66 33337
rect 14 33294 66 33303
rect 174 33337 226 33346
rect 174 33303 183 33337
rect 183 33303 217 33337
rect 217 33303 226 33337
rect 174 33294 226 33303
rect 334 33337 386 33346
rect 334 33303 343 33337
rect 343 33303 377 33337
rect 377 33303 386 33337
rect 334 33294 386 33303
rect 494 33337 546 33346
rect 494 33303 503 33337
rect 503 33303 537 33337
rect 537 33303 546 33337
rect 494 33294 546 33303
rect 654 33337 706 33346
rect 654 33303 663 33337
rect 663 33303 697 33337
rect 697 33303 706 33337
rect 654 33294 706 33303
rect 814 33337 866 33346
rect 814 33303 823 33337
rect 823 33303 857 33337
rect 857 33303 866 33337
rect 814 33294 866 33303
rect 974 33337 1026 33346
rect 974 33303 983 33337
rect 983 33303 1017 33337
rect 1017 33303 1026 33337
rect 974 33294 1026 33303
rect 1134 33337 1186 33346
rect 1134 33303 1143 33337
rect 1143 33303 1177 33337
rect 1177 33303 1186 33337
rect 1134 33294 1186 33303
rect 1294 33337 1346 33346
rect 1294 33303 1303 33337
rect 1303 33303 1337 33337
rect 1337 33303 1346 33337
rect 1294 33294 1346 33303
rect 1454 33337 1506 33346
rect 1454 33303 1463 33337
rect 1463 33303 1497 33337
rect 1497 33303 1506 33337
rect 1454 33294 1506 33303
rect 1614 33337 1666 33346
rect 1614 33303 1623 33337
rect 1623 33303 1657 33337
rect 1657 33303 1666 33337
rect 1614 33294 1666 33303
rect 1774 33337 1826 33346
rect 1774 33303 1783 33337
rect 1783 33303 1817 33337
rect 1817 33303 1826 33337
rect 1774 33294 1826 33303
rect 1934 33337 1986 33346
rect 1934 33303 1943 33337
rect 1943 33303 1977 33337
rect 1977 33303 1986 33337
rect 1934 33294 1986 33303
rect 2094 33337 2146 33346
rect 2094 33303 2103 33337
rect 2103 33303 2137 33337
rect 2137 33303 2146 33337
rect 2094 33294 2146 33303
rect 2254 33337 2306 33346
rect 2254 33303 2263 33337
rect 2263 33303 2297 33337
rect 2297 33303 2306 33337
rect 2254 33294 2306 33303
rect 2414 33337 2466 33346
rect 2414 33303 2423 33337
rect 2423 33303 2457 33337
rect 2457 33303 2466 33337
rect 2414 33294 2466 33303
rect 2574 33337 2626 33346
rect 2574 33303 2583 33337
rect 2583 33303 2617 33337
rect 2617 33303 2626 33337
rect 2574 33294 2626 33303
rect 2734 33337 2786 33346
rect 2734 33303 2743 33337
rect 2743 33303 2777 33337
rect 2777 33303 2786 33337
rect 2734 33294 2786 33303
rect 2894 33337 2946 33346
rect 2894 33303 2903 33337
rect 2903 33303 2937 33337
rect 2937 33303 2946 33337
rect 2894 33294 2946 33303
rect 3054 33337 3106 33346
rect 3054 33303 3063 33337
rect 3063 33303 3097 33337
rect 3097 33303 3106 33337
rect 3054 33294 3106 33303
rect 3214 33337 3266 33346
rect 3214 33303 3223 33337
rect 3223 33303 3257 33337
rect 3257 33303 3266 33337
rect 3214 33294 3266 33303
rect 3374 33337 3426 33346
rect 3374 33303 3383 33337
rect 3383 33303 3417 33337
rect 3417 33303 3426 33337
rect 3374 33294 3426 33303
rect 3534 33337 3586 33346
rect 3534 33303 3543 33337
rect 3543 33303 3577 33337
rect 3577 33303 3586 33337
rect 3534 33294 3586 33303
rect 3694 33337 3746 33346
rect 3694 33303 3703 33337
rect 3703 33303 3737 33337
rect 3737 33303 3746 33337
rect 3694 33294 3746 33303
rect 3854 33337 3906 33346
rect 3854 33303 3863 33337
rect 3863 33303 3897 33337
rect 3897 33303 3906 33337
rect 3854 33294 3906 33303
rect 4014 33337 4066 33346
rect 4014 33303 4023 33337
rect 4023 33303 4057 33337
rect 4057 33303 4066 33337
rect 4014 33294 4066 33303
rect 4174 33337 4226 33346
rect 4174 33303 4183 33337
rect 4183 33303 4217 33337
rect 4217 33303 4226 33337
rect 4174 33294 4226 33303
rect 4334 33337 4386 33346
rect 4334 33303 4343 33337
rect 4343 33303 4377 33337
rect 4377 33303 4386 33337
rect 4334 33294 4386 33303
rect 4494 33337 4546 33346
rect 4494 33303 4503 33337
rect 4503 33303 4537 33337
rect 4537 33303 4546 33337
rect 4494 33294 4546 33303
rect 4654 33337 4706 33346
rect 4654 33303 4663 33337
rect 4663 33303 4697 33337
rect 4697 33303 4706 33337
rect 4654 33294 4706 33303
rect 4814 33337 4866 33346
rect 4814 33303 4823 33337
rect 4823 33303 4857 33337
rect 4857 33303 4866 33337
rect 4814 33294 4866 33303
rect 4974 33337 5026 33346
rect 4974 33303 4983 33337
rect 4983 33303 5017 33337
rect 5017 33303 5026 33337
rect 4974 33294 5026 33303
rect 5134 33337 5186 33346
rect 5134 33303 5143 33337
rect 5143 33303 5177 33337
rect 5177 33303 5186 33337
rect 5134 33294 5186 33303
rect 5294 33337 5346 33346
rect 5294 33303 5303 33337
rect 5303 33303 5337 33337
rect 5337 33303 5346 33337
rect 5294 33294 5346 33303
rect 5454 33337 5506 33346
rect 5454 33303 5463 33337
rect 5463 33303 5497 33337
rect 5497 33303 5506 33337
rect 5454 33294 5506 33303
rect 5614 33337 5666 33346
rect 5614 33303 5623 33337
rect 5623 33303 5657 33337
rect 5657 33303 5666 33337
rect 5614 33294 5666 33303
rect 5774 33337 5826 33346
rect 5774 33303 5783 33337
rect 5783 33303 5817 33337
rect 5817 33303 5826 33337
rect 5774 33294 5826 33303
rect 5934 33337 5986 33346
rect 5934 33303 5943 33337
rect 5943 33303 5977 33337
rect 5977 33303 5986 33337
rect 5934 33294 5986 33303
rect 6094 33337 6146 33346
rect 6094 33303 6103 33337
rect 6103 33303 6137 33337
rect 6137 33303 6146 33337
rect 6094 33294 6146 33303
rect 6254 33337 6306 33346
rect 6254 33303 6263 33337
rect 6263 33303 6297 33337
rect 6297 33303 6306 33337
rect 6254 33294 6306 33303
rect 6414 33337 6466 33346
rect 6414 33303 6423 33337
rect 6423 33303 6457 33337
rect 6457 33303 6466 33337
rect 6414 33294 6466 33303
rect 6574 33337 6626 33346
rect 6574 33303 6583 33337
rect 6583 33303 6617 33337
rect 6617 33303 6626 33337
rect 6574 33294 6626 33303
rect 6734 33337 6786 33346
rect 6734 33303 6743 33337
rect 6743 33303 6777 33337
rect 6777 33303 6786 33337
rect 6734 33294 6786 33303
rect 6894 33337 6946 33346
rect 6894 33303 6903 33337
rect 6903 33303 6937 33337
rect 6937 33303 6946 33337
rect 6894 33294 6946 33303
rect 7054 33337 7106 33346
rect 7054 33303 7063 33337
rect 7063 33303 7097 33337
rect 7097 33303 7106 33337
rect 7054 33294 7106 33303
rect 7214 33337 7266 33346
rect 7214 33303 7223 33337
rect 7223 33303 7257 33337
rect 7257 33303 7266 33337
rect 7214 33294 7266 33303
rect 7374 33337 7426 33346
rect 7374 33303 7383 33337
rect 7383 33303 7417 33337
rect 7417 33303 7426 33337
rect 7374 33294 7426 33303
rect 7534 33337 7586 33346
rect 7534 33303 7543 33337
rect 7543 33303 7577 33337
rect 7577 33303 7586 33337
rect 7534 33294 7586 33303
rect 7694 33337 7746 33346
rect 7694 33303 7703 33337
rect 7703 33303 7737 33337
rect 7737 33303 7746 33337
rect 7694 33294 7746 33303
rect 7854 33337 7906 33346
rect 7854 33303 7863 33337
rect 7863 33303 7897 33337
rect 7897 33303 7906 33337
rect 7854 33294 7906 33303
rect 8014 33337 8066 33346
rect 8014 33303 8023 33337
rect 8023 33303 8057 33337
rect 8057 33303 8066 33337
rect 8014 33294 8066 33303
rect 8174 33337 8226 33346
rect 8174 33303 8183 33337
rect 8183 33303 8217 33337
rect 8217 33303 8226 33337
rect 8174 33294 8226 33303
rect 8334 33337 8386 33346
rect 8334 33303 8343 33337
rect 8343 33303 8377 33337
rect 8377 33303 8386 33337
rect 8334 33294 8386 33303
rect 12494 33337 12546 33346
rect 12494 33303 12503 33337
rect 12503 33303 12537 33337
rect 12537 33303 12546 33337
rect 12494 33294 12546 33303
rect 12654 33337 12706 33346
rect 12654 33303 12663 33337
rect 12663 33303 12697 33337
rect 12697 33303 12706 33337
rect 12654 33294 12706 33303
rect 12814 33337 12866 33346
rect 12814 33303 12823 33337
rect 12823 33303 12857 33337
rect 12857 33303 12866 33337
rect 12814 33294 12866 33303
rect 12974 33337 13026 33346
rect 12974 33303 12983 33337
rect 12983 33303 13017 33337
rect 13017 33303 13026 33337
rect 12974 33294 13026 33303
rect 13134 33337 13186 33346
rect 13134 33303 13143 33337
rect 13143 33303 13177 33337
rect 13177 33303 13186 33337
rect 13134 33294 13186 33303
rect 13294 33337 13346 33346
rect 13294 33303 13303 33337
rect 13303 33303 13337 33337
rect 13337 33303 13346 33337
rect 13294 33294 13346 33303
rect 13454 33337 13506 33346
rect 13454 33303 13463 33337
rect 13463 33303 13497 33337
rect 13497 33303 13506 33337
rect 13454 33294 13506 33303
rect 13614 33337 13666 33346
rect 13614 33303 13623 33337
rect 13623 33303 13657 33337
rect 13657 33303 13666 33337
rect 13614 33294 13666 33303
rect 13774 33337 13826 33346
rect 13774 33303 13783 33337
rect 13783 33303 13817 33337
rect 13817 33303 13826 33337
rect 13774 33294 13826 33303
rect 13934 33337 13986 33346
rect 13934 33303 13943 33337
rect 13943 33303 13977 33337
rect 13977 33303 13986 33337
rect 13934 33294 13986 33303
rect 14094 33337 14146 33346
rect 14094 33303 14103 33337
rect 14103 33303 14137 33337
rect 14137 33303 14146 33337
rect 14094 33294 14146 33303
rect 14254 33337 14306 33346
rect 14254 33303 14263 33337
rect 14263 33303 14297 33337
rect 14297 33303 14306 33337
rect 14254 33294 14306 33303
rect 14414 33337 14466 33346
rect 14414 33303 14423 33337
rect 14423 33303 14457 33337
rect 14457 33303 14466 33337
rect 14414 33294 14466 33303
rect 14574 33337 14626 33346
rect 14574 33303 14583 33337
rect 14583 33303 14617 33337
rect 14617 33303 14626 33337
rect 14574 33294 14626 33303
rect 14734 33337 14786 33346
rect 14734 33303 14743 33337
rect 14743 33303 14777 33337
rect 14777 33303 14786 33337
rect 14734 33294 14786 33303
rect 14894 33337 14946 33346
rect 14894 33303 14903 33337
rect 14903 33303 14937 33337
rect 14937 33303 14946 33337
rect 14894 33294 14946 33303
rect 15054 33337 15106 33346
rect 15054 33303 15063 33337
rect 15063 33303 15097 33337
rect 15097 33303 15106 33337
rect 15054 33294 15106 33303
rect 15214 33337 15266 33346
rect 15214 33303 15223 33337
rect 15223 33303 15257 33337
rect 15257 33303 15266 33337
rect 15214 33294 15266 33303
rect 15374 33337 15426 33346
rect 15374 33303 15383 33337
rect 15383 33303 15417 33337
rect 15417 33303 15426 33337
rect 15374 33294 15426 33303
rect 15534 33337 15586 33346
rect 15534 33303 15543 33337
rect 15543 33303 15577 33337
rect 15577 33303 15586 33337
rect 15534 33294 15586 33303
rect 15694 33337 15746 33346
rect 15694 33303 15703 33337
rect 15703 33303 15737 33337
rect 15737 33303 15746 33337
rect 15694 33294 15746 33303
rect 15854 33337 15906 33346
rect 15854 33303 15863 33337
rect 15863 33303 15897 33337
rect 15897 33303 15906 33337
rect 15854 33294 15906 33303
rect 16014 33337 16066 33346
rect 16014 33303 16023 33337
rect 16023 33303 16057 33337
rect 16057 33303 16066 33337
rect 16014 33294 16066 33303
rect 16174 33337 16226 33346
rect 16174 33303 16183 33337
rect 16183 33303 16217 33337
rect 16217 33303 16226 33337
rect 16174 33294 16226 33303
rect 16334 33337 16386 33346
rect 16334 33303 16343 33337
rect 16343 33303 16377 33337
rect 16377 33303 16386 33337
rect 16334 33294 16386 33303
rect 16494 33337 16546 33346
rect 16494 33303 16503 33337
rect 16503 33303 16537 33337
rect 16537 33303 16546 33337
rect 16494 33294 16546 33303
rect 16654 33337 16706 33346
rect 16654 33303 16663 33337
rect 16663 33303 16697 33337
rect 16697 33303 16706 33337
rect 16654 33294 16706 33303
rect 16814 33337 16866 33346
rect 16814 33303 16823 33337
rect 16823 33303 16857 33337
rect 16857 33303 16866 33337
rect 16814 33294 16866 33303
rect 16974 33337 17026 33346
rect 16974 33303 16983 33337
rect 16983 33303 17017 33337
rect 17017 33303 17026 33337
rect 16974 33294 17026 33303
rect 17134 33337 17186 33346
rect 17134 33303 17143 33337
rect 17143 33303 17177 33337
rect 17177 33303 17186 33337
rect 17134 33294 17186 33303
rect 17294 33337 17346 33346
rect 17294 33303 17303 33337
rect 17303 33303 17337 33337
rect 17337 33303 17346 33337
rect 17294 33294 17346 33303
rect 17454 33337 17506 33346
rect 17454 33303 17463 33337
rect 17463 33303 17497 33337
rect 17497 33303 17506 33337
rect 17454 33294 17506 33303
rect 17614 33337 17666 33346
rect 17614 33303 17623 33337
rect 17623 33303 17657 33337
rect 17657 33303 17666 33337
rect 17614 33294 17666 33303
rect 17774 33337 17826 33346
rect 17774 33303 17783 33337
rect 17783 33303 17817 33337
rect 17817 33303 17826 33337
rect 17774 33294 17826 33303
rect 17934 33337 17986 33346
rect 17934 33303 17943 33337
rect 17943 33303 17977 33337
rect 17977 33303 17986 33337
rect 17934 33294 17986 33303
rect 18094 33337 18146 33346
rect 18094 33303 18103 33337
rect 18103 33303 18137 33337
rect 18137 33303 18146 33337
rect 18094 33294 18146 33303
rect 18254 33337 18306 33346
rect 18254 33303 18263 33337
rect 18263 33303 18297 33337
rect 18297 33303 18306 33337
rect 18254 33294 18306 33303
rect 18414 33337 18466 33346
rect 18414 33303 18423 33337
rect 18423 33303 18457 33337
rect 18457 33303 18466 33337
rect 18414 33294 18466 33303
rect 18574 33337 18626 33346
rect 18574 33303 18583 33337
rect 18583 33303 18617 33337
rect 18617 33303 18626 33337
rect 18574 33294 18626 33303
rect 18734 33337 18786 33346
rect 18734 33303 18743 33337
rect 18743 33303 18777 33337
rect 18777 33303 18786 33337
rect 18734 33294 18786 33303
rect 18894 33337 18946 33346
rect 18894 33303 18903 33337
rect 18903 33303 18937 33337
rect 18937 33303 18946 33337
rect 18894 33294 18946 33303
rect 23134 33337 23186 33346
rect 23134 33303 23143 33337
rect 23143 33303 23177 33337
rect 23177 33303 23186 33337
rect 23134 33294 23186 33303
rect 23294 33337 23346 33346
rect 23294 33303 23303 33337
rect 23303 33303 23337 33337
rect 23337 33303 23346 33337
rect 23294 33294 23346 33303
rect 23454 33337 23506 33346
rect 23454 33303 23463 33337
rect 23463 33303 23497 33337
rect 23497 33303 23506 33337
rect 23454 33294 23506 33303
rect 23614 33337 23666 33346
rect 23614 33303 23623 33337
rect 23623 33303 23657 33337
rect 23657 33303 23666 33337
rect 23614 33294 23666 33303
rect 23774 33337 23826 33346
rect 23774 33303 23783 33337
rect 23783 33303 23817 33337
rect 23817 33303 23826 33337
rect 23774 33294 23826 33303
rect 23934 33337 23986 33346
rect 23934 33303 23943 33337
rect 23943 33303 23977 33337
rect 23977 33303 23986 33337
rect 23934 33294 23986 33303
rect 24094 33337 24146 33346
rect 24094 33303 24103 33337
rect 24103 33303 24137 33337
rect 24137 33303 24146 33337
rect 24094 33294 24146 33303
rect 24254 33337 24306 33346
rect 24254 33303 24263 33337
rect 24263 33303 24297 33337
rect 24297 33303 24306 33337
rect 24254 33294 24306 33303
rect 24414 33337 24466 33346
rect 24414 33303 24423 33337
rect 24423 33303 24457 33337
rect 24457 33303 24466 33337
rect 24414 33294 24466 33303
rect 24574 33337 24626 33346
rect 24574 33303 24583 33337
rect 24583 33303 24617 33337
rect 24617 33303 24626 33337
rect 24574 33294 24626 33303
rect 24734 33337 24786 33346
rect 24734 33303 24743 33337
rect 24743 33303 24777 33337
rect 24777 33303 24786 33337
rect 24734 33294 24786 33303
rect 24894 33337 24946 33346
rect 24894 33303 24903 33337
rect 24903 33303 24937 33337
rect 24937 33303 24946 33337
rect 24894 33294 24946 33303
rect 25054 33337 25106 33346
rect 25054 33303 25063 33337
rect 25063 33303 25097 33337
rect 25097 33303 25106 33337
rect 25054 33294 25106 33303
rect 25214 33337 25266 33346
rect 25214 33303 25223 33337
rect 25223 33303 25257 33337
rect 25257 33303 25266 33337
rect 25214 33294 25266 33303
rect 25374 33337 25426 33346
rect 25374 33303 25383 33337
rect 25383 33303 25417 33337
rect 25417 33303 25426 33337
rect 25374 33294 25426 33303
rect 25534 33337 25586 33346
rect 25534 33303 25543 33337
rect 25543 33303 25577 33337
rect 25577 33303 25586 33337
rect 25534 33294 25586 33303
rect 25694 33337 25746 33346
rect 25694 33303 25703 33337
rect 25703 33303 25737 33337
rect 25737 33303 25746 33337
rect 25694 33294 25746 33303
rect 25854 33337 25906 33346
rect 25854 33303 25863 33337
rect 25863 33303 25897 33337
rect 25897 33303 25906 33337
rect 25854 33294 25906 33303
rect 26014 33337 26066 33346
rect 26014 33303 26023 33337
rect 26023 33303 26057 33337
rect 26057 33303 26066 33337
rect 26014 33294 26066 33303
rect 26174 33337 26226 33346
rect 26174 33303 26183 33337
rect 26183 33303 26217 33337
rect 26217 33303 26226 33337
rect 26174 33294 26226 33303
rect 26334 33337 26386 33346
rect 26334 33303 26343 33337
rect 26343 33303 26377 33337
rect 26377 33303 26386 33337
rect 26334 33294 26386 33303
rect 26494 33337 26546 33346
rect 26494 33303 26503 33337
rect 26503 33303 26537 33337
rect 26537 33303 26546 33337
rect 26494 33294 26546 33303
rect 26654 33337 26706 33346
rect 26654 33303 26663 33337
rect 26663 33303 26697 33337
rect 26697 33303 26706 33337
rect 26654 33294 26706 33303
rect 26814 33337 26866 33346
rect 26814 33303 26823 33337
rect 26823 33303 26857 33337
rect 26857 33303 26866 33337
rect 26814 33294 26866 33303
rect 26974 33337 27026 33346
rect 26974 33303 26983 33337
rect 26983 33303 27017 33337
rect 27017 33303 27026 33337
rect 26974 33294 27026 33303
rect 27134 33337 27186 33346
rect 27134 33303 27143 33337
rect 27143 33303 27177 33337
rect 27177 33303 27186 33337
rect 27134 33294 27186 33303
rect 27294 33337 27346 33346
rect 27294 33303 27303 33337
rect 27303 33303 27337 33337
rect 27337 33303 27346 33337
rect 27294 33294 27346 33303
rect 27454 33337 27506 33346
rect 27454 33303 27463 33337
rect 27463 33303 27497 33337
rect 27497 33303 27506 33337
rect 27454 33294 27506 33303
rect 27614 33337 27666 33346
rect 27614 33303 27623 33337
rect 27623 33303 27657 33337
rect 27657 33303 27666 33337
rect 27614 33294 27666 33303
rect 27774 33337 27826 33346
rect 27774 33303 27783 33337
rect 27783 33303 27817 33337
rect 27817 33303 27826 33337
rect 27774 33294 27826 33303
rect 27934 33337 27986 33346
rect 27934 33303 27943 33337
rect 27943 33303 27977 33337
rect 27977 33303 27986 33337
rect 27934 33294 27986 33303
rect 28094 33337 28146 33346
rect 28094 33303 28103 33337
rect 28103 33303 28137 33337
rect 28137 33303 28146 33337
rect 28094 33294 28146 33303
rect 28254 33337 28306 33346
rect 28254 33303 28263 33337
rect 28263 33303 28297 33337
rect 28297 33303 28306 33337
rect 28254 33294 28306 33303
rect 28414 33337 28466 33346
rect 28414 33303 28423 33337
rect 28423 33303 28457 33337
rect 28457 33303 28466 33337
rect 28414 33294 28466 33303
rect 28574 33337 28626 33346
rect 28574 33303 28583 33337
rect 28583 33303 28617 33337
rect 28617 33303 28626 33337
rect 28574 33294 28626 33303
rect 28734 33337 28786 33346
rect 28734 33303 28743 33337
rect 28743 33303 28777 33337
rect 28777 33303 28786 33337
rect 28734 33294 28786 33303
rect 28894 33337 28946 33346
rect 28894 33303 28903 33337
rect 28903 33303 28937 33337
rect 28937 33303 28946 33337
rect 28894 33294 28946 33303
rect 29054 33337 29106 33346
rect 29054 33303 29063 33337
rect 29063 33303 29097 33337
rect 29097 33303 29106 33337
rect 29054 33294 29106 33303
rect 29214 33337 29266 33346
rect 29214 33303 29223 33337
rect 29223 33303 29257 33337
rect 29257 33303 29266 33337
rect 29214 33294 29266 33303
rect 29374 33337 29426 33346
rect 29374 33303 29383 33337
rect 29383 33303 29417 33337
rect 29417 33303 29426 33337
rect 29374 33294 29426 33303
rect 33534 33337 33586 33346
rect 33534 33303 33543 33337
rect 33543 33303 33577 33337
rect 33577 33303 33586 33337
rect 33534 33294 33586 33303
rect 33694 33337 33746 33346
rect 33694 33303 33703 33337
rect 33703 33303 33737 33337
rect 33737 33303 33746 33337
rect 33694 33294 33746 33303
rect 33854 33337 33906 33346
rect 33854 33303 33863 33337
rect 33863 33303 33897 33337
rect 33897 33303 33906 33337
rect 33854 33294 33906 33303
rect 34014 33337 34066 33346
rect 34014 33303 34023 33337
rect 34023 33303 34057 33337
rect 34057 33303 34066 33337
rect 34014 33294 34066 33303
rect 34174 33337 34226 33346
rect 34174 33303 34183 33337
rect 34183 33303 34217 33337
rect 34217 33303 34226 33337
rect 34174 33294 34226 33303
rect 34334 33337 34386 33346
rect 34334 33303 34343 33337
rect 34343 33303 34377 33337
rect 34377 33303 34386 33337
rect 34334 33294 34386 33303
rect 34494 33337 34546 33346
rect 34494 33303 34503 33337
rect 34503 33303 34537 33337
rect 34537 33303 34546 33337
rect 34494 33294 34546 33303
rect 34654 33337 34706 33346
rect 34654 33303 34663 33337
rect 34663 33303 34697 33337
rect 34697 33303 34706 33337
rect 34654 33294 34706 33303
rect 34814 33337 34866 33346
rect 34814 33303 34823 33337
rect 34823 33303 34857 33337
rect 34857 33303 34866 33337
rect 34814 33294 34866 33303
rect 34974 33337 35026 33346
rect 34974 33303 34983 33337
rect 34983 33303 35017 33337
rect 35017 33303 35026 33337
rect 34974 33294 35026 33303
rect 35134 33337 35186 33346
rect 35134 33303 35143 33337
rect 35143 33303 35177 33337
rect 35177 33303 35186 33337
rect 35134 33294 35186 33303
rect 35294 33337 35346 33346
rect 35294 33303 35303 33337
rect 35303 33303 35337 33337
rect 35337 33303 35346 33337
rect 35294 33294 35346 33303
rect 35454 33337 35506 33346
rect 35454 33303 35463 33337
rect 35463 33303 35497 33337
rect 35497 33303 35506 33337
rect 35454 33294 35506 33303
rect 35614 33337 35666 33346
rect 35614 33303 35623 33337
rect 35623 33303 35657 33337
rect 35657 33303 35666 33337
rect 35614 33294 35666 33303
rect 35774 33337 35826 33346
rect 35774 33303 35783 33337
rect 35783 33303 35817 33337
rect 35817 33303 35826 33337
rect 35774 33294 35826 33303
rect 35934 33337 35986 33346
rect 35934 33303 35943 33337
rect 35943 33303 35977 33337
rect 35977 33303 35986 33337
rect 35934 33294 35986 33303
rect 36094 33337 36146 33346
rect 36094 33303 36103 33337
rect 36103 33303 36137 33337
rect 36137 33303 36146 33337
rect 36094 33294 36146 33303
rect 36254 33337 36306 33346
rect 36254 33303 36263 33337
rect 36263 33303 36297 33337
rect 36297 33303 36306 33337
rect 36254 33294 36306 33303
rect 36414 33337 36466 33346
rect 36414 33303 36423 33337
rect 36423 33303 36457 33337
rect 36457 33303 36466 33337
rect 36414 33294 36466 33303
rect 36574 33337 36626 33346
rect 36574 33303 36583 33337
rect 36583 33303 36617 33337
rect 36617 33303 36626 33337
rect 36574 33294 36626 33303
rect 36734 33337 36786 33346
rect 36734 33303 36743 33337
rect 36743 33303 36777 33337
rect 36777 33303 36786 33337
rect 36734 33294 36786 33303
rect 36894 33337 36946 33346
rect 36894 33303 36903 33337
rect 36903 33303 36937 33337
rect 36937 33303 36946 33337
rect 36894 33294 36946 33303
rect 37054 33337 37106 33346
rect 37054 33303 37063 33337
rect 37063 33303 37097 33337
rect 37097 33303 37106 33337
rect 37054 33294 37106 33303
rect 37214 33337 37266 33346
rect 37214 33303 37223 33337
rect 37223 33303 37257 33337
rect 37257 33303 37266 33337
rect 37214 33294 37266 33303
rect 37374 33337 37426 33346
rect 37374 33303 37383 33337
rect 37383 33303 37417 33337
rect 37417 33303 37426 33337
rect 37374 33294 37426 33303
rect 37534 33337 37586 33346
rect 37534 33303 37543 33337
rect 37543 33303 37577 33337
rect 37577 33303 37586 33337
rect 37534 33294 37586 33303
rect 37694 33337 37746 33346
rect 37694 33303 37703 33337
rect 37703 33303 37737 33337
rect 37737 33303 37746 33337
rect 37694 33294 37746 33303
rect 37854 33337 37906 33346
rect 37854 33303 37863 33337
rect 37863 33303 37897 33337
rect 37897 33303 37906 33337
rect 37854 33294 37906 33303
rect 38014 33337 38066 33346
rect 38014 33303 38023 33337
rect 38023 33303 38057 33337
rect 38057 33303 38066 33337
rect 38014 33294 38066 33303
rect 38174 33337 38226 33346
rect 38174 33303 38183 33337
rect 38183 33303 38217 33337
rect 38217 33303 38226 33337
rect 38174 33294 38226 33303
rect 38334 33337 38386 33346
rect 38334 33303 38343 33337
rect 38343 33303 38377 33337
rect 38377 33303 38386 33337
rect 38334 33294 38386 33303
rect 38494 33337 38546 33346
rect 38494 33303 38503 33337
rect 38503 33303 38537 33337
rect 38537 33303 38546 33337
rect 38494 33294 38546 33303
rect 38654 33337 38706 33346
rect 38654 33303 38663 33337
rect 38663 33303 38697 33337
rect 38697 33303 38706 33337
rect 38654 33294 38706 33303
rect 38814 33337 38866 33346
rect 38814 33303 38823 33337
rect 38823 33303 38857 33337
rect 38857 33303 38866 33337
rect 38814 33294 38866 33303
rect 38974 33337 39026 33346
rect 38974 33303 38983 33337
rect 38983 33303 39017 33337
rect 39017 33303 39026 33337
rect 38974 33294 39026 33303
rect 39134 33337 39186 33346
rect 39134 33303 39143 33337
rect 39143 33303 39177 33337
rect 39177 33303 39186 33337
rect 39134 33294 39186 33303
rect 39294 33337 39346 33346
rect 39294 33303 39303 33337
rect 39303 33303 39337 33337
rect 39337 33303 39346 33337
rect 39294 33294 39346 33303
rect 39454 33337 39506 33346
rect 39454 33303 39463 33337
rect 39463 33303 39497 33337
rect 39497 33303 39506 33337
rect 39454 33294 39506 33303
rect 39614 33337 39666 33346
rect 39614 33303 39623 33337
rect 39623 33303 39657 33337
rect 39657 33303 39666 33337
rect 39614 33294 39666 33303
rect 39774 33337 39826 33346
rect 39774 33303 39783 33337
rect 39783 33303 39817 33337
rect 39817 33303 39826 33337
rect 39774 33294 39826 33303
rect 39934 33337 39986 33346
rect 39934 33303 39943 33337
rect 39943 33303 39977 33337
rect 39977 33303 39986 33337
rect 39934 33294 39986 33303
rect 40094 33337 40146 33346
rect 40094 33303 40103 33337
rect 40103 33303 40137 33337
rect 40137 33303 40146 33337
rect 40094 33294 40146 33303
rect 40254 33337 40306 33346
rect 40254 33303 40263 33337
rect 40263 33303 40297 33337
rect 40297 33303 40306 33337
rect 40254 33294 40306 33303
rect 40414 33337 40466 33346
rect 40414 33303 40423 33337
rect 40423 33303 40457 33337
rect 40457 33303 40466 33337
rect 40414 33294 40466 33303
rect 40574 33337 40626 33346
rect 40574 33303 40583 33337
rect 40583 33303 40617 33337
rect 40617 33303 40626 33337
rect 40574 33294 40626 33303
rect 40734 33337 40786 33346
rect 40734 33303 40743 33337
rect 40743 33303 40777 33337
rect 40777 33303 40786 33337
rect 40734 33294 40786 33303
rect 40894 33337 40946 33346
rect 40894 33303 40903 33337
rect 40903 33303 40937 33337
rect 40937 33303 40946 33337
rect 40894 33294 40946 33303
rect 41054 33337 41106 33346
rect 41054 33303 41063 33337
rect 41063 33303 41097 33337
rect 41097 33303 41106 33337
rect 41054 33294 41106 33303
rect 41214 33337 41266 33346
rect 41214 33303 41223 33337
rect 41223 33303 41257 33337
rect 41257 33303 41266 33337
rect 41214 33294 41266 33303
rect 41374 33337 41426 33346
rect 41374 33303 41383 33337
rect 41383 33303 41417 33337
rect 41417 33303 41426 33337
rect 41374 33294 41426 33303
rect 41534 33337 41586 33346
rect 41534 33303 41543 33337
rect 41543 33303 41577 33337
rect 41577 33303 41586 33337
rect 41534 33294 41586 33303
rect 41694 33337 41746 33346
rect 41694 33303 41703 33337
rect 41703 33303 41737 33337
rect 41737 33303 41746 33337
rect 41694 33294 41746 33303
rect 41854 33337 41906 33346
rect 41854 33303 41863 33337
rect 41863 33303 41897 33337
rect 41897 33303 41906 33337
rect 41854 33294 41906 33303
rect 14 33017 66 33026
rect 14 32983 23 33017
rect 23 32983 57 33017
rect 57 32983 66 33017
rect 14 32974 66 32983
rect 174 33017 226 33026
rect 174 32983 183 33017
rect 183 32983 217 33017
rect 217 32983 226 33017
rect 174 32974 226 32983
rect 334 33017 386 33026
rect 334 32983 343 33017
rect 343 32983 377 33017
rect 377 32983 386 33017
rect 334 32974 386 32983
rect 494 33017 546 33026
rect 494 32983 503 33017
rect 503 32983 537 33017
rect 537 32983 546 33017
rect 494 32974 546 32983
rect 654 33017 706 33026
rect 654 32983 663 33017
rect 663 32983 697 33017
rect 697 32983 706 33017
rect 654 32974 706 32983
rect 814 33017 866 33026
rect 814 32983 823 33017
rect 823 32983 857 33017
rect 857 32983 866 33017
rect 814 32974 866 32983
rect 974 33017 1026 33026
rect 974 32983 983 33017
rect 983 32983 1017 33017
rect 1017 32983 1026 33017
rect 974 32974 1026 32983
rect 1134 33017 1186 33026
rect 1134 32983 1143 33017
rect 1143 32983 1177 33017
rect 1177 32983 1186 33017
rect 1134 32974 1186 32983
rect 1294 33017 1346 33026
rect 1294 32983 1303 33017
rect 1303 32983 1337 33017
rect 1337 32983 1346 33017
rect 1294 32974 1346 32983
rect 1454 33017 1506 33026
rect 1454 32983 1463 33017
rect 1463 32983 1497 33017
rect 1497 32983 1506 33017
rect 1454 32974 1506 32983
rect 1614 33017 1666 33026
rect 1614 32983 1623 33017
rect 1623 32983 1657 33017
rect 1657 32983 1666 33017
rect 1614 32974 1666 32983
rect 1774 33017 1826 33026
rect 1774 32983 1783 33017
rect 1783 32983 1817 33017
rect 1817 32983 1826 33017
rect 1774 32974 1826 32983
rect 1934 33017 1986 33026
rect 1934 32983 1943 33017
rect 1943 32983 1977 33017
rect 1977 32983 1986 33017
rect 1934 32974 1986 32983
rect 2094 33017 2146 33026
rect 2094 32983 2103 33017
rect 2103 32983 2137 33017
rect 2137 32983 2146 33017
rect 2094 32974 2146 32983
rect 2254 33017 2306 33026
rect 2254 32983 2263 33017
rect 2263 32983 2297 33017
rect 2297 32983 2306 33017
rect 2254 32974 2306 32983
rect 2414 33017 2466 33026
rect 2414 32983 2423 33017
rect 2423 32983 2457 33017
rect 2457 32983 2466 33017
rect 2414 32974 2466 32983
rect 2574 33017 2626 33026
rect 2574 32983 2583 33017
rect 2583 32983 2617 33017
rect 2617 32983 2626 33017
rect 2574 32974 2626 32983
rect 2734 33017 2786 33026
rect 2734 32983 2743 33017
rect 2743 32983 2777 33017
rect 2777 32983 2786 33017
rect 2734 32974 2786 32983
rect 2894 33017 2946 33026
rect 2894 32983 2903 33017
rect 2903 32983 2937 33017
rect 2937 32983 2946 33017
rect 2894 32974 2946 32983
rect 3054 33017 3106 33026
rect 3054 32983 3063 33017
rect 3063 32983 3097 33017
rect 3097 32983 3106 33017
rect 3054 32974 3106 32983
rect 3214 33017 3266 33026
rect 3214 32983 3223 33017
rect 3223 32983 3257 33017
rect 3257 32983 3266 33017
rect 3214 32974 3266 32983
rect 3374 33017 3426 33026
rect 3374 32983 3383 33017
rect 3383 32983 3417 33017
rect 3417 32983 3426 33017
rect 3374 32974 3426 32983
rect 3534 33017 3586 33026
rect 3534 32983 3543 33017
rect 3543 32983 3577 33017
rect 3577 32983 3586 33017
rect 3534 32974 3586 32983
rect 3694 33017 3746 33026
rect 3694 32983 3703 33017
rect 3703 32983 3737 33017
rect 3737 32983 3746 33017
rect 3694 32974 3746 32983
rect 3854 33017 3906 33026
rect 3854 32983 3863 33017
rect 3863 32983 3897 33017
rect 3897 32983 3906 33017
rect 3854 32974 3906 32983
rect 4014 33017 4066 33026
rect 4014 32983 4023 33017
rect 4023 32983 4057 33017
rect 4057 32983 4066 33017
rect 4014 32974 4066 32983
rect 4174 33017 4226 33026
rect 4174 32983 4183 33017
rect 4183 32983 4217 33017
rect 4217 32983 4226 33017
rect 4174 32974 4226 32983
rect 4334 33017 4386 33026
rect 4334 32983 4343 33017
rect 4343 32983 4377 33017
rect 4377 32983 4386 33017
rect 4334 32974 4386 32983
rect 4494 33017 4546 33026
rect 4494 32983 4503 33017
rect 4503 32983 4537 33017
rect 4537 32983 4546 33017
rect 4494 32974 4546 32983
rect 4654 33017 4706 33026
rect 4654 32983 4663 33017
rect 4663 32983 4697 33017
rect 4697 32983 4706 33017
rect 4654 32974 4706 32983
rect 4814 33017 4866 33026
rect 4814 32983 4823 33017
rect 4823 32983 4857 33017
rect 4857 32983 4866 33017
rect 4814 32974 4866 32983
rect 4974 33017 5026 33026
rect 4974 32983 4983 33017
rect 4983 32983 5017 33017
rect 5017 32983 5026 33017
rect 4974 32974 5026 32983
rect 5134 33017 5186 33026
rect 5134 32983 5143 33017
rect 5143 32983 5177 33017
rect 5177 32983 5186 33017
rect 5134 32974 5186 32983
rect 5294 33017 5346 33026
rect 5294 32983 5303 33017
rect 5303 32983 5337 33017
rect 5337 32983 5346 33017
rect 5294 32974 5346 32983
rect 5454 33017 5506 33026
rect 5454 32983 5463 33017
rect 5463 32983 5497 33017
rect 5497 32983 5506 33017
rect 5454 32974 5506 32983
rect 5614 33017 5666 33026
rect 5614 32983 5623 33017
rect 5623 32983 5657 33017
rect 5657 32983 5666 33017
rect 5614 32974 5666 32983
rect 5774 33017 5826 33026
rect 5774 32983 5783 33017
rect 5783 32983 5817 33017
rect 5817 32983 5826 33017
rect 5774 32974 5826 32983
rect 5934 33017 5986 33026
rect 5934 32983 5943 33017
rect 5943 32983 5977 33017
rect 5977 32983 5986 33017
rect 5934 32974 5986 32983
rect 6094 33017 6146 33026
rect 6094 32983 6103 33017
rect 6103 32983 6137 33017
rect 6137 32983 6146 33017
rect 6094 32974 6146 32983
rect 6254 33017 6306 33026
rect 6254 32983 6263 33017
rect 6263 32983 6297 33017
rect 6297 32983 6306 33017
rect 6254 32974 6306 32983
rect 6414 33017 6466 33026
rect 6414 32983 6423 33017
rect 6423 32983 6457 33017
rect 6457 32983 6466 33017
rect 6414 32974 6466 32983
rect 6574 33017 6626 33026
rect 6574 32983 6583 33017
rect 6583 32983 6617 33017
rect 6617 32983 6626 33017
rect 6574 32974 6626 32983
rect 6734 33017 6786 33026
rect 6734 32983 6743 33017
rect 6743 32983 6777 33017
rect 6777 32983 6786 33017
rect 6734 32974 6786 32983
rect 6894 33017 6946 33026
rect 6894 32983 6903 33017
rect 6903 32983 6937 33017
rect 6937 32983 6946 33017
rect 6894 32974 6946 32983
rect 7054 33017 7106 33026
rect 7054 32983 7063 33017
rect 7063 32983 7097 33017
rect 7097 32983 7106 33017
rect 7054 32974 7106 32983
rect 7214 33017 7266 33026
rect 7214 32983 7223 33017
rect 7223 32983 7257 33017
rect 7257 32983 7266 33017
rect 7214 32974 7266 32983
rect 7374 33017 7426 33026
rect 7374 32983 7383 33017
rect 7383 32983 7417 33017
rect 7417 32983 7426 33017
rect 7374 32974 7426 32983
rect 7534 33017 7586 33026
rect 7534 32983 7543 33017
rect 7543 32983 7577 33017
rect 7577 32983 7586 33017
rect 7534 32974 7586 32983
rect 7694 33017 7746 33026
rect 7694 32983 7703 33017
rect 7703 32983 7737 33017
rect 7737 32983 7746 33017
rect 7694 32974 7746 32983
rect 7854 33017 7906 33026
rect 7854 32983 7863 33017
rect 7863 32983 7897 33017
rect 7897 32983 7906 33017
rect 7854 32974 7906 32983
rect 8014 33017 8066 33026
rect 8014 32983 8023 33017
rect 8023 32983 8057 33017
rect 8057 32983 8066 33017
rect 8014 32974 8066 32983
rect 8174 33017 8226 33026
rect 8174 32983 8183 33017
rect 8183 32983 8217 33017
rect 8217 32983 8226 33017
rect 8174 32974 8226 32983
rect 8334 33017 8386 33026
rect 8334 32983 8343 33017
rect 8343 32983 8377 33017
rect 8377 32983 8386 33017
rect 8334 32974 8386 32983
rect 12494 33017 12546 33026
rect 12494 32983 12503 33017
rect 12503 32983 12537 33017
rect 12537 32983 12546 33017
rect 12494 32974 12546 32983
rect 12654 33017 12706 33026
rect 12654 32983 12663 33017
rect 12663 32983 12697 33017
rect 12697 32983 12706 33017
rect 12654 32974 12706 32983
rect 12814 33017 12866 33026
rect 12814 32983 12823 33017
rect 12823 32983 12857 33017
rect 12857 32983 12866 33017
rect 12814 32974 12866 32983
rect 12974 33017 13026 33026
rect 12974 32983 12983 33017
rect 12983 32983 13017 33017
rect 13017 32983 13026 33017
rect 12974 32974 13026 32983
rect 13134 33017 13186 33026
rect 13134 32983 13143 33017
rect 13143 32983 13177 33017
rect 13177 32983 13186 33017
rect 13134 32974 13186 32983
rect 13294 33017 13346 33026
rect 13294 32983 13303 33017
rect 13303 32983 13337 33017
rect 13337 32983 13346 33017
rect 13294 32974 13346 32983
rect 13454 33017 13506 33026
rect 13454 32983 13463 33017
rect 13463 32983 13497 33017
rect 13497 32983 13506 33017
rect 13454 32974 13506 32983
rect 13614 33017 13666 33026
rect 13614 32983 13623 33017
rect 13623 32983 13657 33017
rect 13657 32983 13666 33017
rect 13614 32974 13666 32983
rect 13774 33017 13826 33026
rect 13774 32983 13783 33017
rect 13783 32983 13817 33017
rect 13817 32983 13826 33017
rect 13774 32974 13826 32983
rect 13934 33017 13986 33026
rect 13934 32983 13943 33017
rect 13943 32983 13977 33017
rect 13977 32983 13986 33017
rect 13934 32974 13986 32983
rect 14094 33017 14146 33026
rect 14094 32983 14103 33017
rect 14103 32983 14137 33017
rect 14137 32983 14146 33017
rect 14094 32974 14146 32983
rect 14254 33017 14306 33026
rect 14254 32983 14263 33017
rect 14263 32983 14297 33017
rect 14297 32983 14306 33017
rect 14254 32974 14306 32983
rect 14414 33017 14466 33026
rect 14414 32983 14423 33017
rect 14423 32983 14457 33017
rect 14457 32983 14466 33017
rect 14414 32974 14466 32983
rect 14574 33017 14626 33026
rect 14574 32983 14583 33017
rect 14583 32983 14617 33017
rect 14617 32983 14626 33017
rect 14574 32974 14626 32983
rect 14734 33017 14786 33026
rect 14734 32983 14743 33017
rect 14743 32983 14777 33017
rect 14777 32983 14786 33017
rect 14734 32974 14786 32983
rect 14894 33017 14946 33026
rect 14894 32983 14903 33017
rect 14903 32983 14937 33017
rect 14937 32983 14946 33017
rect 14894 32974 14946 32983
rect 15054 33017 15106 33026
rect 15054 32983 15063 33017
rect 15063 32983 15097 33017
rect 15097 32983 15106 33017
rect 15054 32974 15106 32983
rect 15214 33017 15266 33026
rect 15214 32983 15223 33017
rect 15223 32983 15257 33017
rect 15257 32983 15266 33017
rect 15214 32974 15266 32983
rect 15374 33017 15426 33026
rect 15374 32983 15383 33017
rect 15383 32983 15417 33017
rect 15417 32983 15426 33017
rect 15374 32974 15426 32983
rect 15534 33017 15586 33026
rect 15534 32983 15543 33017
rect 15543 32983 15577 33017
rect 15577 32983 15586 33017
rect 15534 32974 15586 32983
rect 15694 33017 15746 33026
rect 15694 32983 15703 33017
rect 15703 32983 15737 33017
rect 15737 32983 15746 33017
rect 15694 32974 15746 32983
rect 15854 33017 15906 33026
rect 15854 32983 15863 33017
rect 15863 32983 15897 33017
rect 15897 32983 15906 33017
rect 15854 32974 15906 32983
rect 16014 33017 16066 33026
rect 16014 32983 16023 33017
rect 16023 32983 16057 33017
rect 16057 32983 16066 33017
rect 16014 32974 16066 32983
rect 16174 33017 16226 33026
rect 16174 32983 16183 33017
rect 16183 32983 16217 33017
rect 16217 32983 16226 33017
rect 16174 32974 16226 32983
rect 16334 33017 16386 33026
rect 16334 32983 16343 33017
rect 16343 32983 16377 33017
rect 16377 32983 16386 33017
rect 16334 32974 16386 32983
rect 16494 33017 16546 33026
rect 16494 32983 16503 33017
rect 16503 32983 16537 33017
rect 16537 32983 16546 33017
rect 16494 32974 16546 32983
rect 16654 33017 16706 33026
rect 16654 32983 16663 33017
rect 16663 32983 16697 33017
rect 16697 32983 16706 33017
rect 16654 32974 16706 32983
rect 16814 33017 16866 33026
rect 16814 32983 16823 33017
rect 16823 32983 16857 33017
rect 16857 32983 16866 33017
rect 16814 32974 16866 32983
rect 16974 33017 17026 33026
rect 16974 32983 16983 33017
rect 16983 32983 17017 33017
rect 17017 32983 17026 33017
rect 16974 32974 17026 32983
rect 17134 33017 17186 33026
rect 17134 32983 17143 33017
rect 17143 32983 17177 33017
rect 17177 32983 17186 33017
rect 17134 32974 17186 32983
rect 17294 33017 17346 33026
rect 17294 32983 17303 33017
rect 17303 32983 17337 33017
rect 17337 32983 17346 33017
rect 17294 32974 17346 32983
rect 17454 33017 17506 33026
rect 17454 32983 17463 33017
rect 17463 32983 17497 33017
rect 17497 32983 17506 33017
rect 17454 32974 17506 32983
rect 17614 33017 17666 33026
rect 17614 32983 17623 33017
rect 17623 32983 17657 33017
rect 17657 32983 17666 33017
rect 17614 32974 17666 32983
rect 17774 33017 17826 33026
rect 17774 32983 17783 33017
rect 17783 32983 17817 33017
rect 17817 32983 17826 33017
rect 17774 32974 17826 32983
rect 17934 33017 17986 33026
rect 17934 32983 17943 33017
rect 17943 32983 17977 33017
rect 17977 32983 17986 33017
rect 17934 32974 17986 32983
rect 18094 33017 18146 33026
rect 18094 32983 18103 33017
rect 18103 32983 18137 33017
rect 18137 32983 18146 33017
rect 18094 32974 18146 32983
rect 18254 33017 18306 33026
rect 18254 32983 18263 33017
rect 18263 32983 18297 33017
rect 18297 32983 18306 33017
rect 18254 32974 18306 32983
rect 18414 33017 18466 33026
rect 18414 32983 18423 33017
rect 18423 32983 18457 33017
rect 18457 32983 18466 33017
rect 18414 32974 18466 32983
rect 18574 33017 18626 33026
rect 18574 32983 18583 33017
rect 18583 32983 18617 33017
rect 18617 32983 18626 33017
rect 18574 32974 18626 32983
rect 18734 33017 18786 33026
rect 18734 32983 18743 33017
rect 18743 32983 18777 33017
rect 18777 32983 18786 33017
rect 18734 32974 18786 32983
rect 18894 33017 18946 33026
rect 18894 32983 18903 33017
rect 18903 32983 18937 33017
rect 18937 32983 18946 33017
rect 18894 32974 18946 32983
rect 23134 33017 23186 33026
rect 23134 32983 23143 33017
rect 23143 32983 23177 33017
rect 23177 32983 23186 33017
rect 23134 32974 23186 32983
rect 23294 33017 23346 33026
rect 23294 32983 23303 33017
rect 23303 32983 23337 33017
rect 23337 32983 23346 33017
rect 23294 32974 23346 32983
rect 23454 33017 23506 33026
rect 23454 32983 23463 33017
rect 23463 32983 23497 33017
rect 23497 32983 23506 33017
rect 23454 32974 23506 32983
rect 23614 33017 23666 33026
rect 23614 32983 23623 33017
rect 23623 32983 23657 33017
rect 23657 32983 23666 33017
rect 23614 32974 23666 32983
rect 23774 33017 23826 33026
rect 23774 32983 23783 33017
rect 23783 32983 23817 33017
rect 23817 32983 23826 33017
rect 23774 32974 23826 32983
rect 23934 33017 23986 33026
rect 23934 32983 23943 33017
rect 23943 32983 23977 33017
rect 23977 32983 23986 33017
rect 23934 32974 23986 32983
rect 24094 33017 24146 33026
rect 24094 32983 24103 33017
rect 24103 32983 24137 33017
rect 24137 32983 24146 33017
rect 24094 32974 24146 32983
rect 24254 33017 24306 33026
rect 24254 32983 24263 33017
rect 24263 32983 24297 33017
rect 24297 32983 24306 33017
rect 24254 32974 24306 32983
rect 24414 33017 24466 33026
rect 24414 32983 24423 33017
rect 24423 32983 24457 33017
rect 24457 32983 24466 33017
rect 24414 32974 24466 32983
rect 24574 33017 24626 33026
rect 24574 32983 24583 33017
rect 24583 32983 24617 33017
rect 24617 32983 24626 33017
rect 24574 32974 24626 32983
rect 24734 33017 24786 33026
rect 24734 32983 24743 33017
rect 24743 32983 24777 33017
rect 24777 32983 24786 33017
rect 24734 32974 24786 32983
rect 24894 33017 24946 33026
rect 24894 32983 24903 33017
rect 24903 32983 24937 33017
rect 24937 32983 24946 33017
rect 24894 32974 24946 32983
rect 25054 33017 25106 33026
rect 25054 32983 25063 33017
rect 25063 32983 25097 33017
rect 25097 32983 25106 33017
rect 25054 32974 25106 32983
rect 25214 33017 25266 33026
rect 25214 32983 25223 33017
rect 25223 32983 25257 33017
rect 25257 32983 25266 33017
rect 25214 32974 25266 32983
rect 25374 33017 25426 33026
rect 25374 32983 25383 33017
rect 25383 32983 25417 33017
rect 25417 32983 25426 33017
rect 25374 32974 25426 32983
rect 25534 33017 25586 33026
rect 25534 32983 25543 33017
rect 25543 32983 25577 33017
rect 25577 32983 25586 33017
rect 25534 32974 25586 32983
rect 25694 33017 25746 33026
rect 25694 32983 25703 33017
rect 25703 32983 25737 33017
rect 25737 32983 25746 33017
rect 25694 32974 25746 32983
rect 25854 33017 25906 33026
rect 25854 32983 25863 33017
rect 25863 32983 25897 33017
rect 25897 32983 25906 33017
rect 25854 32974 25906 32983
rect 26014 33017 26066 33026
rect 26014 32983 26023 33017
rect 26023 32983 26057 33017
rect 26057 32983 26066 33017
rect 26014 32974 26066 32983
rect 26174 33017 26226 33026
rect 26174 32983 26183 33017
rect 26183 32983 26217 33017
rect 26217 32983 26226 33017
rect 26174 32974 26226 32983
rect 26334 33017 26386 33026
rect 26334 32983 26343 33017
rect 26343 32983 26377 33017
rect 26377 32983 26386 33017
rect 26334 32974 26386 32983
rect 26494 33017 26546 33026
rect 26494 32983 26503 33017
rect 26503 32983 26537 33017
rect 26537 32983 26546 33017
rect 26494 32974 26546 32983
rect 26654 33017 26706 33026
rect 26654 32983 26663 33017
rect 26663 32983 26697 33017
rect 26697 32983 26706 33017
rect 26654 32974 26706 32983
rect 26814 33017 26866 33026
rect 26814 32983 26823 33017
rect 26823 32983 26857 33017
rect 26857 32983 26866 33017
rect 26814 32974 26866 32983
rect 26974 33017 27026 33026
rect 26974 32983 26983 33017
rect 26983 32983 27017 33017
rect 27017 32983 27026 33017
rect 26974 32974 27026 32983
rect 27134 33017 27186 33026
rect 27134 32983 27143 33017
rect 27143 32983 27177 33017
rect 27177 32983 27186 33017
rect 27134 32974 27186 32983
rect 27294 33017 27346 33026
rect 27294 32983 27303 33017
rect 27303 32983 27337 33017
rect 27337 32983 27346 33017
rect 27294 32974 27346 32983
rect 27454 33017 27506 33026
rect 27454 32983 27463 33017
rect 27463 32983 27497 33017
rect 27497 32983 27506 33017
rect 27454 32974 27506 32983
rect 27614 33017 27666 33026
rect 27614 32983 27623 33017
rect 27623 32983 27657 33017
rect 27657 32983 27666 33017
rect 27614 32974 27666 32983
rect 27774 33017 27826 33026
rect 27774 32983 27783 33017
rect 27783 32983 27817 33017
rect 27817 32983 27826 33017
rect 27774 32974 27826 32983
rect 27934 33017 27986 33026
rect 27934 32983 27943 33017
rect 27943 32983 27977 33017
rect 27977 32983 27986 33017
rect 27934 32974 27986 32983
rect 28094 33017 28146 33026
rect 28094 32983 28103 33017
rect 28103 32983 28137 33017
rect 28137 32983 28146 33017
rect 28094 32974 28146 32983
rect 28254 33017 28306 33026
rect 28254 32983 28263 33017
rect 28263 32983 28297 33017
rect 28297 32983 28306 33017
rect 28254 32974 28306 32983
rect 28414 33017 28466 33026
rect 28414 32983 28423 33017
rect 28423 32983 28457 33017
rect 28457 32983 28466 33017
rect 28414 32974 28466 32983
rect 28574 33017 28626 33026
rect 28574 32983 28583 33017
rect 28583 32983 28617 33017
rect 28617 32983 28626 33017
rect 28574 32974 28626 32983
rect 28734 33017 28786 33026
rect 28734 32983 28743 33017
rect 28743 32983 28777 33017
rect 28777 32983 28786 33017
rect 28734 32974 28786 32983
rect 28894 33017 28946 33026
rect 28894 32983 28903 33017
rect 28903 32983 28937 33017
rect 28937 32983 28946 33017
rect 28894 32974 28946 32983
rect 29054 33017 29106 33026
rect 29054 32983 29063 33017
rect 29063 32983 29097 33017
rect 29097 32983 29106 33017
rect 29054 32974 29106 32983
rect 29214 33017 29266 33026
rect 29214 32983 29223 33017
rect 29223 32983 29257 33017
rect 29257 32983 29266 33017
rect 29214 32974 29266 32983
rect 29374 33017 29426 33026
rect 29374 32983 29383 33017
rect 29383 32983 29417 33017
rect 29417 32983 29426 33017
rect 29374 32974 29426 32983
rect 33534 33017 33586 33026
rect 33534 32983 33543 33017
rect 33543 32983 33577 33017
rect 33577 32983 33586 33017
rect 33534 32974 33586 32983
rect 33694 33017 33746 33026
rect 33694 32983 33703 33017
rect 33703 32983 33737 33017
rect 33737 32983 33746 33017
rect 33694 32974 33746 32983
rect 33854 33017 33906 33026
rect 33854 32983 33863 33017
rect 33863 32983 33897 33017
rect 33897 32983 33906 33017
rect 33854 32974 33906 32983
rect 34014 33017 34066 33026
rect 34014 32983 34023 33017
rect 34023 32983 34057 33017
rect 34057 32983 34066 33017
rect 34014 32974 34066 32983
rect 34174 33017 34226 33026
rect 34174 32983 34183 33017
rect 34183 32983 34217 33017
rect 34217 32983 34226 33017
rect 34174 32974 34226 32983
rect 34334 33017 34386 33026
rect 34334 32983 34343 33017
rect 34343 32983 34377 33017
rect 34377 32983 34386 33017
rect 34334 32974 34386 32983
rect 34494 33017 34546 33026
rect 34494 32983 34503 33017
rect 34503 32983 34537 33017
rect 34537 32983 34546 33017
rect 34494 32974 34546 32983
rect 34654 33017 34706 33026
rect 34654 32983 34663 33017
rect 34663 32983 34697 33017
rect 34697 32983 34706 33017
rect 34654 32974 34706 32983
rect 34814 33017 34866 33026
rect 34814 32983 34823 33017
rect 34823 32983 34857 33017
rect 34857 32983 34866 33017
rect 34814 32974 34866 32983
rect 34974 33017 35026 33026
rect 34974 32983 34983 33017
rect 34983 32983 35017 33017
rect 35017 32983 35026 33017
rect 34974 32974 35026 32983
rect 35134 33017 35186 33026
rect 35134 32983 35143 33017
rect 35143 32983 35177 33017
rect 35177 32983 35186 33017
rect 35134 32974 35186 32983
rect 35294 33017 35346 33026
rect 35294 32983 35303 33017
rect 35303 32983 35337 33017
rect 35337 32983 35346 33017
rect 35294 32974 35346 32983
rect 35454 33017 35506 33026
rect 35454 32983 35463 33017
rect 35463 32983 35497 33017
rect 35497 32983 35506 33017
rect 35454 32974 35506 32983
rect 35614 33017 35666 33026
rect 35614 32983 35623 33017
rect 35623 32983 35657 33017
rect 35657 32983 35666 33017
rect 35614 32974 35666 32983
rect 35774 33017 35826 33026
rect 35774 32983 35783 33017
rect 35783 32983 35817 33017
rect 35817 32983 35826 33017
rect 35774 32974 35826 32983
rect 35934 33017 35986 33026
rect 35934 32983 35943 33017
rect 35943 32983 35977 33017
rect 35977 32983 35986 33017
rect 35934 32974 35986 32983
rect 36094 33017 36146 33026
rect 36094 32983 36103 33017
rect 36103 32983 36137 33017
rect 36137 32983 36146 33017
rect 36094 32974 36146 32983
rect 36254 33017 36306 33026
rect 36254 32983 36263 33017
rect 36263 32983 36297 33017
rect 36297 32983 36306 33017
rect 36254 32974 36306 32983
rect 36414 33017 36466 33026
rect 36414 32983 36423 33017
rect 36423 32983 36457 33017
rect 36457 32983 36466 33017
rect 36414 32974 36466 32983
rect 36574 33017 36626 33026
rect 36574 32983 36583 33017
rect 36583 32983 36617 33017
rect 36617 32983 36626 33017
rect 36574 32974 36626 32983
rect 36734 33017 36786 33026
rect 36734 32983 36743 33017
rect 36743 32983 36777 33017
rect 36777 32983 36786 33017
rect 36734 32974 36786 32983
rect 36894 33017 36946 33026
rect 36894 32983 36903 33017
rect 36903 32983 36937 33017
rect 36937 32983 36946 33017
rect 36894 32974 36946 32983
rect 37054 33017 37106 33026
rect 37054 32983 37063 33017
rect 37063 32983 37097 33017
rect 37097 32983 37106 33017
rect 37054 32974 37106 32983
rect 37214 33017 37266 33026
rect 37214 32983 37223 33017
rect 37223 32983 37257 33017
rect 37257 32983 37266 33017
rect 37214 32974 37266 32983
rect 37374 33017 37426 33026
rect 37374 32983 37383 33017
rect 37383 32983 37417 33017
rect 37417 32983 37426 33017
rect 37374 32974 37426 32983
rect 37534 33017 37586 33026
rect 37534 32983 37543 33017
rect 37543 32983 37577 33017
rect 37577 32983 37586 33017
rect 37534 32974 37586 32983
rect 37694 33017 37746 33026
rect 37694 32983 37703 33017
rect 37703 32983 37737 33017
rect 37737 32983 37746 33017
rect 37694 32974 37746 32983
rect 37854 33017 37906 33026
rect 37854 32983 37863 33017
rect 37863 32983 37897 33017
rect 37897 32983 37906 33017
rect 37854 32974 37906 32983
rect 38014 33017 38066 33026
rect 38014 32983 38023 33017
rect 38023 32983 38057 33017
rect 38057 32983 38066 33017
rect 38014 32974 38066 32983
rect 38174 33017 38226 33026
rect 38174 32983 38183 33017
rect 38183 32983 38217 33017
rect 38217 32983 38226 33017
rect 38174 32974 38226 32983
rect 38334 33017 38386 33026
rect 38334 32983 38343 33017
rect 38343 32983 38377 33017
rect 38377 32983 38386 33017
rect 38334 32974 38386 32983
rect 38494 33017 38546 33026
rect 38494 32983 38503 33017
rect 38503 32983 38537 33017
rect 38537 32983 38546 33017
rect 38494 32974 38546 32983
rect 38654 33017 38706 33026
rect 38654 32983 38663 33017
rect 38663 32983 38697 33017
rect 38697 32983 38706 33017
rect 38654 32974 38706 32983
rect 38814 33017 38866 33026
rect 38814 32983 38823 33017
rect 38823 32983 38857 33017
rect 38857 32983 38866 33017
rect 38814 32974 38866 32983
rect 38974 33017 39026 33026
rect 38974 32983 38983 33017
rect 38983 32983 39017 33017
rect 39017 32983 39026 33017
rect 38974 32974 39026 32983
rect 39134 33017 39186 33026
rect 39134 32983 39143 33017
rect 39143 32983 39177 33017
rect 39177 32983 39186 33017
rect 39134 32974 39186 32983
rect 39294 33017 39346 33026
rect 39294 32983 39303 33017
rect 39303 32983 39337 33017
rect 39337 32983 39346 33017
rect 39294 32974 39346 32983
rect 39454 33017 39506 33026
rect 39454 32983 39463 33017
rect 39463 32983 39497 33017
rect 39497 32983 39506 33017
rect 39454 32974 39506 32983
rect 39614 33017 39666 33026
rect 39614 32983 39623 33017
rect 39623 32983 39657 33017
rect 39657 32983 39666 33017
rect 39614 32974 39666 32983
rect 39774 33017 39826 33026
rect 39774 32983 39783 33017
rect 39783 32983 39817 33017
rect 39817 32983 39826 33017
rect 39774 32974 39826 32983
rect 39934 33017 39986 33026
rect 39934 32983 39943 33017
rect 39943 32983 39977 33017
rect 39977 32983 39986 33017
rect 39934 32974 39986 32983
rect 40094 33017 40146 33026
rect 40094 32983 40103 33017
rect 40103 32983 40137 33017
rect 40137 32983 40146 33017
rect 40094 32974 40146 32983
rect 40254 33017 40306 33026
rect 40254 32983 40263 33017
rect 40263 32983 40297 33017
rect 40297 32983 40306 33017
rect 40254 32974 40306 32983
rect 40414 33017 40466 33026
rect 40414 32983 40423 33017
rect 40423 32983 40457 33017
rect 40457 32983 40466 33017
rect 40414 32974 40466 32983
rect 40574 33017 40626 33026
rect 40574 32983 40583 33017
rect 40583 32983 40617 33017
rect 40617 32983 40626 33017
rect 40574 32974 40626 32983
rect 40734 33017 40786 33026
rect 40734 32983 40743 33017
rect 40743 32983 40777 33017
rect 40777 32983 40786 33017
rect 40734 32974 40786 32983
rect 40894 33017 40946 33026
rect 40894 32983 40903 33017
rect 40903 32983 40937 33017
rect 40937 32983 40946 33017
rect 40894 32974 40946 32983
rect 41054 33017 41106 33026
rect 41054 32983 41063 33017
rect 41063 32983 41097 33017
rect 41097 32983 41106 33017
rect 41054 32974 41106 32983
rect 41214 33017 41266 33026
rect 41214 32983 41223 33017
rect 41223 32983 41257 33017
rect 41257 32983 41266 33017
rect 41214 32974 41266 32983
rect 41374 33017 41426 33026
rect 41374 32983 41383 33017
rect 41383 32983 41417 33017
rect 41417 32983 41426 33017
rect 41374 32974 41426 32983
rect 41534 33017 41586 33026
rect 41534 32983 41543 33017
rect 41543 32983 41577 33017
rect 41577 32983 41586 33017
rect 41534 32974 41586 32983
rect 41694 33017 41746 33026
rect 41694 32983 41703 33017
rect 41703 32983 41737 33017
rect 41737 32983 41746 33017
rect 41694 32974 41746 32983
rect 41854 33017 41906 33026
rect 41854 32983 41863 33017
rect 41863 32983 41897 33017
rect 41897 32983 41906 33017
rect 41854 32974 41906 32983
rect 14 32857 66 32866
rect 14 32823 23 32857
rect 23 32823 57 32857
rect 57 32823 66 32857
rect 14 32814 66 32823
rect 174 32857 226 32866
rect 174 32823 183 32857
rect 183 32823 217 32857
rect 217 32823 226 32857
rect 174 32814 226 32823
rect 334 32857 386 32866
rect 334 32823 343 32857
rect 343 32823 377 32857
rect 377 32823 386 32857
rect 334 32814 386 32823
rect 494 32857 546 32866
rect 494 32823 503 32857
rect 503 32823 537 32857
rect 537 32823 546 32857
rect 494 32814 546 32823
rect 654 32857 706 32866
rect 654 32823 663 32857
rect 663 32823 697 32857
rect 697 32823 706 32857
rect 654 32814 706 32823
rect 814 32857 866 32866
rect 814 32823 823 32857
rect 823 32823 857 32857
rect 857 32823 866 32857
rect 814 32814 866 32823
rect 974 32857 1026 32866
rect 974 32823 983 32857
rect 983 32823 1017 32857
rect 1017 32823 1026 32857
rect 974 32814 1026 32823
rect 1134 32857 1186 32866
rect 1134 32823 1143 32857
rect 1143 32823 1177 32857
rect 1177 32823 1186 32857
rect 1134 32814 1186 32823
rect 1294 32857 1346 32866
rect 1294 32823 1303 32857
rect 1303 32823 1337 32857
rect 1337 32823 1346 32857
rect 1294 32814 1346 32823
rect 1454 32857 1506 32866
rect 1454 32823 1463 32857
rect 1463 32823 1497 32857
rect 1497 32823 1506 32857
rect 1454 32814 1506 32823
rect 1614 32857 1666 32866
rect 1614 32823 1623 32857
rect 1623 32823 1657 32857
rect 1657 32823 1666 32857
rect 1614 32814 1666 32823
rect 1774 32857 1826 32866
rect 1774 32823 1783 32857
rect 1783 32823 1817 32857
rect 1817 32823 1826 32857
rect 1774 32814 1826 32823
rect 1934 32857 1986 32866
rect 1934 32823 1943 32857
rect 1943 32823 1977 32857
rect 1977 32823 1986 32857
rect 1934 32814 1986 32823
rect 2094 32857 2146 32866
rect 2094 32823 2103 32857
rect 2103 32823 2137 32857
rect 2137 32823 2146 32857
rect 2094 32814 2146 32823
rect 2254 32857 2306 32866
rect 2254 32823 2263 32857
rect 2263 32823 2297 32857
rect 2297 32823 2306 32857
rect 2254 32814 2306 32823
rect 2414 32857 2466 32866
rect 2414 32823 2423 32857
rect 2423 32823 2457 32857
rect 2457 32823 2466 32857
rect 2414 32814 2466 32823
rect 2574 32857 2626 32866
rect 2574 32823 2583 32857
rect 2583 32823 2617 32857
rect 2617 32823 2626 32857
rect 2574 32814 2626 32823
rect 2734 32857 2786 32866
rect 2734 32823 2743 32857
rect 2743 32823 2777 32857
rect 2777 32823 2786 32857
rect 2734 32814 2786 32823
rect 2894 32857 2946 32866
rect 2894 32823 2903 32857
rect 2903 32823 2937 32857
rect 2937 32823 2946 32857
rect 2894 32814 2946 32823
rect 3054 32857 3106 32866
rect 3054 32823 3063 32857
rect 3063 32823 3097 32857
rect 3097 32823 3106 32857
rect 3054 32814 3106 32823
rect 3214 32857 3266 32866
rect 3214 32823 3223 32857
rect 3223 32823 3257 32857
rect 3257 32823 3266 32857
rect 3214 32814 3266 32823
rect 3374 32857 3426 32866
rect 3374 32823 3383 32857
rect 3383 32823 3417 32857
rect 3417 32823 3426 32857
rect 3374 32814 3426 32823
rect 3534 32857 3586 32866
rect 3534 32823 3543 32857
rect 3543 32823 3577 32857
rect 3577 32823 3586 32857
rect 3534 32814 3586 32823
rect 3694 32857 3746 32866
rect 3694 32823 3703 32857
rect 3703 32823 3737 32857
rect 3737 32823 3746 32857
rect 3694 32814 3746 32823
rect 3854 32857 3906 32866
rect 3854 32823 3863 32857
rect 3863 32823 3897 32857
rect 3897 32823 3906 32857
rect 3854 32814 3906 32823
rect 4014 32857 4066 32866
rect 4014 32823 4023 32857
rect 4023 32823 4057 32857
rect 4057 32823 4066 32857
rect 4014 32814 4066 32823
rect 4174 32857 4226 32866
rect 4174 32823 4183 32857
rect 4183 32823 4217 32857
rect 4217 32823 4226 32857
rect 4174 32814 4226 32823
rect 4334 32857 4386 32866
rect 4334 32823 4343 32857
rect 4343 32823 4377 32857
rect 4377 32823 4386 32857
rect 4334 32814 4386 32823
rect 4494 32857 4546 32866
rect 4494 32823 4503 32857
rect 4503 32823 4537 32857
rect 4537 32823 4546 32857
rect 4494 32814 4546 32823
rect 4654 32857 4706 32866
rect 4654 32823 4663 32857
rect 4663 32823 4697 32857
rect 4697 32823 4706 32857
rect 4654 32814 4706 32823
rect 4814 32857 4866 32866
rect 4814 32823 4823 32857
rect 4823 32823 4857 32857
rect 4857 32823 4866 32857
rect 4814 32814 4866 32823
rect 4974 32857 5026 32866
rect 4974 32823 4983 32857
rect 4983 32823 5017 32857
rect 5017 32823 5026 32857
rect 4974 32814 5026 32823
rect 5134 32857 5186 32866
rect 5134 32823 5143 32857
rect 5143 32823 5177 32857
rect 5177 32823 5186 32857
rect 5134 32814 5186 32823
rect 5294 32857 5346 32866
rect 5294 32823 5303 32857
rect 5303 32823 5337 32857
rect 5337 32823 5346 32857
rect 5294 32814 5346 32823
rect 5454 32857 5506 32866
rect 5454 32823 5463 32857
rect 5463 32823 5497 32857
rect 5497 32823 5506 32857
rect 5454 32814 5506 32823
rect 5614 32857 5666 32866
rect 5614 32823 5623 32857
rect 5623 32823 5657 32857
rect 5657 32823 5666 32857
rect 5614 32814 5666 32823
rect 5774 32857 5826 32866
rect 5774 32823 5783 32857
rect 5783 32823 5817 32857
rect 5817 32823 5826 32857
rect 5774 32814 5826 32823
rect 5934 32857 5986 32866
rect 5934 32823 5943 32857
rect 5943 32823 5977 32857
rect 5977 32823 5986 32857
rect 5934 32814 5986 32823
rect 6094 32857 6146 32866
rect 6094 32823 6103 32857
rect 6103 32823 6137 32857
rect 6137 32823 6146 32857
rect 6094 32814 6146 32823
rect 6254 32857 6306 32866
rect 6254 32823 6263 32857
rect 6263 32823 6297 32857
rect 6297 32823 6306 32857
rect 6254 32814 6306 32823
rect 6414 32857 6466 32866
rect 6414 32823 6423 32857
rect 6423 32823 6457 32857
rect 6457 32823 6466 32857
rect 6414 32814 6466 32823
rect 6574 32857 6626 32866
rect 6574 32823 6583 32857
rect 6583 32823 6617 32857
rect 6617 32823 6626 32857
rect 6574 32814 6626 32823
rect 6734 32857 6786 32866
rect 6734 32823 6743 32857
rect 6743 32823 6777 32857
rect 6777 32823 6786 32857
rect 6734 32814 6786 32823
rect 6894 32857 6946 32866
rect 6894 32823 6903 32857
rect 6903 32823 6937 32857
rect 6937 32823 6946 32857
rect 6894 32814 6946 32823
rect 7054 32857 7106 32866
rect 7054 32823 7063 32857
rect 7063 32823 7097 32857
rect 7097 32823 7106 32857
rect 7054 32814 7106 32823
rect 7214 32857 7266 32866
rect 7214 32823 7223 32857
rect 7223 32823 7257 32857
rect 7257 32823 7266 32857
rect 7214 32814 7266 32823
rect 7374 32857 7426 32866
rect 7374 32823 7383 32857
rect 7383 32823 7417 32857
rect 7417 32823 7426 32857
rect 7374 32814 7426 32823
rect 7534 32857 7586 32866
rect 7534 32823 7543 32857
rect 7543 32823 7577 32857
rect 7577 32823 7586 32857
rect 7534 32814 7586 32823
rect 7694 32857 7746 32866
rect 7694 32823 7703 32857
rect 7703 32823 7737 32857
rect 7737 32823 7746 32857
rect 7694 32814 7746 32823
rect 7854 32857 7906 32866
rect 7854 32823 7863 32857
rect 7863 32823 7897 32857
rect 7897 32823 7906 32857
rect 7854 32814 7906 32823
rect 8014 32857 8066 32866
rect 8014 32823 8023 32857
rect 8023 32823 8057 32857
rect 8057 32823 8066 32857
rect 8014 32814 8066 32823
rect 8174 32857 8226 32866
rect 8174 32823 8183 32857
rect 8183 32823 8217 32857
rect 8217 32823 8226 32857
rect 8174 32814 8226 32823
rect 8334 32857 8386 32866
rect 8334 32823 8343 32857
rect 8343 32823 8377 32857
rect 8377 32823 8386 32857
rect 8334 32814 8386 32823
rect 12494 32857 12546 32866
rect 12494 32823 12503 32857
rect 12503 32823 12537 32857
rect 12537 32823 12546 32857
rect 12494 32814 12546 32823
rect 12654 32857 12706 32866
rect 12654 32823 12663 32857
rect 12663 32823 12697 32857
rect 12697 32823 12706 32857
rect 12654 32814 12706 32823
rect 12814 32857 12866 32866
rect 12814 32823 12823 32857
rect 12823 32823 12857 32857
rect 12857 32823 12866 32857
rect 12814 32814 12866 32823
rect 12974 32857 13026 32866
rect 12974 32823 12983 32857
rect 12983 32823 13017 32857
rect 13017 32823 13026 32857
rect 12974 32814 13026 32823
rect 13134 32857 13186 32866
rect 13134 32823 13143 32857
rect 13143 32823 13177 32857
rect 13177 32823 13186 32857
rect 13134 32814 13186 32823
rect 13294 32857 13346 32866
rect 13294 32823 13303 32857
rect 13303 32823 13337 32857
rect 13337 32823 13346 32857
rect 13294 32814 13346 32823
rect 13454 32857 13506 32866
rect 13454 32823 13463 32857
rect 13463 32823 13497 32857
rect 13497 32823 13506 32857
rect 13454 32814 13506 32823
rect 13614 32857 13666 32866
rect 13614 32823 13623 32857
rect 13623 32823 13657 32857
rect 13657 32823 13666 32857
rect 13614 32814 13666 32823
rect 13774 32857 13826 32866
rect 13774 32823 13783 32857
rect 13783 32823 13817 32857
rect 13817 32823 13826 32857
rect 13774 32814 13826 32823
rect 13934 32857 13986 32866
rect 13934 32823 13943 32857
rect 13943 32823 13977 32857
rect 13977 32823 13986 32857
rect 13934 32814 13986 32823
rect 14094 32857 14146 32866
rect 14094 32823 14103 32857
rect 14103 32823 14137 32857
rect 14137 32823 14146 32857
rect 14094 32814 14146 32823
rect 14254 32857 14306 32866
rect 14254 32823 14263 32857
rect 14263 32823 14297 32857
rect 14297 32823 14306 32857
rect 14254 32814 14306 32823
rect 14414 32857 14466 32866
rect 14414 32823 14423 32857
rect 14423 32823 14457 32857
rect 14457 32823 14466 32857
rect 14414 32814 14466 32823
rect 14574 32857 14626 32866
rect 14574 32823 14583 32857
rect 14583 32823 14617 32857
rect 14617 32823 14626 32857
rect 14574 32814 14626 32823
rect 14734 32857 14786 32866
rect 14734 32823 14743 32857
rect 14743 32823 14777 32857
rect 14777 32823 14786 32857
rect 14734 32814 14786 32823
rect 14894 32857 14946 32866
rect 14894 32823 14903 32857
rect 14903 32823 14937 32857
rect 14937 32823 14946 32857
rect 14894 32814 14946 32823
rect 15054 32857 15106 32866
rect 15054 32823 15063 32857
rect 15063 32823 15097 32857
rect 15097 32823 15106 32857
rect 15054 32814 15106 32823
rect 15214 32857 15266 32866
rect 15214 32823 15223 32857
rect 15223 32823 15257 32857
rect 15257 32823 15266 32857
rect 15214 32814 15266 32823
rect 15374 32857 15426 32866
rect 15374 32823 15383 32857
rect 15383 32823 15417 32857
rect 15417 32823 15426 32857
rect 15374 32814 15426 32823
rect 15534 32857 15586 32866
rect 15534 32823 15543 32857
rect 15543 32823 15577 32857
rect 15577 32823 15586 32857
rect 15534 32814 15586 32823
rect 15694 32857 15746 32866
rect 15694 32823 15703 32857
rect 15703 32823 15737 32857
rect 15737 32823 15746 32857
rect 15694 32814 15746 32823
rect 15854 32857 15906 32866
rect 15854 32823 15863 32857
rect 15863 32823 15897 32857
rect 15897 32823 15906 32857
rect 15854 32814 15906 32823
rect 16014 32857 16066 32866
rect 16014 32823 16023 32857
rect 16023 32823 16057 32857
rect 16057 32823 16066 32857
rect 16014 32814 16066 32823
rect 16174 32857 16226 32866
rect 16174 32823 16183 32857
rect 16183 32823 16217 32857
rect 16217 32823 16226 32857
rect 16174 32814 16226 32823
rect 16334 32857 16386 32866
rect 16334 32823 16343 32857
rect 16343 32823 16377 32857
rect 16377 32823 16386 32857
rect 16334 32814 16386 32823
rect 16494 32857 16546 32866
rect 16494 32823 16503 32857
rect 16503 32823 16537 32857
rect 16537 32823 16546 32857
rect 16494 32814 16546 32823
rect 16654 32857 16706 32866
rect 16654 32823 16663 32857
rect 16663 32823 16697 32857
rect 16697 32823 16706 32857
rect 16654 32814 16706 32823
rect 16814 32857 16866 32866
rect 16814 32823 16823 32857
rect 16823 32823 16857 32857
rect 16857 32823 16866 32857
rect 16814 32814 16866 32823
rect 16974 32857 17026 32866
rect 16974 32823 16983 32857
rect 16983 32823 17017 32857
rect 17017 32823 17026 32857
rect 16974 32814 17026 32823
rect 17134 32857 17186 32866
rect 17134 32823 17143 32857
rect 17143 32823 17177 32857
rect 17177 32823 17186 32857
rect 17134 32814 17186 32823
rect 17294 32857 17346 32866
rect 17294 32823 17303 32857
rect 17303 32823 17337 32857
rect 17337 32823 17346 32857
rect 17294 32814 17346 32823
rect 17454 32857 17506 32866
rect 17454 32823 17463 32857
rect 17463 32823 17497 32857
rect 17497 32823 17506 32857
rect 17454 32814 17506 32823
rect 17614 32857 17666 32866
rect 17614 32823 17623 32857
rect 17623 32823 17657 32857
rect 17657 32823 17666 32857
rect 17614 32814 17666 32823
rect 17774 32857 17826 32866
rect 17774 32823 17783 32857
rect 17783 32823 17817 32857
rect 17817 32823 17826 32857
rect 17774 32814 17826 32823
rect 17934 32857 17986 32866
rect 17934 32823 17943 32857
rect 17943 32823 17977 32857
rect 17977 32823 17986 32857
rect 17934 32814 17986 32823
rect 18094 32857 18146 32866
rect 18094 32823 18103 32857
rect 18103 32823 18137 32857
rect 18137 32823 18146 32857
rect 18094 32814 18146 32823
rect 18254 32857 18306 32866
rect 18254 32823 18263 32857
rect 18263 32823 18297 32857
rect 18297 32823 18306 32857
rect 18254 32814 18306 32823
rect 18414 32857 18466 32866
rect 18414 32823 18423 32857
rect 18423 32823 18457 32857
rect 18457 32823 18466 32857
rect 18414 32814 18466 32823
rect 18574 32857 18626 32866
rect 18574 32823 18583 32857
rect 18583 32823 18617 32857
rect 18617 32823 18626 32857
rect 18574 32814 18626 32823
rect 18734 32857 18786 32866
rect 18734 32823 18743 32857
rect 18743 32823 18777 32857
rect 18777 32823 18786 32857
rect 18734 32814 18786 32823
rect 18894 32857 18946 32866
rect 18894 32823 18903 32857
rect 18903 32823 18937 32857
rect 18937 32823 18946 32857
rect 18894 32814 18946 32823
rect 23134 32857 23186 32866
rect 23134 32823 23143 32857
rect 23143 32823 23177 32857
rect 23177 32823 23186 32857
rect 23134 32814 23186 32823
rect 23294 32857 23346 32866
rect 23294 32823 23303 32857
rect 23303 32823 23337 32857
rect 23337 32823 23346 32857
rect 23294 32814 23346 32823
rect 23454 32857 23506 32866
rect 23454 32823 23463 32857
rect 23463 32823 23497 32857
rect 23497 32823 23506 32857
rect 23454 32814 23506 32823
rect 23614 32857 23666 32866
rect 23614 32823 23623 32857
rect 23623 32823 23657 32857
rect 23657 32823 23666 32857
rect 23614 32814 23666 32823
rect 23774 32857 23826 32866
rect 23774 32823 23783 32857
rect 23783 32823 23817 32857
rect 23817 32823 23826 32857
rect 23774 32814 23826 32823
rect 23934 32857 23986 32866
rect 23934 32823 23943 32857
rect 23943 32823 23977 32857
rect 23977 32823 23986 32857
rect 23934 32814 23986 32823
rect 24094 32857 24146 32866
rect 24094 32823 24103 32857
rect 24103 32823 24137 32857
rect 24137 32823 24146 32857
rect 24094 32814 24146 32823
rect 24254 32857 24306 32866
rect 24254 32823 24263 32857
rect 24263 32823 24297 32857
rect 24297 32823 24306 32857
rect 24254 32814 24306 32823
rect 24414 32857 24466 32866
rect 24414 32823 24423 32857
rect 24423 32823 24457 32857
rect 24457 32823 24466 32857
rect 24414 32814 24466 32823
rect 24574 32857 24626 32866
rect 24574 32823 24583 32857
rect 24583 32823 24617 32857
rect 24617 32823 24626 32857
rect 24574 32814 24626 32823
rect 24734 32857 24786 32866
rect 24734 32823 24743 32857
rect 24743 32823 24777 32857
rect 24777 32823 24786 32857
rect 24734 32814 24786 32823
rect 24894 32857 24946 32866
rect 24894 32823 24903 32857
rect 24903 32823 24937 32857
rect 24937 32823 24946 32857
rect 24894 32814 24946 32823
rect 25054 32857 25106 32866
rect 25054 32823 25063 32857
rect 25063 32823 25097 32857
rect 25097 32823 25106 32857
rect 25054 32814 25106 32823
rect 25214 32857 25266 32866
rect 25214 32823 25223 32857
rect 25223 32823 25257 32857
rect 25257 32823 25266 32857
rect 25214 32814 25266 32823
rect 25374 32857 25426 32866
rect 25374 32823 25383 32857
rect 25383 32823 25417 32857
rect 25417 32823 25426 32857
rect 25374 32814 25426 32823
rect 25534 32857 25586 32866
rect 25534 32823 25543 32857
rect 25543 32823 25577 32857
rect 25577 32823 25586 32857
rect 25534 32814 25586 32823
rect 25694 32857 25746 32866
rect 25694 32823 25703 32857
rect 25703 32823 25737 32857
rect 25737 32823 25746 32857
rect 25694 32814 25746 32823
rect 25854 32857 25906 32866
rect 25854 32823 25863 32857
rect 25863 32823 25897 32857
rect 25897 32823 25906 32857
rect 25854 32814 25906 32823
rect 26014 32857 26066 32866
rect 26014 32823 26023 32857
rect 26023 32823 26057 32857
rect 26057 32823 26066 32857
rect 26014 32814 26066 32823
rect 26174 32857 26226 32866
rect 26174 32823 26183 32857
rect 26183 32823 26217 32857
rect 26217 32823 26226 32857
rect 26174 32814 26226 32823
rect 26334 32857 26386 32866
rect 26334 32823 26343 32857
rect 26343 32823 26377 32857
rect 26377 32823 26386 32857
rect 26334 32814 26386 32823
rect 26494 32857 26546 32866
rect 26494 32823 26503 32857
rect 26503 32823 26537 32857
rect 26537 32823 26546 32857
rect 26494 32814 26546 32823
rect 26654 32857 26706 32866
rect 26654 32823 26663 32857
rect 26663 32823 26697 32857
rect 26697 32823 26706 32857
rect 26654 32814 26706 32823
rect 26814 32857 26866 32866
rect 26814 32823 26823 32857
rect 26823 32823 26857 32857
rect 26857 32823 26866 32857
rect 26814 32814 26866 32823
rect 26974 32857 27026 32866
rect 26974 32823 26983 32857
rect 26983 32823 27017 32857
rect 27017 32823 27026 32857
rect 26974 32814 27026 32823
rect 27134 32857 27186 32866
rect 27134 32823 27143 32857
rect 27143 32823 27177 32857
rect 27177 32823 27186 32857
rect 27134 32814 27186 32823
rect 27294 32857 27346 32866
rect 27294 32823 27303 32857
rect 27303 32823 27337 32857
rect 27337 32823 27346 32857
rect 27294 32814 27346 32823
rect 27454 32857 27506 32866
rect 27454 32823 27463 32857
rect 27463 32823 27497 32857
rect 27497 32823 27506 32857
rect 27454 32814 27506 32823
rect 27614 32857 27666 32866
rect 27614 32823 27623 32857
rect 27623 32823 27657 32857
rect 27657 32823 27666 32857
rect 27614 32814 27666 32823
rect 27774 32857 27826 32866
rect 27774 32823 27783 32857
rect 27783 32823 27817 32857
rect 27817 32823 27826 32857
rect 27774 32814 27826 32823
rect 27934 32857 27986 32866
rect 27934 32823 27943 32857
rect 27943 32823 27977 32857
rect 27977 32823 27986 32857
rect 27934 32814 27986 32823
rect 28094 32857 28146 32866
rect 28094 32823 28103 32857
rect 28103 32823 28137 32857
rect 28137 32823 28146 32857
rect 28094 32814 28146 32823
rect 28254 32857 28306 32866
rect 28254 32823 28263 32857
rect 28263 32823 28297 32857
rect 28297 32823 28306 32857
rect 28254 32814 28306 32823
rect 28414 32857 28466 32866
rect 28414 32823 28423 32857
rect 28423 32823 28457 32857
rect 28457 32823 28466 32857
rect 28414 32814 28466 32823
rect 28574 32857 28626 32866
rect 28574 32823 28583 32857
rect 28583 32823 28617 32857
rect 28617 32823 28626 32857
rect 28574 32814 28626 32823
rect 28734 32857 28786 32866
rect 28734 32823 28743 32857
rect 28743 32823 28777 32857
rect 28777 32823 28786 32857
rect 28734 32814 28786 32823
rect 28894 32857 28946 32866
rect 28894 32823 28903 32857
rect 28903 32823 28937 32857
rect 28937 32823 28946 32857
rect 28894 32814 28946 32823
rect 29054 32857 29106 32866
rect 29054 32823 29063 32857
rect 29063 32823 29097 32857
rect 29097 32823 29106 32857
rect 29054 32814 29106 32823
rect 29214 32857 29266 32866
rect 29214 32823 29223 32857
rect 29223 32823 29257 32857
rect 29257 32823 29266 32857
rect 29214 32814 29266 32823
rect 29374 32857 29426 32866
rect 29374 32823 29383 32857
rect 29383 32823 29417 32857
rect 29417 32823 29426 32857
rect 29374 32814 29426 32823
rect 33534 32857 33586 32866
rect 33534 32823 33543 32857
rect 33543 32823 33577 32857
rect 33577 32823 33586 32857
rect 33534 32814 33586 32823
rect 33694 32857 33746 32866
rect 33694 32823 33703 32857
rect 33703 32823 33737 32857
rect 33737 32823 33746 32857
rect 33694 32814 33746 32823
rect 33854 32857 33906 32866
rect 33854 32823 33863 32857
rect 33863 32823 33897 32857
rect 33897 32823 33906 32857
rect 33854 32814 33906 32823
rect 34014 32857 34066 32866
rect 34014 32823 34023 32857
rect 34023 32823 34057 32857
rect 34057 32823 34066 32857
rect 34014 32814 34066 32823
rect 34174 32857 34226 32866
rect 34174 32823 34183 32857
rect 34183 32823 34217 32857
rect 34217 32823 34226 32857
rect 34174 32814 34226 32823
rect 34334 32857 34386 32866
rect 34334 32823 34343 32857
rect 34343 32823 34377 32857
rect 34377 32823 34386 32857
rect 34334 32814 34386 32823
rect 34494 32857 34546 32866
rect 34494 32823 34503 32857
rect 34503 32823 34537 32857
rect 34537 32823 34546 32857
rect 34494 32814 34546 32823
rect 34654 32857 34706 32866
rect 34654 32823 34663 32857
rect 34663 32823 34697 32857
rect 34697 32823 34706 32857
rect 34654 32814 34706 32823
rect 34814 32857 34866 32866
rect 34814 32823 34823 32857
rect 34823 32823 34857 32857
rect 34857 32823 34866 32857
rect 34814 32814 34866 32823
rect 34974 32857 35026 32866
rect 34974 32823 34983 32857
rect 34983 32823 35017 32857
rect 35017 32823 35026 32857
rect 34974 32814 35026 32823
rect 35134 32857 35186 32866
rect 35134 32823 35143 32857
rect 35143 32823 35177 32857
rect 35177 32823 35186 32857
rect 35134 32814 35186 32823
rect 35294 32857 35346 32866
rect 35294 32823 35303 32857
rect 35303 32823 35337 32857
rect 35337 32823 35346 32857
rect 35294 32814 35346 32823
rect 35454 32857 35506 32866
rect 35454 32823 35463 32857
rect 35463 32823 35497 32857
rect 35497 32823 35506 32857
rect 35454 32814 35506 32823
rect 35614 32857 35666 32866
rect 35614 32823 35623 32857
rect 35623 32823 35657 32857
rect 35657 32823 35666 32857
rect 35614 32814 35666 32823
rect 35774 32857 35826 32866
rect 35774 32823 35783 32857
rect 35783 32823 35817 32857
rect 35817 32823 35826 32857
rect 35774 32814 35826 32823
rect 35934 32857 35986 32866
rect 35934 32823 35943 32857
rect 35943 32823 35977 32857
rect 35977 32823 35986 32857
rect 35934 32814 35986 32823
rect 36094 32857 36146 32866
rect 36094 32823 36103 32857
rect 36103 32823 36137 32857
rect 36137 32823 36146 32857
rect 36094 32814 36146 32823
rect 36254 32857 36306 32866
rect 36254 32823 36263 32857
rect 36263 32823 36297 32857
rect 36297 32823 36306 32857
rect 36254 32814 36306 32823
rect 36414 32857 36466 32866
rect 36414 32823 36423 32857
rect 36423 32823 36457 32857
rect 36457 32823 36466 32857
rect 36414 32814 36466 32823
rect 36574 32857 36626 32866
rect 36574 32823 36583 32857
rect 36583 32823 36617 32857
rect 36617 32823 36626 32857
rect 36574 32814 36626 32823
rect 36734 32857 36786 32866
rect 36734 32823 36743 32857
rect 36743 32823 36777 32857
rect 36777 32823 36786 32857
rect 36734 32814 36786 32823
rect 36894 32857 36946 32866
rect 36894 32823 36903 32857
rect 36903 32823 36937 32857
rect 36937 32823 36946 32857
rect 36894 32814 36946 32823
rect 37054 32857 37106 32866
rect 37054 32823 37063 32857
rect 37063 32823 37097 32857
rect 37097 32823 37106 32857
rect 37054 32814 37106 32823
rect 37214 32857 37266 32866
rect 37214 32823 37223 32857
rect 37223 32823 37257 32857
rect 37257 32823 37266 32857
rect 37214 32814 37266 32823
rect 37374 32857 37426 32866
rect 37374 32823 37383 32857
rect 37383 32823 37417 32857
rect 37417 32823 37426 32857
rect 37374 32814 37426 32823
rect 37534 32857 37586 32866
rect 37534 32823 37543 32857
rect 37543 32823 37577 32857
rect 37577 32823 37586 32857
rect 37534 32814 37586 32823
rect 37694 32857 37746 32866
rect 37694 32823 37703 32857
rect 37703 32823 37737 32857
rect 37737 32823 37746 32857
rect 37694 32814 37746 32823
rect 37854 32857 37906 32866
rect 37854 32823 37863 32857
rect 37863 32823 37897 32857
rect 37897 32823 37906 32857
rect 37854 32814 37906 32823
rect 38014 32857 38066 32866
rect 38014 32823 38023 32857
rect 38023 32823 38057 32857
rect 38057 32823 38066 32857
rect 38014 32814 38066 32823
rect 38174 32857 38226 32866
rect 38174 32823 38183 32857
rect 38183 32823 38217 32857
rect 38217 32823 38226 32857
rect 38174 32814 38226 32823
rect 38334 32857 38386 32866
rect 38334 32823 38343 32857
rect 38343 32823 38377 32857
rect 38377 32823 38386 32857
rect 38334 32814 38386 32823
rect 38494 32857 38546 32866
rect 38494 32823 38503 32857
rect 38503 32823 38537 32857
rect 38537 32823 38546 32857
rect 38494 32814 38546 32823
rect 38654 32857 38706 32866
rect 38654 32823 38663 32857
rect 38663 32823 38697 32857
rect 38697 32823 38706 32857
rect 38654 32814 38706 32823
rect 38814 32857 38866 32866
rect 38814 32823 38823 32857
rect 38823 32823 38857 32857
rect 38857 32823 38866 32857
rect 38814 32814 38866 32823
rect 38974 32857 39026 32866
rect 38974 32823 38983 32857
rect 38983 32823 39017 32857
rect 39017 32823 39026 32857
rect 38974 32814 39026 32823
rect 39134 32857 39186 32866
rect 39134 32823 39143 32857
rect 39143 32823 39177 32857
rect 39177 32823 39186 32857
rect 39134 32814 39186 32823
rect 39294 32857 39346 32866
rect 39294 32823 39303 32857
rect 39303 32823 39337 32857
rect 39337 32823 39346 32857
rect 39294 32814 39346 32823
rect 39454 32857 39506 32866
rect 39454 32823 39463 32857
rect 39463 32823 39497 32857
rect 39497 32823 39506 32857
rect 39454 32814 39506 32823
rect 39614 32857 39666 32866
rect 39614 32823 39623 32857
rect 39623 32823 39657 32857
rect 39657 32823 39666 32857
rect 39614 32814 39666 32823
rect 39774 32857 39826 32866
rect 39774 32823 39783 32857
rect 39783 32823 39817 32857
rect 39817 32823 39826 32857
rect 39774 32814 39826 32823
rect 39934 32857 39986 32866
rect 39934 32823 39943 32857
rect 39943 32823 39977 32857
rect 39977 32823 39986 32857
rect 39934 32814 39986 32823
rect 40094 32857 40146 32866
rect 40094 32823 40103 32857
rect 40103 32823 40137 32857
rect 40137 32823 40146 32857
rect 40094 32814 40146 32823
rect 40254 32857 40306 32866
rect 40254 32823 40263 32857
rect 40263 32823 40297 32857
rect 40297 32823 40306 32857
rect 40254 32814 40306 32823
rect 40414 32857 40466 32866
rect 40414 32823 40423 32857
rect 40423 32823 40457 32857
rect 40457 32823 40466 32857
rect 40414 32814 40466 32823
rect 40574 32857 40626 32866
rect 40574 32823 40583 32857
rect 40583 32823 40617 32857
rect 40617 32823 40626 32857
rect 40574 32814 40626 32823
rect 40734 32857 40786 32866
rect 40734 32823 40743 32857
rect 40743 32823 40777 32857
rect 40777 32823 40786 32857
rect 40734 32814 40786 32823
rect 40894 32857 40946 32866
rect 40894 32823 40903 32857
rect 40903 32823 40937 32857
rect 40937 32823 40946 32857
rect 40894 32814 40946 32823
rect 41054 32857 41106 32866
rect 41054 32823 41063 32857
rect 41063 32823 41097 32857
rect 41097 32823 41106 32857
rect 41054 32814 41106 32823
rect 41214 32857 41266 32866
rect 41214 32823 41223 32857
rect 41223 32823 41257 32857
rect 41257 32823 41266 32857
rect 41214 32814 41266 32823
rect 41374 32857 41426 32866
rect 41374 32823 41383 32857
rect 41383 32823 41417 32857
rect 41417 32823 41426 32857
rect 41374 32814 41426 32823
rect 41534 32857 41586 32866
rect 41534 32823 41543 32857
rect 41543 32823 41577 32857
rect 41577 32823 41586 32857
rect 41534 32814 41586 32823
rect 41694 32857 41746 32866
rect 41694 32823 41703 32857
rect 41703 32823 41737 32857
rect 41737 32823 41746 32857
rect 41694 32814 41746 32823
rect 41854 32857 41906 32866
rect 41854 32823 41863 32857
rect 41863 32823 41897 32857
rect 41897 32823 41906 32857
rect 41854 32814 41906 32823
rect 14 32537 66 32546
rect 14 32503 23 32537
rect 23 32503 57 32537
rect 57 32503 66 32537
rect 14 32494 66 32503
rect 174 32537 226 32546
rect 174 32503 183 32537
rect 183 32503 217 32537
rect 217 32503 226 32537
rect 174 32494 226 32503
rect 334 32537 386 32546
rect 334 32503 343 32537
rect 343 32503 377 32537
rect 377 32503 386 32537
rect 334 32494 386 32503
rect 494 32537 546 32546
rect 494 32503 503 32537
rect 503 32503 537 32537
rect 537 32503 546 32537
rect 494 32494 546 32503
rect 654 32537 706 32546
rect 654 32503 663 32537
rect 663 32503 697 32537
rect 697 32503 706 32537
rect 654 32494 706 32503
rect 814 32537 866 32546
rect 814 32503 823 32537
rect 823 32503 857 32537
rect 857 32503 866 32537
rect 814 32494 866 32503
rect 974 32537 1026 32546
rect 974 32503 983 32537
rect 983 32503 1017 32537
rect 1017 32503 1026 32537
rect 974 32494 1026 32503
rect 1134 32537 1186 32546
rect 1134 32503 1143 32537
rect 1143 32503 1177 32537
rect 1177 32503 1186 32537
rect 1134 32494 1186 32503
rect 1294 32537 1346 32546
rect 1294 32503 1303 32537
rect 1303 32503 1337 32537
rect 1337 32503 1346 32537
rect 1294 32494 1346 32503
rect 1454 32537 1506 32546
rect 1454 32503 1463 32537
rect 1463 32503 1497 32537
rect 1497 32503 1506 32537
rect 1454 32494 1506 32503
rect 1614 32537 1666 32546
rect 1614 32503 1623 32537
rect 1623 32503 1657 32537
rect 1657 32503 1666 32537
rect 1614 32494 1666 32503
rect 1774 32537 1826 32546
rect 1774 32503 1783 32537
rect 1783 32503 1817 32537
rect 1817 32503 1826 32537
rect 1774 32494 1826 32503
rect 1934 32537 1986 32546
rect 1934 32503 1943 32537
rect 1943 32503 1977 32537
rect 1977 32503 1986 32537
rect 1934 32494 1986 32503
rect 2094 32537 2146 32546
rect 2094 32503 2103 32537
rect 2103 32503 2137 32537
rect 2137 32503 2146 32537
rect 2094 32494 2146 32503
rect 2254 32537 2306 32546
rect 2254 32503 2263 32537
rect 2263 32503 2297 32537
rect 2297 32503 2306 32537
rect 2254 32494 2306 32503
rect 2414 32537 2466 32546
rect 2414 32503 2423 32537
rect 2423 32503 2457 32537
rect 2457 32503 2466 32537
rect 2414 32494 2466 32503
rect 2574 32537 2626 32546
rect 2574 32503 2583 32537
rect 2583 32503 2617 32537
rect 2617 32503 2626 32537
rect 2574 32494 2626 32503
rect 2734 32537 2786 32546
rect 2734 32503 2743 32537
rect 2743 32503 2777 32537
rect 2777 32503 2786 32537
rect 2734 32494 2786 32503
rect 2894 32537 2946 32546
rect 2894 32503 2903 32537
rect 2903 32503 2937 32537
rect 2937 32503 2946 32537
rect 2894 32494 2946 32503
rect 3054 32537 3106 32546
rect 3054 32503 3063 32537
rect 3063 32503 3097 32537
rect 3097 32503 3106 32537
rect 3054 32494 3106 32503
rect 3214 32537 3266 32546
rect 3214 32503 3223 32537
rect 3223 32503 3257 32537
rect 3257 32503 3266 32537
rect 3214 32494 3266 32503
rect 3374 32537 3426 32546
rect 3374 32503 3383 32537
rect 3383 32503 3417 32537
rect 3417 32503 3426 32537
rect 3374 32494 3426 32503
rect 3534 32537 3586 32546
rect 3534 32503 3543 32537
rect 3543 32503 3577 32537
rect 3577 32503 3586 32537
rect 3534 32494 3586 32503
rect 3694 32537 3746 32546
rect 3694 32503 3703 32537
rect 3703 32503 3737 32537
rect 3737 32503 3746 32537
rect 3694 32494 3746 32503
rect 3854 32537 3906 32546
rect 3854 32503 3863 32537
rect 3863 32503 3897 32537
rect 3897 32503 3906 32537
rect 3854 32494 3906 32503
rect 4014 32537 4066 32546
rect 4014 32503 4023 32537
rect 4023 32503 4057 32537
rect 4057 32503 4066 32537
rect 4014 32494 4066 32503
rect 4174 32537 4226 32546
rect 4174 32503 4183 32537
rect 4183 32503 4217 32537
rect 4217 32503 4226 32537
rect 4174 32494 4226 32503
rect 4334 32537 4386 32546
rect 4334 32503 4343 32537
rect 4343 32503 4377 32537
rect 4377 32503 4386 32537
rect 4334 32494 4386 32503
rect 4494 32537 4546 32546
rect 4494 32503 4503 32537
rect 4503 32503 4537 32537
rect 4537 32503 4546 32537
rect 4494 32494 4546 32503
rect 4654 32537 4706 32546
rect 4654 32503 4663 32537
rect 4663 32503 4697 32537
rect 4697 32503 4706 32537
rect 4654 32494 4706 32503
rect 4814 32537 4866 32546
rect 4814 32503 4823 32537
rect 4823 32503 4857 32537
rect 4857 32503 4866 32537
rect 4814 32494 4866 32503
rect 4974 32537 5026 32546
rect 4974 32503 4983 32537
rect 4983 32503 5017 32537
rect 5017 32503 5026 32537
rect 4974 32494 5026 32503
rect 5134 32537 5186 32546
rect 5134 32503 5143 32537
rect 5143 32503 5177 32537
rect 5177 32503 5186 32537
rect 5134 32494 5186 32503
rect 5294 32537 5346 32546
rect 5294 32503 5303 32537
rect 5303 32503 5337 32537
rect 5337 32503 5346 32537
rect 5294 32494 5346 32503
rect 5454 32537 5506 32546
rect 5454 32503 5463 32537
rect 5463 32503 5497 32537
rect 5497 32503 5506 32537
rect 5454 32494 5506 32503
rect 5614 32537 5666 32546
rect 5614 32503 5623 32537
rect 5623 32503 5657 32537
rect 5657 32503 5666 32537
rect 5614 32494 5666 32503
rect 5774 32537 5826 32546
rect 5774 32503 5783 32537
rect 5783 32503 5817 32537
rect 5817 32503 5826 32537
rect 5774 32494 5826 32503
rect 5934 32537 5986 32546
rect 5934 32503 5943 32537
rect 5943 32503 5977 32537
rect 5977 32503 5986 32537
rect 5934 32494 5986 32503
rect 6094 32537 6146 32546
rect 6094 32503 6103 32537
rect 6103 32503 6137 32537
rect 6137 32503 6146 32537
rect 6094 32494 6146 32503
rect 6254 32537 6306 32546
rect 6254 32503 6263 32537
rect 6263 32503 6297 32537
rect 6297 32503 6306 32537
rect 6254 32494 6306 32503
rect 6414 32537 6466 32546
rect 6414 32503 6423 32537
rect 6423 32503 6457 32537
rect 6457 32503 6466 32537
rect 6414 32494 6466 32503
rect 6574 32537 6626 32546
rect 6574 32503 6583 32537
rect 6583 32503 6617 32537
rect 6617 32503 6626 32537
rect 6574 32494 6626 32503
rect 6734 32537 6786 32546
rect 6734 32503 6743 32537
rect 6743 32503 6777 32537
rect 6777 32503 6786 32537
rect 6734 32494 6786 32503
rect 6894 32537 6946 32546
rect 6894 32503 6903 32537
rect 6903 32503 6937 32537
rect 6937 32503 6946 32537
rect 6894 32494 6946 32503
rect 7054 32537 7106 32546
rect 7054 32503 7063 32537
rect 7063 32503 7097 32537
rect 7097 32503 7106 32537
rect 7054 32494 7106 32503
rect 7214 32537 7266 32546
rect 7214 32503 7223 32537
rect 7223 32503 7257 32537
rect 7257 32503 7266 32537
rect 7214 32494 7266 32503
rect 7374 32537 7426 32546
rect 7374 32503 7383 32537
rect 7383 32503 7417 32537
rect 7417 32503 7426 32537
rect 7374 32494 7426 32503
rect 7534 32537 7586 32546
rect 7534 32503 7543 32537
rect 7543 32503 7577 32537
rect 7577 32503 7586 32537
rect 7534 32494 7586 32503
rect 7694 32537 7746 32546
rect 7694 32503 7703 32537
rect 7703 32503 7737 32537
rect 7737 32503 7746 32537
rect 7694 32494 7746 32503
rect 7854 32537 7906 32546
rect 7854 32503 7863 32537
rect 7863 32503 7897 32537
rect 7897 32503 7906 32537
rect 7854 32494 7906 32503
rect 8014 32537 8066 32546
rect 8014 32503 8023 32537
rect 8023 32503 8057 32537
rect 8057 32503 8066 32537
rect 8014 32494 8066 32503
rect 8174 32537 8226 32546
rect 8174 32503 8183 32537
rect 8183 32503 8217 32537
rect 8217 32503 8226 32537
rect 8174 32494 8226 32503
rect 8334 32537 8386 32546
rect 8334 32503 8343 32537
rect 8343 32503 8377 32537
rect 8377 32503 8386 32537
rect 8334 32494 8386 32503
rect 12494 32537 12546 32546
rect 12494 32503 12503 32537
rect 12503 32503 12537 32537
rect 12537 32503 12546 32537
rect 12494 32494 12546 32503
rect 12654 32537 12706 32546
rect 12654 32503 12663 32537
rect 12663 32503 12697 32537
rect 12697 32503 12706 32537
rect 12654 32494 12706 32503
rect 12814 32537 12866 32546
rect 12814 32503 12823 32537
rect 12823 32503 12857 32537
rect 12857 32503 12866 32537
rect 12814 32494 12866 32503
rect 12974 32537 13026 32546
rect 12974 32503 12983 32537
rect 12983 32503 13017 32537
rect 13017 32503 13026 32537
rect 12974 32494 13026 32503
rect 13134 32537 13186 32546
rect 13134 32503 13143 32537
rect 13143 32503 13177 32537
rect 13177 32503 13186 32537
rect 13134 32494 13186 32503
rect 13294 32537 13346 32546
rect 13294 32503 13303 32537
rect 13303 32503 13337 32537
rect 13337 32503 13346 32537
rect 13294 32494 13346 32503
rect 13454 32537 13506 32546
rect 13454 32503 13463 32537
rect 13463 32503 13497 32537
rect 13497 32503 13506 32537
rect 13454 32494 13506 32503
rect 13614 32537 13666 32546
rect 13614 32503 13623 32537
rect 13623 32503 13657 32537
rect 13657 32503 13666 32537
rect 13614 32494 13666 32503
rect 13774 32537 13826 32546
rect 13774 32503 13783 32537
rect 13783 32503 13817 32537
rect 13817 32503 13826 32537
rect 13774 32494 13826 32503
rect 13934 32537 13986 32546
rect 13934 32503 13943 32537
rect 13943 32503 13977 32537
rect 13977 32503 13986 32537
rect 13934 32494 13986 32503
rect 14094 32537 14146 32546
rect 14094 32503 14103 32537
rect 14103 32503 14137 32537
rect 14137 32503 14146 32537
rect 14094 32494 14146 32503
rect 14254 32537 14306 32546
rect 14254 32503 14263 32537
rect 14263 32503 14297 32537
rect 14297 32503 14306 32537
rect 14254 32494 14306 32503
rect 14414 32537 14466 32546
rect 14414 32503 14423 32537
rect 14423 32503 14457 32537
rect 14457 32503 14466 32537
rect 14414 32494 14466 32503
rect 14574 32537 14626 32546
rect 14574 32503 14583 32537
rect 14583 32503 14617 32537
rect 14617 32503 14626 32537
rect 14574 32494 14626 32503
rect 14734 32537 14786 32546
rect 14734 32503 14743 32537
rect 14743 32503 14777 32537
rect 14777 32503 14786 32537
rect 14734 32494 14786 32503
rect 14894 32537 14946 32546
rect 14894 32503 14903 32537
rect 14903 32503 14937 32537
rect 14937 32503 14946 32537
rect 14894 32494 14946 32503
rect 15054 32537 15106 32546
rect 15054 32503 15063 32537
rect 15063 32503 15097 32537
rect 15097 32503 15106 32537
rect 15054 32494 15106 32503
rect 15214 32537 15266 32546
rect 15214 32503 15223 32537
rect 15223 32503 15257 32537
rect 15257 32503 15266 32537
rect 15214 32494 15266 32503
rect 15374 32537 15426 32546
rect 15374 32503 15383 32537
rect 15383 32503 15417 32537
rect 15417 32503 15426 32537
rect 15374 32494 15426 32503
rect 15534 32537 15586 32546
rect 15534 32503 15543 32537
rect 15543 32503 15577 32537
rect 15577 32503 15586 32537
rect 15534 32494 15586 32503
rect 15694 32537 15746 32546
rect 15694 32503 15703 32537
rect 15703 32503 15737 32537
rect 15737 32503 15746 32537
rect 15694 32494 15746 32503
rect 15854 32537 15906 32546
rect 15854 32503 15863 32537
rect 15863 32503 15897 32537
rect 15897 32503 15906 32537
rect 15854 32494 15906 32503
rect 16014 32537 16066 32546
rect 16014 32503 16023 32537
rect 16023 32503 16057 32537
rect 16057 32503 16066 32537
rect 16014 32494 16066 32503
rect 16174 32537 16226 32546
rect 16174 32503 16183 32537
rect 16183 32503 16217 32537
rect 16217 32503 16226 32537
rect 16174 32494 16226 32503
rect 16334 32537 16386 32546
rect 16334 32503 16343 32537
rect 16343 32503 16377 32537
rect 16377 32503 16386 32537
rect 16334 32494 16386 32503
rect 16494 32537 16546 32546
rect 16494 32503 16503 32537
rect 16503 32503 16537 32537
rect 16537 32503 16546 32537
rect 16494 32494 16546 32503
rect 16654 32537 16706 32546
rect 16654 32503 16663 32537
rect 16663 32503 16697 32537
rect 16697 32503 16706 32537
rect 16654 32494 16706 32503
rect 16814 32537 16866 32546
rect 16814 32503 16823 32537
rect 16823 32503 16857 32537
rect 16857 32503 16866 32537
rect 16814 32494 16866 32503
rect 16974 32537 17026 32546
rect 16974 32503 16983 32537
rect 16983 32503 17017 32537
rect 17017 32503 17026 32537
rect 16974 32494 17026 32503
rect 17134 32537 17186 32546
rect 17134 32503 17143 32537
rect 17143 32503 17177 32537
rect 17177 32503 17186 32537
rect 17134 32494 17186 32503
rect 17294 32537 17346 32546
rect 17294 32503 17303 32537
rect 17303 32503 17337 32537
rect 17337 32503 17346 32537
rect 17294 32494 17346 32503
rect 17454 32537 17506 32546
rect 17454 32503 17463 32537
rect 17463 32503 17497 32537
rect 17497 32503 17506 32537
rect 17454 32494 17506 32503
rect 17614 32537 17666 32546
rect 17614 32503 17623 32537
rect 17623 32503 17657 32537
rect 17657 32503 17666 32537
rect 17614 32494 17666 32503
rect 17774 32537 17826 32546
rect 17774 32503 17783 32537
rect 17783 32503 17817 32537
rect 17817 32503 17826 32537
rect 17774 32494 17826 32503
rect 17934 32537 17986 32546
rect 17934 32503 17943 32537
rect 17943 32503 17977 32537
rect 17977 32503 17986 32537
rect 17934 32494 17986 32503
rect 18094 32537 18146 32546
rect 18094 32503 18103 32537
rect 18103 32503 18137 32537
rect 18137 32503 18146 32537
rect 18094 32494 18146 32503
rect 18254 32537 18306 32546
rect 18254 32503 18263 32537
rect 18263 32503 18297 32537
rect 18297 32503 18306 32537
rect 18254 32494 18306 32503
rect 18414 32537 18466 32546
rect 18414 32503 18423 32537
rect 18423 32503 18457 32537
rect 18457 32503 18466 32537
rect 18414 32494 18466 32503
rect 18574 32537 18626 32546
rect 18574 32503 18583 32537
rect 18583 32503 18617 32537
rect 18617 32503 18626 32537
rect 18574 32494 18626 32503
rect 18734 32537 18786 32546
rect 18734 32503 18743 32537
rect 18743 32503 18777 32537
rect 18777 32503 18786 32537
rect 18734 32494 18786 32503
rect 18894 32537 18946 32546
rect 18894 32503 18903 32537
rect 18903 32503 18937 32537
rect 18937 32503 18946 32537
rect 18894 32494 18946 32503
rect 23134 32537 23186 32546
rect 23134 32503 23143 32537
rect 23143 32503 23177 32537
rect 23177 32503 23186 32537
rect 23134 32494 23186 32503
rect 23294 32537 23346 32546
rect 23294 32503 23303 32537
rect 23303 32503 23337 32537
rect 23337 32503 23346 32537
rect 23294 32494 23346 32503
rect 23454 32537 23506 32546
rect 23454 32503 23463 32537
rect 23463 32503 23497 32537
rect 23497 32503 23506 32537
rect 23454 32494 23506 32503
rect 23614 32537 23666 32546
rect 23614 32503 23623 32537
rect 23623 32503 23657 32537
rect 23657 32503 23666 32537
rect 23614 32494 23666 32503
rect 23774 32537 23826 32546
rect 23774 32503 23783 32537
rect 23783 32503 23817 32537
rect 23817 32503 23826 32537
rect 23774 32494 23826 32503
rect 23934 32537 23986 32546
rect 23934 32503 23943 32537
rect 23943 32503 23977 32537
rect 23977 32503 23986 32537
rect 23934 32494 23986 32503
rect 24094 32537 24146 32546
rect 24094 32503 24103 32537
rect 24103 32503 24137 32537
rect 24137 32503 24146 32537
rect 24094 32494 24146 32503
rect 24254 32537 24306 32546
rect 24254 32503 24263 32537
rect 24263 32503 24297 32537
rect 24297 32503 24306 32537
rect 24254 32494 24306 32503
rect 24414 32537 24466 32546
rect 24414 32503 24423 32537
rect 24423 32503 24457 32537
rect 24457 32503 24466 32537
rect 24414 32494 24466 32503
rect 24574 32537 24626 32546
rect 24574 32503 24583 32537
rect 24583 32503 24617 32537
rect 24617 32503 24626 32537
rect 24574 32494 24626 32503
rect 24734 32537 24786 32546
rect 24734 32503 24743 32537
rect 24743 32503 24777 32537
rect 24777 32503 24786 32537
rect 24734 32494 24786 32503
rect 24894 32537 24946 32546
rect 24894 32503 24903 32537
rect 24903 32503 24937 32537
rect 24937 32503 24946 32537
rect 24894 32494 24946 32503
rect 25054 32537 25106 32546
rect 25054 32503 25063 32537
rect 25063 32503 25097 32537
rect 25097 32503 25106 32537
rect 25054 32494 25106 32503
rect 25214 32537 25266 32546
rect 25214 32503 25223 32537
rect 25223 32503 25257 32537
rect 25257 32503 25266 32537
rect 25214 32494 25266 32503
rect 25374 32537 25426 32546
rect 25374 32503 25383 32537
rect 25383 32503 25417 32537
rect 25417 32503 25426 32537
rect 25374 32494 25426 32503
rect 25534 32537 25586 32546
rect 25534 32503 25543 32537
rect 25543 32503 25577 32537
rect 25577 32503 25586 32537
rect 25534 32494 25586 32503
rect 25694 32537 25746 32546
rect 25694 32503 25703 32537
rect 25703 32503 25737 32537
rect 25737 32503 25746 32537
rect 25694 32494 25746 32503
rect 25854 32537 25906 32546
rect 25854 32503 25863 32537
rect 25863 32503 25897 32537
rect 25897 32503 25906 32537
rect 25854 32494 25906 32503
rect 26014 32537 26066 32546
rect 26014 32503 26023 32537
rect 26023 32503 26057 32537
rect 26057 32503 26066 32537
rect 26014 32494 26066 32503
rect 26174 32537 26226 32546
rect 26174 32503 26183 32537
rect 26183 32503 26217 32537
rect 26217 32503 26226 32537
rect 26174 32494 26226 32503
rect 26334 32537 26386 32546
rect 26334 32503 26343 32537
rect 26343 32503 26377 32537
rect 26377 32503 26386 32537
rect 26334 32494 26386 32503
rect 26494 32537 26546 32546
rect 26494 32503 26503 32537
rect 26503 32503 26537 32537
rect 26537 32503 26546 32537
rect 26494 32494 26546 32503
rect 26654 32537 26706 32546
rect 26654 32503 26663 32537
rect 26663 32503 26697 32537
rect 26697 32503 26706 32537
rect 26654 32494 26706 32503
rect 26814 32537 26866 32546
rect 26814 32503 26823 32537
rect 26823 32503 26857 32537
rect 26857 32503 26866 32537
rect 26814 32494 26866 32503
rect 26974 32537 27026 32546
rect 26974 32503 26983 32537
rect 26983 32503 27017 32537
rect 27017 32503 27026 32537
rect 26974 32494 27026 32503
rect 27134 32537 27186 32546
rect 27134 32503 27143 32537
rect 27143 32503 27177 32537
rect 27177 32503 27186 32537
rect 27134 32494 27186 32503
rect 27294 32537 27346 32546
rect 27294 32503 27303 32537
rect 27303 32503 27337 32537
rect 27337 32503 27346 32537
rect 27294 32494 27346 32503
rect 27454 32537 27506 32546
rect 27454 32503 27463 32537
rect 27463 32503 27497 32537
rect 27497 32503 27506 32537
rect 27454 32494 27506 32503
rect 27614 32537 27666 32546
rect 27614 32503 27623 32537
rect 27623 32503 27657 32537
rect 27657 32503 27666 32537
rect 27614 32494 27666 32503
rect 27774 32537 27826 32546
rect 27774 32503 27783 32537
rect 27783 32503 27817 32537
rect 27817 32503 27826 32537
rect 27774 32494 27826 32503
rect 27934 32537 27986 32546
rect 27934 32503 27943 32537
rect 27943 32503 27977 32537
rect 27977 32503 27986 32537
rect 27934 32494 27986 32503
rect 28094 32537 28146 32546
rect 28094 32503 28103 32537
rect 28103 32503 28137 32537
rect 28137 32503 28146 32537
rect 28094 32494 28146 32503
rect 28254 32537 28306 32546
rect 28254 32503 28263 32537
rect 28263 32503 28297 32537
rect 28297 32503 28306 32537
rect 28254 32494 28306 32503
rect 28414 32537 28466 32546
rect 28414 32503 28423 32537
rect 28423 32503 28457 32537
rect 28457 32503 28466 32537
rect 28414 32494 28466 32503
rect 28574 32537 28626 32546
rect 28574 32503 28583 32537
rect 28583 32503 28617 32537
rect 28617 32503 28626 32537
rect 28574 32494 28626 32503
rect 28734 32537 28786 32546
rect 28734 32503 28743 32537
rect 28743 32503 28777 32537
rect 28777 32503 28786 32537
rect 28734 32494 28786 32503
rect 28894 32537 28946 32546
rect 28894 32503 28903 32537
rect 28903 32503 28937 32537
rect 28937 32503 28946 32537
rect 28894 32494 28946 32503
rect 29054 32537 29106 32546
rect 29054 32503 29063 32537
rect 29063 32503 29097 32537
rect 29097 32503 29106 32537
rect 29054 32494 29106 32503
rect 29214 32537 29266 32546
rect 29214 32503 29223 32537
rect 29223 32503 29257 32537
rect 29257 32503 29266 32537
rect 29214 32494 29266 32503
rect 29374 32537 29426 32546
rect 29374 32503 29383 32537
rect 29383 32503 29417 32537
rect 29417 32503 29426 32537
rect 29374 32494 29426 32503
rect 33534 32537 33586 32546
rect 33534 32503 33543 32537
rect 33543 32503 33577 32537
rect 33577 32503 33586 32537
rect 33534 32494 33586 32503
rect 33694 32537 33746 32546
rect 33694 32503 33703 32537
rect 33703 32503 33737 32537
rect 33737 32503 33746 32537
rect 33694 32494 33746 32503
rect 33854 32537 33906 32546
rect 33854 32503 33863 32537
rect 33863 32503 33897 32537
rect 33897 32503 33906 32537
rect 33854 32494 33906 32503
rect 34014 32537 34066 32546
rect 34014 32503 34023 32537
rect 34023 32503 34057 32537
rect 34057 32503 34066 32537
rect 34014 32494 34066 32503
rect 34174 32537 34226 32546
rect 34174 32503 34183 32537
rect 34183 32503 34217 32537
rect 34217 32503 34226 32537
rect 34174 32494 34226 32503
rect 34334 32537 34386 32546
rect 34334 32503 34343 32537
rect 34343 32503 34377 32537
rect 34377 32503 34386 32537
rect 34334 32494 34386 32503
rect 34494 32537 34546 32546
rect 34494 32503 34503 32537
rect 34503 32503 34537 32537
rect 34537 32503 34546 32537
rect 34494 32494 34546 32503
rect 34654 32537 34706 32546
rect 34654 32503 34663 32537
rect 34663 32503 34697 32537
rect 34697 32503 34706 32537
rect 34654 32494 34706 32503
rect 34814 32537 34866 32546
rect 34814 32503 34823 32537
rect 34823 32503 34857 32537
rect 34857 32503 34866 32537
rect 34814 32494 34866 32503
rect 34974 32537 35026 32546
rect 34974 32503 34983 32537
rect 34983 32503 35017 32537
rect 35017 32503 35026 32537
rect 34974 32494 35026 32503
rect 35134 32537 35186 32546
rect 35134 32503 35143 32537
rect 35143 32503 35177 32537
rect 35177 32503 35186 32537
rect 35134 32494 35186 32503
rect 35294 32537 35346 32546
rect 35294 32503 35303 32537
rect 35303 32503 35337 32537
rect 35337 32503 35346 32537
rect 35294 32494 35346 32503
rect 35454 32537 35506 32546
rect 35454 32503 35463 32537
rect 35463 32503 35497 32537
rect 35497 32503 35506 32537
rect 35454 32494 35506 32503
rect 35614 32537 35666 32546
rect 35614 32503 35623 32537
rect 35623 32503 35657 32537
rect 35657 32503 35666 32537
rect 35614 32494 35666 32503
rect 35774 32537 35826 32546
rect 35774 32503 35783 32537
rect 35783 32503 35817 32537
rect 35817 32503 35826 32537
rect 35774 32494 35826 32503
rect 35934 32537 35986 32546
rect 35934 32503 35943 32537
rect 35943 32503 35977 32537
rect 35977 32503 35986 32537
rect 35934 32494 35986 32503
rect 36094 32537 36146 32546
rect 36094 32503 36103 32537
rect 36103 32503 36137 32537
rect 36137 32503 36146 32537
rect 36094 32494 36146 32503
rect 36254 32537 36306 32546
rect 36254 32503 36263 32537
rect 36263 32503 36297 32537
rect 36297 32503 36306 32537
rect 36254 32494 36306 32503
rect 36414 32537 36466 32546
rect 36414 32503 36423 32537
rect 36423 32503 36457 32537
rect 36457 32503 36466 32537
rect 36414 32494 36466 32503
rect 36574 32537 36626 32546
rect 36574 32503 36583 32537
rect 36583 32503 36617 32537
rect 36617 32503 36626 32537
rect 36574 32494 36626 32503
rect 36734 32537 36786 32546
rect 36734 32503 36743 32537
rect 36743 32503 36777 32537
rect 36777 32503 36786 32537
rect 36734 32494 36786 32503
rect 36894 32537 36946 32546
rect 36894 32503 36903 32537
rect 36903 32503 36937 32537
rect 36937 32503 36946 32537
rect 36894 32494 36946 32503
rect 37054 32537 37106 32546
rect 37054 32503 37063 32537
rect 37063 32503 37097 32537
rect 37097 32503 37106 32537
rect 37054 32494 37106 32503
rect 37214 32537 37266 32546
rect 37214 32503 37223 32537
rect 37223 32503 37257 32537
rect 37257 32503 37266 32537
rect 37214 32494 37266 32503
rect 37374 32537 37426 32546
rect 37374 32503 37383 32537
rect 37383 32503 37417 32537
rect 37417 32503 37426 32537
rect 37374 32494 37426 32503
rect 37534 32537 37586 32546
rect 37534 32503 37543 32537
rect 37543 32503 37577 32537
rect 37577 32503 37586 32537
rect 37534 32494 37586 32503
rect 37694 32537 37746 32546
rect 37694 32503 37703 32537
rect 37703 32503 37737 32537
rect 37737 32503 37746 32537
rect 37694 32494 37746 32503
rect 37854 32537 37906 32546
rect 37854 32503 37863 32537
rect 37863 32503 37897 32537
rect 37897 32503 37906 32537
rect 37854 32494 37906 32503
rect 38014 32537 38066 32546
rect 38014 32503 38023 32537
rect 38023 32503 38057 32537
rect 38057 32503 38066 32537
rect 38014 32494 38066 32503
rect 38174 32537 38226 32546
rect 38174 32503 38183 32537
rect 38183 32503 38217 32537
rect 38217 32503 38226 32537
rect 38174 32494 38226 32503
rect 38334 32537 38386 32546
rect 38334 32503 38343 32537
rect 38343 32503 38377 32537
rect 38377 32503 38386 32537
rect 38334 32494 38386 32503
rect 38494 32537 38546 32546
rect 38494 32503 38503 32537
rect 38503 32503 38537 32537
rect 38537 32503 38546 32537
rect 38494 32494 38546 32503
rect 38654 32537 38706 32546
rect 38654 32503 38663 32537
rect 38663 32503 38697 32537
rect 38697 32503 38706 32537
rect 38654 32494 38706 32503
rect 38814 32537 38866 32546
rect 38814 32503 38823 32537
rect 38823 32503 38857 32537
rect 38857 32503 38866 32537
rect 38814 32494 38866 32503
rect 38974 32537 39026 32546
rect 38974 32503 38983 32537
rect 38983 32503 39017 32537
rect 39017 32503 39026 32537
rect 38974 32494 39026 32503
rect 39134 32537 39186 32546
rect 39134 32503 39143 32537
rect 39143 32503 39177 32537
rect 39177 32503 39186 32537
rect 39134 32494 39186 32503
rect 39294 32537 39346 32546
rect 39294 32503 39303 32537
rect 39303 32503 39337 32537
rect 39337 32503 39346 32537
rect 39294 32494 39346 32503
rect 39454 32537 39506 32546
rect 39454 32503 39463 32537
rect 39463 32503 39497 32537
rect 39497 32503 39506 32537
rect 39454 32494 39506 32503
rect 39614 32537 39666 32546
rect 39614 32503 39623 32537
rect 39623 32503 39657 32537
rect 39657 32503 39666 32537
rect 39614 32494 39666 32503
rect 39774 32537 39826 32546
rect 39774 32503 39783 32537
rect 39783 32503 39817 32537
rect 39817 32503 39826 32537
rect 39774 32494 39826 32503
rect 39934 32537 39986 32546
rect 39934 32503 39943 32537
rect 39943 32503 39977 32537
rect 39977 32503 39986 32537
rect 39934 32494 39986 32503
rect 40094 32537 40146 32546
rect 40094 32503 40103 32537
rect 40103 32503 40137 32537
rect 40137 32503 40146 32537
rect 40094 32494 40146 32503
rect 40254 32537 40306 32546
rect 40254 32503 40263 32537
rect 40263 32503 40297 32537
rect 40297 32503 40306 32537
rect 40254 32494 40306 32503
rect 40414 32537 40466 32546
rect 40414 32503 40423 32537
rect 40423 32503 40457 32537
rect 40457 32503 40466 32537
rect 40414 32494 40466 32503
rect 40574 32537 40626 32546
rect 40574 32503 40583 32537
rect 40583 32503 40617 32537
rect 40617 32503 40626 32537
rect 40574 32494 40626 32503
rect 40734 32537 40786 32546
rect 40734 32503 40743 32537
rect 40743 32503 40777 32537
rect 40777 32503 40786 32537
rect 40734 32494 40786 32503
rect 40894 32537 40946 32546
rect 40894 32503 40903 32537
rect 40903 32503 40937 32537
rect 40937 32503 40946 32537
rect 40894 32494 40946 32503
rect 41054 32537 41106 32546
rect 41054 32503 41063 32537
rect 41063 32503 41097 32537
rect 41097 32503 41106 32537
rect 41054 32494 41106 32503
rect 41214 32537 41266 32546
rect 41214 32503 41223 32537
rect 41223 32503 41257 32537
rect 41257 32503 41266 32537
rect 41214 32494 41266 32503
rect 41374 32537 41426 32546
rect 41374 32503 41383 32537
rect 41383 32503 41417 32537
rect 41417 32503 41426 32537
rect 41374 32494 41426 32503
rect 41534 32537 41586 32546
rect 41534 32503 41543 32537
rect 41543 32503 41577 32537
rect 41577 32503 41586 32537
rect 41534 32494 41586 32503
rect 41694 32537 41746 32546
rect 41694 32503 41703 32537
rect 41703 32503 41737 32537
rect 41737 32503 41746 32537
rect 41694 32494 41746 32503
rect 41854 32537 41906 32546
rect 41854 32503 41863 32537
rect 41863 32503 41897 32537
rect 41897 32503 41906 32537
rect 41854 32494 41906 32503
rect 14 32377 66 32386
rect 14 32343 23 32377
rect 23 32343 57 32377
rect 57 32343 66 32377
rect 14 32334 66 32343
rect 174 32377 226 32386
rect 174 32343 183 32377
rect 183 32343 217 32377
rect 217 32343 226 32377
rect 174 32334 226 32343
rect 334 32377 386 32386
rect 334 32343 343 32377
rect 343 32343 377 32377
rect 377 32343 386 32377
rect 334 32334 386 32343
rect 494 32377 546 32386
rect 494 32343 503 32377
rect 503 32343 537 32377
rect 537 32343 546 32377
rect 494 32334 546 32343
rect 654 32377 706 32386
rect 654 32343 663 32377
rect 663 32343 697 32377
rect 697 32343 706 32377
rect 654 32334 706 32343
rect 814 32377 866 32386
rect 814 32343 823 32377
rect 823 32343 857 32377
rect 857 32343 866 32377
rect 814 32334 866 32343
rect 974 32377 1026 32386
rect 974 32343 983 32377
rect 983 32343 1017 32377
rect 1017 32343 1026 32377
rect 974 32334 1026 32343
rect 1134 32377 1186 32386
rect 1134 32343 1143 32377
rect 1143 32343 1177 32377
rect 1177 32343 1186 32377
rect 1134 32334 1186 32343
rect 1294 32377 1346 32386
rect 1294 32343 1303 32377
rect 1303 32343 1337 32377
rect 1337 32343 1346 32377
rect 1294 32334 1346 32343
rect 1454 32377 1506 32386
rect 1454 32343 1463 32377
rect 1463 32343 1497 32377
rect 1497 32343 1506 32377
rect 1454 32334 1506 32343
rect 1614 32377 1666 32386
rect 1614 32343 1623 32377
rect 1623 32343 1657 32377
rect 1657 32343 1666 32377
rect 1614 32334 1666 32343
rect 1774 32377 1826 32386
rect 1774 32343 1783 32377
rect 1783 32343 1817 32377
rect 1817 32343 1826 32377
rect 1774 32334 1826 32343
rect 1934 32377 1986 32386
rect 1934 32343 1943 32377
rect 1943 32343 1977 32377
rect 1977 32343 1986 32377
rect 1934 32334 1986 32343
rect 2094 32377 2146 32386
rect 2094 32343 2103 32377
rect 2103 32343 2137 32377
rect 2137 32343 2146 32377
rect 2094 32334 2146 32343
rect 2254 32377 2306 32386
rect 2254 32343 2263 32377
rect 2263 32343 2297 32377
rect 2297 32343 2306 32377
rect 2254 32334 2306 32343
rect 2414 32377 2466 32386
rect 2414 32343 2423 32377
rect 2423 32343 2457 32377
rect 2457 32343 2466 32377
rect 2414 32334 2466 32343
rect 2574 32377 2626 32386
rect 2574 32343 2583 32377
rect 2583 32343 2617 32377
rect 2617 32343 2626 32377
rect 2574 32334 2626 32343
rect 2734 32377 2786 32386
rect 2734 32343 2743 32377
rect 2743 32343 2777 32377
rect 2777 32343 2786 32377
rect 2734 32334 2786 32343
rect 2894 32377 2946 32386
rect 2894 32343 2903 32377
rect 2903 32343 2937 32377
rect 2937 32343 2946 32377
rect 2894 32334 2946 32343
rect 3054 32377 3106 32386
rect 3054 32343 3063 32377
rect 3063 32343 3097 32377
rect 3097 32343 3106 32377
rect 3054 32334 3106 32343
rect 3214 32377 3266 32386
rect 3214 32343 3223 32377
rect 3223 32343 3257 32377
rect 3257 32343 3266 32377
rect 3214 32334 3266 32343
rect 3374 32377 3426 32386
rect 3374 32343 3383 32377
rect 3383 32343 3417 32377
rect 3417 32343 3426 32377
rect 3374 32334 3426 32343
rect 3534 32377 3586 32386
rect 3534 32343 3543 32377
rect 3543 32343 3577 32377
rect 3577 32343 3586 32377
rect 3534 32334 3586 32343
rect 3694 32377 3746 32386
rect 3694 32343 3703 32377
rect 3703 32343 3737 32377
rect 3737 32343 3746 32377
rect 3694 32334 3746 32343
rect 3854 32377 3906 32386
rect 3854 32343 3863 32377
rect 3863 32343 3897 32377
rect 3897 32343 3906 32377
rect 3854 32334 3906 32343
rect 4014 32377 4066 32386
rect 4014 32343 4023 32377
rect 4023 32343 4057 32377
rect 4057 32343 4066 32377
rect 4014 32334 4066 32343
rect 4174 32377 4226 32386
rect 4174 32343 4183 32377
rect 4183 32343 4217 32377
rect 4217 32343 4226 32377
rect 4174 32334 4226 32343
rect 4334 32377 4386 32386
rect 4334 32343 4343 32377
rect 4343 32343 4377 32377
rect 4377 32343 4386 32377
rect 4334 32334 4386 32343
rect 4494 32377 4546 32386
rect 4494 32343 4503 32377
rect 4503 32343 4537 32377
rect 4537 32343 4546 32377
rect 4494 32334 4546 32343
rect 4654 32377 4706 32386
rect 4654 32343 4663 32377
rect 4663 32343 4697 32377
rect 4697 32343 4706 32377
rect 4654 32334 4706 32343
rect 4814 32377 4866 32386
rect 4814 32343 4823 32377
rect 4823 32343 4857 32377
rect 4857 32343 4866 32377
rect 4814 32334 4866 32343
rect 4974 32377 5026 32386
rect 4974 32343 4983 32377
rect 4983 32343 5017 32377
rect 5017 32343 5026 32377
rect 4974 32334 5026 32343
rect 5134 32377 5186 32386
rect 5134 32343 5143 32377
rect 5143 32343 5177 32377
rect 5177 32343 5186 32377
rect 5134 32334 5186 32343
rect 5294 32377 5346 32386
rect 5294 32343 5303 32377
rect 5303 32343 5337 32377
rect 5337 32343 5346 32377
rect 5294 32334 5346 32343
rect 5454 32377 5506 32386
rect 5454 32343 5463 32377
rect 5463 32343 5497 32377
rect 5497 32343 5506 32377
rect 5454 32334 5506 32343
rect 5614 32377 5666 32386
rect 5614 32343 5623 32377
rect 5623 32343 5657 32377
rect 5657 32343 5666 32377
rect 5614 32334 5666 32343
rect 5774 32377 5826 32386
rect 5774 32343 5783 32377
rect 5783 32343 5817 32377
rect 5817 32343 5826 32377
rect 5774 32334 5826 32343
rect 5934 32377 5986 32386
rect 5934 32343 5943 32377
rect 5943 32343 5977 32377
rect 5977 32343 5986 32377
rect 5934 32334 5986 32343
rect 6094 32377 6146 32386
rect 6094 32343 6103 32377
rect 6103 32343 6137 32377
rect 6137 32343 6146 32377
rect 6094 32334 6146 32343
rect 6254 32377 6306 32386
rect 6254 32343 6263 32377
rect 6263 32343 6297 32377
rect 6297 32343 6306 32377
rect 6254 32334 6306 32343
rect 6414 32377 6466 32386
rect 6414 32343 6423 32377
rect 6423 32343 6457 32377
rect 6457 32343 6466 32377
rect 6414 32334 6466 32343
rect 6574 32377 6626 32386
rect 6574 32343 6583 32377
rect 6583 32343 6617 32377
rect 6617 32343 6626 32377
rect 6574 32334 6626 32343
rect 6734 32377 6786 32386
rect 6734 32343 6743 32377
rect 6743 32343 6777 32377
rect 6777 32343 6786 32377
rect 6734 32334 6786 32343
rect 6894 32377 6946 32386
rect 6894 32343 6903 32377
rect 6903 32343 6937 32377
rect 6937 32343 6946 32377
rect 6894 32334 6946 32343
rect 7054 32377 7106 32386
rect 7054 32343 7063 32377
rect 7063 32343 7097 32377
rect 7097 32343 7106 32377
rect 7054 32334 7106 32343
rect 7214 32377 7266 32386
rect 7214 32343 7223 32377
rect 7223 32343 7257 32377
rect 7257 32343 7266 32377
rect 7214 32334 7266 32343
rect 7374 32377 7426 32386
rect 7374 32343 7383 32377
rect 7383 32343 7417 32377
rect 7417 32343 7426 32377
rect 7374 32334 7426 32343
rect 7534 32377 7586 32386
rect 7534 32343 7543 32377
rect 7543 32343 7577 32377
rect 7577 32343 7586 32377
rect 7534 32334 7586 32343
rect 7694 32377 7746 32386
rect 7694 32343 7703 32377
rect 7703 32343 7737 32377
rect 7737 32343 7746 32377
rect 7694 32334 7746 32343
rect 7854 32377 7906 32386
rect 7854 32343 7863 32377
rect 7863 32343 7897 32377
rect 7897 32343 7906 32377
rect 7854 32334 7906 32343
rect 8014 32377 8066 32386
rect 8014 32343 8023 32377
rect 8023 32343 8057 32377
rect 8057 32343 8066 32377
rect 8014 32334 8066 32343
rect 8174 32377 8226 32386
rect 8174 32343 8183 32377
rect 8183 32343 8217 32377
rect 8217 32343 8226 32377
rect 8174 32334 8226 32343
rect 8334 32377 8386 32386
rect 8334 32343 8343 32377
rect 8343 32343 8377 32377
rect 8377 32343 8386 32377
rect 8334 32334 8386 32343
rect 12494 32377 12546 32386
rect 12494 32343 12503 32377
rect 12503 32343 12537 32377
rect 12537 32343 12546 32377
rect 12494 32334 12546 32343
rect 12654 32377 12706 32386
rect 12654 32343 12663 32377
rect 12663 32343 12697 32377
rect 12697 32343 12706 32377
rect 12654 32334 12706 32343
rect 12814 32377 12866 32386
rect 12814 32343 12823 32377
rect 12823 32343 12857 32377
rect 12857 32343 12866 32377
rect 12814 32334 12866 32343
rect 12974 32377 13026 32386
rect 12974 32343 12983 32377
rect 12983 32343 13017 32377
rect 13017 32343 13026 32377
rect 12974 32334 13026 32343
rect 13134 32377 13186 32386
rect 13134 32343 13143 32377
rect 13143 32343 13177 32377
rect 13177 32343 13186 32377
rect 13134 32334 13186 32343
rect 13294 32377 13346 32386
rect 13294 32343 13303 32377
rect 13303 32343 13337 32377
rect 13337 32343 13346 32377
rect 13294 32334 13346 32343
rect 13454 32377 13506 32386
rect 13454 32343 13463 32377
rect 13463 32343 13497 32377
rect 13497 32343 13506 32377
rect 13454 32334 13506 32343
rect 13614 32377 13666 32386
rect 13614 32343 13623 32377
rect 13623 32343 13657 32377
rect 13657 32343 13666 32377
rect 13614 32334 13666 32343
rect 13774 32377 13826 32386
rect 13774 32343 13783 32377
rect 13783 32343 13817 32377
rect 13817 32343 13826 32377
rect 13774 32334 13826 32343
rect 13934 32377 13986 32386
rect 13934 32343 13943 32377
rect 13943 32343 13977 32377
rect 13977 32343 13986 32377
rect 13934 32334 13986 32343
rect 14094 32377 14146 32386
rect 14094 32343 14103 32377
rect 14103 32343 14137 32377
rect 14137 32343 14146 32377
rect 14094 32334 14146 32343
rect 14254 32377 14306 32386
rect 14254 32343 14263 32377
rect 14263 32343 14297 32377
rect 14297 32343 14306 32377
rect 14254 32334 14306 32343
rect 14414 32377 14466 32386
rect 14414 32343 14423 32377
rect 14423 32343 14457 32377
rect 14457 32343 14466 32377
rect 14414 32334 14466 32343
rect 14574 32377 14626 32386
rect 14574 32343 14583 32377
rect 14583 32343 14617 32377
rect 14617 32343 14626 32377
rect 14574 32334 14626 32343
rect 14734 32377 14786 32386
rect 14734 32343 14743 32377
rect 14743 32343 14777 32377
rect 14777 32343 14786 32377
rect 14734 32334 14786 32343
rect 14894 32377 14946 32386
rect 14894 32343 14903 32377
rect 14903 32343 14937 32377
rect 14937 32343 14946 32377
rect 14894 32334 14946 32343
rect 15054 32377 15106 32386
rect 15054 32343 15063 32377
rect 15063 32343 15097 32377
rect 15097 32343 15106 32377
rect 15054 32334 15106 32343
rect 15214 32377 15266 32386
rect 15214 32343 15223 32377
rect 15223 32343 15257 32377
rect 15257 32343 15266 32377
rect 15214 32334 15266 32343
rect 15374 32377 15426 32386
rect 15374 32343 15383 32377
rect 15383 32343 15417 32377
rect 15417 32343 15426 32377
rect 15374 32334 15426 32343
rect 15534 32377 15586 32386
rect 15534 32343 15543 32377
rect 15543 32343 15577 32377
rect 15577 32343 15586 32377
rect 15534 32334 15586 32343
rect 15694 32377 15746 32386
rect 15694 32343 15703 32377
rect 15703 32343 15737 32377
rect 15737 32343 15746 32377
rect 15694 32334 15746 32343
rect 15854 32377 15906 32386
rect 15854 32343 15863 32377
rect 15863 32343 15897 32377
rect 15897 32343 15906 32377
rect 15854 32334 15906 32343
rect 16014 32377 16066 32386
rect 16014 32343 16023 32377
rect 16023 32343 16057 32377
rect 16057 32343 16066 32377
rect 16014 32334 16066 32343
rect 16174 32377 16226 32386
rect 16174 32343 16183 32377
rect 16183 32343 16217 32377
rect 16217 32343 16226 32377
rect 16174 32334 16226 32343
rect 16334 32377 16386 32386
rect 16334 32343 16343 32377
rect 16343 32343 16377 32377
rect 16377 32343 16386 32377
rect 16334 32334 16386 32343
rect 16494 32377 16546 32386
rect 16494 32343 16503 32377
rect 16503 32343 16537 32377
rect 16537 32343 16546 32377
rect 16494 32334 16546 32343
rect 16654 32377 16706 32386
rect 16654 32343 16663 32377
rect 16663 32343 16697 32377
rect 16697 32343 16706 32377
rect 16654 32334 16706 32343
rect 16814 32377 16866 32386
rect 16814 32343 16823 32377
rect 16823 32343 16857 32377
rect 16857 32343 16866 32377
rect 16814 32334 16866 32343
rect 16974 32377 17026 32386
rect 16974 32343 16983 32377
rect 16983 32343 17017 32377
rect 17017 32343 17026 32377
rect 16974 32334 17026 32343
rect 17134 32377 17186 32386
rect 17134 32343 17143 32377
rect 17143 32343 17177 32377
rect 17177 32343 17186 32377
rect 17134 32334 17186 32343
rect 17294 32377 17346 32386
rect 17294 32343 17303 32377
rect 17303 32343 17337 32377
rect 17337 32343 17346 32377
rect 17294 32334 17346 32343
rect 17454 32377 17506 32386
rect 17454 32343 17463 32377
rect 17463 32343 17497 32377
rect 17497 32343 17506 32377
rect 17454 32334 17506 32343
rect 17614 32377 17666 32386
rect 17614 32343 17623 32377
rect 17623 32343 17657 32377
rect 17657 32343 17666 32377
rect 17614 32334 17666 32343
rect 17774 32377 17826 32386
rect 17774 32343 17783 32377
rect 17783 32343 17817 32377
rect 17817 32343 17826 32377
rect 17774 32334 17826 32343
rect 17934 32377 17986 32386
rect 17934 32343 17943 32377
rect 17943 32343 17977 32377
rect 17977 32343 17986 32377
rect 17934 32334 17986 32343
rect 18094 32377 18146 32386
rect 18094 32343 18103 32377
rect 18103 32343 18137 32377
rect 18137 32343 18146 32377
rect 18094 32334 18146 32343
rect 18254 32377 18306 32386
rect 18254 32343 18263 32377
rect 18263 32343 18297 32377
rect 18297 32343 18306 32377
rect 18254 32334 18306 32343
rect 18414 32377 18466 32386
rect 18414 32343 18423 32377
rect 18423 32343 18457 32377
rect 18457 32343 18466 32377
rect 18414 32334 18466 32343
rect 18574 32377 18626 32386
rect 18574 32343 18583 32377
rect 18583 32343 18617 32377
rect 18617 32343 18626 32377
rect 18574 32334 18626 32343
rect 18734 32377 18786 32386
rect 18734 32343 18743 32377
rect 18743 32343 18777 32377
rect 18777 32343 18786 32377
rect 18734 32334 18786 32343
rect 18894 32377 18946 32386
rect 18894 32343 18903 32377
rect 18903 32343 18937 32377
rect 18937 32343 18946 32377
rect 18894 32334 18946 32343
rect 23134 32377 23186 32386
rect 23134 32343 23143 32377
rect 23143 32343 23177 32377
rect 23177 32343 23186 32377
rect 23134 32334 23186 32343
rect 23294 32377 23346 32386
rect 23294 32343 23303 32377
rect 23303 32343 23337 32377
rect 23337 32343 23346 32377
rect 23294 32334 23346 32343
rect 23454 32377 23506 32386
rect 23454 32343 23463 32377
rect 23463 32343 23497 32377
rect 23497 32343 23506 32377
rect 23454 32334 23506 32343
rect 23614 32377 23666 32386
rect 23614 32343 23623 32377
rect 23623 32343 23657 32377
rect 23657 32343 23666 32377
rect 23614 32334 23666 32343
rect 23774 32377 23826 32386
rect 23774 32343 23783 32377
rect 23783 32343 23817 32377
rect 23817 32343 23826 32377
rect 23774 32334 23826 32343
rect 23934 32377 23986 32386
rect 23934 32343 23943 32377
rect 23943 32343 23977 32377
rect 23977 32343 23986 32377
rect 23934 32334 23986 32343
rect 24094 32377 24146 32386
rect 24094 32343 24103 32377
rect 24103 32343 24137 32377
rect 24137 32343 24146 32377
rect 24094 32334 24146 32343
rect 24254 32377 24306 32386
rect 24254 32343 24263 32377
rect 24263 32343 24297 32377
rect 24297 32343 24306 32377
rect 24254 32334 24306 32343
rect 24414 32377 24466 32386
rect 24414 32343 24423 32377
rect 24423 32343 24457 32377
rect 24457 32343 24466 32377
rect 24414 32334 24466 32343
rect 24574 32377 24626 32386
rect 24574 32343 24583 32377
rect 24583 32343 24617 32377
rect 24617 32343 24626 32377
rect 24574 32334 24626 32343
rect 24734 32377 24786 32386
rect 24734 32343 24743 32377
rect 24743 32343 24777 32377
rect 24777 32343 24786 32377
rect 24734 32334 24786 32343
rect 24894 32377 24946 32386
rect 24894 32343 24903 32377
rect 24903 32343 24937 32377
rect 24937 32343 24946 32377
rect 24894 32334 24946 32343
rect 25054 32377 25106 32386
rect 25054 32343 25063 32377
rect 25063 32343 25097 32377
rect 25097 32343 25106 32377
rect 25054 32334 25106 32343
rect 25214 32377 25266 32386
rect 25214 32343 25223 32377
rect 25223 32343 25257 32377
rect 25257 32343 25266 32377
rect 25214 32334 25266 32343
rect 25374 32377 25426 32386
rect 25374 32343 25383 32377
rect 25383 32343 25417 32377
rect 25417 32343 25426 32377
rect 25374 32334 25426 32343
rect 25534 32377 25586 32386
rect 25534 32343 25543 32377
rect 25543 32343 25577 32377
rect 25577 32343 25586 32377
rect 25534 32334 25586 32343
rect 25694 32377 25746 32386
rect 25694 32343 25703 32377
rect 25703 32343 25737 32377
rect 25737 32343 25746 32377
rect 25694 32334 25746 32343
rect 25854 32377 25906 32386
rect 25854 32343 25863 32377
rect 25863 32343 25897 32377
rect 25897 32343 25906 32377
rect 25854 32334 25906 32343
rect 26014 32377 26066 32386
rect 26014 32343 26023 32377
rect 26023 32343 26057 32377
rect 26057 32343 26066 32377
rect 26014 32334 26066 32343
rect 26174 32377 26226 32386
rect 26174 32343 26183 32377
rect 26183 32343 26217 32377
rect 26217 32343 26226 32377
rect 26174 32334 26226 32343
rect 26334 32377 26386 32386
rect 26334 32343 26343 32377
rect 26343 32343 26377 32377
rect 26377 32343 26386 32377
rect 26334 32334 26386 32343
rect 26494 32377 26546 32386
rect 26494 32343 26503 32377
rect 26503 32343 26537 32377
rect 26537 32343 26546 32377
rect 26494 32334 26546 32343
rect 26654 32377 26706 32386
rect 26654 32343 26663 32377
rect 26663 32343 26697 32377
rect 26697 32343 26706 32377
rect 26654 32334 26706 32343
rect 26814 32377 26866 32386
rect 26814 32343 26823 32377
rect 26823 32343 26857 32377
rect 26857 32343 26866 32377
rect 26814 32334 26866 32343
rect 26974 32377 27026 32386
rect 26974 32343 26983 32377
rect 26983 32343 27017 32377
rect 27017 32343 27026 32377
rect 26974 32334 27026 32343
rect 27134 32377 27186 32386
rect 27134 32343 27143 32377
rect 27143 32343 27177 32377
rect 27177 32343 27186 32377
rect 27134 32334 27186 32343
rect 27294 32377 27346 32386
rect 27294 32343 27303 32377
rect 27303 32343 27337 32377
rect 27337 32343 27346 32377
rect 27294 32334 27346 32343
rect 27454 32377 27506 32386
rect 27454 32343 27463 32377
rect 27463 32343 27497 32377
rect 27497 32343 27506 32377
rect 27454 32334 27506 32343
rect 27614 32377 27666 32386
rect 27614 32343 27623 32377
rect 27623 32343 27657 32377
rect 27657 32343 27666 32377
rect 27614 32334 27666 32343
rect 27774 32377 27826 32386
rect 27774 32343 27783 32377
rect 27783 32343 27817 32377
rect 27817 32343 27826 32377
rect 27774 32334 27826 32343
rect 27934 32377 27986 32386
rect 27934 32343 27943 32377
rect 27943 32343 27977 32377
rect 27977 32343 27986 32377
rect 27934 32334 27986 32343
rect 28094 32377 28146 32386
rect 28094 32343 28103 32377
rect 28103 32343 28137 32377
rect 28137 32343 28146 32377
rect 28094 32334 28146 32343
rect 28254 32377 28306 32386
rect 28254 32343 28263 32377
rect 28263 32343 28297 32377
rect 28297 32343 28306 32377
rect 28254 32334 28306 32343
rect 28414 32377 28466 32386
rect 28414 32343 28423 32377
rect 28423 32343 28457 32377
rect 28457 32343 28466 32377
rect 28414 32334 28466 32343
rect 28574 32377 28626 32386
rect 28574 32343 28583 32377
rect 28583 32343 28617 32377
rect 28617 32343 28626 32377
rect 28574 32334 28626 32343
rect 28734 32377 28786 32386
rect 28734 32343 28743 32377
rect 28743 32343 28777 32377
rect 28777 32343 28786 32377
rect 28734 32334 28786 32343
rect 28894 32377 28946 32386
rect 28894 32343 28903 32377
rect 28903 32343 28937 32377
rect 28937 32343 28946 32377
rect 28894 32334 28946 32343
rect 29054 32377 29106 32386
rect 29054 32343 29063 32377
rect 29063 32343 29097 32377
rect 29097 32343 29106 32377
rect 29054 32334 29106 32343
rect 29214 32377 29266 32386
rect 29214 32343 29223 32377
rect 29223 32343 29257 32377
rect 29257 32343 29266 32377
rect 29214 32334 29266 32343
rect 29374 32377 29426 32386
rect 29374 32343 29383 32377
rect 29383 32343 29417 32377
rect 29417 32343 29426 32377
rect 29374 32334 29426 32343
rect 33534 32377 33586 32386
rect 33534 32343 33543 32377
rect 33543 32343 33577 32377
rect 33577 32343 33586 32377
rect 33534 32334 33586 32343
rect 33694 32377 33746 32386
rect 33694 32343 33703 32377
rect 33703 32343 33737 32377
rect 33737 32343 33746 32377
rect 33694 32334 33746 32343
rect 33854 32377 33906 32386
rect 33854 32343 33863 32377
rect 33863 32343 33897 32377
rect 33897 32343 33906 32377
rect 33854 32334 33906 32343
rect 34014 32377 34066 32386
rect 34014 32343 34023 32377
rect 34023 32343 34057 32377
rect 34057 32343 34066 32377
rect 34014 32334 34066 32343
rect 34174 32377 34226 32386
rect 34174 32343 34183 32377
rect 34183 32343 34217 32377
rect 34217 32343 34226 32377
rect 34174 32334 34226 32343
rect 34334 32377 34386 32386
rect 34334 32343 34343 32377
rect 34343 32343 34377 32377
rect 34377 32343 34386 32377
rect 34334 32334 34386 32343
rect 34494 32377 34546 32386
rect 34494 32343 34503 32377
rect 34503 32343 34537 32377
rect 34537 32343 34546 32377
rect 34494 32334 34546 32343
rect 34654 32377 34706 32386
rect 34654 32343 34663 32377
rect 34663 32343 34697 32377
rect 34697 32343 34706 32377
rect 34654 32334 34706 32343
rect 34814 32377 34866 32386
rect 34814 32343 34823 32377
rect 34823 32343 34857 32377
rect 34857 32343 34866 32377
rect 34814 32334 34866 32343
rect 34974 32377 35026 32386
rect 34974 32343 34983 32377
rect 34983 32343 35017 32377
rect 35017 32343 35026 32377
rect 34974 32334 35026 32343
rect 35134 32377 35186 32386
rect 35134 32343 35143 32377
rect 35143 32343 35177 32377
rect 35177 32343 35186 32377
rect 35134 32334 35186 32343
rect 35294 32377 35346 32386
rect 35294 32343 35303 32377
rect 35303 32343 35337 32377
rect 35337 32343 35346 32377
rect 35294 32334 35346 32343
rect 35454 32377 35506 32386
rect 35454 32343 35463 32377
rect 35463 32343 35497 32377
rect 35497 32343 35506 32377
rect 35454 32334 35506 32343
rect 35614 32377 35666 32386
rect 35614 32343 35623 32377
rect 35623 32343 35657 32377
rect 35657 32343 35666 32377
rect 35614 32334 35666 32343
rect 35774 32377 35826 32386
rect 35774 32343 35783 32377
rect 35783 32343 35817 32377
rect 35817 32343 35826 32377
rect 35774 32334 35826 32343
rect 35934 32377 35986 32386
rect 35934 32343 35943 32377
rect 35943 32343 35977 32377
rect 35977 32343 35986 32377
rect 35934 32334 35986 32343
rect 36094 32377 36146 32386
rect 36094 32343 36103 32377
rect 36103 32343 36137 32377
rect 36137 32343 36146 32377
rect 36094 32334 36146 32343
rect 36254 32377 36306 32386
rect 36254 32343 36263 32377
rect 36263 32343 36297 32377
rect 36297 32343 36306 32377
rect 36254 32334 36306 32343
rect 36414 32377 36466 32386
rect 36414 32343 36423 32377
rect 36423 32343 36457 32377
rect 36457 32343 36466 32377
rect 36414 32334 36466 32343
rect 36574 32377 36626 32386
rect 36574 32343 36583 32377
rect 36583 32343 36617 32377
rect 36617 32343 36626 32377
rect 36574 32334 36626 32343
rect 36734 32377 36786 32386
rect 36734 32343 36743 32377
rect 36743 32343 36777 32377
rect 36777 32343 36786 32377
rect 36734 32334 36786 32343
rect 36894 32377 36946 32386
rect 36894 32343 36903 32377
rect 36903 32343 36937 32377
rect 36937 32343 36946 32377
rect 36894 32334 36946 32343
rect 37054 32377 37106 32386
rect 37054 32343 37063 32377
rect 37063 32343 37097 32377
rect 37097 32343 37106 32377
rect 37054 32334 37106 32343
rect 37214 32377 37266 32386
rect 37214 32343 37223 32377
rect 37223 32343 37257 32377
rect 37257 32343 37266 32377
rect 37214 32334 37266 32343
rect 37374 32377 37426 32386
rect 37374 32343 37383 32377
rect 37383 32343 37417 32377
rect 37417 32343 37426 32377
rect 37374 32334 37426 32343
rect 37534 32377 37586 32386
rect 37534 32343 37543 32377
rect 37543 32343 37577 32377
rect 37577 32343 37586 32377
rect 37534 32334 37586 32343
rect 37694 32377 37746 32386
rect 37694 32343 37703 32377
rect 37703 32343 37737 32377
rect 37737 32343 37746 32377
rect 37694 32334 37746 32343
rect 37854 32377 37906 32386
rect 37854 32343 37863 32377
rect 37863 32343 37897 32377
rect 37897 32343 37906 32377
rect 37854 32334 37906 32343
rect 38014 32377 38066 32386
rect 38014 32343 38023 32377
rect 38023 32343 38057 32377
rect 38057 32343 38066 32377
rect 38014 32334 38066 32343
rect 38174 32377 38226 32386
rect 38174 32343 38183 32377
rect 38183 32343 38217 32377
rect 38217 32343 38226 32377
rect 38174 32334 38226 32343
rect 38334 32377 38386 32386
rect 38334 32343 38343 32377
rect 38343 32343 38377 32377
rect 38377 32343 38386 32377
rect 38334 32334 38386 32343
rect 38494 32377 38546 32386
rect 38494 32343 38503 32377
rect 38503 32343 38537 32377
rect 38537 32343 38546 32377
rect 38494 32334 38546 32343
rect 38654 32377 38706 32386
rect 38654 32343 38663 32377
rect 38663 32343 38697 32377
rect 38697 32343 38706 32377
rect 38654 32334 38706 32343
rect 38814 32377 38866 32386
rect 38814 32343 38823 32377
rect 38823 32343 38857 32377
rect 38857 32343 38866 32377
rect 38814 32334 38866 32343
rect 38974 32377 39026 32386
rect 38974 32343 38983 32377
rect 38983 32343 39017 32377
rect 39017 32343 39026 32377
rect 38974 32334 39026 32343
rect 39134 32377 39186 32386
rect 39134 32343 39143 32377
rect 39143 32343 39177 32377
rect 39177 32343 39186 32377
rect 39134 32334 39186 32343
rect 39294 32377 39346 32386
rect 39294 32343 39303 32377
rect 39303 32343 39337 32377
rect 39337 32343 39346 32377
rect 39294 32334 39346 32343
rect 39454 32377 39506 32386
rect 39454 32343 39463 32377
rect 39463 32343 39497 32377
rect 39497 32343 39506 32377
rect 39454 32334 39506 32343
rect 39614 32377 39666 32386
rect 39614 32343 39623 32377
rect 39623 32343 39657 32377
rect 39657 32343 39666 32377
rect 39614 32334 39666 32343
rect 39774 32377 39826 32386
rect 39774 32343 39783 32377
rect 39783 32343 39817 32377
rect 39817 32343 39826 32377
rect 39774 32334 39826 32343
rect 39934 32377 39986 32386
rect 39934 32343 39943 32377
rect 39943 32343 39977 32377
rect 39977 32343 39986 32377
rect 39934 32334 39986 32343
rect 40094 32377 40146 32386
rect 40094 32343 40103 32377
rect 40103 32343 40137 32377
rect 40137 32343 40146 32377
rect 40094 32334 40146 32343
rect 40254 32377 40306 32386
rect 40254 32343 40263 32377
rect 40263 32343 40297 32377
rect 40297 32343 40306 32377
rect 40254 32334 40306 32343
rect 40414 32377 40466 32386
rect 40414 32343 40423 32377
rect 40423 32343 40457 32377
rect 40457 32343 40466 32377
rect 40414 32334 40466 32343
rect 40574 32377 40626 32386
rect 40574 32343 40583 32377
rect 40583 32343 40617 32377
rect 40617 32343 40626 32377
rect 40574 32334 40626 32343
rect 40734 32377 40786 32386
rect 40734 32343 40743 32377
rect 40743 32343 40777 32377
rect 40777 32343 40786 32377
rect 40734 32334 40786 32343
rect 40894 32377 40946 32386
rect 40894 32343 40903 32377
rect 40903 32343 40937 32377
rect 40937 32343 40946 32377
rect 40894 32334 40946 32343
rect 41054 32377 41106 32386
rect 41054 32343 41063 32377
rect 41063 32343 41097 32377
rect 41097 32343 41106 32377
rect 41054 32334 41106 32343
rect 41214 32377 41266 32386
rect 41214 32343 41223 32377
rect 41223 32343 41257 32377
rect 41257 32343 41266 32377
rect 41214 32334 41266 32343
rect 41374 32377 41426 32386
rect 41374 32343 41383 32377
rect 41383 32343 41417 32377
rect 41417 32343 41426 32377
rect 41374 32334 41426 32343
rect 41534 32377 41586 32386
rect 41534 32343 41543 32377
rect 41543 32343 41577 32377
rect 41577 32343 41586 32377
rect 41534 32334 41586 32343
rect 41694 32377 41746 32386
rect 41694 32343 41703 32377
rect 41703 32343 41737 32377
rect 41737 32343 41746 32377
rect 41694 32334 41746 32343
rect 41854 32377 41906 32386
rect 41854 32343 41863 32377
rect 41863 32343 41897 32377
rect 41897 32343 41906 32377
rect 41854 32334 41906 32343
rect 14 32057 66 32066
rect 14 32023 23 32057
rect 23 32023 57 32057
rect 57 32023 66 32057
rect 14 32014 66 32023
rect 174 32057 226 32066
rect 174 32023 183 32057
rect 183 32023 217 32057
rect 217 32023 226 32057
rect 174 32014 226 32023
rect 334 32057 386 32066
rect 334 32023 343 32057
rect 343 32023 377 32057
rect 377 32023 386 32057
rect 334 32014 386 32023
rect 494 32057 546 32066
rect 494 32023 503 32057
rect 503 32023 537 32057
rect 537 32023 546 32057
rect 494 32014 546 32023
rect 654 32057 706 32066
rect 654 32023 663 32057
rect 663 32023 697 32057
rect 697 32023 706 32057
rect 654 32014 706 32023
rect 814 32057 866 32066
rect 814 32023 823 32057
rect 823 32023 857 32057
rect 857 32023 866 32057
rect 814 32014 866 32023
rect 974 32057 1026 32066
rect 974 32023 983 32057
rect 983 32023 1017 32057
rect 1017 32023 1026 32057
rect 974 32014 1026 32023
rect 1134 32057 1186 32066
rect 1134 32023 1143 32057
rect 1143 32023 1177 32057
rect 1177 32023 1186 32057
rect 1134 32014 1186 32023
rect 1294 32057 1346 32066
rect 1294 32023 1303 32057
rect 1303 32023 1337 32057
rect 1337 32023 1346 32057
rect 1294 32014 1346 32023
rect 1454 32057 1506 32066
rect 1454 32023 1463 32057
rect 1463 32023 1497 32057
rect 1497 32023 1506 32057
rect 1454 32014 1506 32023
rect 1614 32057 1666 32066
rect 1614 32023 1623 32057
rect 1623 32023 1657 32057
rect 1657 32023 1666 32057
rect 1614 32014 1666 32023
rect 1774 32057 1826 32066
rect 1774 32023 1783 32057
rect 1783 32023 1817 32057
rect 1817 32023 1826 32057
rect 1774 32014 1826 32023
rect 1934 32057 1986 32066
rect 1934 32023 1943 32057
rect 1943 32023 1977 32057
rect 1977 32023 1986 32057
rect 1934 32014 1986 32023
rect 2094 32057 2146 32066
rect 2094 32023 2103 32057
rect 2103 32023 2137 32057
rect 2137 32023 2146 32057
rect 2094 32014 2146 32023
rect 2254 32057 2306 32066
rect 2254 32023 2263 32057
rect 2263 32023 2297 32057
rect 2297 32023 2306 32057
rect 2254 32014 2306 32023
rect 2414 32057 2466 32066
rect 2414 32023 2423 32057
rect 2423 32023 2457 32057
rect 2457 32023 2466 32057
rect 2414 32014 2466 32023
rect 2574 32057 2626 32066
rect 2574 32023 2583 32057
rect 2583 32023 2617 32057
rect 2617 32023 2626 32057
rect 2574 32014 2626 32023
rect 2734 32057 2786 32066
rect 2734 32023 2743 32057
rect 2743 32023 2777 32057
rect 2777 32023 2786 32057
rect 2734 32014 2786 32023
rect 2894 32057 2946 32066
rect 2894 32023 2903 32057
rect 2903 32023 2937 32057
rect 2937 32023 2946 32057
rect 2894 32014 2946 32023
rect 3054 32057 3106 32066
rect 3054 32023 3063 32057
rect 3063 32023 3097 32057
rect 3097 32023 3106 32057
rect 3054 32014 3106 32023
rect 3214 32057 3266 32066
rect 3214 32023 3223 32057
rect 3223 32023 3257 32057
rect 3257 32023 3266 32057
rect 3214 32014 3266 32023
rect 3374 32057 3426 32066
rect 3374 32023 3383 32057
rect 3383 32023 3417 32057
rect 3417 32023 3426 32057
rect 3374 32014 3426 32023
rect 3534 32057 3586 32066
rect 3534 32023 3543 32057
rect 3543 32023 3577 32057
rect 3577 32023 3586 32057
rect 3534 32014 3586 32023
rect 3694 32057 3746 32066
rect 3694 32023 3703 32057
rect 3703 32023 3737 32057
rect 3737 32023 3746 32057
rect 3694 32014 3746 32023
rect 3854 32057 3906 32066
rect 3854 32023 3863 32057
rect 3863 32023 3897 32057
rect 3897 32023 3906 32057
rect 3854 32014 3906 32023
rect 4014 32057 4066 32066
rect 4014 32023 4023 32057
rect 4023 32023 4057 32057
rect 4057 32023 4066 32057
rect 4014 32014 4066 32023
rect 4174 32057 4226 32066
rect 4174 32023 4183 32057
rect 4183 32023 4217 32057
rect 4217 32023 4226 32057
rect 4174 32014 4226 32023
rect 4334 32057 4386 32066
rect 4334 32023 4343 32057
rect 4343 32023 4377 32057
rect 4377 32023 4386 32057
rect 4334 32014 4386 32023
rect 4494 32057 4546 32066
rect 4494 32023 4503 32057
rect 4503 32023 4537 32057
rect 4537 32023 4546 32057
rect 4494 32014 4546 32023
rect 4654 32057 4706 32066
rect 4654 32023 4663 32057
rect 4663 32023 4697 32057
rect 4697 32023 4706 32057
rect 4654 32014 4706 32023
rect 4814 32057 4866 32066
rect 4814 32023 4823 32057
rect 4823 32023 4857 32057
rect 4857 32023 4866 32057
rect 4814 32014 4866 32023
rect 4974 32057 5026 32066
rect 4974 32023 4983 32057
rect 4983 32023 5017 32057
rect 5017 32023 5026 32057
rect 4974 32014 5026 32023
rect 5134 32057 5186 32066
rect 5134 32023 5143 32057
rect 5143 32023 5177 32057
rect 5177 32023 5186 32057
rect 5134 32014 5186 32023
rect 5294 32057 5346 32066
rect 5294 32023 5303 32057
rect 5303 32023 5337 32057
rect 5337 32023 5346 32057
rect 5294 32014 5346 32023
rect 5454 32057 5506 32066
rect 5454 32023 5463 32057
rect 5463 32023 5497 32057
rect 5497 32023 5506 32057
rect 5454 32014 5506 32023
rect 5614 32057 5666 32066
rect 5614 32023 5623 32057
rect 5623 32023 5657 32057
rect 5657 32023 5666 32057
rect 5614 32014 5666 32023
rect 5774 32057 5826 32066
rect 5774 32023 5783 32057
rect 5783 32023 5817 32057
rect 5817 32023 5826 32057
rect 5774 32014 5826 32023
rect 5934 32057 5986 32066
rect 5934 32023 5943 32057
rect 5943 32023 5977 32057
rect 5977 32023 5986 32057
rect 5934 32014 5986 32023
rect 6094 32057 6146 32066
rect 6094 32023 6103 32057
rect 6103 32023 6137 32057
rect 6137 32023 6146 32057
rect 6094 32014 6146 32023
rect 6254 32057 6306 32066
rect 6254 32023 6263 32057
rect 6263 32023 6297 32057
rect 6297 32023 6306 32057
rect 6254 32014 6306 32023
rect 6414 32057 6466 32066
rect 6414 32023 6423 32057
rect 6423 32023 6457 32057
rect 6457 32023 6466 32057
rect 6414 32014 6466 32023
rect 6574 32057 6626 32066
rect 6574 32023 6583 32057
rect 6583 32023 6617 32057
rect 6617 32023 6626 32057
rect 6574 32014 6626 32023
rect 6734 32057 6786 32066
rect 6734 32023 6743 32057
rect 6743 32023 6777 32057
rect 6777 32023 6786 32057
rect 6734 32014 6786 32023
rect 6894 32057 6946 32066
rect 6894 32023 6903 32057
rect 6903 32023 6937 32057
rect 6937 32023 6946 32057
rect 6894 32014 6946 32023
rect 7054 32057 7106 32066
rect 7054 32023 7063 32057
rect 7063 32023 7097 32057
rect 7097 32023 7106 32057
rect 7054 32014 7106 32023
rect 7214 32057 7266 32066
rect 7214 32023 7223 32057
rect 7223 32023 7257 32057
rect 7257 32023 7266 32057
rect 7214 32014 7266 32023
rect 7374 32057 7426 32066
rect 7374 32023 7383 32057
rect 7383 32023 7417 32057
rect 7417 32023 7426 32057
rect 7374 32014 7426 32023
rect 7534 32057 7586 32066
rect 7534 32023 7543 32057
rect 7543 32023 7577 32057
rect 7577 32023 7586 32057
rect 7534 32014 7586 32023
rect 7694 32057 7746 32066
rect 7694 32023 7703 32057
rect 7703 32023 7737 32057
rect 7737 32023 7746 32057
rect 7694 32014 7746 32023
rect 7854 32057 7906 32066
rect 7854 32023 7863 32057
rect 7863 32023 7897 32057
rect 7897 32023 7906 32057
rect 7854 32014 7906 32023
rect 8014 32057 8066 32066
rect 8014 32023 8023 32057
rect 8023 32023 8057 32057
rect 8057 32023 8066 32057
rect 8014 32014 8066 32023
rect 8174 32057 8226 32066
rect 8174 32023 8183 32057
rect 8183 32023 8217 32057
rect 8217 32023 8226 32057
rect 8174 32014 8226 32023
rect 8334 32057 8386 32066
rect 8334 32023 8343 32057
rect 8343 32023 8377 32057
rect 8377 32023 8386 32057
rect 8334 32014 8386 32023
rect 12494 32057 12546 32066
rect 12494 32023 12503 32057
rect 12503 32023 12537 32057
rect 12537 32023 12546 32057
rect 12494 32014 12546 32023
rect 12654 32057 12706 32066
rect 12654 32023 12663 32057
rect 12663 32023 12697 32057
rect 12697 32023 12706 32057
rect 12654 32014 12706 32023
rect 12814 32057 12866 32066
rect 12814 32023 12823 32057
rect 12823 32023 12857 32057
rect 12857 32023 12866 32057
rect 12814 32014 12866 32023
rect 12974 32057 13026 32066
rect 12974 32023 12983 32057
rect 12983 32023 13017 32057
rect 13017 32023 13026 32057
rect 12974 32014 13026 32023
rect 13134 32057 13186 32066
rect 13134 32023 13143 32057
rect 13143 32023 13177 32057
rect 13177 32023 13186 32057
rect 13134 32014 13186 32023
rect 13294 32057 13346 32066
rect 13294 32023 13303 32057
rect 13303 32023 13337 32057
rect 13337 32023 13346 32057
rect 13294 32014 13346 32023
rect 13454 32057 13506 32066
rect 13454 32023 13463 32057
rect 13463 32023 13497 32057
rect 13497 32023 13506 32057
rect 13454 32014 13506 32023
rect 13614 32057 13666 32066
rect 13614 32023 13623 32057
rect 13623 32023 13657 32057
rect 13657 32023 13666 32057
rect 13614 32014 13666 32023
rect 13774 32057 13826 32066
rect 13774 32023 13783 32057
rect 13783 32023 13817 32057
rect 13817 32023 13826 32057
rect 13774 32014 13826 32023
rect 13934 32057 13986 32066
rect 13934 32023 13943 32057
rect 13943 32023 13977 32057
rect 13977 32023 13986 32057
rect 13934 32014 13986 32023
rect 14094 32057 14146 32066
rect 14094 32023 14103 32057
rect 14103 32023 14137 32057
rect 14137 32023 14146 32057
rect 14094 32014 14146 32023
rect 14254 32057 14306 32066
rect 14254 32023 14263 32057
rect 14263 32023 14297 32057
rect 14297 32023 14306 32057
rect 14254 32014 14306 32023
rect 14414 32057 14466 32066
rect 14414 32023 14423 32057
rect 14423 32023 14457 32057
rect 14457 32023 14466 32057
rect 14414 32014 14466 32023
rect 14574 32057 14626 32066
rect 14574 32023 14583 32057
rect 14583 32023 14617 32057
rect 14617 32023 14626 32057
rect 14574 32014 14626 32023
rect 14734 32057 14786 32066
rect 14734 32023 14743 32057
rect 14743 32023 14777 32057
rect 14777 32023 14786 32057
rect 14734 32014 14786 32023
rect 14894 32057 14946 32066
rect 14894 32023 14903 32057
rect 14903 32023 14937 32057
rect 14937 32023 14946 32057
rect 14894 32014 14946 32023
rect 15054 32057 15106 32066
rect 15054 32023 15063 32057
rect 15063 32023 15097 32057
rect 15097 32023 15106 32057
rect 15054 32014 15106 32023
rect 15214 32057 15266 32066
rect 15214 32023 15223 32057
rect 15223 32023 15257 32057
rect 15257 32023 15266 32057
rect 15214 32014 15266 32023
rect 15374 32057 15426 32066
rect 15374 32023 15383 32057
rect 15383 32023 15417 32057
rect 15417 32023 15426 32057
rect 15374 32014 15426 32023
rect 15534 32057 15586 32066
rect 15534 32023 15543 32057
rect 15543 32023 15577 32057
rect 15577 32023 15586 32057
rect 15534 32014 15586 32023
rect 15694 32057 15746 32066
rect 15694 32023 15703 32057
rect 15703 32023 15737 32057
rect 15737 32023 15746 32057
rect 15694 32014 15746 32023
rect 15854 32057 15906 32066
rect 15854 32023 15863 32057
rect 15863 32023 15897 32057
rect 15897 32023 15906 32057
rect 15854 32014 15906 32023
rect 16014 32057 16066 32066
rect 16014 32023 16023 32057
rect 16023 32023 16057 32057
rect 16057 32023 16066 32057
rect 16014 32014 16066 32023
rect 16174 32057 16226 32066
rect 16174 32023 16183 32057
rect 16183 32023 16217 32057
rect 16217 32023 16226 32057
rect 16174 32014 16226 32023
rect 16334 32057 16386 32066
rect 16334 32023 16343 32057
rect 16343 32023 16377 32057
rect 16377 32023 16386 32057
rect 16334 32014 16386 32023
rect 16494 32057 16546 32066
rect 16494 32023 16503 32057
rect 16503 32023 16537 32057
rect 16537 32023 16546 32057
rect 16494 32014 16546 32023
rect 16654 32057 16706 32066
rect 16654 32023 16663 32057
rect 16663 32023 16697 32057
rect 16697 32023 16706 32057
rect 16654 32014 16706 32023
rect 16814 32057 16866 32066
rect 16814 32023 16823 32057
rect 16823 32023 16857 32057
rect 16857 32023 16866 32057
rect 16814 32014 16866 32023
rect 16974 32057 17026 32066
rect 16974 32023 16983 32057
rect 16983 32023 17017 32057
rect 17017 32023 17026 32057
rect 16974 32014 17026 32023
rect 17134 32057 17186 32066
rect 17134 32023 17143 32057
rect 17143 32023 17177 32057
rect 17177 32023 17186 32057
rect 17134 32014 17186 32023
rect 17294 32057 17346 32066
rect 17294 32023 17303 32057
rect 17303 32023 17337 32057
rect 17337 32023 17346 32057
rect 17294 32014 17346 32023
rect 17454 32057 17506 32066
rect 17454 32023 17463 32057
rect 17463 32023 17497 32057
rect 17497 32023 17506 32057
rect 17454 32014 17506 32023
rect 17614 32057 17666 32066
rect 17614 32023 17623 32057
rect 17623 32023 17657 32057
rect 17657 32023 17666 32057
rect 17614 32014 17666 32023
rect 17774 32057 17826 32066
rect 17774 32023 17783 32057
rect 17783 32023 17817 32057
rect 17817 32023 17826 32057
rect 17774 32014 17826 32023
rect 17934 32057 17986 32066
rect 17934 32023 17943 32057
rect 17943 32023 17977 32057
rect 17977 32023 17986 32057
rect 17934 32014 17986 32023
rect 18094 32057 18146 32066
rect 18094 32023 18103 32057
rect 18103 32023 18137 32057
rect 18137 32023 18146 32057
rect 18094 32014 18146 32023
rect 18254 32057 18306 32066
rect 18254 32023 18263 32057
rect 18263 32023 18297 32057
rect 18297 32023 18306 32057
rect 18254 32014 18306 32023
rect 18414 32057 18466 32066
rect 18414 32023 18423 32057
rect 18423 32023 18457 32057
rect 18457 32023 18466 32057
rect 18414 32014 18466 32023
rect 18574 32057 18626 32066
rect 18574 32023 18583 32057
rect 18583 32023 18617 32057
rect 18617 32023 18626 32057
rect 18574 32014 18626 32023
rect 18734 32057 18786 32066
rect 18734 32023 18743 32057
rect 18743 32023 18777 32057
rect 18777 32023 18786 32057
rect 18734 32014 18786 32023
rect 18894 32057 18946 32066
rect 18894 32023 18903 32057
rect 18903 32023 18937 32057
rect 18937 32023 18946 32057
rect 18894 32014 18946 32023
rect 23134 32057 23186 32066
rect 23134 32023 23143 32057
rect 23143 32023 23177 32057
rect 23177 32023 23186 32057
rect 23134 32014 23186 32023
rect 23294 32057 23346 32066
rect 23294 32023 23303 32057
rect 23303 32023 23337 32057
rect 23337 32023 23346 32057
rect 23294 32014 23346 32023
rect 23454 32057 23506 32066
rect 23454 32023 23463 32057
rect 23463 32023 23497 32057
rect 23497 32023 23506 32057
rect 23454 32014 23506 32023
rect 23614 32057 23666 32066
rect 23614 32023 23623 32057
rect 23623 32023 23657 32057
rect 23657 32023 23666 32057
rect 23614 32014 23666 32023
rect 23774 32057 23826 32066
rect 23774 32023 23783 32057
rect 23783 32023 23817 32057
rect 23817 32023 23826 32057
rect 23774 32014 23826 32023
rect 23934 32057 23986 32066
rect 23934 32023 23943 32057
rect 23943 32023 23977 32057
rect 23977 32023 23986 32057
rect 23934 32014 23986 32023
rect 24094 32057 24146 32066
rect 24094 32023 24103 32057
rect 24103 32023 24137 32057
rect 24137 32023 24146 32057
rect 24094 32014 24146 32023
rect 24254 32057 24306 32066
rect 24254 32023 24263 32057
rect 24263 32023 24297 32057
rect 24297 32023 24306 32057
rect 24254 32014 24306 32023
rect 24414 32057 24466 32066
rect 24414 32023 24423 32057
rect 24423 32023 24457 32057
rect 24457 32023 24466 32057
rect 24414 32014 24466 32023
rect 24574 32057 24626 32066
rect 24574 32023 24583 32057
rect 24583 32023 24617 32057
rect 24617 32023 24626 32057
rect 24574 32014 24626 32023
rect 24734 32057 24786 32066
rect 24734 32023 24743 32057
rect 24743 32023 24777 32057
rect 24777 32023 24786 32057
rect 24734 32014 24786 32023
rect 24894 32057 24946 32066
rect 24894 32023 24903 32057
rect 24903 32023 24937 32057
rect 24937 32023 24946 32057
rect 24894 32014 24946 32023
rect 25054 32057 25106 32066
rect 25054 32023 25063 32057
rect 25063 32023 25097 32057
rect 25097 32023 25106 32057
rect 25054 32014 25106 32023
rect 25214 32057 25266 32066
rect 25214 32023 25223 32057
rect 25223 32023 25257 32057
rect 25257 32023 25266 32057
rect 25214 32014 25266 32023
rect 25374 32057 25426 32066
rect 25374 32023 25383 32057
rect 25383 32023 25417 32057
rect 25417 32023 25426 32057
rect 25374 32014 25426 32023
rect 25534 32057 25586 32066
rect 25534 32023 25543 32057
rect 25543 32023 25577 32057
rect 25577 32023 25586 32057
rect 25534 32014 25586 32023
rect 25694 32057 25746 32066
rect 25694 32023 25703 32057
rect 25703 32023 25737 32057
rect 25737 32023 25746 32057
rect 25694 32014 25746 32023
rect 25854 32057 25906 32066
rect 25854 32023 25863 32057
rect 25863 32023 25897 32057
rect 25897 32023 25906 32057
rect 25854 32014 25906 32023
rect 26014 32057 26066 32066
rect 26014 32023 26023 32057
rect 26023 32023 26057 32057
rect 26057 32023 26066 32057
rect 26014 32014 26066 32023
rect 26174 32057 26226 32066
rect 26174 32023 26183 32057
rect 26183 32023 26217 32057
rect 26217 32023 26226 32057
rect 26174 32014 26226 32023
rect 26334 32057 26386 32066
rect 26334 32023 26343 32057
rect 26343 32023 26377 32057
rect 26377 32023 26386 32057
rect 26334 32014 26386 32023
rect 26494 32057 26546 32066
rect 26494 32023 26503 32057
rect 26503 32023 26537 32057
rect 26537 32023 26546 32057
rect 26494 32014 26546 32023
rect 26654 32057 26706 32066
rect 26654 32023 26663 32057
rect 26663 32023 26697 32057
rect 26697 32023 26706 32057
rect 26654 32014 26706 32023
rect 26814 32057 26866 32066
rect 26814 32023 26823 32057
rect 26823 32023 26857 32057
rect 26857 32023 26866 32057
rect 26814 32014 26866 32023
rect 26974 32057 27026 32066
rect 26974 32023 26983 32057
rect 26983 32023 27017 32057
rect 27017 32023 27026 32057
rect 26974 32014 27026 32023
rect 27134 32057 27186 32066
rect 27134 32023 27143 32057
rect 27143 32023 27177 32057
rect 27177 32023 27186 32057
rect 27134 32014 27186 32023
rect 27294 32057 27346 32066
rect 27294 32023 27303 32057
rect 27303 32023 27337 32057
rect 27337 32023 27346 32057
rect 27294 32014 27346 32023
rect 27454 32057 27506 32066
rect 27454 32023 27463 32057
rect 27463 32023 27497 32057
rect 27497 32023 27506 32057
rect 27454 32014 27506 32023
rect 27614 32057 27666 32066
rect 27614 32023 27623 32057
rect 27623 32023 27657 32057
rect 27657 32023 27666 32057
rect 27614 32014 27666 32023
rect 27774 32057 27826 32066
rect 27774 32023 27783 32057
rect 27783 32023 27817 32057
rect 27817 32023 27826 32057
rect 27774 32014 27826 32023
rect 27934 32057 27986 32066
rect 27934 32023 27943 32057
rect 27943 32023 27977 32057
rect 27977 32023 27986 32057
rect 27934 32014 27986 32023
rect 28094 32057 28146 32066
rect 28094 32023 28103 32057
rect 28103 32023 28137 32057
rect 28137 32023 28146 32057
rect 28094 32014 28146 32023
rect 28254 32057 28306 32066
rect 28254 32023 28263 32057
rect 28263 32023 28297 32057
rect 28297 32023 28306 32057
rect 28254 32014 28306 32023
rect 28414 32057 28466 32066
rect 28414 32023 28423 32057
rect 28423 32023 28457 32057
rect 28457 32023 28466 32057
rect 28414 32014 28466 32023
rect 28574 32057 28626 32066
rect 28574 32023 28583 32057
rect 28583 32023 28617 32057
rect 28617 32023 28626 32057
rect 28574 32014 28626 32023
rect 28734 32057 28786 32066
rect 28734 32023 28743 32057
rect 28743 32023 28777 32057
rect 28777 32023 28786 32057
rect 28734 32014 28786 32023
rect 28894 32057 28946 32066
rect 28894 32023 28903 32057
rect 28903 32023 28937 32057
rect 28937 32023 28946 32057
rect 28894 32014 28946 32023
rect 29054 32057 29106 32066
rect 29054 32023 29063 32057
rect 29063 32023 29097 32057
rect 29097 32023 29106 32057
rect 29054 32014 29106 32023
rect 29214 32057 29266 32066
rect 29214 32023 29223 32057
rect 29223 32023 29257 32057
rect 29257 32023 29266 32057
rect 29214 32014 29266 32023
rect 29374 32057 29426 32066
rect 29374 32023 29383 32057
rect 29383 32023 29417 32057
rect 29417 32023 29426 32057
rect 29374 32014 29426 32023
rect 33534 32057 33586 32066
rect 33534 32023 33543 32057
rect 33543 32023 33577 32057
rect 33577 32023 33586 32057
rect 33534 32014 33586 32023
rect 33694 32057 33746 32066
rect 33694 32023 33703 32057
rect 33703 32023 33737 32057
rect 33737 32023 33746 32057
rect 33694 32014 33746 32023
rect 33854 32057 33906 32066
rect 33854 32023 33863 32057
rect 33863 32023 33897 32057
rect 33897 32023 33906 32057
rect 33854 32014 33906 32023
rect 34014 32057 34066 32066
rect 34014 32023 34023 32057
rect 34023 32023 34057 32057
rect 34057 32023 34066 32057
rect 34014 32014 34066 32023
rect 34174 32057 34226 32066
rect 34174 32023 34183 32057
rect 34183 32023 34217 32057
rect 34217 32023 34226 32057
rect 34174 32014 34226 32023
rect 34334 32057 34386 32066
rect 34334 32023 34343 32057
rect 34343 32023 34377 32057
rect 34377 32023 34386 32057
rect 34334 32014 34386 32023
rect 34494 32057 34546 32066
rect 34494 32023 34503 32057
rect 34503 32023 34537 32057
rect 34537 32023 34546 32057
rect 34494 32014 34546 32023
rect 34654 32057 34706 32066
rect 34654 32023 34663 32057
rect 34663 32023 34697 32057
rect 34697 32023 34706 32057
rect 34654 32014 34706 32023
rect 34814 32057 34866 32066
rect 34814 32023 34823 32057
rect 34823 32023 34857 32057
rect 34857 32023 34866 32057
rect 34814 32014 34866 32023
rect 34974 32057 35026 32066
rect 34974 32023 34983 32057
rect 34983 32023 35017 32057
rect 35017 32023 35026 32057
rect 34974 32014 35026 32023
rect 35134 32057 35186 32066
rect 35134 32023 35143 32057
rect 35143 32023 35177 32057
rect 35177 32023 35186 32057
rect 35134 32014 35186 32023
rect 35294 32057 35346 32066
rect 35294 32023 35303 32057
rect 35303 32023 35337 32057
rect 35337 32023 35346 32057
rect 35294 32014 35346 32023
rect 35454 32057 35506 32066
rect 35454 32023 35463 32057
rect 35463 32023 35497 32057
rect 35497 32023 35506 32057
rect 35454 32014 35506 32023
rect 35614 32057 35666 32066
rect 35614 32023 35623 32057
rect 35623 32023 35657 32057
rect 35657 32023 35666 32057
rect 35614 32014 35666 32023
rect 35774 32057 35826 32066
rect 35774 32023 35783 32057
rect 35783 32023 35817 32057
rect 35817 32023 35826 32057
rect 35774 32014 35826 32023
rect 35934 32057 35986 32066
rect 35934 32023 35943 32057
rect 35943 32023 35977 32057
rect 35977 32023 35986 32057
rect 35934 32014 35986 32023
rect 36094 32057 36146 32066
rect 36094 32023 36103 32057
rect 36103 32023 36137 32057
rect 36137 32023 36146 32057
rect 36094 32014 36146 32023
rect 36254 32057 36306 32066
rect 36254 32023 36263 32057
rect 36263 32023 36297 32057
rect 36297 32023 36306 32057
rect 36254 32014 36306 32023
rect 36414 32057 36466 32066
rect 36414 32023 36423 32057
rect 36423 32023 36457 32057
rect 36457 32023 36466 32057
rect 36414 32014 36466 32023
rect 36574 32057 36626 32066
rect 36574 32023 36583 32057
rect 36583 32023 36617 32057
rect 36617 32023 36626 32057
rect 36574 32014 36626 32023
rect 36734 32057 36786 32066
rect 36734 32023 36743 32057
rect 36743 32023 36777 32057
rect 36777 32023 36786 32057
rect 36734 32014 36786 32023
rect 36894 32057 36946 32066
rect 36894 32023 36903 32057
rect 36903 32023 36937 32057
rect 36937 32023 36946 32057
rect 36894 32014 36946 32023
rect 37054 32057 37106 32066
rect 37054 32023 37063 32057
rect 37063 32023 37097 32057
rect 37097 32023 37106 32057
rect 37054 32014 37106 32023
rect 37214 32057 37266 32066
rect 37214 32023 37223 32057
rect 37223 32023 37257 32057
rect 37257 32023 37266 32057
rect 37214 32014 37266 32023
rect 37374 32057 37426 32066
rect 37374 32023 37383 32057
rect 37383 32023 37417 32057
rect 37417 32023 37426 32057
rect 37374 32014 37426 32023
rect 37534 32057 37586 32066
rect 37534 32023 37543 32057
rect 37543 32023 37577 32057
rect 37577 32023 37586 32057
rect 37534 32014 37586 32023
rect 37694 32057 37746 32066
rect 37694 32023 37703 32057
rect 37703 32023 37737 32057
rect 37737 32023 37746 32057
rect 37694 32014 37746 32023
rect 37854 32057 37906 32066
rect 37854 32023 37863 32057
rect 37863 32023 37897 32057
rect 37897 32023 37906 32057
rect 37854 32014 37906 32023
rect 38014 32057 38066 32066
rect 38014 32023 38023 32057
rect 38023 32023 38057 32057
rect 38057 32023 38066 32057
rect 38014 32014 38066 32023
rect 38174 32057 38226 32066
rect 38174 32023 38183 32057
rect 38183 32023 38217 32057
rect 38217 32023 38226 32057
rect 38174 32014 38226 32023
rect 38334 32057 38386 32066
rect 38334 32023 38343 32057
rect 38343 32023 38377 32057
rect 38377 32023 38386 32057
rect 38334 32014 38386 32023
rect 38494 32057 38546 32066
rect 38494 32023 38503 32057
rect 38503 32023 38537 32057
rect 38537 32023 38546 32057
rect 38494 32014 38546 32023
rect 38654 32057 38706 32066
rect 38654 32023 38663 32057
rect 38663 32023 38697 32057
rect 38697 32023 38706 32057
rect 38654 32014 38706 32023
rect 38814 32057 38866 32066
rect 38814 32023 38823 32057
rect 38823 32023 38857 32057
rect 38857 32023 38866 32057
rect 38814 32014 38866 32023
rect 38974 32057 39026 32066
rect 38974 32023 38983 32057
rect 38983 32023 39017 32057
rect 39017 32023 39026 32057
rect 38974 32014 39026 32023
rect 39134 32057 39186 32066
rect 39134 32023 39143 32057
rect 39143 32023 39177 32057
rect 39177 32023 39186 32057
rect 39134 32014 39186 32023
rect 39294 32057 39346 32066
rect 39294 32023 39303 32057
rect 39303 32023 39337 32057
rect 39337 32023 39346 32057
rect 39294 32014 39346 32023
rect 39454 32057 39506 32066
rect 39454 32023 39463 32057
rect 39463 32023 39497 32057
rect 39497 32023 39506 32057
rect 39454 32014 39506 32023
rect 39614 32057 39666 32066
rect 39614 32023 39623 32057
rect 39623 32023 39657 32057
rect 39657 32023 39666 32057
rect 39614 32014 39666 32023
rect 39774 32057 39826 32066
rect 39774 32023 39783 32057
rect 39783 32023 39817 32057
rect 39817 32023 39826 32057
rect 39774 32014 39826 32023
rect 39934 32057 39986 32066
rect 39934 32023 39943 32057
rect 39943 32023 39977 32057
rect 39977 32023 39986 32057
rect 39934 32014 39986 32023
rect 40094 32057 40146 32066
rect 40094 32023 40103 32057
rect 40103 32023 40137 32057
rect 40137 32023 40146 32057
rect 40094 32014 40146 32023
rect 40254 32057 40306 32066
rect 40254 32023 40263 32057
rect 40263 32023 40297 32057
rect 40297 32023 40306 32057
rect 40254 32014 40306 32023
rect 40414 32057 40466 32066
rect 40414 32023 40423 32057
rect 40423 32023 40457 32057
rect 40457 32023 40466 32057
rect 40414 32014 40466 32023
rect 40574 32057 40626 32066
rect 40574 32023 40583 32057
rect 40583 32023 40617 32057
rect 40617 32023 40626 32057
rect 40574 32014 40626 32023
rect 40734 32057 40786 32066
rect 40734 32023 40743 32057
rect 40743 32023 40777 32057
rect 40777 32023 40786 32057
rect 40734 32014 40786 32023
rect 40894 32057 40946 32066
rect 40894 32023 40903 32057
rect 40903 32023 40937 32057
rect 40937 32023 40946 32057
rect 40894 32014 40946 32023
rect 41054 32057 41106 32066
rect 41054 32023 41063 32057
rect 41063 32023 41097 32057
rect 41097 32023 41106 32057
rect 41054 32014 41106 32023
rect 41214 32057 41266 32066
rect 41214 32023 41223 32057
rect 41223 32023 41257 32057
rect 41257 32023 41266 32057
rect 41214 32014 41266 32023
rect 41374 32057 41426 32066
rect 41374 32023 41383 32057
rect 41383 32023 41417 32057
rect 41417 32023 41426 32057
rect 41374 32014 41426 32023
rect 41534 32057 41586 32066
rect 41534 32023 41543 32057
rect 41543 32023 41577 32057
rect 41577 32023 41586 32057
rect 41534 32014 41586 32023
rect 41694 32057 41746 32066
rect 41694 32023 41703 32057
rect 41703 32023 41737 32057
rect 41737 32023 41746 32057
rect 41694 32014 41746 32023
rect 41854 32057 41906 32066
rect 41854 32023 41863 32057
rect 41863 32023 41897 32057
rect 41897 32023 41906 32057
rect 41854 32014 41906 32023
rect 14 31737 66 31746
rect 14 31703 23 31737
rect 23 31703 57 31737
rect 57 31703 66 31737
rect 14 31694 66 31703
rect 174 31737 226 31746
rect 174 31703 183 31737
rect 183 31703 217 31737
rect 217 31703 226 31737
rect 174 31694 226 31703
rect 334 31737 386 31746
rect 334 31703 343 31737
rect 343 31703 377 31737
rect 377 31703 386 31737
rect 334 31694 386 31703
rect 494 31737 546 31746
rect 494 31703 503 31737
rect 503 31703 537 31737
rect 537 31703 546 31737
rect 494 31694 546 31703
rect 654 31737 706 31746
rect 654 31703 663 31737
rect 663 31703 697 31737
rect 697 31703 706 31737
rect 654 31694 706 31703
rect 814 31737 866 31746
rect 814 31703 823 31737
rect 823 31703 857 31737
rect 857 31703 866 31737
rect 814 31694 866 31703
rect 974 31737 1026 31746
rect 974 31703 983 31737
rect 983 31703 1017 31737
rect 1017 31703 1026 31737
rect 974 31694 1026 31703
rect 1134 31737 1186 31746
rect 1134 31703 1143 31737
rect 1143 31703 1177 31737
rect 1177 31703 1186 31737
rect 1134 31694 1186 31703
rect 1294 31737 1346 31746
rect 1294 31703 1303 31737
rect 1303 31703 1337 31737
rect 1337 31703 1346 31737
rect 1294 31694 1346 31703
rect 1454 31737 1506 31746
rect 1454 31703 1463 31737
rect 1463 31703 1497 31737
rect 1497 31703 1506 31737
rect 1454 31694 1506 31703
rect 1614 31737 1666 31746
rect 1614 31703 1623 31737
rect 1623 31703 1657 31737
rect 1657 31703 1666 31737
rect 1614 31694 1666 31703
rect 1774 31737 1826 31746
rect 1774 31703 1783 31737
rect 1783 31703 1817 31737
rect 1817 31703 1826 31737
rect 1774 31694 1826 31703
rect 1934 31737 1986 31746
rect 1934 31703 1943 31737
rect 1943 31703 1977 31737
rect 1977 31703 1986 31737
rect 1934 31694 1986 31703
rect 2094 31737 2146 31746
rect 2094 31703 2103 31737
rect 2103 31703 2137 31737
rect 2137 31703 2146 31737
rect 2094 31694 2146 31703
rect 2254 31737 2306 31746
rect 2254 31703 2263 31737
rect 2263 31703 2297 31737
rect 2297 31703 2306 31737
rect 2254 31694 2306 31703
rect 2414 31737 2466 31746
rect 2414 31703 2423 31737
rect 2423 31703 2457 31737
rect 2457 31703 2466 31737
rect 2414 31694 2466 31703
rect 2574 31737 2626 31746
rect 2574 31703 2583 31737
rect 2583 31703 2617 31737
rect 2617 31703 2626 31737
rect 2574 31694 2626 31703
rect 2734 31737 2786 31746
rect 2734 31703 2743 31737
rect 2743 31703 2777 31737
rect 2777 31703 2786 31737
rect 2734 31694 2786 31703
rect 2894 31737 2946 31746
rect 2894 31703 2903 31737
rect 2903 31703 2937 31737
rect 2937 31703 2946 31737
rect 2894 31694 2946 31703
rect 3054 31737 3106 31746
rect 3054 31703 3063 31737
rect 3063 31703 3097 31737
rect 3097 31703 3106 31737
rect 3054 31694 3106 31703
rect 3214 31737 3266 31746
rect 3214 31703 3223 31737
rect 3223 31703 3257 31737
rect 3257 31703 3266 31737
rect 3214 31694 3266 31703
rect 3374 31737 3426 31746
rect 3374 31703 3383 31737
rect 3383 31703 3417 31737
rect 3417 31703 3426 31737
rect 3374 31694 3426 31703
rect 3534 31737 3586 31746
rect 3534 31703 3543 31737
rect 3543 31703 3577 31737
rect 3577 31703 3586 31737
rect 3534 31694 3586 31703
rect 3694 31737 3746 31746
rect 3694 31703 3703 31737
rect 3703 31703 3737 31737
rect 3737 31703 3746 31737
rect 3694 31694 3746 31703
rect 3854 31737 3906 31746
rect 3854 31703 3863 31737
rect 3863 31703 3897 31737
rect 3897 31703 3906 31737
rect 3854 31694 3906 31703
rect 4014 31737 4066 31746
rect 4014 31703 4023 31737
rect 4023 31703 4057 31737
rect 4057 31703 4066 31737
rect 4014 31694 4066 31703
rect 4174 31737 4226 31746
rect 4174 31703 4183 31737
rect 4183 31703 4217 31737
rect 4217 31703 4226 31737
rect 4174 31694 4226 31703
rect 4334 31737 4386 31746
rect 4334 31703 4343 31737
rect 4343 31703 4377 31737
rect 4377 31703 4386 31737
rect 4334 31694 4386 31703
rect 4494 31737 4546 31746
rect 4494 31703 4503 31737
rect 4503 31703 4537 31737
rect 4537 31703 4546 31737
rect 4494 31694 4546 31703
rect 4654 31737 4706 31746
rect 4654 31703 4663 31737
rect 4663 31703 4697 31737
rect 4697 31703 4706 31737
rect 4654 31694 4706 31703
rect 4814 31737 4866 31746
rect 4814 31703 4823 31737
rect 4823 31703 4857 31737
rect 4857 31703 4866 31737
rect 4814 31694 4866 31703
rect 4974 31737 5026 31746
rect 4974 31703 4983 31737
rect 4983 31703 5017 31737
rect 5017 31703 5026 31737
rect 4974 31694 5026 31703
rect 5134 31737 5186 31746
rect 5134 31703 5143 31737
rect 5143 31703 5177 31737
rect 5177 31703 5186 31737
rect 5134 31694 5186 31703
rect 5294 31737 5346 31746
rect 5294 31703 5303 31737
rect 5303 31703 5337 31737
rect 5337 31703 5346 31737
rect 5294 31694 5346 31703
rect 5454 31737 5506 31746
rect 5454 31703 5463 31737
rect 5463 31703 5497 31737
rect 5497 31703 5506 31737
rect 5454 31694 5506 31703
rect 5614 31737 5666 31746
rect 5614 31703 5623 31737
rect 5623 31703 5657 31737
rect 5657 31703 5666 31737
rect 5614 31694 5666 31703
rect 5774 31737 5826 31746
rect 5774 31703 5783 31737
rect 5783 31703 5817 31737
rect 5817 31703 5826 31737
rect 5774 31694 5826 31703
rect 5934 31737 5986 31746
rect 5934 31703 5943 31737
rect 5943 31703 5977 31737
rect 5977 31703 5986 31737
rect 5934 31694 5986 31703
rect 6094 31737 6146 31746
rect 6094 31703 6103 31737
rect 6103 31703 6137 31737
rect 6137 31703 6146 31737
rect 6094 31694 6146 31703
rect 6254 31737 6306 31746
rect 6254 31703 6263 31737
rect 6263 31703 6297 31737
rect 6297 31703 6306 31737
rect 6254 31694 6306 31703
rect 6414 31737 6466 31746
rect 6414 31703 6423 31737
rect 6423 31703 6457 31737
rect 6457 31703 6466 31737
rect 6414 31694 6466 31703
rect 6574 31737 6626 31746
rect 6574 31703 6583 31737
rect 6583 31703 6617 31737
rect 6617 31703 6626 31737
rect 6574 31694 6626 31703
rect 6734 31737 6786 31746
rect 6734 31703 6743 31737
rect 6743 31703 6777 31737
rect 6777 31703 6786 31737
rect 6734 31694 6786 31703
rect 6894 31737 6946 31746
rect 6894 31703 6903 31737
rect 6903 31703 6937 31737
rect 6937 31703 6946 31737
rect 6894 31694 6946 31703
rect 7054 31737 7106 31746
rect 7054 31703 7063 31737
rect 7063 31703 7097 31737
rect 7097 31703 7106 31737
rect 7054 31694 7106 31703
rect 7214 31737 7266 31746
rect 7214 31703 7223 31737
rect 7223 31703 7257 31737
rect 7257 31703 7266 31737
rect 7214 31694 7266 31703
rect 7374 31737 7426 31746
rect 7374 31703 7383 31737
rect 7383 31703 7417 31737
rect 7417 31703 7426 31737
rect 7374 31694 7426 31703
rect 7534 31737 7586 31746
rect 7534 31703 7543 31737
rect 7543 31703 7577 31737
rect 7577 31703 7586 31737
rect 7534 31694 7586 31703
rect 7694 31737 7746 31746
rect 7694 31703 7703 31737
rect 7703 31703 7737 31737
rect 7737 31703 7746 31737
rect 7694 31694 7746 31703
rect 7854 31737 7906 31746
rect 7854 31703 7863 31737
rect 7863 31703 7897 31737
rect 7897 31703 7906 31737
rect 7854 31694 7906 31703
rect 8014 31737 8066 31746
rect 8014 31703 8023 31737
rect 8023 31703 8057 31737
rect 8057 31703 8066 31737
rect 8014 31694 8066 31703
rect 8174 31737 8226 31746
rect 8174 31703 8183 31737
rect 8183 31703 8217 31737
rect 8217 31703 8226 31737
rect 8174 31694 8226 31703
rect 8334 31737 8386 31746
rect 8334 31703 8343 31737
rect 8343 31703 8377 31737
rect 8377 31703 8386 31737
rect 8334 31694 8386 31703
rect 12494 31737 12546 31746
rect 12494 31703 12503 31737
rect 12503 31703 12537 31737
rect 12537 31703 12546 31737
rect 12494 31694 12546 31703
rect 12654 31737 12706 31746
rect 12654 31703 12663 31737
rect 12663 31703 12697 31737
rect 12697 31703 12706 31737
rect 12654 31694 12706 31703
rect 12814 31737 12866 31746
rect 12814 31703 12823 31737
rect 12823 31703 12857 31737
rect 12857 31703 12866 31737
rect 12814 31694 12866 31703
rect 12974 31737 13026 31746
rect 12974 31703 12983 31737
rect 12983 31703 13017 31737
rect 13017 31703 13026 31737
rect 12974 31694 13026 31703
rect 13134 31737 13186 31746
rect 13134 31703 13143 31737
rect 13143 31703 13177 31737
rect 13177 31703 13186 31737
rect 13134 31694 13186 31703
rect 13294 31737 13346 31746
rect 13294 31703 13303 31737
rect 13303 31703 13337 31737
rect 13337 31703 13346 31737
rect 13294 31694 13346 31703
rect 13454 31737 13506 31746
rect 13454 31703 13463 31737
rect 13463 31703 13497 31737
rect 13497 31703 13506 31737
rect 13454 31694 13506 31703
rect 13614 31737 13666 31746
rect 13614 31703 13623 31737
rect 13623 31703 13657 31737
rect 13657 31703 13666 31737
rect 13614 31694 13666 31703
rect 13774 31737 13826 31746
rect 13774 31703 13783 31737
rect 13783 31703 13817 31737
rect 13817 31703 13826 31737
rect 13774 31694 13826 31703
rect 13934 31737 13986 31746
rect 13934 31703 13943 31737
rect 13943 31703 13977 31737
rect 13977 31703 13986 31737
rect 13934 31694 13986 31703
rect 14094 31737 14146 31746
rect 14094 31703 14103 31737
rect 14103 31703 14137 31737
rect 14137 31703 14146 31737
rect 14094 31694 14146 31703
rect 14254 31737 14306 31746
rect 14254 31703 14263 31737
rect 14263 31703 14297 31737
rect 14297 31703 14306 31737
rect 14254 31694 14306 31703
rect 14414 31737 14466 31746
rect 14414 31703 14423 31737
rect 14423 31703 14457 31737
rect 14457 31703 14466 31737
rect 14414 31694 14466 31703
rect 14574 31737 14626 31746
rect 14574 31703 14583 31737
rect 14583 31703 14617 31737
rect 14617 31703 14626 31737
rect 14574 31694 14626 31703
rect 14734 31737 14786 31746
rect 14734 31703 14743 31737
rect 14743 31703 14777 31737
rect 14777 31703 14786 31737
rect 14734 31694 14786 31703
rect 14894 31737 14946 31746
rect 14894 31703 14903 31737
rect 14903 31703 14937 31737
rect 14937 31703 14946 31737
rect 14894 31694 14946 31703
rect 15054 31737 15106 31746
rect 15054 31703 15063 31737
rect 15063 31703 15097 31737
rect 15097 31703 15106 31737
rect 15054 31694 15106 31703
rect 15214 31737 15266 31746
rect 15214 31703 15223 31737
rect 15223 31703 15257 31737
rect 15257 31703 15266 31737
rect 15214 31694 15266 31703
rect 15374 31737 15426 31746
rect 15374 31703 15383 31737
rect 15383 31703 15417 31737
rect 15417 31703 15426 31737
rect 15374 31694 15426 31703
rect 15534 31737 15586 31746
rect 15534 31703 15543 31737
rect 15543 31703 15577 31737
rect 15577 31703 15586 31737
rect 15534 31694 15586 31703
rect 15694 31737 15746 31746
rect 15694 31703 15703 31737
rect 15703 31703 15737 31737
rect 15737 31703 15746 31737
rect 15694 31694 15746 31703
rect 15854 31737 15906 31746
rect 15854 31703 15863 31737
rect 15863 31703 15897 31737
rect 15897 31703 15906 31737
rect 15854 31694 15906 31703
rect 16014 31737 16066 31746
rect 16014 31703 16023 31737
rect 16023 31703 16057 31737
rect 16057 31703 16066 31737
rect 16014 31694 16066 31703
rect 16174 31737 16226 31746
rect 16174 31703 16183 31737
rect 16183 31703 16217 31737
rect 16217 31703 16226 31737
rect 16174 31694 16226 31703
rect 16334 31737 16386 31746
rect 16334 31703 16343 31737
rect 16343 31703 16377 31737
rect 16377 31703 16386 31737
rect 16334 31694 16386 31703
rect 16494 31737 16546 31746
rect 16494 31703 16503 31737
rect 16503 31703 16537 31737
rect 16537 31703 16546 31737
rect 16494 31694 16546 31703
rect 16654 31737 16706 31746
rect 16654 31703 16663 31737
rect 16663 31703 16697 31737
rect 16697 31703 16706 31737
rect 16654 31694 16706 31703
rect 16814 31737 16866 31746
rect 16814 31703 16823 31737
rect 16823 31703 16857 31737
rect 16857 31703 16866 31737
rect 16814 31694 16866 31703
rect 16974 31737 17026 31746
rect 16974 31703 16983 31737
rect 16983 31703 17017 31737
rect 17017 31703 17026 31737
rect 16974 31694 17026 31703
rect 17134 31737 17186 31746
rect 17134 31703 17143 31737
rect 17143 31703 17177 31737
rect 17177 31703 17186 31737
rect 17134 31694 17186 31703
rect 17294 31737 17346 31746
rect 17294 31703 17303 31737
rect 17303 31703 17337 31737
rect 17337 31703 17346 31737
rect 17294 31694 17346 31703
rect 17454 31737 17506 31746
rect 17454 31703 17463 31737
rect 17463 31703 17497 31737
rect 17497 31703 17506 31737
rect 17454 31694 17506 31703
rect 17614 31737 17666 31746
rect 17614 31703 17623 31737
rect 17623 31703 17657 31737
rect 17657 31703 17666 31737
rect 17614 31694 17666 31703
rect 17774 31737 17826 31746
rect 17774 31703 17783 31737
rect 17783 31703 17817 31737
rect 17817 31703 17826 31737
rect 17774 31694 17826 31703
rect 17934 31737 17986 31746
rect 17934 31703 17943 31737
rect 17943 31703 17977 31737
rect 17977 31703 17986 31737
rect 17934 31694 17986 31703
rect 18094 31737 18146 31746
rect 18094 31703 18103 31737
rect 18103 31703 18137 31737
rect 18137 31703 18146 31737
rect 18094 31694 18146 31703
rect 18254 31737 18306 31746
rect 18254 31703 18263 31737
rect 18263 31703 18297 31737
rect 18297 31703 18306 31737
rect 18254 31694 18306 31703
rect 18414 31737 18466 31746
rect 18414 31703 18423 31737
rect 18423 31703 18457 31737
rect 18457 31703 18466 31737
rect 18414 31694 18466 31703
rect 18574 31737 18626 31746
rect 18574 31703 18583 31737
rect 18583 31703 18617 31737
rect 18617 31703 18626 31737
rect 18574 31694 18626 31703
rect 18734 31737 18786 31746
rect 18734 31703 18743 31737
rect 18743 31703 18777 31737
rect 18777 31703 18786 31737
rect 18734 31694 18786 31703
rect 18894 31737 18946 31746
rect 18894 31703 18903 31737
rect 18903 31703 18937 31737
rect 18937 31703 18946 31737
rect 18894 31694 18946 31703
rect 23134 31737 23186 31746
rect 23134 31703 23143 31737
rect 23143 31703 23177 31737
rect 23177 31703 23186 31737
rect 23134 31694 23186 31703
rect 23294 31737 23346 31746
rect 23294 31703 23303 31737
rect 23303 31703 23337 31737
rect 23337 31703 23346 31737
rect 23294 31694 23346 31703
rect 23454 31737 23506 31746
rect 23454 31703 23463 31737
rect 23463 31703 23497 31737
rect 23497 31703 23506 31737
rect 23454 31694 23506 31703
rect 23614 31737 23666 31746
rect 23614 31703 23623 31737
rect 23623 31703 23657 31737
rect 23657 31703 23666 31737
rect 23614 31694 23666 31703
rect 23774 31737 23826 31746
rect 23774 31703 23783 31737
rect 23783 31703 23817 31737
rect 23817 31703 23826 31737
rect 23774 31694 23826 31703
rect 23934 31737 23986 31746
rect 23934 31703 23943 31737
rect 23943 31703 23977 31737
rect 23977 31703 23986 31737
rect 23934 31694 23986 31703
rect 24094 31737 24146 31746
rect 24094 31703 24103 31737
rect 24103 31703 24137 31737
rect 24137 31703 24146 31737
rect 24094 31694 24146 31703
rect 24254 31737 24306 31746
rect 24254 31703 24263 31737
rect 24263 31703 24297 31737
rect 24297 31703 24306 31737
rect 24254 31694 24306 31703
rect 24414 31737 24466 31746
rect 24414 31703 24423 31737
rect 24423 31703 24457 31737
rect 24457 31703 24466 31737
rect 24414 31694 24466 31703
rect 24574 31737 24626 31746
rect 24574 31703 24583 31737
rect 24583 31703 24617 31737
rect 24617 31703 24626 31737
rect 24574 31694 24626 31703
rect 24734 31737 24786 31746
rect 24734 31703 24743 31737
rect 24743 31703 24777 31737
rect 24777 31703 24786 31737
rect 24734 31694 24786 31703
rect 24894 31737 24946 31746
rect 24894 31703 24903 31737
rect 24903 31703 24937 31737
rect 24937 31703 24946 31737
rect 24894 31694 24946 31703
rect 25054 31737 25106 31746
rect 25054 31703 25063 31737
rect 25063 31703 25097 31737
rect 25097 31703 25106 31737
rect 25054 31694 25106 31703
rect 25214 31737 25266 31746
rect 25214 31703 25223 31737
rect 25223 31703 25257 31737
rect 25257 31703 25266 31737
rect 25214 31694 25266 31703
rect 25374 31737 25426 31746
rect 25374 31703 25383 31737
rect 25383 31703 25417 31737
rect 25417 31703 25426 31737
rect 25374 31694 25426 31703
rect 25534 31737 25586 31746
rect 25534 31703 25543 31737
rect 25543 31703 25577 31737
rect 25577 31703 25586 31737
rect 25534 31694 25586 31703
rect 25694 31737 25746 31746
rect 25694 31703 25703 31737
rect 25703 31703 25737 31737
rect 25737 31703 25746 31737
rect 25694 31694 25746 31703
rect 25854 31737 25906 31746
rect 25854 31703 25863 31737
rect 25863 31703 25897 31737
rect 25897 31703 25906 31737
rect 25854 31694 25906 31703
rect 26014 31737 26066 31746
rect 26014 31703 26023 31737
rect 26023 31703 26057 31737
rect 26057 31703 26066 31737
rect 26014 31694 26066 31703
rect 26174 31737 26226 31746
rect 26174 31703 26183 31737
rect 26183 31703 26217 31737
rect 26217 31703 26226 31737
rect 26174 31694 26226 31703
rect 26334 31737 26386 31746
rect 26334 31703 26343 31737
rect 26343 31703 26377 31737
rect 26377 31703 26386 31737
rect 26334 31694 26386 31703
rect 26494 31737 26546 31746
rect 26494 31703 26503 31737
rect 26503 31703 26537 31737
rect 26537 31703 26546 31737
rect 26494 31694 26546 31703
rect 26654 31737 26706 31746
rect 26654 31703 26663 31737
rect 26663 31703 26697 31737
rect 26697 31703 26706 31737
rect 26654 31694 26706 31703
rect 26814 31737 26866 31746
rect 26814 31703 26823 31737
rect 26823 31703 26857 31737
rect 26857 31703 26866 31737
rect 26814 31694 26866 31703
rect 26974 31737 27026 31746
rect 26974 31703 26983 31737
rect 26983 31703 27017 31737
rect 27017 31703 27026 31737
rect 26974 31694 27026 31703
rect 27134 31737 27186 31746
rect 27134 31703 27143 31737
rect 27143 31703 27177 31737
rect 27177 31703 27186 31737
rect 27134 31694 27186 31703
rect 27294 31737 27346 31746
rect 27294 31703 27303 31737
rect 27303 31703 27337 31737
rect 27337 31703 27346 31737
rect 27294 31694 27346 31703
rect 27454 31737 27506 31746
rect 27454 31703 27463 31737
rect 27463 31703 27497 31737
rect 27497 31703 27506 31737
rect 27454 31694 27506 31703
rect 27614 31737 27666 31746
rect 27614 31703 27623 31737
rect 27623 31703 27657 31737
rect 27657 31703 27666 31737
rect 27614 31694 27666 31703
rect 27774 31737 27826 31746
rect 27774 31703 27783 31737
rect 27783 31703 27817 31737
rect 27817 31703 27826 31737
rect 27774 31694 27826 31703
rect 27934 31737 27986 31746
rect 27934 31703 27943 31737
rect 27943 31703 27977 31737
rect 27977 31703 27986 31737
rect 27934 31694 27986 31703
rect 28094 31737 28146 31746
rect 28094 31703 28103 31737
rect 28103 31703 28137 31737
rect 28137 31703 28146 31737
rect 28094 31694 28146 31703
rect 28254 31737 28306 31746
rect 28254 31703 28263 31737
rect 28263 31703 28297 31737
rect 28297 31703 28306 31737
rect 28254 31694 28306 31703
rect 28414 31737 28466 31746
rect 28414 31703 28423 31737
rect 28423 31703 28457 31737
rect 28457 31703 28466 31737
rect 28414 31694 28466 31703
rect 28574 31737 28626 31746
rect 28574 31703 28583 31737
rect 28583 31703 28617 31737
rect 28617 31703 28626 31737
rect 28574 31694 28626 31703
rect 28734 31737 28786 31746
rect 28734 31703 28743 31737
rect 28743 31703 28777 31737
rect 28777 31703 28786 31737
rect 28734 31694 28786 31703
rect 28894 31737 28946 31746
rect 28894 31703 28903 31737
rect 28903 31703 28937 31737
rect 28937 31703 28946 31737
rect 28894 31694 28946 31703
rect 29054 31737 29106 31746
rect 29054 31703 29063 31737
rect 29063 31703 29097 31737
rect 29097 31703 29106 31737
rect 29054 31694 29106 31703
rect 29214 31737 29266 31746
rect 29214 31703 29223 31737
rect 29223 31703 29257 31737
rect 29257 31703 29266 31737
rect 29214 31694 29266 31703
rect 29374 31737 29426 31746
rect 29374 31703 29383 31737
rect 29383 31703 29417 31737
rect 29417 31703 29426 31737
rect 29374 31694 29426 31703
rect 33534 31737 33586 31746
rect 33534 31703 33543 31737
rect 33543 31703 33577 31737
rect 33577 31703 33586 31737
rect 33534 31694 33586 31703
rect 33694 31737 33746 31746
rect 33694 31703 33703 31737
rect 33703 31703 33737 31737
rect 33737 31703 33746 31737
rect 33694 31694 33746 31703
rect 33854 31737 33906 31746
rect 33854 31703 33863 31737
rect 33863 31703 33897 31737
rect 33897 31703 33906 31737
rect 33854 31694 33906 31703
rect 34014 31737 34066 31746
rect 34014 31703 34023 31737
rect 34023 31703 34057 31737
rect 34057 31703 34066 31737
rect 34014 31694 34066 31703
rect 34174 31737 34226 31746
rect 34174 31703 34183 31737
rect 34183 31703 34217 31737
rect 34217 31703 34226 31737
rect 34174 31694 34226 31703
rect 34334 31737 34386 31746
rect 34334 31703 34343 31737
rect 34343 31703 34377 31737
rect 34377 31703 34386 31737
rect 34334 31694 34386 31703
rect 34494 31737 34546 31746
rect 34494 31703 34503 31737
rect 34503 31703 34537 31737
rect 34537 31703 34546 31737
rect 34494 31694 34546 31703
rect 34654 31737 34706 31746
rect 34654 31703 34663 31737
rect 34663 31703 34697 31737
rect 34697 31703 34706 31737
rect 34654 31694 34706 31703
rect 34814 31737 34866 31746
rect 34814 31703 34823 31737
rect 34823 31703 34857 31737
rect 34857 31703 34866 31737
rect 34814 31694 34866 31703
rect 34974 31737 35026 31746
rect 34974 31703 34983 31737
rect 34983 31703 35017 31737
rect 35017 31703 35026 31737
rect 34974 31694 35026 31703
rect 35134 31737 35186 31746
rect 35134 31703 35143 31737
rect 35143 31703 35177 31737
rect 35177 31703 35186 31737
rect 35134 31694 35186 31703
rect 35294 31737 35346 31746
rect 35294 31703 35303 31737
rect 35303 31703 35337 31737
rect 35337 31703 35346 31737
rect 35294 31694 35346 31703
rect 35454 31737 35506 31746
rect 35454 31703 35463 31737
rect 35463 31703 35497 31737
rect 35497 31703 35506 31737
rect 35454 31694 35506 31703
rect 35614 31737 35666 31746
rect 35614 31703 35623 31737
rect 35623 31703 35657 31737
rect 35657 31703 35666 31737
rect 35614 31694 35666 31703
rect 35774 31737 35826 31746
rect 35774 31703 35783 31737
rect 35783 31703 35817 31737
rect 35817 31703 35826 31737
rect 35774 31694 35826 31703
rect 35934 31737 35986 31746
rect 35934 31703 35943 31737
rect 35943 31703 35977 31737
rect 35977 31703 35986 31737
rect 35934 31694 35986 31703
rect 36094 31737 36146 31746
rect 36094 31703 36103 31737
rect 36103 31703 36137 31737
rect 36137 31703 36146 31737
rect 36094 31694 36146 31703
rect 36254 31737 36306 31746
rect 36254 31703 36263 31737
rect 36263 31703 36297 31737
rect 36297 31703 36306 31737
rect 36254 31694 36306 31703
rect 36414 31737 36466 31746
rect 36414 31703 36423 31737
rect 36423 31703 36457 31737
rect 36457 31703 36466 31737
rect 36414 31694 36466 31703
rect 36574 31737 36626 31746
rect 36574 31703 36583 31737
rect 36583 31703 36617 31737
rect 36617 31703 36626 31737
rect 36574 31694 36626 31703
rect 36734 31737 36786 31746
rect 36734 31703 36743 31737
rect 36743 31703 36777 31737
rect 36777 31703 36786 31737
rect 36734 31694 36786 31703
rect 36894 31737 36946 31746
rect 36894 31703 36903 31737
rect 36903 31703 36937 31737
rect 36937 31703 36946 31737
rect 36894 31694 36946 31703
rect 37054 31737 37106 31746
rect 37054 31703 37063 31737
rect 37063 31703 37097 31737
rect 37097 31703 37106 31737
rect 37054 31694 37106 31703
rect 37214 31737 37266 31746
rect 37214 31703 37223 31737
rect 37223 31703 37257 31737
rect 37257 31703 37266 31737
rect 37214 31694 37266 31703
rect 37374 31737 37426 31746
rect 37374 31703 37383 31737
rect 37383 31703 37417 31737
rect 37417 31703 37426 31737
rect 37374 31694 37426 31703
rect 37534 31737 37586 31746
rect 37534 31703 37543 31737
rect 37543 31703 37577 31737
rect 37577 31703 37586 31737
rect 37534 31694 37586 31703
rect 37694 31737 37746 31746
rect 37694 31703 37703 31737
rect 37703 31703 37737 31737
rect 37737 31703 37746 31737
rect 37694 31694 37746 31703
rect 37854 31737 37906 31746
rect 37854 31703 37863 31737
rect 37863 31703 37897 31737
rect 37897 31703 37906 31737
rect 37854 31694 37906 31703
rect 38014 31737 38066 31746
rect 38014 31703 38023 31737
rect 38023 31703 38057 31737
rect 38057 31703 38066 31737
rect 38014 31694 38066 31703
rect 38174 31737 38226 31746
rect 38174 31703 38183 31737
rect 38183 31703 38217 31737
rect 38217 31703 38226 31737
rect 38174 31694 38226 31703
rect 38334 31737 38386 31746
rect 38334 31703 38343 31737
rect 38343 31703 38377 31737
rect 38377 31703 38386 31737
rect 38334 31694 38386 31703
rect 38494 31737 38546 31746
rect 38494 31703 38503 31737
rect 38503 31703 38537 31737
rect 38537 31703 38546 31737
rect 38494 31694 38546 31703
rect 38654 31737 38706 31746
rect 38654 31703 38663 31737
rect 38663 31703 38697 31737
rect 38697 31703 38706 31737
rect 38654 31694 38706 31703
rect 38814 31737 38866 31746
rect 38814 31703 38823 31737
rect 38823 31703 38857 31737
rect 38857 31703 38866 31737
rect 38814 31694 38866 31703
rect 38974 31737 39026 31746
rect 38974 31703 38983 31737
rect 38983 31703 39017 31737
rect 39017 31703 39026 31737
rect 38974 31694 39026 31703
rect 39134 31737 39186 31746
rect 39134 31703 39143 31737
rect 39143 31703 39177 31737
rect 39177 31703 39186 31737
rect 39134 31694 39186 31703
rect 39294 31737 39346 31746
rect 39294 31703 39303 31737
rect 39303 31703 39337 31737
rect 39337 31703 39346 31737
rect 39294 31694 39346 31703
rect 39454 31737 39506 31746
rect 39454 31703 39463 31737
rect 39463 31703 39497 31737
rect 39497 31703 39506 31737
rect 39454 31694 39506 31703
rect 39614 31737 39666 31746
rect 39614 31703 39623 31737
rect 39623 31703 39657 31737
rect 39657 31703 39666 31737
rect 39614 31694 39666 31703
rect 39774 31737 39826 31746
rect 39774 31703 39783 31737
rect 39783 31703 39817 31737
rect 39817 31703 39826 31737
rect 39774 31694 39826 31703
rect 39934 31737 39986 31746
rect 39934 31703 39943 31737
rect 39943 31703 39977 31737
rect 39977 31703 39986 31737
rect 39934 31694 39986 31703
rect 40094 31737 40146 31746
rect 40094 31703 40103 31737
rect 40103 31703 40137 31737
rect 40137 31703 40146 31737
rect 40094 31694 40146 31703
rect 40254 31737 40306 31746
rect 40254 31703 40263 31737
rect 40263 31703 40297 31737
rect 40297 31703 40306 31737
rect 40254 31694 40306 31703
rect 40414 31737 40466 31746
rect 40414 31703 40423 31737
rect 40423 31703 40457 31737
rect 40457 31703 40466 31737
rect 40414 31694 40466 31703
rect 40574 31737 40626 31746
rect 40574 31703 40583 31737
rect 40583 31703 40617 31737
rect 40617 31703 40626 31737
rect 40574 31694 40626 31703
rect 40734 31737 40786 31746
rect 40734 31703 40743 31737
rect 40743 31703 40777 31737
rect 40777 31703 40786 31737
rect 40734 31694 40786 31703
rect 40894 31737 40946 31746
rect 40894 31703 40903 31737
rect 40903 31703 40937 31737
rect 40937 31703 40946 31737
rect 40894 31694 40946 31703
rect 41054 31737 41106 31746
rect 41054 31703 41063 31737
rect 41063 31703 41097 31737
rect 41097 31703 41106 31737
rect 41054 31694 41106 31703
rect 41214 31737 41266 31746
rect 41214 31703 41223 31737
rect 41223 31703 41257 31737
rect 41257 31703 41266 31737
rect 41214 31694 41266 31703
rect 41374 31737 41426 31746
rect 41374 31703 41383 31737
rect 41383 31703 41417 31737
rect 41417 31703 41426 31737
rect 41374 31694 41426 31703
rect 41534 31737 41586 31746
rect 41534 31703 41543 31737
rect 41543 31703 41577 31737
rect 41577 31703 41586 31737
rect 41534 31694 41586 31703
rect 41694 31737 41746 31746
rect 41694 31703 41703 31737
rect 41703 31703 41737 31737
rect 41737 31703 41746 31737
rect 41694 31694 41746 31703
rect 41854 31737 41906 31746
rect 41854 31703 41863 31737
rect 41863 31703 41897 31737
rect 41897 31703 41906 31737
rect 41854 31694 41906 31703
rect 14 31417 66 31426
rect 14 31383 23 31417
rect 23 31383 57 31417
rect 57 31383 66 31417
rect 14 31374 66 31383
rect 174 31417 226 31426
rect 174 31383 183 31417
rect 183 31383 217 31417
rect 217 31383 226 31417
rect 174 31374 226 31383
rect 334 31417 386 31426
rect 334 31383 343 31417
rect 343 31383 377 31417
rect 377 31383 386 31417
rect 334 31374 386 31383
rect 494 31417 546 31426
rect 494 31383 503 31417
rect 503 31383 537 31417
rect 537 31383 546 31417
rect 494 31374 546 31383
rect 654 31417 706 31426
rect 654 31383 663 31417
rect 663 31383 697 31417
rect 697 31383 706 31417
rect 654 31374 706 31383
rect 814 31417 866 31426
rect 814 31383 823 31417
rect 823 31383 857 31417
rect 857 31383 866 31417
rect 814 31374 866 31383
rect 974 31417 1026 31426
rect 974 31383 983 31417
rect 983 31383 1017 31417
rect 1017 31383 1026 31417
rect 974 31374 1026 31383
rect 1134 31417 1186 31426
rect 1134 31383 1143 31417
rect 1143 31383 1177 31417
rect 1177 31383 1186 31417
rect 1134 31374 1186 31383
rect 1294 31417 1346 31426
rect 1294 31383 1303 31417
rect 1303 31383 1337 31417
rect 1337 31383 1346 31417
rect 1294 31374 1346 31383
rect 1454 31417 1506 31426
rect 1454 31383 1463 31417
rect 1463 31383 1497 31417
rect 1497 31383 1506 31417
rect 1454 31374 1506 31383
rect 1614 31417 1666 31426
rect 1614 31383 1623 31417
rect 1623 31383 1657 31417
rect 1657 31383 1666 31417
rect 1614 31374 1666 31383
rect 1774 31417 1826 31426
rect 1774 31383 1783 31417
rect 1783 31383 1817 31417
rect 1817 31383 1826 31417
rect 1774 31374 1826 31383
rect 1934 31417 1986 31426
rect 1934 31383 1943 31417
rect 1943 31383 1977 31417
rect 1977 31383 1986 31417
rect 1934 31374 1986 31383
rect 2094 31417 2146 31426
rect 2094 31383 2103 31417
rect 2103 31383 2137 31417
rect 2137 31383 2146 31417
rect 2094 31374 2146 31383
rect 2254 31417 2306 31426
rect 2254 31383 2263 31417
rect 2263 31383 2297 31417
rect 2297 31383 2306 31417
rect 2254 31374 2306 31383
rect 2414 31417 2466 31426
rect 2414 31383 2423 31417
rect 2423 31383 2457 31417
rect 2457 31383 2466 31417
rect 2414 31374 2466 31383
rect 2574 31417 2626 31426
rect 2574 31383 2583 31417
rect 2583 31383 2617 31417
rect 2617 31383 2626 31417
rect 2574 31374 2626 31383
rect 2734 31417 2786 31426
rect 2734 31383 2743 31417
rect 2743 31383 2777 31417
rect 2777 31383 2786 31417
rect 2734 31374 2786 31383
rect 2894 31417 2946 31426
rect 2894 31383 2903 31417
rect 2903 31383 2937 31417
rect 2937 31383 2946 31417
rect 2894 31374 2946 31383
rect 3054 31417 3106 31426
rect 3054 31383 3063 31417
rect 3063 31383 3097 31417
rect 3097 31383 3106 31417
rect 3054 31374 3106 31383
rect 3214 31417 3266 31426
rect 3214 31383 3223 31417
rect 3223 31383 3257 31417
rect 3257 31383 3266 31417
rect 3214 31374 3266 31383
rect 3374 31417 3426 31426
rect 3374 31383 3383 31417
rect 3383 31383 3417 31417
rect 3417 31383 3426 31417
rect 3374 31374 3426 31383
rect 3534 31417 3586 31426
rect 3534 31383 3543 31417
rect 3543 31383 3577 31417
rect 3577 31383 3586 31417
rect 3534 31374 3586 31383
rect 3694 31417 3746 31426
rect 3694 31383 3703 31417
rect 3703 31383 3737 31417
rect 3737 31383 3746 31417
rect 3694 31374 3746 31383
rect 3854 31417 3906 31426
rect 3854 31383 3863 31417
rect 3863 31383 3897 31417
rect 3897 31383 3906 31417
rect 3854 31374 3906 31383
rect 4014 31417 4066 31426
rect 4014 31383 4023 31417
rect 4023 31383 4057 31417
rect 4057 31383 4066 31417
rect 4014 31374 4066 31383
rect 4174 31417 4226 31426
rect 4174 31383 4183 31417
rect 4183 31383 4217 31417
rect 4217 31383 4226 31417
rect 4174 31374 4226 31383
rect 4334 31417 4386 31426
rect 4334 31383 4343 31417
rect 4343 31383 4377 31417
rect 4377 31383 4386 31417
rect 4334 31374 4386 31383
rect 4494 31417 4546 31426
rect 4494 31383 4503 31417
rect 4503 31383 4537 31417
rect 4537 31383 4546 31417
rect 4494 31374 4546 31383
rect 4654 31417 4706 31426
rect 4654 31383 4663 31417
rect 4663 31383 4697 31417
rect 4697 31383 4706 31417
rect 4654 31374 4706 31383
rect 4814 31417 4866 31426
rect 4814 31383 4823 31417
rect 4823 31383 4857 31417
rect 4857 31383 4866 31417
rect 4814 31374 4866 31383
rect 4974 31417 5026 31426
rect 4974 31383 4983 31417
rect 4983 31383 5017 31417
rect 5017 31383 5026 31417
rect 4974 31374 5026 31383
rect 5134 31417 5186 31426
rect 5134 31383 5143 31417
rect 5143 31383 5177 31417
rect 5177 31383 5186 31417
rect 5134 31374 5186 31383
rect 5294 31417 5346 31426
rect 5294 31383 5303 31417
rect 5303 31383 5337 31417
rect 5337 31383 5346 31417
rect 5294 31374 5346 31383
rect 5454 31417 5506 31426
rect 5454 31383 5463 31417
rect 5463 31383 5497 31417
rect 5497 31383 5506 31417
rect 5454 31374 5506 31383
rect 5614 31417 5666 31426
rect 5614 31383 5623 31417
rect 5623 31383 5657 31417
rect 5657 31383 5666 31417
rect 5614 31374 5666 31383
rect 5774 31417 5826 31426
rect 5774 31383 5783 31417
rect 5783 31383 5817 31417
rect 5817 31383 5826 31417
rect 5774 31374 5826 31383
rect 5934 31417 5986 31426
rect 5934 31383 5943 31417
rect 5943 31383 5977 31417
rect 5977 31383 5986 31417
rect 5934 31374 5986 31383
rect 6094 31417 6146 31426
rect 6094 31383 6103 31417
rect 6103 31383 6137 31417
rect 6137 31383 6146 31417
rect 6094 31374 6146 31383
rect 6254 31417 6306 31426
rect 6254 31383 6263 31417
rect 6263 31383 6297 31417
rect 6297 31383 6306 31417
rect 6254 31374 6306 31383
rect 6414 31417 6466 31426
rect 6414 31383 6423 31417
rect 6423 31383 6457 31417
rect 6457 31383 6466 31417
rect 6414 31374 6466 31383
rect 6574 31417 6626 31426
rect 6574 31383 6583 31417
rect 6583 31383 6617 31417
rect 6617 31383 6626 31417
rect 6574 31374 6626 31383
rect 6734 31417 6786 31426
rect 6734 31383 6743 31417
rect 6743 31383 6777 31417
rect 6777 31383 6786 31417
rect 6734 31374 6786 31383
rect 6894 31417 6946 31426
rect 6894 31383 6903 31417
rect 6903 31383 6937 31417
rect 6937 31383 6946 31417
rect 6894 31374 6946 31383
rect 7054 31417 7106 31426
rect 7054 31383 7063 31417
rect 7063 31383 7097 31417
rect 7097 31383 7106 31417
rect 7054 31374 7106 31383
rect 7214 31417 7266 31426
rect 7214 31383 7223 31417
rect 7223 31383 7257 31417
rect 7257 31383 7266 31417
rect 7214 31374 7266 31383
rect 7374 31417 7426 31426
rect 7374 31383 7383 31417
rect 7383 31383 7417 31417
rect 7417 31383 7426 31417
rect 7374 31374 7426 31383
rect 7534 31417 7586 31426
rect 7534 31383 7543 31417
rect 7543 31383 7577 31417
rect 7577 31383 7586 31417
rect 7534 31374 7586 31383
rect 7694 31417 7746 31426
rect 7694 31383 7703 31417
rect 7703 31383 7737 31417
rect 7737 31383 7746 31417
rect 7694 31374 7746 31383
rect 7854 31417 7906 31426
rect 7854 31383 7863 31417
rect 7863 31383 7897 31417
rect 7897 31383 7906 31417
rect 7854 31374 7906 31383
rect 8014 31417 8066 31426
rect 8014 31383 8023 31417
rect 8023 31383 8057 31417
rect 8057 31383 8066 31417
rect 8014 31374 8066 31383
rect 8174 31417 8226 31426
rect 8174 31383 8183 31417
rect 8183 31383 8217 31417
rect 8217 31383 8226 31417
rect 8174 31374 8226 31383
rect 8334 31417 8386 31426
rect 8334 31383 8343 31417
rect 8343 31383 8377 31417
rect 8377 31383 8386 31417
rect 8334 31374 8386 31383
rect 12494 31417 12546 31426
rect 12494 31383 12503 31417
rect 12503 31383 12537 31417
rect 12537 31383 12546 31417
rect 12494 31374 12546 31383
rect 12654 31417 12706 31426
rect 12654 31383 12663 31417
rect 12663 31383 12697 31417
rect 12697 31383 12706 31417
rect 12654 31374 12706 31383
rect 12814 31417 12866 31426
rect 12814 31383 12823 31417
rect 12823 31383 12857 31417
rect 12857 31383 12866 31417
rect 12814 31374 12866 31383
rect 12974 31417 13026 31426
rect 12974 31383 12983 31417
rect 12983 31383 13017 31417
rect 13017 31383 13026 31417
rect 12974 31374 13026 31383
rect 13134 31417 13186 31426
rect 13134 31383 13143 31417
rect 13143 31383 13177 31417
rect 13177 31383 13186 31417
rect 13134 31374 13186 31383
rect 13294 31417 13346 31426
rect 13294 31383 13303 31417
rect 13303 31383 13337 31417
rect 13337 31383 13346 31417
rect 13294 31374 13346 31383
rect 13454 31417 13506 31426
rect 13454 31383 13463 31417
rect 13463 31383 13497 31417
rect 13497 31383 13506 31417
rect 13454 31374 13506 31383
rect 13614 31417 13666 31426
rect 13614 31383 13623 31417
rect 13623 31383 13657 31417
rect 13657 31383 13666 31417
rect 13614 31374 13666 31383
rect 13774 31417 13826 31426
rect 13774 31383 13783 31417
rect 13783 31383 13817 31417
rect 13817 31383 13826 31417
rect 13774 31374 13826 31383
rect 13934 31417 13986 31426
rect 13934 31383 13943 31417
rect 13943 31383 13977 31417
rect 13977 31383 13986 31417
rect 13934 31374 13986 31383
rect 14094 31417 14146 31426
rect 14094 31383 14103 31417
rect 14103 31383 14137 31417
rect 14137 31383 14146 31417
rect 14094 31374 14146 31383
rect 14254 31417 14306 31426
rect 14254 31383 14263 31417
rect 14263 31383 14297 31417
rect 14297 31383 14306 31417
rect 14254 31374 14306 31383
rect 14414 31417 14466 31426
rect 14414 31383 14423 31417
rect 14423 31383 14457 31417
rect 14457 31383 14466 31417
rect 14414 31374 14466 31383
rect 14574 31417 14626 31426
rect 14574 31383 14583 31417
rect 14583 31383 14617 31417
rect 14617 31383 14626 31417
rect 14574 31374 14626 31383
rect 14734 31417 14786 31426
rect 14734 31383 14743 31417
rect 14743 31383 14777 31417
rect 14777 31383 14786 31417
rect 14734 31374 14786 31383
rect 14894 31417 14946 31426
rect 14894 31383 14903 31417
rect 14903 31383 14937 31417
rect 14937 31383 14946 31417
rect 14894 31374 14946 31383
rect 15054 31417 15106 31426
rect 15054 31383 15063 31417
rect 15063 31383 15097 31417
rect 15097 31383 15106 31417
rect 15054 31374 15106 31383
rect 15214 31417 15266 31426
rect 15214 31383 15223 31417
rect 15223 31383 15257 31417
rect 15257 31383 15266 31417
rect 15214 31374 15266 31383
rect 15374 31417 15426 31426
rect 15374 31383 15383 31417
rect 15383 31383 15417 31417
rect 15417 31383 15426 31417
rect 15374 31374 15426 31383
rect 15534 31417 15586 31426
rect 15534 31383 15543 31417
rect 15543 31383 15577 31417
rect 15577 31383 15586 31417
rect 15534 31374 15586 31383
rect 15694 31417 15746 31426
rect 15694 31383 15703 31417
rect 15703 31383 15737 31417
rect 15737 31383 15746 31417
rect 15694 31374 15746 31383
rect 15854 31417 15906 31426
rect 15854 31383 15863 31417
rect 15863 31383 15897 31417
rect 15897 31383 15906 31417
rect 15854 31374 15906 31383
rect 16014 31417 16066 31426
rect 16014 31383 16023 31417
rect 16023 31383 16057 31417
rect 16057 31383 16066 31417
rect 16014 31374 16066 31383
rect 16174 31417 16226 31426
rect 16174 31383 16183 31417
rect 16183 31383 16217 31417
rect 16217 31383 16226 31417
rect 16174 31374 16226 31383
rect 16334 31417 16386 31426
rect 16334 31383 16343 31417
rect 16343 31383 16377 31417
rect 16377 31383 16386 31417
rect 16334 31374 16386 31383
rect 16494 31417 16546 31426
rect 16494 31383 16503 31417
rect 16503 31383 16537 31417
rect 16537 31383 16546 31417
rect 16494 31374 16546 31383
rect 16654 31417 16706 31426
rect 16654 31383 16663 31417
rect 16663 31383 16697 31417
rect 16697 31383 16706 31417
rect 16654 31374 16706 31383
rect 16814 31417 16866 31426
rect 16814 31383 16823 31417
rect 16823 31383 16857 31417
rect 16857 31383 16866 31417
rect 16814 31374 16866 31383
rect 16974 31417 17026 31426
rect 16974 31383 16983 31417
rect 16983 31383 17017 31417
rect 17017 31383 17026 31417
rect 16974 31374 17026 31383
rect 17134 31417 17186 31426
rect 17134 31383 17143 31417
rect 17143 31383 17177 31417
rect 17177 31383 17186 31417
rect 17134 31374 17186 31383
rect 17294 31417 17346 31426
rect 17294 31383 17303 31417
rect 17303 31383 17337 31417
rect 17337 31383 17346 31417
rect 17294 31374 17346 31383
rect 17454 31417 17506 31426
rect 17454 31383 17463 31417
rect 17463 31383 17497 31417
rect 17497 31383 17506 31417
rect 17454 31374 17506 31383
rect 17614 31417 17666 31426
rect 17614 31383 17623 31417
rect 17623 31383 17657 31417
rect 17657 31383 17666 31417
rect 17614 31374 17666 31383
rect 17774 31417 17826 31426
rect 17774 31383 17783 31417
rect 17783 31383 17817 31417
rect 17817 31383 17826 31417
rect 17774 31374 17826 31383
rect 17934 31417 17986 31426
rect 17934 31383 17943 31417
rect 17943 31383 17977 31417
rect 17977 31383 17986 31417
rect 17934 31374 17986 31383
rect 18094 31417 18146 31426
rect 18094 31383 18103 31417
rect 18103 31383 18137 31417
rect 18137 31383 18146 31417
rect 18094 31374 18146 31383
rect 18254 31417 18306 31426
rect 18254 31383 18263 31417
rect 18263 31383 18297 31417
rect 18297 31383 18306 31417
rect 18254 31374 18306 31383
rect 18414 31417 18466 31426
rect 18414 31383 18423 31417
rect 18423 31383 18457 31417
rect 18457 31383 18466 31417
rect 18414 31374 18466 31383
rect 18574 31417 18626 31426
rect 18574 31383 18583 31417
rect 18583 31383 18617 31417
rect 18617 31383 18626 31417
rect 18574 31374 18626 31383
rect 18734 31417 18786 31426
rect 18734 31383 18743 31417
rect 18743 31383 18777 31417
rect 18777 31383 18786 31417
rect 18734 31374 18786 31383
rect 18894 31417 18946 31426
rect 18894 31383 18903 31417
rect 18903 31383 18937 31417
rect 18937 31383 18946 31417
rect 18894 31374 18946 31383
rect 23134 31417 23186 31426
rect 23134 31383 23143 31417
rect 23143 31383 23177 31417
rect 23177 31383 23186 31417
rect 23134 31374 23186 31383
rect 23294 31417 23346 31426
rect 23294 31383 23303 31417
rect 23303 31383 23337 31417
rect 23337 31383 23346 31417
rect 23294 31374 23346 31383
rect 23454 31417 23506 31426
rect 23454 31383 23463 31417
rect 23463 31383 23497 31417
rect 23497 31383 23506 31417
rect 23454 31374 23506 31383
rect 23614 31417 23666 31426
rect 23614 31383 23623 31417
rect 23623 31383 23657 31417
rect 23657 31383 23666 31417
rect 23614 31374 23666 31383
rect 23774 31417 23826 31426
rect 23774 31383 23783 31417
rect 23783 31383 23817 31417
rect 23817 31383 23826 31417
rect 23774 31374 23826 31383
rect 23934 31417 23986 31426
rect 23934 31383 23943 31417
rect 23943 31383 23977 31417
rect 23977 31383 23986 31417
rect 23934 31374 23986 31383
rect 24094 31417 24146 31426
rect 24094 31383 24103 31417
rect 24103 31383 24137 31417
rect 24137 31383 24146 31417
rect 24094 31374 24146 31383
rect 24254 31417 24306 31426
rect 24254 31383 24263 31417
rect 24263 31383 24297 31417
rect 24297 31383 24306 31417
rect 24254 31374 24306 31383
rect 24414 31417 24466 31426
rect 24414 31383 24423 31417
rect 24423 31383 24457 31417
rect 24457 31383 24466 31417
rect 24414 31374 24466 31383
rect 24574 31417 24626 31426
rect 24574 31383 24583 31417
rect 24583 31383 24617 31417
rect 24617 31383 24626 31417
rect 24574 31374 24626 31383
rect 24734 31417 24786 31426
rect 24734 31383 24743 31417
rect 24743 31383 24777 31417
rect 24777 31383 24786 31417
rect 24734 31374 24786 31383
rect 24894 31417 24946 31426
rect 24894 31383 24903 31417
rect 24903 31383 24937 31417
rect 24937 31383 24946 31417
rect 24894 31374 24946 31383
rect 25054 31417 25106 31426
rect 25054 31383 25063 31417
rect 25063 31383 25097 31417
rect 25097 31383 25106 31417
rect 25054 31374 25106 31383
rect 25214 31417 25266 31426
rect 25214 31383 25223 31417
rect 25223 31383 25257 31417
rect 25257 31383 25266 31417
rect 25214 31374 25266 31383
rect 25374 31417 25426 31426
rect 25374 31383 25383 31417
rect 25383 31383 25417 31417
rect 25417 31383 25426 31417
rect 25374 31374 25426 31383
rect 25534 31417 25586 31426
rect 25534 31383 25543 31417
rect 25543 31383 25577 31417
rect 25577 31383 25586 31417
rect 25534 31374 25586 31383
rect 25694 31417 25746 31426
rect 25694 31383 25703 31417
rect 25703 31383 25737 31417
rect 25737 31383 25746 31417
rect 25694 31374 25746 31383
rect 25854 31417 25906 31426
rect 25854 31383 25863 31417
rect 25863 31383 25897 31417
rect 25897 31383 25906 31417
rect 25854 31374 25906 31383
rect 26014 31417 26066 31426
rect 26014 31383 26023 31417
rect 26023 31383 26057 31417
rect 26057 31383 26066 31417
rect 26014 31374 26066 31383
rect 26174 31417 26226 31426
rect 26174 31383 26183 31417
rect 26183 31383 26217 31417
rect 26217 31383 26226 31417
rect 26174 31374 26226 31383
rect 26334 31417 26386 31426
rect 26334 31383 26343 31417
rect 26343 31383 26377 31417
rect 26377 31383 26386 31417
rect 26334 31374 26386 31383
rect 26494 31417 26546 31426
rect 26494 31383 26503 31417
rect 26503 31383 26537 31417
rect 26537 31383 26546 31417
rect 26494 31374 26546 31383
rect 26654 31417 26706 31426
rect 26654 31383 26663 31417
rect 26663 31383 26697 31417
rect 26697 31383 26706 31417
rect 26654 31374 26706 31383
rect 26814 31417 26866 31426
rect 26814 31383 26823 31417
rect 26823 31383 26857 31417
rect 26857 31383 26866 31417
rect 26814 31374 26866 31383
rect 26974 31417 27026 31426
rect 26974 31383 26983 31417
rect 26983 31383 27017 31417
rect 27017 31383 27026 31417
rect 26974 31374 27026 31383
rect 27134 31417 27186 31426
rect 27134 31383 27143 31417
rect 27143 31383 27177 31417
rect 27177 31383 27186 31417
rect 27134 31374 27186 31383
rect 27294 31417 27346 31426
rect 27294 31383 27303 31417
rect 27303 31383 27337 31417
rect 27337 31383 27346 31417
rect 27294 31374 27346 31383
rect 27454 31417 27506 31426
rect 27454 31383 27463 31417
rect 27463 31383 27497 31417
rect 27497 31383 27506 31417
rect 27454 31374 27506 31383
rect 27614 31417 27666 31426
rect 27614 31383 27623 31417
rect 27623 31383 27657 31417
rect 27657 31383 27666 31417
rect 27614 31374 27666 31383
rect 27774 31417 27826 31426
rect 27774 31383 27783 31417
rect 27783 31383 27817 31417
rect 27817 31383 27826 31417
rect 27774 31374 27826 31383
rect 27934 31417 27986 31426
rect 27934 31383 27943 31417
rect 27943 31383 27977 31417
rect 27977 31383 27986 31417
rect 27934 31374 27986 31383
rect 28094 31417 28146 31426
rect 28094 31383 28103 31417
rect 28103 31383 28137 31417
rect 28137 31383 28146 31417
rect 28094 31374 28146 31383
rect 28254 31417 28306 31426
rect 28254 31383 28263 31417
rect 28263 31383 28297 31417
rect 28297 31383 28306 31417
rect 28254 31374 28306 31383
rect 28414 31417 28466 31426
rect 28414 31383 28423 31417
rect 28423 31383 28457 31417
rect 28457 31383 28466 31417
rect 28414 31374 28466 31383
rect 28574 31417 28626 31426
rect 28574 31383 28583 31417
rect 28583 31383 28617 31417
rect 28617 31383 28626 31417
rect 28574 31374 28626 31383
rect 28734 31417 28786 31426
rect 28734 31383 28743 31417
rect 28743 31383 28777 31417
rect 28777 31383 28786 31417
rect 28734 31374 28786 31383
rect 28894 31417 28946 31426
rect 28894 31383 28903 31417
rect 28903 31383 28937 31417
rect 28937 31383 28946 31417
rect 28894 31374 28946 31383
rect 29054 31417 29106 31426
rect 29054 31383 29063 31417
rect 29063 31383 29097 31417
rect 29097 31383 29106 31417
rect 29054 31374 29106 31383
rect 29214 31417 29266 31426
rect 29214 31383 29223 31417
rect 29223 31383 29257 31417
rect 29257 31383 29266 31417
rect 29214 31374 29266 31383
rect 29374 31417 29426 31426
rect 29374 31383 29383 31417
rect 29383 31383 29417 31417
rect 29417 31383 29426 31417
rect 29374 31374 29426 31383
rect 33534 31417 33586 31426
rect 33534 31383 33543 31417
rect 33543 31383 33577 31417
rect 33577 31383 33586 31417
rect 33534 31374 33586 31383
rect 33694 31417 33746 31426
rect 33694 31383 33703 31417
rect 33703 31383 33737 31417
rect 33737 31383 33746 31417
rect 33694 31374 33746 31383
rect 33854 31417 33906 31426
rect 33854 31383 33863 31417
rect 33863 31383 33897 31417
rect 33897 31383 33906 31417
rect 33854 31374 33906 31383
rect 34014 31417 34066 31426
rect 34014 31383 34023 31417
rect 34023 31383 34057 31417
rect 34057 31383 34066 31417
rect 34014 31374 34066 31383
rect 34174 31417 34226 31426
rect 34174 31383 34183 31417
rect 34183 31383 34217 31417
rect 34217 31383 34226 31417
rect 34174 31374 34226 31383
rect 34334 31417 34386 31426
rect 34334 31383 34343 31417
rect 34343 31383 34377 31417
rect 34377 31383 34386 31417
rect 34334 31374 34386 31383
rect 34494 31417 34546 31426
rect 34494 31383 34503 31417
rect 34503 31383 34537 31417
rect 34537 31383 34546 31417
rect 34494 31374 34546 31383
rect 34654 31417 34706 31426
rect 34654 31383 34663 31417
rect 34663 31383 34697 31417
rect 34697 31383 34706 31417
rect 34654 31374 34706 31383
rect 34814 31417 34866 31426
rect 34814 31383 34823 31417
rect 34823 31383 34857 31417
rect 34857 31383 34866 31417
rect 34814 31374 34866 31383
rect 34974 31417 35026 31426
rect 34974 31383 34983 31417
rect 34983 31383 35017 31417
rect 35017 31383 35026 31417
rect 34974 31374 35026 31383
rect 35134 31417 35186 31426
rect 35134 31383 35143 31417
rect 35143 31383 35177 31417
rect 35177 31383 35186 31417
rect 35134 31374 35186 31383
rect 35294 31417 35346 31426
rect 35294 31383 35303 31417
rect 35303 31383 35337 31417
rect 35337 31383 35346 31417
rect 35294 31374 35346 31383
rect 35454 31417 35506 31426
rect 35454 31383 35463 31417
rect 35463 31383 35497 31417
rect 35497 31383 35506 31417
rect 35454 31374 35506 31383
rect 35614 31417 35666 31426
rect 35614 31383 35623 31417
rect 35623 31383 35657 31417
rect 35657 31383 35666 31417
rect 35614 31374 35666 31383
rect 35774 31417 35826 31426
rect 35774 31383 35783 31417
rect 35783 31383 35817 31417
rect 35817 31383 35826 31417
rect 35774 31374 35826 31383
rect 35934 31417 35986 31426
rect 35934 31383 35943 31417
rect 35943 31383 35977 31417
rect 35977 31383 35986 31417
rect 35934 31374 35986 31383
rect 36094 31417 36146 31426
rect 36094 31383 36103 31417
rect 36103 31383 36137 31417
rect 36137 31383 36146 31417
rect 36094 31374 36146 31383
rect 36254 31417 36306 31426
rect 36254 31383 36263 31417
rect 36263 31383 36297 31417
rect 36297 31383 36306 31417
rect 36254 31374 36306 31383
rect 36414 31417 36466 31426
rect 36414 31383 36423 31417
rect 36423 31383 36457 31417
rect 36457 31383 36466 31417
rect 36414 31374 36466 31383
rect 36574 31417 36626 31426
rect 36574 31383 36583 31417
rect 36583 31383 36617 31417
rect 36617 31383 36626 31417
rect 36574 31374 36626 31383
rect 36734 31417 36786 31426
rect 36734 31383 36743 31417
rect 36743 31383 36777 31417
rect 36777 31383 36786 31417
rect 36734 31374 36786 31383
rect 36894 31417 36946 31426
rect 36894 31383 36903 31417
rect 36903 31383 36937 31417
rect 36937 31383 36946 31417
rect 36894 31374 36946 31383
rect 37054 31417 37106 31426
rect 37054 31383 37063 31417
rect 37063 31383 37097 31417
rect 37097 31383 37106 31417
rect 37054 31374 37106 31383
rect 37214 31417 37266 31426
rect 37214 31383 37223 31417
rect 37223 31383 37257 31417
rect 37257 31383 37266 31417
rect 37214 31374 37266 31383
rect 37374 31417 37426 31426
rect 37374 31383 37383 31417
rect 37383 31383 37417 31417
rect 37417 31383 37426 31417
rect 37374 31374 37426 31383
rect 37534 31417 37586 31426
rect 37534 31383 37543 31417
rect 37543 31383 37577 31417
rect 37577 31383 37586 31417
rect 37534 31374 37586 31383
rect 37694 31417 37746 31426
rect 37694 31383 37703 31417
rect 37703 31383 37737 31417
rect 37737 31383 37746 31417
rect 37694 31374 37746 31383
rect 37854 31417 37906 31426
rect 37854 31383 37863 31417
rect 37863 31383 37897 31417
rect 37897 31383 37906 31417
rect 37854 31374 37906 31383
rect 38014 31417 38066 31426
rect 38014 31383 38023 31417
rect 38023 31383 38057 31417
rect 38057 31383 38066 31417
rect 38014 31374 38066 31383
rect 38174 31417 38226 31426
rect 38174 31383 38183 31417
rect 38183 31383 38217 31417
rect 38217 31383 38226 31417
rect 38174 31374 38226 31383
rect 38334 31417 38386 31426
rect 38334 31383 38343 31417
rect 38343 31383 38377 31417
rect 38377 31383 38386 31417
rect 38334 31374 38386 31383
rect 38494 31417 38546 31426
rect 38494 31383 38503 31417
rect 38503 31383 38537 31417
rect 38537 31383 38546 31417
rect 38494 31374 38546 31383
rect 38654 31417 38706 31426
rect 38654 31383 38663 31417
rect 38663 31383 38697 31417
rect 38697 31383 38706 31417
rect 38654 31374 38706 31383
rect 38814 31417 38866 31426
rect 38814 31383 38823 31417
rect 38823 31383 38857 31417
rect 38857 31383 38866 31417
rect 38814 31374 38866 31383
rect 38974 31417 39026 31426
rect 38974 31383 38983 31417
rect 38983 31383 39017 31417
rect 39017 31383 39026 31417
rect 38974 31374 39026 31383
rect 39134 31417 39186 31426
rect 39134 31383 39143 31417
rect 39143 31383 39177 31417
rect 39177 31383 39186 31417
rect 39134 31374 39186 31383
rect 39294 31417 39346 31426
rect 39294 31383 39303 31417
rect 39303 31383 39337 31417
rect 39337 31383 39346 31417
rect 39294 31374 39346 31383
rect 39454 31417 39506 31426
rect 39454 31383 39463 31417
rect 39463 31383 39497 31417
rect 39497 31383 39506 31417
rect 39454 31374 39506 31383
rect 39614 31417 39666 31426
rect 39614 31383 39623 31417
rect 39623 31383 39657 31417
rect 39657 31383 39666 31417
rect 39614 31374 39666 31383
rect 39774 31417 39826 31426
rect 39774 31383 39783 31417
rect 39783 31383 39817 31417
rect 39817 31383 39826 31417
rect 39774 31374 39826 31383
rect 39934 31417 39986 31426
rect 39934 31383 39943 31417
rect 39943 31383 39977 31417
rect 39977 31383 39986 31417
rect 39934 31374 39986 31383
rect 40094 31417 40146 31426
rect 40094 31383 40103 31417
rect 40103 31383 40137 31417
rect 40137 31383 40146 31417
rect 40094 31374 40146 31383
rect 40254 31417 40306 31426
rect 40254 31383 40263 31417
rect 40263 31383 40297 31417
rect 40297 31383 40306 31417
rect 40254 31374 40306 31383
rect 40414 31417 40466 31426
rect 40414 31383 40423 31417
rect 40423 31383 40457 31417
rect 40457 31383 40466 31417
rect 40414 31374 40466 31383
rect 40574 31417 40626 31426
rect 40574 31383 40583 31417
rect 40583 31383 40617 31417
rect 40617 31383 40626 31417
rect 40574 31374 40626 31383
rect 40734 31417 40786 31426
rect 40734 31383 40743 31417
rect 40743 31383 40777 31417
rect 40777 31383 40786 31417
rect 40734 31374 40786 31383
rect 40894 31417 40946 31426
rect 40894 31383 40903 31417
rect 40903 31383 40937 31417
rect 40937 31383 40946 31417
rect 40894 31374 40946 31383
rect 41054 31417 41106 31426
rect 41054 31383 41063 31417
rect 41063 31383 41097 31417
rect 41097 31383 41106 31417
rect 41054 31374 41106 31383
rect 41214 31417 41266 31426
rect 41214 31383 41223 31417
rect 41223 31383 41257 31417
rect 41257 31383 41266 31417
rect 41214 31374 41266 31383
rect 41374 31417 41426 31426
rect 41374 31383 41383 31417
rect 41383 31383 41417 31417
rect 41417 31383 41426 31417
rect 41374 31374 41426 31383
rect 41534 31417 41586 31426
rect 41534 31383 41543 31417
rect 41543 31383 41577 31417
rect 41577 31383 41586 31417
rect 41534 31374 41586 31383
rect 41694 31417 41746 31426
rect 41694 31383 41703 31417
rect 41703 31383 41737 31417
rect 41737 31383 41746 31417
rect 41694 31374 41746 31383
rect 41854 31417 41906 31426
rect 41854 31383 41863 31417
rect 41863 31383 41897 31417
rect 41897 31383 41906 31417
rect 41854 31374 41906 31383
rect 14 31097 66 31106
rect 14 31063 23 31097
rect 23 31063 57 31097
rect 57 31063 66 31097
rect 14 31054 66 31063
rect 174 31097 226 31106
rect 174 31063 183 31097
rect 183 31063 217 31097
rect 217 31063 226 31097
rect 174 31054 226 31063
rect 334 31097 386 31106
rect 334 31063 343 31097
rect 343 31063 377 31097
rect 377 31063 386 31097
rect 334 31054 386 31063
rect 494 31097 546 31106
rect 494 31063 503 31097
rect 503 31063 537 31097
rect 537 31063 546 31097
rect 494 31054 546 31063
rect 654 31097 706 31106
rect 654 31063 663 31097
rect 663 31063 697 31097
rect 697 31063 706 31097
rect 654 31054 706 31063
rect 814 31097 866 31106
rect 814 31063 823 31097
rect 823 31063 857 31097
rect 857 31063 866 31097
rect 814 31054 866 31063
rect 974 31097 1026 31106
rect 974 31063 983 31097
rect 983 31063 1017 31097
rect 1017 31063 1026 31097
rect 974 31054 1026 31063
rect 1134 31097 1186 31106
rect 1134 31063 1143 31097
rect 1143 31063 1177 31097
rect 1177 31063 1186 31097
rect 1134 31054 1186 31063
rect 1294 31097 1346 31106
rect 1294 31063 1303 31097
rect 1303 31063 1337 31097
rect 1337 31063 1346 31097
rect 1294 31054 1346 31063
rect 1454 31097 1506 31106
rect 1454 31063 1463 31097
rect 1463 31063 1497 31097
rect 1497 31063 1506 31097
rect 1454 31054 1506 31063
rect 1614 31097 1666 31106
rect 1614 31063 1623 31097
rect 1623 31063 1657 31097
rect 1657 31063 1666 31097
rect 1614 31054 1666 31063
rect 1774 31097 1826 31106
rect 1774 31063 1783 31097
rect 1783 31063 1817 31097
rect 1817 31063 1826 31097
rect 1774 31054 1826 31063
rect 1934 31097 1986 31106
rect 1934 31063 1943 31097
rect 1943 31063 1977 31097
rect 1977 31063 1986 31097
rect 1934 31054 1986 31063
rect 2094 31097 2146 31106
rect 2094 31063 2103 31097
rect 2103 31063 2137 31097
rect 2137 31063 2146 31097
rect 2094 31054 2146 31063
rect 2254 31097 2306 31106
rect 2254 31063 2263 31097
rect 2263 31063 2297 31097
rect 2297 31063 2306 31097
rect 2254 31054 2306 31063
rect 2414 31097 2466 31106
rect 2414 31063 2423 31097
rect 2423 31063 2457 31097
rect 2457 31063 2466 31097
rect 2414 31054 2466 31063
rect 2574 31097 2626 31106
rect 2574 31063 2583 31097
rect 2583 31063 2617 31097
rect 2617 31063 2626 31097
rect 2574 31054 2626 31063
rect 2734 31097 2786 31106
rect 2734 31063 2743 31097
rect 2743 31063 2777 31097
rect 2777 31063 2786 31097
rect 2734 31054 2786 31063
rect 2894 31097 2946 31106
rect 2894 31063 2903 31097
rect 2903 31063 2937 31097
rect 2937 31063 2946 31097
rect 2894 31054 2946 31063
rect 3054 31097 3106 31106
rect 3054 31063 3063 31097
rect 3063 31063 3097 31097
rect 3097 31063 3106 31097
rect 3054 31054 3106 31063
rect 3214 31097 3266 31106
rect 3214 31063 3223 31097
rect 3223 31063 3257 31097
rect 3257 31063 3266 31097
rect 3214 31054 3266 31063
rect 3374 31097 3426 31106
rect 3374 31063 3383 31097
rect 3383 31063 3417 31097
rect 3417 31063 3426 31097
rect 3374 31054 3426 31063
rect 3534 31097 3586 31106
rect 3534 31063 3543 31097
rect 3543 31063 3577 31097
rect 3577 31063 3586 31097
rect 3534 31054 3586 31063
rect 3694 31097 3746 31106
rect 3694 31063 3703 31097
rect 3703 31063 3737 31097
rect 3737 31063 3746 31097
rect 3694 31054 3746 31063
rect 3854 31097 3906 31106
rect 3854 31063 3863 31097
rect 3863 31063 3897 31097
rect 3897 31063 3906 31097
rect 3854 31054 3906 31063
rect 4014 31097 4066 31106
rect 4014 31063 4023 31097
rect 4023 31063 4057 31097
rect 4057 31063 4066 31097
rect 4014 31054 4066 31063
rect 4174 31097 4226 31106
rect 4174 31063 4183 31097
rect 4183 31063 4217 31097
rect 4217 31063 4226 31097
rect 4174 31054 4226 31063
rect 4334 31097 4386 31106
rect 4334 31063 4343 31097
rect 4343 31063 4377 31097
rect 4377 31063 4386 31097
rect 4334 31054 4386 31063
rect 4494 31097 4546 31106
rect 4494 31063 4503 31097
rect 4503 31063 4537 31097
rect 4537 31063 4546 31097
rect 4494 31054 4546 31063
rect 4654 31097 4706 31106
rect 4654 31063 4663 31097
rect 4663 31063 4697 31097
rect 4697 31063 4706 31097
rect 4654 31054 4706 31063
rect 4814 31097 4866 31106
rect 4814 31063 4823 31097
rect 4823 31063 4857 31097
rect 4857 31063 4866 31097
rect 4814 31054 4866 31063
rect 4974 31097 5026 31106
rect 4974 31063 4983 31097
rect 4983 31063 5017 31097
rect 5017 31063 5026 31097
rect 4974 31054 5026 31063
rect 5134 31097 5186 31106
rect 5134 31063 5143 31097
rect 5143 31063 5177 31097
rect 5177 31063 5186 31097
rect 5134 31054 5186 31063
rect 5294 31097 5346 31106
rect 5294 31063 5303 31097
rect 5303 31063 5337 31097
rect 5337 31063 5346 31097
rect 5294 31054 5346 31063
rect 5454 31097 5506 31106
rect 5454 31063 5463 31097
rect 5463 31063 5497 31097
rect 5497 31063 5506 31097
rect 5454 31054 5506 31063
rect 5614 31097 5666 31106
rect 5614 31063 5623 31097
rect 5623 31063 5657 31097
rect 5657 31063 5666 31097
rect 5614 31054 5666 31063
rect 5774 31097 5826 31106
rect 5774 31063 5783 31097
rect 5783 31063 5817 31097
rect 5817 31063 5826 31097
rect 5774 31054 5826 31063
rect 5934 31097 5986 31106
rect 5934 31063 5943 31097
rect 5943 31063 5977 31097
rect 5977 31063 5986 31097
rect 5934 31054 5986 31063
rect 6094 31097 6146 31106
rect 6094 31063 6103 31097
rect 6103 31063 6137 31097
rect 6137 31063 6146 31097
rect 6094 31054 6146 31063
rect 6254 31097 6306 31106
rect 6254 31063 6263 31097
rect 6263 31063 6297 31097
rect 6297 31063 6306 31097
rect 6254 31054 6306 31063
rect 6414 31097 6466 31106
rect 6414 31063 6423 31097
rect 6423 31063 6457 31097
rect 6457 31063 6466 31097
rect 6414 31054 6466 31063
rect 6574 31097 6626 31106
rect 6574 31063 6583 31097
rect 6583 31063 6617 31097
rect 6617 31063 6626 31097
rect 6574 31054 6626 31063
rect 6734 31097 6786 31106
rect 6734 31063 6743 31097
rect 6743 31063 6777 31097
rect 6777 31063 6786 31097
rect 6734 31054 6786 31063
rect 6894 31097 6946 31106
rect 6894 31063 6903 31097
rect 6903 31063 6937 31097
rect 6937 31063 6946 31097
rect 6894 31054 6946 31063
rect 7054 31097 7106 31106
rect 7054 31063 7063 31097
rect 7063 31063 7097 31097
rect 7097 31063 7106 31097
rect 7054 31054 7106 31063
rect 7214 31097 7266 31106
rect 7214 31063 7223 31097
rect 7223 31063 7257 31097
rect 7257 31063 7266 31097
rect 7214 31054 7266 31063
rect 7374 31097 7426 31106
rect 7374 31063 7383 31097
rect 7383 31063 7417 31097
rect 7417 31063 7426 31097
rect 7374 31054 7426 31063
rect 7534 31097 7586 31106
rect 7534 31063 7543 31097
rect 7543 31063 7577 31097
rect 7577 31063 7586 31097
rect 7534 31054 7586 31063
rect 7694 31097 7746 31106
rect 7694 31063 7703 31097
rect 7703 31063 7737 31097
rect 7737 31063 7746 31097
rect 7694 31054 7746 31063
rect 7854 31097 7906 31106
rect 7854 31063 7863 31097
rect 7863 31063 7897 31097
rect 7897 31063 7906 31097
rect 7854 31054 7906 31063
rect 8014 31097 8066 31106
rect 8014 31063 8023 31097
rect 8023 31063 8057 31097
rect 8057 31063 8066 31097
rect 8014 31054 8066 31063
rect 8174 31097 8226 31106
rect 8174 31063 8183 31097
rect 8183 31063 8217 31097
rect 8217 31063 8226 31097
rect 8174 31054 8226 31063
rect 8334 31097 8386 31106
rect 8334 31063 8343 31097
rect 8343 31063 8377 31097
rect 8377 31063 8386 31097
rect 8334 31054 8386 31063
rect 12494 31097 12546 31106
rect 12494 31063 12503 31097
rect 12503 31063 12537 31097
rect 12537 31063 12546 31097
rect 12494 31054 12546 31063
rect 12654 31097 12706 31106
rect 12654 31063 12663 31097
rect 12663 31063 12697 31097
rect 12697 31063 12706 31097
rect 12654 31054 12706 31063
rect 12814 31097 12866 31106
rect 12814 31063 12823 31097
rect 12823 31063 12857 31097
rect 12857 31063 12866 31097
rect 12814 31054 12866 31063
rect 12974 31097 13026 31106
rect 12974 31063 12983 31097
rect 12983 31063 13017 31097
rect 13017 31063 13026 31097
rect 12974 31054 13026 31063
rect 13134 31097 13186 31106
rect 13134 31063 13143 31097
rect 13143 31063 13177 31097
rect 13177 31063 13186 31097
rect 13134 31054 13186 31063
rect 13294 31097 13346 31106
rect 13294 31063 13303 31097
rect 13303 31063 13337 31097
rect 13337 31063 13346 31097
rect 13294 31054 13346 31063
rect 13454 31097 13506 31106
rect 13454 31063 13463 31097
rect 13463 31063 13497 31097
rect 13497 31063 13506 31097
rect 13454 31054 13506 31063
rect 13614 31097 13666 31106
rect 13614 31063 13623 31097
rect 13623 31063 13657 31097
rect 13657 31063 13666 31097
rect 13614 31054 13666 31063
rect 13774 31097 13826 31106
rect 13774 31063 13783 31097
rect 13783 31063 13817 31097
rect 13817 31063 13826 31097
rect 13774 31054 13826 31063
rect 13934 31097 13986 31106
rect 13934 31063 13943 31097
rect 13943 31063 13977 31097
rect 13977 31063 13986 31097
rect 13934 31054 13986 31063
rect 14094 31097 14146 31106
rect 14094 31063 14103 31097
rect 14103 31063 14137 31097
rect 14137 31063 14146 31097
rect 14094 31054 14146 31063
rect 14254 31097 14306 31106
rect 14254 31063 14263 31097
rect 14263 31063 14297 31097
rect 14297 31063 14306 31097
rect 14254 31054 14306 31063
rect 14414 31097 14466 31106
rect 14414 31063 14423 31097
rect 14423 31063 14457 31097
rect 14457 31063 14466 31097
rect 14414 31054 14466 31063
rect 14574 31097 14626 31106
rect 14574 31063 14583 31097
rect 14583 31063 14617 31097
rect 14617 31063 14626 31097
rect 14574 31054 14626 31063
rect 14734 31097 14786 31106
rect 14734 31063 14743 31097
rect 14743 31063 14777 31097
rect 14777 31063 14786 31097
rect 14734 31054 14786 31063
rect 14894 31097 14946 31106
rect 14894 31063 14903 31097
rect 14903 31063 14937 31097
rect 14937 31063 14946 31097
rect 14894 31054 14946 31063
rect 15054 31097 15106 31106
rect 15054 31063 15063 31097
rect 15063 31063 15097 31097
rect 15097 31063 15106 31097
rect 15054 31054 15106 31063
rect 15214 31097 15266 31106
rect 15214 31063 15223 31097
rect 15223 31063 15257 31097
rect 15257 31063 15266 31097
rect 15214 31054 15266 31063
rect 15374 31097 15426 31106
rect 15374 31063 15383 31097
rect 15383 31063 15417 31097
rect 15417 31063 15426 31097
rect 15374 31054 15426 31063
rect 15534 31097 15586 31106
rect 15534 31063 15543 31097
rect 15543 31063 15577 31097
rect 15577 31063 15586 31097
rect 15534 31054 15586 31063
rect 15694 31097 15746 31106
rect 15694 31063 15703 31097
rect 15703 31063 15737 31097
rect 15737 31063 15746 31097
rect 15694 31054 15746 31063
rect 15854 31097 15906 31106
rect 15854 31063 15863 31097
rect 15863 31063 15897 31097
rect 15897 31063 15906 31097
rect 15854 31054 15906 31063
rect 16014 31097 16066 31106
rect 16014 31063 16023 31097
rect 16023 31063 16057 31097
rect 16057 31063 16066 31097
rect 16014 31054 16066 31063
rect 16174 31097 16226 31106
rect 16174 31063 16183 31097
rect 16183 31063 16217 31097
rect 16217 31063 16226 31097
rect 16174 31054 16226 31063
rect 16334 31097 16386 31106
rect 16334 31063 16343 31097
rect 16343 31063 16377 31097
rect 16377 31063 16386 31097
rect 16334 31054 16386 31063
rect 16494 31097 16546 31106
rect 16494 31063 16503 31097
rect 16503 31063 16537 31097
rect 16537 31063 16546 31097
rect 16494 31054 16546 31063
rect 16654 31097 16706 31106
rect 16654 31063 16663 31097
rect 16663 31063 16697 31097
rect 16697 31063 16706 31097
rect 16654 31054 16706 31063
rect 16814 31097 16866 31106
rect 16814 31063 16823 31097
rect 16823 31063 16857 31097
rect 16857 31063 16866 31097
rect 16814 31054 16866 31063
rect 16974 31097 17026 31106
rect 16974 31063 16983 31097
rect 16983 31063 17017 31097
rect 17017 31063 17026 31097
rect 16974 31054 17026 31063
rect 17134 31097 17186 31106
rect 17134 31063 17143 31097
rect 17143 31063 17177 31097
rect 17177 31063 17186 31097
rect 17134 31054 17186 31063
rect 17294 31097 17346 31106
rect 17294 31063 17303 31097
rect 17303 31063 17337 31097
rect 17337 31063 17346 31097
rect 17294 31054 17346 31063
rect 17454 31097 17506 31106
rect 17454 31063 17463 31097
rect 17463 31063 17497 31097
rect 17497 31063 17506 31097
rect 17454 31054 17506 31063
rect 17614 31097 17666 31106
rect 17614 31063 17623 31097
rect 17623 31063 17657 31097
rect 17657 31063 17666 31097
rect 17614 31054 17666 31063
rect 17774 31097 17826 31106
rect 17774 31063 17783 31097
rect 17783 31063 17817 31097
rect 17817 31063 17826 31097
rect 17774 31054 17826 31063
rect 17934 31097 17986 31106
rect 17934 31063 17943 31097
rect 17943 31063 17977 31097
rect 17977 31063 17986 31097
rect 17934 31054 17986 31063
rect 18094 31097 18146 31106
rect 18094 31063 18103 31097
rect 18103 31063 18137 31097
rect 18137 31063 18146 31097
rect 18094 31054 18146 31063
rect 18254 31097 18306 31106
rect 18254 31063 18263 31097
rect 18263 31063 18297 31097
rect 18297 31063 18306 31097
rect 18254 31054 18306 31063
rect 18414 31097 18466 31106
rect 18414 31063 18423 31097
rect 18423 31063 18457 31097
rect 18457 31063 18466 31097
rect 18414 31054 18466 31063
rect 18574 31097 18626 31106
rect 18574 31063 18583 31097
rect 18583 31063 18617 31097
rect 18617 31063 18626 31097
rect 18574 31054 18626 31063
rect 18734 31097 18786 31106
rect 18734 31063 18743 31097
rect 18743 31063 18777 31097
rect 18777 31063 18786 31097
rect 18734 31054 18786 31063
rect 18894 31097 18946 31106
rect 18894 31063 18903 31097
rect 18903 31063 18937 31097
rect 18937 31063 18946 31097
rect 18894 31054 18946 31063
rect 23134 31097 23186 31106
rect 23134 31063 23143 31097
rect 23143 31063 23177 31097
rect 23177 31063 23186 31097
rect 23134 31054 23186 31063
rect 23294 31097 23346 31106
rect 23294 31063 23303 31097
rect 23303 31063 23337 31097
rect 23337 31063 23346 31097
rect 23294 31054 23346 31063
rect 23454 31097 23506 31106
rect 23454 31063 23463 31097
rect 23463 31063 23497 31097
rect 23497 31063 23506 31097
rect 23454 31054 23506 31063
rect 23614 31097 23666 31106
rect 23614 31063 23623 31097
rect 23623 31063 23657 31097
rect 23657 31063 23666 31097
rect 23614 31054 23666 31063
rect 23774 31097 23826 31106
rect 23774 31063 23783 31097
rect 23783 31063 23817 31097
rect 23817 31063 23826 31097
rect 23774 31054 23826 31063
rect 23934 31097 23986 31106
rect 23934 31063 23943 31097
rect 23943 31063 23977 31097
rect 23977 31063 23986 31097
rect 23934 31054 23986 31063
rect 24094 31097 24146 31106
rect 24094 31063 24103 31097
rect 24103 31063 24137 31097
rect 24137 31063 24146 31097
rect 24094 31054 24146 31063
rect 24254 31097 24306 31106
rect 24254 31063 24263 31097
rect 24263 31063 24297 31097
rect 24297 31063 24306 31097
rect 24254 31054 24306 31063
rect 24414 31097 24466 31106
rect 24414 31063 24423 31097
rect 24423 31063 24457 31097
rect 24457 31063 24466 31097
rect 24414 31054 24466 31063
rect 24574 31097 24626 31106
rect 24574 31063 24583 31097
rect 24583 31063 24617 31097
rect 24617 31063 24626 31097
rect 24574 31054 24626 31063
rect 24734 31097 24786 31106
rect 24734 31063 24743 31097
rect 24743 31063 24777 31097
rect 24777 31063 24786 31097
rect 24734 31054 24786 31063
rect 24894 31097 24946 31106
rect 24894 31063 24903 31097
rect 24903 31063 24937 31097
rect 24937 31063 24946 31097
rect 24894 31054 24946 31063
rect 25054 31097 25106 31106
rect 25054 31063 25063 31097
rect 25063 31063 25097 31097
rect 25097 31063 25106 31097
rect 25054 31054 25106 31063
rect 25214 31097 25266 31106
rect 25214 31063 25223 31097
rect 25223 31063 25257 31097
rect 25257 31063 25266 31097
rect 25214 31054 25266 31063
rect 25374 31097 25426 31106
rect 25374 31063 25383 31097
rect 25383 31063 25417 31097
rect 25417 31063 25426 31097
rect 25374 31054 25426 31063
rect 25534 31097 25586 31106
rect 25534 31063 25543 31097
rect 25543 31063 25577 31097
rect 25577 31063 25586 31097
rect 25534 31054 25586 31063
rect 25694 31097 25746 31106
rect 25694 31063 25703 31097
rect 25703 31063 25737 31097
rect 25737 31063 25746 31097
rect 25694 31054 25746 31063
rect 25854 31097 25906 31106
rect 25854 31063 25863 31097
rect 25863 31063 25897 31097
rect 25897 31063 25906 31097
rect 25854 31054 25906 31063
rect 26014 31097 26066 31106
rect 26014 31063 26023 31097
rect 26023 31063 26057 31097
rect 26057 31063 26066 31097
rect 26014 31054 26066 31063
rect 26174 31097 26226 31106
rect 26174 31063 26183 31097
rect 26183 31063 26217 31097
rect 26217 31063 26226 31097
rect 26174 31054 26226 31063
rect 26334 31097 26386 31106
rect 26334 31063 26343 31097
rect 26343 31063 26377 31097
rect 26377 31063 26386 31097
rect 26334 31054 26386 31063
rect 26494 31097 26546 31106
rect 26494 31063 26503 31097
rect 26503 31063 26537 31097
rect 26537 31063 26546 31097
rect 26494 31054 26546 31063
rect 26654 31097 26706 31106
rect 26654 31063 26663 31097
rect 26663 31063 26697 31097
rect 26697 31063 26706 31097
rect 26654 31054 26706 31063
rect 26814 31097 26866 31106
rect 26814 31063 26823 31097
rect 26823 31063 26857 31097
rect 26857 31063 26866 31097
rect 26814 31054 26866 31063
rect 26974 31097 27026 31106
rect 26974 31063 26983 31097
rect 26983 31063 27017 31097
rect 27017 31063 27026 31097
rect 26974 31054 27026 31063
rect 27134 31097 27186 31106
rect 27134 31063 27143 31097
rect 27143 31063 27177 31097
rect 27177 31063 27186 31097
rect 27134 31054 27186 31063
rect 27294 31097 27346 31106
rect 27294 31063 27303 31097
rect 27303 31063 27337 31097
rect 27337 31063 27346 31097
rect 27294 31054 27346 31063
rect 27454 31097 27506 31106
rect 27454 31063 27463 31097
rect 27463 31063 27497 31097
rect 27497 31063 27506 31097
rect 27454 31054 27506 31063
rect 27614 31097 27666 31106
rect 27614 31063 27623 31097
rect 27623 31063 27657 31097
rect 27657 31063 27666 31097
rect 27614 31054 27666 31063
rect 27774 31097 27826 31106
rect 27774 31063 27783 31097
rect 27783 31063 27817 31097
rect 27817 31063 27826 31097
rect 27774 31054 27826 31063
rect 27934 31097 27986 31106
rect 27934 31063 27943 31097
rect 27943 31063 27977 31097
rect 27977 31063 27986 31097
rect 27934 31054 27986 31063
rect 28094 31097 28146 31106
rect 28094 31063 28103 31097
rect 28103 31063 28137 31097
rect 28137 31063 28146 31097
rect 28094 31054 28146 31063
rect 28254 31097 28306 31106
rect 28254 31063 28263 31097
rect 28263 31063 28297 31097
rect 28297 31063 28306 31097
rect 28254 31054 28306 31063
rect 28414 31097 28466 31106
rect 28414 31063 28423 31097
rect 28423 31063 28457 31097
rect 28457 31063 28466 31097
rect 28414 31054 28466 31063
rect 28574 31097 28626 31106
rect 28574 31063 28583 31097
rect 28583 31063 28617 31097
rect 28617 31063 28626 31097
rect 28574 31054 28626 31063
rect 28734 31097 28786 31106
rect 28734 31063 28743 31097
rect 28743 31063 28777 31097
rect 28777 31063 28786 31097
rect 28734 31054 28786 31063
rect 28894 31097 28946 31106
rect 28894 31063 28903 31097
rect 28903 31063 28937 31097
rect 28937 31063 28946 31097
rect 28894 31054 28946 31063
rect 29054 31097 29106 31106
rect 29054 31063 29063 31097
rect 29063 31063 29097 31097
rect 29097 31063 29106 31097
rect 29054 31054 29106 31063
rect 29214 31097 29266 31106
rect 29214 31063 29223 31097
rect 29223 31063 29257 31097
rect 29257 31063 29266 31097
rect 29214 31054 29266 31063
rect 29374 31097 29426 31106
rect 29374 31063 29383 31097
rect 29383 31063 29417 31097
rect 29417 31063 29426 31097
rect 29374 31054 29426 31063
rect 33534 31097 33586 31106
rect 33534 31063 33543 31097
rect 33543 31063 33577 31097
rect 33577 31063 33586 31097
rect 33534 31054 33586 31063
rect 33694 31097 33746 31106
rect 33694 31063 33703 31097
rect 33703 31063 33737 31097
rect 33737 31063 33746 31097
rect 33694 31054 33746 31063
rect 33854 31097 33906 31106
rect 33854 31063 33863 31097
rect 33863 31063 33897 31097
rect 33897 31063 33906 31097
rect 33854 31054 33906 31063
rect 34014 31097 34066 31106
rect 34014 31063 34023 31097
rect 34023 31063 34057 31097
rect 34057 31063 34066 31097
rect 34014 31054 34066 31063
rect 34174 31097 34226 31106
rect 34174 31063 34183 31097
rect 34183 31063 34217 31097
rect 34217 31063 34226 31097
rect 34174 31054 34226 31063
rect 34334 31097 34386 31106
rect 34334 31063 34343 31097
rect 34343 31063 34377 31097
rect 34377 31063 34386 31097
rect 34334 31054 34386 31063
rect 34494 31097 34546 31106
rect 34494 31063 34503 31097
rect 34503 31063 34537 31097
rect 34537 31063 34546 31097
rect 34494 31054 34546 31063
rect 34654 31097 34706 31106
rect 34654 31063 34663 31097
rect 34663 31063 34697 31097
rect 34697 31063 34706 31097
rect 34654 31054 34706 31063
rect 34814 31097 34866 31106
rect 34814 31063 34823 31097
rect 34823 31063 34857 31097
rect 34857 31063 34866 31097
rect 34814 31054 34866 31063
rect 34974 31097 35026 31106
rect 34974 31063 34983 31097
rect 34983 31063 35017 31097
rect 35017 31063 35026 31097
rect 34974 31054 35026 31063
rect 35134 31097 35186 31106
rect 35134 31063 35143 31097
rect 35143 31063 35177 31097
rect 35177 31063 35186 31097
rect 35134 31054 35186 31063
rect 35294 31097 35346 31106
rect 35294 31063 35303 31097
rect 35303 31063 35337 31097
rect 35337 31063 35346 31097
rect 35294 31054 35346 31063
rect 35454 31097 35506 31106
rect 35454 31063 35463 31097
rect 35463 31063 35497 31097
rect 35497 31063 35506 31097
rect 35454 31054 35506 31063
rect 35614 31097 35666 31106
rect 35614 31063 35623 31097
rect 35623 31063 35657 31097
rect 35657 31063 35666 31097
rect 35614 31054 35666 31063
rect 35774 31097 35826 31106
rect 35774 31063 35783 31097
rect 35783 31063 35817 31097
rect 35817 31063 35826 31097
rect 35774 31054 35826 31063
rect 35934 31097 35986 31106
rect 35934 31063 35943 31097
rect 35943 31063 35977 31097
rect 35977 31063 35986 31097
rect 35934 31054 35986 31063
rect 36094 31097 36146 31106
rect 36094 31063 36103 31097
rect 36103 31063 36137 31097
rect 36137 31063 36146 31097
rect 36094 31054 36146 31063
rect 36254 31097 36306 31106
rect 36254 31063 36263 31097
rect 36263 31063 36297 31097
rect 36297 31063 36306 31097
rect 36254 31054 36306 31063
rect 36414 31097 36466 31106
rect 36414 31063 36423 31097
rect 36423 31063 36457 31097
rect 36457 31063 36466 31097
rect 36414 31054 36466 31063
rect 36574 31097 36626 31106
rect 36574 31063 36583 31097
rect 36583 31063 36617 31097
rect 36617 31063 36626 31097
rect 36574 31054 36626 31063
rect 36734 31097 36786 31106
rect 36734 31063 36743 31097
rect 36743 31063 36777 31097
rect 36777 31063 36786 31097
rect 36734 31054 36786 31063
rect 36894 31097 36946 31106
rect 36894 31063 36903 31097
rect 36903 31063 36937 31097
rect 36937 31063 36946 31097
rect 36894 31054 36946 31063
rect 37054 31097 37106 31106
rect 37054 31063 37063 31097
rect 37063 31063 37097 31097
rect 37097 31063 37106 31097
rect 37054 31054 37106 31063
rect 37214 31097 37266 31106
rect 37214 31063 37223 31097
rect 37223 31063 37257 31097
rect 37257 31063 37266 31097
rect 37214 31054 37266 31063
rect 37374 31097 37426 31106
rect 37374 31063 37383 31097
rect 37383 31063 37417 31097
rect 37417 31063 37426 31097
rect 37374 31054 37426 31063
rect 37534 31097 37586 31106
rect 37534 31063 37543 31097
rect 37543 31063 37577 31097
rect 37577 31063 37586 31097
rect 37534 31054 37586 31063
rect 37694 31097 37746 31106
rect 37694 31063 37703 31097
rect 37703 31063 37737 31097
rect 37737 31063 37746 31097
rect 37694 31054 37746 31063
rect 37854 31097 37906 31106
rect 37854 31063 37863 31097
rect 37863 31063 37897 31097
rect 37897 31063 37906 31097
rect 37854 31054 37906 31063
rect 38014 31097 38066 31106
rect 38014 31063 38023 31097
rect 38023 31063 38057 31097
rect 38057 31063 38066 31097
rect 38014 31054 38066 31063
rect 38174 31097 38226 31106
rect 38174 31063 38183 31097
rect 38183 31063 38217 31097
rect 38217 31063 38226 31097
rect 38174 31054 38226 31063
rect 38334 31097 38386 31106
rect 38334 31063 38343 31097
rect 38343 31063 38377 31097
rect 38377 31063 38386 31097
rect 38334 31054 38386 31063
rect 38494 31097 38546 31106
rect 38494 31063 38503 31097
rect 38503 31063 38537 31097
rect 38537 31063 38546 31097
rect 38494 31054 38546 31063
rect 38654 31097 38706 31106
rect 38654 31063 38663 31097
rect 38663 31063 38697 31097
rect 38697 31063 38706 31097
rect 38654 31054 38706 31063
rect 38814 31097 38866 31106
rect 38814 31063 38823 31097
rect 38823 31063 38857 31097
rect 38857 31063 38866 31097
rect 38814 31054 38866 31063
rect 38974 31097 39026 31106
rect 38974 31063 38983 31097
rect 38983 31063 39017 31097
rect 39017 31063 39026 31097
rect 38974 31054 39026 31063
rect 39134 31097 39186 31106
rect 39134 31063 39143 31097
rect 39143 31063 39177 31097
rect 39177 31063 39186 31097
rect 39134 31054 39186 31063
rect 39294 31097 39346 31106
rect 39294 31063 39303 31097
rect 39303 31063 39337 31097
rect 39337 31063 39346 31097
rect 39294 31054 39346 31063
rect 39454 31097 39506 31106
rect 39454 31063 39463 31097
rect 39463 31063 39497 31097
rect 39497 31063 39506 31097
rect 39454 31054 39506 31063
rect 39614 31097 39666 31106
rect 39614 31063 39623 31097
rect 39623 31063 39657 31097
rect 39657 31063 39666 31097
rect 39614 31054 39666 31063
rect 39774 31097 39826 31106
rect 39774 31063 39783 31097
rect 39783 31063 39817 31097
rect 39817 31063 39826 31097
rect 39774 31054 39826 31063
rect 39934 31097 39986 31106
rect 39934 31063 39943 31097
rect 39943 31063 39977 31097
rect 39977 31063 39986 31097
rect 39934 31054 39986 31063
rect 40094 31097 40146 31106
rect 40094 31063 40103 31097
rect 40103 31063 40137 31097
rect 40137 31063 40146 31097
rect 40094 31054 40146 31063
rect 40254 31097 40306 31106
rect 40254 31063 40263 31097
rect 40263 31063 40297 31097
rect 40297 31063 40306 31097
rect 40254 31054 40306 31063
rect 40414 31097 40466 31106
rect 40414 31063 40423 31097
rect 40423 31063 40457 31097
rect 40457 31063 40466 31097
rect 40414 31054 40466 31063
rect 40574 31097 40626 31106
rect 40574 31063 40583 31097
rect 40583 31063 40617 31097
rect 40617 31063 40626 31097
rect 40574 31054 40626 31063
rect 40734 31097 40786 31106
rect 40734 31063 40743 31097
rect 40743 31063 40777 31097
rect 40777 31063 40786 31097
rect 40734 31054 40786 31063
rect 40894 31097 40946 31106
rect 40894 31063 40903 31097
rect 40903 31063 40937 31097
rect 40937 31063 40946 31097
rect 40894 31054 40946 31063
rect 41054 31097 41106 31106
rect 41054 31063 41063 31097
rect 41063 31063 41097 31097
rect 41097 31063 41106 31097
rect 41054 31054 41106 31063
rect 41214 31097 41266 31106
rect 41214 31063 41223 31097
rect 41223 31063 41257 31097
rect 41257 31063 41266 31097
rect 41214 31054 41266 31063
rect 41374 31097 41426 31106
rect 41374 31063 41383 31097
rect 41383 31063 41417 31097
rect 41417 31063 41426 31097
rect 41374 31054 41426 31063
rect 41534 31097 41586 31106
rect 41534 31063 41543 31097
rect 41543 31063 41577 31097
rect 41577 31063 41586 31097
rect 41534 31054 41586 31063
rect 41694 31097 41746 31106
rect 41694 31063 41703 31097
rect 41703 31063 41737 31097
rect 41737 31063 41746 31097
rect 41694 31054 41746 31063
rect 41854 31097 41906 31106
rect 41854 31063 41863 31097
rect 41863 31063 41897 31097
rect 41897 31063 41906 31097
rect 41854 31054 41906 31063
rect 14 30777 66 30786
rect 14 30743 23 30777
rect 23 30743 57 30777
rect 57 30743 66 30777
rect 14 30734 66 30743
rect 174 30777 226 30786
rect 174 30743 183 30777
rect 183 30743 217 30777
rect 217 30743 226 30777
rect 174 30734 226 30743
rect 334 30777 386 30786
rect 334 30743 343 30777
rect 343 30743 377 30777
rect 377 30743 386 30777
rect 334 30734 386 30743
rect 494 30777 546 30786
rect 494 30743 503 30777
rect 503 30743 537 30777
rect 537 30743 546 30777
rect 494 30734 546 30743
rect 654 30777 706 30786
rect 654 30743 663 30777
rect 663 30743 697 30777
rect 697 30743 706 30777
rect 654 30734 706 30743
rect 814 30777 866 30786
rect 814 30743 823 30777
rect 823 30743 857 30777
rect 857 30743 866 30777
rect 814 30734 866 30743
rect 974 30777 1026 30786
rect 974 30743 983 30777
rect 983 30743 1017 30777
rect 1017 30743 1026 30777
rect 974 30734 1026 30743
rect 1134 30777 1186 30786
rect 1134 30743 1143 30777
rect 1143 30743 1177 30777
rect 1177 30743 1186 30777
rect 1134 30734 1186 30743
rect 1294 30777 1346 30786
rect 1294 30743 1303 30777
rect 1303 30743 1337 30777
rect 1337 30743 1346 30777
rect 1294 30734 1346 30743
rect 1454 30777 1506 30786
rect 1454 30743 1463 30777
rect 1463 30743 1497 30777
rect 1497 30743 1506 30777
rect 1454 30734 1506 30743
rect 1614 30777 1666 30786
rect 1614 30743 1623 30777
rect 1623 30743 1657 30777
rect 1657 30743 1666 30777
rect 1614 30734 1666 30743
rect 1774 30777 1826 30786
rect 1774 30743 1783 30777
rect 1783 30743 1817 30777
rect 1817 30743 1826 30777
rect 1774 30734 1826 30743
rect 1934 30777 1986 30786
rect 1934 30743 1943 30777
rect 1943 30743 1977 30777
rect 1977 30743 1986 30777
rect 1934 30734 1986 30743
rect 2094 30777 2146 30786
rect 2094 30743 2103 30777
rect 2103 30743 2137 30777
rect 2137 30743 2146 30777
rect 2094 30734 2146 30743
rect 2254 30777 2306 30786
rect 2254 30743 2263 30777
rect 2263 30743 2297 30777
rect 2297 30743 2306 30777
rect 2254 30734 2306 30743
rect 2414 30777 2466 30786
rect 2414 30743 2423 30777
rect 2423 30743 2457 30777
rect 2457 30743 2466 30777
rect 2414 30734 2466 30743
rect 2574 30777 2626 30786
rect 2574 30743 2583 30777
rect 2583 30743 2617 30777
rect 2617 30743 2626 30777
rect 2574 30734 2626 30743
rect 2734 30777 2786 30786
rect 2734 30743 2743 30777
rect 2743 30743 2777 30777
rect 2777 30743 2786 30777
rect 2734 30734 2786 30743
rect 2894 30777 2946 30786
rect 2894 30743 2903 30777
rect 2903 30743 2937 30777
rect 2937 30743 2946 30777
rect 2894 30734 2946 30743
rect 3054 30777 3106 30786
rect 3054 30743 3063 30777
rect 3063 30743 3097 30777
rect 3097 30743 3106 30777
rect 3054 30734 3106 30743
rect 3214 30777 3266 30786
rect 3214 30743 3223 30777
rect 3223 30743 3257 30777
rect 3257 30743 3266 30777
rect 3214 30734 3266 30743
rect 3374 30777 3426 30786
rect 3374 30743 3383 30777
rect 3383 30743 3417 30777
rect 3417 30743 3426 30777
rect 3374 30734 3426 30743
rect 3534 30777 3586 30786
rect 3534 30743 3543 30777
rect 3543 30743 3577 30777
rect 3577 30743 3586 30777
rect 3534 30734 3586 30743
rect 3694 30777 3746 30786
rect 3694 30743 3703 30777
rect 3703 30743 3737 30777
rect 3737 30743 3746 30777
rect 3694 30734 3746 30743
rect 3854 30777 3906 30786
rect 3854 30743 3863 30777
rect 3863 30743 3897 30777
rect 3897 30743 3906 30777
rect 3854 30734 3906 30743
rect 4014 30777 4066 30786
rect 4014 30743 4023 30777
rect 4023 30743 4057 30777
rect 4057 30743 4066 30777
rect 4014 30734 4066 30743
rect 4174 30777 4226 30786
rect 4174 30743 4183 30777
rect 4183 30743 4217 30777
rect 4217 30743 4226 30777
rect 4174 30734 4226 30743
rect 4334 30777 4386 30786
rect 4334 30743 4343 30777
rect 4343 30743 4377 30777
rect 4377 30743 4386 30777
rect 4334 30734 4386 30743
rect 4494 30777 4546 30786
rect 4494 30743 4503 30777
rect 4503 30743 4537 30777
rect 4537 30743 4546 30777
rect 4494 30734 4546 30743
rect 4654 30777 4706 30786
rect 4654 30743 4663 30777
rect 4663 30743 4697 30777
rect 4697 30743 4706 30777
rect 4654 30734 4706 30743
rect 4814 30777 4866 30786
rect 4814 30743 4823 30777
rect 4823 30743 4857 30777
rect 4857 30743 4866 30777
rect 4814 30734 4866 30743
rect 4974 30777 5026 30786
rect 4974 30743 4983 30777
rect 4983 30743 5017 30777
rect 5017 30743 5026 30777
rect 4974 30734 5026 30743
rect 5134 30777 5186 30786
rect 5134 30743 5143 30777
rect 5143 30743 5177 30777
rect 5177 30743 5186 30777
rect 5134 30734 5186 30743
rect 5294 30777 5346 30786
rect 5294 30743 5303 30777
rect 5303 30743 5337 30777
rect 5337 30743 5346 30777
rect 5294 30734 5346 30743
rect 5454 30777 5506 30786
rect 5454 30743 5463 30777
rect 5463 30743 5497 30777
rect 5497 30743 5506 30777
rect 5454 30734 5506 30743
rect 5614 30777 5666 30786
rect 5614 30743 5623 30777
rect 5623 30743 5657 30777
rect 5657 30743 5666 30777
rect 5614 30734 5666 30743
rect 5774 30777 5826 30786
rect 5774 30743 5783 30777
rect 5783 30743 5817 30777
rect 5817 30743 5826 30777
rect 5774 30734 5826 30743
rect 5934 30777 5986 30786
rect 5934 30743 5943 30777
rect 5943 30743 5977 30777
rect 5977 30743 5986 30777
rect 5934 30734 5986 30743
rect 6094 30777 6146 30786
rect 6094 30743 6103 30777
rect 6103 30743 6137 30777
rect 6137 30743 6146 30777
rect 6094 30734 6146 30743
rect 6254 30777 6306 30786
rect 6254 30743 6263 30777
rect 6263 30743 6297 30777
rect 6297 30743 6306 30777
rect 6254 30734 6306 30743
rect 6414 30777 6466 30786
rect 6414 30743 6423 30777
rect 6423 30743 6457 30777
rect 6457 30743 6466 30777
rect 6414 30734 6466 30743
rect 6574 30777 6626 30786
rect 6574 30743 6583 30777
rect 6583 30743 6617 30777
rect 6617 30743 6626 30777
rect 6574 30734 6626 30743
rect 6734 30777 6786 30786
rect 6734 30743 6743 30777
rect 6743 30743 6777 30777
rect 6777 30743 6786 30777
rect 6734 30734 6786 30743
rect 6894 30777 6946 30786
rect 6894 30743 6903 30777
rect 6903 30743 6937 30777
rect 6937 30743 6946 30777
rect 6894 30734 6946 30743
rect 7054 30777 7106 30786
rect 7054 30743 7063 30777
rect 7063 30743 7097 30777
rect 7097 30743 7106 30777
rect 7054 30734 7106 30743
rect 7214 30777 7266 30786
rect 7214 30743 7223 30777
rect 7223 30743 7257 30777
rect 7257 30743 7266 30777
rect 7214 30734 7266 30743
rect 7374 30777 7426 30786
rect 7374 30743 7383 30777
rect 7383 30743 7417 30777
rect 7417 30743 7426 30777
rect 7374 30734 7426 30743
rect 7534 30777 7586 30786
rect 7534 30743 7543 30777
rect 7543 30743 7577 30777
rect 7577 30743 7586 30777
rect 7534 30734 7586 30743
rect 7694 30777 7746 30786
rect 7694 30743 7703 30777
rect 7703 30743 7737 30777
rect 7737 30743 7746 30777
rect 7694 30734 7746 30743
rect 7854 30777 7906 30786
rect 7854 30743 7863 30777
rect 7863 30743 7897 30777
rect 7897 30743 7906 30777
rect 7854 30734 7906 30743
rect 8014 30777 8066 30786
rect 8014 30743 8023 30777
rect 8023 30743 8057 30777
rect 8057 30743 8066 30777
rect 8014 30734 8066 30743
rect 8174 30777 8226 30786
rect 8174 30743 8183 30777
rect 8183 30743 8217 30777
rect 8217 30743 8226 30777
rect 8174 30734 8226 30743
rect 8334 30777 8386 30786
rect 8334 30743 8343 30777
rect 8343 30743 8377 30777
rect 8377 30743 8386 30777
rect 8334 30734 8386 30743
rect 12494 30777 12546 30786
rect 12494 30743 12503 30777
rect 12503 30743 12537 30777
rect 12537 30743 12546 30777
rect 12494 30734 12546 30743
rect 12654 30777 12706 30786
rect 12654 30743 12663 30777
rect 12663 30743 12697 30777
rect 12697 30743 12706 30777
rect 12654 30734 12706 30743
rect 12814 30777 12866 30786
rect 12814 30743 12823 30777
rect 12823 30743 12857 30777
rect 12857 30743 12866 30777
rect 12814 30734 12866 30743
rect 12974 30777 13026 30786
rect 12974 30743 12983 30777
rect 12983 30743 13017 30777
rect 13017 30743 13026 30777
rect 12974 30734 13026 30743
rect 13134 30777 13186 30786
rect 13134 30743 13143 30777
rect 13143 30743 13177 30777
rect 13177 30743 13186 30777
rect 13134 30734 13186 30743
rect 13294 30777 13346 30786
rect 13294 30743 13303 30777
rect 13303 30743 13337 30777
rect 13337 30743 13346 30777
rect 13294 30734 13346 30743
rect 13454 30777 13506 30786
rect 13454 30743 13463 30777
rect 13463 30743 13497 30777
rect 13497 30743 13506 30777
rect 13454 30734 13506 30743
rect 13614 30777 13666 30786
rect 13614 30743 13623 30777
rect 13623 30743 13657 30777
rect 13657 30743 13666 30777
rect 13614 30734 13666 30743
rect 13774 30777 13826 30786
rect 13774 30743 13783 30777
rect 13783 30743 13817 30777
rect 13817 30743 13826 30777
rect 13774 30734 13826 30743
rect 13934 30777 13986 30786
rect 13934 30743 13943 30777
rect 13943 30743 13977 30777
rect 13977 30743 13986 30777
rect 13934 30734 13986 30743
rect 14094 30777 14146 30786
rect 14094 30743 14103 30777
rect 14103 30743 14137 30777
rect 14137 30743 14146 30777
rect 14094 30734 14146 30743
rect 14254 30777 14306 30786
rect 14254 30743 14263 30777
rect 14263 30743 14297 30777
rect 14297 30743 14306 30777
rect 14254 30734 14306 30743
rect 14414 30777 14466 30786
rect 14414 30743 14423 30777
rect 14423 30743 14457 30777
rect 14457 30743 14466 30777
rect 14414 30734 14466 30743
rect 14574 30777 14626 30786
rect 14574 30743 14583 30777
rect 14583 30743 14617 30777
rect 14617 30743 14626 30777
rect 14574 30734 14626 30743
rect 14734 30777 14786 30786
rect 14734 30743 14743 30777
rect 14743 30743 14777 30777
rect 14777 30743 14786 30777
rect 14734 30734 14786 30743
rect 14894 30777 14946 30786
rect 14894 30743 14903 30777
rect 14903 30743 14937 30777
rect 14937 30743 14946 30777
rect 14894 30734 14946 30743
rect 15054 30777 15106 30786
rect 15054 30743 15063 30777
rect 15063 30743 15097 30777
rect 15097 30743 15106 30777
rect 15054 30734 15106 30743
rect 15214 30777 15266 30786
rect 15214 30743 15223 30777
rect 15223 30743 15257 30777
rect 15257 30743 15266 30777
rect 15214 30734 15266 30743
rect 15374 30777 15426 30786
rect 15374 30743 15383 30777
rect 15383 30743 15417 30777
rect 15417 30743 15426 30777
rect 15374 30734 15426 30743
rect 15534 30777 15586 30786
rect 15534 30743 15543 30777
rect 15543 30743 15577 30777
rect 15577 30743 15586 30777
rect 15534 30734 15586 30743
rect 15694 30777 15746 30786
rect 15694 30743 15703 30777
rect 15703 30743 15737 30777
rect 15737 30743 15746 30777
rect 15694 30734 15746 30743
rect 15854 30777 15906 30786
rect 15854 30743 15863 30777
rect 15863 30743 15897 30777
rect 15897 30743 15906 30777
rect 15854 30734 15906 30743
rect 16014 30777 16066 30786
rect 16014 30743 16023 30777
rect 16023 30743 16057 30777
rect 16057 30743 16066 30777
rect 16014 30734 16066 30743
rect 16174 30777 16226 30786
rect 16174 30743 16183 30777
rect 16183 30743 16217 30777
rect 16217 30743 16226 30777
rect 16174 30734 16226 30743
rect 16334 30777 16386 30786
rect 16334 30743 16343 30777
rect 16343 30743 16377 30777
rect 16377 30743 16386 30777
rect 16334 30734 16386 30743
rect 16494 30777 16546 30786
rect 16494 30743 16503 30777
rect 16503 30743 16537 30777
rect 16537 30743 16546 30777
rect 16494 30734 16546 30743
rect 16654 30777 16706 30786
rect 16654 30743 16663 30777
rect 16663 30743 16697 30777
rect 16697 30743 16706 30777
rect 16654 30734 16706 30743
rect 16814 30777 16866 30786
rect 16814 30743 16823 30777
rect 16823 30743 16857 30777
rect 16857 30743 16866 30777
rect 16814 30734 16866 30743
rect 16974 30777 17026 30786
rect 16974 30743 16983 30777
rect 16983 30743 17017 30777
rect 17017 30743 17026 30777
rect 16974 30734 17026 30743
rect 17134 30777 17186 30786
rect 17134 30743 17143 30777
rect 17143 30743 17177 30777
rect 17177 30743 17186 30777
rect 17134 30734 17186 30743
rect 17294 30777 17346 30786
rect 17294 30743 17303 30777
rect 17303 30743 17337 30777
rect 17337 30743 17346 30777
rect 17294 30734 17346 30743
rect 17454 30777 17506 30786
rect 17454 30743 17463 30777
rect 17463 30743 17497 30777
rect 17497 30743 17506 30777
rect 17454 30734 17506 30743
rect 17614 30777 17666 30786
rect 17614 30743 17623 30777
rect 17623 30743 17657 30777
rect 17657 30743 17666 30777
rect 17614 30734 17666 30743
rect 17774 30777 17826 30786
rect 17774 30743 17783 30777
rect 17783 30743 17817 30777
rect 17817 30743 17826 30777
rect 17774 30734 17826 30743
rect 17934 30777 17986 30786
rect 17934 30743 17943 30777
rect 17943 30743 17977 30777
rect 17977 30743 17986 30777
rect 17934 30734 17986 30743
rect 18094 30777 18146 30786
rect 18094 30743 18103 30777
rect 18103 30743 18137 30777
rect 18137 30743 18146 30777
rect 18094 30734 18146 30743
rect 18254 30777 18306 30786
rect 18254 30743 18263 30777
rect 18263 30743 18297 30777
rect 18297 30743 18306 30777
rect 18254 30734 18306 30743
rect 18414 30777 18466 30786
rect 18414 30743 18423 30777
rect 18423 30743 18457 30777
rect 18457 30743 18466 30777
rect 18414 30734 18466 30743
rect 18574 30777 18626 30786
rect 18574 30743 18583 30777
rect 18583 30743 18617 30777
rect 18617 30743 18626 30777
rect 18574 30734 18626 30743
rect 18734 30777 18786 30786
rect 18734 30743 18743 30777
rect 18743 30743 18777 30777
rect 18777 30743 18786 30777
rect 18734 30734 18786 30743
rect 18894 30777 18946 30786
rect 18894 30743 18903 30777
rect 18903 30743 18937 30777
rect 18937 30743 18946 30777
rect 18894 30734 18946 30743
rect 23134 30777 23186 30786
rect 23134 30743 23143 30777
rect 23143 30743 23177 30777
rect 23177 30743 23186 30777
rect 23134 30734 23186 30743
rect 23294 30777 23346 30786
rect 23294 30743 23303 30777
rect 23303 30743 23337 30777
rect 23337 30743 23346 30777
rect 23294 30734 23346 30743
rect 23454 30777 23506 30786
rect 23454 30743 23463 30777
rect 23463 30743 23497 30777
rect 23497 30743 23506 30777
rect 23454 30734 23506 30743
rect 23614 30777 23666 30786
rect 23614 30743 23623 30777
rect 23623 30743 23657 30777
rect 23657 30743 23666 30777
rect 23614 30734 23666 30743
rect 23774 30777 23826 30786
rect 23774 30743 23783 30777
rect 23783 30743 23817 30777
rect 23817 30743 23826 30777
rect 23774 30734 23826 30743
rect 23934 30777 23986 30786
rect 23934 30743 23943 30777
rect 23943 30743 23977 30777
rect 23977 30743 23986 30777
rect 23934 30734 23986 30743
rect 24094 30777 24146 30786
rect 24094 30743 24103 30777
rect 24103 30743 24137 30777
rect 24137 30743 24146 30777
rect 24094 30734 24146 30743
rect 24254 30777 24306 30786
rect 24254 30743 24263 30777
rect 24263 30743 24297 30777
rect 24297 30743 24306 30777
rect 24254 30734 24306 30743
rect 24414 30777 24466 30786
rect 24414 30743 24423 30777
rect 24423 30743 24457 30777
rect 24457 30743 24466 30777
rect 24414 30734 24466 30743
rect 24574 30777 24626 30786
rect 24574 30743 24583 30777
rect 24583 30743 24617 30777
rect 24617 30743 24626 30777
rect 24574 30734 24626 30743
rect 24734 30777 24786 30786
rect 24734 30743 24743 30777
rect 24743 30743 24777 30777
rect 24777 30743 24786 30777
rect 24734 30734 24786 30743
rect 24894 30777 24946 30786
rect 24894 30743 24903 30777
rect 24903 30743 24937 30777
rect 24937 30743 24946 30777
rect 24894 30734 24946 30743
rect 25054 30777 25106 30786
rect 25054 30743 25063 30777
rect 25063 30743 25097 30777
rect 25097 30743 25106 30777
rect 25054 30734 25106 30743
rect 25214 30777 25266 30786
rect 25214 30743 25223 30777
rect 25223 30743 25257 30777
rect 25257 30743 25266 30777
rect 25214 30734 25266 30743
rect 25374 30777 25426 30786
rect 25374 30743 25383 30777
rect 25383 30743 25417 30777
rect 25417 30743 25426 30777
rect 25374 30734 25426 30743
rect 25534 30777 25586 30786
rect 25534 30743 25543 30777
rect 25543 30743 25577 30777
rect 25577 30743 25586 30777
rect 25534 30734 25586 30743
rect 25694 30777 25746 30786
rect 25694 30743 25703 30777
rect 25703 30743 25737 30777
rect 25737 30743 25746 30777
rect 25694 30734 25746 30743
rect 25854 30777 25906 30786
rect 25854 30743 25863 30777
rect 25863 30743 25897 30777
rect 25897 30743 25906 30777
rect 25854 30734 25906 30743
rect 26014 30777 26066 30786
rect 26014 30743 26023 30777
rect 26023 30743 26057 30777
rect 26057 30743 26066 30777
rect 26014 30734 26066 30743
rect 26174 30777 26226 30786
rect 26174 30743 26183 30777
rect 26183 30743 26217 30777
rect 26217 30743 26226 30777
rect 26174 30734 26226 30743
rect 26334 30777 26386 30786
rect 26334 30743 26343 30777
rect 26343 30743 26377 30777
rect 26377 30743 26386 30777
rect 26334 30734 26386 30743
rect 26494 30777 26546 30786
rect 26494 30743 26503 30777
rect 26503 30743 26537 30777
rect 26537 30743 26546 30777
rect 26494 30734 26546 30743
rect 26654 30777 26706 30786
rect 26654 30743 26663 30777
rect 26663 30743 26697 30777
rect 26697 30743 26706 30777
rect 26654 30734 26706 30743
rect 26814 30777 26866 30786
rect 26814 30743 26823 30777
rect 26823 30743 26857 30777
rect 26857 30743 26866 30777
rect 26814 30734 26866 30743
rect 26974 30777 27026 30786
rect 26974 30743 26983 30777
rect 26983 30743 27017 30777
rect 27017 30743 27026 30777
rect 26974 30734 27026 30743
rect 27134 30777 27186 30786
rect 27134 30743 27143 30777
rect 27143 30743 27177 30777
rect 27177 30743 27186 30777
rect 27134 30734 27186 30743
rect 27294 30777 27346 30786
rect 27294 30743 27303 30777
rect 27303 30743 27337 30777
rect 27337 30743 27346 30777
rect 27294 30734 27346 30743
rect 27454 30777 27506 30786
rect 27454 30743 27463 30777
rect 27463 30743 27497 30777
rect 27497 30743 27506 30777
rect 27454 30734 27506 30743
rect 27614 30777 27666 30786
rect 27614 30743 27623 30777
rect 27623 30743 27657 30777
rect 27657 30743 27666 30777
rect 27614 30734 27666 30743
rect 27774 30777 27826 30786
rect 27774 30743 27783 30777
rect 27783 30743 27817 30777
rect 27817 30743 27826 30777
rect 27774 30734 27826 30743
rect 27934 30777 27986 30786
rect 27934 30743 27943 30777
rect 27943 30743 27977 30777
rect 27977 30743 27986 30777
rect 27934 30734 27986 30743
rect 28094 30777 28146 30786
rect 28094 30743 28103 30777
rect 28103 30743 28137 30777
rect 28137 30743 28146 30777
rect 28094 30734 28146 30743
rect 28254 30777 28306 30786
rect 28254 30743 28263 30777
rect 28263 30743 28297 30777
rect 28297 30743 28306 30777
rect 28254 30734 28306 30743
rect 28414 30777 28466 30786
rect 28414 30743 28423 30777
rect 28423 30743 28457 30777
rect 28457 30743 28466 30777
rect 28414 30734 28466 30743
rect 28574 30777 28626 30786
rect 28574 30743 28583 30777
rect 28583 30743 28617 30777
rect 28617 30743 28626 30777
rect 28574 30734 28626 30743
rect 28734 30777 28786 30786
rect 28734 30743 28743 30777
rect 28743 30743 28777 30777
rect 28777 30743 28786 30777
rect 28734 30734 28786 30743
rect 28894 30777 28946 30786
rect 28894 30743 28903 30777
rect 28903 30743 28937 30777
rect 28937 30743 28946 30777
rect 28894 30734 28946 30743
rect 29054 30777 29106 30786
rect 29054 30743 29063 30777
rect 29063 30743 29097 30777
rect 29097 30743 29106 30777
rect 29054 30734 29106 30743
rect 29214 30777 29266 30786
rect 29214 30743 29223 30777
rect 29223 30743 29257 30777
rect 29257 30743 29266 30777
rect 29214 30734 29266 30743
rect 29374 30777 29426 30786
rect 29374 30743 29383 30777
rect 29383 30743 29417 30777
rect 29417 30743 29426 30777
rect 29374 30734 29426 30743
rect 33534 30777 33586 30786
rect 33534 30743 33543 30777
rect 33543 30743 33577 30777
rect 33577 30743 33586 30777
rect 33534 30734 33586 30743
rect 33694 30777 33746 30786
rect 33694 30743 33703 30777
rect 33703 30743 33737 30777
rect 33737 30743 33746 30777
rect 33694 30734 33746 30743
rect 33854 30777 33906 30786
rect 33854 30743 33863 30777
rect 33863 30743 33897 30777
rect 33897 30743 33906 30777
rect 33854 30734 33906 30743
rect 34014 30777 34066 30786
rect 34014 30743 34023 30777
rect 34023 30743 34057 30777
rect 34057 30743 34066 30777
rect 34014 30734 34066 30743
rect 34174 30777 34226 30786
rect 34174 30743 34183 30777
rect 34183 30743 34217 30777
rect 34217 30743 34226 30777
rect 34174 30734 34226 30743
rect 34334 30777 34386 30786
rect 34334 30743 34343 30777
rect 34343 30743 34377 30777
rect 34377 30743 34386 30777
rect 34334 30734 34386 30743
rect 34494 30777 34546 30786
rect 34494 30743 34503 30777
rect 34503 30743 34537 30777
rect 34537 30743 34546 30777
rect 34494 30734 34546 30743
rect 34654 30777 34706 30786
rect 34654 30743 34663 30777
rect 34663 30743 34697 30777
rect 34697 30743 34706 30777
rect 34654 30734 34706 30743
rect 34814 30777 34866 30786
rect 34814 30743 34823 30777
rect 34823 30743 34857 30777
rect 34857 30743 34866 30777
rect 34814 30734 34866 30743
rect 34974 30777 35026 30786
rect 34974 30743 34983 30777
rect 34983 30743 35017 30777
rect 35017 30743 35026 30777
rect 34974 30734 35026 30743
rect 35134 30777 35186 30786
rect 35134 30743 35143 30777
rect 35143 30743 35177 30777
rect 35177 30743 35186 30777
rect 35134 30734 35186 30743
rect 35294 30777 35346 30786
rect 35294 30743 35303 30777
rect 35303 30743 35337 30777
rect 35337 30743 35346 30777
rect 35294 30734 35346 30743
rect 35454 30777 35506 30786
rect 35454 30743 35463 30777
rect 35463 30743 35497 30777
rect 35497 30743 35506 30777
rect 35454 30734 35506 30743
rect 35614 30777 35666 30786
rect 35614 30743 35623 30777
rect 35623 30743 35657 30777
rect 35657 30743 35666 30777
rect 35614 30734 35666 30743
rect 35774 30777 35826 30786
rect 35774 30743 35783 30777
rect 35783 30743 35817 30777
rect 35817 30743 35826 30777
rect 35774 30734 35826 30743
rect 35934 30777 35986 30786
rect 35934 30743 35943 30777
rect 35943 30743 35977 30777
rect 35977 30743 35986 30777
rect 35934 30734 35986 30743
rect 36094 30777 36146 30786
rect 36094 30743 36103 30777
rect 36103 30743 36137 30777
rect 36137 30743 36146 30777
rect 36094 30734 36146 30743
rect 36254 30777 36306 30786
rect 36254 30743 36263 30777
rect 36263 30743 36297 30777
rect 36297 30743 36306 30777
rect 36254 30734 36306 30743
rect 36414 30777 36466 30786
rect 36414 30743 36423 30777
rect 36423 30743 36457 30777
rect 36457 30743 36466 30777
rect 36414 30734 36466 30743
rect 36574 30777 36626 30786
rect 36574 30743 36583 30777
rect 36583 30743 36617 30777
rect 36617 30743 36626 30777
rect 36574 30734 36626 30743
rect 36734 30777 36786 30786
rect 36734 30743 36743 30777
rect 36743 30743 36777 30777
rect 36777 30743 36786 30777
rect 36734 30734 36786 30743
rect 36894 30777 36946 30786
rect 36894 30743 36903 30777
rect 36903 30743 36937 30777
rect 36937 30743 36946 30777
rect 36894 30734 36946 30743
rect 37054 30777 37106 30786
rect 37054 30743 37063 30777
rect 37063 30743 37097 30777
rect 37097 30743 37106 30777
rect 37054 30734 37106 30743
rect 37214 30777 37266 30786
rect 37214 30743 37223 30777
rect 37223 30743 37257 30777
rect 37257 30743 37266 30777
rect 37214 30734 37266 30743
rect 37374 30777 37426 30786
rect 37374 30743 37383 30777
rect 37383 30743 37417 30777
rect 37417 30743 37426 30777
rect 37374 30734 37426 30743
rect 37534 30777 37586 30786
rect 37534 30743 37543 30777
rect 37543 30743 37577 30777
rect 37577 30743 37586 30777
rect 37534 30734 37586 30743
rect 37694 30777 37746 30786
rect 37694 30743 37703 30777
rect 37703 30743 37737 30777
rect 37737 30743 37746 30777
rect 37694 30734 37746 30743
rect 37854 30777 37906 30786
rect 37854 30743 37863 30777
rect 37863 30743 37897 30777
rect 37897 30743 37906 30777
rect 37854 30734 37906 30743
rect 38014 30777 38066 30786
rect 38014 30743 38023 30777
rect 38023 30743 38057 30777
rect 38057 30743 38066 30777
rect 38014 30734 38066 30743
rect 38174 30777 38226 30786
rect 38174 30743 38183 30777
rect 38183 30743 38217 30777
rect 38217 30743 38226 30777
rect 38174 30734 38226 30743
rect 38334 30777 38386 30786
rect 38334 30743 38343 30777
rect 38343 30743 38377 30777
rect 38377 30743 38386 30777
rect 38334 30734 38386 30743
rect 38494 30777 38546 30786
rect 38494 30743 38503 30777
rect 38503 30743 38537 30777
rect 38537 30743 38546 30777
rect 38494 30734 38546 30743
rect 38654 30777 38706 30786
rect 38654 30743 38663 30777
rect 38663 30743 38697 30777
rect 38697 30743 38706 30777
rect 38654 30734 38706 30743
rect 38814 30777 38866 30786
rect 38814 30743 38823 30777
rect 38823 30743 38857 30777
rect 38857 30743 38866 30777
rect 38814 30734 38866 30743
rect 38974 30777 39026 30786
rect 38974 30743 38983 30777
rect 38983 30743 39017 30777
rect 39017 30743 39026 30777
rect 38974 30734 39026 30743
rect 39134 30777 39186 30786
rect 39134 30743 39143 30777
rect 39143 30743 39177 30777
rect 39177 30743 39186 30777
rect 39134 30734 39186 30743
rect 39294 30777 39346 30786
rect 39294 30743 39303 30777
rect 39303 30743 39337 30777
rect 39337 30743 39346 30777
rect 39294 30734 39346 30743
rect 39454 30777 39506 30786
rect 39454 30743 39463 30777
rect 39463 30743 39497 30777
rect 39497 30743 39506 30777
rect 39454 30734 39506 30743
rect 39614 30777 39666 30786
rect 39614 30743 39623 30777
rect 39623 30743 39657 30777
rect 39657 30743 39666 30777
rect 39614 30734 39666 30743
rect 39774 30777 39826 30786
rect 39774 30743 39783 30777
rect 39783 30743 39817 30777
rect 39817 30743 39826 30777
rect 39774 30734 39826 30743
rect 39934 30777 39986 30786
rect 39934 30743 39943 30777
rect 39943 30743 39977 30777
rect 39977 30743 39986 30777
rect 39934 30734 39986 30743
rect 40094 30777 40146 30786
rect 40094 30743 40103 30777
rect 40103 30743 40137 30777
rect 40137 30743 40146 30777
rect 40094 30734 40146 30743
rect 40254 30777 40306 30786
rect 40254 30743 40263 30777
rect 40263 30743 40297 30777
rect 40297 30743 40306 30777
rect 40254 30734 40306 30743
rect 40414 30777 40466 30786
rect 40414 30743 40423 30777
rect 40423 30743 40457 30777
rect 40457 30743 40466 30777
rect 40414 30734 40466 30743
rect 40574 30777 40626 30786
rect 40574 30743 40583 30777
rect 40583 30743 40617 30777
rect 40617 30743 40626 30777
rect 40574 30734 40626 30743
rect 40734 30777 40786 30786
rect 40734 30743 40743 30777
rect 40743 30743 40777 30777
rect 40777 30743 40786 30777
rect 40734 30734 40786 30743
rect 40894 30777 40946 30786
rect 40894 30743 40903 30777
rect 40903 30743 40937 30777
rect 40937 30743 40946 30777
rect 40894 30734 40946 30743
rect 41054 30777 41106 30786
rect 41054 30743 41063 30777
rect 41063 30743 41097 30777
rect 41097 30743 41106 30777
rect 41054 30734 41106 30743
rect 41214 30777 41266 30786
rect 41214 30743 41223 30777
rect 41223 30743 41257 30777
rect 41257 30743 41266 30777
rect 41214 30734 41266 30743
rect 41374 30777 41426 30786
rect 41374 30743 41383 30777
rect 41383 30743 41417 30777
rect 41417 30743 41426 30777
rect 41374 30734 41426 30743
rect 41534 30777 41586 30786
rect 41534 30743 41543 30777
rect 41543 30743 41577 30777
rect 41577 30743 41586 30777
rect 41534 30734 41586 30743
rect 41694 30777 41746 30786
rect 41694 30743 41703 30777
rect 41703 30743 41737 30777
rect 41737 30743 41746 30777
rect 41694 30734 41746 30743
rect 41854 30777 41906 30786
rect 41854 30743 41863 30777
rect 41863 30743 41897 30777
rect 41897 30743 41906 30777
rect 41854 30734 41906 30743
rect 14 30457 66 30466
rect 14 30423 23 30457
rect 23 30423 57 30457
rect 57 30423 66 30457
rect 14 30414 66 30423
rect 174 30457 226 30466
rect 174 30423 183 30457
rect 183 30423 217 30457
rect 217 30423 226 30457
rect 174 30414 226 30423
rect 334 30457 386 30466
rect 334 30423 343 30457
rect 343 30423 377 30457
rect 377 30423 386 30457
rect 334 30414 386 30423
rect 494 30457 546 30466
rect 494 30423 503 30457
rect 503 30423 537 30457
rect 537 30423 546 30457
rect 494 30414 546 30423
rect 654 30457 706 30466
rect 654 30423 663 30457
rect 663 30423 697 30457
rect 697 30423 706 30457
rect 654 30414 706 30423
rect 814 30457 866 30466
rect 814 30423 823 30457
rect 823 30423 857 30457
rect 857 30423 866 30457
rect 814 30414 866 30423
rect 974 30457 1026 30466
rect 974 30423 983 30457
rect 983 30423 1017 30457
rect 1017 30423 1026 30457
rect 974 30414 1026 30423
rect 1134 30457 1186 30466
rect 1134 30423 1143 30457
rect 1143 30423 1177 30457
rect 1177 30423 1186 30457
rect 1134 30414 1186 30423
rect 1294 30457 1346 30466
rect 1294 30423 1303 30457
rect 1303 30423 1337 30457
rect 1337 30423 1346 30457
rect 1294 30414 1346 30423
rect 1454 30457 1506 30466
rect 1454 30423 1463 30457
rect 1463 30423 1497 30457
rect 1497 30423 1506 30457
rect 1454 30414 1506 30423
rect 1614 30457 1666 30466
rect 1614 30423 1623 30457
rect 1623 30423 1657 30457
rect 1657 30423 1666 30457
rect 1614 30414 1666 30423
rect 1774 30457 1826 30466
rect 1774 30423 1783 30457
rect 1783 30423 1817 30457
rect 1817 30423 1826 30457
rect 1774 30414 1826 30423
rect 1934 30457 1986 30466
rect 1934 30423 1943 30457
rect 1943 30423 1977 30457
rect 1977 30423 1986 30457
rect 1934 30414 1986 30423
rect 2094 30457 2146 30466
rect 2094 30423 2103 30457
rect 2103 30423 2137 30457
rect 2137 30423 2146 30457
rect 2094 30414 2146 30423
rect 2254 30457 2306 30466
rect 2254 30423 2263 30457
rect 2263 30423 2297 30457
rect 2297 30423 2306 30457
rect 2254 30414 2306 30423
rect 2414 30457 2466 30466
rect 2414 30423 2423 30457
rect 2423 30423 2457 30457
rect 2457 30423 2466 30457
rect 2414 30414 2466 30423
rect 2574 30457 2626 30466
rect 2574 30423 2583 30457
rect 2583 30423 2617 30457
rect 2617 30423 2626 30457
rect 2574 30414 2626 30423
rect 2734 30457 2786 30466
rect 2734 30423 2743 30457
rect 2743 30423 2777 30457
rect 2777 30423 2786 30457
rect 2734 30414 2786 30423
rect 2894 30457 2946 30466
rect 2894 30423 2903 30457
rect 2903 30423 2937 30457
rect 2937 30423 2946 30457
rect 2894 30414 2946 30423
rect 3054 30457 3106 30466
rect 3054 30423 3063 30457
rect 3063 30423 3097 30457
rect 3097 30423 3106 30457
rect 3054 30414 3106 30423
rect 3214 30457 3266 30466
rect 3214 30423 3223 30457
rect 3223 30423 3257 30457
rect 3257 30423 3266 30457
rect 3214 30414 3266 30423
rect 3374 30457 3426 30466
rect 3374 30423 3383 30457
rect 3383 30423 3417 30457
rect 3417 30423 3426 30457
rect 3374 30414 3426 30423
rect 3534 30457 3586 30466
rect 3534 30423 3543 30457
rect 3543 30423 3577 30457
rect 3577 30423 3586 30457
rect 3534 30414 3586 30423
rect 3694 30457 3746 30466
rect 3694 30423 3703 30457
rect 3703 30423 3737 30457
rect 3737 30423 3746 30457
rect 3694 30414 3746 30423
rect 3854 30457 3906 30466
rect 3854 30423 3863 30457
rect 3863 30423 3897 30457
rect 3897 30423 3906 30457
rect 3854 30414 3906 30423
rect 4014 30457 4066 30466
rect 4014 30423 4023 30457
rect 4023 30423 4057 30457
rect 4057 30423 4066 30457
rect 4014 30414 4066 30423
rect 4174 30457 4226 30466
rect 4174 30423 4183 30457
rect 4183 30423 4217 30457
rect 4217 30423 4226 30457
rect 4174 30414 4226 30423
rect 4334 30457 4386 30466
rect 4334 30423 4343 30457
rect 4343 30423 4377 30457
rect 4377 30423 4386 30457
rect 4334 30414 4386 30423
rect 4494 30457 4546 30466
rect 4494 30423 4503 30457
rect 4503 30423 4537 30457
rect 4537 30423 4546 30457
rect 4494 30414 4546 30423
rect 4654 30457 4706 30466
rect 4654 30423 4663 30457
rect 4663 30423 4697 30457
rect 4697 30423 4706 30457
rect 4654 30414 4706 30423
rect 4814 30457 4866 30466
rect 4814 30423 4823 30457
rect 4823 30423 4857 30457
rect 4857 30423 4866 30457
rect 4814 30414 4866 30423
rect 4974 30457 5026 30466
rect 4974 30423 4983 30457
rect 4983 30423 5017 30457
rect 5017 30423 5026 30457
rect 4974 30414 5026 30423
rect 5134 30457 5186 30466
rect 5134 30423 5143 30457
rect 5143 30423 5177 30457
rect 5177 30423 5186 30457
rect 5134 30414 5186 30423
rect 5294 30457 5346 30466
rect 5294 30423 5303 30457
rect 5303 30423 5337 30457
rect 5337 30423 5346 30457
rect 5294 30414 5346 30423
rect 5454 30457 5506 30466
rect 5454 30423 5463 30457
rect 5463 30423 5497 30457
rect 5497 30423 5506 30457
rect 5454 30414 5506 30423
rect 5614 30457 5666 30466
rect 5614 30423 5623 30457
rect 5623 30423 5657 30457
rect 5657 30423 5666 30457
rect 5614 30414 5666 30423
rect 5774 30457 5826 30466
rect 5774 30423 5783 30457
rect 5783 30423 5817 30457
rect 5817 30423 5826 30457
rect 5774 30414 5826 30423
rect 5934 30457 5986 30466
rect 5934 30423 5943 30457
rect 5943 30423 5977 30457
rect 5977 30423 5986 30457
rect 5934 30414 5986 30423
rect 6094 30457 6146 30466
rect 6094 30423 6103 30457
rect 6103 30423 6137 30457
rect 6137 30423 6146 30457
rect 6094 30414 6146 30423
rect 6254 30457 6306 30466
rect 6254 30423 6263 30457
rect 6263 30423 6297 30457
rect 6297 30423 6306 30457
rect 6254 30414 6306 30423
rect 6414 30457 6466 30466
rect 6414 30423 6423 30457
rect 6423 30423 6457 30457
rect 6457 30423 6466 30457
rect 6414 30414 6466 30423
rect 6574 30457 6626 30466
rect 6574 30423 6583 30457
rect 6583 30423 6617 30457
rect 6617 30423 6626 30457
rect 6574 30414 6626 30423
rect 6734 30457 6786 30466
rect 6734 30423 6743 30457
rect 6743 30423 6777 30457
rect 6777 30423 6786 30457
rect 6734 30414 6786 30423
rect 6894 30457 6946 30466
rect 6894 30423 6903 30457
rect 6903 30423 6937 30457
rect 6937 30423 6946 30457
rect 6894 30414 6946 30423
rect 7054 30457 7106 30466
rect 7054 30423 7063 30457
rect 7063 30423 7097 30457
rect 7097 30423 7106 30457
rect 7054 30414 7106 30423
rect 7214 30457 7266 30466
rect 7214 30423 7223 30457
rect 7223 30423 7257 30457
rect 7257 30423 7266 30457
rect 7214 30414 7266 30423
rect 7374 30457 7426 30466
rect 7374 30423 7383 30457
rect 7383 30423 7417 30457
rect 7417 30423 7426 30457
rect 7374 30414 7426 30423
rect 7534 30457 7586 30466
rect 7534 30423 7543 30457
rect 7543 30423 7577 30457
rect 7577 30423 7586 30457
rect 7534 30414 7586 30423
rect 7694 30457 7746 30466
rect 7694 30423 7703 30457
rect 7703 30423 7737 30457
rect 7737 30423 7746 30457
rect 7694 30414 7746 30423
rect 7854 30457 7906 30466
rect 7854 30423 7863 30457
rect 7863 30423 7897 30457
rect 7897 30423 7906 30457
rect 7854 30414 7906 30423
rect 8014 30457 8066 30466
rect 8014 30423 8023 30457
rect 8023 30423 8057 30457
rect 8057 30423 8066 30457
rect 8014 30414 8066 30423
rect 8174 30457 8226 30466
rect 8174 30423 8183 30457
rect 8183 30423 8217 30457
rect 8217 30423 8226 30457
rect 8174 30414 8226 30423
rect 8334 30457 8386 30466
rect 8334 30423 8343 30457
rect 8343 30423 8377 30457
rect 8377 30423 8386 30457
rect 8334 30414 8386 30423
rect 12494 30457 12546 30466
rect 12494 30423 12503 30457
rect 12503 30423 12537 30457
rect 12537 30423 12546 30457
rect 12494 30414 12546 30423
rect 12654 30457 12706 30466
rect 12654 30423 12663 30457
rect 12663 30423 12697 30457
rect 12697 30423 12706 30457
rect 12654 30414 12706 30423
rect 12814 30457 12866 30466
rect 12814 30423 12823 30457
rect 12823 30423 12857 30457
rect 12857 30423 12866 30457
rect 12814 30414 12866 30423
rect 12974 30457 13026 30466
rect 12974 30423 12983 30457
rect 12983 30423 13017 30457
rect 13017 30423 13026 30457
rect 12974 30414 13026 30423
rect 13134 30457 13186 30466
rect 13134 30423 13143 30457
rect 13143 30423 13177 30457
rect 13177 30423 13186 30457
rect 13134 30414 13186 30423
rect 13294 30457 13346 30466
rect 13294 30423 13303 30457
rect 13303 30423 13337 30457
rect 13337 30423 13346 30457
rect 13294 30414 13346 30423
rect 13454 30457 13506 30466
rect 13454 30423 13463 30457
rect 13463 30423 13497 30457
rect 13497 30423 13506 30457
rect 13454 30414 13506 30423
rect 13614 30457 13666 30466
rect 13614 30423 13623 30457
rect 13623 30423 13657 30457
rect 13657 30423 13666 30457
rect 13614 30414 13666 30423
rect 13774 30457 13826 30466
rect 13774 30423 13783 30457
rect 13783 30423 13817 30457
rect 13817 30423 13826 30457
rect 13774 30414 13826 30423
rect 13934 30457 13986 30466
rect 13934 30423 13943 30457
rect 13943 30423 13977 30457
rect 13977 30423 13986 30457
rect 13934 30414 13986 30423
rect 14094 30457 14146 30466
rect 14094 30423 14103 30457
rect 14103 30423 14137 30457
rect 14137 30423 14146 30457
rect 14094 30414 14146 30423
rect 14254 30457 14306 30466
rect 14254 30423 14263 30457
rect 14263 30423 14297 30457
rect 14297 30423 14306 30457
rect 14254 30414 14306 30423
rect 14414 30457 14466 30466
rect 14414 30423 14423 30457
rect 14423 30423 14457 30457
rect 14457 30423 14466 30457
rect 14414 30414 14466 30423
rect 14574 30457 14626 30466
rect 14574 30423 14583 30457
rect 14583 30423 14617 30457
rect 14617 30423 14626 30457
rect 14574 30414 14626 30423
rect 14734 30457 14786 30466
rect 14734 30423 14743 30457
rect 14743 30423 14777 30457
rect 14777 30423 14786 30457
rect 14734 30414 14786 30423
rect 14894 30457 14946 30466
rect 14894 30423 14903 30457
rect 14903 30423 14937 30457
rect 14937 30423 14946 30457
rect 14894 30414 14946 30423
rect 15054 30457 15106 30466
rect 15054 30423 15063 30457
rect 15063 30423 15097 30457
rect 15097 30423 15106 30457
rect 15054 30414 15106 30423
rect 15214 30457 15266 30466
rect 15214 30423 15223 30457
rect 15223 30423 15257 30457
rect 15257 30423 15266 30457
rect 15214 30414 15266 30423
rect 15374 30457 15426 30466
rect 15374 30423 15383 30457
rect 15383 30423 15417 30457
rect 15417 30423 15426 30457
rect 15374 30414 15426 30423
rect 15534 30457 15586 30466
rect 15534 30423 15543 30457
rect 15543 30423 15577 30457
rect 15577 30423 15586 30457
rect 15534 30414 15586 30423
rect 15694 30457 15746 30466
rect 15694 30423 15703 30457
rect 15703 30423 15737 30457
rect 15737 30423 15746 30457
rect 15694 30414 15746 30423
rect 15854 30457 15906 30466
rect 15854 30423 15863 30457
rect 15863 30423 15897 30457
rect 15897 30423 15906 30457
rect 15854 30414 15906 30423
rect 16014 30457 16066 30466
rect 16014 30423 16023 30457
rect 16023 30423 16057 30457
rect 16057 30423 16066 30457
rect 16014 30414 16066 30423
rect 16174 30457 16226 30466
rect 16174 30423 16183 30457
rect 16183 30423 16217 30457
rect 16217 30423 16226 30457
rect 16174 30414 16226 30423
rect 16334 30457 16386 30466
rect 16334 30423 16343 30457
rect 16343 30423 16377 30457
rect 16377 30423 16386 30457
rect 16334 30414 16386 30423
rect 16494 30457 16546 30466
rect 16494 30423 16503 30457
rect 16503 30423 16537 30457
rect 16537 30423 16546 30457
rect 16494 30414 16546 30423
rect 16654 30457 16706 30466
rect 16654 30423 16663 30457
rect 16663 30423 16697 30457
rect 16697 30423 16706 30457
rect 16654 30414 16706 30423
rect 16814 30457 16866 30466
rect 16814 30423 16823 30457
rect 16823 30423 16857 30457
rect 16857 30423 16866 30457
rect 16814 30414 16866 30423
rect 16974 30457 17026 30466
rect 16974 30423 16983 30457
rect 16983 30423 17017 30457
rect 17017 30423 17026 30457
rect 16974 30414 17026 30423
rect 17134 30457 17186 30466
rect 17134 30423 17143 30457
rect 17143 30423 17177 30457
rect 17177 30423 17186 30457
rect 17134 30414 17186 30423
rect 17294 30457 17346 30466
rect 17294 30423 17303 30457
rect 17303 30423 17337 30457
rect 17337 30423 17346 30457
rect 17294 30414 17346 30423
rect 17454 30457 17506 30466
rect 17454 30423 17463 30457
rect 17463 30423 17497 30457
rect 17497 30423 17506 30457
rect 17454 30414 17506 30423
rect 17614 30457 17666 30466
rect 17614 30423 17623 30457
rect 17623 30423 17657 30457
rect 17657 30423 17666 30457
rect 17614 30414 17666 30423
rect 17774 30457 17826 30466
rect 17774 30423 17783 30457
rect 17783 30423 17817 30457
rect 17817 30423 17826 30457
rect 17774 30414 17826 30423
rect 17934 30457 17986 30466
rect 17934 30423 17943 30457
rect 17943 30423 17977 30457
rect 17977 30423 17986 30457
rect 17934 30414 17986 30423
rect 18094 30457 18146 30466
rect 18094 30423 18103 30457
rect 18103 30423 18137 30457
rect 18137 30423 18146 30457
rect 18094 30414 18146 30423
rect 18254 30457 18306 30466
rect 18254 30423 18263 30457
rect 18263 30423 18297 30457
rect 18297 30423 18306 30457
rect 18254 30414 18306 30423
rect 18414 30457 18466 30466
rect 18414 30423 18423 30457
rect 18423 30423 18457 30457
rect 18457 30423 18466 30457
rect 18414 30414 18466 30423
rect 18574 30457 18626 30466
rect 18574 30423 18583 30457
rect 18583 30423 18617 30457
rect 18617 30423 18626 30457
rect 18574 30414 18626 30423
rect 18734 30457 18786 30466
rect 18734 30423 18743 30457
rect 18743 30423 18777 30457
rect 18777 30423 18786 30457
rect 18734 30414 18786 30423
rect 18894 30457 18946 30466
rect 18894 30423 18903 30457
rect 18903 30423 18937 30457
rect 18937 30423 18946 30457
rect 18894 30414 18946 30423
rect 23134 30457 23186 30466
rect 23134 30423 23143 30457
rect 23143 30423 23177 30457
rect 23177 30423 23186 30457
rect 23134 30414 23186 30423
rect 23294 30457 23346 30466
rect 23294 30423 23303 30457
rect 23303 30423 23337 30457
rect 23337 30423 23346 30457
rect 23294 30414 23346 30423
rect 23454 30457 23506 30466
rect 23454 30423 23463 30457
rect 23463 30423 23497 30457
rect 23497 30423 23506 30457
rect 23454 30414 23506 30423
rect 23614 30457 23666 30466
rect 23614 30423 23623 30457
rect 23623 30423 23657 30457
rect 23657 30423 23666 30457
rect 23614 30414 23666 30423
rect 23774 30457 23826 30466
rect 23774 30423 23783 30457
rect 23783 30423 23817 30457
rect 23817 30423 23826 30457
rect 23774 30414 23826 30423
rect 23934 30457 23986 30466
rect 23934 30423 23943 30457
rect 23943 30423 23977 30457
rect 23977 30423 23986 30457
rect 23934 30414 23986 30423
rect 24094 30457 24146 30466
rect 24094 30423 24103 30457
rect 24103 30423 24137 30457
rect 24137 30423 24146 30457
rect 24094 30414 24146 30423
rect 24254 30457 24306 30466
rect 24254 30423 24263 30457
rect 24263 30423 24297 30457
rect 24297 30423 24306 30457
rect 24254 30414 24306 30423
rect 24414 30457 24466 30466
rect 24414 30423 24423 30457
rect 24423 30423 24457 30457
rect 24457 30423 24466 30457
rect 24414 30414 24466 30423
rect 24574 30457 24626 30466
rect 24574 30423 24583 30457
rect 24583 30423 24617 30457
rect 24617 30423 24626 30457
rect 24574 30414 24626 30423
rect 24734 30457 24786 30466
rect 24734 30423 24743 30457
rect 24743 30423 24777 30457
rect 24777 30423 24786 30457
rect 24734 30414 24786 30423
rect 24894 30457 24946 30466
rect 24894 30423 24903 30457
rect 24903 30423 24937 30457
rect 24937 30423 24946 30457
rect 24894 30414 24946 30423
rect 25054 30457 25106 30466
rect 25054 30423 25063 30457
rect 25063 30423 25097 30457
rect 25097 30423 25106 30457
rect 25054 30414 25106 30423
rect 25214 30457 25266 30466
rect 25214 30423 25223 30457
rect 25223 30423 25257 30457
rect 25257 30423 25266 30457
rect 25214 30414 25266 30423
rect 25374 30457 25426 30466
rect 25374 30423 25383 30457
rect 25383 30423 25417 30457
rect 25417 30423 25426 30457
rect 25374 30414 25426 30423
rect 25534 30457 25586 30466
rect 25534 30423 25543 30457
rect 25543 30423 25577 30457
rect 25577 30423 25586 30457
rect 25534 30414 25586 30423
rect 25694 30457 25746 30466
rect 25694 30423 25703 30457
rect 25703 30423 25737 30457
rect 25737 30423 25746 30457
rect 25694 30414 25746 30423
rect 25854 30457 25906 30466
rect 25854 30423 25863 30457
rect 25863 30423 25897 30457
rect 25897 30423 25906 30457
rect 25854 30414 25906 30423
rect 26014 30457 26066 30466
rect 26014 30423 26023 30457
rect 26023 30423 26057 30457
rect 26057 30423 26066 30457
rect 26014 30414 26066 30423
rect 26174 30457 26226 30466
rect 26174 30423 26183 30457
rect 26183 30423 26217 30457
rect 26217 30423 26226 30457
rect 26174 30414 26226 30423
rect 26334 30457 26386 30466
rect 26334 30423 26343 30457
rect 26343 30423 26377 30457
rect 26377 30423 26386 30457
rect 26334 30414 26386 30423
rect 26494 30457 26546 30466
rect 26494 30423 26503 30457
rect 26503 30423 26537 30457
rect 26537 30423 26546 30457
rect 26494 30414 26546 30423
rect 26654 30457 26706 30466
rect 26654 30423 26663 30457
rect 26663 30423 26697 30457
rect 26697 30423 26706 30457
rect 26654 30414 26706 30423
rect 26814 30457 26866 30466
rect 26814 30423 26823 30457
rect 26823 30423 26857 30457
rect 26857 30423 26866 30457
rect 26814 30414 26866 30423
rect 26974 30457 27026 30466
rect 26974 30423 26983 30457
rect 26983 30423 27017 30457
rect 27017 30423 27026 30457
rect 26974 30414 27026 30423
rect 27134 30457 27186 30466
rect 27134 30423 27143 30457
rect 27143 30423 27177 30457
rect 27177 30423 27186 30457
rect 27134 30414 27186 30423
rect 27294 30457 27346 30466
rect 27294 30423 27303 30457
rect 27303 30423 27337 30457
rect 27337 30423 27346 30457
rect 27294 30414 27346 30423
rect 27454 30457 27506 30466
rect 27454 30423 27463 30457
rect 27463 30423 27497 30457
rect 27497 30423 27506 30457
rect 27454 30414 27506 30423
rect 27614 30457 27666 30466
rect 27614 30423 27623 30457
rect 27623 30423 27657 30457
rect 27657 30423 27666 30457
rect 27614 30414 27666 30423
rect 27774 30457 27826 30466
rect 27774 30423 27783 30457
rect 27783 30423 27817 30457
rect 27817 30423 27826 30457
rect 27774 30414 27826 30423
rect 27934 30457 27986 30466
rect 27934 30423 27943 30457
rect 27943 30423 27977 30457
rect 27977 30423 27986 30457
rect 27934 30414 27986 30423
rect 28094 30457 28146 30466
rect 28094 30423 28103 30457
rect 28103 30423 28137 30457
rect 28137 30423 28146 30457
rect 28094 30414 28146 30423
rect 28254 30457 28306 30466
rect 28254 30423 28263 30457
rect 28263 30423 28297 30457
rect 28297 30423 28306 30457
rect 28254 30414 28306 30423
rect 28414 30457 28466 30466
rect 28414 30423 28423 30457
rect 28423 30423 28457 30457
rect 28457 30423 28466 30457
rect 28414 30414 28466 30423
rect 28574 30457 28626 30466
rect 28574 30423 28583 30457
rect 28583 30423 28617 30457
rect 28617 30423 28626 30457
rect 28574 30414 28626 30423
rect 28734 30457 28786 30466
rect 28734 30423 28743 30457
rect 28743 30423 28777 30457
rect 28777 30423 28786 30457
rect 28734 30414 28786 30423
rect 28894 30457 28946 30466
rect 28894 30423 28903 30457
rect 28903 30423 28937 30457
rect 28937 30423 28946 30457
rect 28894 30414 28946 30423
rect 29054 30457 29106 30466
rect 29054 30423 29063 30457
rect 29063 30423 29097 30457
rect 29097 30423 29106 30457
rect 29054 30414 29106 30423
rect 29214 30457 29266 30466
rect 29214 30423 29223 30457
rect 29223 30423 29257 30457
rect 29257 30423 29266 30457
rect 29214 30414 29266 30423
rect 29374 30457 29426 30466
rect 29374 30423 29383 30457
rect 29383 30423 29417 30457
rect 29417 30423 29426 30457
rect 29374 30414 29426 30423
rect 33534 30457 33586 30466
rect 33534 30423 33543 30457
rect 33543 30423 33577 30457
rect 33577 30423 33586 30457
rect 33534 30414 33586 30423
rect 33694 30457 33746 30466
rect 33694 30423 33703 30457
rect 33703 30423 33737 30457
rect 33737 30423 33746 30457
rect 33694 30414 33746 30423
rect 33854 30457 33906 30466
rect 33854 30423 33863 30457
rect 33863 30423 33897 30457
rect 33897 30423 33906 30457
rect 33854 30414 33906 30423
rect 34014 30457 34066 30466
rect 34014 30423 34023 30457
rect 34023 30423 34057 30457
rect 34057 30423 34066 30457
rect 34014 30414 34066 30423
rect 34174 30457 34226 30466
rect 34174 30423 34183 30457
rect 34183 30423 34217 30457
rect 34217 30423 34226 30457
rect 34174 30414 34226 30423
rect 34334 30457 34386 30466
rect 34334 30423 34343 30457
rect 34343 30423 34377 30457
rect 34377 30423 34386 30457
rect 34334 30414 34386 30423
rect 34494 30457 34546 30466
rect 34494 30423 34503 30457
rect 34503 30423 34537 30457
rect 34537 30423 34546 30457
rect 34494 30414 34546 30423
rect 34654 30457 34706 30466
rect 34654 30423 34663 30457
rect 34663 30423 34697 30457
rect 34697 30423 34706 30457
rect 34654 30414 34706 30423
rect 34814 30457 34866 30466
rect 34814 30423 34823 30457
rect 34823 30423 34857 30457
rect 34857 30423 34866 30457
rect 34814 30414 34866 30423
rect 34974 30457 35026 30466
rect 34974 30423 34983 30457
rect 34983 30423 35017 30457
rect 35017 30423 35026 30457
rect 34974 30414 35026 30423
rect 35134 30457 35186 30466
rect 35134 30423 35143 30457
rect 35143 30423 35177 30457
rect 35177 30423 35186 30457
rect 35134 30414 35186 30423
rect 35294 30457 35346 30466
rect 35294 30423 35303 30457
rect 35303 30423 35337 30457
rect 35337 30423 35346 30457
rect 35294 30414 35346 30423
rect 35454 30457 35506 30466
rect 35454 30423 35463 30457
rect 35463 30423 35497 30457
rect 35497 30423 35506 30457
rect 35454 30414 35506 30423
rect 35614 30457 35666 30466
rect 35614 30423 35623 30457
rect 35623 30423 35657 30457
rect 35657 30423 35666 30457
rect 35614 30414 35666 30423
rect 35774 30457 35826 30466
rect 35774 30423 35783 30457
rect 35783 30423 35817 30457
rect 35817 30423 35826 30457
rect 35774 30414 35826 30423
rect 35934 30457 35986 30466
rect 35934 30423 35943 30457
rect 35943 30423 35977 30457
rect 35977 30423 35986 30457
rect 35934 30414 35986 30423
rect 36094 30457 36146 30466
rect 36094 30423 36103 30457
rect 36103 30423 36137 30457
rect 36137 30423 36146 30457
rect 36094 30414 36146 30423
rect 36254 30457 36306 30466
rect 36254 30423 36263 30457
rect 36263 30423 36297 30457
rect 36297 30423 36306 30457
rect 36254 30414 36306 30423
rect 36414 30457 36466 30466
rect 36414 30423 36423 30457
rect 36423 30423 36457 30457
rect 36457 30423 36466 30457
rect 36414 30414 36466 30423
rect 36574 30457 36626 30466
rect 36574 30423 36583 30457
rect 36583 30423 36617 30457
rect 36617 30423 36626 30457
rect 36574 30414 36626 30423
rect 36734 30457 36786 30466
rect 36734 30423 36743 30457
rect 36743 30423 36777 30457
rect 36777 30423 36786 30457
rect 36734 30414 36786 30423
rect 36894 30457 36946 30466
rect 36894 30423 36903 30457
rect 36903 30423 36937 30457
rect 36937 30423 36946 30457
rect 36894 30414 36946 30423
rect 37054 30457 37106 30466
rect 37054 30423 37063 30457
rect 37063 30423 37097 30457
rect 37097 30423 37106 30457
rect 37054 30414 37106 30423
rect 37214 30457 37266 30466
rect 37214 30423 37223 30457
rect 37223 30423 37257 30457
rect 37257 30423 37266 30457
rect 37214 30414 37266 30423
rect 37374 30457 37426 30466
rect 37374 30423 37383 30457
rect 37383 30423 37417 30457
rect 37417 30423 37426 30457
rect 37374 30414 37426 30423
rect 37534 30457 37586 30466
rect 37534 30423 37543 30457
rect 37543 30423 37577 30457
rect 37577 30423 37586 30457
rect 37534 30414 37586 30423
rect 37694 30457 37746 30466
rect 37694 30423 37703 30457
rect 37703 30423 37737 30457
rect 37737 30423 37746 30457
rect 37694 30414 37746 30423
rect 37854 30457 37906 30466
rect 37854 30423 37863 30457
rect 37863 30423 37897 30457
rect 37897 30423 37906 30457
rect 37854 30414 37906 30423
rect 38014 30457 38066 30466
rect 38014 30423 38023 30457
rect 38023 30423 38057 30457
rect 38057 30423 38066 30457
rect 38014 30414 38066 30423
rect 38174 30457 38226 30466
rect 38174 30423 38183 30457
rect 38183 30423 38217 30457
rect 38217 30423 38226 30457
rect 38174 30414 38226 30423
rect 38334 30457 38386 30466
rect 38334 30423 38343 30457
rect 38343 30423 38377 30457
rect 38377 30423 38386 30457
rect 38334 30414 38386 30423
rect 38494 30457 38546 30466
rect 38494 30423 38503 30457
rect 38503 30423 38537 30457
rect 38537 30423 38546 30457
rect 38494 30414 38546 30423
rect 38654 30457 38706 30466
rect 38654 30423 38663 30457
rect 38663 30423 38697 30457
rect 38697 30423 38706 30457
rect 38654 30414 38706 30423
rect 38814 30457 38866 30466
rect 38814 30423 38823 30457
rect 38823 30423 38857 30457
rect 38857 30423 38866 30457
rect 38814 30414 38866 30423
rect 38974 30457 39026 30466
rect 38974 30423 38983 30457
rect 38983 30423 39017 30457
rect 39017 30423 39026 30457
rect 38974 30414 39026 30423
rect 39134 30457 39186 30466
rect 39134 30423 39143 30457
rect 39143 30423 39177 30457
rect 39177 30423 39186 30457
rect 39134 30414 39186 30423
rect 39294 30457 39346 30466
rect 39294 30423 39303 30457
rect 39303 30423 39337 30457
rect 39337 30423 39346 30457
rect 39294 30414 39346 30423
rect 39454 30457 39506 30466
rect 39454 30423 39463 30457
rect 39463 30423 39497 30457
rect 39497 30423 39506 30457
rect 39454 30414 39506 30423
rect 39614 30457 39666 30466
rect 39614 30423 39623 30457
rect 39623 30423 39657 30457
rect 39657 30423 39666 30457
rect 39614 30414 39666 30423
rect 39774 30457 39826 30466
rect 39774 30423 39783 30457
rect 39783 30423 39817 30457
rect 39817 30423 39826 30457
rect 39774 30414 39826 30423
rect 39934 30457 39986 30466
rect 39934 30423 39943 30457
rect 39943 30423 39977 30457
rect 39977 30423 39986 30457
rect 39934 30414 39986 30423
rect 40094 30457 40146 30466
rect 40094 30423 40103 30457
rect 40103 30423 40137 30457
rect 40137 30423 40146 30457
rect 40094 30414 40146 30423
rect 40254 30457 40306 30466
rect 40254 30423 40263 30457
rect 40263 30423 40297 30457
rect 40297 30423 40306 30457
rect 40254 30414 40306 30423
rect 40414 30457 40466 30466
rect 40414 30423 40423 30457
rect 40423 30423 40457 30457
rect 40457 30423 40466 30457
rect 40414 30414 40466 30423
rect 40574 30457 40626 30466
rect 40574 30423 40583 30457
rect 40583 30423 40617 30457
rect 40617 30423 40626 30457
rect 40574 30414 40626 30423
rect 40734 30457 40786 30466
rect 40734 30423 40743 30457
rect 40743 30423 40777 30457
rect 40777 30423 40786 30457
rect 40734 30414 40786 30423
rect 40894 30457 40946 30466
rect 40894 30423 40903 30457
rect 40903 30423 40937 30457
rect 40937 30423 40946 30457
rect 40894 30414 40946 30423
rect 41054 30457 41106 30466
rect 41054 30423 41063 30457
rect 41063 30423 41097 30457
rect 41097 30423 41106 30457
rect 41054 30414 41106 30423
rect 41214 30457 41266 30466
rect 41214 30423 41223 30457
rect 41223 30423 41257 30457
rect 41257 30423 41266 30457
rect 41214 30414 41266 30423
rect 41374 30457 41426 30466
rect 41374 30423 41383 30457
rect 41383 30423 41417 30457
rect 41417 30423 41426 30457
rect 41374 30414 41426 30423
rect 41534 30457 41586 30466
rect 41534 30423 41543 30457
rect 41543 30423 41577 30457
rect 41577 30423 41586 30457
rect 41534 30414 41586 30423
rect 41694 30457 41746 30466
rect 41694 30423 41703 30457
rect 41703 30423 41737 30457
rect 41737 30423 41746 30457
rect 41694 30414 41746 30423
rect 41854 30457 41906 30466
rect 41854 30423 41863 30457
rect 41863 30423 41897 30457
rect 41897 30423 41906 30457
rect 41854 30414 41906 30423
rect 14 30297 66 30306
rect 14 30263 23 30297
rect 23 30263 57 30297
rect 57 30263 66 30297
rect 14 30254 66 30263
rect 174 30297 226 30306
rect 174 30263 183 30297
rect 183 30263 217 30297
rect 217 30263 226 30297
rect 174 30254 226 30263
rect 334 30297 386 30306
rect 334 30263 343 30297
rect 343 30263 377 30297
rect 377 30263 386 30297
rect 334 30254 386 30263
rect 494 30297 546 30306
rect 494 30263 503 30297
rect 503 30263 537 30297
rect 537 30263 546 30297
rect 494 30254 546 30263
rect 654 30297 706 30306
rect 654 30263 663 30297
rect 663 30263 697 30297
rect 697 30263 706 30297
rect 654 30254 706 30263
rect 814 30297 866 30306
rect 814 30263 823 30297
rect 823 30263 857 30297
rect 857 30263 866 30297
rect 814 30254 866 30263
rect 974 30297 1026 30306
rect 974 30263 983 30297
rect 983 30263 1017 30297
rect 1017 30263 1026 30297
rect 974 30254 1026 30263
rect 1134 30297 1186 30306
rect 1134 30263 1143 30297
rect 1143 30263 1177 30297
rect 1177 30263 1186 30297
rect 1134 30254 1186 30263
rect 1294 30297 1346 30306
rect 1294 30263 1303 30297
rect 1303 30263 1337 30297
rect 1337 30263 1346 30297
rect 1294 30254 1346 30263
rect 1454 30297 1506 30306
rect 1454 30263 1463 30297
rect 1463 30263 1497 30297
rect 1497 30263 1506 30297
rect 1454 30254 1506 30263
rect 1614 30297 1666 30306
rect 1614 30263 1623 30297
rect 1623 30263 1657 30297
rect 1657 30263 1666 30297
rect 1614 30254 1666 30263
rect 1774 30297 1826 30306
rect 1774 30263 1783 30297
rect 1783 30263 1817 30297
rect 1817 30263 1826 30297
rect 1774 30254 1826 30263
rect 1934 30297 1986 30306
rect 1934 30263 1943 30297
rect 1943 30263 1977 30297
rect 1977 30263 1986 30297
rect 1934 30254 1986 30263
rect 2094 30297 2146 30306
rect 2094 30263 2103 30297
rect 2103 30263 2137 30297
rect 2137 30263 2146 30297
rect 2094 30254 2146 30263
rect 2254 30297 2306 30306
rect 2254 30263 2263 30297
rect 2263 30263 2297 30297
rect 2297 30263 2306 30297
rect 2254 30254 2306 30263
rect 2414 30297 2466 30306
rect 2414 30263 2423 30297
rect 2423 30263 2457 30297
rect 2457 30263 2466 30297
rect 2414 30254 2466 30263
rect 2574 30297 2626 30306
rect 2574 30263 2583 30297
rect 2583 30263 2617 30297
rect 2617 30263 2626 30297
rect 2574 30254 2626 30263
rect 2734 30297 2786 30306
rect 2734 30263 2743 30297
rect 2743 30263 2777 30297
rect 2777 30263 2786 30297
rect 2734 30254 2786 30263
rect 2894 30297 2946 30306
rect 2894 30263 2903 30297
rect 2903 30263 2937 30297
rect 2937 30263 2946 30297
rect 2894 30254 2946 30263
rect 3054 30297 3106 30306
rect 3054 30263 3063 30297
rect 3063 30263 3097 30297
rect 3097 30263 3106 30297
rect 3054 30254 3106 30263
rect 3214 30297 3266 30306
rect 3214 30263 3223 30297
rect 3223 30263 3257 30297
rect 3257 30263 3266 30297
rect 3214 30254 3266 30263
rect 3374 30297 3426 30306
rect 3374 30263 3383 30297
rect 3383 30263 3417 30297
rect 3417 30263 3426 30297
rect 3374 30254 3426 30263
rect 3534 30297 3586 30306
rect 3534 30263 3543 30297
rect 3543 30263 3577 30297
rect 3577 30263 3586 30297
rect 3534 30254 3586 30263
rect 3694 30297 3746 30306
rect 3694 30263 3703 30297
rect 3703 30263 3737 30297
rect 3737 30263 3746 30297
rect 3694 30254 3746 30263
rect 3854 30297 3906 30306
rect 3854 30263 3863 30297
rect 3863 30263 3897 30297
rect 3897 30263 3906 30297
rect 3854 30254 3906 30263
rect 4014 30297 4066 30306
rect 4014 30263 4023 30297
rect 4023 30263 4057 30297
rect 4057 30263 4066 30297
rect 4014 30254 4066 30263
rect 4174 30297 4226 30306
rect 4174 30263 4183 30297
rect 4183 30263 4217 30297
rect 4217 30263 4226 30297
rect 4174 30254 4226 30263
rect 4334 30297 4386 30306
rect 4334 30263 4343 30297
rect 4343 30263 4377 30297
rect 4377 30263 4386 30297
rect 4334 30254 4386 30263
rect 4494 30297 4546 30306
rect 4494 30263 4503 30297
rect 4503 30263 4537 30297
rect 4537 30263 4546 30297
rect 4494 30254 4546 30263
rect 4654 30297 4706 30306
rect 4654 30263 4663 30297
rect 4663 30263 4697 30297
rect 4697 30263 4706 30297
rect 4654 30254 4706 30263
rect 4814 30297 4866 30306
rect 4814 30263 4823 30297
rect 4823 30263 4857 30297
rect 4857 30263 4866 30297
rect 4814 30254 4866 30263
rect 4974 30297 5026 30306
rect 4974 30263 4983 30297
rect 4983 30263 5017 30297
rect 5017 30263 5026 30297
rect 4974 30254 5026 30263
rect 5134 30297 5186 30306
rect 5134 30263 5143 30297
rect 5143 30263 5177 30297
rect 5177 30263 5186 30297
rect 5134 30254 5186 30263
rect 5294 30297 5346 30306
rect 5294 30263 5303 30297
rect 5303 30263 5337 30297
rect 5337 30263 5346 30297
rect 5294 30254 5346 30263
rect 5454 30297 5506 30306
rect 5454 30263 5463 30297
rect 5463 30263 5497 30297
rect 5497 30263 5506 30297
rect 5454 30254 5506 30263
rect 5614 30297 5666 30306
rect 5614 30263 5623 30297
rect 5623 30263 5657 30297
rect 5657 30263 5666 30297
rect 5614 30254 5666 30263
rect 5774 30297 5826 30306
rect 5774 30263 5783 30297
rect 5783 30263 5817 30297
rect 5817 30263 5826 30297
rect 5774 30254 5826 30263
rect 5934 30297 5986 30306
rect 5934 30263 5943 30297
rect 5943 30263 5977 30297
rect 5977 30263 5986 30297
rect 5934 30254 5986 30263
rect 6094 30297 6146 30306
rect 6094 30263 6103 30297
rect 6103 30263 6137 30297
rect 6137 30263 6146 30297
rect 6094 30254 6146 30263
rect 6254 30297 6306 30306
rect 6254 30263 6263 30297
rect 6263 30263 6297 30297
rect 6297 30263 6306 30297
rect 6254 30254 6306 30263
rect 6414 30297 6466 30306
rect 6414 30263 6423 30297
rect 6423 30263 6457 30297
rect 6457 30263 6466 30297
rect 6414 30254 6466 30263
rect 6574 30297 6626 30306
rect 6574 30263 6583 30297
rect 6583 30263 6617 30297
rect 6617 30263 6626 30297
rect 6574 30254 6626 30263
rect 6734 30297 6786 30306
rect 6734 30263 6743 30297
rect 6743 30263 6777 30297
rect 6777 30263 6786 30297
rect 6734 30254 6786 30263
rect 6894 30297 6946 30306
rect 6894 30263 6903 30297
rect 6903 30263 6937 30297
rect 6937 30263 6946 30297
rect 6894 30254 6946 30263
rect 7054 30297 7106 30306
rect 7054 30263 7063 30297
rect 7063 30263 7097 30297
rect 7097 30263 7106 30297
rect 7054 30254 7106 30263
rect 7214 30297 7266 30306
rect 7214 30263 7223 30297
rect 7223 30263 7257 30297
rect 7257 30263 7266 30297
rect 7214 30254 7266 30263
rect 7374 30297 7426 30306
rect 7374 30263 7383 30297
rect 7383 30263 7417 30297
rect 7417 30263 7426 30297
rect 7374 30254 7426 30263
rect 7534 30297 7586 30306
rect 7534 30263 7543 30297
rect 7543 30263 7577 30297
rect 7577 30263 7586 30297
rect 7534 30254 7586 30263
rect 7694 30297 7746 30306
rect 7694 30263 7703 30297
rect 7703 30263 7737 30297
rect 7737 30263 7746 30297
rect 7694 30254 7746 30263
rect 7854 30297 7906 30306
rect 7854 30263 7863 30297
rect 7863 30263 7897 30297
rect 7897 30263 7906 30297
rect 7854 30254 7906 30263
rect 8014 30297 8066 30306
rect 8014 30263 8023 30297
rect 8023 30263 8057 30297
rect 8057 30263 8066 30297
rect 8014 30254 8066 30263
rect 8174 30297 8226 30306
rect 8174 30263 8183 30297
rect 8183 30263 8217 30297
rect 8217 30263 8226 30297
rect 8174 30254 8226 30263
rect 8334 30297 8386 30306
rect 8334 30263 8343 30297
rect 8343 30263 8377 30297
rect 8377 30263 8386 30297
rect 8334 30254 8386 30263
rect 12494 30297 12546 30306
rect 12494 30263 12503 30297
rect 12503 30263 12537 30297
rect 12537 30263 12546 30297
rect 12494 30254 12546 30263
rect 12654 30297 12706 30306
rect 12654 30263 12663 30297
rect 12663 30263 12697 30297
rect 12697 30263 12706 30297
rect 12654 30254 12706 30263
rect 12814 30297 12866 30306
rect 12814 30263 12823 30297
rect 12823 30263 12857 30297
rect 12857 30263 12866 30297
rect 12814 30254 12866 30263
rect 12974 30297 13026 30306
rect 12974 30263 12983 30297
rect 12983 30263 13017 30297
rect 13017 30263 13026 30297
rect 12974 30254 13026 30263
rect 13134 30297 13186 30306
rect 13134 30263 13143 30297
rect 13143 30263 13177 30297
rect 13177 30263 13186 30297
rect 13134 30254 13186 30263
rect 13294 30297 13346 30306
rect 13294 30263 13303 30297
rect 13303 30263 13337 30297
rect 13337 30263 13346 30297
rect 13294 30254 13346 30263
rect 13454 30297 13506 30306
rect 13454 30263 13463 30297
rect 13463 30263 13497 30297
rect 13497 30263 13506 30297
rect 13454 30254 13506 30263
rect 13614 30297 13666 30306
rect 13614 30263 13623 30297
rect 13623 30263 13657 30297
rect 13657 30263 13666 30297
rect 13614 30254 13666 30263
rect 13774 30297 13826 30306
rect 13774 30263 13783 30297
rect 13783 30263 13817 30297
rect 13817 30263 13826 30297
rect 13774 30254 13826 30263
rect 13934 30297 13986 30306
rect 13934 30263 13943 30297
rect 13943 30263 13977 30297
rect 13977 30263 13986 30297
rect 13934 30254 13986 30263
rect 14094 30297 14146 30306
rect 14094 30263 14103 30297
rect 14103 30263 14137 30297
rect 14137 30263 14146 30297
rect 14094 30254 14146 30263
rect 14254 30297 14306 30306
rect 14254 30263 14263 30297
rect 14263 30263 14297 30297
rect 14297 30263 14306 30297
rect 14254 30254 14306 30263
rect 14414 30297 14466 30306
rect 14414 30263 14423 30297
rect 14423 30263 14457 30297
rect 14457 30263 14466 30297
rect 14414 30254 14466 30263
rect 14574 30297 14626 30306
rect 14574 30263 14583 30297
rect 14583 30263 14617 30297
rect 14617 30263 14626 30297
rect 14574 30254 14626 30263
rect 14734 30297 14786 30306
rect 14734 30263 14743 30297
rect 14743 30263 14777 30297
rect 14777 30263 14786 30297
rect 14734 30254 14786 30263
rect 14894 30297 14946 30306
rect 14894 30263 14903 30297
rect 14903 30263 14937 30297
rect 14937 30263 14946 30297
rect 14894 30254 14946 30263
rect 15054 30297 15106 30306
rect 15054 30263 15063 30297
rect 15063 30263 15097 30297
rect 15097 30263 15106 30297
rect 15054 30254 15106 30263
rect 15214 30297 15266 30306
rect 15214 30263 15223 30297
rect 15223 30263 15257 30297
rect 15257 30263 15266 30297
rect 15214 30254 15266 30263
rect 15374 30297 15426 30306
rect 15374 30263 15383 30297
rect 15383 30263 15417 30297
rect 15417 30263 15426 30297
rect 15374 30254 15426 30263
rect 15534 30297 15586 30306
rect 15534 30263 15543 30297
rect 15543 30263 15577 30297
rect 15577 30263 15586 30297
rect 15534 30254 15586 30263
rect 15694 30297 15746 30306
rect 15694 30263 15703 30297
rect 15703 30263 15737 30297
rect 15737 30263 15746 30297
rect 15694 30254 15746 30263
rect 15854 30297 15906 30306
rect 15854 30263 15863 30297
rect 15863 30263 15897 30297
rect 15897 30263 15906 30297
rect 15854 30254 15906 30263
rect 16014 30297 16066 30306
rect 16014 30263 16023 30297
rect 16023 30263 16057 30297
rect 16057 30263 16066 30297
rect 16014 30254 16066 30263
rect 16174 30297 16226 30306
rect 16174 30263 16183 30297
rect 16183 30263 16217 30297
rect 16217 30263 16226 30297
rect 16174 30254 16226 30263
rect 16334 30297 16386 30306
rect 16334 30263 16343 30297
rect 16343 30263 16377 30297
rect 16377 30263 16386 30297
rect 16334 30254 16386 30263
rect 16494 30297 16546 30306
rect 16494 30263 16503 30297
rect 16503 30263 16537 30297
rect 16537 30263 16546 30297
rect 16494 30254 16546 30263
rect 16654 30297 16706 30306
rect 16654 30263 16663 30297
rect 16663 30263 16697 30297
rect 16697 30263 16706 30297
rect 16654 30254 16706 30263
rect 16814 30297 16866 30306
rect 16814 30263 16823 30297
rect 16823 30263 16857 30297
rect 16857 30263 16866 30297
rect 16814 30254 16866 30263
rect 16974 30297 17026 30306
rect 16974 30263 16983 30297
rect 16983 30263 17017 30297
rect 17017 30263 17026 30297
rect 16974 30254 17026 30263
rect 17134 30297 17186 30306
rect 17134 30263 17143 30297
rect 17143 30263 17177 30297
rect 17177 30263 17186 30297
rect 17134 30254 17186 30263
rect 17294 30297 17346 30306
rect 17294 30263 17303 30297
rect 17303 30263 17337 30297
rect 17337 30263 17346 30297
rect 17294 30254 17346 30263
rect 17454 30297 17506 30306
rect 17454 30263 17463 30297
rect 17463 30263 17497 30297
rect 17497 30263 17506 30297
rect 17454 30254 17506 30263
rect 17614 30297 17666 30306
rect 17614 30263 17623 30297
rect 17623 30263 17657 30297
rect 17657 30263 17666 30297
rect 17614 30254 17666 30263
rect 17774 30297 17826 30306
rect 17774 30263 17783 30297
rect 17783 30263 17817 30297
rect 17817 30263 17826 30297
rect 17774 30254 17826 30263
rect 17934 30297 17986 30306
rect 17934 30263 17943 30297
rect 17943 30263 17977 30297
rect 17977 30263 17986 30297
rect 17934 30254 17986 30263
rect 18094 30297 18146 30306
rect 18094 30263 18103 30297
rect 18103 30263 18137 30297
rect 18137 30263 18146 30297
rect 18094 30254 18146 30263
rect 18254 30297 18306 30306
rect 18254 30263 18263 30297
rect 18263 30263 18297 30297
rect 18297 30263 18306 30297
rect 18254 30254 18306 30263
rect 18414 30297 18466 30306
rect 18414 30263 18423 30297
rect 18423 30263 18457 30297
rect 18457 30263 18466 30297
rect 18414 30254 18466 30263
rect 18574 30297 18626 30306
rect 18574 30263 18583 30297
rect 18583 30263 18617 30297
rect 18617 30263 18626 30297
rect 18574 30254 18626 30263
rect 18734 30297 18786 30306
rect 18734 30263 18743 30297
rect 18743 30263 18777 30297
rect 18777 30263 18786 30297
rect 18734 30254 18786 30263
rect 18894 30297 18946 30306
rect 18894 30263 18903 30297
rect 18903 30263 18937 30297
rect 18937 30263 18946 30297
rect 18894 30254 18946 30263
rect 23134 30297 23186 30306
rect 23134 30263 23143 30297
rect 23143 30263 23177 30297
rect 23177 30263 23186 30297
rect 23134 30254 23186 30263
rect 23294 30297 23346 30306
rect 23294 30263 23303 30297
rect 23303 30263 23337 30297
rect 23337 30263 23346 30297
rect 23294 30254 23346 30263
rect 23454 30297 23506 30306
rect 23454 30263 23463 30297
rect 23463 30263 23497 30297
rect 23497 30263 23506 30297
rect 23454 30254 23506 30263
rect 23614 30297 23666 30306
rect 23614 30263 23623 30297
rect 23623 30263 23657 30297
rect 23657 30263 23666 30297
rect 23614 30254 23666 30263
rect 23774 30297 23826 30306
rect 23774 30263 23783 30297
rect 23783 30263 23817 30297
rect 23817 30263 23826 30297
rect 23774 30254 23826 30263
rect 23934 30297 23986 30306
rect 23934 30263 23943 30297
rect 23943 30263 23977 30297
rect 23977 30263 23986 30297
rect 23934 30254 23986 30263
rect 24094 30297 24146 30306
rect 24094 30263 24103 30297
rect 24103 30263 24137 30297
rect 24137 30263 24146 30297
rect 24094 30254 24146 30263
rect 24254 30297 24306 30306
rect 24254 30263 24263 30297
rect 24263 30263 24297 30297
rect 24297 30263 24306 30297
rect 24254 30254 24306 30263
rect 24414 30297 24466 30306
rect 24414 30263 24423 30297
rect 24423 30263 24457 30297
rect 24457 30263 24466 30297
rect 24414 30254 24466 30263
rect 24574 30297 24626 30306
rect 24574 30263 24583 30297
rect 24583 30263 24617 30297
rect 24617 30263 24626 30297
rect 24574 30254 24626 30263
rect 24734 30297 24786 30306
rect 24734 30263 24743 30297
rect 24743 30263 24777 30297
rect 24777 30263 24786 30297
rect 24734 30254 24786 30263
rect 24894 30297 24946 30306
rect 24894 30263 24903 30297
rect 24903 30263 24937 30297
rect 24937 30263 24946 30297
rect 24894 30254 24946 30263
rect 25054 30297 25106 30306
rect 25054 30263 25063 30297
rect 25063 30263 25097 30297
rect 25097 30263 25106 30297
rect 25054 30254 25106 30263
rect 25214 30297 25266 30306
rect 25214 30263 25223 30297
rect 25223 30263 25257 30297
rect 25257 30263 25266 30297
rect 25214 30254 25266 30263
rect 25374 30297 25426 30306
rect 25374 30263 25383 30297
rect 25383 30263 25417 30297
rect 25417 30263 25426 30297
rect 25374 30254 25426 30263
rect 25534 30297 25586 30306
rect 25534 30263 25543 30297
rect 25543 30263 25577 30297
rect 25577 30263 25586 30297
rect 25534 30254 25586 30263
rect 25694 30297 25746 30306
rect 25694 30263 25703 30297
rect 25703 30263 25737 30297
rect 25737 30263 25746 30297
rect 25694 30254 25746 30263
rect 25854 30297 25906 30306
rect 25854 30263 25863 30297
rect 25863 30263 25897 30297
rect 25897 30263 25906 30297
rect 25854 30254 25906 30263
rect 26014 30297 26066 30306
rect 26014 30263 26023 30297
rect 26023 30263 26057 30297
rect 26057 30263 26066 30297
rect 26014 30254 26066 30263
rect 26174 30297 26226 30306
rect 26174 30263 26183 30297
rect 26183 30263 26217 30297
rect 26217 30263 26226 30297
rect 26174 30254 26226 30263
rect 26334 30297 26386 30306
rect 26334 30263 26343 30297
rect 26343 30263 26377 30297
rect 26377 30263 26386 30297
rect 26334 30254 26386 30263
rect 26494 30297 26546 30306
rect 26494 30263 26503 30297
rect 26503 30263 26537 30297
rect 26537 30263 26546 30297
rect 26494 30254 26546 30263
rect 26654 30297 26706 30306
rect 26654 30263 26663 30297
rect 26663 30263 26697 30297
rect 26697 30263 26706 30297
rect 26654 30254 26706 30263
rect 26814 30297 26866 30306
rect 26814 30263 26823 30297
rect 26823 30263 26857 30297
rect 26857 30263 26866 30297
rect 26814 30254 26866 30263
rect 26974 30297 27026 30306
rect 26974 30263 26983 30297
rect 26983 30263 27017 30297
rect 27017 30263 27026 30297
rect 26974 30254 27026 30263
rect 27134 30297 27186 30306
rect 27134 30263 27143 30297
rect 27143 30263 27177 30297
rect 27177 30263 27186 30297
rect 27134 30254 27186 30263
rect 27294 30297 27346 30306
rect 27294 30263 27303 30297
rect 27303 30263 27337 30297
rect 27337 30263 27346 30297
rect 27294 30254 27346 30263
rect 27454 30297 27506 30306
rect 27454 30263 27463 30297
rect 27463 30263 27497 30297
rect 27497 30263 27506 30297
rect 27454 30254 27506 30263
rect 27614 30297 27666 30306
rect 27614 30263 27623 30297
rect 27623 30263 27657 30297
rect 27657 30263 27666 30297
rect 27614 30254 27666 30263
rect 27774 30297 27826 30306
rect 27774 30263 27783 30297
rect 27783 30263 27817 30297
rect 27817 30263 27826 30297
rect 27774 30254 27826 30263
rect 27934 30297 27986 30306
rect 27934 30263 27943 30297
rect 27943 30263 27977 30297
rect 27977 30263 27986 30297
rect 27934 30254 27986 30263
rect 28094 30297 28146 30306
rect 28094 30263 28103 30297
rect 28103 30263 28137 30297
rect 28137 30263 28146 30297
rect 28094 30254 28146 30263
rect 28254 30297 28306 30306
rect 28254 30263 28263 30297
rect 28263 30263 28297 30297
rect 28297 30263 28306 30297
rect 28254 30254 28306 30263
rect 28414 30297 28466 30306
rect 28414 30263 28423 30297
rect 28423 30263 28457 30297
rect 28457 30263 28466 30297
rect 28414 30254 28466 30263
rect 28574 30297 28626 30306
rect 28574 30263 28583 30297
rect 28583 30263 28617 30297
rect 28617 30263 28626 30297
rect 28574 30254 28626 30263
rect 28734 30297 28786 30306
rect 28734 30263 28743 30297
rect 28743 30263 28777 30297
rect 28777 30263 28786 30297
rect 28734 30254 28786 30263
rect 28894 30297 28946 30306
rect 28894 30263 28903 30297
rect 28903 30263 28937 30297
rect 28937 30263 28946 30297
rect 28894 30254 28946 30263
rect 29054 30297 29106 30306
rect 29054 30263 29063 30297
rect 29063 30263 29097 30297
rect 29097 30263 29106 30297
rect 29054 30254 29106 30263
rect 29214 30297 29266 30306
rect 29214 30263 29223 30297
rect 29223 30263 29257 30297
rect 29257 30263 29266 30297
rect 29214 30254 29266 30263
rect 29374 30297 29426 30306
rect 29374 30263 29383 30297
rect 29383 30263 29417 30297
rect 29417 30263 29426 30297
rect 29374 30254 29426 30263
rect 33534 30297 33586 30306
rect 33534 30263 33543 30297
rect 33543 30263 33577 30297
rect 33577 30263 33586 30297
rect 33534 30254 33586 30263
rect 33694 30297 33746 30306
rect 33694 30263 33703 30297
rect 33703 30263 33737 30297
rect 33737 30263 33746 30297
rect 33694 30254 33746 30263
rect 33854 30297 33906 30306
rect 33854 30263 33863 30297
rect 33863 30263 33897 30297
rect 33897 30263 33906 30297
rect 33854 30254 33906 30263
rect 34014 30297 34066 30306
rect 34014 30263 34023 30297
rect 34023 30263 34057 30297
rect 34057 30263 34066 30297
rect 34014 30254 34066 30263
rect 34174 30297 34226 30306
rect 34174 30263 34183 30297
rect 34183 30263 34217 30297
rect 34217 30263 34226 30297
rect 34174 30254 34226 30263
rect 34334 30297 34386 30306
rect 34334 30263 34343 30297
rect 34343 30263 34377 30297
rect 34377 30263 34386 30297
rect 34334 30254 34386 30263
rect 34494 30297 34546 30306
rect 34494 30263 34503 30297
rect 34503 30263 34537 30297
rect 34537 30263 34546 30297
rect 34494 30254 34546 30263
rect 34654 30297 34706 30306
rect 34654 30263 34663 30297
rect 34663 30263 34697 30297
rect 34697 30263 34706 30297
rect 34654 30254 34706 30263
rect 34814 30297 34866 30306
rect 34814 30263 34823 30297
rect 34823 30263 34857 30297
rect 34857 30263 34866 30297
rect 34814 30254 34866 30263
rect 34974 30297 35026 30306
rect 34974 30263 34983 30297
rect 34983 30263 35017 30297
rect 35017 30263 35026 30297
rect 34974 30254 35026 30263
rect 35134 30297 35186 30306
rect 35134 30263 35143 30297
rect 35143 30263 35177 30297
rect 35177 30263 35186 30297
rect 35134 30254 35186 30263
rect 35294 30297 35346 30306
rect 35294 30263 35303 30297
rect 35303 30263 35337 30297
rect 35337 30263 35346 30297
rect 35294 30254 35346 30263
rect 35454 30297 35506 30306
rect 35454 30263 35463 30297
rect 35463 30263 35497 30297
rect 35497 30263 35506 30297
rect 35454 30254 35506 30263
rect 35614 30297 35666 30306
rect 35614 30263 35623 30297
rect 35623 30263 35657 30297
rect 35657 30263 35666 30297
rect 35614 30254 35666 30263
rect 35774 30297 35826 30306
rect 35774 30263 35783 30297
rect 35783 30263 35817 30297
rect 35817 30263 35826 30297
rect 35774 30254 35826 30263
rect 35934 30297 35986 30306
rect 35934 30263 35943 30297
rect 35943 30263 35977 30297
rect 35977 30263 35986 30297
rect 35934 30254 35986 30263
rect 36094 30297 36146 30306
rect 36094 30263 36103 30297
rect 36103 30263 36137 30297
rect 36137 30263 36146 30297
rect 36094 30254 36146 30263
rect 36254 30297 36306 30306
rect 36254 30263 36263 30297
rect 36263 30263 36297 30297
rect 36297 30263 36306 30297
rect 36254 30254 36306 30263
rect 36414 30297 36466 30306
rect 36414 30263 36423 30297
rect 36423 30263 36457 30297
rect 36457 30263 36466 30297
rect 36414 30254 36466 30263
rect 36574 30297 36626 30306
rect 36574 30263 36583 30297
rect 36583 30263 36617 30297
rect 36617 30263 36626 30297
rect 36574 30254 36626 30263
rect 36734 30297 36786 30306
rect 36734 30263 36743 30297
rect 36743 30263 36777 30297
rect 36777 30263 36786 30297
rect 36734 30254 36786 30263
rect 36894 30297 36946 30306
rect 36894 30263 36903 30297
rect 36903 30263 36937 30297
rect 36937 30263 36946 30297
rect 36894 30254 36946 30263
rect 37054 30297 37106 30306
rect 37054 30263 37063 30297
rect 37063 30263 37097 30297
rect 37097 30263 37106 30297
rect 37054 30254 37106 30263
rect 37214 30297 37266 30306
rect 37214 30263 37223 30297
rect 37223 30263 37257 30297
rect 37257 30263 37266 30297
rect 37214 30254 37266 30263
rect 37374 30297 37426 30306
rect 37374 30263 37383 30297
rect 37383 30263 37417 30297
rect 37417 30263 37426 30297
rect 37374 30254 37426 30263
rect 37534 30297 37586 30306
rect 37534 30263 37543 30297
rect 37543 30263 37577 30297
rect 37577 30263 37586 30297
rect 37534 30254 37586 30263
rect 37694 30297 37746 30306
rect 37694 30263 37703 30297
rect 37703 30263 37737 30297
rect 37737 30263 37746 30297
rect 37694 30254 37746 30263
rect 37854 30297 37906 30306
rect 37854 30263 37863 30297
rect 37863 30263 37897 30297
rect 37897 30263 37906 30297
rect 37854 30254 37906 30263
rect 38014 30297 38066 30306
rect 38014 30263 38023 30297
rect 38023 30263 38057 30297
rect 38057 30263 38066 30297
rect 38014 30254 38066 30263
rect 38174 30297 38226 30306
rect 38174 30263 38183 30297
rect 38183 30263 38217 30297
rect 38217 30263 38226 30297
rect 38174 30254 38226 30263
rect 38334 30297 38386 30306
rect 38334 30263 38343 30297
rect 38343 30263 38377 30297
rect 38377 30263 38386 30297
rect 38334 30254 38386 30263
rect 38494 30297 38546 30306
rect 38494 30263 38503 30297
rect 38503 30263 38537 30297
rect 38537 30263 38546 30297
rect 38494 30254 38546 30263
rect 38654 30297 38706 30306
rect 38654 30263 38663 30297
rect 38663 30263 38697 30297
rect 38697 30263 38706 30297
rect 38654 30254 38706 30263
rect 38814 30297 38866 30306
rect 38814 30263 38823 30297
rect 38823 30263 38857 30297
rect 38857 30263 38866 30297
rect 38814 30254 38866 30263
rect 38974 30297 39026 30306
rect 38974 30263 38983 30297
rect 38983 30263 39017 30297
rect 39017 30263 39026 30297
rect 38974 30254 39026 30263
rect 39134 30297 39186 30306
rect 39134 30263 39143 30297
rect 39143 30263 39177 30297
rect 39177 30263 39186 30297
rect 39134 30254 39186 30263
rect 39294 30297 39346 30306
rect 39294 30263 39303 30297
rect 39303 30263 39337 30297
rect 39337 30263 39346 30297
rect 39294 30254 39346 30263
rect 39454 30297 39506 30306
rect 39454 30263 39463 30297
rect 39463 30263 39497 30297
rect 39497 30263 39506 30297
rect 39454 30254 39506 30263
rect 39614 30297 39666 30306
rect 39614 30263 39623 30297
rect 39623 30263 39657 30297
rect 39657 30263 39666 30297
rect 39614 30254 39666 30263
rect 39774 30297 39826 30306
rect 39774 30263 39783 30297
rect 39783 30263 39817 30297
rect 39817 30263 39826 30297
rect 39774 30254 39826 30263
rect 39934 30297 39986 30306
rect 39934 30263 39943 30297
rect 39943 30263 39977 30297
rect 39977 30263 39986 30297
rect 39934 30254 39986 30263
rect 40094 30297 40146 30306
rect 40094 30263 40103 30297
rect 40103 30263 40137 30297
rect 40137 30263 40146 30297
rect 40094 30254 40146 30263
rect 40254 30297 40306 30306
rect 40254 30263 40263 30297
rect 40263 30263 40297 30297
rect 40297 30263 40306 30297
rect 40254 30254 40306 30263
rect 40414 30297 40466 30306
rect 40414 30263 40423 30297
rect 40423 30263 40457 30297
rect 40457 30263 40466 30297
rect 40414 30254 40466 30263
rect 40574 30297 40626 30306
rect 40574 30263 40583 30297
rect 40583 30263 40617 30297
rect 40617 30263 40626 30297
rect 40574 30254 40626 30263
rect 40734 30297 40786 30306
rect 40734 30263 40743 30297
rect 40743 30263 40777 30297
rect 40777 30263 40786 30297
rect 40734 30254 40786 30263
rect 40894 30297 40946 30306
rect 40894 30263 40903 30297
rect 40903 30263 40937 30297
rect 40937 30263 40946 30297
rect 40894 30254 40946 30263
rect 41054 30297 41106 30306
rect 41054 30263 41063 30297
rect 41063 30263 41097 30297
rect 41097 30263 41106 30297
rect 41054 30254 41106 30263
rect 41214 30297 41266 30306
rect 41214 30263 41223 30297
rect 41223 30263 41257 30297
rect 41257 30263 41266 30297
rect 41214 30254 41266 30263
rect 41374 30297 41426 30306
rect 41374 30263 41383 30297
rect 41383 30263 41417 30297
rect 41417 30263 41426 30297
rect 41374 30254 41426 30263
rect 41534 30297 41586 30306
rect 41534 30263 41543 30297
rect 41543 30263 41577 30297
rect 41577 30263 41586 30297
rect 41534 30254 41586 30263
rect 41694 30297 41746 30306
rect 41694 30263 41703 30297
rect 41703 30263 41737 30297
rect 41737 30263 41746 30297
rect 41694 30254 41746 30263
rect 41854 30297 41906 30306
rect 41854 30263 41863 30297
rect 41863 30263 41897 30297
rect 41897 30263 41906 30297
rect 41854 30254 41906 30263
rect 14 29977 66 29986
rect 14 29943 23 29977
rect 23 29943 57 29977
rect 57 29943 66 29977
rect 14 29934 66 29943
rect 174 29977 226 29986
rect 174 29943 183 29977
rect 183 29943 217 29977
rect 217 29943 226 29977
rect 174 29934 226 29943
rect 334 29977 386 29986
rect 334 29943 343 29977
rect 343 29943 377 29977
rect 377 29943 386 29977
rect 334 29934 386 29943
rect 494 29977 546 29986
rect 494 29943 503 29977
rect 503 29943 537 29977
rect 537 29943 546 29977
rect 494 29934 546 29943
rect 654 29977 706 29986
rect 654 29943 663 29977
rect 663 29943 697 29977
rect 697 29943 706 29977
rect 654 29934 706 29943
rect 814 29977 866 29986
rect 814 29943 823 29977
rect 823 29943 857 29977
rect 857 29943 866 29977
rect 814 29934 866 29943
rect 974 29977 1026 29986
rect 974 29943 983 29977
rect 983 29943 1017 29977
rect 1017 29943 1026 29977
rect 974 29934 1026 29943
rect 1134 29977 1186 29986
rect 1134 29943 1143 29977
rect 1143 29943 1177 29977
rect 1177 29943 1186 29977
rect 1134 29934 1186 29943
rect 1294 29977 1346 29986
rect 1294 29943 1303 29977
rect 1303 29943 1337 29977
rect 1337 29943 1346 29977
rect 1294 29934 1346 29943
rect 1454 29977 1506 29986
rect 1454 29943 1463 29977
rect 1463 29943 1497 29977
rect 1497 29943 1506 29977
rect 1454 29934 1506 29943
rect 1614 29977 1666 29986
rect 1614 29943 1623 29977
rect 1623 29943 1657 29977
rect 1657 29943 1666 29977
rect 1614 29934 1666 29943
rect 1774 29977 1826 29986
rect 1774 29943 1783 29977
rect 1783 29943 1817 29977
rect 1817 29943 1826 29977
rect 1774 29934 1826 29943
rect 1934 29977 1986 29986
rect 1934 29943 1943 29977
rect 1943 29943 1977 29977
rect 1977 29943 1986 29977
rect 1934 29934 1986 29943
rect 2094 29977 2146 29986
rect 2094 29943 2103 29977
rect 2103 29943 2137 29977
rect 2137 29943 2146 29977
rect 2094 29934 2146 29943
rect 2254 29977 2306 29986
rect 2254 29943 2263 29977
rect 2263 29943 2297 29977
rect 2297 29943 2306 29977
rect 2254 29934 2306 29943
rect 2414 29977 2466 29986
rect 2414 29943 2423 29977
rect 2423 29943 2457 29977
rect 2457 29943 2466 29977
rect 2414 29934 2466 29943
rect 2574 29977 2626 29986
rect 2574 29943 2583 29977
rect 2583 29943 2617 29977
rect 2617 29943 2626 29977
rect 2574 29934 2626 29943
rect 2734 29977 2786 29986
rect 2734 29943 2743 29977
rect 2743 29943 2777 29977
rect 2777 29943 2786 29977
rect 2734 29934 2786 29943
rect 2894 29977 2946 29986
rect 2894 29943 2903 29977
rect 2903 29943 2937 29977
rect 2937 29943 2946 29977
rect 2894 29934 2946 29943
rect 3054 29977 3106 29986
rect 3054 29943 3063 29977
rect 3063 29943 3097 29977
rect 3097 29943 3106 29977
rect 3054 29934 3106 29943
rect 3214 29977 3266 29986
rect 3214 29943 3223 29977
rect 3223 29943 3257 29977
rect 3257 29943 3266 29977
rect 3214 29934 3266 29943
rect 3374 29977 3426 29986
rect 3374 29943 3383 29977
rect 3383 29943 3417 29977
rect 3417 29943 3426 29977
rect 3374 29934 3426 29943
rect 3534 29977 3586 29986
rect 3534 29943 3543 29977
rect 3543 29943 3577 29977
rect 3577 29943 3586 29977
rect 3534 29934 3586 29943
rect 3694 29977 3746 29986
rect 3694 29943 3703 29977
rect 3703 29943 3737 29977
rect 3737 29943 3746 29977
rect 3694 29934 3746 29943
rect 3854 29977 3906 29986
rect 3854 29943 3863 29977
rect 3863 29943 3897 29977
rect 3897 29943 3906 29977
rect 3854 29934 3906 29943
rect 4014 29977 4066 29986
rect 4014 29943 4023 29977
rect 4023 29943 4057 29977
rect 4057 29943 4066 29977
rect 4014 29934 4066 29943
rect 4174 29977 4226 29986
rect 4174 29943 4183 29977
rect 4183 29943 4217 29977
rect 4217 29943 4226 29977
rect 4174 29934 4226 29943
rect 4334 29977 4386 29986
rect 4334 29943 4343 29977
rect 4343 29943 4377 29977
rect 4377 29943 4386 29977
rect 4334 29934 4386 29943
rect 4494 29977 4546 29986
rect 4494 29943 4503 29977
rect 4503 29943 4537 29977
rect 4537 29943 4546 29977
rect 4494 29934 4546 29943
rect 4654 29977 4706 29986
rect 4654 29943 4663 29977
rect 4663 29943 4697 29977
rect 4697 29943 4706 29977
rect 4654 29934 4706 29943
rect 4814 29977 4866 29986
rect 4814 29943 4823 29977
rect 4823 29943 4857 29977
rect 4857 29943 4866 29977
rect 4814 29934 4866 29943
rect 4974 29977 5026 29986
rect 4974 29943 4983 29977
rect 4983 29943 5017 29977
rect 5017 29943 5026 29977
rect 4974 29934 5026 29943
rect 5134 29977 5186 29986
rect 5134 29943 5143 29977
rect 5143 29943 5177 29977
rect 5177 29943 5186 29977
rect 5134 29934 5186 29943
rect 5294 29977 5346 29986
rect 5294 29943 5303 29977
rect 5303 29943 5337 29977
rect 5337 29943 5346 29977
rect 5294 29934 5346 29943
rect 5454 29977 5506 29986
rect 5454 29943 5463 29977
rect 5463 29943 5497 29977
rect 5497 29943 5506 29977
rect 5454 29934 5506 29943
rect 5614 29977 5666 29986
rect 5614 29943 5623 29977
rect 5623 29943 5657 29977
rect 5657 29943 5666 29977
rect 5614 29934 5666 29943
rect 5774 29977 5826 29986
rect 5774 29943 5783 29977
rect 5783 29943 5817 29977
rect 5817 29943 5826 29977
rect 5774 29934 5826 29943
rect 5934 29977 5986 29986
rect 5934 29943 5943 29977
rect 5943 29943 5977 29977
rect 5977 29943 5986 29977
rect 5934 29934 5986 29943
rect 6094 29977 6146 29986
rect 6094 29943 6103 29977
rect 6103 29943 6137 29977
rect 6137 29943 6146 29977
rect 6094 29934 6146 29943
rect 6254 29977 6306 29986
rect 6254 29943 6263 29977
rect 6263 29943 6297 29977
rect 6297 29943 6306 29977
rect 6254 29934 6306 29943
rect 6414 29977 6466 29986
rect 6414 29943 6423 29977
rect 6423 29943 6457 29977
rect 6457 29943 6466 29977
rect 6414 29934 6466 29943
rect 6574 29977 6626 29986
rect 6574 29943 6583 29977
rect 6583 29943 6617 29977
rect 6617 29943 6626 29977
rect 6574 29934 6626 29943
rect 6734 29977 6786 29986
rect 6734 29943 6743 29977
rect 6743 29943 6777 29977
rect 6777 29943 6786 29977
rect 6734 29934 6786 29943
rect 6894 29977 6946 29986
rect 6894 29943 6903 29977
rect 6903 29943 6937 29977
rect 6937 29943 6946 29977
rect 6894 29934 6946 29943
rect 7054 29977 7106 29986
rect 7054 29943 7063 29977
rect 7063 29943 7097 29977
rect 7097 29943 7106 29977
rect 7054 29934 7106 29943
rect 7214 29977 7266 29986
rect 7214 29943 7223 29977
rect 7223 29943 7257 29977
rect 7257 29943 7266 29977
rect 7214 29934 7266 29943
rect 7374 29977 7426 29986
rect 7374 29943 7383 29977
rect 7383 29943 7417 29977
rect 7417 29943 7426 29977
rect 7374 29934 7426 29943
rect 7534 29977 7586 29986
rect 7534 29943 7543 29977
rect 7543 29943 7577 29977
rect 7577 29943 7586 29977
rect 7534 29934 7586 29943
rect 7694 29977 7746 29986
rect 7694 29943 7703 29977
rect 7703 29943 7737 29977
rect 7737 29943 7746 29977
rect 7694 29934 7746 29943
rect 7854 29977 7906 29986
rect 7854 29943 7863 29977
rect 7863 29943 7897 29977
rect 7897 29943 7906 29977
rect 7854 29934 7906 29943
rect 8014 29977 8066 29986
rect 8014 29943 8023 29977
rect 8023 29943 8057 29977
rect 8057 29943 8066 29977
rect 8014 29934 8066 29943
rect 8174 29977 8226 29986
rect 8174 29943 8183 29977
rect 8183 29943 8217 29977
rect 8217 29943 8226 29977
rect 8174 29934 8226 29943
rect 8334 29977 8386 29986
rect 8334 29943 8343 29977
rect 8343 29943 8377 29977
rect 8377 29943 8386 29977
rect 8334 29934 8386 29943
rect 12494 29977 12546 29986
rect 12494 29943 12503 29977
rect 12503 29943 12537 29977
rect 12537 29943 12546 29977
rect 12494 29934 12546 29943
rect 12654 29977 12706 29986
rect 12654 29943 12663 29977
rect 12663 29943 12697 29977
rect 12697 29943 12706 29977
rect 12654 29934 12706 29943
rect 12814 29977 12866 29986
rect 12814 29943 12823 29977
rect 12823 29943 12857 29977
rect 12857 29943 12866 29977
rect 12814 29934 12866 29943
rect 12974 29977 13026 29986
rect 12974 29943 12983 29977
rect 12983 29943 13017 29977
rect 13017 29943 13026 29977
rect 12974 29934 13026 29943
rect 13134 29977 13186 29986
rect 13134 29943 13143 29977
rect 13143 29943 13177 29977
rect 13177 29943 13186 29977
rect 13134 29934 13186 29943
rect 13294 29977 13346 29986
rect 13294 29943 13303 29977
rect 13303 29943 13337 29977
rect 13337 29943 13346 29977
rect 13294 29934 13346 29943
rect 13454 29977 13506 29986
rect 13454 29943 13463 29977
rect 13463 29943 13497 29977
rect 13497 29943 13506 29977
rect 13454 29934 13506 29943
rect 13614 29977 13666 29986
rect 13614 29943 13623 29977
rect 13623 29943 13657 29977
rect 13657 29943 13666 29977
rect 13614 29934 13666 29943
rect 13774 29977 13826 29986
rect 13774 29943 13783 29977
rect 13783 29943 13817 29977
rect 13817 29943 13826 29977
rect 13774 29934 13826 29943
rect 13934 29977 13986 29986
rect 13934 29943 13943 29977
rect 13943 29943 13977 29977
rect 13977 29943 13986 29977
rect 13934 29934 13986 29943
rect 14094 29977 14146 29986
rect 14094 29943 14103 29977
rect 14103 29943 14137 29977
rect 14137 29943 14146 29977
rect 14094 29934 14146 29943
rect 14254 29977 14306 29986
rect 14254 29943 14263 29977
rect 14263 29943 14297 29977
rect 14297 29943 14306 29977
rect 14254 29934 14306 29943
rect 14414 29977 14466 29986
rect 14414 29943 14423 29977
rect 14423 29943 14457 29977
rect 14457 29943 14466 29977
rect 14414 29934 14466 29943
rect 14574 29977 14626 29986
rect 14574 29943 14583 29977
rect 14583 29943 14617 29977
rect 14617 29943 14626 29977
rect 14574 29934 14626 29943
rect 14734 29977 14786 29986
rect 14734 29943 14743 29977
rect 14743 29943 14777 29977
rect 14777 29943 14786 29977
rect 14734 29934 14786 29943
rect 14894 29977 14946 29986
rect 14894 29943 14903 29977
rect 14903 29943 14937 29977
rect 14937 29943 14946 29977
rect 14894 29934 14946 29943
rect 15054 29977 15106 29986
rect 15054 29943 15063 29977
rect 15063 29943 15097 29977
rect 15097 29943 15106 29977
rect 15054 29934 15106 29943
rect 15214 29977 15266 29986
rect 15214 29943 15223 29977
rect 15223 29943 15257 29977
rect 15257 29943 15266 29977
rect 15214 29934 15266 29943
rect 15374 29977 15426 29986
rect 15374 29943 15383 29977
rect 15383 29943 15417 29977
rect 15417 29943 15426 29977
rect 15374 29934 15426 29943
rect 15534 29977 15586 29986
rect 15534 29943 15543 29977
rect 15543 29943 15577 29977
rect 15577 29943 15586 29977
rect 15534 29934 15586 29943
rect 15694 29977 15746 29986
rect 15694 29943 15703 29977
rect 15703 29943 15737 29977
rect 15737 29943 15746 29977
rect 15694 29934 15746 29943
rect 15854 29977 15906 29986
rect 15854 29943 15863 29977
rect 15863 29943 15897 29977
rect 15897 29943 15906 29977
rect 15854 29934 15906 29943
rect 16014 29977 16066 29986
rect 16014 29943 16023 29977
rect 16023 29943 16057 29977
rect 16057 29943 16066 29977
rect 16014 29934 16066 29943
rect 16174 29977 16226 29986
rect 16174 29943 16183 29977
rect 16183 29943 16217 29977
rect 16217 29943 16226 29977
rect 16174 29934 16226 29943
rect 16334 29977 16386 29986
rect 16334 29943 16343 29977
rect 16343 29943 16377 29977
rect 16377 29943 16386 29977
rect 16334 29934 16386 29943
rect 16494 29977 16546 29986
rect 16494 29943 16503 29977
rect 16503 29943 16537 29977
rect 16537 29943 16546 29977
rect 16494 29934 16546 29943
rect 16654 29977 16706 29986
rect 16654 29943 16663 29977
rect 16663 29943 16697 29977
rect 16697 29943 16706 29977
rect 16654 29934 16706 29943
rect 16814 29977 16866 29986
rect 16814 29943 16823 29977
rect 16823 29943 16857 29977
rect 16857 29943 16866 29977
rect 16814 29934 16866 29943
rect 16974 29977 17026 29986
rect 16974 29943 16983 29977
rect 16983 29943 17017 29977
rect 17017 29943 17026 29977
rect 16974 29934 17026 29943
rect 17134 29977 17186 29986
rect 17134 29943 17143 29977
rect 17143 29943 17177 29977
rect 17177 29943 17186 29977
rect 17134 29934 17186 29943
rect 17294 29977 17346 29986
rect 17294 29943 17303 29977
rect 17303 29943 17337 29977
rect 17337 29943 17346 29977
rect 17294 29934 17346 29943
rect 17454 29977 17506 29986
rect 17454 29943 17463 29977
rect 17463 29943 17497 29977
rect 17497 29943 17506 29977
rect 17454 29934 17506 29943
rect 17614 29977 17666 29986
rect 17614 29943 17623 29977
rect 17623 29943 17657 29977
rect 17657 29943 17666 29977
rect 17614 29934 17666 29943
rect 17774 29977 17826 29986
rect 17774 29943 17783 29977
rect 17783 29943 17817 29977
rect 17817 29943 17826 29977
rect 17774 29934 17826 29943
rect 17934 29977 17986 29986
rect 17934 29943 17943 29977
rect 17943 29943 17977 29977
rect 17977 29943 17986 29977
rect 17934 29934 17986 29943
rect 18094 29977 18146 29986
rect 18094 29943 18103 29977
rect 18103 29943 18137 29977
rect 18137 29943 18146 29977
rect 18094 29934 18146 29943
rect 18254 29977 18306 29986
rect 18254 29943 18263 29977
rect 18263 29943 18297 29977
rect 18297 29943 18306 29977
rect 18254 29934 18306 29943
rect 18414 29977 18466 29986
rect 18414 29943 18423 29977
rect 18423 29943 18457 29977
rect 18457 29943 18466 29977
rect 18414 29934 18466 29943
rect 18574 29977 18626 29986
rect 18574 29943 18583 29977
rect 18583 29943 18617 29977
rect 18617 29943 18626 29977
rect 18574 29934 18626 29943
rect 18734 29977 18786 29986
rect 18734 29943 18743 29977
rect 18743 29943 18777 29977
rect 18777 29943 18786 29977
rect 18734 29934 18786 29943
rect 18894 29977 18946 29986
rect 18894 29943 18903 29977
rect 18903 29943 18937 29977
rect 18937 29943 18946 29977
rect 18894 29934 18946 29943
rect 23134 29977 23186 29986
rect 23134 29943 23143 29977
rect 23143 29943 23177 29977
rect 23177 29943 23186 29977
rect 23134 29934 23186 29943
rect 23294 29977 23346 29986
rect 23294 29943 23303 29977
rect 23303 29943 23337 29977
rect 23337 29943 23346 29977
rect 23294 29934 23346 29943
rect 23454 29977 23506 29986
rect 23454 29943 23463 29977
rect 23463 29943 23497 29977
rect 23497 29943 23506 29977
rect 23454 29934 23506 29943
rect 23614 29977 23666 29986
rect 23614 29943 23623 29977
rect 23623 29943 23657 29977
rect 23657 29943 23666 29977
rect 23614 29934 23666 29943
rect 23774 29977 23826 29986
rect 23774 29943 23783 29977
rect 23783 29943 23817 29977
rect 23817 29943 23826 29977
rect 23774 29934 23826 29943
rect 23934 29977 23986 29986
rect 23934 29943 23943 29977
rect 23943 29943 23977 29977
rect 23977 29943 23986 29977
rect 23934 29934 23986 29943
rect 24094 29977 24146 29986
rect 24094 29943 24103 29977
rect 24103 29943 24137 29977
rect 24137 29943 24146 29977
rect 24094 29934 24146 29943
rect 24254 29977 24306 29986
rect 24254 29943 24263 29977
rect 24263 29943 24297 29977
rect 24297 29943 24306 29977
rect 24254 29934 24306 29943
rect 24414 29977 24466 29986
rect 24414 29943 24423 29977
rect 24423 29943 24457 29977
rect 24457 29943 24466 29977
rect 24414 29934 24466 29943
rect 24574 29977 24626 29986
rect 24574 29943 24583 29977
rect 24583 29943 24617 29977
rect 24617 29943 24626 29977
rect 24574 29934 24626 29943
rect 24734 29977 24786 29986
rect 24734 29943 24743 29977
rect 24743 29943 24777 29977
rect 24777 29943 24786 29977
rect 24734 29934 24786 29943
rect 24894 29977 24946 29986
rect 24894 29943 24903 29977
rect 24903 29943 24937 29977
rect 24937 29943 24946 29977
rect 24894 29934 24946 29943
rect 25054 29977 25106 29986
rect 25054 29943 25063 29977
rect 25063 29943 25097 29977
rect 25097 29943 25106 29977
rect 25054 29934 25106 29943
rect 25214 29977 25266 29986
rect 25214 29943 25223 29977
rect 25223 29943 25257 29977
rect 25257 29943 25266 29977
rect 25214 29934 25266 29943
rect 25374 29977 25426 29986
rect 25374 29943 25383 29977
rect 25383 29943 25417 29977
rect 25417 29943 25426 29977
rect 25374 29934 25426 29943
rect 25534 29977 25586 29986
rect 25534 29943 25543 29977
rect 25543 29943 25577 29977
rect 25577 29943 25586 29977
rect 25534 29934 25586 29943
rect 25694 29977 25746 29986
rect 25694 29943 25703 29977
rect 25703 29943 25737 29977
rect 25737 29943 25746 29977
rect 25694 29934 25746 29943
rect 25854 29977 25906 29986
rect 25854 29943 25863 29977
rect 25863 29943 25897 29977
rect 25897 29943 25906 29977
rect 25854 29934 25906 29943
rect 26014 29977 26066 29986
rect 26014 29943 26023 29977
rect 26023 29943 26057 29977
rect 26057 29943 26066 29977
rect 26014 29934 26066 29943
rect 26174 29977 26226 29986
rect 26174 29943 26183 29977
rect 26183 29943 26217 29977
rect 26217 29943 26226 29977
rect 26174 29934 26226 29943
rect 26334 29977 26386 29986
rect 26334 29943 26343 29977
rect 26343 29943 26377 29977
rect 26377 29943 26386 29977
rect 26334 29934 26386 29943
rect 26494 29977 26546 29986
rect 26494 29943 26503 29977
rect 26503 29943 26537 29977
rect 26537 29943 26546 29977
rect 26494 29934 26546 29943
rect 26654 29977 26706 29986
rect 26654 29943 26663 29977
rect 26663 29943 26697 29977
rect 26697 29943 26706 29977
rect 26654 29934 26706 29943
rect 26814 29977 26866 29986
rect 26814 29943 26823 29977
rect 26823 29943 26857 29977
rect 26857 29943 26866 29977
rect 26814 29934 26866 29943
rect 26974 29977 27026 29986
rect 26974 29943 26983 29977
rect 26983 29943 27017 29977
rect 27017 29943 27026 29977
rect 26974 29934 27026 29943
rect 27134 29977 27186 29986
rect 27134 29943 27143 29977
rect 27143 29943 27177 29977
rect 27177 29943 27186 29977
rect 27134 29934 27186 29943
rect 27294 29977 27346 29986
rect 27294 29943 27303 29977
rect 27303 29943 27337 29977
rect 27337 29943 27346 29977
rect 27294 29934 27346 29943
rect 27454 29977 27506 29986
rect 27454 29943 27463 29977
rect 27463 29943 27497 29977
rect 27497 29943 27506 29977
rect 27454 29934 27506 29943
rect 27614 29977 27666 29986
rect 27614 29943 27623 29977
rect 27623 29943 27657 29977
rect 27657 29943 27666 29977
rect 27614 29934 27666 29943
rect 27774 29977 27826 29986
rect 27774 29943 27783 29977
rect 27783 29943 27817 29977
rect 27817 29943 27826 29977
rect 27774 29934 27826 29943
rect 27934 29977 27986 29986
rect 27934 29943 27943 29977
rect 27943 29943 27977 29977
rect 27977 29943 27986 29977
rect 27934 29934 27986 29943
rect 28094 29977 28146 29986
rect 28094 29943 28103 29977
rect 28103 29943 28137 29977
rect 28137 29943 28146 29977
rect 28094 29934 28146 29943
rect 28254 29977 28306 29986
rect 28254 29943 28263 29977
rect 28263 29943 28297 29977
rect 28297 29943 28306 29977
rect 28254 29934 28306 29943
rect 28414 29977 28466 29986
rect 28414 29943 28423 29977
rect 28423 29943 28457 29977
rect 28457 29943 28466 29977
rect 28414 29934 28466 29943
rect 28574 29977 28626 29986
rect 28574 29943 28583 29977
rect 28583 29943 28617 29977
rect 28617 29943 28626 29977
rect 28574 29934 28626 29943
rect 28734 29977 28786 29986
rect 28734 29943 28743 29977
rect 28743 29943 28777 29977
rect 28777 29943 28786 29977
rect 28734 29934 28786 29943
rect 28894 29977 28946 29986
rect 28894 29943 28903 29977
rect 28903 29943 28937 29977
rect 28937 29943 28946 29977
rect 28894 29934 28946 29943
rect 29054 29977 29106 29986
rect 29054 29943 29063 29977
rect 29063 29943 29097 29977
rect 29097 29943 29106 29977
rect 29054 29934 29106 29943
rect 29214 29977 29266 29986
rect 29214 29943 29223 29977
rect 29223 29943 29257 29977
rect 29257 29943 29266 29977
rect 29214 29934 29266 29943
rect 29374 29977 29426 29986
rect 29374 29943 29383 29977
rect 29383 29943 29417 29977
rect 29417 29943 29426 29977
rect 29374 29934 29426 29943
rect 33534 29977 33586 29986
rect 33534 29943 33543 29977
rect 33543 29943 33577 29977
rect 33577 29943 33586 29977
rect 33534 29934 33586 29943
rect 33694 29977 33746 29986
rect 33694 29943 33703 29977
rect 33703 29943 33737 29977
rect 33737 29943 33746 29977
rect 33694 29934 33746 29943
rect 33854 29977 33906 29986
rect 33854 29943 33863 29977
rect 33863 29943 33897 29977
rect 33897 29943 33906 29977
rect 33854 29934 33906 29943
rect 34014 29977 34066 29986
rect 34014 29943 34023 29977
rect 34023 29943 34057 29977
rect 34057 29943 34066 29977
rect 34014 29934 34066 29943
rect 34174 29977 34226 29986
rect 34174 29943 34183 29977
rect 34183 29943 34217 29977
rect 34217 29943 34226 29977
rect 34174 29934 34226 29943
rect 34334 29977 34386 29986
rect 34334 29943 34343 29977
rect 34343 29943 34377 29977
rect 34377 29943 34386 29977
rect 34334 29934 34386 29943
rect 34494 29977 34546 29986
rect 34494 29943 34503 29977
rect 34503 29943 34537 29977
rect 34537 29943 34546 29977
rect 34494 29934 34546 29943
rect 34654 29977 34706 29986
rect 34654 29943 34663 29977
rect 34663 29943 34697 29977
rect 34697 29943 34706 29977
rect 34654 29934 34706 29943
rect 34814 29977 34866 29986
rect 34814 29943 34823 29977
rect 34823 29943 34857 29977
rect 34857 29943 34866 29977
rect 34814 29934 34866 29943
rect 34974 29977 35026 29986
rect 34974 29943 34983 29977
rect 34983 29943 35017 29977
rect 35017 29943 35026 29977
rect 34974 29934 35026 29943
rect 35134 29977 35186 29986
rect 35134 29943 35143 29977
rect 35143 29943 35177 29977
rect 35177 29943 35186 29977
rect 35134 29934 35186 29943
rect 35294 29977 35346 29986
rect 35294 29943 35303 29977
rect 35303 29943 35337 29977
rect 35337 29943 35346 29977
rect 35294 29934 35346 29943
rect 35454 29977 35506 29986
rect 35454 29943 35463 29977
rect 35463 29943 35497 29977
rect 35497 29943 35506 29977
rect 35454 29934 35506 29943
rect 35614 29977 35666 29986
rect 35614 29943 35623 29977
rect 35623 29943 35657 29977
rect 35657 29943 35666 29977
rect 35614 29934 35666 29943
rect 35774 29977 35826 29986
rect 35774 29943 35783 29977
rect 35783 29943 35817 29977
rect 35817 29943 35826 29977
rect 35774 29934 35826 29943
rect 35934 29977 35986 29986
rect 35934 29943 35943 29977
rect 35943 29943 35977 29977
rect 35977 29943 35986 29977
rect 35934 29934 35986 29943
rect 36094 29977 36146 29986
rect 36094 29943 36103 29977
rect 36103 29943 36137 29977
rect 36137 29943 36146 29977
rect 36094 29934 36146 29943
rect 36254 29977 36306 29986
rect 36254 29943 36263 29977
rect 36263 29943 36297 29977
rect 36297 29943 36306 29977
rect 36254 29934 36306 29943
rect 36414 29977 36466 29986
rect 36414 29943 36423 29977
rect 36423 29943 36457 29977
rect 36457 29943 36466 29977
rect 36414 29934 36466 29943
rect 36574 29977 36626 29986
rect 36574 29943 36583 29977
rect 36583 29943 36617 29977
rect 36617 29943 36626 29977
rect 36574 29934 36626 29943
rect 36734 29977 36786 29986
rect 36734 29943 36743 29977
rect 36743 29943 36777 29977
rect 36777 29943 36786 29977
rect 36734 29934 36786 29943
rect 36894 29977 36946 29986
rect 36894 29943 36903 29977
rect 36903 29943 36937 29977
rect 36937 29943 36946 29977
rect 36894 29934 36946 29943
rect 37054 29977 37106 29986
rect 37054 29943 37063 29977
rect 37063 29943 37097 29977
rect 37097 29943 37106 29977
rect 37054 29934 37106 29943
rect 37214 29977 37266 29986
rect 37214 29943 37223 29977
rect 37223 29943 37257 29977
rect 37257 29943 37266 29977
rect 37214 29934 37266 29943
rect 37374 29977 37426 29986
rect 37374 29943 37383 29977
rect 37383 29943 37417 29977
rect 37417 29943 37426 29977
rect 37374 29934 37426 29943
rect 37534 29977 37586 29986
rect 37534 29943 37543 29977
rect 37543 29943 37577 29977
rect 37577 29943 37586 29977
rect 37534 29934 37586 29943
rect 37694 29977 37746 29986
rect 37694 29943 37703 29977
rect 37703 29943 37737 29977
rect 37737 29943 37746 29977
rect 37694 29934 37746 29943
rect 37854 29977 37906 29986
rect 37854 29943 37863 29977
rect 37863 29943 37897 29977
rect 37897 29943 37906 29977
rect 37854 29934 37906 29943
rect 38014 29977 38066 29986
rect 38014 29943 38023 29977
rect 38023 29943 38057 29977
rect 38057 29943 38066 29977
rect 38014 29934 38066 29943
rect 38174 29977 38226 29986
rect 38174 29943 38183 29977
rect 38183 29943 38217 29977
rect 38217 29943 38226 29977
rect 38174 29934 38226 29943
rect 38334 29977 38386 29986
rect 38334 29943 38343 29977
rect 38343 29943 38377 29977
rect 38377 29943 38386 29977
rect 38334 29934 38386 29943
rect 38494 29977 38546 29986
rect 38494 29943 38503 29977
rect 38503 29943 38537 29977
rect 38537 29943 38546 29977
rect 38494 29934 38546 29943
rect 38654 29977 38706 29986
rect 38654 29943 38663 29977
rect 38663 29943 38697 29977
rect 38697 29943 38706 29977
rect 38654 29934 38706 29943
rect 38814 29977 38866 29986
rect 38814 29943 38823 29977
rect 38823 29943 38857 29977
rect 38857 29943 38866 29977
rect 38814 29934 38866 29943
rect 38974 29977 39026 29986
rect 38974 29943 38983 29977
rect 38983 29943 39017 29977
rect 39017 29943 39026 29977
rect 38974 29934 39026 29943
rect 39134 29977 39186 29986
rect 39134 29943 39143 29977
rect 39143 29943 39177 29977
rect 39177 29943 39186 29977
rect 39134 29934 39186 29943
rect 39294 29977 39346 29986
rect 39294 29943 39303 29977
rect 39303 29943 39337 29977
rect 39337 29943 39346 29977
rect 39294 29934 39346 29943
rect 39454 29977 39506 29986
rect 39454 29943 39463 29977
rect 39463 29943 39497 29977
rect 39497 29943 39506 29977
rect 39454 29934 39506 29943
rect 39614 29977 39666 29986
rect 39614 29943 39623 29977
rect 39623 29943 39657 29977
rect 39657 29943 39666 29977
rect 39614 29934 39666 29943
rect 39774 29977 39826 29986
rect 39774 29943 39783 29977
rect 39783 29943 39817 29977
rect 39817 29943 39826 29977
rect 39774 29934 39826 29943
rect 39934 29977 39986 29986
rect 39934 29943 39943 29977
rect 39943 29943 39977 29977
rect 39977 29943 39986 29977
rect 39934 29934 39986 29943
rect 40094 29977 40146 29986
rect 40094 29943 40103 29977
rect 40103 29943 40137 29977
rect 40137 29943 40146 29977
rect 40094 29934 40146 29943
rect 40254 29977 40306 29986
rect 40254 29943 40263 29977
rect 40263 29943 40297 29977
rect 40297 29943 40306 29977
rect 40254 29934 40306 29943
rect 40414 29977 40466 29986
rect 40414 29943 40423 29977
rect 40423 29943 40457 29977
rect 40457 29943 40466 29977
rect 40414 29934 40466 29943
rect 40574 29977 40626 29986
rect 40574 29943 40583 29977
rect 40583 29943 40617 29977
rect 40617 29943 40626 29977
rect 40574 29934 40626 29943
rect 40734 29977 40786 29986
rect 40734 29943 40743 29977
rect 40743 29943 40777 29977
rect 40777 29943 40786 29977
rect 40734 29934 40786 29943
rect 40894 29977 40946 29986
rect 40894 29943 40903 29977
rect 40903 29943 40937 29977
rect 40937 29943 40946 29977
rect 40894 29934 40946 29943
rect 41054 29977 41106 29986
rect 41054 29943 41063 29977
rect 41063 29943 41097 29977
rect 41097 29943 41106 29977
rect 41054 29934 41106 29943
rect 41214 29977 41266 29986
rect 41214 29943 41223 29977
rect 41223 29943 41257 29977
rect 41257 29943 41266 29977
rect 41214 29934 41266 29943
rect 41374 29977 41426 29986
rect 41374 29943 41383 29977
rect 41383 29943 41417 29977
rect 41417 29943 41426 29977
rect 41374 29934 41426 29943
rect 41534 29977 41586 29986
rect 41534 29943 41543 29977
rect 41543 29943 41577 29977
rect 41577 29943 41586 29977
rect 41534 29934 41586 29943
rect 41694 29977 41746 29986
rect 41694 29943 41703 29977
rect 41703 29943 41737 29977
rect 41737 29943 41746 29977
rect 41694 29934 41746 29943
rect 41854 29977 41906 29986
rect 41854 29943 41863 29977
rect 41863 29943 41897 29977
rect 41897 29943 41906 29977
rect 41854 29934 41906 29943
rect 14 29817 66 29826
rect 14 29783 23 29817
rect 23 29783 57 29817
rect 57 29783 66 29817
rect 14 29774 66 29783
rect 174 29817 226 29826
rect 174 29783 183 29817
rect 183 29783 217 29817
rect 217 29783 226 29817
rect 174 29774 226 29783
rect 334 29817 386 29826
rect 334 29783 343 29817
rect 343 29783 377 29817
rect 377 29783 386 29817
rect 334 29774 386 29783
rect 494 29817 546 29826
rect 494 29783 503 29817
rect 503 29783 537 29817
rect 537 29783 546 29817
rect 494 29774 546 29783
rect 654 29817 706 29826
rect 654 29783 663 29817
rect 663 29783 697 29817
rect 697 29783 706 29817
rect 654 29774 706 29783
rect 814 29817 866 29826
rect 814 29783 823 29817
rect 823 29783 857 29817
rect 857 29783 866 29817
rect 814 29774 866 29783
rect 974 29817 1026 29826
rect 974 29783 983 29817
rect 983 29783 1017 29817
rect 1017 29783 1026 29817
rect 974 29774 1026 29783
rect 1134 29817 1186 29826
rect 1134 29783 1143 29817
rect 1143 29783 1177 29817
rect 1177 29783 1186 29817
rect 1134 29774 1186 29783
rect 1294 29817 1346 29826
rect 1294 29783 1303 29817
rect 1303 29783 1337 29817
rect 1337 29783 1346 29817
rect 1294 29774 1346 29783
rect 1454 29817 1506 29826
rect 1454 29783 1463 29817
rect 1463 29783 1497 29817
rect 1497 29783 1506 29817
rect 1454 29774 1506 29783
rect 1614 29817 1666 29826
rect 1614 29783 1623 29817
rect 1623 29783 1657 29817
rect 1657 29783 1666 29817
rect 1614 29774 1666 29783
rect 1774 29817 1826 29826
rect 1774 29783 1783 29817
rect 1783 29783 1817 29817
rect 1817 29783 1826 29817
rect 1774 29774 1826 29783
rect 1934 29817 1986 29826
rect 1934 29783 1943 29817
rect 1943 29783 1977 29817
rect 1977 29783 1986 29817
rect 1934 29774 1986 29783
rect 2094 29817 2146 29826
rect 2094 29783 2103 29817
rect 2103 29783 2137 29817
rect 2137 29783 2146 29817
rect 2094 29774 2146 29783
rect 2254 29817 2306 29826
rect 2254 29783 2263 29817
rect 2263 29783 2297 29817
rect 2297 29783 2306 29817
rect 2254 29774 2306 29783
rect 2414 29817 2466 29826
rect 2414 29783 2423 29817
rect 2423 29783 2457 29817
rect 2457 29783 2466 29817
rect 2414 29774 2466 29783
rect 2574 29817 2626 29826
rect 2574 29783 2583 29817
rect 2583 29783 2617 29817
rect 2617 29783 2626 29817
rect 2574 29774 2626 29783
rect 2734 29817 2786 29826
rect 2734 29783 2743 29817
rect 2743 29783 2777 29817
rect 2777 29783 2786 29817
rect 2734 29774 2786 29783
rect 2894 29817 2946 29826
rect 2894 29783 2903 29817
rect 2903 29783 2937 29817
rect 2937 29783 2946 29817
rect 2894 29774 2946 29783
rect 3054 29817 3106 29826
rect 3054 29783 3063 29817
rect 3063 29783 3097 29817
rect 3097 29783 3106 29817
rect 3054 29774 3106 29783
rect 3214 29817 3266 29826
rect 3214 29783 3223 29817
rect 3223 29783 3257 29817
rect 3257 29783 3266 29817
rect 3214 29774 3266 29783
rect 3374 29817 3426 29826
rect 3374 29783 3383 29817
rect 3383 29783 3417 29817
rect 3417 29783 3426 29817
rect 3374 29774 3426 29783
rect 3534 29817 3586 29826
rect 3534 29783 3543 29817
rect 3543 29783 3577 29817
rect 3577 29783 3586 29817
rect 3534 29774 3586 29783
rect 3694 29817 3746 29826
rect 3694 29783 3703 29817
rect 3703 29783 3737 29817
rect 3737 29783 3746 29817
rect 3694 29774 3746 29783
rect 3854 29817 3906 29826
rect 3854 29783 3863 29817
rect 3863 29783 3897 29817
rect 3897 29783 3906 29817
rect 3854 29774 3906 29783
rect 4014 29817 4066 29826
rect 4014 29783 4023 29817
rect 4023 29783 4057 29817
rect 4057 29783 4066 29817
rect 4014 29774 4066 29783
rect 4174 29817 4226 29826
rect 4174 29783 4183 29817
rect 4183 29783 4217 29817
rect 4217 29783 4226 29817
rect 4174 29774 4226 29783
rect 4334 29817 4386 29826
rect 4334 29783 4343 29817
rect 4343 29783 4377 29817
rect 4377 29783 4386 29817
rect 4334 29774 4386 29783
rect 4494 29817 4546 29826
rect 4494 29783 4503 29817
rect 4503 29783 4537 29817
rect 4537 29783 4546 29817
rect 4494 29774 4546 29783
rect 4654 29817 4706 29826
rect 4654 29783 4663 29817
rect 4663 29783 4697 29817
rect 4697 29783 4706 29817
rect 4654 29774 4706 29783
rect 4814 29817 4866 29826
rect 4814 29783 4823 29817
rect 4823 29783 4857 29817
rect 4857 29783 4866 29817
rect 4814 29774 4866 29783
rect 4974 29817 5026 29826
rect 4974 29783 4983 29817
rect 4983 29783 5017 29817
rect 5017 29783 5026 29817
rect 4974 29774 5026 29783
rect 5134 29817 5186 29826
rect 5134 29783 5143 29817
rect 5143 29783 5177 29817
rect 5177 29783 5186 29817
rect 5134 29774 5186 29783
rect 5294 29817 5346 29826
rect 5294 29783 5303 29817
rect 5303 29783 5337 29817
rect 5337 29783 5346 29817
rect 5294 29774 5346 29783
rect 5454 29817 5506 29826
rect 5454 29783 5463 29817
rect 5463 29783 5497 29817
rect 5497 29783 5506 29817
rect 5454 29774 5506 29783
rect 5614 29817 5666 29826
rect 5614 29783 5623 29817
rect 5623 29783 5657 29817
rect 5657 29783 5666 29817
rect 5614 29774 5666 29783
rect 5774 29817 5826 29826
rect 5774 29783 5783 29817
rect 5783 29783 5817 29817
rect 5817 29783 5826 29817
rect 5774 29774 5826 29783
rect 5934 29817 5986 29826
rect 5934 29783 5943 29817
rect 5943 29783 5977 29817
rect 5977 29783 5986 29817
rect 5934 29774 5986 29783
rect 6094 29817 6146 29826
rect 6094 29783 6103 29817
rect 6103 29783 6137 29817
rect 6137 29783 6146 29817
rect 6094 29774 6146 29783
rect 6254 29817 6306 29826
rect 6254 29783 6263 29817
rect 6263 29783 6297 29817
rect 6297 29783 6306 29817
rect 6254 29774 6306 29783
rect 6414 29817 6466 29826
rect 6414 29783 6423 29817
rect 6423 29783 6457 29817
rect 6457 29783 6466 29817
rect 6414 29774 6466 29783
rect 6574 29817 6626 29826
rect 6574 29783 6583 29817
rect 6583 29783 6617 29817
rect 6617 29783 6626 29817
rect 6574 29774 6626 29783
rect 6734 29817 6786 29826
rect 6734 29783 6743 29817
rect 6743 29783 6777 29817
rect 6777 29783 6786 29817
rect 6734 29774 6786 29783
rect 6894 29817 6946 29826
rect 6894 29783 6903 29817
rect 6903 29783 6937 29817
rect 6937 29783 6946 29817
rect 6894 29774 6946 29783
rect 7054 29817 7106 29826
rect 7054 29783 7063 29817
rect 7063 29783 7097 29817
rect 7097 29783 7106 29817
rect 7054 29774 7106 29783
rect 7214 29817 7266 29826
rect 7214 29783 7223 29817
rect 7223 29783 7257 29817
rect 7257 29783 7266 29817
rect 7214 29774 7266 29783
rect 7374 29817 7426 29826
rect 7374 29783 7383 29817
rect 7383 29783 7417 29817
rect 7417 29783 7426 29817
rect 7374 29774 7426 29783
rect 7534 29817 7586 29826
rect 7534 29783 7543 29817
rect 7543 29783 7577 29817
rect 7577 29783 7586 29817
rect 7534 29774 7586 29783
rect 7694 29817 7746 29826
rect 7694 29783 7703 29817
rect 7703 29783 7737 29817
rect 7737 29783 7746 29817
rect 7694 29774 7746 29783
rect 7854 29817 7906 29826
rect 7854 29783 7863 29817
rect 7863 29783 7897 29817
rect 7897 29783 7906 29817
rect 7854 29774 7906 29783
rect 8014 29817 8066 29826
rect 8014 29783 8023 29817
rect 8023 29783 8057 29817
rect 8057 29783 8066 29817
rect 8014 29774 8066 29783
rect 8174 29817 8226 29826
rect 8174 29783 8183 29817
rect 8183 29783 8217 29817
rect 8217 29783 8226 29817
rect 8174 29774 8226 29783
rect 8334 29817 8386 29826
rect 8334 29783 8343 29817
rect 8343 29783 8377 29817
rect 8377 29783 8386 29817
rect 8334 29774 8386 29783
rect 12494 29817 12546 29826
rect 12494 29783 12503 29817
rect 12503 29783 12537 29817
rect 12537 29783 12546 29817
rect 12494 29774 12546 29783
rect 12654 29817 12706 29826
rect 12654 29783 12663 29817
rect 12663 29783 12697 29817
rect 12697 29783 12706 29817
rect 12654 29774 12706 29783
rect 12814 29817 12866 29826
rect 12814 29783 12823 29817
rect 12823 29783 12857 29817
rect 12857 29783 12866 29817
rect 12814 29774 12866 29783
rect 12974 29817 13026 29826
rect 12974 29783 12983 29817
rect 12983 29783 13017 29817
rect 13017 29783 13026 29817
rect 12974 29774 13026 29783
rect 13134 29817 13186 29826
rect 13134 29783 13143 29817
rect 13143 29783 13177 29817
rect 13177 29783 13186 29817
rect 13134 29774 13186 29783
rect 13294 29817 13346 29826
rect 13294 29783 13303 29817
rect 13303 29783 13337 29817
rect 13337 29783 13346 29817
rect 13294 29774 13346 29783
rect 13454 29817 13506 29826
rect 13454 29783 13463 29817
rect 13463 29783 13497 29817
rect 13497 29783 13506 29817
rect 13454 29774 13506 29783
rect 13614 29817 13666 29826
rect 13614 29783 13623 29817
rect 13623 29783 13657 29817
rect 13657 29783 13666 29817
rect 13614 29774 13666 29783
rect 13774 29817 13826 29826
rect 13774 29783 13783 29817
rect 13783 29783 13817 29817
rect 13817 29783 13826 29817
rect 13774 29774 13826 29783
rect 13934 29817 13986 29826
rect 13934 29783 13943 29817
rect 13943 29783 13977 29817
rect 13977 29783 13986 29817
rect 13934 29774 13986 29783
rect 14094 29817 14146 29826
rect 14094 29783 14103 29817
rect 14103 29783 14137 29817
rect 14137 29783 14146 29817
rect 14094 29774 14146 29783
rect 14254 29817 14306 29826
rect 14254 29783 14263 29817
rect 14263 29783 14297 29817
rect 14297 29783 14306 29817
rect 14254 29774 14306 29783
rect 14414 29817 14466 29826
rect 14414 29783 14423 29817
rect 14423 29783 14457 29817
rect 14457 29783 14466 29817
rect 14414 29774 14466 29783
rect 14574 29817 14626 29826
rect 14574 29783 14583 29817
rect 14583 29783 14617 29817
rect 14617 29783 14626 29817
rect 14574 29774 14626 29783
rect 14734 29817 14786 29826
rect 14734 29783 14743 29817
rect 14743 29783 14777 29817
rect 14777 29783 14786 29817
rect 14734 29774 14786 29783
rect 14894 29817 14946 29826
rect 14894 29783 14903 29817
rect 14903 29783 14937 29817
rect 14937 29783 14946 29817
rect 14894 29774 14946 29783
rect 15054 29817 15106 29826
rect 15054 29783 15063 29817
rect 15063 29783 15097 29817
rect 15097 29783 15106 29817
rect 15054 29774 15106 29783
rect 15214 29817 15266 29826
rect 15214 29783 15223 29817
rect 15223 29783 15257 29817
rect 15257 29783 15266 29817
rect 15214 29774 15266 29783
rect 15374 29817 15426 29826
rect 15374 29783 15383 29817
rect 15383 29783 15417 29817
rect 15417 29783 15426 29817
rect 15374 29774 15426 29783
rect 15534 29817 15586 29826
rect 15534 29783 15543 29817
rect 15543 29783 15577 29817
rect 15577 29783 15586 29817
rect 15534 29774 15586 29783
rect 15694 29817 15746 29826
rect 15694 29783 15703 29817
rect 15703 29783 15737 29817
rect 15737 29783 15746 29817
rect 15694 29774 15746 29783
rect 15854 29817 15906 29826
rect 15854 29783 15863 29817
rect 15863 29783 15897 29817
rect 15897 29783 15906 29817
rect 15854 29774 15906 29783
rect 16014 29817 16066 29826
rect 16014 29783 16023 29817
rect 16023 29783 16057 29817
rect 16057 29783 16066 29817
rect 16014 29774 16066 29783
rect 16174 29817 16226 29826
rect 16174 29783 16183 29817
rect 16183 29783 16217 29817
rect 16217 29783 16226 29817
rect 16174 29774 16226 29783
rect 16334 29817 16386 29826
rect 16334 29783 16343 29817
rect 16343 29783 16377 29817
rect 16377 29783 16386 29817
rect 16334 29774 16386 29783
rect 16494 29817 16546 29826
rect 16494 29783 16503 29817
rect 16503 29783 16537 29817
rect 16537 29783 16546 29817
rect 16494 29774 16546 29783
rect 16654 29817 16706 29826
rect 16654 29783 16663 29817
rect 16663 29783 16697 29817
rect 16697 29783 16706 29817
rect 16654 29774 16706 29783
rect 16814 29817 16866 29826
rect 16814 29783 16823 29817
rect 16823 29783 16857 29817
rect 16857 29783 16866 29817
rect 16814 29774 16866 29783
rect 16974 29817 17026 29826
rect 16974 29783 16983 29817
rect 16983 29783 17017 29817
rect 17017 29783 17026 29817
rect 16974 29774 17026 29783
rect 17134 29817 17186 29826
rect 17134 29783 17143 29817
rect 17143 29783 17177 29817
rect 17177 29783 17186 29817
rect 17134 29774 17186 29783
rect 17294 29817 17346 29826
rect 17294 29783 17303 29817
rect 17303 29783 17337 29817
rect 17337 29783 17346 29817
rect 17294 29774 17346 29783
rect 17454 29817 17506 29826
rect 17454 29783 17463 29817
rect 17463 29783 17497 29817
rect 17497 29783 17506 29817
rect 17454 29774 17506 29783
rect 17614 29817 17666 29826
rect 17614 29783 17623 29817
rect 17623 29783 17657 29817
rect 17657 29783 17666 29817
rect 17614 29774 17666 29783
rect 17774 29817 17826 29826
rect 17774 29783 17783 29817
rect 17783 29783 17817 29817
rect 17817 29783 17826 29817
rect 17774 29774 17826 29783
rect 17934 29817 17986 29826
rect 17934 29783 17943 29817
rect 17943 29783 17977 29817
rect 17977 29783 17986 29817
rect 17934 29774 17986 29783
rect 18094 29817 18146 29826
rect 18094 29783 18103 29817
rect 18103 29783 18137 29817
rect 18137 29783 18146 29817
rect 18094 29774 18146 29783
rect 18254 29817 18306 29826
rect 18254 29783 18263 29817
rect 18263 29783 18297 29817
rect 18297 29783 18306 29817
rect 18254 29774 18306 29783
rect 18414 29817 18466 29826
rect 18414 29783 18423 29817
rect 18423 29783 18457 29817
rect 18457 29783 18466 29817
rect 18414 29774 18466 29783
rect 18574 29817 18626 29826
rect 18574 29783 18583 29817
rect 18583 29783 18617 29817
rect 18617 29783 18626 29817
rect 18574 29774 18626 29783
rect 18734 29817 18786 29826
rect 18734 29783 18743 29817
rect 18743 29783 18777 29817
rect 18777 29783 18786 29817
rect 18734 29774 18786 29783
rect 18894 29817 18946 29826
rect 18894 29783 18903 29817
rect 18903 29783 18937 29817
rect 18937 29783 18946 29817
rect 18894 29774 18946 29783
rect 23134 29817 23186 29826
rect 23134 29783 23143 29817
rect 23143 29783 23177 29817
rect 23177 29783 23186 29817
rect 23134 29774 23186 29783
rect 23294 29817 23346 29826
rect 23294 29783 23303 29817
rect 23303 29783 23337 29817
rect 23337 29783 23346 29817
rect 23294 29774 23346 29783
rect 23454 29817 23506 29826
rect 23454 29783 23463 29817
rect 23463 29783 23497 29817
rect 23497 29783 23506 29817
rect 23454 29774 23506 29783
rect 23614 29817 23666 29826
rect 23614 29783 23623 29817
rect 23623 29783 23657 29817
rect 23657 29783 23666 29817
rect 23614 29774 23666 29783
rect 23774 29817 23826 29826
rect 23774 29783 23783 29817
rect 23783 29783 23817 29817
rect 23817 29783 23826 29817
rect 23774 29774 23826 29783
rect 23934 29817 23986 29826
rect 23934 29783 23943 29817
rect 23943 29783 23977 29817
rect 23977 29783 23986 29817
rect 23934 29774 23986 29783
rect 24094 29817 24146 29826
rect 24094 29783 24103 29817
rect 24103 29783 24137 29817
rect 24137 29783 24146 29817
rect 24094 29774 24146 29783
rect 24254 29817 24306 29826
rect 24254 29783 24263 29817
rect 24263 29783 24297 29817
rect 24297 29783 24306 29817
rect 24254 29774 24306 29783
rect 24414 29817 24466 29826
rect 24414 29783 24423 29817
rect 24423 29783 24457 29817
rect 24457 29783 24466 29817
rect 24414 29774 24466 29783
rect 24574 29817 24626 29826
rect 24574 29783 24583 29817
rect 24583 29783 24617 29817
rect 24617 29783 24626 29817
rect 24574 29774 24626 29783
rect 24734 29817 24786 29826
rect 24734 29783 24743 29817
rect 24743 29783 24777 29817
rect 24777 29783 24786 29817
rect 24734 29774 24786 29783
rect 24894 29817 24946 29826
rect 24894 29783 24903 29817
rect 24903 29783 24937 29817
rect 24937 29783 24946 29817
rect 24894 29774 24946 29783
rect 25054 29817 25106 29826
rect 25054 29783 25063 29817
rect 25063 29783 25097 29817
rect 25097 29783 25106 29817
rect 25054 29774 25106 29783
rect 25214 29817 25266 29826
rect 25214 29783 25223 29817
rect 25223 29783 25257 29817
rect 25257 29783 25266 29817
rect 25214 29774 25266 29783
rect 25374 29817 25426 29826
rect 25374 29783 25383 29817
rect 25383 29783 25417 29817
rect 25417 29783 25426 29817
rect 25374 29774 25426 29783
rect 25534 29817 25586 29826
rect 25534 29783 25543 29817
rect 25543 29783 25577 29817
rect 25577 29783 25586 29817
rect 25534 29774 25586 29783
rect 25694 29817 25746 29826
rect 25694 29783 25703 29817
rect 25703 29783 25737 29817
rect 25737 29783 25746 29817
rect 25694 29774 25746 29783
rect 25854 29817 25906 29826
rect 25854 29783 25863 29817
rect 25863 29783 25897 29817
rect 25897 29783 25906 29817
rect 25854 29774 25906 29783
rect 26014 29817 26066 29826
rect 26014 29783 26023 29817
rect 26023 29783 26057 29817
rect 26057 29783 26066 29817
rect 26014 29774 26066 29783
rect 26174 29817 26226 29826
rect 26174 29783 26183 29817
rect 26183 29783 26217 29817
rect 26217 29783 26226 29817
rect 26174 29774 26226 29783
rect 26334 29817 26386 29826
rect 26334 29783 26343 29817
rect 26343 29783 26377 29817
rect 26377 29783 26386 29817
rect 26334 29774 26386 29783
rect 26494 29817 26546 29826
rect 26494 29783 26503 29817
rect 26503 29783 26537 29817
rect 26537 29783 26546 29817
rect 26494 29774 26546 29783
rect 26654 29817 26706 29826
rect 26654 29783 26663 29817
rect 26663 29783 26697 29817
rect 26697 29783 26706 29817
rect 26654 29774 26706 29783
rect 26814 29817 26866 29826
rect 26814 29783 26823 29817
rect 26823 29783 26857 29817
rect 26857 29783 26866 29817
rect 26814 29774 26866 29783
rect 26974 29817 27026 29826
rect 26974 29783 26983 29817
rect 26983 29783 27017 29817
rect 27017 29783 27026 29817
rect 26974 29774 27026 29783
rect 27134 29817 27186 29826
rect 27134 29783 27143 29817
rect 27143 29783 27177 29817
rect 27177 29783 27186 29817
rect 27134 29774 27186 29783
rect 27294 29817 27346 29826
rect 27294 29783 27303 29817
rect 27303 29783 27337 29817
rect 27337 29783 27346 29817
rect 27294 29774 27346 29783
rect 27454 29817 27506 29826
rect 27454 29783 27463 29817
rect 27463 29783 27497 29817
rect 27497 29783 27506 29817
rect 27454 29774 27506 29783
rect 27614 29817 27666 29826
rect 27614 29783 27623 29817
rect 27623 29783 27657 29817
rect 27657 29783 27666 29817
rect 27614 29774 27666 29783
rect 27774 29817 27826 29826
rect 27774 29783 27783 29817
rect 27783 29783 27817 29817
rect 27817 29783 27826 29817
rect 27774 29774 27826 29783
rect 27934 29817 27986 29826
rect 27934 29783 27943 29817
rect 27943 29783 27977 29817
rect 27977 29783 27986 29817
rect 27934 29774 27986 29783
rect 28094 29817 28146 29826
rect 28094 29783 28103 29817
rect 28103 29783 28137 29817
rect 28137 29783 28146 29817
rect 28094 29774 28146 29783
rect 28254 29817 28306 29826
rect 28254 29783 28263 29817
rect 28263 29783 28297 29817
rect 28297 29783 28306 29817
rect 28254 29774 28306 29783
rect 28414 29817 28466 29826
rect 28414 29783 28423 29817
rect 28423 29783 28457 29817
rect 28457 29783 28466 29817
rect 28414 29774 28466 29783
rect 28574 29817 28626 29826
rect 28574 29783 28583 29817
rect 28583 29783 28617 29817
rect 28617 29783 28626 29817
rect 28574 29774 28626 29783
rect 28734 29817 28786 29826
rect 28734 29783 28743 29817
rect 28743 29783 28777 29817
rect 28777 29783 28786 29817
rect 28734 29774 28786 29783
rect 28894 29817 28946 29826
rect 28894 29783 28903 29817
rect 28903 29783 28937 29817
rect 28937 29783 28946 29817
rect 28894 29774 28946 29783
rect 29054 29817 29106 29826
rect 29054 29783 29063 29817
rect 29063 29783 29097 29817
rect 29097 29783 29106 29817
rect 29054 29774 29106 29783
rect 29214 29817 29266 29826
rect 29214 29783 29223 29817
rect 29223 29783 29257 29817
rect 29257 29783 29266 29817
rect 29214 29774 29266 29783
rect 29374 29817 29426 29826
rect 29374 29783 29383 29817
rect 29383 29783 29417 29817
rect 29417 29783 29426 29817
rect 29374 29774 29426 29783
rect 33534 29817 33586 29826
rect 33534 29783 33543 29817
rect 33543 29783 33577 29817
rect 33577 29783 33586 29817
rect 33534 29774 33586 29783
rect 33694 29817 33746 29826
rect 33694 29783 33703 29817
rect 33703 29783 33737 29817
rect 33737 29783 33746 29817
rect 33694 29774 33746 29783
rect 33854 29817 33906 29826
rect 33854 29783 33863 29817
rect 33863 29783 33897 29817
rect 33897 29783 33906 29817
rect 33854 29774 33906 29783
rect 34014 29817 34066 29826
rect 34014 29783 34023 29817
rect 34023 29783 34057 29817
rect 34057 29783 34066 29817
rect 34014 29774 34066 29783
rect 34174 29817 34226 29826
rect 34174 29783 34183 29817
rect 34183 29783 34217 29817
rect 34217 29783 34226 29817
rect 34174 29774 34226 29783
rect 34334 29817 34386 29826
rect 34334 29783 34343 29817
rect 34343 29783 34377 29817
rect 34377 29783 34386 29817
rect 34334 29774 34386 29783
rect 34494 29817 34546 29826
rect 34494 29783 34503 29817
rect 34503 29783 34537 29817
rect 34537 29783 34546 29817
rect 34494 29774 34546 29783
rect 34654 29817 34706 29826
rect 34654 29783 34663 29817
rect 34663 29783 34697 29817
rect 34697 29783 34706 29817
rect 34654 29774 34706 29783
rect 34814 29817 34866 29826
rect 34814 29783 34823 29817
rect 34823 29783 34857 29817
rect 34857 29783 34866 29817
rect 34814 29774 34866 29783
rect 34974 29817 35026 29826
rect 34974 29783 34983 29817
rect 34983 29783 35017 29817
rect 35017 29783 35026 29817
rect 34974 29774 35026 29783
rect 35134 29817 35186 29826
rect 35134 29783 35143 29817
rect 35143 29783 35177 29817
rect 35177 29783 35186 29817
rect 35134 29774 35186 29783
rect 35294 29817 35346 29826
rect 35294 29783 35303 29817
rect 35303 29783 35337 29817
rect 35337 29783 35346 29817
rect 35294 29774 35346 29783
rect 35454 29817 35506 29826
rect 35454 29783 35463 29817
rect 35463 29783 35497 29817
rect 35497 29783 35506 29817
rect 35454 29774 35506 29783
rect 35614 29817 35666 29826
rect 35614 29783 35623 29817
rect 35623 29783 35657 29817
rect 35657 29783 35666 29817
rect 35614 29774 35666 29783
rect 35774 29817 35826 29826
rect 35774 29783 35783 29817
rect 35783 29783 35817 29817
rect 35817 29783 35826 29817
rect 35774 29774 35826 29783
rect 35934 29817 35986 29826
rect 35934 29783 35943 29817
rect 35943 29783 35977 29817
rect 35977 29783 35986 29817
rect 35934 29774 35986 29783
rect 36094 29817 36146 29826
rect 36094 29783 36103 29817
rect 36103 29783 36137 29817
rect 36137 29783 36146 29817
rect 36094 29774 36146 29783
rect 36254 29817 36306 29826
rect 36254 29783 36263 29817
rect 36263 29783 36297 29817
rect 36297 29783 36306 29817
rect 36254 29774 36306 29783
rect 36414 29817 36466 29826
rect 36414 29783 36423 29817
rect 36423 29783 36457 29817
rect 36457 29783 36466 29817
rect 36414 29774 36466 29783
rect 36574 29817 36626 29826
rect 36574 29783 36583 29817
rect 36583 29783 36617 29817
rect 36617 29783 36626 29817
rect 36574 29774 36626 29783
rect 36734 29817 36786 29826
rect 36734 29783 36743 29817
rect 36743 29783 36777 29817
rect 36777 29783 36786 29817
rect 36734 29774 36786 29783
rect 36894 29817 36946 29826
rect 36894 29783 36903 29817
rect 36903 29783 36937 29817
rect 36937 29783 36946 29817
rect 36894 29774 36946 29783
rect 37054 29817 37106 29826
rect 37054 29783 37063 29817
rect 37063 29783 37097 29817
rect 37097 29783 37106 29817
rect 37054 29774 37106 29783
rect 37214 29817 37266 29826
rect 37214 29783 37223 29817
rect 37223 29783 37257 29817
rect 37257 29783 37266 29817
rect 37214 29774 37266 29783
rect 37374 29817 37426 29826
rect 37374 29783 37383 29817
rect 37383 29783 37417 29817
rect 37417 29783 37426 29817
rect 37374 29774 37426 29783
rect 37534 29817 37586 29826
rect 37534 29783 37543 29817
rect 37543 29783 37577 29817
rect 37577 29783 37586 29817
rect 37534 29774 37586 29783
rect 37694 29817 37746 29826
rect 37694 29783 37703 29817
rect 37703 29783 37737 29817
rect 37737 29783 37746 29817
rect 37694 29774 37746 29783
rect 37854 29817 37906 29826
rect 37854 29783 37863 29817
rect 37863 29783 37897 29817
rect 37897 29783 37906 29817
rect 37854 29774 37906 29783
rect 38014 29817 38066 29826
rect 38014 29783 38023 29817
rect 38023 29783 38057 29817
rect 38057 29783 38066 29817
rect 38014 29774 38066 29783
rect 38174 29817 38226 29826
rect 38174 29783 38183 29817
rect 38183 29783 38217 29817
rect 38217 29783 38226 29817
rect 38174 29774 38226 29783
rect 38334 29817 38386 29826
rect 38334 29783 38343 29817
rect 38343 29783 38377 29817
rect 38377 29783 38386 29817
rect 38334 29774 38386 29783
rect 38494 29817 38546 29826
rect 38494 29783 38503 29817
rect 38503 29783 38537 29817
rect 38537 29783 38546 29817
rect 38494 29774 38546 29783
rect 38654 29817 38706 29826
rect 38654 29783 38663 29817
rect 38663 29783 38697 29817
rect 38697 29783 38706 29817
rect 38654 29774 38706 29783
rect 38814 29817 38866 29826
rect 38814 29783 38823 29817
rect 38823 29783 38857 29817
rect 38857 29783 38866 29817
rect 38814 29774 38866 29783
rect 38974 29817 39026 29826
rect 38974 29783 38983 29817
rect 38983 29783 39017 29817
rect 39017 29783 39026 29817
rect 38974 29774 39026 29783
rect 39134 29817 39186 29826
rect 39134 29783 39143 29817
rect 39143 29783 39177 29817
rect 39177 29783 39186 29817
rect 39134 29774 39186 29783
rect 39294 29817 39346 29826
rect 39294 29783 39303 29817
rect 39303 29783 39337 29817
rect 39337 29783 39346 29817
rect 39294 29774 39346 29783
rect 39454 29817 39506 29826
rect 39454 29783 39463 29817
rect 39463 29783 39497 29817
rect 39497 29783 39506 29817
rect 39454 29774 39506 29783
rect 39614 29817 39666 29826
rect 39614 29783 39623 29817
rect 39623 29783 39657 29817
rect 39657 29783 39666 29817
rect 39614 29774 39666 29783
rect 39774 29817 39826 29826
rect 39774 29783 39783 29817
rect 39783 29783 39817 29817
rect 39817 29783 39826 29817
rect 39774 29774 39826 29783
rect 39934 29817 39986 29826
rect 39934 29783 39943 29817
rect 39943 29783 39977 29817
rect 39977 29783 39986 29817
rect 39934 29774 39986 29783
rect 40094 29817 40146 29826
rect 40094 29783 40103 29817
rect 40103 29783 40137 29817
rect 40137 29783 40146 29817
rect 40094 29774 40146 29783
rect 40254 29817 40306 29826
rect 40254 29783 40263 29817
rect 40263 29783 40297 29817
rect 40297 29783 40306 29817
rect 40254 29774 40306 29783
rect 40414 29817 40466 29826
rect 40414 29783 40423 29817
rect 40423 29783 40457 29817
rect 40457 29783 40466 29817
rect 40414 29774 40466 29783
rect 40574 29817 40626 29826
rect 40574 29783 40583 29817
rect 40583 29783 40617 29817
rect 40617 29783 40626 29817
rect 40574 29774 40626 29783
rect 40734 29817 40786 29826
rect 40734 29783 40743 29817
rect 40743 29783 40777 29817
rect 40777 29783 40786 29817
rect 40734 29774 40786 29783
rect 40894 29817 40946 29826
rect 40894 29783 40903 29817
rect 40903 29783 40937 29817
rect 40937 29783 40946 29817
rect 40894 29774 40946 29783
rect 41054 29817 41106 29826
rect 41054 29783 41063 29817
rect 41063 29783 41097 29817
rect 41097 29783 41106 29817
rect 41054 29774 41106 29783
rect 41214 29817 41266 29826
rect 41214 29783 41223 29817
rect 41223 29783 41257 29817
rect 41257 29783 41266 29817
rect 41214 29774 41266 29783
rect 41374 29817 41426 29826
rect 41374 29783 41383 29817
rect 41383 29783 41417 29817
rect 41417 29783 41426 29817
rect 41374 29774 41426 29783
rect 41534 29817 41586 29826
rect 41534 29783 41543 29817
rect 41543 29783 41577 29817
rect 41577 29783 41586 29817
rect 41534 29774 41586 29783
rect 41694 29817 41746 29826
rect 41694 29783 41703 29817
rect 41703 29783 41737 29817
rect 41737 29783 41746 29817
rect 41694 29774 41746 29783
rect 41854 29817 41906 29826
rect 41854 29783 41863 29817
rect 41863 29783 41897 29817
rect 41897 29783 41906 29817
rect 41854 29774 41906 29783
rect 14 29497 66 29506
rect 14 29463 23 29497
rect 23 29463 57 29497
rect 57 29463 66 29497
rect 14 29454 66 29463
rect 174 29497 226 29506
rect 174 29463 183 29497
rect 183 29463 217 29497
rect 217 29463 226 29497
rect 174 29454 226 29463
rect 334 29497 386 29506
rect 334 29463 343 29497
rect 343 29463 377 29497
rect 377 29463 386 29497
rect 334 29454 386 29463
rect 494 29497 546 29506
rect 494 29463 503 29497
rect 503 29463 537 29497
rect 537 29463 546 29497
rect 494 29454 546 29463
rect 654 29497 706 29506
rect 654 29463 663 29497
rect 663 29463 697 29497
rect 697 29463 706 29497
rect 654 29454 706 29463
rect 814 29497 866 29506
rect 814 29463 823 29497
rect 823 29463 857 29497
rect 857 29463 866 29497
rect 814 29454 866 29463
rect 974 29497 1026 29506
rect 974 29463 983 29497
rect 983 29463 1017 29497
rect 1017 29463 1026 29497
rect 974 29454 1026 29463
rect 1134 29497 1186 29506
rect 1134 29463 1143 29497
rect 1143 29463 1177 29497
rect 1177 29463 1186 29497
rect 1134 29454 1186 29463
rect 1294 29497 1346 29506
rect 1294 29463 1303 29497
rect 1303 29463 1337 29497
rect 1337 29463 1346 29497
rect 1294 29454 1346 29463
rect 1454 29497 1506 29506
rect 1454 29463 1463 29497
rect 1463 29463 1497 29497
rect 1497 29463 1506 29497
rect 1454 29454 1506 29463
rect 1614 29497 1666 29506
rect 1614 29463 1623 29497
rect 1623 29463 1657 29497
rect 1657 29463 1666 29497
rect 1614 29454 1666 29463
rect 1774 29497 1826 29506
rect 1774 29463 1783 29497
rect 1783 29463 1817 29497
rect 1817 29463 1826 29497
rect 1774 29454 1826 29463
rect 1934 29497 1986 29506
rect 1934 29463 1943 29497
rect 1943 29463 1977 29497
rect 1977 29463 1986 29497
rect 1934 29454 1986 29463
rect 2094 29497 2146 29506
rect 2094 29463 2103 29497
rect 2103 29463 2137 29497
rect 2137 29463 2146 29497
rect 2094 29454 2146 29463
rect 2254 29497 2306 29506
rect 2254 29463 2263 29497
rect 2263 29463 2297 29497
rect 2297 29463 2306 29497
rect 2254 29454 2306 29463
rect 2414 29497 2466 29506
rect 2414 29463 2423 29497
rect 2423 29463 2457 29497
rect 2457 29463 2466 29497
rect 2414 29454 2466 29463
rect 2574 29497 2626 29506
rect 2574 29463 2583 29497
rect 2583 29463 2617 29497
rect 2617 29463 2626 29497
rect 2574 29454 2626 29463
rect 2734 29497 2786 29506
rect 2734 29463 2743 29497
rect 2743 29463 2777 29497
rect 2777 29463 2786 29497
rect 2734 29454 2786 29463
rect 2894 29497 2946 29506
rect 2894 29463 2903 29497
rect 2903 29463 2937 29497
rect 2937 29463 2946 29497
rect 2894 29454 2946 29463
rect 3054 29497 3106 29506
rect 3054 29463 3063 29497
rect 3063 29463 3097 29497
rect 3097 29463 3106 29497
rect 3054 29454 3106 29463
rect 3214 29497 3266 29506
rect 3214 29463 3223 29497
rect 3223 29463 3257 29497
rect 3257 29463 3266 29497
rect 3214 29454 3266 29463
rect 3374 29497 3426 29506
rect 3374 29463 3383 29497
rect 3383 29463 3417 29497
rect 3417 29463 3426 29497
rect 3374 29454 3426 29463
rect 3534 29497 3586 29506
rect 3534 29463 3543 29497
rect 3543 29463 3577 29497
rect 3577 29463 3586 29497
rect 3534 29454 3586 29463
rect 3694 29497 3746 29506
rect 3694 29463 3703 29497
rect 3703 29463 3737 29497
rect 3737 29463 3746 29497
rect 3694 29454 3746 29463
rect 3854 29497 3906 29506
rect 3854 29463 3863 29497
rect 3863 29463 3897 29497
rect 3897 29463 3906 29497
rect 3854 29454 3906 29463
rect 4014 29497 4066 29506
rect 4014 29463 4023 29497
rect 4023 29463 4057 29497
rect 4057 29463 4066 29497
rect 4014 29454 4066 29463
rect 4174 29497 4226 29506
rect 4174 29463 4183 29497
rect 4183 29463 4217 29497
rect 4217 29463 4226 29497
rect 4174 29454 4226 29463
rect 4334 29497 4386 29506
rect 4334 29463 4343 29497
rect 4343 29463 4377 29497
rect 4377 29463 4386 29497
rect 4334 29454 4386 29463
rect 4494 29497 4546 29506
rect 4494 29463 4503 29497
rect 4503 29463 4537 29497
rect 4537 29463 4546 29497
rect 4494 29454 4546 29463
rect 4654 29497 4706 29506
rect 4654 29463 4663 29497
rect 4663 29463 4697 29497
rect 4697 29463 4706 29497
rect 4654 29454 4706 29463
rect 4814 29497 4866 29506
rect 4814 29463 4823 29497
rect 4823 29463 4857 29497
rect 4857 29463 4866 29497
rect 4814 29454 4866 29463
rect 4974 29497 5026 29506
rect 4974 29463 4983 29497
rect 4983 29463 5017 29497
rect 5017 29463 5026 29497
rect 4974 29454 5026 29463
rect 5134 29497 5186 29506
rect 5134 29463 5143 29497
rect 5143 29463 5177 29497
rect 5177 29463 5186 29497
rect 5134 29454 5186 29463
rect 5294 29497 5346 29506
rect 5294 29463 5303 29497
rect 5303 29463 5337 29497
rect 5337 29463 5346 29497
rect 5294 29454 5346 29463
rect 5454 29497 5506 29506
rect 5454 29463 5463 29497
rect 5463 29463 5497 29497
rect 5497 29463 5506 29497
rect 5454 29454 5506 29463
rect 5614 29497 5666 29506
rect 5614 29463 5623 29497
rect 5623 29463 5657 29497
rect 5657 29463 5666 29497
rect 5614 29454 5666 29463
rect 5774 29497 5826 29506
rect 5774 29463 5783 29497
rect 5783 29463 5817 29497
rect 5817 29463 5826 29497
rect 5774 29454 5826 29463
rect 5934 29497 5986 29506
rect 5934 29463 5943 29497
rect 5943 29463 5977 29497
rect 5977 29463 5986 29497
rect 5934 29454 5986 29463
rect 6094 29497 6146 29506
rect 6094 29463 6103 29497
rect 6103 29463 6137 29497
rect 6137 29463 6146 29497
rect 6094 29454 6146 29463
rect 6254 29497 6306 29506
rect 6254 29463 6263 29497
rect 6263 29463 6297 29497
rect 6297 29463 6306 29497
rect 6254 29454 6306 29463
rect 6414 29497 6466 29506
rect 6414 29463 6423 29497
rect 6423 29463 6457 29497
rect 6457 29463 6466 29497
rect 6414 29454 6466 29463
rect 6574 29497 6626 29506
rect 6574 29463 6583 29497
rect 6583 29463 6617 29497
rect 6617 29463 6626 29497
rect 6574 29454 6626 29463
rect 6734 29497 6786 29506
rect 6734 29463 6743 29497
rect 6743 29463 6777 29497
rect 6777 29463 6786 29497
rect 6734 29454 6786 29463
rect 6894 29497 6946 29506
rect 6894 29463 6903 29497
rect 6903 29463 6937 29497
rect 6937 29463 6946 29497
rect 6894 29454 6946 29463
rect 7054 29497 7106 29506
rect 7054 29463 7063 29497
rect 7063 29463 7097 29497
rect 7097 29463 7106 29497
rect 7054 29454 7106 29463
rect 7214 29497 7266 29506
rect 7214 29463 7223 29497
rect 7223 29463 7257 29497
rect 7257 29463 7266 29497
rect 7214 29454 7266 29463
rect 7374 29497 7426 29506
rect 7374 29463 7383 29497
rect 7383 29463 7417 29497
rect 7417 29463 7426 29497
rect 7374 29454 7426 29463
rect 7534 29497 7586 29506
rect 7534 29463 7543 29497
rect 7543 29463 7577 29497
rect 7577 29463 7586 29497
rect 7534 29454 7586 29463
rect 7694 29497 7746 29506
rect 7694 29463 7703 29497
rect 7703 29463 7737 29497
rect 7737 29463 7746 29497
rect 7694 29454 7746 29463
rect 7854 29497 7906 29506
rect 7854 29463 7863 29497
rect 7863 29463 7897 29497
rect 7897 29463 7906 29497
rect 7854 29454 7906 29463
rect 8014 29497 8066 29506
rect 8014 29463 8023 29497
rect 8023 29463 8057 29497
rect 8057 29463 8066 29497
rect 8014 29454 8066 29463
rect 8174 29497 8226 29506
rect 8174 29463 8183 29497
rect 8183 29463 8217 29497
rect 8217 29463 8226 29497
rect 8174 29454 8226 29463
rect 8334 29497 8386 29506
rect 8334 29463 8343 29497
rect 8343 29463 8377 29497
rect 8377 29463 8386 29497
rect 8334 29454 8386 29463
rect 12494 29497 12546 29506
rect 12494 29463 12503 29497
rect 12503 29463 12537 29497
rect 12537 29463 12546 29497
rect 12494 29454 12546 29463
rect 12654 29497 12706 29506
rect 12654 29463 12663 29497
rect 12663 29463 12697 29497
rect 12697 29463 12706 29497
rect 12654 29454 12706 29463
rect 12814 29497 12866 29506
rect 12814 29463 12823 29497
rect 12823 29463 12857 29497
rect 12857 29463 12866 29497
rect 12814 29454 12866 29463
rect 12974 29497 13026 29506
rect 12974 29463 12983 29497
rect 12983 29463 13017 29497
rect 13017 29463 13026 29497
rect 12974 29454 13026 29463
rect 13134 29497 13186 29506
rect 13134 29463 13143 29497
rect 13143 29463 13177 29497
rect 13177 29463 13186 29497
rect 13134 29454 13186 29463
rect 13294 29497 13346 29506
rect 13294 29463 13303 29497
rect 13303 29463 13337 29497
rect 13337 29463 13346 29497
rect 13294 29454 13346 29463
rect 13454 29497 13506 29506
rect 13454 29463 13463 29497
rect 13463 29463 13497 29497
rect 13497 29463 13506 29497
rect 13454 29454 13506 29463
rect 13614 29497 13666 29506
rect 13614 29463 13623 29497
rect 13623 29463 13657 29497
rect 13657 29463 13666 29497
rect 13614 29454 13666 29463
rect 13774 29497 13826 29506
rect 13774 29463 13783 29497
rect 13783 29463 13817 29497
rect 13817 29463 13826 29497
rect 13774 29454 13826 29463
rect 13934 29497 13986 29506
rect 13934 29463 13943 29497
rect 13943 29463 13977 29497
rect 13977 29463 13986 29497
rect 13934 29454 13986 29463
rect 14094 29497 14146 29506
rect 14094 29463 14103 29497
rect 14103 29463 14137 29497
rect 14137 29463 14146 29497
rect 14094 29454 14146 29463
rect 14254 29497 14306 29506
rect 14254 29463 14263 29497
rect 14263 29463 14297 29497
rect 14297 29463 14306 29497
rect 14254 29454 14306 29463
rect 14414 29497 14466 29506
rect 14414 29463 14423 29497
rect 14423 29463 14457 29497
rect 14457 29463 14466 29497
rect 14414 29454 14466 29463
rect 14574 29497 14626 29506
rect 14574 29463 14583 29497
rect 14583 29463 14617 29497
rect 14617 29463 14626 29497
rect 14574 29454 14626 29463
rect 14734 29497 14786 29506
rect 14734 29463 14743 29497
rect 14743 29463 14777 29497
rect 14777 29463 14786 29497
rect 14734 29454 14786 29463
rect 14894 29497 14946 29506
rect 14894 29463 14903 29497
rect 14903 29463 14937 29497
rect 14937 29463 14946 29497
rect 14894 29454 14946 29463
rect 15054 29497 15106 29506
rect 15054 29463 15063 29497
rect 15063 29463 15097 29497
rect 15097 29463 15106 29497
rect 15054 29454 15106 29463
rect 15214 29497 15266 29506
rect 15214 29463 15223 29497
rect 15223 29463 15257 29497
rect 15257 29463 15266 29497
rect 15214 29454 15266 29463
rect 15374 29497 15426 29506
rect 15374 29463 15383 29497
rect 15383 29463 15417 29497
rect 15417 29463 15426 29497
rect 15374 29454 15426 29463
rect 15534 29497 15586 29506
rect 15534 29463 15543 29497
rect 15543 29463 15577 29497
rect 15577 29463 15586 29497
rect 15534 29454 15586 29463
rect 15694 29497 15746 29506
rect 15694 29463 15703 29497
rect 15703 29463 15737 29497
rect 15737 29463 15746 29497
rect 15694 29454 15746 29463
rect 15854 29497 15906 29506
rect 15854 29463 15863 29497
rect 15863 29463 15897 29497
rect 15897 29463 15906 29497
rect 15854 29454 15906 29463
rect 16014 29497 16066 29506
rect 16014 29463 16023 29497
rect 16023 29463 16057 29497
rect 16057 29463 16066 29497
rect 16014 29454 16066 29463
rect 16174 29497 16226 29506
rect 16174 29463 16183 29497
rect 16183 29463 16217 29497
rect 16217 29463 16226 29497
rect 16174 29454 16226 29463
rect 16334 29497 16386 29506
rect 16334 29463 16343 29497
rect 16343 29463 16377 29497
rect 16377 29463 16386 29497
rect 16334 29454 16386 29463
rect 16494 29497 16546 29506
rect 16494 29463 16503 29497
rect 16503 29463 16537 29497
rect 16537 29463 16546 29497
rect 16494 29454 16546 29463
rect 16654 29497 16706 29506
rect 16654 29463 16663 29497
rect 16663 29463 16697 29497
rect 16697 29463 16706 29497
rect 16654 29454 16706 29463
rect 16814 29497 16866 29506
rect 16814 29463 16823 29497
rect 16823 29463 16857 29497
rect 16857 29463 16866 29497
rect 16814 29454 16866 29463
rect 16974 29497 17026 29506
rect 16974 29463 16983 29497
rect 16983 29463 17017 29497
rect 17017 29463 17026 29497
rect 16974 29454 17026 29463
rect 17134 29497 17186 29506
rect 17134 29463 17143 29497
rect 17143 29463 17177 29497
rect 17177 29463 17186 29497
rect 17134 29454 17186 29463
rect 17294 29497 17346 29506
rect 17294 29463 17303 29497
rect 17303 29463 17337 29497
rect 17337 29463 17346 29497
rect 17294 29454 17346 29463
rect 17454 29497 17506 29506
rect 17454 29463 17463 29497
rect 17463 29463 17497 29497
rect 17497 29463 17506 29497
rect 17454 29454 17506 29463
rect 17614 29497 17666 29506
rect 17614 29463 17623 29497
rect 17623 29463 17657 29497
rect 17657 29463 17666 29497
rect 17614 29454 17666 29463
rect 17774 29497 17826 29506
rect 17774 29463 17783 29497
rect 17783 29463 17817 29497
rect 17817 29463 17826 29497
rect 17774 29454 17826 29463
rect 17934 29497 17986 29506
rect 17934 29463 17943 29497
rect 17943 29463 17977 29497
rect 17977 29463 17986 29497
rect 17934 29454 17986 29463
rect 18094 29497 18146 29506
rect 18094 29463 18103 29497
rect 18103 29463 18137 29497
rect 18137 29463 18146 29497
rect 18094 29454 18146 29463
rect 18254 29497 18306 29506
rect 18254 29463 18263 29497
rect 18263 29463 18297 29497
rect 18297 29463 18306 29497
rect 18254 29454 18306 29463
rect 18414 29497 18466 29506
rect 18414 29463 18423 29497
rect 18423 29463 18457 29497
rect 18457 29463 18466 29497
rect 18414 29454 18466 29463
rect 18574 29497 18626 29506
rect 18574 29463 18583 29497
rect 18583 29463 18617 29497
rect 18617 29463 18626 29497
rect 18574 29454 18626 29463
rect 18734 29497 18786 29506
rect 18734 29463 18743 29497
rect 18743 29463 18777 29497
rect 18777 29463 18786 29497
rect 18734 29454 18786 29463
rect 18894 29497 18946 29506
rect 18894 29463 18903 29497
rect 18903 29463 18937 29497
rect 18937 29463 18946 29497
rect 18894 29454 18946 29463
rect 23134 29497 23186 29506
rect 23134 29463 23143 29497
rect 23143 29463 23177 29497
rect 23177 29463 23186 29497
rect 23134 29454 23186 29463
rect 23294 29497 23346 29506
rect 23294 29463 23303 29497
rect 23303 29463 23337 29497
rect 23337 29463 23346 29497
rect 23294 29454 23346 29463
rect 23454 29497 23506 29506
rect 23454 29463 23463 29497
rect 23463 29463 23497 29497
rect 23497 29463 23506 29497
rect 23454 29454 23506 29463
rect 23614 29497 23666 29506
rect 23614 29463 23623 29497
rect 23623 29463 23657 29497
rect 23657 29463 23666 29497
rect 23614 29454 23666 29463
rect 23774 29497 23826 29506
rect 23774 29463 23783 29497
rect 23783 29463 23817 29497
rect 23817 29463 23826 29497
rect 23774 29454 23826 29463
rect 23934 29497 23986 29506
rect 23934 29463 23943 29497
rect 23943 29463 23977 29497
rect 23977 29463 23986 29497
rect 23934 29454 23986 29463
rect 24094 29497 24146 29506
rect 24094 29463 24103 29497
rect 24103 29463 24137 29497
rect 24137 29463 24146 29497
rect 24094 29454 24146 29463
rect 24254 29497 24306 29506
rect 24254 29463 24263 29497
rect 24263 29463 24297 29497
rect 24297 29463 24306 29497
rect 24254 29454 24306 29463
rect 24414 29497 24466 29506
rect 24414 29463 24423 29497
rect 24423 29463 24457 29497
rect 24457 29463 24466 29497
rect 24414 29454 24466 29463
rect 24574 29497 24626 29506
rect 24574 29463 24583 29497
rect 24583 29463 24617 29497
rect 24617 29463 24626 29497
rect 24574 29454 24626 29463
rect 24734 29497 24786 29506
rect 24734 29463 24743 29497
rect 24743 29463 24777 29497
rect 24777 29463 24786 29497
rect 24734 29454 24786 29463
rect 24894 29497 24946 29506
rect 24894 29463 24903 29497
rect 24903 29463 24937 29497
rect 24937 29463 24946 29497
rect 24894 29454 24946 29463
rect 25054 29497 25106 29506
rect 25054 29463 25063 29497
rect 25063 29463 25097 29497
rect 25097 29463 25106 29497
rect 25054 29454 25106 29463
rect 25214 29497 25266 29506
rect 25214 29463 25223 29497
rect 25223 29463 25257 29497
rect 25257 29463 25266 29497
rect 25214 29454 25266 29463
rect 25374 29497 25426 29506
rect 25374 29463 25383 29497
rect 25383 29463 25417 29497
rect 25417 29463 25426 29497
rect 25374 29454 25426 29463
rect 25534 29497 25586 29506
rect 25534 29463 25543 29497
rect 25543 29463 25577 29497
rect 25577 29463 25586 29497
rect 25534 29454 25586 29463
rect 25694 29497 25746 29506
rect 25694 29463 25703 29497
rect 25703 29463 25737 29497
rect 25737 29463 25746 29497
rect 25694 29454 25746 29463
rect 25854 29497 25906 29506
rect 25854 29463 25863 29497
rect 25863 29463 25897 29497
rect 25897 29463 25906 29497
rect 25854 29454 25906 29463
rect 26014 29497 26066 29506
rect 26014 29463 26023 29497
rect 26023 29463 26057 29497
rect 26057 29463 26066 29497
rect 26014 29454 26066 29463
rect 26174 29497 26226 29506
rect 26174 29463 26183 29497
rect 26183 29463 26217 29497
rect 26217 29463 26226 29497
rect 26174 29454 26226 29463
rect 26334 29497 26386 29506
rect 26334 29463 26343 29497
rect 26343 29463 26377 29497
rect 26377 29463 26386 29497
rect 26334 29454 26386 29463
rect 26494 29497 26546 29506
rect 26494 29463 26503 29497
rect 26503 29463 26537 29497
rect 26537 29463 26546 29497
rect 26494 29454 26546 29463
rect 26654 29497 26706 29506
rect 26654 29463 26663 29497
rect 26663 29463 26697 29497
rect 26697 29463 26706 29497
rect 26654 29454 26706 29463
rect 26814 29497 26866 29506
rect 26814 29463 26823 29497
rect 26823 29463 26857 29497
rect 26857 29463 26866 29497
rect 26814 29454 26866 29463
rect 26974 29497 27026 29506
rect 26974 29463 26983 29497
rect 26983 29463 27017 29497
rect 27017 29463 27026 29497
rect 26974 29454 27026 29463
rect 27134 29497 27186 29506
rect 27134 29463 27143 29497
rect 27143 29463 27177 29497
rect 27177 29463 27186 29497
rect 27134 29454 27186 29463
rect 27294 29497 27346 29506
rect 27294 29463 27303 29497
rect 27303 29463 27337 29497
rect 27337 29463 27346 29497
rect 27294 29454 27346 29463
rect 27454 29497 27506 29506
rect 27454 29463 27463 29497
rect 27463 29463 27497 29497
rect 27497 29463 27506 29497
rect 27454 29454 27506 29463
rect 27614 29497 27666 29506
rect 27614 29463 27623 29497
rect 27623 29463 27657 29497
rect 27657 29463 27666 29497
rect 27614 29454 27666 29463
rect 27774 29497 27826 29506
rect 27774 29463 27783 29497
rect 27783 29463 27817 29497
rect 27817 29463 27826 29497
rect 27774 29454 27826 29463
rect 27934 29497 27986 29506
rect 27934 29463 27943 29497
rect 27943 29463 27977 29497
rect 27977 29463 27986 29497
rect 27934 29454 27986 29463
rect 28094 29497 28146 29506
rect 28094 29463 28103 29497
rect 28103 29463 28137 29497
rect 28137 29463 28146 29497
rect 28094 29454 28146 29463
rect 28254 29497 28306 29506
rect 28254 29463 28263 29497
rect 28263 29463 28297 29497
rect 28297 29463 28306 29497
rect 28254 29454 28306 29463
rect 28414 29497 28466 29506
rect 28414 29463 28423 29497
rect 28423 29463 28457 29497
rect 28457 29463 28466 29497
rect 28414 29454 28466 29463
rect 28574 29497 28626 29506
rect 28574 29463 28583 29497
rect 28583 29463 28617 29497
rect 28617 29463 28626 29497
rect 28574 29454 28626 29463
rect 28734 29497 28786 29506
rect 28734 29463 28743 29497
rect 28743 29463 28777 29497
rect 28777 29463 28786 29497
rect 28734 29454 28786 29463
rect 28894 29497 28946 29506
rect 28894 29463 28903 29497
rect 28903 29463 28937 29497
rect 28937 29463 28946 29497
rect 28894 29454 28946 29463
rect 29054 29497 29106 29506
rect 29054 29463 29063 29497
rect 29063 29463 29097 29497
rect 29097 29463 29106 29497
rect 29054 29454 29106 29463
rect 29214 29497 29266 29506
rect 29214 29463 29223 29497
rect 29223 29463 29257 29497
rect 29257 29463 29266 29497
rect 29214 29454 29266 29463
rect 29374 29497 29426 29506
rect 29374 29463 29383 29497
rect 29383 29463 29417 29497
rect 29417 29463 29426 29497
rect 29374 29454 29426 29463
rect 33534 29497 33586 29506
rect 33534 29463 33543 29497
rect 33543 29463 33577 29497
rect 33577 29463 33586 29497
rect 33534 29454 33586 29463
rect 33694 29497 33746 29506
rect 33694 29463 33703 29497
rect 33703 29463 33737 29497
rect 33737 29463 33746 29497
rect 33694 29454 33746 29463
rect 33854 29497 33906 29506
rect 33854 29463 33863 29497
rect 33863 29463 33897 29497
rect 33897 29463 33906 29497
rect 33854 29454 33906 29463
rect 34014 29497 34066 29506
rect 34014 29463 34023 29497
rect 34023 29463 34057 29497
rect 34057 29463 34066 29497
rect 34014 29454 34066 29463
rect 34174 29497 34226 29506
rect 34174 29463 34183 29497
rect 34183 29463 34217 29497
rect 34217 29463 34226 29497
rect 34174 29454 34226 29463
rect 34334 29497 34386 29506
rect 34334 29463 34343 29497
rect 34343 29463 34377 29497
rect 34377 29463 34386 29497
rect 34334 29454 34386 29463
rect 34494 29497 34546 29506
rect 34494 29463 34503 29497
rect 34503 29463 34537 29497
rect 34537 29463 34546 29497
rect 34494 29454 34546 29463
rect 34654 29497 34706 29506
rect 34654 29463 34663 29497
rect 34663 29463 34697 29497
rect 34697 29463 34706 29497
rect 34654 29454 34706 29463
rect 34814 29497 34866 29506
rect 34814 29463 34823 29497
rect 34823 29463 34857 29497
rect 34857 29463 34866 29497
rect 34814 29454 34866 29463
rect 34974 29497 35026 29506
rect 34974 29463 34983 29497
rect 34983 29463 35017 29497
rect 35017 29463 35026 29497
rect 34974 29454 35026 29463
rect 35134 29497 35186 29506
rect 35134 29463 35143 29497
rect 35143 29463 35177 29497
rect 35177 29463 35186 29497
rect 35134 29454 35186 29463
rect 35294 29497 35346 29506
rect 35294 29463 35303 29497
rect 35303 29463 35337 29497
rect 35337 29463 35346 29497
rect 35294 29454 35346 29463
rect 35454 29497 35506 29506
rect 35454 29463 35463 29497
rect 35463 29463 35497 29497
rect 35497 29463 35506 29497
rect 35454 29454 35506 29463
rect 35614 29497 35666 29506
rect 35614 29463 35623 29497
rect 35623 29463 35657 29497
rect 35657 29463 35666 29497
rect 35614 29454 35666 29463
rect 35774 29497 35826 29506
rect 35774 29463 35783 29497
rect 35783 29463 35817 29497
rect 35817 29463 35826 29497
rect 35774 29454 35826 29463
rect 35934 29497 35986 29506
rect 35934 29463 35943 29497
rect 35943 29463 35977 29497
rect 35977 29463 35986 29497
rect 35934 29454 35986 29463
rect 36094 29497 36146 29506
rect 36094 29463 36103 29497
rect 36103 29463 36137 29497
rect 36137 29463 36146 29497
rect 36094 29454 36146 29463
rect 36254 29497 36306 29506
rect 36254 29463 36263 29497
rect 36263 29463 36297 29497
rect 36297 29463 36306 29497
rect 36254 29454 36306 29463
rect 36414 29497 36466 29506
rect 36414 29463 36423 29497
rect 36423 29463 36457 29497
rect 36457 29463 36466 29497
rect 36414 29454 36466 29463
rect 36574 29497 36626 29506
rect 36574 29463 36583 29497
rect 36583 29463 36617 29497
rect 36617 29463 36626 29497
rect 36574 29454 36626 29463
rect 36734 29497 36786 29506
rect 36734 29463 36743 29497
rect 36743 29463 36777 29497
rect 36777 29463 36786 29497
rect 36734 29454 36786 29463
rect 36894 29497 36946 29506
rect 36894 29463 36903 29497
rect 36903 29463 36937 29497
rect 36937 29463 36946 29497
rect 36894 29454 36946 29463
rect 37054 29497 37106 29506
rect 37054 29463 37063 29497
rect 37063 29463 37097 29497
rect 37097 29463 37106 29497
rect 37054 29454 37106 29463
rect 37214 29497 37266 29506
rect 37214 29463 37223 29497
rect 37223 29463 37257 29497
rect 37257 29463 37266 29497
rect 37214 29454 37266 29463
rect 37374 29497 37426 29506
rect 37374 29463 37383 29497
rect 37383 29463 37417 29497
rect 37417 29463 37426 29497
rect 37374 29454 37426 29463
rect 37534 29497 37586 29506
rect 37534 29463 37543 29497
rect 37543 29463 37577 29497
rect 37577 29463 37586 29497
rect 37534 29454 37586 29463
rect 37694 29497 37746 29506
rect 37694 29463 37703 29497
rect 37703 29463 37737 29497
rect 37737 29463 37746 29497
rect 37694 29454 37746 29463
rect 37854 29497 37906 29506
rect 37854 29463 37863 29497
rect 37863 29463 37897 29497
rect 37897 29463 37906 29497
rect 37854 29454 37906 29463
rect 38014 29497 38066 29506
rect 38014 29463 38023 29497
rect 38023 29463 38057 29497
rect 38057 29463 38066 29497
rect 38014 29454 38066 29463
rect 38174 29497 38226 29506
rect 38174 29463 38183 29497
rect 38183 29463 38217 29497
rect 38217 29463 38226 29497
rect 38174 29454 38226 29463
rect 38334 29497 38386 29506
rect 38334 29463 38343 29497
rect 38343 29463 38377 29497
rect 38377 29463 38386 29497
rect 38334 29454 38386 29463
rect 38494 29497 38546 29506
rect 38494 29463 38503 29497
rect 38503 29463 38537 29497
rect 38537 29463 38546 29497
rect 38494 29454 38546 29463
rect 38654 29497 38706 29506
rect 38654 29463 38663 29497
rect 38663 29463 38697 29497
rect 38697 29463 38706 29497
rect 38654 29454 38706 29463
rect 38814 29497 38866 29506
rect 38814 29463 38823 29497
rect 38823 29463 38857 29497
rect 38857 29463 38866 29497
rect 38814 29454 38866 29463
rect 38974 29497 39026 29506
rect 38974 29463 38983 29497
rect 38983 29463 39017 29497
rect 39017 29463 39026 29497
rect 38974 29454 39026 29463
rect 39134 29497 39186 29506
rect 39134 29463 39143 29497
rect 39143 29463 39177 29497
rect 39177 29463 39186 29497
rect 39134 29454 39186 29463
rect 39294 29497 39346 29506
rect 39294 29463 39303 29497
rect 39303 29463 39337 29497
rect 39337 29463 39346 29497
rect 39294 29454 39346 29463
rect 39454 29497 39506 29506
rect 39454 29463 39463 29497
rect 39463 29463 39497 29497
rect 39497 29463 39506 29497
rect 39454 29454 39506 29463
rect 39614 29497 39666 29506
rect 39614 29463 39623 29497
rect 39623 29463 39657 29497
rect 39657 29463 39666 29497
rect 39614 29454 39666 29463
rect 39774 29497 39826 29506
rect 39774 29463 39783 29497
rect 39783 29463 39817 29497
rect 39817 29463 39826 29497
rect 39774 29454 39826 29463
rect 39934 29497 39986 29506
rect 39934 29463 39943 29497
rect 39943 29463 39977 29497
rect 39977 29463 39986 29497
rect 39934 29454 39986 29463
rect 40094 29497 40146 29506
rect 40094 29463 40103 29497
rect 40103 29463 40137 29497
rect 40137 29463 40146 29497
rect 40094 29454 40146 29463
rect 40254 29497 40306 29506
rect 40254 29463 40263 29497
rect 40263 29463 40297 29497
rect 40297 29463 40306 29497
rect 40254 29454 40306 29463
rect 40414 29497 40466 29506
rect 40414 29463 40423 29497
rect 40423 29463 40457 29497
rect 40457 29463 40466 29497
rect 40414 29454 40466 29463
rect 40574 29497 40626 29506
rect 40574 29463 40583 29497
rect 40583 29463 40617 29497
rect 40617 29463 40626 29497
rect 40574 29454 40626 29463
rect 40734 29497 40786 29506
rect 40734 29463 40743 29497
rect 40743 29463 40777 29497
rect 40777 29463 40786 29497
rect 40734 29454 40786 29463
rect 40894 29497 40946 29506
rect 40894 29463 40903 29497
rect 40903 29463 40937 29497
rect 40937 29463 40946 29497
rect 40894 29454 40946 29463
rect 41054 29497 41106 29506
rect 41054 29463 41063 29497
rect 41063 29463 41097 29497
rect 41097 29463 41106 29497
rect 41054 29454 41106 29463
rect 41214 29497 41266 29506
rect 41214 29463 41223 29497
rect 41223 29463 41257 29497
rect 41257 29463 41266 29497
rect 41214 29454 41266 29463
rect 41374 29497 41426 29506
rect 41374 29463 41383 29497
rect 41383 29463 41417 29497
rect 41417 29463 41426 29497
rect 41374 29454 41426 29463
rect 41534 29497 41586 29506
rect 41534 29463 41543 29497
rect 41543 29463 41577 29497
rect 41577 29463 41586 29497
rect 41534 29454 41586 29463
rect 41694 29497 41746 29506
rect 41694 29463 41703 29497
rect 41703 29463 41737 29497
rect 41737 29463 41746 29497
rect 41694 29454 41746 29463
rect 41854 29497 41906 29506
rect 41854 29463 41863 29497
rect 41863 29463 41897 29497
rect 41897 29463 41906 29497
rect 41854 29454 41906 29463
<< metal2 >>
rect 0 37348 41920 37360
rect 0 37292 12 37348
rect 68 37292 172 37348
rect 228 37292 332 37348
rect 388 37292 492 37348
rect 548 37292 652 37348
rect 708 37292 812 37348
rect 868 37292 972 37348
rect 1028 37292 1132 37348
rect 1188 37292 1292 37348
rect 1348 37292 1452 37348
rect 1508 37292 1612 37348
rect 1668 37292 1772 37348
rect 1828 37292 1932 37348
rect 1988 37292 2092 37348
rect 2148 37292 2252 37348
rect 2308 37292 2412 37348
rect 2468 37292 2572 37348
rect 2628 37292 2732 37348
rect 2788 37292 2892 37348
rect 2948 37292 3052 37348
rect 3108 37292 3212 37348
rect 3268 37292 3372 37348
rect 3428 37292 3532 37348
rect 3588 37292 3692 37348
rect 3748 37292 3852 37348
rect 3908 37292 4012 37348
rect 4068 37292 4172 37348
rect 4228 37292 4332 37348
rect 4388 37292 4492 37348
rect 4548 37292 4652 37348
rect 4708 37292 4812 37348
rect 4868 37292 4972 37348
rect 5028 37292 5132 37348
rect 5188 37292 5292 37348
rect 5348 37292 5452 37348
rect 5508 37292 5612 37348
rect 5668 37292 5772 37348
rect 5828 37292 5932 37348
rect 5988 37292 6092 37348
rect 6148 37292 6252 37348
rect 6308 37292 6412 37348
rect 6468 37292 6572 37348
rect 6628 37292 6732 37348
rect 6788 37292 6892 37348
rect 6948 37292 7052 37348
rect 7108 37292 7212 37348
rect 7268 37292 7372 37348
rect 7428 37292 7532 37348
rect 7588 37292 7692 37348
rect 7748 37292 7852 37348
rect 7908 37292 8012 37348
rect 8068 37292 8172 37348
rect 8228 37292 8332 37348
rect 8388 37292 8492 37348
rect 8548 37292 8812 37348
rect 8868 37292 12492 37348
rect 12548 37292 12652 37348
rect 12708 37292 12812 37348
rect 12868 37292 12972 37348
rect 13028 37292 13132 37348
rect 13188 37292 13292 37348
rect 13348 37292 13452 37348
rect 13508 37292 13612 37348
rect 13668 37292 13772 37348
rect 13828 37292 13932 37348
rect 13988 37292 14092 37348
rect 14148 37292 14252 37348
rect 14308 37292 14412 37348
rect 14468 37292 14572 37348
rect 14628 37292 14732 37348
rect 14788 37292 14892 37348
rect 14948 37292 15052 37348
rect 15108 37292 15212 37348
rect 15268 37292 15372 37348
rect 15428 37292 15532 37348
rect 15588 37292 15692 37348
rect 15748 37292 15852 37348
rect 15908 37292 16012 37348
rect 16068 37292 16172 37348
rect 16228 37292 16332 37348
rect 16388 37292 16492 37348
rect 16548 37292 16652 37348
rect 16708 37292 16812 37348
rect 16868 37292 16972 37348
rect 17028 37292 17132 37348
rect 17188 37292 17292 37348
rect 17348 37292 17452 37348
rect 17508 37292 17612 37348
rect 17668 37292 17772 37348
rect 17828 37292 17932 37348
rect 17988 37292 18092 37348
rect 18148 37292 18252 37348
rect 18308 37292 18412 37348
rect 18468 37292 18572 37348
rect 18628 37292 18732 37348
rect 18788 37292 18892 37348
rect 18948 37292 22572 37348
rect 22628 37292 22892 37348
rect 22948 37292 23132 37348
rect 23188 37292 23292 37348
rect 23348 37292 23452 37348
rect 23508 37292 23612 37348
rect 23668 37292 23772 37348
rect 23828 37292 23932 37348
rect 23988 37292 24092 37348
rect 24148 37292 24252 37348
rect 24308 37292 24412 37348
rect 24468 37292 24572 37348
rect 24628 37292 24732 37348
rect 24788 37292 24892 37348
rect 24948 37292 25052 37348
rect 25108 37292 25212 37348
rect 25268 37292 25372 37348
rect 25428 37292 25532 37348
rect 25588 37292 25692 37348
rect 25748 37292 25852 37348
rect 25908 37292 26012 37348
rect 26068 37292 26172 37348
rect 26228 37292 26332 37348
rect 26388 37292 26492 37348
rect 26548 37292 26652 37348
rect 26708 37292 26812 37348
rect 26868 37292 26972 37348
rect 27028 37292 27132 37348
rect 27188 37292 27292 37348
rect 27348 37292 27452 37348
rect 27508 37292 27612 37348
rect 27668 37292 27772 37348
rect 27828 37292 27932 37348
rect 27988 37292 28092 37348
rect 28148 37292 28252 37348
rect 28308 37292 28412 37348
rect 28468 37292 28572 37348
rect 28628 37292 28732 37348
rect 28788 37292 28892 37348
rect 28948 37292 29052 37348
rect 29108 37292 29212 37348
rect 29268 37292 29372 37348
rect 29428 37292 33052 37348
rect 33108 37292 33372 37348
rect 33428 37292 33532 37348
rect 33588 37292 33692 37348
rect 33748 37292 33852 37348
rect 33908 37292 34012 37348
rect 34068 37292 34172 37348
rect 34228 37292 34332 37348
rect 34388 37292 34492 37348
rect 34548 37292 34652 37348
rect 34708 37292 34812 37348
rect 34868 37292 34972 37348
rect 35028 37292 35132 37348
rect 35188 37292 35292 37348
rect 35348 37292 35452 37348
rect 35508 37292 35612 37348
rect 35668 37292 35772 37348
rect 35828 37292 35932 37348
rect 35988 37292 36092 37348
rect 36148 37292 36252 37348
rect 36308 37292 36412 37348
rect 36468 37292 36572 37348
rect 36628 37292 36732 37348
rect 36788 37292 36892 37348
rect 36948 37292 37052 37348
rect 37108 37292 37212 37348
rect 37268 37292 37372 37348
rect 37428 37292 37532 37348
rect 37588 37292 37692 37348
rect 37748 37292 37852 37348
rect 37908 37292 38012 37348
rect 38068 37292 38172 37348
rect 38228 37292 38332 37348
rect 38388 37292 38492 37348
rect 38548 37292 38652 37348
rect 38708 37292 38812 37348
rect 38868 37292 38972 37348
rect 39028 37292 39132 37348
rect 39188 37292 39292 37348
rect 39348 37292 39452 37348
rect 39508 37292 39612 37348
rect 39668 37292 39772 37348
rect 39828 37292 39932 37348
rect 39988 37292 40092 37348
rect 40148 37292 40252 37348
rect 40308 37292 40412 37348
rect 40468 37292 40572 37348
rect 40628 37292 40732 37348
rect 40788 37292 40892 37348
rect 40948 37292 41052 37348
rect 41108 37292 41212 37348
rect 41268 37292 41372 37348
rect 41428 37292 41532 37348
rect 41588 37292 41692 37348
rect 41748 37292 41852 37348
rect 41908 37292 41920 37348
rect 0 37280 41920 37292
rect 0 37188 41920 37200
rect 0 37132 8652 37188
rect 8708 37132 22732 37188
rect 22788 37132 33212 37188
rect 33268 37132 41920 37188
rect 0 37120 41920 37132
rect 0 37028 41920 37040
rect 0 36972 12 37028
rect 68 36972 172 37028
rect 228 36972 332 37028
rect 388 36972 492 37028
rect 548 36972 652 37028
rect 708 36972 812 37028
rect 868 36972 972 37028
rect 1028 36972 1132 37028
rect 1188 36972 1292 37028
rect 1348 36972 1452 37028
rect 1508 36972 1612 37028
rect 1668 36972 1772 37028
rect 1828 36972 1932 37028
rect 1988 36972 2092 37028
rect 2148 36972 2252 37028
rect 2308 36972 2412 37028
rect 2468 36972 2572 37028
rect 2628 36972 2732 37028
rect 2788 36972 2892 37028
rect 2948 36972 3052 37028
rect 3108 36972 3212 37028
rect 3268 36972 3372 37028
rect 3428 36972 3532 37028
rect 3588 36972 3692 37028
rect 3748 36972 3852 37028
rect 3908 36972 4012 37028
rect 4068 36972 4172 37028
rect 4228 36972 4332 37028
rect 4388 36972 4492 37028
rect 4548 36972 4652 37028
rect 4708 36972 4812 37028
rect 4868 36972 4972 37028
rect 5028 36972 5132 37028
rect 5188 36972 5292 37028
rect 5348 36972 5452 37028
rect 5508 36972 5612 37028
rect 5668 36972 5772 37028
rect 5828 36972 5932 37028
rect 5988 36972 6092 37028
rect 6148 36972 6252 37028
rect 6308 36972 6412 37028
rect 6468 36972 6572 37028
rect 6628 36972 6732 37028
rect 6788 36972 6892 37028
rect 6948 36972 7052 37028
rect 7108 36972 7212 37028
rect 7268 36972 7372 37028
rect 7428 36972 7532 37028
rect 7588 36972 7692 37028
rect 7748 36972 7852 37028
rect 7908 36972 8012 37028
rect 8068 36972 8172 37028
rect 8228 36972 8332 37028
rect 8388 36972 8492 37028
rect 8548 36972 8812 37028
rect 8868 36972 12492 37028
rect 12548 36972 12652 37028
rect 12708 36972 12812 37028
rect 12868 36972 12972 37028
rect 13028 36972 13132 37028
rect 13188 36972 13292 37028
rect 13348 36972 13452 37028
rect 13508 36972 13612 37028
rect 13668 36972 13772 37028
rect 13828 36972 13932 37028
rect 13988 36972 14092 37028
rect 14148 36972 14252 37028
rect 14308 36972 14412 37028
rect 14468 36972 14572 37028
rect 14628 36972 14732 37028
rect 14788 36972 14892 37028
rect 14948 36972 15052 37028
rect 15108 36972 15212 37028
rect 15268 36972 15372 37028
rect 15428 36972 15532 37028
rect 15588 36972 15692 37028
rect 15748 36972 15852 37028
rect 15908 36972 16012 37028
rect 16068 36972 16172 37028
rect 16228 36972 16332 37028
rect 16388 36972 16492 37028
rect 16548 36972 16652 37028
rect 16708 36972 16812 37028
rect 16868 36972 16972 37028
rect 17028 36972 17132 37028
rect 17188 36972 17292 37028
rect 17348 36972 17452 37028
rect 17508 36972 17612 37028
rect 17668 36972 17772 37028
rect 17828 36972 17932 37028
rect 17988 36972 18092 37028
rect 18148 36972 18252 37028
rect 18308 36972 18412 37028
rect 18468 36972 18572 37028
rect 18628 36972 18732 37028
rect 18788 36972 18892 37028
rect 18948 36972 22572 37028
rect 22628 36972 22892 37028
rect 22948 36972 23132 37028
rect 23188 36972 23292 37028
rect 23348 36972 23452 37028
rect 23508 36972 23612 37028
rect 23668 36972 23772 37028
rect 23828 36972 23932 37028
rect 23988 36972 24092 37028
rect 24148 36972 24252 37028
rect 24308 36972 24412 37028
rect 24468 36972 24572 37028
rect 24628 36972 24732 37028
rect 24788 36972 24892 37028
rect 24948 36972 25052 37028
rect 25108 36972 25212 37028
rect 25268 36972 25372 37028
rect 25428 36972 25532 37028
rect 25588 36972 25692 37028
rect 25748 36972 25852 37028
rect 25908 36972 26012 37028
rect 26068 36972 26172 37028
rect 26228 36972 26332 37028
rect 26388 36972 26492 37028
rect 26548 36972 26652 37028
rect 26708 36972 26812 37028
rect 26868 36972 26972 37028
rect 27028 36972 27132 37028
rect 27188 36972 27292 37028
rect 27348 36972 27452 37028
rect 27508 36972 27612 37028
rect 27668 36972 27772 37028
rect 27828 36972 27932 37028
rect 27988 36972 28092 37028
rect 28148 36972 28252 37028
rect 28308 36972 28412 37028
rect 28468 36972 28572 37028
rect 28628 36972 28732 37028
rect 28788 36972 28892 37028
rect 28948 36972 29052 37028
rect 29108 36972 29212 37028
rect 29268 36972 29372 37028
rect 29428 36972 33052 37028
rect 33108 36972 33372 37028
rect 33428 36972 33532 37028
rect 33588 36972 33692 37028
rect 33748 36972 33852 37028
rect 33908 36972 34012 37028
rect 34068 36972 34172 37028
rect 34228 36972 34332 37028
rect 34388 36972 34492 37028
rect 34548 36972 34652 37028
rect 34708 36972 34812 37028
rect 34868 36972 34972 37028
rect 35028 36972 35132 37028
rect 35188 36972 35292 37028
rect 35348 36972 35452 37028
rect 35508 36972 35612 37028
rect 35668 36972 35772 37028
rect 35828 36972 35932 37028
rect 35988 36972 36092 37028
rect 36148 36972 36252 37028
rect 36308 36972 36412 37028
rect 36468 36972 36572 37028
rect 36628 36972 36732 37028
rect 36788 36972 36892 37028
rect 36948 36972 37052 37028
rect 37108 36972 37212 37028
rect 37268 36972 37372 37028
rect 37428 36972 37532 37028
rect 37588 36972 37692 37028
rect 37748 36972 37852 37028
rect 37908 36972 38012 37028
rect 38068 36972 38172 37028
rect 38228 36972 38332 37028
rect 38388 36972 38492 37028
rect 38548 36972 38652 37028
rect 38708 36972 38812 37028
rect 38868 36972 38972 37028
rect 39028 36972 39132 37028
rect 39188 36972 39292 37028
rect 39348 36972 39452 37028
rect 39508 36972 39612 37028
rect 39668 36972 39772 37028
rect 39828 36972 39932 37028
rect 39988 36972 40092 37028
rect 40148 36972 40252 37028
rect 40308 36972 40412 37028
rect 40468 36972 40572 37028
rect 40628 36972 40732 37028
rect 40788 36972 40892 37028
rect 40948 36972 41052 37028
rect 41108 36972 41212 37028
rect 41268 36972 41372 37028
rect 41428 36972 41532 37028
rect 41588 36972 41692 37028
rect 41748 36972 41852 37028
rect 41908 36972 41920 37028
rect 0 36960 41920 36972
rect 0 36868 41920 36880
rect 0 36812 12 36868
rect 68 36812 172 36868
rect 228 36812 332 36868
rect 388 36812 492 36868
rect 548 36812 652 36868
rect 708 36812 812 36868
rect 868 36812 972 36868
rect 1028 36812 1132 36868
rect 1188 36812 1292 36868
rect 1348 36812 1452 36868
rect 1508 36812 1612 36868
rect 1668 36812 1772 36868
rect 1828 36812 1932 36868
rect 1988 36812 2092 36868
rect 2148 36812 2252 36868
rect 2308 36812 2412 36868
rect 2468 36812 2572 36868
rect 2628 36812 2732 36868
rect 2788 36812 2892 36868
rect 2948 36812 3052 36868
rect 3108 36812 3212 36868
rect 3268 36812 3372 36868
rect 3428 36812 3532 36868
rect 3588 36812 3692 36868
rect 3748 36812 3852 36868
rect 3908 36812 4012 36868
rect 4068 36812 4172 36868
rect 4228 36812 4332 36868
rect 4388 36812 4492 36868
rect 4548 36812 4652 36868
rect 4708 36812 4812 36868
rect 4868 36812 4972 36868
rect 5028 36812 5132 36868
rect 5188 36812 5292 36868
rect 5348 36812 5452 36868
rect 5508 36812 5612 36868
rect 5668 36812 5772 36868
rect 5828 36812 5932 36868
rect 5988 36812 6092 36868
rect 6148 36812 6252 36868
rect 6308 36812 6412 36868
rect 6468 36812 6572 36868
rect 6628 36812 6732 36868
rect 6788 36812 6892 36868
rect 6948 36812 7052 36868
rect 7108 36812 7212 36868
rect 7268 36812 7372 36868
rect 7428 36812 7532 36868
rect 7588 36812 7692 36868
rect 7748 36812 7852 36868
rect 7908 36812 8012 36868
rect 8068 36812 8172 36868
rect 8228 36812 8332 36868
rect 8388 36812 8972 36868
rect 9028 36812 9292 36868
rect 9348 36812 12492 36868
rect 12548 36812 12652 36868
rect 12708 36812 12812 36868
rect 12868 36812 12972 36868
rect 13028 36812 13132 36868
rect 13188 36812 13292 36868
rect 13348 36812 13452 36868
rect 13508 36812 13612 36868
rect 13668 36812 13772 36868
rect 13828 36812 13932 36868
rect 13988 36812 14092 36868
rect 14148 36812 14252 36868
rect 14308 36812 14412 36868
rect 14468 36812 14572 36868
rect 14628 36812 14732 36868
rect 14788 36812 14892 36868
rect 14948 36812 15052 36868
rect 15108 36812 15212 36868
rect 15268 36812 15372 36868
rect 15428 36812 15532 36868
rect 15588 36812 15692 36868
rect 15748 36812 15852 36868
rect 15908 36812 16012 36868
rect 16068 36812 16172 36868
rect 16228 36812 16332 36868
rect 16388 36812 16492 36868
rect 16548 36812 16652 36868
rect 16708 36812 16812 36868
rect 16868 36812 16972 36868
rect 17028 36812 17132 36868
rect 17188 36812 17292 36868
rect 17348 36812 17452 36868
rect 17508 36812 17612 36868
rect 17668 36812 17772 36868
rect 17828 36812 17932 36868
rect 17988 36812 18092 36868
rect 18148 36812 18252 36868
rect 18308 36812 18412 36868
rect 18468 36812 18572 36868
rect 18628 36812 18732 36868
rect 18788 36812 18892 36868
rect 18948 36812 22092 36868
rect 22148 36812 22412 36868
rect 22468 36812 23132 36868
rect 23188 36812 23292 36868
rect 23348 36812 23452 36868
rect 23508 36812 23612 36868
rect 23668 36812 23772 36868
rect 23828 36812 23932 36868
rect 23988 36812 24092 36868
rect 24148 36812 24252 36868
rect 24308 36812 24412 36868
rect 24468 36812 24572 36868
rect 24628 36812 24732 36868
rect 24788 36812 24892 36868
rect 24948 36812 25052 36868
rect 25108 36812 25212 36868
rect 25268 36812 25372 36868
rect 25428 36812 25532 36868
rect 25588 36812 25692 36868
rect 25748 36812 25852 36868
rect 25908 36812 26012 36868
rect 26068 36812 26172 36868
rect 26228 36812 26332 36868
rect 26388 36812 26492 36868
rect 26548 36812 26652 36868
rect 26708 36812 26812 36868
rect 26868 36812 26972 36868
rect 27028 36812 27132 36868
rect 27188 36812 27292 36868
rect 27348 36812 27452 36868
rect 27508 36812 27612 36868
rect 27668 36812 27772 36868
rect 27828 36812 27932 36868
rect 27988 36812 28092 36868
rect 28148 36812 28252 36868
rect 28308 36812 28412 36868
rect 28468 36812 28572 36868
rect 28628 36812 28732 36868
rect 28788 36812 28892 36868
rect 28948 36812 29052 36868
rect 29108 36812 29212 36868
rect 29268 36812 29372 36868
rect 29428 36812 32572 36868
rect 32628 36812 32892 36868
rect 32948 36812 33532 36868
rect 33588 36812 33692 36868
rect 33748 36812 33852 36868
rect 33908 36812 34012 36868
rect 34068 36812 34172 36868
rect 34228 36812 34332 36868
rect 34388 36812 34492 36868
rect 34548 36812 34652 36868
rect 34708 36812 34812 36868
rect 34868 36812 34972 36868
rect 35028 36812 35132 36868
rect 35188 36812 35292 36868
rect 35348 36812 35452 36868
rect 35508 36812 35612 36868
rect 35668 36812 35772 36868
rect 35828 36812 35932 36868
rect 35988 36812 36092 36868
rect 36148 36812 36252 36868
rect 36308 36812 36412 36868
rect 36468 36812 36572 36868
rect 36628 36812 36732 36868
rect 36788 36812 36892 36868
rect 36948 36812 37052 36868
rect 37108 36812 37212 36868
rect 37268 36812 37372 36868
rect 37428 36812 37532 36868
rect 37588 36812 37692 36868
rect 37748 36812 37852 36868
rect 37908 36812 38012 36868
rect 38068 36812 38172 36868
rect 38228 36812 38332 36868
rect 38388 36812 38492 36868
rect 38548 36812 38652 36868
rect 38708 36812 38812 36868
rect 38868 36812 38972 36868
rect 39028 36812 39132 36868
rect 39188 36812 39292 36868
rect 39348 36812 39452 36868
rect 39508 36812 39612 36868
rect 39668 36812 39772 36868
rect 39828 36812 39932 36868
rect 39988 36812 40092 36868
rect 40148 36812 40252 36868
rect 40308 36812 40412 36868
rect 40468 36812 40572 36868
rect 40628 36812 40732 36868
rect 40788 36812 40892 36868
rect 40948 36812 41052 36868
rect 41108 36812 41212 36868
rect 41268 36812 41372 36868
rect 41428 36812 41532 36868
rect 41588 36812 41692 36868
rect 41748 36812 41852 36868
rect 41908 36812 41920 36868
rect 0 36800 41920 36812
rect 0 36708 41920 36720
rect 0 36652 9132 36708
rect 9188 36652 22252 36708
rect 22308 36652 32732 36708
rect 32788 36652 41920 36708
rect 0 36640 41920 36652
rect 0 36548 41920 36560
rect 0 36492 12 36548
rect 68 36492 172 36548
rect 228 36492 332 36548
rect 388 36492 492 36548
rect 548 36492 652 36548
rect 708 36492 812 36548
rect 868 36492 972 36548
rect 1028 36492 1132 36548
rect 1188 36492 1292 36548
rect 1348 36492 1452 36548
rect 1508 36492 1612 36548
rect 1668 36492 1772 36548
rect 1828 36492 1932 36548
rect 1988 36492 2092 36548
rect 2148 36492 2252 36548
rect 2308 36492 2412 36548
rect 2468 36492 2572 36548
rect 2628 36492 2732 36548
rect 2788 36492 2892 36548
rect 2948 36492 3052 36548
rect 3108 36492 3212 36548
rect 3268 36492 3372 36548
rect 3428 36492 3532 36548
rect 3588 36492 3692 36548
rect 3748 36492 3852 36548
rect 3908 36492 4012 36548
rect 4068 36492 4172 36548
rect 4228 36492 4332 36548
rect 4388 36492 4492 36548
rect 4548 36492 4652 36548
rect 4708 36492 4812 36548
rect 4868 36492 4972 36548
rect 5028 36492 5132 36548
rect 5188 36492 5292 36548
rect 5348 36492 5452 36548
rect 5508 36492 5612 36548
rect 5668 36492 5772 36548
rect 5828 36492 5932 36548
rect 5988 36492 6092 36548
rect 6148 36492 6252 36548
rect 6308 36492 6412 36548
rect 6468 36492 6572 36548
rect 6628 36492 6732 36548
rect 6788 36492 6892 36548
rect 6948 36492 7052 36548
rect 7108 36492 7212 36548
rect 7268 36492 7372 36548
rect 7428 36492 7532 36548
rect 7588 36492 7692 36548
rect 7748 36492 7852 36548
rect 7908 36492 8012 36548
rect 8068 36492 8172 36548
rect 8228 36492 8332 36548
rect 8388 36492 8972 36548
rect 9028 36492 9292 36548
rect 9348 36492 12492 36548
rect 12548 36492 12652 36548
rect 12708 36492 12812 36548
rect 12868 36492 12972 36548
rect 13028 36492 13132 36548
rect 13188 36492 13292 36548
rect 13348 36492 13452 36548
rect 13508 36492 13612 36548
rect 13668 36492 13772 36548
rect 13828 36492 13932 36548
rect 13988 36492 14092 36548
rect 14148 36492 14252 36548
rect 14308 36492 14412 36548
rect 14468 36492 14572 36548
rect 14628 36492 14732 36548
rect 14788 36492 14892 36548
rect 14948 36492 15052 36548
rect 15108 36492 15212 36548
rect 15268 36492 15372 36548
rect 15428 36492 15532 36548
rect 15588 36492 15692 36548
rect 15748 36492 15852 36548
rect 15908 36492 16012 36548
rect 16068 36492 16172 36548
rect 16228 36492 16332 36548
rect 16388 36492 16492 36548
rect 16548 36492 16652 36548
rect 16708 36492 16812 36548
rect 16868 36492 16972 36548
rect 17028 36492 17132 36548
rect 17188 36492 17292 36548
rect 17348 36492 17452 36548
rect 17508 36492 17612 36548
rect 17668 36492 17772 36548
rect 17828 36492 17932 36548
rect 17988 36492 18092 36548
rect 18148 36492 18252 36548
rect 18308 36492 18412 36548
rect 18468 36492 18572 36548
rect 18628 36492 18732 36548
rect 18788 36492 18892 36548
rect 18948 36492 22092 36548
rect 22148 36492 22412 36548
rect 22468 36492 23132 36548
rect 23188 36492 23292 36548
rect 23348 36492 23452 36548
rect 23508 36492 23612 36548
rect 23668 36492 23772 36548
rect 23828 36492 23932 36548
rect 23988 36492 24092 36548
rect 24148 36492 24252 36548
rect 24308 36492 24412 36548
rect 24468 36492 24572 36548
rect 24628 36492 24732 36548
rect 24788 36492 24892 36548
rect 24948 36492 25052 36548
rect 25108 36492 25212 36548
rect 25268 36492 25372 36548
rect 25428 36492 25532 36548
rect 25588 36492 25692 36548
rect 25748 36492 25852 36548
rect 25908 36492 26012 36548
rect 26068 36492 26172 36548
rect 26228 36492 26332 36548
rect 26388 36492 26492 36548
rect 26548 36492 26652 36548
rect 26708 36492 26812 36548
rect 26868 36492 26972 36548
rect 27028 36492 27132 36548
rect 27188 36492 27292 36548
rect 27348 36492 27452 36548
rect 27508 36492 27612 36548
rect 27668 36492 27772 36548
rect 27828 36492 27932 36548
rect 27988 36492 28092 36548
rect 28148 36492 28252 36548
rect 28308 36492 28412 36548
rect 28468 36492 28572 36548
rect 28628 36492 28732 36548
rect 28788 36492 28892 36548
rect 28948 36492 29052 36548
rect 29108 36492 29212 36548
rect 29268 36492 29372 36548
rect 29428 36492 32572 36548
rect 32628 36492 32892 36548
rect 32948 36492 33532 36548
rect 33588 36492 33692 36548
rect 33748 36492 33852 36548
rect 33908 36492 34012 36548
rect 34068 36492 34172 36548
rect 34228 36492 34332 36548
rect 34388 36492 34492 36548
rect 34548 36492 34652 36548
rect 34708 36492 34812 36548
rect 34868 36492 34972 36548
rect 35028 36492 35132 36548
rect 35188 36492 35292 36548
rect 35348 36492 35452 36548
rect 35508 36492 35612 36548
rect 35668 36492 35772 36548
rect 35828 36492 35932 36548
rect 35988 36492 36092 36548
rect 36148 36492 36252 36548
rect 36308 36492 36412 36548
rect 36468 36492 36572 36548
rect 36628 36492 36732 36548
rect 36788 36492 36892 36548
rect 36948 36492 37052 36548
rect 37108 36492 37212 36548
rect 37268 36492 37372 36548
rect 37428 36492 37532 36548
rect 37588 36492 37692 36548
rect 37748 36492 37852 36548
rect 37908 36492 38012 36548
rect 38068 36492 38172 36548
rect 38228 36492 38332 36548
rect 38388 36492 38492 36548
rect 38548 36492 38652 36548
rect 38708 36492 38812 36548
rect 38868 36492 38972 36548
rect 39028 36492 39132 36548
rect 39188 36492 39292 36548
rect 39348 36492 39452 36548
rect 39508 36492 39612 36548
rect 39668 36492 39772 36548
rect 39828 36492 39932 36548
rect 39988 36492 40092 36548
rect 40148 36492 40252 36548
rect 40308 36492 40412 36548
rect 40468 36492 40572 36548
rect 40628 36492 40732 36548
rect 40788 36492 40892 36548
rect 40948 36492 41052 36548
rect 41108 36492 41212 36548
rect 41268 36492 41372 36548
rect 41428 36492 41532 36548
rect 41588 36492 41692 36548
rect 41748 36492 41852 36548
rect 41908 36492 41920 36548
rect 0 36480 41920 36492
rect 0 36388 41920 36400
rect 0 36332 12 36388
rect 68 36332 172 36388
rect 228 36332 332 36388
rect 388 36332 492 36388
rect 548 36332 652 36388
rect 708 36332 812 36388
rect 868 36332 972 36388
rect 1028 36332 1132 36388
rect 1188 36332 1292 36388
rect 1348 36332 1452 36388
rect 1508 36332 1612 36388
rect 1668 36332 1772 36388
rect 1828 36332 1932 36388
rect 1988 36332 2092 36388
rect 2148 36332 2252 36388
rect 2308 36332 2412 36388
rect 2468 36332 2572 36388
rect 2628 36332 2732 36388
rect 2788 36332 2892 36388
rect 2948 36332 3052 36388
rect 3108 36332 3212 36388
rect 3268 36332 3372 36388
rect 3428 36332 3532 36388
rect 3588 36332 3692 36388
rect 3748 36332 3852 36388
rect 3908 36332 4012 36388
rect 4068 36332 4172 36388
rect 4228 36332 4332 36388
rect 4388 36332 4492 36388
rect 4548 36332 4652 36388
rect 4708 36332 4812 36388
rect 4868 36332 4972 36388
rect 5028 36332 5132 36388
rect 5188 36332 5292 36388
rect 5348 36332 5452 36388
rect 5508 36332 5612 36388
rect 5668 36332 5772 36388
rect 5828 36332 5932 36388
rect 5988 36332 6092 36388
rect 6148 36332 6252 36388
rect 6308 36332 6412 36388
rect 6468 36332 6572 36388
rect 6628 36332 6732 36388
rect 6788 36332 6892 36388
rect 6948 36332 7052 36388
rect 7108 36332 7212 36388
rect 7268 36332 7372 36388
rect 7428 36332 7532 36388
rect 7588 36332 7692 36388
rect 7748 36332 7852 36388
rect 7908 36332 8012 36388
rect 8068 36332 8172 36388
rect 8228 36332 8332 36388
rect 8388 36332 9452 36388
rect 9508 36332 9772 36388
rect 9828 36332 10092 36388
rect 10148 36332 10412 36388
rect 10468 36332 10732 36388
rect 10788 36332 11052 36388
rect 11108 36332 11372 36388
rect 11428 36332 12492 36388
rect 12548 36332 12652 36388
rect 12708 36332 12812 36388
rect 12868 36332 12972 36388
rect 13028 36332 13132 36388
rect 13188 36332 13292 36388
rect 13348 36332 13452 36388
rect 13508 36332 13612 36388
rect 13668 36332 13772 36388
rect 13828 36332 13932 36388
rect 13988 36332 14092 36388
rect 14148 36332 14252 36388
rect 14308 36332 14412 36388
rect 14468 36332 14572 36388
rect 14628 36332 14732 36388
rect 14788 36332 14892 36388
rect 14948 36332 15052 36388
rect 15108 36332 15212 36388
rect 15268 36332 15372 36388
rect 15428 36332 15532 36388
rect 15588 36332 15692 36388
rect 15748 36332 15852 36388
rect 15908 36332 16012 36388
rect 16068 36332 16172 36388
rect 16228 36332 16332 36388
rect 16388 36332 16492 36388
rect 16548 36332 16652 36388
rect 16708 36332 16812 36388
rect 16868 36332 16972 36388
rect 17028 36332 17132 36388
rect 17188 36332 17292 36388
rect 17348 36332 17452 36388
rect 17508 36332 17612 36388
rect 17668 36332 17772 36388
rect 17828 36332 17932 36388
rect 17988 36332 18092 36388
rect 18148 36332 18252 36388
rect 18308 36332 18412 36388
rect 18468 36332 18572 36388
rect 18628 36332 18732 36388
rect 18788 36332 18892 36388
rect 18948 36332 20012 36388
rect 20068 36332 20332 36388
rect 20388 36332 20652 36388
rect 20708 36332 20972 36388
rect 21028 36332 21292 36388
rect 21348 36332 21612 36388
rect 21668 36332 21932 36388
rect 21988 36332 23132 36388
rect 23188 36332 23292 36388
rect 23348 36332 23452 36388
rect 23508 36332 23612 36388
rect 23668 36332 23772 36388
rect 23828 36332 23932 36388
rect 23988 36332 24092 36388
rect 24148 36332 24252 36388
rect 24308 36332 24412 36388
rect 24468 36332 24572 36388
rect 24628 36332 24732 36388
rect 24788 36332 24892 36388
rect 24948 36332 25052 36388
rect 25108 36332 25212 36388
rect 25268 36332 25372 36388
rect 25428 36332 25532 36388
rect 25588 36332 25692 36388
rect 25748 36332 25852 36388
rect 25908 36332 26012 36388
rect 26068 36332 26172 36388
rect 26228 36332 26332 36388
rect 26388 36332 26492 36388
rect 26548 36332 26652 36388
rect 26708 36332 26812 36388
rect 26868 36332 26972 36388
rect 27028 36332 27132 36388
rect 27188 36332 27292 36388
rect 27348 36332 27452 36388
rect 27508 36332 27612 36388
rect 27668 36332 27772 36388
rect 27828 36332 27932 36388
rect 27988 36332 28092 36388
rect 28148 36332 28252 36388
rect 28308 36332 28412 36388
rect 28468 36332 28572 36388
rect 28628 36332 28732 36388
rect 28788 36332 28892 36388
rect 28948 36332 29052 36388
rect 29108 36332 29212 36388
rect 29268 36332 29372 36388
rect 29428 36332 30492 36388
rect 30548 36332 30812 36388
rect 30868 36332 31132 36388
rect 31188 36332 31452 36388
rect 31508 36332 31772 36388
rect 31828 36332 32092 36388
rect 32148 36332 32412 36388
rect 32468 36332 33532 36388
rect 33588 36332 33692 36388
rect 33748 36332 33852 36388
rect 33908 36332 34012 36388
rect 34068 36332 34172 36388
rect 34228 36332 34332 36388
rect 34388 36332 34492 36388
rect 34548 36332 34652 36388
rect 34708 36332 34812 36388
rect 34868 36332 34972 36388
rect 35028 36332 35132 36388
rect 35188 36332 35292 36388
rect 35348 36332 35452 36388
rect 35508 36332 35612 36388
rect 35668 36332 35772 36388
rect 35828 36332 35932 36388
rect 35988 36332 36092 36388
rect 36148 36332 36252 36388
rect 36308 36332 36412 36388
rect 36468 36332 36572 36388
rect 36628 36332 36732 36388
rect 36788 36332 36892 36388
rect 36948 36332 37052 36388
rect 37108 36332 37212 36388
rect 37268 36332 37372 36388
rect 37428 36332 37532 36388
rect 37588 36332 37692 36388
rect 37748 36332 37852 36388
rect 37908 36332 38012 36388
rect 38068 36332 38172 36388
rect 38228 36332 38332 36388
rect 38388 36332 38492 36388
rect 38548 36332 38652 36388
rect 38708 36332 38812 36388
rect 38868 36332 38972 36388
rect 39028 36332 39132 36388
rect 39188 36332 39292 36388
rect 39348 36332 39452 36388
rect 39508 36332 39612 36388
rect 39668 36332 39772 36388
rect 39828 36332 39932 36388
rect 39988 36332 40092 36388
rect 40148 36332 40252 36388
rect 40308 36332 40412 36388
rect 40468 36332 40572 36388
rect 40628 36332 40732 36388
rect 40788 36332 40892 36388
rect 40948 36332 41052 36388
rect 41108 36332 41212 36388
rect 41268 36332 41372 36388
rect 41428 36332 41532 36388
rect 41588 36332 41692 36388
rect 41748 36332 41852 36388
rect 41908 36332 41920 36388
rect 0 36320 41920 36332
rect 0 36228 41920 36240
rect 0 36172 9612 36228
rect 9668 36172 21772 36228
rect 21828 36172 32252 36228
rect 32308 36172 41920 36228
rect 0 36160 41920 36172
rect 0 36068 41920 36080
rect 0 36012 12 36068
rect 68 36012 172 36068
rect 228 36012 332 36068
rect 388 36012 492 36068
rect 548 36012 652 36068
rect 708 36012 812 36068
rect 868 36012 972 36068
rect 1028 36012 1132 36068
rect 1188 36012 1292 36068
rect 1348 36012 1452 36068
rect 1508 36012 1612 36068
rect 1668 36012 1772 36068
rect 1828 36012 1932 36068
rect 1988 36012 2092 36068
rect 2148 36012 2252 36068
rect 2308 36012 2412 36068
rect 2468 36012 2572 36068
rect 2628 36012 2732 36068
rect 2788 36012 2892 36068
rect 2948 36012 3052 36068
rect 3108 36012 3212 36068
rect 3268 36012 3372 36068
rect 3428 36012 3532 36068
rect 3588 36012 3692 36068
rect 3748 36012 3852 36068
rect 3908 36012 4012 36068
rect 4068 36012 4172 36068
rect 4228 36012 4332 36068
rect 4388 36012 4492 36068
rect 4548 36012 4652 36068
rect 4708 36012 4812 36068
rect 4868 36012 4972 36068
rect 5028 36012 5132 36068
rect 5188 36012 5292 36068
rect 5348 36012 5452 36068
rect 5508 36012 5612 36068
rect 5668 36012 5772 36068
rect 5828 36012 5932 36068
rect 5988 36012 6092 36068
rect 6148 36012 6252 36068
rect 6308 36012 6412 36068
rect 6468 36012 6572 36068
rect 6628 36012 6732 36068
rect 6788 36012 6892 36068
rect 6948 36012 7052 36068
rect 7108 36012 7212 36068
rect 7268 36012 7372 36068
rect 7428 36012 7532 36068
rect 7588 36012 7692 36068
rect 7748 36012 7852 36068
rect 7908 36012 8012 36068
rect 8068 36012 8172 36068
rect 8228 36012 8332 36068
rect 8388 36012 9452 36068
rect 9508 36012 9772 36068
rect 9828 36012 10092 36068
rect 10148 36012 10412 36068
rect 10468 36012 10732 36068
rect 10788 36012 11052 36068
rect 11108 36012 11372 36068
rect 11428 36012 12492 36068
rect 12548 36012 12652 36068
rect 12708 36012 12812 36068
rect 12868 36012 12972 36068
rect 13028 36012 13132 36068
rect 13188 36012 13292 36068
rect 13348 36012 13452 36068
rect 13508 36012 13612 36068
rect 13668 36012 13772 36068
rect 13828 36012 13932 36068
rect 13988 36012 14092 36068
rect 14148 36012 14252 36068
rect 14308 36012 14412 36068
rect 14468 36012 14572 36068
rect 14628 36012 14732 36068
rect 14788 36012 14892 36068
rect 14948 36012 15052 36068
rect 15108 36012 15212 36068
rect 15268 36012 15372 36068
rect 15428 36012 15532 36068
rect 15588 36012 15692 36068
rect 15748 36012 15852 36068
rect 15908 36012 16012 36068
rect 16068 36012 16172 36068
rect 16228 36012 16332 36068
rect 16388 36012 16492 36068
rect 16548 36012 16652 36068
rect 16708 36012 16812 36068
rect 16868 36012 16972 36068
rect 17028 36012 17132 36068
rect 17188 36012 17292 36068
rect 17348 36012 17452 36068
rect 17508 36012 17612 36068
rect 17668 36012 17772 36068
rect 17828 36012 17932 36068
rect 17988 36012 18092 36068
rect 18148 36012 18252 36068
rect 18308 36012 18412 36068
rect 18468 36012 18572 36068
rect 18628 36012 18732 36068
rect 18788 36012 18892 36068
rect 18948 36012 20012 36068
rect 20068 36012 20332 36068
rect 20388 36012 20652 36068
rect 20708 36012 20972 36068
rect 21028 36012 21292 36068
rect 21348 36012 21612 36068
rect 21668 36012 21932 36068
rect 21988 36012 23132 36068
rect 23188 36012 23292 36068
rect 23348 36012 23452 36068
rect 23508 36012 23612 36068
rect 23668 36012 23772 36068
rect 23828 36012 23932 36068
rect 23988 36012 24092 36068
rect 24148 36012 24252 36068
rect 24308 36012 24412 36068
rect 24468 36012 24572 36068
rect 24628 36012 24732 36068
rect 24788 36012 24892 36068
rect 24948 36012 25052 36068
rect 25108 36012 25212 36068
rect 25268 36012 25372 36068
rect 25428 36012 25532 36068
rect 25588 36012 25692 36068
rect 25748 36012 25852 36068
rect 25908 36012 26012 36068
rect 26068 36012 26172 36068
rect 26228 36012 26332 36068
rect 26388 36012 26492 36068
rect 26548 36012 26652 36068
rect 26708 36012 26812 36068
rect 26868 36012 26972 36068
rect 27028 36012 27132 36068
rect 27188 36012 27292 36068
rect 27348 36012 27452 36068
rect 27508 36012 27612 36068
rect 27668 36012 27772 36068
rect 27828 36012 27932 36068
rect 27988 36012 28092 36068
rect 28148 36012 28252 36068
rect 28308 36012 28412 36068
rect 28468 36012 28572 36068
rect 28628 36012 28732 36068
rect 28788 36012 28892 36068
rect 28948 36012 29052 36068
rect 29108 36012 29212 36068
rect 29268 36012 29372 36068
rect 29428 36012 30492 36068
rect 30548 36012 30812 36068
rect 30868 36012 31132 36068
rect 31188 36012 31452 36068
rect 31508 36012 31772 36068
rect 31828 36012 32092 36068
rect 32148 36012 32412 36068
rect 32468 36012 33532 36068
rect 33588 36012 33692 36068
rect 33748 36012 33852 36068
rect 33908 36012 34012 36068
rect 34068 36012 34172 36068
rect 34228 36012 34332 36068
rect 34388 36012 34492 36068
rect 34548 36012 34652 36068
rect 34708 36012 34812 36068
rect 34868 36012 34972 36068
rect 35028 36012 35132 36068
rect 35188 36012 35292 36068
rect 35348 36012 35452 36068
rect 35508 36012 35612 36068
rect 35668 36012 35772 36068
rect 35828 36012 35932 36068
rect 35988 36012 36092 36068
rect 36148 36012 36252 36068
rect 36308 36012 36412 36068
rect 36468 36012 36572 36068
rect 36628 36012 36732 36068
rect 36788 36012 36892 36068
rect 36948 36012 37052 36068
rect 37108 36012 37212 36068
rect 37268 36012 37372 36068
rect 37428 36012 37532 36068
rect 37588 36012 37692 36068
rect 37748 36012 37852 36068
rect 37908 36012 38012 36068
rect 38068 36012 38172 36068
rect 38228 36012 38332 36068
rect 38388 36012 38492 36068
rect 38548 36012 38652 36068
rect 38708 36012 38812 36068
rect 38868 36012 38972 36068
rect 39028 36012 39132 36068
rect 39188 36012 39292 36068
rect 39348 36012 39452 36068
rect 39508 36012 39612 36068
rect 39668 36012 39772 36068
rect 39828 36012 39932 36068
rect 39988 36012 40092 36068
rect 40148 36012 40252 36068
rect 40308 36012 40412 36068
rect 40468 36012 40572 36068
rect 40628 36012 40732 36068
rect 40788 36012 40892 36068
rect 40948 36012 41052 36068
rect 41108 36012 41212 36068
rect 41268 36012 41372 36068
rect 41428 36012 41532 36068
rect 41588 36012 41692 36068
rect 41748 36012 41852 36068
rect 41908 36012 41920 36068
rect 0 36000 41920 36012
rect 0 35908 41920 35920
rect 0 35852 9932 35908
rect 9988 35852 21452 35908
rect 21508 35852 31932 35908
rect 31988 35852 41920 35908
rect 0 35840 41920 35852
rect 0 35748 41920 35760
rect 0 35692 12 35748
rect 68 35692 172 35748
rect 228 35692 332 35748
rect 388 35692 492 35748
rect 548 35692 652 35748
rect 708 35692 812 35748
rect 868 35692 972 35748
rect 1028 35692 1132 35748
rect 1188 35692 1292 35748
rect 1348 35692 1452 35748
rect 1508 35692 1612 35748
rect 1668 35692 1772 35748
rect 1828 35692 1932 35748
rect 1988 35692 2092 35748
rect 2148 35692 2252 35748
rect 2308 35692 2412 35748
rect 2468 35692 2572 35748
rect 2628 35692 2732 35748
rect 2788 35692 2892 35748
rect 2948 35692 3052 35748
rect 3108 35692 3212 35748
rect 3268 35692 3372 35748
rect 3428 35692 3532 35748
rect 3588 35692 3692 35748
rect 3748 35692 3852 35748
rect 3908 35692 4012 35748
rect 4068 35692 4172 35748
rect 4228 35692 4332 35748
rect 4388 35692 4492 35748
rect 4548 35692 4652 35748
rect 4708 35692 4812 35748
rect 4868 35692 4972 35748
rect 5028 35692 5132 35748
rect 5188 35692 5292 35748
rect 5348 35692 5452 35748
rect 5508 35692 5612 35748
rect 5668 35692 5772 35748
rect 5828 35692 5932 35748
rect 5988 35692 6092 35748
rect 6148 35692 6252 35748
rect 6308 35692 6412 35748
rect 6468 35692 6572 35748
rect 6628 35692 6732 35748
rect 6788 35692 6892 35748
rect 6948 35692 7052 35748
rect 7108 35692 7212 35748
rect 7268 35692 7372 35748
rect 7428 35692 7532 35748
rect 7588 35692 7692 35748
rect 7748 35692 7852 35748
rect 7908 35692 8012 35748
rect 8068 35692 8172 35748
rect 8228 35692 8332 35748
rect 8388 35692 9452 35748
rect 9508 35692 9772 35748
rect 9828 35692 10092 35748
rect 10148 35692 10412 35748
rect 10468 35692 10732 35748
rect 10788 35692 11052 35748
rect 11108 35692 11372 35748
rect 11428 35692 12492 35748
rect 12548 35692 12652 35748
rect 12708 35692 12812 35748
rect 12868 35692 12972 35748
rect 13028 35692 13132 35748
rect 13188 35692 13292 35748
rect 13348 35692 13452 35748
rect 13508 35692 13612 35748
rect 13668 35692 13772 35748
rect 13828 35692 13932 35748
rect 13988 35692 14092 35748
rect 14148 35692 14252 35748
rect 14308 35692 14412 35748
rect 14468 35692 14572 35748
rect 14628 35692 14732 35748
rect 14788 35692 14892 35748
rect 14948 35692 15052 35748
rect 15108 35692 15212 35748
rect 15268 35692 15372 35748
rect 15428 35692 15532 35748
rect 15588 35692 15692 35748
rect 15748 35692 15852 35748
rect 15908 35692 16012 35748
rect 16068 35692 16172 35748
rect 16228 35692 16332 35748
rect 16388 35692 16492 35748
rect 16548 35692 16652 35748
rect 16708 35692 16812 35748
rect 16868 35692 16972 35748
rect 17028 35692 17132 35748
rect 17188 35692 17292 35748
rect 17348 35692 17452 35748
rect 17508 35692 17612 35748
rect 17668 35692 17772 35748
rect 17828 35692 17932 35748
rect 17988 35692 18092 35748
rect 18148 35692 18252 35748
rect 18308 35692 18412 35748
rect 18468 35692 18572 35748
rect 18628 35692 18732 35748
rect 18788 35692 18892 35748
rect 18948 35692 20012 35748
rect 20068 35692 20332 35748
rect 20388 35692 20652 35748
rect 20708 35692 20972 35748
rect 21028 35692 21292 35748
rect 21348 35692 21612 35748
rect 21668 35692 21932 35748
rect 21988 35692 23132 35748
rect 23188 35692 23292 35748
rect 23348 35692 23452 35748
rect 23508 35692 23612 35748
rect 23668 35692 23772 35748
rect 23828 35692 23932 35748
rect 23988 35692 24092 35748
rect 24148 35692 24252 35748
rect 24308 35692 24412 35748
rect 24468 35692 24572 35748
rect 24628 35692 24732 35748
rect 24788 35692 24892 35748
rect 24948 35692 25052 35748
rect 25108 35692 25212 35748
rect 25268 35692 25372 35748
rect 25428 35692 25532 35748
rect 25588 35692 25692 35748
rect 25748 35692 25852 35748
rect 25908 35692 26012 35748
rect 26068 35692 26172 35748
rect 26228 35692 26332 35748
rect 26388 35692 26492 35748
rect 26548 35692 26652 35748
rect 26708 35692 26812 35748
rect 26868 35692 26972 35748
rect 27028 35692 27132 35748
rect 27188 35692 27292 35748
rect 27348 35692 27452 35748
rect 27508 35692 27612 35748
rect 27668 35692 27772 35748
rect 27828 35692 27932 35748
rect 27988 35692 28092 35748
rect 28148 35692 28252 35748
rect 28308 35692 28412 35748
rect 28468 35692 28572 35748
rect 28628 35692 28732 35748
rect 28788 35692 28892 35748
rect 28948 35692 29052 35748
rect 29108 35692 29212 35748
rect 29268 35692 29372 35748
rect 29428 35692 30492 35748
rect 30548 35692 30812 35748
rect 30868 35692 31132 35748
rect 31188 35692 31452 35748
rect 31508 35692 31772 35748
rect 31828 35692 32092 35748
rect 32148 35692 32412 35748
rect 32468 35692 33532 35748
rect 33588 35692 33692 35748
rect 33748 35692 33852 35748
rect 33908 35692 34012 35748
rect 34068 35692 34172 35748
rect 34228 35692 34332 35748
rect 34388 35692 34492 35748
rect 34548 35692 34652 35748
rect 34708 35692 34812 35748
rect 34868 35692 34972 35748
rect 35028 35692 35132 35748
rect 35188 35692 35292 35748
rect 35348 35692 35452 35748
rect 35508 35692 35612 35748
rect 35668 35692 35772 35748
rect 35828 35692 35932 35748
rect 35988 35692 36092 35748
rect 36148 35692 36252 35748
rect 36308 35692 36412 35748
rect 36468 35692 36572 35748
rect 36628 35692 36732 35748
rect 36788 35692 36892 35748
rect 36948 35692 37052 35748
rect 37108 35692 37212 35748
rect 37268 35692 37372 35748
rect 37428 35692 37532 35748
rect 37588 35692 37692 35748
rect 37748 35692 37852 35748
rect 37908 35692 38012 35748
rect 38068 35692 38172 35748
rect 38228 35692 38332 35748
rect 38388 35692 38492 35748
rect 38548 35692 38652 35748
rect 38708 35692 38812 35748
rect 38868 35692 38972 35748
rect 39028 35692 39132 35748
rect 39188 35692 39292 35748
rect 39348 35692 39452 35748
rect 39508 35692 39612 35748
rect 39668 35692 39772 35748
rect 39828 35692 39932 35748
rect 39988 35692 40092 35748
rect 40148 35692 40252 35748
rect 40308 35692 40412 35748
rect 40468 35692 40572 35748
rect 40628 35692 40732 35748
rect 40788 35692 40892 35748
rect 40948 35692 41052 35748
rect 41108 35692 41212 35748
rect 41268 35692 41372 35748
rect 41428 35692 41532 35748
rect 41588 35692 41692 35748
rect 41748 35692 41852 35748
rect 41908 35692 41920 35748
rect 0 35680 41920 35692
rect 0 35588 41920 35600
rect 0 35532 10252 35588
rect 10308 35532 21132 35588
rect 21188 35532 31612 35588
rect 31668 35532 41920 35588
rect 0 35520 41920 35532
rect 0 35428 41920 35440
rect 0 35372 12 35428
rect 68 35372 172 35428
rect 228 35372 332 35428
rect 388 35372 492 35428
rect 548 35372 652 35428
rect 708 35372 812 35428
rect 868 35372 972 35428
rect 1028 35372 1132 35428
rect 1188 35372 1292 35428
rect 1348 35372 1452 35428
rect 1508 35372 1612 35428
rect 1668 35372 1772 35428
rect 1828 35372 1932 35428
rect 1988 35372 2092 35428
rect 2148 35372 2252 35428
rect 2308 35372 2412 35428
rect 2468 35372 2572 35428
rect 2628 35372 2732 35428
rect 2788 35372 2892 35428
rect 2948 35372 3052 35428
rect 3108 35372 3212 35428
rect 3268 35372 3372 35428
rect 3428 35372 3532 35428
rect 3588 35372 3692 35428
rect 3748 35372 3852 35428
rect 3908 35372 4012 35428
rect 4068 35372 4172 35428
rect 4228 35372 4332 35428
rect 4388 35372 4492 35428
rect 4548 35372 4652 35428
rect 4708 35372 4812 35428
rect 4868 35372 4972 35428
rect 5028 35372 5132 35428
rect 5188 35372 5292 35428
rect 5348 35372 5452 35428
rect 5508 35372 5612 35428
rect 5668 35372 5772 35428
rect 5828 35372 5932 35428
rect 5988 35372 6092 35428
rect 6148 35372 6252 35428
rect 6308 35372 6412 35428
rect 6468 35372 6572 35428
rect 6628 35372 6732 35428
rect 6788 35372 6892 35428
rect 6948 35372 7052 35428
rect 7108 35372 7212 35428
rect 7268 35372 7372 35428
rect 7428 35372 7532 35428
rect 7588 35372 7692 35428
rect 7748 35372 7852 35428
rect 7908 35372 8012 35428
rect 8068 35372 8172 35428
rect 8228 35372 8332 35428
rect 8388 35372 9452 35428
rect 9508 35372 9772 35428
rect 9828 35372 10092 35428
rect 10148 35372 10412 35428
rect 10468 35372 10732 35428
rect 10788 35372 11052 35428
rect 11108 35372 11372 35428
rect 11428 35372 12492 35428
rect 12548 35372 12652 35428
rect 12708 35372 12812 35428
rect 12868 35372 12972 35428
rect 13028 35372 13132 35428
rect 13188 35372 13292 35428
rect 13348 35372 13452 35428
rect 13508 35372 13612 35428
rect 13668 35372 13772 35428
rect 13828 35372 13932 35428
rect 13988 35372 14092 35428
rect 14148 35372 14252 35428
rect 14308 35372 14412 35428
rect 14468 35372 14572 35428
rect 14628 35372 14732 35428
rect 14788 35372 14892 35428
rect 14948 35372 15052 35428
rect 15108 35372 15212 35428
rect 15268 35372 15372 35428
rect 15428 35372 15532 35428
rect 15588 35372 15692 35428
rect 15748 35372 15852 35428
rect 15908 35372 16012 35428
rect 16068 35372 16172 35428
rect 16228 35372 16332 35428
rect 16388 35372 16492 35428
rect 16548 35372 16652 35428
rect 16708 35372 16812 35428
rect 16868 35372 16972 35428
rect 17028 35372 17132 35428
rect 17188 35372 17292 35428
rect 17348 35372 17452 35428
rect 17508 35372 17612 35428
rect 17668 35372 17772 35428
rect 17828 35372 17932 35428
rect 17988 35372 18092 35428
rect 18148 35372 18252 35428
rect 18308 35372 18412 35428
rect 18468 35372 18572 35428
rect 18628 35372 18732 35428
rect 18788 35372 18892 35428
rect 18948 35372 20012 35428
rect 20068 35372 20332 35428
rect 20388 35372 20652 35428
rect 20708 35372 20972 35428
rect 21028 35372 21292 35428
rect 21348 35372 21612 35428
rect 21668 35372 21932 35428
rect 21988 35372 23132 35428
rect 23188 35372 23292 35428
rect 23348 35372 23452 35428
rect 23508 35372 23612 35428
rect 23668 35372 23772 35428
rect 23828 35372 23932 35428
rect 23988 35372 24092 35428
rect 24148 35372 24252 35428
rect 24308 35372 24412 35428
rect 24468 35372 24572 35428
rect 24628 35372 24732 35428
rect 24788 35372 24892 35428
rect 24948 35372 25052 35428
rect 25108 35372 25212 35428
rect 25268 35372 25372 35428
rect 25428 35372 25532 35428
rect 25588 35372 25692 35428
rect 25748 35372 25852 35428
rect 25908 35372 26012 35428
rect 26068 35372 26172 35428
rect 26228 35372 26332 35428
rect 26388 35372 26492 35428
rect 26548 35372 26652 35428
rect 26708 35372 26812 35428
rect 26868 35372 26972 35428
rect 27028 35372 27132 35428
rect 27188 35372 27292 35428
rect 27348 35372 27452 35428
rect 27508 35372 27612 35428
rect 27668 35372 27772 35428
rect 27828 35372 27932 35428
rect 27988 35372 28092 35428
rect 28148 35372 28252 35428
rect 28308 35372 28412 35428
rect 28468 35372 28572 35428
rect 28628 35372 28732 35428
rect 28788 35372 28892 35428
rect 28948 35372 29052 35428
rect 29108 35372 29212 35428
rect 29268 35372 29372 35428
rect 29428 35372 30492 35428
rect 30548 35372 30812 35428
rect 30868 35372 31132 35428
rect 31188 35372 31452 35428
rect 31508 35372 31772 35428
rect 31828 35372 32092 35428
rect 32148 35372 32412 35428
rect 32468 35372 33532 35428
rect 33588 35372 33692 35428
rect 33748 35372 33852 35428
rect 33908 35372 34012 35428
rect 34068 35372 34172 35428
rect 34228 35372 34332 35428
rect 34388 35372 34492 35428
rect 34548 35372 34652 35428
rect 34708 35372 34812 35428
rect 34868 35372 34972 35428
rect 35028 35372 35132 35428
rect 35188 35372 35292 35428
rect 35348 35372 35452 35428
rect 35508 35372 35612 35428
rect 35668 35372 35772 35428
rect 35828 35372 35932 35428
rect 35988 35372 36092 35428
rect 36148 35372 36252 35428
rect 36308 35372 36412 35428
rect 36468 35372 36572 35428
rect 36628 35372 36732 35428
rect 36788 35372 36892 35428
rect 36948 35372 37052 35428
rect 37108 35372 37212 35428
rect 37268 35372 37372 35428
rect 37428 35372 37532 35428
rect 37588 35372 37692 35428
rect 37748 35372 37852 35428
rect 37908 35372 38012 35428
rect 38068 35372 38172 35428
rect 38228 35372 38332 35428
rect 38388 35372 38492 35428
rect 38548 35372 38652 35428
rect 38708 35372 38812 35428
rect 38868 35372 38972 35428
rect 39028 35372 39132 35428
rect 39188 35372 39292 35428
rect 39348 35372 39452 35428
rect 39508 35372 39612 35428
rect 39668 35372 39772 35428
rect 39828 35372 39932 35428
rect 39988 35372 40092 35428
rect 40148 35372 40252 35428
rect 40308 35372 40412 35428
rect 40468 35372 40572 35428
rect 40628 35372 40732 35428
rect 40788 35372 40892 35428
rect 40948 35372 41052 35428
rect 41108 35372 41212 35428
rect 41268 35372 41372 35428
rect 41428 35372 41532 35428
rect 41588 35372 41692 35428
rect 41748 35372 41852 35428
rect 41908 35372 41920 35428
rect 0 35360 41920 35372
rect 0 35268 41920 35280
rect 0 35212 10572 35268
rect 10628 35212 20812 35268
rect 20868 35212 31292 35268
rect 31348 35212 41920 35268
rect 0 35200 41920 35212
rect 0 35108 41920 35120
rect 0 35052 12 35108
rect 68 35052 172 35108
rect 228 35052 332 35108
rect 388 35052 492 35108
rect 548 35052 652 35108
rect 708 35052 812 35108
rect 868 35052 972 35108
rect 1028 35052 1132 35108
rect 1188 35052 1292 35108
rect 1348 35052 1452 35108
rect 1508 35052 1612 35108
rect 1668 35052 1772 35108
rect 1828 35052 1932 35108
rect 1988 35052 2092 35108
rect 2148 35052 2252 35108
rect 2308 35052 2412 35108
rect 2468 35052 2572 35108
rect 2628 35052 2732 35108
rect 2788 35052 2892 35108
rect 2948 35052 3052 35108
rect 3108 35052 3212 35108
rect 3268 35052 3372 35108
rect 3428 35052 3532 35108
rect 3588 35052 3692 35108
rect 3748 35052 3852 35108
rect 3908 35052 4012 35108
rect 4068 35052 4172 35108
rect 4228 35052 4332 35108
rect 4388 35052 4492 35108
rect 4548 35052 4652 35108
rect 4708 35052 4812 35108
rect 4868 35052 4972 35108
rect 5028 35052 5132 35108
rect 5188 35052 5292 35108
rect 5348 35052 5452 35108
rect 5508 35052 5612 35108
rect 5668 35052 5772 35108
rect 5828 35052 5932 35108
rect 5988 35052 6092 35108
rect 6148 35052 6252 35108
rect 6308 35052 6412 35108
rect 6468 35052 6572 35108
rect 6628 35052 6732 35108
rect 6788 35052 6892 35108
rect 6948 35052 7052 35108
rect 7108 35052 7212 35108
rect 7268 35052 7372 35108
rect 7428 35052 7532 35108
rect 7588 35052 7692 35108
rect 7748 35052 7852 35108
rect 7908 35052 8012 35108
rect 8068 35052 8172 35108
rect 8228 35052 8332 35108
rect 8388 35052 9452 35108
rect 9508 35052 9772 35108
rect 9828 35052 10092 35108
rect 10148 35052 10412 35108
rect 10468 35052 10732 35108
rect 10788 35052 11052 35108
rect 11108 35052 11372 35108
rect 11428 35052 12492 35108
rect 12548 35052 12652 35108
rect 12708 35052 12812 35108
rect 12868 35052 12972 35108
rect 13028 35052 13132 35108
rect 13188 35052 13292 35108
rect 13348 35052 13452 35108
rect 13508 35052 13612 35108
rect 13668 35052 13772 35108
rect 13828 35052 13932 35108
rect 13988 35052 14092 35108
rect 14148 35052 14252 35108
rect 14308 35052 14412 35108
rect 14468 35052 14572 35108
rect 14628 35052 14732 35108
rect 14788 35052 14892 35108
rect 14948 35052 15052 35108
rect 15108 35052 15212 35108
rect 15268 35052 15372 35108
rect 15428 35052 15532 35108
rect 15588 35052 15692 35108
rect 15748 35052 15852 35108
rect 15908 35052 16012 35108
rect 16068 35052 16172 35108
rect 16228 35052 16332 35108
rect 16388 35052 16492 35108
rect 16548 35052 16652 35108
rect 16708 35052 16812 35108
rect 16868 35052 16972 35108
rect 17028 35052 17132 35108
rect 17188 35052 17292 35108
rect 17348 35052 17452 35108
rect 17508 35052 17612 35108
rect 17668 35052 17772 35108
rect 17828 35052 17932 35108
rect 17988 35052 18092 35108
rect 18148 35052 18252 35108
rect 18308 35052 18412 35108
rect 18468 35052 18572 35108
rect 18628 35052 18732 35108
rect 18788 35052 18892 35108
rect 18948 35052 20012 35108
rect 20068 35052 20332 35108
rect 20388 35052 20652 35108
rect 20708 35052 20972 35108
rect 21028 35052 21292 35108
rect 21348 35052 21612 35108
rect 21668 35052 21932 35108
rect 21988 35052 23132 35108
rect 23188 35052 23292 35108
rect 23348 35052 23452 35108
rect 23508 35052 23612 35108
rect 23668 35052 23772 35108
rect 23828 35052 23932 35108
rect 23988 35052 24092 35108
rect 24148 35052 24252 35108
rect 24308 35052 24412 35108
rect 24468 35052 24572 35108
rect 24628 35052 24732 35108
rect 24788 35052 24892 35108
rect 24948 35052 25052 35108
rect 25108 35052 25212 35108
rect 25268 35052 25372 35108
rect 25428 35052 25532 35108
rect 25588 35052 25692 35108
rect 25748 35052 25852 35108
rect 25908 35052 26012 35108
rect 26068 35052 26172 35108
rect 26228 35052 26332 35108
rect 26388 35052 26492 35108
rect 26548 35052 26652 35108
rect 26708 35052 26812 35108
rect 26868 35052 26972 35108
rect 27028 35052 27132 35108
rect 27188 35052 27292 35108
rect 27348 35052 27452 35108
rect 27508 35052 27612 35108
rect 27668 35052 27772 35108
rect 27828 35052 27932 35108
rect 27988 35052 28092 35108
rect 28148 35052 28252 35108
rect 28308 35052 28412 35108
rect 28468 35052 28572 35108
rect 28628 35052 28732 35108
rect 28788 35052 28892 35108
rect 28948 35052 29052 35108
rect 29108 35052 29212 35108
rect 29268 35052 29372 35108
rect 29428 35052 30492 35108
rect 30548 35052 30812 35108
rect 30868 35052 31132 35108
rect 31188 35052 31452 35108
rect 31508 35052 31772 35108
rect 31828 35052 32092 35108
rect 32148 35052 32412 35108
rect 32468 35052 33532 35108
rect 33588 35052 33692 35108
rect 33748 35052 33852 35108
rect 33908 35052 34012 35108
rect 34068 35052 34172 35108
rect 34228 35052 34332 35108
rect 34388 35052 34492 35108
rect 34548 35052 34652 35108
rect 34708 35052 34812 35108
rect 34868 35052 34972 35108
rect 35028 35052 35132 35108
rect 35188 35052 35292 35108
rect 35348 35052 35452 35108
rect 35508 35052 35612 35108
rect 35668 35052 35772 35108
rect 35828 35052 35932 35108
rect 35988 35052 36092 35108
rect 36148 35052 36252 35108
rect 36308 35052 36412 35108
rect 36468 35052 36572 35108
rect 36628 35052 36732 35108
rect 36788 35052 36892 35108
rect 36948 35052 37052 35108
rect 37108 35052 37212 35108
rect 37268 35052 37372 35108
rect 37428 35052 37532 35108
rect 37588 35052 37692 35108
rect 37748 35052 37852 35108
rect 37908 35052 38012 35108
rect 38068 35052 38172 35108
rect 38228 35052 38332 35108
rect 38388 35052 38492 35108
rect 38548 35052 38652 35108
rect 38708 35052 38812 35108
rect 38868 35052 38972 35108
rect 39028 35052 39132 35108
rect 39188 35052 39292 35108
rect 39348 35052 39452 35108
rect 39508 35052 39612 35108
rect 39668 35052 39772 35108
rect 39828 35052 39932 35108
rect 39988 35052 40092 35108
rect 40148 35052 40252 35108
rect 40308 35052 40412 35108
rect 40468 35052 40572 35108
rect 40628 35052 40732 35108
rect 40788 35052 40892 35108
rect 40948 35052 41052 35108
rect 41108 35052 41212 35108
rect 41268 35052 41372 35108
rect 41428 35052 41532 35108
rect 41588 35052 41692 35108
rect 41748 35052 41852 35108
rect 41908 35052 41920 35108
rect 0 35040 41920 35052
rect 0 34948 41920 34960
rect 0 34892 10892 34948
rect 10948 34892 20492 34948
rect 20548 34892 30972 34948
rect 31028 34892 41920 34948
rect 0 34880 41920 34892
rect 0 34788 41920 34800
rect 0 34732 12 34788
rect 68 34732 172 34788
rect 228 34732 332 34788
rect 388 34732 492 34788
rect 548 34732 652 34788
rect 708 34732 812 34788
rect 868 34732 972 34788
rect 1028 34732 1132 34788
rect 1188 34732 1292 34788
rect 1348 34732 1452 34788
rect 1508 34732 1612 34788
rect 1668 34732 1772 34788
rect 1828 34732 1932 34788
rect 1988 34732 2092 34788
rect 2148 34732 2252 34788
rect 2308 34732 2412 34788
rect 2468 34732 2572 34788
rect 2628 34732 2732 34788
rect 2788 34732 2892 34788
rect 2948 34732 3052 34788
rect 3108 34732 3212 34788
rect 3268 34732 3372 34788
rect 3428 34732 3532 34788
rect 3588 34732 3692 34788
rect 3748 34732 3852 34788
rect 3908 34732 4012 34788
rect 4068 34732 4172 34788
rect 4228 34732 4332 34788
rect 4388 34732 4492 34788
rect 4548 34732 4652 34788
rect 4708 34732 4812 34788
rect 4868 34732 4972 34788
rect 5028 34732 5132 34788
rect 5188 34732 5292 34788
rect 5348 34732 5452 34788
rect 5508 34732 5612 34788
rect 5668 34732 5772 34788
rect 5828 34732 5932 34788
rect 5988 34732 6092 34788
rect 6148 34732 6252 34788
rect 6308 34732 6412 34788
rect 6468 34732 6572 34788
rect 6628 34732 6732 34788
rect 6788 34732 6892 34788
rect 6948 34732 7052 34788
rect 7108 34732 7212 34788
rect 7268 34732 7372 34788
rect 7428 34732 7532 34788
rect 7588 34732 7692 34788
rect 7748 34732 7852 34788
rect 7908 34732 8012 34788
rect 8068 34732 8172 34788
rect 8228 34732 8332 34788
rect 8388 34732 9452 34788
rect 9508 34732 9772 34788
rect 9828 34732 10092 34788
rect 10148 34732 10412 34788
rect 10468 34732 10732 34788
rect 10788 34732 11052 34788
rect 11108 34732 11372 34788
rect 11428 34732 12492 34788
rect 12548 34732 12652 34788
rect 12708 34732 12812 34788
rect 12868 34732 12972 34788
rect 13028 34732 13132 34788
rect 13188 34732 13292 34788
rect 13348 34732 13452 34788
rect 13508 34732 13612 34788
rect 13668 34732 13772 34788
rect 13828 34732 13932 34788
rect 13988 34732 14092 34788
rect 14148 34732 14252 34788
rect 14308 34732 14412 34788
rect 14468 34732 14572 34788
rect 14628 34732 14732 34788
rect 14788 34732 14892 34788
rect 14948 34732 15052 34788
rect 15108 34732 15212 34788
rect 15268 34732 15372 34788
rect 15428 34732 15532 34788
rect 15588 34732 15692 34788
rect 15748 34732 15852 34788
rect 15908 34732 16012 34788
rect 16068 34732 16172 34788
rect 16228 34732 16332 34788
rect 16388 34732 16492 34788
rect 16548 34732 16652 34788
rect 16708 34732 16812 34788
rect 16868 34732 16972 34788
rect 17028 34732 17132 34788
rect 17188 34732 17292 34788
rect 17348 34732 17452 34788
rect 17508 34732 17612 34788
rect 17668 34732 17772 34788
rect 17828 34732 17932 34788
rect 17988 34732 18092 34788
rect 18148 34732 18252 34788
rect 18308 34732 18412 34788
rect 18468 34732 18572 34788
rect 18628 34732 18732 34788
rect 18788 34732 18892 34788
rect 18948 34732 20012 34788
rect 20068 34732 20332 34788
rect 20388 34732 20652 34788
rect 20708 34732 20972 34788
rect 21028 34732 21292 34788
rect 21348 34732 21612 34788
rect 21668 34732 21932 34788
rect 21988 34732 23132 34788
rect 23188 34732 23292 34788
rect 23348 34732 23452 34788
rect 23508 34732 23612 34788
rect 23668 34732 23772 34788
rect 23828 34732 23932 34788
rect 23988 34732 24092 34788
rect 24148 34732 24252 34788
rect 24308 34732 24412 34788
rect 24468 34732 24572 34788
rect 24628 34732 24732 34788
rect 24788 34732 24892 34788
rect 24948 34732 25052 34788
rect 25108 34732 25212 34788
rect 25268 34732 25372 34788
rect 25428 34732 25532 34788
rect 25588 34732 25692 34788
rect 25748 34732 25852 34788
rect 25908 34732 26012 34788
rect 26068 34732 26172 34788
rect 26228 34732 26332 34788
rect 26388 34732 26492 34788
rect 26548 34732 26652 34788
rect 26708 34732 26812 34788
rect 26868 34732 26972 34788
rect 27028 34732 27132 34788
rect 27188 34732 27292 34788
rect 27348 34732 27452 34788
rect 27508 34732 27612 34788
rect 27668 34732 27772 34788
rect 27828 34732 27932 34788
rect 27988 34732 28092 34788
rect 28148 34732 28252 34788
rect 28308 34732 28412 34788
rect 28468 34732 28572 34788
rect 28628 34732 28732 34788
rect 28788 34732 28892 34788
rect 28948 34732 29052 34788
rect 29108 34732 29212 34788
rect 29268 34732 29372 34788
rect 29428 34732 30492 34788
rect 30548 34732 30812 34788
rect 30868 34732 31132 34788
rect 31188 34732 31452 34788
rect 31508 34732 31772 34788
rect 31828 34732 32092 34788
rect 32148 34732 32412 34788
rect 32468 34732 33532 34788
rect 33588 34732 33692 34788
rect 33748 34732 33852 34788
rect 33908 34732 34012 34788
rect 34068 34732 34172 34788
rect 34228 34732 34332 34788
rect 34388 34732 34492 34788
rect 34548 34732 34652 34788
rect 34708 34732 34812 34788
rect 34868 34732 34972 34788
rect 35028 34732 35132 34788
rect 35188 34732 35292 34788
rect 35348 34732 35452 34788
rect 35508 34732 35612 34788
rect 35668 34732 35772 34788
rect 35828 34732 35932 34788
rect 35988 34732 36092 34788
rect 36148 34732 36252 34788
rect 36308 34732 36412 34788
rect 36468 34732 36572 34788
rect 36628 34732 36732 34788
rect 36788 34732 36892 34788
rect 36948 34732 37052 34788
rect 37108 34732 37212 34788
rect 37268 34732 37372 34788
rect 37428 34732 37532 34788
rect 37588 34732 37692 34788
rect 37748 34732 37852 34788
rect 37908 34732 38012 34788
rect 38068 34732 38172 34788
rect 38228 34732 38332 34788
rect 38388 34732 38492 34788
rect 38548 34732 38652 34788
rect 38708 34732 38812 34788
rect 38868 34732 38972 34788
rect 39028 34732 39132 34788
rect 39188 34732 39292 34788
rect 39348 34732 39452 34788
rect 39508 34732 39612 34788
rect 39668 34732 39772 34788
rect 39828 34732 39932 34788
rect 39988 34732 40092 34788
rect 40148 34732 40252 34788
rect 40308 34732 40412 34788
rect 40468 34732 40572 34788
rect 40628 34732 40732 34788
rect 40788 34732 40892 34788
rect 40948 34732 41052 34788
rect 41108 34732 41212 34788
rect 41268 34732 41372 34788
rect 41428 34732 41532 34788
rect 41588 34732 41692 34788
rect 41748 34732 41852 34788
rect 41908 34732 41920 34788
rect 0 34720 41920 34732
rect 0 34628 41920 34640
rect 0 34572 11212 34628
rect 11268 34572 20172 34628
rect 20228 34572 30652 34628
rect 30708 34572 41920 34628
rect 0 34560 41920 34572
rect 0 34468 41920 34480
rect 0 34412 12 34468
rect 68 34412 172 34468
rect 228 34412 332 34468
rect 388 34412 492 34468
rect 548 34412 652 34468
rect 708 34412 812 34468
rect 868 34412 972 34468
rect 1028 34412 1132 34468
rect 1188 34412 1292 34468
rect 1348 34412 1452 34468
rect 1508 34412 1612 34468
rect 1668 34412 1772 34468
rect 1828 34412 1932 34468
rect 1988 34412 2092 34468
rect 2148 34412 2252 34468
rect 2308 34412 2412 34468
rect 2468 34412 2572 34468
rect 2628 34412 2732 34468
rect 2788 34412 2892 34468
rect 2948 34412 3052 34468
rect 3108 34412 3212 34468
rect 3268 34412 3372 34468
rect 3428 34412 3532 34468
rect 3588 34412 3692 34468
rect 3748 34412 3852 34468
rect 3908 34412 4012 34468
rect 4068 34412 4172 34468
rect 4228 34412 4332 34468
rect 4388 34412 4492 34468
rect 4548 34412 4652 34468
rect 4708 34412 4812 34468
rect 4868 34412 4972 34468
rect 5028 34412 5132 34468
rect 5188 34412 5292 34468
rect 5348 34412 5452 34468
rect 5508 34412 5612 34468
rect 5668 34412 5772 34468
rect 5828 34412 5932 34468
rect 5988 34412 6092 34468
rect 6148 34412 6252 34468
rect 6308 34412 6412 34468
rect 6468 34412 6572 34468
rect 6628 34412 6732 34468
rect 6788 34412 6892 34468
rect 6948 34412 7052 34468
rect 7108 34412 7212 34468
rect 7268 34412 7372 34468
rect 7428 34412 7532 34468
rect 7588 34412 7692 34468
rect 7748 34412 7852 34468
rect 7908 34412 8012 34468
rect 8068 34412 8172 34468
rect 8228 34412 8332 34468
rect 8388 34412 9452 34468
rect 9508 34412 9772 34468
rect 9828 34412 10092 34468
rect 10148 34412 10412 34468
rect 10468 34412 10732 34468
rect 10788 34412 11052 34468
rect 11108 34412 11372 34468
rect 11428 34412 12492 34468
rect 12548 34412 12652 34468
rect 12708 34412 12812 34468
rect 12868 34412 12972 34468
rect 13028 34412 13132 34468
rect 13188 34412 13292 34468
rect 13348 34412 13452 34468
rect 13508 34412 13612 34468
rect 13668 34412 13772 34468
rect 13828 34412 13932 34468
rect 13988 34412 14092 34468
rect 14148 34412 14252 34468
rect 14308 34412 14412 34468
rect 14468 34412 14572 34468
rect 14628 34412 14732 34468
rect 14788 34412 14892 34468
rect 14948 34412 15052 34468
rect 15108 34412 15212 34468
rect 15268 34412 15372 34468
rect 15428 34412 15532 34468
rect 15588 34412 15692 34468
rect 15748 34412 15852 34468
rect 15908 34412 16012 34468
rect 16068 34412 16172 34468
rect 16228 34412 16332 34468
rect 16388 34412 16492 34468
rect 16548 34412 16652 34468
rect 16708 34412 16812 34468
rect 16868 34412 16972 34468
rect 17028 34412 17132 34468
rect 17188 34412 17292 34468
rect 17348 34412 17452 34468
rect 17508 34412 17612 34468
rect 17668 34412 17772 34468
rect 17828 34412 17932 34468
rect 17988 34412 18092 34468
rect 18148 34412 18252 34468
rect 18308 34412 18412 34468
rect 18468 34412 18572 34468
rect 18628 34412 18732 34468
rect 18788 34412 18892 34468
rect 18948 34412 20012 34468
rect 20068 34412 20332 34468
rect 20388 34412 20652 34468
rect 20708 34412 20972 34468
rect 21028 34412 21292 34468
rect 21348 34412 21612 34468
rect 21668 34412 21932 34468
rect 21988 34412 23132 34468
rect 23188 34412 23292 34468
rect 23348 34412 23452 34468
rect 23508 34412 23612 34468
rect 23668 34412 23772 34468
rect 23828 34412 23932 34468
rect 23988 34412 24092 34468
rect 24148 34412 24252 34468
rect 24308 34412 24412 34468
rect 24468 34412 24572 34468
rect 24628 34412 24732 34468
rect 24788 34412 24892 34468
rect 24948 34412 25052 34468
rect 25108 34412 25212 34468
rect 25268 34412 25372 34468
rect 25428 34412 25532 34468
rect 25588 34412 25692 34468
rect 25748 34412 25852 34468
rect 25908 34412 26012 34468
rect 26068 34412 26172 34468
rect 26228 34412 26332 34468
rect 26388 34412 26492 34468
rect 26548 34412 26652 34468
rect 26708 34412 26812 34468
rect 26868 34412 26972 34468
rect 27028 34412 27132 34468
rect 27188 34412 27292 34468
rect 27348 34412 27452 34468
rect 27508 34412 27612 34468
rect 27668 34412 27772 34468
rect 27828 34412 27932 34468
rect 27988 34412 28092 34468
rect 28148 34412 28252 34468
rect 28308 34412 28412 34468
rect 28468 34412 28572 34468
rect 28628 34412 28732 34468
rect 28788 34412 28892 34468
rect 28948 34412 29052 34468
rect 29108 34412 29212 34468
rect 29268 34412 29372 34468
rect 29428 34412 30492 34468
rect 30548 34412 30812 34468
rect 30868 34412 31132 34468
rect 31188 34412 31452 34468
rect 31508 34412 31772 34468
rect 31828 34412 32092 34468
rect 32148 34412 32412 34468
rect 32468 34412 33532 34468
rect 33588 34412 33692 34468
rect 33748 34412 33852 34468
rect 33908 34412 34012 34468
rect 34068 34412 34172 34468
rect 34228 34412 34332 34468
rect 34388 34412 34492 34468
rect 34548 34412 34652 34468
rect 34708 34412 34812 34468
rect 34868 34412 34972 34468
rect 35028 34412 35132 34468
rect 35188 34412 35292 34468
rect 35348 34412 35452 34468
rect 35508 34412 35612 34468
rect 35668 34412 35772 34468
rect 35828 34412 35932 34468
rect 35988 34412 36092 34468
rect 36148 34412 36252 34468
rect 36308 34412 36412 34468
rect 36468 34412 36572 34468
rect 36628 34412 36732 34468
rect 36788 34412 36892 34468
rect 36948 34412 37052 34468
rect 37108 34412 37212 34468
rect 37268 34412 37372 34468
rect 37428 34412 37532 34468
rect 37588 34412 37692 34468
rect 37748 34412 37852 34468
rect 37908 34412 38012 34468
rect 38068 34412 38172 34468
rect 38228 34412 38332 34468
rect 38388 34412 38492 34468
rect 38548 34412 38652 34468
rect 38708 34412 38812 34468
rect 38868 34412 38972 34468
rect 39028 34412 39132 34468
rect 39188 34412 39292 34468
rect 39348 34412 39452 34468
rect 39508 34412 39612 34468
rect 39668 34412 39772 34468
rect 39828 34412 39932 34468
rect 39988 34412 40092 34468
rect 40148 34412 40252 34468
rect 40308 34412 40412 34468
rect 40468 34412 40572 34468
rect 40628 34412 40732 34468
rect 40788 34412 40892 34468
rect 40948 34412 41052 34468
rect 41108 34412 41212 34468
rect 41268 34412 41372 34468
rect 41428 34412 41532 34468
rect 41588 34412 41692 34468
rect 41748 34412 41852 34468
rect 41908 34412 41920 34468
rect 0 34400 41920 34412
rect 0 34308 41920 34320
rect 0 34252 12 34308
rect 68 34252 172 34308
rect 228 34252 332 34308
rect 388 34252 492 34308
rect 548 34252 652 34308
rect 708 34252 812 34308
rect 868 34252 972 34308
rect 1028 34252 1132 34308
rect 1188 34252 1292 34308
rect 1348 34252 1452 34308
rect 1508 34252 1612 34308
rect 1668 34252 1772 34308
rect 1828 34252 1932 34308
rect 1988 34252 2092 34308
rect 2148 34252 2252 34308
rect 2308 34252 2412 34308
rect 2468 34252 2572 34308
rect 2628 34252 2732 34308
rect 2788 34252 2892 34308
rect 2948 34252 3052 34308
rect 3108 34252 3212 34308
rect 3268 34252 3372 34308
rect 3428 34252 3532 34308
rect 3588 34252 3692 34308
rect 3748 34252 3852 34308
rect 3908 34252 4012 34308
rect 4068 34252 4172 34308
rect 4228 34252 4332 34308
rect 4388 34252 4492 34308
rect 4548 34252 4652 34308
rect 4708 34252 4812 34308
rect 4868 34252 4972 34308
rect 5028 34252 5132 34308
rect 5188 34252 5292 34308
rect 5348 34252 5452 34308
rect 5508 34252 5612 34308
rect 5668 34252 5772 34308
rect 5828 34252 5932 34308
rect 5988 34252 6092 34308
rect 6148 34252 6252 34308
rect 6308 34252 6412 34308
rect 6468 34252 6572 34308
rect 6628 34252 6732 34308
rect 6788 34252 6892 34308
rect 6948 34252 7052 34308
rect 7108 34252 7212 34308
rect 7268 34252 7372 34308
rect 7428 34252 7532 34308
rect 7588 34252 7692 34308
rect 7748 34252 7852 34308
rect 7908 34252 8012 34308
rect 8068 34252 8172 34308
rect 8228 34252 8332 34308
rect 8388 34252 11532 34308
rect 11588 34252 11852 34308
rect 11908 34252 12492 34308
rect 12548 34252 12652 34308
rect 12708 34252 12812 34308
rect 12868 34252 12972 34308
rect 13028 34252 13132 34308
rect 13188 34252 13292 34308
rect 13348 34252 13452 34308
rect 13508 34252 13612 34308
rect 13668 34252 13772 34308
rect 13828 34252 13932 34308
rect 13988 34252 14092 34308
rect 14148 34252 14252 34308
rect 14308 34252 14412 34308
rect 14468 34252 14572 34308
rect 14628 34252 14732 34308
rect 14788 34252 14892 34308
rect 14948 34252 15052 34308
rect 15108 34252 15212 34308
rect 15268 34252 15372 34308
rect 15428 34252 15532 34308
rect 15588 34252 15692 34308
rect 15748 34252 15852 34308
rect 15908 34252 16012 34308
rect 16068 34252 16172 34308
rect 16228 34252 16332 34308
rect 16388 34252 16492 34308
rect 16548 34252 16652 34308
rect 16708 34252 16812 34308
rect 16868 34252 16972 34308
rect 17028 34252 17132 34308
rect 17188 34252 17292 34308
rect 17348 34252 17452 34308
rect 17508 34252 17612 34308
rect 17668 34252 17772 34308
rect 17828 34252 17932 34308
rect 17988 34252 18092 34308
rect 18148 34252 18252 34308
rect 18308 34252 18412 34308
rect 18468 34252 18572 34308
rect 18628 34252 18732 34308
rect 18788 34252 18892 34308
rect 18948 34252 19532 34308
rect 19588 34252 19852 34308
rect 19908 34252 23132 34308
rect 23188 34252 23292 34308
rect 23348 34252 23452 34308
rect 23508 34252 23612 34308
rect 23668 34252 23772 34308
rect 23828 34252 23932 34308
rect 23988 34252 24092 34308
rect 24148 34252 24252 34308
rect 24308 34252 24412 34308
rect 24468 34252 24572 34308
rect 24628 34252 24732 34308
rect 24788 34252 24892 34308
rect 24948 34252 25052 34308
rect 25108 34252 25212 34308
rect 25268 34252 25372 34308
rect 25428 34252 25532 34308
rect 25588 34252 25692 34308
rect 25748 34252 25852 34308
rect 25908 34252 26012 34308
rect 26068 34252 26172 34308
rect 26228 34252 26332 34308
rect 26388 34252 26492 34308
rect 26548 34252 26652 34308
rect 26708 34252 26812 34308
rect 26868 34252 26972 34308
rect 27028 34252 27132 34308
rect 27188 34252 27292 34308
rect 27348 34252 27452 34308
rect 27508 34252 27612 34308
rect 27668 34252 27772 34308
rect 27828 34252 27932 34308
rect 27988 34252 28092 34308
rect 28148 34252 28252 34308
rect 28308 34252 28412 34308
rect 28468 34252 28572 34308
rect 28628 34252 28732 34308
rect 28788 34252 28892 34308
rect 28948 34252 29052 34308
rect 29108 34252 29212 34308
rect 29268 34252 29372 34308
rect 29428 34252 30012 34308
rect 30068 34252 30332 34308
rect 30388 34252 33532 34308
rect 33588 34252 33692 34308
rect 33748 34252 33852 34308
rect 33908 34252 34012 34308
rect 34068 34252 34172 34308
rect 34228 34252 34332 34308
rect 34388 34252 34492 34308
rect 34548 34252 34652 34308
rect 34708 34252 34812 34308
rect 34868 34252 34972 34308
rect 35028 34252 35132 34308
rect 35188 34252 35292 34308
rect 35348 34252 35452 34308
rect 35508 34252 35612 34308
rect 35668 34252 35772 34308
rect 35828 34252 35932 34308
rect 35988 34252 36092 34308
rect 36148 34252 36252 34308
rect 36308 34252 36412 34308
rect 36468 34252 36572 34308
rect 36628 34252 36732 34308
rect 36788 34252 36892 34308
rect 36948 34252 37052 34308
rect 37108 34252 37212 34308
rect 37268 34252 37372 34308
rect 37428 34252 37532 34308
rect 37588 34252 37692 34308
rect 37748 34252 37852 34308
rect 37908 34252 38012 34308
rect 38068 34252 38172 34308
rect 38228 34252 38332 34308
rect 38388 34252 38492 34308
rect 38548 34252 38652 34308
rect 38708 34252 38812 34308
rect 38868 34252 38972 34308
rect 39028 34252 39132 34308
rect 39188 34252 39292 34308
rect 39348 34252 39452 34308
rect 39508 34252 39612 34308
rect 39668 34252 39772 34308
rect 39828 34252 39932 34308
rect 39988 34252 40092 34308
rect 40148 34252 40252 34308
rect 40308 34252 40412 34308
rect 40468 34252 40572 34308
rect 40628 34252 40732 34308
rect 40788 34252 40892 34308
rect 40948 34252 41052 34308
rect 41108 34252 41212 34308
rect 41268 34252 41372 34308
rect 41428 34252 41532 34308
rect 41588 34252 41692 34308
rect 41748 34252 41852 34308
rect 41908 34252 41920 34308
rect 0 34240 41920 34252
rect 0 34148 41920 34160
rect 0 34092 11692 34148
rect 11748 34092 19692 34148
rect 19748 34092 30172 34148
rect 30228 34092 41920 34148
rect 0 34080 41920 34092
rect 0 33988 41920 34000
rect 0 33932 12 33988
rect 68 33932 172 33988
rect 228 33932 332 33988
rect 388 33932 492 33988
rect 548 33932 652 33988
rect 708 33932 812 33988
rect 868 33932 972 33988
rect 1028 33932 1132 33988
rect 1188 33932 1292 33988
rect 1348 33932 1452 33988
rect 1508 33932 1612 33988
rect 1668 33932 1772 33988
rect 1828 33932 1932 33988
rect 1988 33932 2092 33988
rect 2148 33932 2252 33988
rect 2308 33932 2412 33988
rect 2468 33932 2572 33988
rect 2628 33932 2732 33988
rect 2788 33932 2892 33988
rect 2948 33932 3052 33988
rect 3108 33932 3212 33988
rect 3268 33932 3372 33988
rect 3428 33932 3532 33988
rect 3588 33932 3692 33988
rect 3748 33932 3852 33988
rect 3908 33932 4012 33988
rect 4068 33932 4172 33988
rect 4228 33932 4332 33988
rect 4388 33932 4492 33988
rect 4548 33932 4652 33988
rect 4708 33932 4812 33988
rect 4868 33932 4972 33988
rect 5028 33932 5132 33988
rect 5188 33932 5292 33988
rect 5348 33932 5452 33988
rect 5508 33932 5612 33988
rect 5668 33932 5772 33988
rect 5828 33932 5932 33988
rect 5988 33932 6092 33988
rect 6148 33932 6252 33988
rect 6308 33932 6412 33988
rect 6468 33932 6572 33988
rect 6628 33932 6732 33988
rect 6788 33932 6892 33988
rect 6948 33932 7052 33988
rect 7108 33932 7212 33988
rect 7268 33932 7372 33988
rect 7428 33932 7532 33988
rect 7588 33932 7692 33988
rect 7748 33932 7852 33988
rect 7908 33932 8012 33988
rect 8068 33932 8172 33988
rect 8228 33932 8332 33988
rect 8388 33932 11532 33988
rect 11588 33932 11852 33988
rect 11908 33932 12492 33988
rect 12548 33932 12652 33988
rect 12708 33932 12812 33988
rect 12868 33932 12972 33988
rect 13028 33932 13132 33988
rect 13188 33932 13292 33988
rect 13348 33932 13452 33988
rect 13508 33932 13612 33988
rect 13668 33932 13772 33988
rect 13828 33932 13932 33988
rect 13988 33932 14092 33988
rect 14148 33932 14252 33988
rect 14308 33932 14412 33988
rect 14468 33932 14572 33988
rect 14628 33932 14732 33988
rect 14788 33932 14892 33988
rect 14948 33932 15052 33988
rect 15108 33932 15212 33988
rect 15268 33932 15372 33988
rect 15428 33932 15532 33988
rect 15588 33932 15692 33988
rect 15748 33932 15852 33988
rect 15908 33932 16012 33988
rect 16068 33932 16172 33988
rect 16228 33932 16332 33988
rect 16388 33932 16492 33988
rect 16548 33932 16652 33988
rect 16708 33932 16812 33988
rect 16868 33932 16972 33988
rect 17028 33932 17132 33988
rect 17188 33932 17292 33988
rect 17348 33932 17452 33988
rect 17508 33932 17612 33988
rect 17668 33932 17772 33988
rect 17828 33932 17932 33988
rect 17988 33932 18092 33988
rect 18148 33932 18252 33988
rect 18308 33932 18412 33988
rect 18468 33932 18572 33988
rect 18628 33932 18732 33988
rect 18788 33932 18892 33988
rect 18948 33932 19532 33988
rect 19588 33932 19852 33988
rect 19908 33932 23132 33988
rect 23188 33932 23292 33988
rect 23348 33932 23452 33988
rect 23508 33932 23612 33988
rect 23668 33932 23772 33988
rect 23828 33932 23932 33988
rect 23988 33932 24092 33988
rect 24148 33932 24252 33988
rect 24308 33932 24412 33988
rect 24468 33932 24572 33988
rect 24628 33932 24732 33988
rect 24788 33932 24892 33988
rect 24948 33932 25052 33988
rect 25108 33932 25212 33988
rect 25268 33932 25372 33988
rect 25428 33932 25532 33988
rect 25588 33932 25692 33988
rect 25748 33932 25852 33988
rect 25908 33932 26012 33988
rect 26068 33932 26172 33988
rect 26228 33932 26332 33988
rect 26388 33932 26492 33988
rect 26548 33932 26652 33988
rect 26708 33932 26812 33988
rect 26868 33932 26972 33988
rect 27028 33932 27132 33988
rect 27188 33932 27292 33988
rect 27348 33932 27452 33988
rect 27508 33932 27612 33988
rect 27668 33932 27772 33988
rect 27828 33932 27932 33988
rect 27988 33932 28092 33988
rect 28148 33932 28252 33988
rect 28308 33932 28412 33988
rect 28468 33932 28572 33988
rect 28628 33932 28732 33988
rect 28788 33932 28892 33988
rect 28948 33932 29052 33988
rect 29108 33932 29212 33988
rect 29268 33932 29372 33988
rect 29428 33932 30012 33988
rect 30068 33932 30332 33988
rect 30388 33932 33532 33988
rect 33588 33932 33692 33988
rect 33748 33932 33852 33988
rect 33908 33932 34012 33988
rect 34068 33932 34172 33988
rect 34228 33932 34332 33988
rect 34388 33932 34492 33988
rect 34548 33932 34652 33988
rect 34708 33932 34812 33988
rect 34868 33932 34972 33988
rect 35028 33932 35132 33988
rect 35188 33932 35292 33988
rect 35348 33932 35452 33988
rect 35508 33932 35612 33988
rect 35668 33932 35772 33988
rect 35828 33932 35932 33988
rect 35988 33932 36092 33988
rect 36148 33932 36252 33988
rect 36308 33932 36412 33988
rect 36468 33932 36572 33988
rect 36628 33932 36732 33988
rect 36788 33932 36892 33988
rect 36948 33932 37052 33988
rect 37108 33932 37212 33988
rect 37268 33932 37372 33988
rect 37428 33932 37532 33988
rect 37588 33932 37692 33988
rect 37748 33932 37852 33988
rect 37908 33932 38012 33988
rect 38068 33932 38172 33988
rect 38228 33932 38332 33988
rect 38388 33932 38492 33988
rect 38548 33932 38652 33988
rect 38708 33932 38812 33988
rect 38868 33932 38972 33988
rect 39028 33932 39132 33988
rect 39188 33932 39292 33988
rect 39348 33932 39452 33988
rect 39508 33932 39612 33988
rect 39668 33932 39772 33988
rect 39828 33932 39932 33988
rect 39988 33932 40092 33988
rect 40148 33932 40252 33988
rect 40308 33932 40412 33988
rect 40468 33932 40572 33988
rect 40628 33932 40732 33988
rect 40788 33932 40892 33988
rect 40948 33932 41052 33988
rect 41108 33932 41212 33988
rect 41268 33932 41372 33988
rect 41428 33932 41532 33988
rect 41588 33932 41692 33988
rect 41748 33932 41852 33988
rect 41908 33932 41920 33988
rect 0 33920 41920 33932
rect 0 33828 41920 33840
rect 0 33772 12 33828
rect 68 33772 172 33828
rect 228 33772 332 33828
rect 388 33772 492 33828
rect 548 33772 652 33828
rect 708 33772 812 33828
rect 868 33772 972 33828
rect 1028 33772 1132 33828
rect 1188 33772 1292 33828
rect 1348 33772 1452 33828
rect 1508 33772 1612 33828
rect 1668 33772 1772 33828
rect 1828 33772 1932 33828
rect 1988 33772 2092 33828
rect 2148 33772 2252 33828
rect 2308 33772 2412 33828
rect 2468 33772 2572 33828
rect 2628 33772 2732 33828
rect 2788 33772 2892 33828
rect 2948 33772 3052 33828
rect 3108 33772 3212 33828
rect 3268 33772 3372 33828
rect 3428 33772 3532 33828
rect 3588 33772 3692 33828
rect 3748 33772 3852 33828
rect 3908 33772 4012 33828
rect 4068 33772 4172 33828
rect 4228 33772 4332 33828
rect 4388 33772 4492 33828
rect 4548 33772 4652 33828
rect 4708 33772 4812 33828
rect 4868 33772 4972 33828
rect 5028 33772 5132 33828
rect 5188 33772 5292 33828
rect 5348 33772 5452 33828
rect 5508 33772 5612 33828
rect 5668 33772 5772 33828
rect 5828 33772 5932 33828
rect 5988 33772 6092 33828
rect 6148 33772 6252 33828
rect 6308 33772 6412 33828
rect 6468 33772 6572 33828
rect 6628 33772 6732 33828
rect 6788 33772 6892 33828
rect 6948 33772 7052 33828
rect 7108 33772 7212 33828
rect 7268 33772 7372 33828
rect 7428 33772 7532 33828
rect 7588 33772 7692 33828
rect 7748 33772 7852 33828
rect 7908 33772 8012 33828
rect 8068 33772 8172 33828
rect 8228 33772 8332 33828
rect 8388 33772 12012 33828
rect 12068 33772 12332 33828
rect 12388 33772 12492 33828
rect 12548 33772 12652 33828
rect 12708 33772 12812 33828
rect 12868 33772 12972 33828
rect 13028 33772 13132 33828
rect 13188 33772 13292 33828
rect 13348 33772 13452 33828
rect 13508 33772 13612 33828
rect 13668 33772 13772 33828
rect 13828 33772 13932 33828
rect 13988 33772 14092 33828
rect 14148 33772 14252 33828
rect 14308 33772 14412 33828
rect 14468 33772 14572 33828
rect 14628 33772 14732 33828
rect 14788 33772 14892 33828
rect 14948 33772 15052 33828
rect 15108 33772 15212 33828
rect 15268 33772 15372 33828
rect 15428 33772 15532 33828
rect 15588 33772 15692 33828
rect 15748 33772 15852 33828
rect 15908 33772 16012 33828
rect 16068 33772 16172 33828
rect 16228 33772 16332 33828
rect 16388 33772 16492 33828
rect 16548 33772 16652 33828
rect 16708 33772 16812 33828
rect 16868 33772 16972 33828
rect 17028 33772 17132 33828
rect 17188 33772 17292 33828
rect 17348 33772 17452 33828
rect 17508 33772 17612 33828
rect 17668 33772 17772 33828
rect 17828 33772 17932 33828
rect 17988 33772 18092 33828
rect 18148 33772 18252 33828
rect 18308 33772 18412 33828
rect 18468 33772 18572 33828
rect 18628 33772 18732 33828
rect 18788 33772 18892 33828
rect 18948 33772 19052 33828
rect 19108 33772 19372 33828
rect 19428 33772 23132 33828
rect 23188 33772 23292 33828
rect 23348 33772 23452 33828
rect 23508 33772 23612 33828
rect 23668 33772 23772 33828
rect 23828 33772 23932 33828
rect 23988 33772 24092 33828
rect 24148 33772 24252 33828
rect 24308 33772 24412 33828
rect 24468 33772 24572 33828
rect 24628 33772 24732 33828
rect 24788 33772 24892 33828
rect 24948 33772 25052 33828
rect 25108 33772 25212 33828
rect 25268 33772 25372 33828
rect 25428 33772 25532 33828
rect 25588 33772 25692 33828
rect 25748 33772 25852 33828
rect 25908 33772 26012 33828
rect 26068 33772 26172 33828
rect 26228 33772 26332 33828
rect 26388 33772 26492 33828
rect 26548 33772 26652 33828
rect 26708 33772 26812 33828
rect 26868 33772 26972 33828
rect 27028 33772 27132 33828
rect 27188 33772 27292 33828
rect 27348 33772 27452 33828
rect 27508 33772 27612 33828
rect 27668 33772 27772 33828
rect 27828 33772 27932 33828
rect 27988 33772 28092 33828
rect 28148 33772 28252 33828
rect 28308 33772 28412 33828
rect 28468 33772 28572 33828
rect 28628 33772 28732 33828
rect 28788 33772 28892 33828
rect 28948 33772 29052 33828
rect 29108 33772 29212 33828
rect 29268 33772 29372 33828
rect 29428 33772 29532 33828
rect 29588 33772 29852 33828
rect 29908 33772 33532 33828
rect 33588 33772 33692 33828
rect 33748 33772 33852 33828
rect 33908 33772 34012 33828
rect 34068 33772 34172 33828
rect 34228 33772 34332 33828
rect 34388 33772 34492 33828
rect 34548 33772 34652 33828
rect 34708 33772 34812 33828
rect 34868 33772 34972 33828
rect 35028 33772 35132 33828
rect 35188 33772 35292 33828
rect 35348 33772 35452 33828
rect 35508 33772 35612 33828
rect 35668 33772 35772 33828
rect 35828 33772 35932 33828
rect 35988 33772 36092 33828
rect 36148 33772 36252 33828
rect 36308 33772 36412 33828
rect 36468 33772 36572 33828
rect 36628 33772 36732 33828
rect 36788 33772 36892 33828
rect 36948 33772 37052 33828
rect 37108 33772 37212 33828
rect 37268 33772 37372 33828
rect 37428 33772 37532 33828
rect 37588 33772 37692 33828
rect 37748 33772 37852 33828
rect 37908 33772 38012 33828
rect 38068 33772 38172 33828
rect 38228 33772 38332 33828
rect 38388 33772 38492 33828
rect 38548 33772 38652 33828
rect 38708 33772 38812 33828
rect 38868 33772 38972 33828
rect 39028 33772 39132 33828
rect 39188 33772 39292 33828
rect 39348 33772 39452 33828
rect 39508 33772 39612 33828
rect 39668 33772 39772 33828
rect 39828 33772 39932 33828
rect 39988 33772 40092 33828
rect 40148 33772 40252 33828
rect 40308 33772 40412 33828
rect 40468 33772 40572 33828
rect 40628 33772 40732 33828
rect 40788 33772 40892 33828
rect 40948 33772 41052 33828
rect 41108 33772 41212 33828
rect 41268 33772 41372 33828
rect 41428 33772 41532 33828
rect 41588 33772 41692 33828
rect 41748 33772 41852 33828
rect 41908 33772 41920 33828
rect 0 33760 41920 33772
rect 0 33668 41920 33680
rect 0 33612 12172 33668
rect 12228 33612 19212 33668
rect 19268 33612 29692 33668
rect 29748 33612 41920 33668
rect 0 33600 41920 33612
rect 0 33508 41920 33520
rect 0 33452 12 33508
rect 68 33452 172 33508
rect 228 33452 332 33508
rect 388 33452 492 33508
rect 548 33452 652 33508
rect 708 33452 812 33508
rect 868 33452 972 33508
rect 1028 33452 1132 33508
rect 1188 33452 1292 33508
rect 1348 33452 1452 33508
rect 1508 33452 1612 33508
rect 1668 33452 1772 33508
rect 1828 33452 1932 33508
rect 1988 33452 2092 33508
rect 2148 33452 2252 33508
rect 2308 33452 2412 33508
rect 2468 33452 2572 33508
rect 2628 33452 2732 33508
rect 2788 33452 2892 33508
rect 2948 33452 3052 33508
rect 3108 33452 3212 33508
rect 3268 33452 3372 33508
rect 3428 33452 3532 33508
rect 3588 33452 3692 33508
rect 3748 33452 3852 33508
rect 3908 33452 4012 33508
rect 4068 33452 4172 33508
rect 4228 33452 4332 33508
rect 4388 33452 4492 33508
rect 4548 33452 4652 33508
rect 4708 33452 4812 33508
rect 4868 33452 4972 33508
rect 5028 33452 5132 33508
rect 5188 33452 5292 33508
rect 5348 33452 5452 33508
rect 5508 33452 5612 33508
rect 5668 33452 5772 33508
rect 5828 33452 5932 33508
rect 5988 33452 6092 33508
rect 6148 33452 6252 33508
rect 6308 33452 6412 33508
rect 6468 33452 6572 33508
rect 6628 33452 6732 33508
rect 6788 33452 6892 33508
rect 6948 33452 7052 33508
rect 7108 33452 7212 33508
rect 7268 33452 7372 33508
rect 7428 33452 7532 33508
rect 7588 33452 7692 33508
rect 7748 33452 7852 33508
rect 7908 33452 8012 33508
rect 8068 33452 8172 33508
rect 8228 33452 8332 33508
rect 8388 33452 12012 33508
rect 12068 33452 12332 33508
rect 12388 33452 12492 33508
rect 12548 33452 12652 33508
rect 12708 33452 12812 33508
rect 12868 33452 12972 33508
rect 13028 33452 13132 33508
rect 13188 33452 13292 33508
rect 13348 33452 13452 33508
rect 13508 33452 13612 33508
rect 13668 33452 13772 33508
rect 13828 33452 13932 33508
rect 13988 33452 14092 33508
rect 14148 33452 14252 33508
rect 14308 33452 14412 33508
rect 14468 33452 14572 33508
rect 14628 33452 14732 33508
rect 14788 33452 14892 33508
rect 14948 33452 15052 33508
rect 15108 33452 15212 33508
rect 15268 33452 15372 33508
rect 15428 33452 15532 33508
rect 15588 33452 15692 33508
rect 15748 33452 15852 33508
rect 15908 33452 16012 33508
rect 16068 33452 16172 33508
rect 16228 33452 16332 33508
rect 16388 33452 16492 33508
rect 16548 33452 16652 33508
rect 16708 33452 16812 33508
rect 16868 33452 16972 33508
rect 17028 33452 17132 33508
rect 17188 33452 17292 33508
rect 17348 33452 17452 33508
rect 17508 33452 17612 33508
rect 17668 33452 17772 33508
rect 17828 33452 17932 33508
rect 17988 33452 18092 33508
rect 18148 33452 18252 33508
rect 18308 33452 18412 33508
rect 18468 33452 18572 33508
rect 18628 33452 18732 33508
rect 18788 33452 18892 33508
rect 18948 33452 19052 33508
rect 19108 33452 19372 33508
rect 19428 33452 23132 33508
rect 23188 33452 23292 33508
rect 23348 33452 23452 33508
rect 23508 33452 23612 33508
rect 23668 33452 23772 33508
rect 23828 33452 23932 33508
rect 23988 33452 24092 33508
rect 24148 33452 24252 33508
rect 24308 33452 24412 33508
rect 24468 33452 24572 33508
rect 24628 33452 24732 33508
rect 24788 33452 24892 33508
rect 24948 33452 25052 33508
rect 25108 33452 25212 33508
rect 25268 33452 25372 33508
rect 25428 33452 25532 33508
rect 25588 33452 25692 33508
rect 25748 33452 25852 33508
rect 25908 33452 26012 33508
rect 26068 33452 26172 33508
rect 26228 33452 26332 33508
rect 26388 33452 26492 33508
rect 26548 33452 26652 33508
rect 26708 33452 26812 33508
rect 26868 33452 26972 33508
rect 27028 33452 27132 33508
rect 27188 33452 27292 33508
rect 27348 33452 27452 33508
rect 27508 33452 27612 33508
rect 27668 33452 27772 33508
rect 27828 33452 27932 33508
rect 27988 33452 28092 33508
rect 28148 33452 28252 33508
rect 28308 33452 28412 33508
rect 28468 33452 28572 33508
rect 28628 33452 28732 33508
rect 28788 33452 28892 33508
rect 28948 33452 29052 33508
rect 29108 33452 29212 33508
rect 29268 33452 29372 33508
rect 29428 33452 29532 33508
rect 29588 33452 29852 33508
rect 29908 33452 33532 33508
rect 33588 33452 33692 33508
rect 33748 33452 33852 33508
rect 33908 33452 34012 33508
rect 34068 33452 34172 33508
rect 34228 33452 34332 33508
rect 34388 33452 34492 33508
rect 34548 33452 34652 33508
rect 34708 33452 34812 33508
rect 34868 33452 34972 33508
rect 35028 33452 35132 33508
rect 35188 33452 35292 33508
rect 35348 33452 35452 33508
rect 35508 33452 35612 33508
rect 35668 33452 35772 33508
rect 35828 33452 35932 33508
rect 35988 33452 36092 33508
rect 36148 33452 36252 33508
rect 36308 33452 36412 33508
rect 36468 33452 36572 33508
rect 36628 33452 36732 33508
rect 36788 33452 36892 33508
rect 36948 33452 37052 33508
rect 37108 33452 37212 33508
rect 37268 33452 37372 33508
rect 37428 33452 37532 33508
rect 37588 33452 37692 33508
rect 37748 33452 37852 33508
rect 37908 33452 38012 33508
rect 38068 33452 38172 33508
rect 38228 33452 38332 33508
rect 38388 33452 38492 33508
rect 38548 33452 38652 33508
rect 38708 33452 38812 33508
rect 38868 33452 38972 33508
rect 39028 33452 39132 33508
rect 39188 33452 39292 33508
rect 39348 33452 39452 33508
rect 39508 33452 39612 33508
rect 39668 33452 39772 33508
rect 39828 33452 39932 33508
rect 39988 33452 40092 33508
rect 40148 33452 40252 33508
rect 40308 33452 40412 33508
rect 40468 33452 40572 33508
rect 40628 33452 40732 33508
rect 40788 33452 40892 33508
rect 40948 33452 41052 33508
rect 41108 33452 41212 33508
rect 41268 33452 41372 33508
rect 41428 33452 41532 33508
rect 41588 33452 41692 33508
rect 41748 33452 41852 33508
rect 41908 33452 41920 33508
rect 0 33440 41920 33452
rect 0 33348 41920 33360
rect 0 33292 12 33348
rect 68 33292 172 33348
rect 228 33292 332 33348
rect 388 33292 492 33348
rect 548 33292 652 33348
rect 708 33292 812 33348
rect 868 33292 972 33348
rect 1028 33292 1132 33348
rect 1188 33292 1292 33348
rect 1348 33292 1452 33348
rect 1508 33292 1612 33348
rect 1668 33292 1772 33348
rect 1828 33292 1932 33348
rect 1988 33292 2092 33348
rect 2148 33292 2252 33348
rect 2308 33292 2412 33348
rect 2468 33292 2572 33348
rect 2628 33292 2732 33348
rect 2788 33292 2892 33348
rect 2948 33292 3052 33348
rect 3108 33292 3212 33348
rect 3268 33292 3372 33348
rect 3428 33292 3532 33348
rect 3588 33292 3692 33348
rect 3748 33292 3852 33348
rect 3908 33292 4012 33348
rect 4068 33292 4172 33348
rect 4228 33292 4332 33348
rect 4388 33292 4492 33348
rect 4548 33292 4652 33348
rect 4708 33292 4812 33348
rect 4868 33292 4972 33348
rect 5028 33292 5132 33348
rect 5188 33292 5292 33348
rect 5348 33292 5452 33348
rect 5508 33292 5612 33348
rect 5668 33292 5772 33348
rect 5828 33292 5932 33348
rect 5988 33292 6092 33348
rect 6148 33292 6252 33348
rect 6308 33292 6412 33348
rect 6468 33292 6572 33348
rect 6628 33292 6732 33348
rect 6788 33292 6892 33348
rect 6948 33292 7052 33348
rect 7108 33292 7212 33348
rect 7268 33292 7372 33348
rect 7428 33292 7532 33348
rect 7588 33292 7692 33348
rect 7748 33292 7852 33348
rect 7908 33292 8012 33348
rect 8068 33292 8172 33348
rect 8228 33292 8332 33348
rect 8388 33292 8492 33348
rect 8548 33292 8812 33348
rect 8868 33292 12492 33348
rect 12548 33292 12652 33348
rect 12708 33292 12812 33348
rect 12868 33292 12972 33348
rect 13028 33292 13132 33348
rect 13188 33292 13292 33348
rect 13348 33292 13452 33348
rect 13508 33292 13612 33348
rect 13668 33292 13772 33348
rect 13828 33292 13932 33348
rect 13988 33292 14092 33348
rect 14148 33292 14252 33348
rect 14308 33292 14412 33348
rect 14468 33292 14572 33348
rect 14628 33292 14732 33348
rect 14788 33292 14892 33348
rect 14948 33292 15052 33348
rect 15108 33292 15212 33348
rect 15268 33292 15372 33348
rect 15428 33292 15532 33348
rect 15588 33292 15692 33348
rect 15748 33292 15852 33348
rect 15908 33292 16012 33348
rect 16068 33292 16172 33348
rect 16228 33292 16332 33348
rect 16388 33292 16492 33348
rect 16548 33292 16652 33348
rect 16708 33292 16812 33348
rect 16868 33292 16972 33348
rect 17028 33292 17132 33348
rect 17188 33292 17292 33348
rect 17348 33292 17452 33348
rect 17508 33292 17612 33348
rect 17668 33292 17772 33348
rect 17828 33292 17932 33348
rect 17988 33292 18092 33348
rect 18148 33292 18252 33348
rect 18308 33292 18412 33348
rect 18468 33292 18572 33348
rect 18628 33292 18732 33348
rect 18788 33292 18892 33348
rect 18948 33292 19052 33348
rect 19108 33292 19372 33348
rect 19428 33292 23132 33348
rect 23188 33292 23292 33348
rect 23348 33292 23452 33348
rect 23508 33292 23612 33348
rect 23668 33292 23772 33348
rect 23828 33292 23932 33348
rect 23988 33292 24092 33348
rect 24148 33292 24252 33348
rect 24308 33292 24412 33348
rect 24468 33292 24572 33348
rect 24628 33292 24732 33348
rect 24788 33292 24892 33348
rect 24948 33292 25052 33348
rect 25108 33292 25212 33348
rect 25268 33292 25372 33348
rect 25428 33292 25532 33348
rect 25588 33292 25692 33348
rect 25748 33292 25852 33348
rect 25908 33292 26012 33348
rect 26068 33292 26172 33348
rect 26228 33292 26332 33348
rect 26388 33292 26492 33348
rect 26548 33292 26652 33348
rect 26708 33292 26812 33348
rect 26868 33292 26972 33348
rect 27028 33292 27132 33348
rect 27188 33292 27292 33348
rect 27348 33292 27452 33348
rect 27508 33292 27612 33348
rect 27668 33292 27772 33348
rect 27828 33292 27932 33348
rect 27988 33292 28092 33348
rect 28148 33292 28252 33348
rect 28308 33292 28412 33348
rect 28468 33292 28572 33348
rect 28628 33292 28732 33348
rect 28788 33292 28892 33348
rect 28948 33292 29052 33348
rect 29108 33292 29212 33348
rect 29268 33292 29372 33348
rect 29428 33292 33052 33348
rect 33108 33292 33372 33348
rect 33428 33292 33532 33348
rect 33588 33292 33692 33348
rect 33748 33292 33852 33348
rect 33908 33292 34012 33348
rect 34068 33292 34172 33348
rect 34228 33292 34332 33348
rect 34388 33292 34492 33348
rect 34548 33292 34652 33348
rect 34708 33292 34812 33348
rect 34868 33292 34972 33348
rect 35028 33292 35132 33348
rect 35188 33292 35292 33348
rect 35348 33292 35452 33348
rect 35508 33292 35612 33348
rect 35668 33292 35772 33348
rect 35828 33292 35932 33348
rect 35988 33292 36092 33348
rect 36148 33292 36252 33348
rect 36308 33292 36412 33348
rect 36468 33292 36572 33348
rect 36628 33292 36732 33348
rect 36788 33292 36892 33348
rect 36948 33292 37052 33348
rect 37108 33292 37212 33348
rect 37268 33292 37372 33348
rect 37428 33292 37532 33348
rect 37588 33292 37692 33348
rect 37748 33292 37852 33348
rect 37908 33292 38012 33348
rect 38068 33292 38172 33348
rect 38228 33292 38332 33348
rect 38388 33292 38492 33348
rect 38548 33292 38652 33348
rect 38708 33292 38812 33348
rect 38868 33292 38972 33348
rect 39028 33292 39132 33348
rect 39188 33292 39292 33348
rect 39348 33292 39452 33348
rect 39508 33292 39612 33348
rect 39668 33292 39772 33348
rect 39828 33292 39932 33348
rect 39988 33292 40092 33348
rect 40148 33292 40252 33348
rect 40308 33292 40412 33348
rect 40468 33292 40572 33348
rect 40628 33292 40732 33348
rect 40788 33292 40892 33348
rect 40948 33292 41052 33348
rect 41108 33292 41212 33348
rect 41268 33292 41372 33348
rect 41428 33292 41532 33348
rect 41588 33292 41692 33348
rect 41748 33292 41852 33348
rect 41908 33292 41920 33348
rect 0 33280 41920 33292
rect 0 33188 41920 33200
rect 0 33132 8652 33188
rect 8708 33132 19212 33188
rect 19268 33132 33212 33188
rect 33268 33132 41920 33188
rect 0 33120 41920 33132
rect 0 33028 41920 33040
rect 0 32972 12 33028
rect 68 32972 172 33028
rect 228 32972 332 33028
rect 388 32972 492 33028
rect 548 32972 652 33028
rect 708 32972 812 33028
rect 868 32972 972 33028
rect 1028 32972 1132 33028
rect 1188 32972 1292 33028
rect 1348 32972 1452 33028
rect 1508 32972 1612 33028
rect 1668 32972 1772 33028
rect 1828 32972 1932 33028
rect 1988 32972 2092 33028
rect 2148 32972 2252 33028
rect 2308 32972 2412 33028
rect 2468 32972 2572 33028
rect 2628 32972 2732 33028
rect 2788 32972 2892 33028
rect 2948 32972 3052 33028
rect 3108 32972 3212 33028
rect 3268 32972 3372 33028
rect 3428 32972 3532 33028
rect 3588 32972 3692 33028
rect 3748 32972 3852 33028
rect 3908 32972 4012 33028
rect 4068 32972 4172 33028
rect 4228 32972 4332 33028
rect 4388 32972 4492 33028
rect 4548 32972 4652 33028
rect 4708 32972 4812 33028
rect 4868 32972 4972 33028
rect 5028 32972 5132 33028
rect 5188 32972 5292 33028
rect 5348 32972 5452 33028
rect 5508 32972 5612 33028
rect 5668 32972 5772 33028
rect 5828 32972 5932 33028
rect 5988 32972 6092 33028
rect 6148 32972 6252 33028
rect 6308 32972 6412 33028
rect 6468 32972 6572 33028
rect 6628 32972 6732 33028
rect 6788 32972 6892 33028
rect 6948 32972 7052 33028
rect 7108 32972 7212 33028
rect 7268 32972 7372 33028
rect 7428 32972 7532 33028
rect 7588 32972 7692 33028
rect 7748 32972 7852 33028
rect 7908 32972 8012 33028
rect 8068 32972 8172 33028
rect 8228 32972 8332 33028
rect 8388 32972 8492 33028
rect 8548 32972 8812 33028
rect 8868 32972 12492 33028
rect 12548 32972 12652 33028
rect 12708 32972 12812 33028
rect 12868 32972 12972 33028
rect 13028 32972 13132 33028
rect 13188 32972 13292 33028
rect 13348 32972 13452 33028
rect 13508 32972 13612 33028
rect 13668 32972 13772 33028
rect 13828 32972 13932 33028
rect 13988 32972 14092 33028
rect 14148 32972 14252 33028
rect 14308 32972 14412 33028
rect 14468 32972 14572 33028
rect 14628 32972 14732 33028
rect 14788 32972 14892 33028
rect 14948 32972 15052 33028
rect 15108 32972 15212 33028
rect 15268 32972 15372 33028
rect 15428 32972 15532 33028
rect 15588 32972 15692 33028
rect 15748 32972 15852 33028
rect 15908 32972 16012 33028
rect 16068 32972 16172 33028
rect 16228 32972 16332 33028
rect 16388 32972 16492 33028
rect 16548 32972 16652 33028
rect 16708 32972 16812 33028
rect 16868 32972 16972 33028
rect 17028 32972 17132 33028
rect 17188 32972 17292 33028
rect 17348 32972 17452 33028
rect 17508 32972 17612 33028
rect 17668 32972 17772 33028
rect 17828 32972 17932 33028
rect 17988 32972 18092 33028
rect 18148 32972 18252 33028
rect 18308 32972 18412 33028
rect 18468 32972 18572 33028
rect 18628 32972 18732 33028
rect 18788 32972 18892 33028
rect 18948 32972 19052 33028
rect 19108 32972 19372 33028
rect 19428 32972 23132 33028
rect 23188 32972 23292 33028
rect 23348 32972 23452 33028
rect 23508 32972 23612 33028
rect 23668 32972 23772 33028
rect 23828 32972 23932 33028
rect 23988 32972 24092 33028
rect 24148 32972 24252 33028
rect 24308 32972 24412 33028
rect 24468 32972 24572 33028
rect 24628 32972 24732 33028
rect 24788 32972 24892 33028
rect 24948 32972 25052 33028
rect 25108 32972 25212 33028
rect 25268 32972 25372 33028
rect 25428 32972 25532 33028
rect 25588 32972 25692 33028
rect 25748 32972 25852 33028
rect 25908 32972 26012 33028
rect 26068 32972 26172 33028
rect 26228 32972 26332 33028
rect 26388 32972 26492 33028
rect 26548 32972 26652 33028
rect 26708 32972 26812 33028
rect 26868 32972 26972 33028
rect 27028 32972 27132 33028
rect 27188 32972 27292 33028
rect 27348 32972 27452 33028
rect 27508 32972 27612 33028
rect 27668 32972 27772 33028
rect 27828 32972 27932 33028
rect 27988 32972 28092 33028
rect 28148 32972 28252 33028
rect 28308 32972 28412 33028
rect 28468 32972 28572 33028
rect 28628 32972 28732 33028
rect 28788 32972 28892 33028
rect 28948 32972 29052 33028
rect 29108 32972 29212 33028
rect 29268 32972 29372 33028
rect 29428 32972 33052 33028
rect 33108 32972 33372 33028
rect 33428 32972 33532 33028
rect 33588 32972 33692 33028
rect 33748 32972 33852 33028
rect 33908 32972 34012 33028
rect 34068 32972 34172 33028
rect 34228 32972 34332 33028
rect 34388 32972 34492 33028
rect 34548 32972 34652 33028
rect 34708 32972 34812 33028
rect 34868 32972 34972 33028
rect 35028 32972 35132 33028
rect 35188 32972 35292 33028
rect 35348 32972 35452 33028
rect 35508 32972 35612 33028
rect 35668 32972 35772 33028
rect 35828 32972 35932 33028
rect 35988 32972 36092 33028
rect 36148 32972 36252 33028
rect 36308 32972 36412 33028
rect 36468 32972 36572 33028
rect 36628 32972 36732 33028
rect 36788 32972 36892 33028
rect 36948 32972 37052 33028
rect 37108 32972 37212 33028
rect 37268 32972 37372 33028
rect 37428 32972 37532 33028
rect 37588 32972 37692 33028
rect 37748 32972 37852 33028
rect 37908 32972 38012 33028
rect 38068 32972 38172 33028
rect 38228 32972 38332 33028
rect 38388 32972 38492 33028
rect 38548 32972 38652 33028
rect 38708 32972 38812 33028
rect 38868 32972 38972 33028
rect 39028 32972 39132 33028
rect 39188 32972 39292 33028
rect 39348 32972 39452 33028
rect 39508 32972 39612 33028
rect 39668 32972 39772 33028
rect 39828 32972 39932 33028
rect 39988 32972 40092 33028
rect 40148 32972 40252 33028
rect 40308 32972 40412 33028
rect 40468 32972 40572 33028
rect 40628 32972 40732 33028
rect 40788 32972 40892 33028
rect 40948 32972 41052 33028
rect 41108 32972 41212 33028
rect 41268 32972 41372 33028
rect 41428 32972 41532 33028
rect 41588 32972 41692 33028
rect 41748 32972 41852 33028
rect 41908 32972 41920 33028
rect 0 32960 41920 32972
rect 0 32868 41920 32880
rect 0 32812 12 32868
rect 68 32812 172 32868
rect 228 32812 332 32868
rect 388 32812 492 32868
rect 548 32812 652 32868
rect 708 32812 812 32868
rect 868 32812 972 32868
rect 1028 32812 1132 32868
rect 1188 32812 1292 32868
rect 1348 32812 1452 32868
rect 1508 32812 1612 32868
rect 1668 32812 1772 32868
rect 1828 32812 1932 32868
rect 1988 32812 2092 32868
rect 2148 32812 2252 32868
rect 2308 32812 2412 32868
rect 2468 32812 2572 32868
rect 2628 32812 2732 32868
rect 2788 32812 2892 32868
rect 2948 32812 3052 32868
rect 3108 32812 3212 32868
rect 3268 32812 3372 32868
rect 3428 32812 3532 32868
rect 3588 32812 3692 32868
rect 3748 32812 3852 32868
rect 3908 32812 4012 32868
rect 4068 32812 4172 32868
rect 4228 32812 4332 32868
rect 4388 32812 4492 32868
rect 4548 32812 4652 32868
rect 4708 32812 4812 32868
rect 4868 32812 4972 32868
rect 5028 32812 5132 32868
rect 5188 32812 5292 32868
rect 5348 32812 5452 32868
rect 5508 32812 5612 32868
rect 5668 32812 5772 32868
rect 5828 32812 5932 32868
rect 5988 32812 6092 32868
rect 6148 32812 6252 32868
rect 6308 32812 6412 32868
rect 6468 32812 6572 32868
rect 6628 32812 6732 32868
rect 6788 32812 6892 32868
rect 6948 32812 7052 32868
rect 7108 32812 7212 32868
rect 7268 32812 7372 32868
rect 7428 32812 7532 32868
rect 7588 32812 7692 32868
rect 7748 32812 7852 32868
rect 7908 32812 8012 32868
rect 8068 32812 8172 32868
rect 8228 32812 8332 32868
rect 8388 32812 8972 32868
rect 9028 32812 9292 32868
rect 9348 32812 12492 32868
rect 12548 32812 12652 32868
rect 12708 32812 12812 32868
rect 12868 32812 12972 32868
rect 13028 32812 13132 32868
rect 13188 32812 13292 32868
rect 13348 32812 13452 32868
rect 13508 32812 13612 32868
rect 13668 32812 13772 32868
rect 13828 32812 13932 32868
rect 13988 32812 14092 32868
rect 14148 32812 14252 32868
rect 14308 32812 14412 32868
rect 14468 32812 14572 32868
rect 14628 32812 14732 32868
rect 14788 32812 14892 32868
rect 14948 32812 15052 32868
rect 15108 32812 15212 32868
rect 15268 32812 15372 32868
rect 15428 32812 15532 32868
rect 15588 32812 15692 32868
rect 15748 32812 15852 32868
rect 15908 32812 16012 32868
rect 16068 32812 16172 32868
rect 16228 32812 16332 32868
rect 16388 32812 16492 32868
rect 16548 32812 16652 32868
rect 16708 32812 16812 32868
rect 16868 32812 16972 32868
rect 17028 32812 17132 32868
rect 17188 32812 17292 32868
rect 17348 32812 17452 32868
rect 17508 32812 17612 32868
rect 17668 32812 17772 32868
rect 17828 32812 17932 32868
rect 17988 32812 18092 32868
rect 18148 32812 18252 32868
rect 18308 32812 18412 32868
rect 18468 32812 18572 32868
rect 18628 32812 18732 32868
rect 18788 32812 18892 32868
rect 18948 32812 19532 32868
rect 19588 32812 19852 32868
rect 19908 32812 23132 32868
rect 23188 32812 23292 32868
rect 23348 32812 23452 32868
rect 23508 32812 23612 32868
rect 23668 32812 23772 32868
rect 23828 32812 23932 32868
rect 23988 32812 24092 32868
rect 24148 32812 24252 32868
rect 24308 32812 24412 32868
rect 24468 32812 24572 32868
rect 24628 32812 24732 32868
rect 24788 32812 24892 32868
rect 24948 32812 25052 32868
rect 25108 32812 25212 32868
rect 25268 32812 25372 32868
rect 25428 32812 25532 32868
rect 25588 32812 25692 32868
rect 25748 32812 25852 32868
rect 25908 32812 26012 32868
rect 26068 32812 26172 32868
rect 26228 32812 26332 32868
rect 26388 32812 26492 32868
rect 26548 32812 26652 32868
rect 26708 32812 26812 32868
rect 26868 32812 26972 32868
rect 27028 32812 27132 32868
rect 27188 32812 27292 32868
rect 27348 32812 27452 32868
rect 27508 32812 27612 32868
rect 27668 32812 27772 32868
rect 27828 32812 27932 32868
rect 27988 32812 28092 32868
rect 28148 32812 28252 32868
rect 28308 32812 28412 32868
rect 28468 32812 28572 32868
rect 28628 32812 28732 32868
rect 28788 32812 28892 32868
rect 28948 32812 29052 32868
rect 29108 32812 29212 32868
rect 29268 32812 29372 32868
rect 29428 32812 32572 32868
rect 32628 32812 32892 32868
rect 32948 32812 33532 32868
rect 33588 32812 33692 32868
rect 33748 32812 33852 32868
rect 33908 32812 34012 32868
rect 34068 32812 34172 32868
rect 34228 32812 34332 32868
rect 34388 32812 34492 32868
rect 34548 32812 34652 32868
rect 34708 32812 34812 32868
rect 34868 32812 34972 32868
rect 35028 32812 35132 32868
rect 35188 32812 35292 32868
rect 35348 32812 35452 32868
rect 35508 32812 35612 32868
rect 35668 32812 35772 32868
rect 35828 32812 35932 32868
rect 35988 32812 36092 32868
rect 36148 32812 36252 32868
rect 36308 32812 36412 32868
rect 36468 32812 36572 32868
rect 36628 32812 36732 32868
rect 36788 32812 36892 32868
rect 36948 32812 37052 32868
rect 37108 32812 37212 32868
rect 37268 32812 37372 32868
rect 37428 32812 37532 32868
rect 37588 32812 37692 32868
rect 37748 32812 37852 32868
rect 37908 32812 38012 32868
rect 38068 32812 38172 32868
rect 38228 32812 38332 32868
rect 38388 32812 38492 32868
rect 38548 32812 38652 32868
rect 38708 32812 38812 32868
rect 38868 32812 38972 32868
rect 39028 32812 39132 32868
rect 39188 32812 39292 32868
rect 39348 32812 39452 32868
rect 39508 32812 39612 32868
rect 39668 32812 39772 32868
rect 39828 32812 39932 32868
rect 39988 32812 40092 32868
rect 40148 32812 40252 32868
rect 40308 32812 40412 32868
rect 40468 32812 40572 32868
rect 40628 32812 40732 32868
rect 40788 32812 40892 32868
rect 40948 32812 41052 32868
rect 41108 32812 41212 32868
rect 41268 32812 41372 32868
rect 41428 32812 41532 32868
rect 41588 32812 41692 32868
rect 41748 32812 41852 32868
rect 41908 32812 41920 32868
rect 0 32800 41920 32812
rect 0 32708 41920 32720
rect 0 32652 9132 32708
rect 9188 32652 19692 32708
rect 19748 32652 32732 32708
rect 32788 32652 41920 32708
rect 0 32640 41920 32652
rect 0 32548 41920 32560
rect 0 32492 12 32548
rect 68 32492 172 32548
rect 228 32492 332 32548
rect 388 32492 492 32548
rect 548 32492 652 32548
rect 708 32492 812 32548
rect 868 32492 972 32548
rect 1028 32492 1132 32548
rect 1188 32492 1292 32548
rect 1348 32492 1452 32548
rect 1508 32492 1612 32548
rect 1668 32492 1772 32548
rect 1828 32492 1932 32548
rect 1988 32492 2092 32548
rect 2148 32492 2252 32548
rect 2308 32492 2412 32548
rect 2468 32492 2572 32548
rect 2628 32492 2732 32548
rect 2788 32492 2892 32548
rect 2948 32492 3052 32548
rect 3108 32492 3212 32548
rect 3268 32492 3372 32548
rect 3428 32492 3532 32548
rect 3588 32492 3692 32548
rect 3748 32492 3852 32548
rect 3908 32492 4012 32548
rect 4068 32492 4172 32548
rect 4228 32492 4332 32548
rect 4388 32492 4492 32548
rect 4548 32492 4652 32548
rect 4708 32492 4812 32548
rect 4868 32492 4972 32548
rect 5028 32492 5132 32548
rect 5188 32492 5292 32548
rect 5348 32492 5452 32548
rect 5508 32492 5612 32548
rect 5668 32492 5772 32548
rect 5828 32492 5932 32548
rect 5988 32492 6092 32548
rect 6148 32492 6252 32548
rect 6308 32492 6412 32548
rect 6468 32492 6572 32548
rect 6628 32492 6732 32548
rect 6788 32492 6892 32548
rect 6948 32492 7052 32548
rect 7108 32492 7212 32548
rect 7268 32492 7372 32548
rect 7428 32492 7532 32548
rect 7588 32492 7692 32548
rect 7748 32492 7852 32548
rect 7908 32492 8012 32548
rect 8068 32492 8172 32548
rect 8228 32492 8332 32548
rect 8388 32492 8972 32548
rect 9028 32492 9292 32548
rect 9348 32492 12492 32548
rect 12548 32492 12652 32548
rect 12708 32492 12812 32548
rect 12868 32492 12972 32548
rect 13028 32492 13132 32548
rect 13188 32492 13292 32548
rect 13348 32492 13452 32548
rect 13508 32492 13612 32548
rect 13668 32492 13772 32548
rect 13828 32492 13932 32548
rect 13988 32492 14092 32548
rect 14148 32492 14252 32548
rect 14308 32492 14412 32548
rect 14468 32492 14572 32548
rect 14628 32492 14732 32548
rect 14788 32492 14892 32548
rect 14948 32492 15052 32548
rect 15108 32492 15212 32548
rect 15268 32492 15372 32548
rect 15428 32492 15532 32548
rect 15588 32492 15692 32548
rect 15748 32492 15852 32548
rect 15908 32492 16012 32548
rect 16068 32492 16172 32548
rect 16228 32492 16332 32548
rect 16388 32492 16492 32548
rect 16548 32492 16652 32548
rect 16708 32492 16812 32548
rect 16868 32492 16972 32548
rect 17028 32492 17132 32548
rect 17188 32492 17292 32548
rect 17348 32492 17452 32548
rect 17508 32492 17612 32548
rect 17668 32492 17772 32548
rect 17828 32492 17932 32548
rect 17988 32492 18092 32548
rect 18148 32492 18252 32548
rect 18308 32492 18412 32548
rect 18468 32492 18572 32548
rect 18628 32492 18732 32548
rect 18788 32492 18892 32548
rect 18948 32492 19532 32548
rect 19588 32492 19852 32548
rect 19908 32492 23132 32548
rect 23188 32492 23292 32548
rect 23348 32492 23452 32548
rect 23508 32492 23612 32548
rect 23668 32492 23772 32548
rect 23828 32492 23932 32548
rect 23988 32492 24092 32548
rect 24148 32492 24252 32548
rect 24308 32492 24412 32548
rect 24468 32492 24572 32548
rect 24628 32492 24732 32548
rect 24788 32492 24892 32548
rect 24948 32492 25052 32548
rect 25108 32492 25212 32548
rect 25268 32492 25372 32548
rect 25428 32492 25532 32548
rect 25588 32492 25692 32548
rect 25748 32492 25852 32548
rect 25908 32492 26012 32548
rect 26068 32492 26172 32548
rect 26228 32492 26332 32548
rect 26388 32492 26492 32548
rect 26548 32492 26652 32548
rect 26708 32492 26812 32548
rect 26868 32492 26972 32548
rect 27028 32492 27132 32548
rect 27188 32492 27292 32548
rect 27348 32492 27452 32548
rect 27508 32492 27612 32548
rect 27668 32492 27772 32548
rect 27828 32492 27932 32548
rect 27988 32492 28092 32548
rect 28148 32492 28252 32548
rect 28308 32492 28412 32548
rect 28468 32492 28572 32548
rect 28628 32492 28732 32548
rect 28788 32492 28892 32548
rect 28948 32492 29052 32548
rect 29108 32492 29212 32548
rect 29268 32492 29372 32548
rect 29428 32492 32572 32548
rect 32628 32492 32892 32548
rect 32948 32492 33532 32548
rect 33588 32492 33692 32548
rect 33748 32492 33852 32548
rect 33908 32492 34012 32548
rect 34068 32492 34172 32548
rect 34228 32492 34332 32548
rect 34388 32492 34492 32548
rect 34548 32492 34652 32548
rect 34708 32492 34812 32548
rect 34868 32492 34972 32548
rect 35028 32492 35132 32548
rect 35188 32492 35292 32548
rect 35348 32492 35452 32548
rect 35508 32492 35612 32548
rect 35668 32492 35772 32548
rect 35828 32492 35932 32548
rect 35988 32492 36092 32548
rect 36148 32492 36252 32548
rect 36308 32492 36412 32548
rect 36468 32492 36572 32548
rect 36628 32492 36732 32548
rect 36788 32492 36892 32548
rect 36948 32492 37052 32548
rect 37108 32492 37212 32548
rect 37268 32492 37372 32548
rect 37428 32492 37532 32548
rect 37588 32492 37692 32548
rect 37748 32492 37852 32548
rect 37908 32492 38012 32548
rect 38068 32492 38172 32548
rect 38228 32492 38332 32548
rect 38388 32492 38492 32548
rect 38548 32492 38652 32548
rect 38708 32492 38812 32548
rect 38868 32492 38972 32548
rect 39028 32492 39132 32548
rect 39188 32492 39292 32548
rect 39348 32492 39452 32548
rect 39508 32492 39612 32548
rect 39668 32492 39772 32548
rect 39828 32492 39932 32548
rect 39988 32492 40092 32548
rect 40148 32492 40252 32548
rect 40308 32492 40412 32548
rect 40468 32492 40572 32548
rect 40628 32492 40732 32548
rect 40788 32492 40892 32548
rect 40948 32492 41052 32548
rect 41108 32492 41212 32548
rect 41268 32492 41372 32548
rect 41428 32492 41532 32548
rect 41588 32492 41692 32548
rect 41748 32492 41852 32548
rect 41908 32492 41920 32548
rect 0 32480 41920 32492
rect 0 32388 41920 32400
rect 0 32332 12 32388
rect 68 32332 172 32388
rect 228 32332 332 32388
rect 388 32332 492 32388
rect 548 32332 652 32388
rect 708 32332 812 32388
rect 868 32332 972 32388
rect 1028 32332 1132 32388
rect 1188 32332 1292 32388
rect 1348 32332 1452 32388
rect 1508 32332 1612 32388
rect 1668 32332 1772 32388
rect 1828 32332 1932 32388
rect 1988 32332 2092 32388
rect 2148 32332 2252 32388
rect 2308 32332 2412 32388
rect 2468 32332 2572 32388
rect 2628 32332 2732 32388
rect 2788 32332 2892 32388
rect 2948 32332 3052 32388
rect 3108 32332 3212 32388
rect 3268 32332 3372 32388
rect 3428 32332 3532 32388
rect 3588 32332 3692 32388
rect 3748 32332 3852 32388
rect 3908 32332 4012 32388
rect 4068 32332 4172 32388
rect 4228 32332 4332 32388
rect 4388 32332 4492 32388
rect 4548 32332 4652 32388
rect 4708 32332 4812 32388
rect 4868 32332 4972 32388
rect 5028 32332 5132 32388
rect 5188 32332 5292 32388
rect 5348 32332 5452 32388
rect 5508 32332 5612 32388
rect 5668 32332 5772 32388
rect 5828 32332 5932 32388
rect 5988 32332 6092 32388
rect 6148 32332 6252 32388
rect 6308 32332 6412 32388
rect 6468 32332 6572 32388
rect 6628 32332 6732 32388
rect 6788 32332 6892 32388
rect 6948 32332 7052 32388
rect 7108 32332 7212 32388
rect 7268 32332 7372 32388
rect 7428 32332 7532 32388
rect 7588 32332 7692 32388
rect 7748 32332 7852 32388
rect 7908 32332 8012 32388
rect 8068 32332 8172 32388
rect 8228 32332 8332 32388
rect 8388 32332 9452 32388
rect 9508 32332 9772 32388
rect 9828 32332 10092 32388
rect 10148 32332 10412 32388
rect 10468 32332 10732 32388
rect 10788 32332 11052 32388
rect 11108 32332 11372 32388
rect 11428 32332 12492 32388
rect 12548 32332 12652 32388
rect 12708 32332 12812 32388
rect 12868 32332 12972 32388
rect 13028 32332 13132 32388
rect 13188 32332 13292 32388
rect 13348 32332 13452 32388
rect 13508 32332 13612 32388
rect 13668 32332 13772 32388
rect 13828 32332 13932 32388
rect 13988 32332 14092 32388
rect 14148 32332 14252 32388
rect 14308 32332 14412 32388
rect 14468 32332 14572 32388
rect 14628 32332 14732 32388
rect 14788 32332 14892 32388
rect 14948 32332 15052 32388
rect 15108 32332 15212 32388
rect 15268 32332 15372 32388
rect 15428 32332 15532 32388
rect 15588 32332 15692 32388
rect 15748 32332 15852 32388
rect 15908 32332 16012 32388
rect 16068 32332 16172 32388
rect 16228 32332 16332 32388
rect 16388 32332 16492 32388
rect 16548 32332 16652 32388
rect 16708 32332 16812 32388
rect 16868 32332 16972 32388
rect 17028 32332 17132 32388
rect 17188 32332 17292 32388
rect 17348 32332 17452 32388
rect 17508 32332 17612 32388
rect 17668 32332 17772 32388
rect 17828 32332 17932 32388
rect 17988 32332 18092 32388
rect 18148 32332 18252 32388
rect 18308 32332 18412 32388
rect 18468 32332 18572 32388
rect 18628 32332 18732 32388
rect 18788 32332 18892 32388
rect 18948 32332 20012 32388
rect 20068 32332 20332 32388
rect 20388 32332 20652 32388
rect 20708 32332 20972 32388
rect 21028 32332 21292 32388
rect 21348 32332 21612 32388
rect 21668 32332 21932 32388
rect 21988 32332 23132 32388
rect 23188 32332 23292 32388
rect 23348 32332 23452 32388
rect 23508 32332 23612 32388
rect 23668 32332 23772 32388
rect 23828 32332 23932 32388
rect 23988 32332 24092 32388
rect 24148 32332 24252 32388
rect 24308 32332 24412 32388
rect 24468 32332 24572 32388
rect 24628 32332 24732 32388
rect 24788 32332 24892 32388
rect 24948 32332 25052 32388
rect 25108 32332 25212 32388
rect 25268 32332 25372 32388
rect 25428 32332 25532 32388
rect 25588 32332 25692 32388
rect 25748 32332 25852 32388
rect 25908 32332 26012 32388
rect 26068 32332 26172 32388
rect 26228 32332 26332 32388
rect 26388 32332 26492 32388
rect 26548 32332 26652 32388
rect 26708 32332 26812 32388
rect 26868 32332 26972 32388
rect 27028 32332 27132 32388
rect 27188 32332 27292 32388
rect 27348 32332 27452 32388
rect 27508 32332 27612 32388
rect 27668 32332 27772 32388
rect 27828 32332 27932 32388
rect 27988 32332 28092 32388
rect 28148 32332 28252 32388
rect 28308 32332 28412 32388
rect 28468 32332 28572 32388
rect 28628 32332 28732 32388
rect 28788 32332 28892 32388
rect 28948 32332 29052 32388
rect 29108 32332 29212 32388
rect 29268 32332 29372 32388
rect 29428 32332 30492 32388
rect 30548 32332 30812 32388
rect 30868 32332 31132 32388
rect 31188 32332 31452 32388
rect 31508 32332 31772 32388
rect 31828 32332 32092 32388
rect 32148 32332 32412 32388
rect 32468 32332 33532 32388
rect 33588 32332 33692 32388
rect 33748 32332 33852 32388
rect 33908 32332 34012 32388
rect 34068 32332 34172 32388
rect 34228 32332 34332 32388
rect 34388 32332 34492 32388
rect 34548 32332 34652 32388
rect 34708 32332 34812 32388
rect 34868 32332 34972 32388
rect 35028 32332 35132 32388
rect 35188 32332 35292 32388
rect 35348 32332 35452 32388
rect 35508 32332 35612 32388
rect 35668 32332 35772 32388
rect 35828 32332 35932 32388
rect 35988 32332 36092 32388
rect 36148 32332 36252 32388
rect 36308 32332 36412 32388
rect 36468 32332 36572 32388
rect 36628 32332 36732 32388
rect 36788 32332 36892 32388
rect 36948 32332 37052 32388
rect 37108 32332 37212 32388
rect 37268 32332 37372 32388
rect 37428 32332 37532 32388
rect 37588 32332 37692 32388
rect 37748 32332 37852 32388
rect 37908 32332 38012 32388
rect 38068 32332 38172 32388
rect 38228 32332 38332 32388
rect 38388 32332 38492 32388
rect 38548 32332 38652 32388
rect 38708 32332 38812 32388
rect 38868 32332 38972 32388
rect 39028 32332 39132 32388
rect 39188 32332 39292 32388
rect 39348 32332 39452 32388
rect 39508 32332 39612 32388
rect 39668 32332 39772 32388
rect 39828 32332 39932 32388
rect 39988 32332 40092 32388
rect 40148 32332 40252 32388
rect 40308 32332 40412 32388
rect 40468 32332 40572 32388
rect 40628 32332 40732 32388
rect 40788 32332 40892 32388
rect 40948 32332 41052 32388
rect 41108 32332 41212 32388
rect 41268 32332 41372 32388
rect 41428 32332 41532 32388
rect 41588 32332 41692 32388
rect 41748 32332 41852 32388
rect 41908 32332 41920 32388
rect 0 32320 41920 32332
rect 0 32228 41920 32240
rect 0 32172 9612 32228
rect 9668 32172 20172 32228
rect 20228 32172 32252 32228
rect 32308 32172 41920 32228
rect 0 32160 41920 32172
rect 0 32068 41920 32080
rect 0 32012 12 32068
rect 68 32012 172 32068
rect 228 32012 332 32068
rect 388 32012 492 32068
rect 548 32012 652 32068
rect 708 32012 812 32068
rect 868 32012 972 32068
rect 1028 32012 1132 32068
rect 1188 32012 1292 32068
rect 1348 32012 1452 32068
rect 1508 32012 1612 32068
rect 1668 32012 1772 32068
rect 1828 32012 1932 32068
rect 1988 32012 2092 32068
rect 2148 32012 2252 32068
rect 2308 32012 2412 32068
rect 2468 32012 2572 32068
rect 2628 32012 2732 32068
rect 2788 32012 2892 32068
rect 2948 32012 3052 32068
rect 3108 32012 3212 32068
rect 3268 32012 3372 32068
rect 3428 32012 3532 32068
rect 3588 32012 3692 32068
rect 3748 32012 3852 32068
rect 3908 32012 4012 32068
rect 4068 32012 4172 32068
rect 4228 32012 4332 32068
rect 4388 32012 4492 32068
rect 4548 32012 4652 32068
rect 4708 32012 4812 32068
rect 4868 32012 4972 32068
rect 5028 32012 5132 32068
rect 5188 32012 5292 32068
rect 5348 32012 5452 32068
rect 5508 32012 5612 32068
rect 5668 32012 5772 32068
rect 5828 32012 5932 32068
rect 5988 32012 6092 32068
rect 6148 32012 6252 32068
rect 6308 32012 6412 32068
rect 6468 32012 6572 32068
rect 6628 32012 6732 32068
rect 6788 32012 6892 32068
rect 6948 32012 7052 32068
rect 7108 32012 7212 32068
rect 7268 32012 7372 32068
rect 7428 32012 7532 32068
rect 7588 32012 7692 32068
rect 7748 32012 7852 32068
rect 7908 32012 8012 32068
rect 8068 32012 8172 32068
rect 8228 32012 8332 32068
rect 8388 32012 9452 32068
rect 9508 32012 9772 32068
rect 9828 32012 10092 32068
rect 10148 32012 10412 32068
rect 10468 32012 10732 32068
rect 10788 32012 11052 32068
rect 11108 32012 11372 32068
rect 11428 32012 12492 32068
rect 12548 32012 12652 32068
rect 12708 32012 12812 32068
rect 12868 32012 12972 32068
rect 13028 32012 13132 32068
rect 13188 32012 13292 32068
rect 13348 32012 13452 32068
rect 13508 32012 13612 32068
rect 13668 32012 13772 32068
rect 13828 32012 13932 32068
rect 13988 32012 14092 32068
rect 14148 32012 14252 32068
rect 14308 32012 14412 32068
rect 14468 32012 14572 32068
rect 14628 32012 14732 32068
rect 14788 32012 14892 32068
rect 14948 32012 15052 32068
rect 15108 32012 15212 32068
rect 15268 32012 15372 32068
rect 15428 32012 15532 32068
rect 15588 32012 15692 32068
rect 15748 32012 15852 32068
rect 15908 32012 16012 32068
rect 16068 32012 16172 32068
rect 16228 32012 16332 32068
rect 16388 32012 16492 32068
rect 16548 32012 16652 32068
rect 16708 32012 16812 32068
rect 16868 32012 16972 32068
rect 17028 32012 17132 32068
rect 17188 32012 17292 32068
rect 17348 32012 17452 32068
rect 17508 32012 17612 32068
rect 17668 32012 17772 32068
rect 17828 32012 17932 32068
rect 17988 32012 18092 32068
rect 18148 32012 18252 32068
rect 18308 32012 18412 32068
rect 18468 32012 18572 32068
rect 18628 32012 18732 32068
rect 18788 32012 18892 32068
rect 18948 32012 20012 32068
rect 20068 32012 20332 32068
rect 20388 32012 20652 32068
rect 20708 32012 20972 32068
rect 21028 32012 21292 32068
rect 21348 32012 21612 32068
rect 21668 32012 21932 32068
rect 21988 32012 23132 32068
rect 23188 32012 23292 32068
rect 23348 32012 23452 32068
rect 23508 32012 23612 32068
rect 23668 32012 23772 32068
rect 23828 32012 23932 32068
rect 23988 32012 24092 32068
rect 24148 32012 24252 32068
rect 24308 32012 24412 32068
rect 24468 32012 24572 32068
rect 24628 32012 24732 32068
rect 24788 32012 24892 32068
rect 24948 32012 25052 32068
rect 25108 32012 25212 32068
rect 25268 32012 25372 32068
rect 25428 32012 25532 32068
rect 25588 32012 25692 32068
rect 25748 32012 25852 32068
rect 25908 32012 26012 32068
rect 26068 32012 26172 32068
rect 26228 32012 26332 32068
rect 26388 32012 26492 32068
rect 26548 32012 26652 32068
rect 26708 32012 26812 32068
rect 26868 32012 26972 32068
rect 27028 32012 27132 32068
rect 27188 32012 27292 32068
rect 27348 32012 27452 32068
rect 27508 32012 27612 32068
rect 27668 32012 27772 32068
rect 27828 32012 27932 32068
rect 27988 32012 28092 32068
rect 28148 32012 28252 32068
rect 28308 32012 28412 32068
rect 28468 32012 28572 32068
rect 28628 32012 28732 32068
rect 28788 32012 28892 32068
rect 28948 32012 29052 32068
rect 29108 32012 29212 32068
rect 29268 32012 29372 32068
rect 29428 32012 30492 32068
rect 30548 32012 30812 32068
rect 30868 32012 31132 32068
rect 31188 32012 31452 32068
rect 31508 32012 31772 32068
rect 31828 32012 32092 32068
rect 32148 32012 32412 32068
rect 32468 32012 33532 32068
rect 33588 32012 33692 32068
rect 33748 32012 33852 32068
rect 33908 32012 34012 32068
rect 34068 32012 34172 32068
rect 34228 32012 34332 32068
rect 34388 32012 34492 32068
rect 34548 32012 34652 32068
rect 34708 32012 34812 32068
rect 34868 32012 34972 32068
rect 35028 32012 35132 32068
rect 35188 32012 35292 32068
rect 35348 32012 35452 32068
rect 35508 32012 35612 32068
rect 35668 32012 35772 32068
rect 35828 32012 35932 32068
rect 35988 32012 36092 32068
rect 36148 32012 36252 32068
rect 36308 32012 36412 32068
rect 36468 32012 36572 32068
rect 36628 32012 36732 32068
rect 36788 32012 36892 32068
rect 36948 32012 37052 32068
rect 37108 32012 37212 32068
rect 37268 32012 37372 32068
rect 37428 32012 37532 32068
rect 37588 32012 37692 32068
rect 37748 32012 37852 32068
rect 37908 32012 38012 32068
rect 38068 32012 38172 32068
rect 38228 32012 38332 32068
rect 38388 32012 38492 32068
rect 38548 32012 38652 32068
rect 38708 32012 38812 32068
rect 38868 32012 38972 32068
rect 39028 32012 39132 32068
rect 39188 32012 39292 32068
rect 39348 32012 39452 32068
rect 39508 32012 39612 32068
rect 39668 32012 39772 32068
rect 39828 32012 39932 32068
rect 39988 32012 40092 32068
rect 40148 32012 40252 32068
rect 40308 32012 40412 32068
rect 40468 32012 40572 32068
rect 40628 32012 40732 32068
rect 40788 32012 40892 32068
rect 40948 32012 41052 32068
rect 41108 32012 41212 32068
rect 41268 32012 41372 32068
rect 41428 32012 41532 32068
rect 41588 32012 41692 32068
rect 41748 32012 41852 32068
rect 41908 32012 41920 32068
rect 0 32000 41920 32012
rect 0 31908 41920 31920
rect 0 31852 9932 31908
rect 9988 31852 20492 31908
rect 20548 31852 31932 31908
rect 31988 31852 41920 31908
rect 0 31840 41920 31852
rect 0 31748 41920 31760
rect 0 31692 12 31748
rect 68 31692 172 31748
rect 228 31692 332 31748
rect 388 31692 492 31748
rect 548 31692 652 31748
rect 708 31692 812 31748
rect 868 31692 972 31748
rect 1028 31692 1132 31748
rect 1188 31692 1292 31748
rect 1348 31692 1452 31748
rect 1508 31692 1612 31748
rect 1668 31692 1772 31748
rect 1828 31692 1932 31748
rect 1988 31692 2092 31748
rect 2148 31692 2252 31748
rect 2308 31692 2412 31748
rect 2468 31692 2572 31748
rect 2628 31692 2732 31748
rect 2788 31692 2892 31748
rect 2948 31692 3052 31748
rect 3108 31692 3212 31748
rect 3268 31692 3372 31748
rect 3428 31692 3532 31748
rect 3588 31692 3692 31748
rect 3748 31692 3852 31748
rect 3908 31692 4012 31748
rect 4068 31692 4172 31748
rect 4228 31692 4332 31748
rect 4388 31692 4492 31748
rect 4548 31692 4652 31748
rect 4708 31692 4812 31748
rect 4868 31692 4972 31748
rect 5028 31692 5132 31748
rect 5188 31692 5292 31748
rect 5348 31692 5452 31748
rect 5508 31692 5612 31748
rect 5668 31692 5772 31748
rect 5828 31692 5932 31748
rect 5988 31692 6092 31748
rect 6148 31692 6252 31748
rect 6308 31692 6412 31748
rect 6468 31692 6572 31748
rect 6628 31692 6732 31748
rect 6788 31692 6892 31748
rect 6948 31692 7052 31748
rect 7108 31692 7212 31748
rect 7268 31692 7372 31748
rect 7428 31692 7532 31748
rect 7588 31692 7692 31748
rect 7748 31692 7852 31748
rect 7908 31692 8012 31748
rect 8068 31692 8172 31748
rect 8228 31692 8332 31748
rect 8388 31692 9452 31748
rect 9508 31692 9772 31748
rect 9828 31692 10092 31748
rect 10148 31692 10412 31748
rect 10468 31692 10732 31748
rect 10788 31692 11052 31748
rect 11108 31692 11372 31748
rect 11428 31692 12492 31748
rect 12548 31692 12652 31748
rect 12708 31692 12812 31748
rect 12868 31692 12972 31748
rect 13028 31692 13132 31748
rect 13188 31692 13292 31748
rect 13348 31692 13452 31748
rect 13508 31692 13612 31748
rect 13668 31692 13772 31748
rect 13828 31692 13932 31748
rect 13988 31692 14092 31748
rect 14148 31692 14252 31748
rect 14308 31692 14412 31748
rect 14468 31692 14572 31748
rect 14628 31692 14732 31748
rect 14788 31692 14892 31748
rect 14948 31692 15052 31748
rect 15108 31692 15212 31748
rect 15268 31692 15372 31748
rect 15428 31692 15532 31748
rect 15588 31692 15692 31748
rect 15748 31692 15852 31748
rect 15908 31692 16012 31748
rect 16068 31692 16172 31748
rect 16228 31692 16332 31748
rect 16388 31692 16492 31748
rect 16548 31692 16652 31748
rect 16708 31692 16812 31748
rect 16868 31692 16972 31748
rect 17028 31692 17132 31748
rect 17188 31692 17292 31748
rect 17348 31692 17452 31748
rect 17508 31692 17612 31748
rect 17668 31692 17772 31748
rect 17828 31692 17932 31748
rect 17988 31692 18092 31748
rect 18148 31692 18252 31748
rect 18308 31692 18412 31748
rect 18468 31692 18572 31748
rect 18628 31692 18732 31748
rect 18788 31692 18892 31748
rect 18948 31692 20012 31748
rect 20068 31692 20332 31748
rect 20388 31692 20652 31748
rect 20708 31692 20972 31748
rect 21028 31692 21292 31748
rect 21348 31692 21612 31748
rect 21668 31692 21932 31748
rect 21988 31692 23132 31748
rect 23188 31692 23292 31748
rect 23348 31692 23452 31748
rect 23508 31692 23612 31748
rect 23668 31692 23772 31748
rect 23828 31692 23932 31748
rect 23988 31692 24092 31748
rect 24148 31692 24252 31748
rect 24308 31692 24412 31748
rect 24468 31692 24572 31748
rect 24628 31692 24732 31748
rect 24788 31692 24892 31748
rect 24948 31692 25052 31748
rect 25108 31692 25212 31748
rect 25268 31692 25372 31748
rect 25428 31692 25532 31748
rect 25588 31692 25692 31748
rect 25748 31692 25852 31748
rect 25908 31692 26012 31748
rect 26068 31692 26172 31748
rect 26228 31692 26332 31748
rect 26388 31692 26492 31748
rect 26548 31692 26652 31748
rect 26708 31692 26812 31748
rect 26868 31692 26972 31748
rect 27028 31692 27132 31748
rect 27188 31692 27292 31748
rect 27348 31692 27452 31748
rect 27508 31692 27612 31748
rect 27668 31692 27772 31748
rect 27828 31692 27932 31748
rect 27988 31692 28092 31748
rect 28148 31692 28252 31748
rect 28308 31692 28412 31748
rect 28468 31692 28572 31748
rect 28628 31692 28732 31748
rect 28788 31692 28892 31748
rect 28948 31692 29052 31748
rect 29108 31692 29212 31748
rect 29268 31692 29372 31748
rect 29428 31692 30492 31748
rect 30548 31692 30812 31748
rect 30868 31692 31132 31748
rect 31188 31692 31452 31748
rect 31508 31692 31772 31748
rect 31828 31692 32092 31748
rect 32148 31692 32412 31748
rect 32468 31692 33532 31748
rect 33588 31692 33692 31748
rect 33748 31692 33852 31748
rect 33908 31692 34012 31748
rect 34068 31692 34172 31748
rect 34228 31692 34332 31748
rect 34388 31692 34492 31748
rect 34548 31692 34652 31748
rect 34708 31692 34812 31748
rect 34868 31692 34972 31748
rect 35028 31692 35132 31748
rect 35188 31692 35292 31748
rect 35348 31692 35452 31748
rect 35508 31692 35612 31748
rect 35668 31692 35772 31748
rect 35828 31692 35932 31748
rect 35988 31692 36092 31748
rect 36148 31692 36252 31748
rect 36308 31692 36412 31748
rect 36468 31692 36572 31748
rect 36628 31692 36732 31748
rect 36788 31692 36892 31748
rect 36948 31692 37052 31748
rect 37108 31692 37212 31748
rect 37268 31692 37372 31748
rect 37428 31692 37532 31748
rect 37588 31692 37692 31748
rect 37748 31692 37852 31748
rect 37908 31692 38012 31748
rect 38068 31692 38172 31748
rect 38228 31692 38332 31748
rect 38388 31692 38492 31748
rect 38548 31692 38652 31748
rect 38708 31692 38812 31748
rect 38868 31692 38972 31748
rect 39028 31692 39132 31748
rect 39188 31692 39292 31748
rect 39348 31692 39452 31748
rect 39508 31692 39612 31748
rect 39668 31692 39772 31748
rect 39828 31692 39932 31748
rect 39988 31692 40092 31748
rect 40148 31692 40252 31748
rect 40308 31692 40412 31748
rect 40468 31692 40572 31748
rect 40628 31692 40732 31748
rect 40788 31692 40892 31748
rect 40948 31692 41052 31748
rect 41108 31692 41212 31748
rect 41268 31692 41372 31748
rect 41428 31692 41532 31748
rect 41588 31692 41692 31748
rect 41748 31692 41852 31748
rect 41908 31692 41920 31748
rect 0 31680 41920 31692
rect 0 31588 41920 31600
rect 0 31532 10252 31588
rect 10308 31532 20812 31588
rect 20868 31532 31612 31588
rect 31668 31532 41920 31588
rect 0 31520 41920 31532
rect 0 31428 41920 31440
rect 0 31372 12 31428
rect 68 31372 172 31428
rect 228 31372 332 31428
rect 388 31372 492 31428
rect 548 31372 652 31428
rect 708 31372 812 31428
rect 868 31372 972 31428
rect 1028 31372 1132 31428
rect 1188 31372 1292 31428
rect 1348 31372 1452 31428
rect 1508 31372 1612 31428
rect 1668 31372 1772 31428
rect 1828 31372 1932 31428
rect 1988 31372 2092 31428
rect 2148 31372 2252 31428
rect 2308 31372 2412 31428
rect 2468 31372 2572 31428
rect 2628 31372 2732 31428
rect 2788 31372 2892 31428
rect 2948 31372 3052 31428
rect 3108 31372 3212 31428
rect 3268 31372 3372 31428
rect 3428 31372 3532 31428
rect 3588 31372 3692 31428
rect 3748 31372 3852 31428
rect 3908 31372 4012 31428
rect 4068 31372 4172 31428
rect 4228 31372 4332 31428
rect 4388 31372 4492 31428
rect 4548 31372 4652 31428
rect 4708 31372 4812 31428
rect 4868 31372 4972 31428
rect 5028 31372 5132 31428
rect 5188 31372 5292 31428
rect 5348 31372 5452 31428
rect 5508 31372 5612 31428
rect 5668 31372 5772 31428
rect 5828 31372 5932 31428
rect 5988 31372 6092 31428
rect 6148 31372 6252 31428
rect 6308 31372 6412 31428
rect 6468 31372 6572 31428
rect 6628 31372 6732 31428
rect 6788 31372 6892 31428
rect 6948 31372 7052 31428
rect 7108 31372 7212 31428
rect 7268 31372 7372 31428
rect 7428 31372 7532 31428
rect 7588 31372 7692 31428
rect 7748 31372 7852 31428
rect 7908 31372 8012 31428
rect 8068 31372 8172 31428
rect 8228 31372 8332 31428
rect 8388 31372 9452 31428
rect 9508 31372 9772 31428
rect 9828 31372 10092 31428
rect 10148 31372 10412 31428
rect 10468 31372 10732 31428
rect 10788 31372 11052 31428
rect 11108 31372 11372 31428
rect 11428 31372 12492 31428
rect 12548 31372 12652 31428
rect 12708 31372 12812 31428
rect 12868 31372 12972 31428
rect 13028 31372 13132 31428
rect 13188 31372 13292 31428
rect 13348 31372 13452 31428
rect 13508 31372 13612 31428
rect 13668 31372 13772 31428
rect 13828 31372 13932 31428
rect 13988 31372 14092 31428
rect 14148 31372 14252 31428
rect 14308 31372 14412 31428
rect 14468 31372 14572 31428
rect 14628 31372 14732 31428
rect 14788 31372 14892 31428
rect 14948 31372 15052 31428
rect 15108 31372 15212 31428
rect 15268 31372 15372 31428
rect 15428 31372 15532 31428
rect 15588 31372 15692 31428
rect 15748 31372 15852 31428
rect 15908 31372 16012 31428
rect 16068 31372 16172 31428
rect 16228 31372 16332 31428
rect 16388 31372 16492 31428
rect 16548 31372 16652 31428
rect 16708 31372 16812 31428
rect 16868 31372 16972 31428
rect 17028 31372 17132 31428
rect 17188 31372 17292 31428
rect 17348 31372 17452 31428
rect 17508 31372 17612 31428
rect 17668 31372 17772 31428
rect 17828 31372 17932 31428
rect 17988 31372 18092 31428
rect 18148 31372 18252 31428
rect 18308 31372 18412 31428
rect 18468 31372 18572 31428
rect 18628 31372 18732 31428
rect 18788 31372 18892 31428
rect 18948 31372 20012 31428
rect 20068 31372 20332 31428
rect 20388 31372 20652 31428
rect 20708 31372 20972 31428
rect 21028 31372 21292 31428
rect 21348 31372 21612 31428
rect 21668 31372 21932 31428
rect 21988 31372 23132 31428
rect 23188 31372 23292 31428
rect 23348 31372 23452 31428
rect 23508 31372 23612 31428
rect 23668 31372 23772 31428
rect 23828 31372 23932 31428
rect 23988 31372 24092 31428
rect 24148 31372 24252 31428
rect 24308 31372 24412 31428
rect 24468 31372 24572 31428
rect 24628 31372 24732 31428
rect 24788 31372 24892 31428
rect 24948 31372 25052 31428
rect 25108 31372 25212 31428
rect 25268 31372 25372 31428
rect 25428 31372 25532 31428
rect 25588 31372 25692 31428
rect 25748 31372 25852 31428
rect 25908 31372 26012 31428
rect 26068 31372 26172 31428
rect 26228 31372 26332 31428
rect 26388 31372 26492 31428
rect 26548 31372 26652 31428
rect 26708 31372 26812 31428
rect 26868 31372 26972 31428
rect 27028 31372 27132 31428
rect 27188 31372 27292 31428
rect 27348 31372 27452 31428
rect 27508 31372 27612 31428
rect 27668 31372 27772 31428
rect 27828 31372 27932 31428
rect 27988 31372 28092 31428
rect 28148 31372 28252 31428
rect 28308 31372 28412 31428
rect 28468 31372 28572 31428
rect 28628 31372 28732 31428
rect 28788 31372 28892 31428
rect 28948 31372 29052 31428
rect 29108 31372 29212 31428
rect 29268 31372 29372 31428
rect 29428 31372 30492 31428
rect 30548 31372 30812 31428
rect 30868 31372 31132 31428
rect 31188 31372 31452 31428
rect 31508 31372 31772 31428
rect 31828 31372 32092 31428
rect 32148 31372 32412 31428
rect 32468 31372 33532 31428
rect 33588 31372 33692 31428
rect 33748 31372 33852 31428
rect 33908 31372 34012 31428
rect 34068 31372 34172 31428
rect 34228 31372 34332 31428
rect 34388 31372 34492 31428
rect 34548 31372 34652 31428
rect 34708 31372 34812 31428
rect 34868 31372 34972 31428
rect 35028 31372 35132 31428
rect 35188 31372 35292 31428
rect 35348 31372 35452 31428
rect 35508 31372 35612 31428
rect 35668 31372 35772 31428
rect 35828 31372 35932 31428
rect 35988 31372 36092 31428
rect 36148 31372 36252 31428
rect 36308 31372 36412 31428
rect 36468 31372 36572 31428
rect 36628 31372 36732 31428
rect 36788 31372 36892 31428
rect 36948 31372 37052 31428
rect 37108 31372 37212 31428
rect 37268 31372 37372 31428
rect 37428 31372 37532 31428
rect 37588 31372 37692 31428
rect 37748 31372 37852 31428
rect 37908 31372 38012 31428
rect 38068 31372 38172 31428
rect 38228 31372 38332 31428
rect 38388 31372 38492 31428
rect 38548 31372 38652 31428
rect 38708 31372 38812 31428
rect 38868 31372 38972 31428
rect 39028 31372 39132 31428
rect 39188 31372 39292 31428
rect 39348 31372 39452 31428
rect 39508 31372 39612 31428
rect 39668 31372 39772 31428
rect 39828 31372 39932 31428
rect 39988 31372 40092 31428
rect 40148 31372 40252 31428
rect 40308 31372 40412 31428
rect 40468 31372 40572 31428
rect 40628 31372 40732 31428
rect 40788 31372 40892 31428
rect 40948 31372 41052 31428
rect 41108 31372 41212 31428
rect 41268 31372 41372 31428
rect 41428 31372 41532 31428
rect 41588 31372 41692 31428
rect 41748 31372 41852 31428
rect 41908 31372 41920 31428
rect 0 31360 41920 31372
rect 0 31268 41920 31280
rect 0 31212 10572 31268
rect 10628 31212 21132 31268
rect 21188 31212 31292 31268
rect 31348 31212 41920 31268
rect 0 31200 41920 31212
rect 0 31108 41920 31120
rect 0 31052 12 31108
rect 68 31052 172 31108
rect 228 31052 332 31108
rect 388 31052 492 31108
rect 548 31052 652 31108
rect 708 31052 812 31108
rect 868 31052 972 31108
rect 1028 31052 1132 31108
rect 1188 31052 1292 31108
rect 1348 31052 1452 31108
rect 1508 31052 1612 31108
rect 1668 31052 1772 31108
rect 1828 31052 1932 31108
rect 1988 31052 2092 31108
rect 2148 31052 2252 31108
rect 2308 31052 2412 31108
rect 2468 31052 2572 31108
rect 2628 31052 2732 31108
rect 2788 31052 2892 31108
rect 2948 31052 3052 31108
rect 3108 31052 3212 31108
rect 3268 31052 3372 31108
rect 3428 31052 3532 31108
rect 3588 31052 3692 31108
rect 3748 31052 3852 31108
rect 3908 31052 4012 31108
rect 4068 31052 4172 31108
rect 4228 31052 4332 31108
rect 4388 31052 4492 31108
rect 4548 31052 4652 31108
rect 4708 31052 4812 31108
rect 4868 31052 4972 31108
rect 5028 31052 5132 31108
rect 5188 31052 5292 31108
rect 5348 31052 5452 31108
rect 5508 31052 5612 31108
rect 5668 31052 5772 31108
rect 5828 31052 5932 31108
rect 5988 31052 6092 31108
rect 6148 31052 6252 31108
rect 6308 31052 6412 31108
rect 6468 31052 6572 31108
rect 6628 31052 6732 31108
rect 6788 31052 6892 31108
rect 6948 31052 7052 31108
rect 7108 31052 7212 31108
rect 7268 31052 7372 31108
rect 7428 31052 7532 31108
rect 7588 31052 7692 31108
rect 7748 31052 7852 31108
rect 7908 31052 8012 31108
rect 8068 31052 8172 31108
rect 8228 31052 8332 31108
rect 8388 31052 9452 31108
rect 9508 31052 9772 31108
rect 9828 31052 10092 31108
rect 10148 31052 10412 31108
rect 10468 31052 10732 31108
rect 10788 31052 11052 31108
rect 11108 31052 11372 31108
rect 11428 31052 12492 31108
rect 12548 31052 12652 31108
rect 12708 31052 12812 31108
rect 12868 31052 12972 31108
rect 13028 31052 13132 31108
rect 13188 31052 13292 31108
rect 13348 31052 13452 31108
rect 13508 31052 13612 31108
rect 13668 31052 13772 31108
rect 13828 31052 13932 31108
rect 13988 31052 14092 31108
rect 14148 31052 14252 31108
rect 14308 31052 14412 31108
rect 14468 31052 14572 31108
rect 14628 31052 14732 31108
rect 14788 31052 14892 31108
rect 14948 31052 15052 31108
rect 15108 31052 15212 31108
rect 15268 31052 15372 31108
rect 15428 31052 15532 31108
rect 15588 31052 15692 31108
rect 15748 31052 15852 31108
rect 15908 31052 16012 31108
rect 16068 31052 16172 31108
rect 16228 31052 16332 31108
rect 16388 31052 16492 31108
rect 16548 31052 16652 31108
rect 16708 31052 16812 31108
rect 16868 31052 16972 31108
rect 17028 31052 17132 31108
rect 17188 31052 17292 31108
rect 17348 31052 17452 31108
rect 17508 31052 17612 31108
rect 17668 31052 17772 31108
rect 17828 31052 17932 31108
rect 17988 31052 18092 31108
rect 18148 31052 18252 31108
rect 18308 31052 18412 31108
rect 18468 31052 18572 31108
rect 18628 31052 18732 31108
rect 18788 31052 18892 31108
rect 18948 31052 20012 31108
rect 20068 31052 20332 31108
rect 20388 31052 20652 31108
rect 20708 31052 20972 31108
rect 21028 31052 21292 31108
rect 21348 31052 21612 31108
rect 21668 31052 21932 31108
rect 21988 31052 23132 31108
rect 23188 31052 23292 31108
rect 23348 31052 23452 31108
rect 23508 31052 23612 31108
rect 23668 31052 23772 31108
rect 23828 31052 23932 31108
rect 23988 31052 24092 31108
rect 24148 31052 24252 31108
rect 24308 31052 24412 31108
rect 24468 31052 24572 31108
rect 24628 31052 24732 31108
rect 24788 31052 24892 31108
rect 24948 31052 25052 31108
rect 25108 31052 25212 31108
rect 25268 31052 25372 31108
rect 25428 31052 25532 31108
rect 25588 31052 25692 31108
rect 25748 31052 25852 31108
rect 25908 31052 26012 31108
rect 26068 31052 26172 31108
rect 26228 31052 26332 31108
rect 26388 31052 26492 31108
rect 26548 31052 26652 31108
rect 26708 31052 26812 31108
rect 26868 31052 26972 31108
rect 27028 31052 27132 31108
rect 27188 31052 27292 31108
rect 27348 31052 27452 31108
rect 27508 31052 27612 31108
rect 27668 31052 27772 31108
rect 27828 31052 27932 31108
rect 27988 31052 28092 31108
rect 28148 31052 28252 31108
rect 28308 31052 28412 31108
rect 28468 31052 28572 31108
rect 28628 31052 28732 31108
rect 28788 31052 28892 31108
rect 28948 31052 29052 31108
rect 29108 31052 29212 31108
rect 29268 31052 29372 31108
rect 29428 31052 30492 31108
rect 30548 31052 30812 31108
rect 30868 31052 31132 31108
rect 31188 31052 31452 31108
rect 31508 31052 31772 31108
rect 31828 31052 32092 31108
rect 32148 31052 32412 31108
rect 32468 31052 33532 31108
rect 33588 31052 33692 31108
rect 33748 31052 33852 31108
rect 33908 31052 34012 31108
rect 34068 31052 34172 31108
rect 34228 31052 34332 31108
rect 34388 31052 34492 31108
rect 34548 31052 34652 31108
rect 34708 31052 34812 31108
rect 34868 31052 34972 31108
rect 35028 31052 35132 31108
rect 35188 31052 35292 31108
rect 35348 31052 35452 31108
rect 35508 31052 35612 31108
rect 35668 31052 35772 31108
rect 35828 31052 35932 31108
rect 35988 31052 36092 31108
rect 36148 31052 36252 31108
rect 36308 31052 36412 31108
rect 36468 31052 36572 31108
rect 36628 31052 36732 31108
rect 36788 31052 36892 31108
rect 36948 31052 37052 31108
rect 37108 31052 37212 31108
rect 37268 31052 37372 31108
rect 37428 31052 37532 31108
rect 37588 31052 37692 31108
rect 37748 31052 37852 31108
rect 37908 31052 38012 31108
rect 38068 31052 38172 31108
rect 38228 31052 38332 31108
rect 38388 31052 38492 31108
rect 38548 31052 38652 31108
rect 38708 31052 38812 31108
rect 38868 31052 38972 31108
rect 39028 31052 39132 31108
rect 39188 31052 39292 31108
rect 39348 31052 39452 31108
rect 39508 31052 39612 31108
rect 39668 31052 39772 31108
rect 39828 31052 39932 31108
rect 39988 31052 40092 31108
rect 40148 31052 40252 31108
rect 40308 31052 40412 31108
rect 40468 31052 40572 31108
rect 40628 31052 40732 31108
rect 40788 31052 40892 31108
rect 40948 31052 41052 31108
rect 41108 31052 41212 31108
rect 41268 31052 41372 31108
rect 41428 31052 41532 31108
rect 41588 31052 41692 31108
rect 41748 31052 41852 31108
rect 41908 31052 41920 31108
rect 0 31040 41920 31052
rect 0 30948 41920 30960
rect 0 30892 10892 30948
rect 10948 30892 21452 30948
rect 21508 30892 30972 30948
rect 31028 30892 41920 30948
rect 0 30880 41920 30892
rect 0 30788 41920 30800
rect 0 30732 12 30788
rect 68 30732 172 30788
rect 228 30732 332 30788
rect 388 30732 492 30788
rect 548 30732 652 30788
rect 708 30732 812 30788
rect 868 30732 972 30788
rect 1028 30732 1132 30788
rect 1188 30732 1292 30788
rect 1348 30732 1452 30788
rect 1508 30732 1612 30788
rect 1668 30732 1772 30788
rect 1828 30732 1932 30788
rect 1988 30732 2092 30788
rect 2148 30732 2252 30788
rect 2308 30732 2412 30788
rect 2468 30732 2572 30788
rect 2628 30732 2732 30788
rect 2788 30732 2892 30788
rect 2948 30732 3052 30788
rect 3108 30732 3212 30788
rect 3268 30732 3372 30788
rect 3428 30732 3532 30788
rect 3588 30732 3692 30788
rect 3748 30732 3852 30788
rect 3908 30732 4012 30788
rect 4068 30732 4172 30788
rect 4228 30732 4332 30788
rect 4388 30732 4492 30788
rect 4548 30732 4652 30788
rect 4708 30732 4812 30788
rect 4868 30732 4972 30788
rect 5028 30732 5132 30788
rect 5188 30732 5292 30788
rect 5348 30732 5452 30788
rect 5508 30732 5612 30788
rect 5668 30732 5772 30788
rect 5828 30732 5932 30788
rect 5988 30732 6092 30788
rect 6148 30732 6252 30788
rect 6308 30732 6412 30788
rect 6468 30732 6572 30788
rect 6628 30732 6732 30788
rect 6788 30732 6892 30788
rect 6948 30732 7052 30788
rect 7108 30732 7212 30788
rect 7268 30732 7372 30788
rect 7428 30732 7532 30788
rect 7588 30732 7692 30788
rect 7748 30732 7852 30788
rect 7908 30732 8012 30788
rect 8068 30732 8172 30788
rect 8228 30732 8332 30788
rect 8388 30732 9452 30788
rect 9508 30732 9772 30788
rect 9828 30732 10092 30788
rect 10148 30732 10412 30788
rect 10468 30732 10732 30788
rect 10788 30732 11052 30788
rect 11108 30732 11372 30788
rect 11428 30732 12492 30788
rect 12548 30732 12652 30788
rect 12708 30732 12812 30788
rect 12868 30732 12972 30788
rect 13028 30732 13132 30788
rect 13188 30732 13292 30788
rect 13348 30732 13452 30788
rect 13508 30732 13612 30788
rect 13668 30732 13772 30788
rect 13828 30732 13932 30788
rect 13988 30732 14092 30788
rect 14148 30732 14252 30788
rect 14308 30732 14412 30788
rect 14468 30732 14572 30788
rect 14628 30732 14732 30788
rect 14788 30732 14892 30788
rect 14948 30732 15052 30788
rect 15108 30732 15212 30788
rect 15268 30732 15372 30788
rect 15428 30732 15532 30788
rect 15588 30732 15692 30788
rect 15748 30732 15852 30788
rect 15908 30732 16012 30788
rect 16068 30732 16172 30788
rect 16228 30732 16332 30788
rect 16388 30732 16492 30788
rect 16548 30732 16652 30788
rect 16708 30732 16812 30788
rect 16868 30732 16972 30788
rect 17028 30732 17132 30788
rect 17188 30732 17292 30788
rect 17348 30732 17452 30788
rect 17508 30732 17612 30788
rect 17668 30732 17772 30788
rect 17828 30732 17932 30788
rect 17988 30732 18092 30788
rect 18148 30732 18252 30788
rect 18308 30732 18412 30788
rect 18468 30732 18572 30788
rect 18628 30732 18732 30788
rect 18788 30732 18892 30788
rect 18948 30732 20012 30788
rect 20068 30732 20332 30788
rect 20388 30732 20652 30788
rect 20708 30732 20972 30788
rect 21028 30732 21292 30788
rect 21348 30732 21612 30788
rect 21668 30732 21932 30788
rect 21988 30732 23132 30788
rect 23188 30732 23292 30788
rect 23348 30732 23452 30788
rect 23508 30732 23612 30788
rect 23668 30732 23772 30788
rect 23828 30732 23932 30788
rect 23988 30732 24092 30788
rect 24148 30732 24252 30788
rect 24308 30732 24412 30788
rect 24468 30732 24572 30788
rect 24628 30732 24732 30788
rect 24788 30732 24892 30788
rect 24948 30732 25052 30788
rect 25108 30732 25212 30788
rect 25268 30732 25372 30788
rect 25428 30732 25532 30788
rect 25588 30732 25692 30788
rect 25748 30732 25852 30788
rect 25908 30732 26012 30788
rect 26068 30732 26172 30788
rect 26228 30732 26332 30788
rect 26388 30732 26492 30788
rect 26548 30732 26652 30788
rect 26708 30732 26812 30788
rect 26868 30732 26972 30788
rect 27028 30732 27132 30788
rect 27188 30732 27292 30788
rect 27348 30732 27452 30788
rect 27508 30732 27612 30788
rect 27668 30732 27772 30788
rect 27828 30732 27932 30788
rect 27988 30732 28092 30788
rect 28148 30732 28252 30788
rect 28308 30732 28412 30788
rect 28468 30732 28572 30788
rect 28628 30732 28732 30788
rect 28788 30732 28892 30788
rect 28948 30732 29052 30788
rect 29108 30732 29212 30788
rect 29268 30732 29372 30788
rect 29428 30732 30492 30788
rect 30548 30732 30812 30788
rect 30868 30732 31132 30788
rect 31188 30732 31452 30788
rect 31508 30732 31772 30788
rect 31828 30732 32092 30788
rect 32148 30732 32412 30788
rect 32468 30732 33532 30788
rect 33588 30732 33692 30788
rect 33748 30732 33852 30788
rect 33908 30732 34012 30788
rect 34068 30732 34172 30788
rect 34228 30732 34332 30788
rect 34388 30732 34492 30788
rect 34548 30732 34652 30788
rect 34708 30732 34812 30788
rect 34868 30732 34972 30788
rect 35028 30732 35132 30788
rect 35188 30732 35292 30788
rect 35348 30732 35452 30788
rect 35508 30732 35612 30788
rect 35668 30732 35772 30788
rect 35828 30732 35932 30788
rect 35988 30732 36092 30788
rect 36148 30732 36252 30788
rect 36308 30732 36412 30788
rect 36468 30732 36572 30788
rect 36628 30732 36732 30788
rect 36788 30732 36892 30788
rect 36948 30732 37052 30788
rect 37108 30732 37212 30788
rect 37268 30732 37372 30788
rect 37428 30732 37532 30788
rect 37588 30732 37692 30788
rect 37748 30732 37852 30788
rect 37908 30732 38012 30788
rect 38068 30732 38172 30788
rect 38228 30732 38332 30788
rect 38388 30732 38492 30788
rect 38548 30732 38652 30788
rect 38708 30732 38812 30788
rect 38868 30732 38972 30788
rect 39028 30732 39132 30788
rect 39188 30732 39292 30788
rect 39348 30732 39452 30788
rect 39508 30732 39612 30788
rect 39668 30732 39772 30788
rect 39828 30732 39932 30788
rect 39988 30732 40092 30788
rect 40148 30732 40252 30788
rect 40308 30732 40412 30788
rect 40468 30732 40572 30788
rect 40628 30732 40732 30788
rect 40788 30732 40892 30788
rect 40948 30732 41052 30788
rect 41108 30732 41212 30788
rect 41268 30732 41372 30788
rect 41428 30732 41532 30788
rect 41588 30732 41692 30788
rect 41748 30732 41852 30788
rect 41908 30732 41920 30788
rect 0 30720 41920 30732
rect 0 30628 41920 30640
rect 0 30572 11212 30628
rect 11268 30572 21772 30628
rect 21828 30572 30652 30628
rect 30708 30572 41920 30628
rect 0 30560 41920 30572
rect 0 30468 41920 30480
rect 0 30412 12 30468
rect 68 30412 172 30468
rect 228 30412 332 30468
rect 388 30412 492 30468
rect 548 30412 652 30468
rect 708 30412 812 30468
rect 868 30412 972 30468
rect 1028 30412 1132 30468
rect 1188 30412 1292 30468
rect 1348 30412 1452 30468
rect 1508 30412 1612 30468
rect 1668 30412 1772 30468
rect 1828 30412 1932 30468
rect 1988 30412 2092 30468
rect 2148 30412 2252 30468
rect 2308 30412 2412 30468
rect 2468 30412 2572 30468
rect 2628 30412 2732 30468
rect 2788 30412 2892 30468
rect 2948 30412 3052 30468
rect 3108 30412 3212 30468
rect 3268 30412 3372 30468
rect 3428 30412 3532 30468
rect 3588 30412 3692 30468
rect 3748 30412 3852 30468
rect 3908 30412 4012 30468
rect 4068 30412 4172 30468
rect 4228 30412 4332 30468
rect 4388 30412 4492 30468
rect 4548 30412 4652 30468
rect 4708 30412 4812 30468
rect 4868 30412 4972 30468
rect 5028 30412 5132 30468
rect 5188 30412 5292 30468
rect 5348 30412 5452 30468
rect 5508 30412 5612 30468
rect 5668 30412 5772 30468
rect 5828 30412 5932 30468
rect 5988 30412 6092 30468
rect 6148 30412 6252 30468
rect 6308 30412 6412 30468
rect 6468 30412 6572 30468
rect 6628 30412 6732 30468
rect 6788 30412 6892 30468
rect 6948 30412 7052 30468
rect 7108 30412 7212 30468
rect 7268 30412 7372 30468
rect 7428 30412 7532 30468
rect 7588 30412 7692 30468
rect 7748 30412 7852 30468
rect 7908 30412 8012 30468
rect 8068 30412 8172 30468
rect 8228 30412 8332 30468
rect 8388 30412 9452 30468
rect 9508 30412 9772 30468
rect 9828 30412 10092 30468
rect 10148 30412 10412 30468
rect 10468 30412 10732 30468
rect 10788 30412 11052 30468
rect 11108 30412 11372 30468
rect 11428 30412 12492 30468
rect 12548 30412 12652 30468
rect 12708 30412 12812 30468
rect 12868 30412 12972 30468
rect 13028 30412 13132 30468
rect 13188 30412 13292 30468
rect 13348 30412 13452 30468
rect 13508 30412 13612 30468
rect 13668 30412 13772 30468
rect 13828 30412 13932 30468
rect 13988 30412 14092 30468
rect 14148 30412 14252 30468
rect 14308 30412 14412 30468
rect 14468 30412 14572 30468
rect 14628 30412 14732 30468
rect 14788 30412 14892 30468
rect 14948 30412 15052 30468
rect 15108 30412 15212 30468
rect 15268 30412 15372 30468
rect 15428 30412 15532 30468
rect 15588 30412 15692 30468
rect 15748 30412 15852 30468
rect 15908 30412 16012 30468
rect 16068 30412 16172 30468
rect 16228 30412 16332 30468
rect 16388 30412 16492 30468
rect 16548 30412 16652 30468
rect 16708 30412 16812 30468
rect 16868 30412 16972 30468
rect 17028 30412 17132 30468
rect 17188 30412 17292 30468
rect 17348 30412 17452 30468
rect 17508 30412 17612 30468
rect 17668 30412 17772 30468
rect 17828 30412 17932 30468
rect 17988 30412 18092 30468
rect 18148 30412 18252 30468
rect 18308 30412 18412 30468
rect 18468 30412 18572 30468
rect 18628 30412 18732 30468
rect 18788 30412 18892 30468
rect 18948 30412 20012 30468
rect 20068 30412 20332 30468
rect 20388 30412 20652 30468
rect 20708 30412 20972 30468
rect 21028 30412 21292 30468
rect 21348 30412 21612 30468
rect 21668 30412 21932 30468
rect 21988 30412 23132 30468
rect 23188 30412 23292 30468
rect 23348 30412 23452 30468
rect 23508 30412 23612 30468
rect 23668 30412 23772 30468
rect 23828 30412 23932 30468
rect 23988 30412 24092 30468
rect 24148 30412 24252 30468
rect 24308 30412 24412 30468
rect 24468 30412 24572 30468
rect 24628 30412 24732 30468
rect 24788 30412 24892 30468
rect 24948 30412 25052 30468
rect 25108 30412 25212 30468
rect 25268 30412 25372 30468
rect 25428 30412 25532 30468
rect 25588 30412 25692 30468
rect 25748 30412 25852 30468
rect 25908 30412 26012 30468
rect 26068 30412 26172 30468
rect 26228 30412 26332 30468
rect 26388 30412 26492 30468
rect 26548 30412 26652 30468
rect 26708 30412 26812 30468
rect 26868 30412 26972 30468
rect 27028 30412 27132 30468
rect 27188 30412 27292 30468
rect 27348 30412 27452 30468
rect 27508 30412 27612 30468
rect 27668 30412 27772 30468
rect 27828 30412 27932 30468
rect 27988 30412 28092 30468
rect 28148 30412 28252 30468
rect 28308 30412 28412 30468
rect 28468 30412 28572 30468
rect 28628 30412 28732 30468
rect 28788 30412 28892 30468
rect 28948 30412 29052 30468
rect 29108 30412 29212 30468
rect 29268 30412 29372 30468
rect 29428 30412 30492 30468
rect 30548 30412 30812 30468
rect 30868 30412 31132 30468
rect 31188 30412 31452 30468
rect 31508 30412 31772 30468
rect 31828 30412 32092 30468
rect 32148 30412 32412 30468
rect 32468 30412 33532 30468
rect 33588 30412 33692 30468
rect 33748 30412 33852 30468
rect 33908 30412 34012 30468
rect 34068 30412 34172 30468
rect 34228 30412 34332 30468
rect 34388 30412 34492 30468
rect 34548 30412 34652 30468
rect 34708 30412 34812 30468
rect 34868 30412 34972 30468
rect 35028 30412 35132 30468
rect 35188 30412 35292 30468
rect 35348 30412 35452 30468
rect 35508 30412 35612 30468
rect 35668 30412 35772 30468
rect 35828 30412 35932 30468
rect 35988 30412 36092 30468
rect 36148 30412 36252 30468
rect 36308 30412 36412 30468
rect 36468 30412 36572 30468
rect 36628 30412 36732 30468
rect 36788 30412 36892 30468
rect 36948 30412 37052 30468
rect 37108 30412 37212 30468
rect 37268 30412 37372 30468
rect 37428 30412 37532 30468
rect 37588 30412 37692 30468
rect 37748 30412 37852 30468
rect 37908 30412 38012 30468
rect 38068 30412 38172 30468
rect 38228 30412 38332 30468
rect 38388 30412 38492 30468
rect 38548 30412 38652 30468
rect 38708 30412 38812 30468
rect 38868 30412 38972 30468
rect 39028 30412 39132 30468
rect 39188 30412 39292 30468
rect 39348 30412 39452 30468
rect 39508 30412 39612 30468
rect 39668 30412 39772 30468
rect 39828 30412 39932 30468
rect 39988 30412 40092 30468
rect 40148 30412 40252 30468
rect 40308 30412 40412 30468
rect 40468 30412 40572 30468
rect 40628 30412 40732 30468
rect 40788 30412 40892 30468
rect 40948 30412 41052 30468
rect 41108 30412 41212 30468
rect 41268 30412 41372 30468
rect 41428 30412 41532 30468
rect 41588 30412 41692 30468
rect 41748 30412 41852 30468
rect 41908 30412 41920 30468
rect 0 30400 41920 30412
rect 0 30308 41920 30320
rect 0 30252 12 30308
rect 68 30252 172 30308
rect 228 30252 332 30308
rect 388 30252 492 30308
rect 548 30252 652 30308
rect 708 30252 812 30308
rect 868 30252 972 30308
rect 1028 30252 1132 30308
rect 1188 30252 1292 30308
rect 1348 30252 1452 30308
rect 1508 30252 1612 30308
rect 1668 30252 1772 30308
rect 1828 30252 1932 30308
rect 1988 30252 2092 30308
rect 2148 30252 2252 30308
rect 2308 30252 2412 30308
rect 2468 30252 2572 30308
rect 2628 30252 2732 30308
rect 2788 30252 2892 30308
rect 2948 30252 3052 30308
rect 3108 30252 3212 30308
rect 3268 30252 3372 30308
rect 3428 30252 3532 30308
rect 3588 30252 3692 30308
rect 3748 30252 3852 30308
rect 3908 30252 4012 30308
rect 4068 30252 4172 30308
rect 4228 30252 4332 30308
rect 4388 30252 4492 30308
rect 4548 30252 4652 30308
rect 4708 30252 4812 30308
rect 4868 30252 4972 30308
rect 5028 30252 5132 30308
rect 5188 30252 5292 30308
rect 5348 30252 5452 30308
rect 5508 30252 5612 30308
rect 5668 30252 5772 30308
rect 5828 30252 5932 30308
rect 5988 30252 6092 30308
rect 6148 30252 6252 30308
rect 6308 30252 6412 30308
rect 6468 30252 6572 30308
rect 6628 30252 6732 30308
rect 6788 30252 6892 30308
rect 6948 30252 7052 30308
rect 7108 30252 7212 30308
rect 7268 30252 7372 30308
rect 7428 30252 7532 30308
rect 7588 30252 7692 30308
rect 7748 30252 7852 30308
rect 7908 30252 8012 30308
rect 8068 30252 8172 30308
rect 8228 30252 8332 30308
rect 8388 30252 11532 30308
rect 11588 30252 11852 30308
rect 11908 30252 12492 30308
rect 12548 30252 12652 30308
rect 12708 30252 12812 30308
rect 12868 30252 12972 30308
rect 13028 30252 13132 30308
rect 13188 30252 13292 30308
rect 13348 30252 13452 30308
rect 13508 30252 13612 30308
rect 13668 30252 13772 30308
rect 13828 30252 13932 30308
rect 13988 30252 14092 30308
rect 14148 30252 14252 30308
rect 14308 30252 14412 30308
rect 14468 30252 14572 30308
rect 14628 30252 14732 30308
rect 14788 30252 14892 30308
rect 14948 30252 15052 30308
rect 15108 30252 15212 30308
rect 15268 30252 15372 30308
rect 15428 30252 15532 30308
rect 15588 30252 15692 30308
rect 15748 30252 15852 30308
rect 15908 30252 16012 30308
rect 16068 30252 16172 30308
rect 16228 30252 16332 30308
rect 16388 30252 16492 30308
rect 16548 30252 16652 30308
rect 16708 30252 16812 30308
rect 16868 30252 16972 30308
rect 17028 30252 17132 30308
rect 17188 30252 17292 30308
rect 17348 30252 17452 30308
rect 17508 30252 17612 30308
rect 17668 30252 17772 30308
rect 17828 30252 17932 30308
rect 17988 30252 18092 30308
rect 18148 30252 18252 30308
rect 18308 30252 18412 30308
rect 18468 30252 18572 30308
rect 18628 30252 18732 30308
rect 18788 30252 18892 30308
rect 18948 30252 22092 30308
rect 22148 30252 22412 30308
rect 22468 30252 23132 30308
rect 23188 30252 23292 30308
rect 23348 30252 23452 30308
rect 23508 30252 23612 30308
rect 23668 30252 23772 30308
rect 23828 30252 23932 30308
rect 23988 30252 24092 30308
rect 24148 30252 24252 30308
rect 24308 30252 24412 30308
rect 24468 30252 24572 30308
rect 24628 30252 24732 30308
rect 24788 30252 24892 30308
rect 24948 30252 25052 30308
rect 25108 30252 25212 30308
rect 25268 30252 25372 30308
rect 25428 30252 25532 30308
rect 25588 30252 25692 30308
rect 25748 30252 25852 30308
rect 25908 30252 26012 30308
rect 26068 30252 26172 30308
rect 26228 30252 26332 30308
rect 26388 30252 26492 30308
rect 26548 30252 26652 30308
rect 26708 30252 26812 30308
rect 26868 30252 26972 30308
rect 27028 30252 27132 30308
rect 27188 30252 27292 30308
rect 27348 30252 27452 30308
rect 27508 30252 27612 30308
rect 27668 30252 27772 30308
rect 27828 30252 27932 30308
rect 27988 30252 28092 30308
rect 28148 30252 28252 30308
rect 28308 30252 28412 30308
rect 28468 30252 28572 30308
rect 28628 30252 28732 30308
rect 28788 30252 28892 30308
rect 28948 30252 29052 30308
rect 29108 30252 29212 30308
rect 29268 30252 29372 30308
rect 29428 30252 30012 30308
rect 30068 30252 30332 30308
rect 30388 30252 33532 30308
rect 33588 30252 33692 30308
rect 33748 30252 33852 30308
rect 33908 30252 34012 30308
rect 34068 30252 34172 30308
rect 34228 30252 34332 30308
rect 34388 30252 34492 30308
rect 34548 30252 34652 30308
rect 34708 30252 34812 30308
rect 34868 30252 34972 30308
rect 35028 30252 35132 30308
rect 35188 30252 35292 30308
rect 35348 30252 35452 30308
rect 35508 30252 35612 30308
rect 35668 30252 35772 30308
rect 35828 30252 35932 30308
rect 35988 30252 36092 30308
rect 36148 30252 36252 30308
rect 36308 30252 36412 30308
rect 36468 30252 36572 30308
rect 36628 30252 36732 30308
rect 36788 30252 36892 30308
rect 36948 30252 37052 30308
rect 37108 30252 37212 30308
rect 37268 30252 37372 30308
rect 37428 30252 37532 30308
rect 37588 30252 37692 30308
rect 37748 30252 37852 30308
rect 37908 30252 38012 30308
rect 38068 30252 38172 30308
rect 38228 30252 38332 30308
rect 38388 30252 38492 30308
rect 38548 30252 38652 30308
rect 38708 30252 38812 30308
rect 38868 30252 38972 30308
rect 39028 30252 39132 30308
rect 39188 30252 39292 30308
rect 39348 30252 39452 30308
rect 39508 30252 39612 30308
rect 39668 30252 39772 30308
rect 39828 30252 39932 30308
rect 39988 30252 40092 30308
rect 40148 30252 40252 30308
rect 40308 30252 40412 30308
rect 40468 30252 40572 30308
rect 40628 30252 40732 30308
rect 40788 30252 40892 30308
rect 40948 30252 41052 30308
rect 41108 30252 41212 30308
rect 41268 30252 41372 30308
rect 41428 30252 41532 30308
rect 41588 30252 41692 30308
rect 41748 30252 41852 30308
rect 41908 30252 41920 30308
rect 0 30240 41920 30252
rect 0 30148 41920 30160
rect 0 30092 11692 30148
rect 11748 30092 22252 30148
rect 22308 30092 30172 30148
rect 30228 30092 41920 30148
rect 0 30080 41920 30092
rect 0 29988 41920 30000
rect 0 29932 12 29988
rect 68 29932 172 29988
rect 228 29932 332 29988
rect 388 29932 492 29988
rect 548 29932 652 29988
rect 708 29932 812 29988
rect 868 29932 972 29988
rect 1028 29932 1132 29988
rect 1188 29932 1292 29988
rect 1348 29932 1452 29988
rect 1508 29932 1612 29988
rect 1668 29932 1772 29988
rect 1828 29932 1932 29988
rect 1988 29932 2092 29988
rect 2148 29932 2252 29988
rect 2308 29932 2412 29988
rect 2468 29932 2572 29988
rect 2628 29932 2732 29988
rect 2788 29932 2892 29988
rect 2948 29932 3052 29988
rect 3108 29932 3212 29988
rect 3268 29932 3372 29988
rect 3428 29932 3532 29988
rect 3588 29932 3692 29988
rect 3748 29932 3852 29988
rect 3908 29932 4012 29988
rect 4068 29932 4172 29988
rect 4228 29932 4332 29988
rect 4388 29932 4492 29988
rect 4548 29932 4652 29988
rect 4708 29932 4812 29988
rect 4868 29932 4972 29988
rect 5028 29932 5132 29988
rect 5188 29932 5292 29988
rect 5348 29932 5452 29988
rect 5508 29932 5612 29988
rect 5668 29932 5772 29988
rect 5828 29932 5932 29988
rect 5988 29932 6092 29988
rect 6148 29932 6252 29988
rect 6308 29932 6412 29988
rect 6468 29932 6572 29988
rect 6628 29932 6732 29988
rect 6788 29932 6892 29988
rect 6948 29932 7052 29988
rect 7108 29932 7212 29988
rect 7268 29932 7372 29988
rect 7428 29932 7532 29988
rect 7588 29932 7692 29988
rect 7748 29932 7852 29988
rect 7908 29932 8012 29988
rect 8068 29932 8172 29988
rect 8228 29932 8332 29988
rect 8388 29932 11532 29988
rect 11588 29932 11852 29988
rect 11908 29932 12492 29988
rect 12548 29932 12652 29988
rect 12708 29932 12812 29988
rect 12868 29932 12972 29988
rect 13028 29932 13132 29988
rect 13188 29932 13292 29988
rect 13348 29932 13452 29988
rect 13508 29932 13612 29988
rect 13668 29932 13772 29988
rect 13828 29932 13932 29988
rect 13988 29932 14092 29988
rect 14148 29932 14252 29988
rect 14308 29932 14412 29988
rect 14468 29932 14572 29988
rect 14628 29932 14732 29988
rect 14788 29932 14892 29988
rect 14948 29932 15052 29988
rect 15108 29932 15212 29988
rect 15268 29932 15372 29988
rect 15428 29932 15532 29988
rect 15588 29932 15692 29988
rect 15748 29932 15852 29988
rect 15908 29932 16012 29988
rect 16068 29932 16172 29988
rect 16228 29932 16332 29988
rect 16388 29932 16492 29988
rect 16548 29932 16652 29988
rect 16708 29932 16812 29988
rect 16868 29932 16972 29988
rect 17028 29932 17132 29988
rect 17188 29932 17292 29988
rect 17348 29932 17452 29988
rect 17508 29932 17612 29988
rect 17668 29932 17772 29988
rect 17828 29932 17932 29988
rect 17988 29932 18092 29988
rect 18148 29932 18252 29988
rect 18308 29932 18412 29988
rect 18468 29932 18572 29988
rect 18628 29932 18732 29988
rect 18788 29932 18892 29988
rect 18948 29932 22092 29988
rect 22148 29932 22412 29988
rect 22468 29932 23132 29988
rect 23188 29932 23292 29988
rect 23348 29932 23452 29988
rect 23508 29932 23612 29988
rect 23668 29932 23772 29988
rect 23828 29932 23932 29988
rect 23988 29932 24092 29988
rect 24148 29932 24252 29988
rect 24308 29932 24412 29988
rect 24468 29932 24572 29988
rect 24628 29932 24732 29988
rect 24788 29932 24892 29988
rect 24948 29932 25052 29988
rect 25108 29932 25212 29988
rect 25268 29932 25372 29988
rect 25428 29932 25532 29988
rect 25588 29932 25692 29988
rect 25748 29932 25852 29988
rect 25908 29932 26012 29988
rect 26068 29932 26172 29988
rect 26228 29932 26332 29988
rect 26388 29932 26492 29988
rect 26548 29932 26652 29988
rect 26708 29932 26812 29988
rect 26868 29932 26972 29988
rect 27028 29932 27132 29988
rect 27188 29932 27292 29988
rect 27348 29932 27452 29988
rect 27508 29932 27612 29988
rect 27668 29932 27772 29988
rect 27828 29932 27932 29988
rect 27988 29932 28092 29988
rect 28148 29932 28252 29988
rect 28308 29932 28412 29988
rect 28468 29932 28572 29988
rect 28628 29932 28732 29988
rect 28788 29932 28892 29988
rect 28948 29932 29052 29988
rect 29108 29932 29212 29988
rect 29268 29932 29372 29988
rect 29428 29932 30012 29988
rect 30068 29932 30332 29988
rect 30388 29932 33532 29988
rect 33588 29932 33692 29988
rect 33748 29932 33852 29988
rect 33908 29932 34012 29988
rect 34068 29932 34172 29988
rect 34228 29932 34332 29988
rect 34388 29932 34492 29988
rect 34548 29932 34652 29988
rect 34708 29932 34812 29988
rect 34868 29932 34972 29988
rect 35028 29932 35132 29988
rect 35188 29932 35292 29988
rect 35348 29932 35452 29988
rect 35508 29932 35612 29988
rect 35668 29932 35772 29988
rect 35828 29932 35932 29988
rect 35988 29932 36092 29988
rect 36148 29932 36252 29988
rect 36308 29932 36412 29988
rect 36468 29932 36572 29988
rect 36628 29932 36732 29988
rect 36788 29932 36892 29988
rect 36948 29932 37052 29988
rect 37108 29932 37212 29988
rect 37268 29932 37372 29988
rect 37428 29932 37532 29988
rect 37588 29932 37692 29988
rect 37748 29932 37852 29988
rect 37908 29932 38012 29988
rect 38068 29932 38172 29988
rect 38228 29932 38332 29988
rect 38388 29932 38492 29988
rect 38548 29932 38652 29988
rect 38708 29932 38812 29988
rect 38868 29932 38972 29988
rect 39028 29932 39132 29988
rect 39188 29932 39292 29988
rect 39348 29932 39452 29988
rect 39508 29932 39612 29988
rect 39668 29932 39772 29988
rect 39828 29932 39932 29988
rect 39988 29932 40092 29988
rect 40148 29932 40252 29988
rect 40308 29932 40412 29988
rect 40468 29932 40572 29988
rect 40628 29932 40732 29988
rect 40788 29932 40892 29988
rect 40948 29932 41052 29988
rect 41108 29932 41212 29988
rect 41268 29932 41372 29988
rect 41428 29932 41532 29988
rect 41588 29932 41692 29988
rect 41748 29932 41852 29988
rect 41908 29932 41920 29988
rect 0 29920 41920 29932
rect 0 29828 41920 29840
rect 0 29772 12 29828
rect 68 29772 172 29828
rect 228 29772 332 29828
rect 388 29772 492 29828
rect 548 29772 652 29828
rect 708 29772 812 29828
rect 868 29772 972 29828
rect 1028 29772 1132 29828
rect 1188 29772 1292 29828
rect 1348 29772 1452 29828
rect 1508 29772 1612 29828
rect 1668 29772 1772 29828
rect 1828 29772 1932 29828
rect 1988 29772 2092 29828
rect 2148 29772 2252 29828
rect 2308 29772 2412 29828
rect 2468 29772 2572 29828
rect 2628 29772 2732 29828
rect 2788 29772 2892 29828
rect 2948 29772 3052 29828
rect 3108 29772 3212 29828
rect 3268 29772 3372 29828
rect 3428 29772 3532 29828
rect 3588 29772 3692 29828
rect 3748 29772 3852 29828
rect 3908 29772 4012 29828
rect 4068 29772 4172 29828
rect 4228 29772 4332 29828
rect 4388 29772 4492 29828
rect 4548 29772 4652 29828
rect 4708 29772 4812 29828
rect 4868 29772 4972 29828
rect 5028 29772 5132 29828
rect 5188 29772 5292 29828
rect 5348 29772 5452 29828
rect 5508 29772 5612 29828
rect 5668 29772 5772 29828
rect 5828 29772 5932 29828
rect 5988 29772 6092 29828
rect 6148 29772 6252 29828
rect 6308 29772 6412 29828
rect 6468 29772 6572 29828
rect 6628 29772 6732 29828
rect 6788 29772 6892 29828
rect 6948 29772 7052 29828
rect 7108 29772 7212 29828
rect 7268 29772 7372 29828
rect 7428 29772 7532 29828
rect 7588 29772 7692 29828
rect 7748 29772 7852 29828
rect 7908 29772 8012 29828
rect 8068 29772 8172 29828
rect 8228 29772 8332 29828
rect 8388 29772 12012 29828
rect 12068 29772 12332 29828
rect 12388 29772 12492 29828
rect 12548 29772 12652 29828
rect 12708 29772 12812 29828
rect 12868 29772 12972 29828
rect 13028 29772 13132 29828
rect 13188 29772 13292 29828
rect 13348 29772 13452 29828
rect 13508 29772 13612 29828
rect 13668 29772 13772 29828
rect 13828 29772 13932 29828
rect 13988 29772 14092 29828
rect 14148 29772 14252 29828
rect 14308 29772 14412 29828
rect 14468 29772 14572 29828
rect 14628 29772 14732 29828
rect 14788 29772 14892 29828
rect 14948 29772 15052 29828
rect 15108 29772 15212 29828
rect 15268 29772 15372 29828
rect 15428 29772 15532 29828
rect 15588 29772 15692 29828
rect 15748 29772 15852 29828
rect 15908 29772 16012 29828
rect 16068 29772 16172 29828
rect 16228 29772 16332 29828
rect 16388 29772 16492 29828
rect 16548 29772 16652 29828
rect 16708 29772 16812 29828
rect 16868 29772 16972 29828
rect 17028 29772 17132 29828
rect 17188 29772 17292 29828
rect 17348 29772 17452 29828
rect 17508 29772 17612 29828
rect 17668 29772 17772 29828
rect 17828 29772 17932 29828
rect 17988 29772 18092 29828
rect 18148 29772 18252 29828
rect 18308 29772 18412 29828
rect 18468 29772 18572 29828
rect 18628 29772 18732 29828
rect 18788 29772 18892 29828
rect 18948 29772 22572 29828
rect 22628 29772 22892 29828
rect 22948 29772 23132 29828
rect 23188 29772 23292 29828
rect 23348 29772 23452 29828
rect 23508 29772 23612 29828
rect 23668 29772 23772 29828
rect 23828 29772 23932 29828
rect 23988 29772 24092 29828
rect 24148 29772 24252 29828
rect 24308 29772 24412 29828
rect 24468 29772 24572 29828
rect 24628 29772 24732 29828
rect 24788 29772 24892 29828
rect 24948 29772 25052 29828
rect 25108 29772 25212 29828
rect 25268 29772 25372 29828
rect 25428 29772 25532 29828
rect 25588 29772 25692 29828
rect 25748 29772 25852 29828
rect 25908 29772 26012 29828
rect 26068 29772 26172 29828
rect 26228 29772 26332 29828
rect 26388 29772 26492 29828
rect 26548 29772 26652 29828
rect 26708 29772 26812 29828
rect 26868 29772 26972 29828
rect 27028 29772 27132 29828
rect 27188 29772 27292 29828
rect 27348 29772 27452 29828
rect 27508 29772 27612 29828
rect 27668 29772 27772 29828
rect 27828 29772 27932 29828
rect 27988 29772 28092 29828
rect 28148 29772 28252 29828
rect 28308 29772 28412 29828
rect 28468 29772 28572 29828
rect 28628 29772 28732 29828
rect 28788 29772 28892 29828
rect 28948 29772 29052 29828
rect 29108 29772 29212 29828
rect 29268 29772 29372 29828
rect 29428 29772 29532 29828
rect 29588 29772 29852 29828
rect 29908 29772 33532 29828
rect 33588 29772 33692 29828
rect 33748 29772 33852 29828
rect 33908 29772 34012 29828
rect 34068 29772 34172 29828
rect 34228 29772 34332 29828
rect 34388 29772 34492 29828
rect 34548 29772 34652 29828
rect 34708 29772 34812 29828
rect 34868 29772 34972 29828
rect 35028 29772 35132 29828
rect 35188 29772 35292 29828
rect 35348 29772 35452 29828
rect 35508 29772 35612 29828
rect 35668 29772 35772 29828
rect 35828 29772 35932 29828
rect 35988 29772 36092 29828
rect 36148 29772 36252 29828
rect 36308 29772 36412 29828
rect 36468 29772 36572 29828
rect 36628 29772 36732 29828
rect 36788 29772 36892 29828
rect 36948 29772 37052 29828
rect 37108 29772 37212 29828
rect 37268 29772 37372 29828
rect 37428 29772 37532 29828
rect 37588 29772 37692 29828
rect 37748 29772 37852 29828
rect 37908 29772 38012 29828
rect 38068 29772 38172 29828
rect 38228 29772 38332 29828
rect 38388 29772 38492 29828
rect 38548 29772 38652 29828
rect 38708 29772 38812 29828
rect 38868 29772 38972 29828
rect 39028 29772 39132 29828
rect 39188 29772 39292 29828
rect 39348 29772 39452 29828
rect 39508 29772 39612 29828
rect 39668 29772 39772 29828
rect 39828 29772 39932 29828
rect 39988 29772 40092 29828
rect 40148 29772 40252 29828
rect 40308 29772 40412 29828
rect 40468 29772 40572 29828
rect 40628 29772 40732 29828
rect 40788 29772 40892 29828
rect 40948 29772 41052 29828
rect 41108 29772 41212 29828
rect 41268 29772 41372 29828
rect 41428 29772 41532 29828
rect 41588 29772 41692 29828
rect 41748 29772 41852 29828
rect 41908 29772 41920 29828
rect 0 29760 41920 29772
rect 0 29668 41920 29680
rect 0 29612 12172 29668
rect 12228 29612 22732 29668
rect 22788 29612 29692 29668
rect 29748 29612 41920 29668
rect 0 29600 41920 29612
rect 0 29508 41920 29520
rect 0 29452 12 29508
rect 68 29452 172 29508
rect 228 29452 332 29508
rect 388 29452 492 29508
rect 548 29452 652 29508
rect 708 29452 812 29508
rect 868 29452 972 29508
rect 1028 29452 1132 29508
rect 1188 29452 1292 29508
rect 1348 29452 1452 29508
rect 1508 29452 1612 29508
rect 1668 29452 1772 29508
rect 1828 29452 1932 29508
rect 1988 29452 2092 29508
rect 2148 29452 2252 29508
rect 2308 29452 2412 29508
rect 2468 29452 2572 29508
rect 2628 29452 2732 29508
rect 2788 29452 2892 29508
rect 2948 29452 3052 29508
rect 3108 29452 3212 29508
rect 3268 29452 3372 29508
rect 3428 29452 3532 29508
rect 3588 29452 3692 29508
rect 3748 29452 3852 29508
rect 3908 29452 4012 29508
rect 4068 29452 4172 29508
rect 4228 29452 4332 29508
rect 4388 29452 4492 29508
rect 4548 29452 4652 29508
rect 4708 29452 4812 29508
rect 4868 29452 4972 29508
rect 5028 29452 5132 29508
rect 5188 29452 5292 29508
rect 5348 29452 5452 29508
rect 5508 29452 5612 29508
rect 5668 29452 5772 29508
rect 5828 29452 5932 29508
rect 5988 29452 6092 29508
rect 6148 29452 6252 29508
rect 6308 29452 6412 29508
rect 6468 29452 6572 29508
rect 6628 29452 6732 29508
rect 6788 29452 6892 29508
rect 6948 29452 7052 29508
rect 7108 29452 7212 29508
rect 7268 29452 7372 29508
rect 7428 29452 7532 29508
rect 7588 29452 7692 29508
rect 7748 29452 7852 29508
rect 7908 29452 8012 29508
rect 8068 29452 8172 29508
rect 8228 29452 8332 29508
rect 8388 29452 12012 29508
rect 12068 29452 12332 29508
rect 12388 29452 12492 29508
rect 12548 29452 12652 29508
rect 12708 29452 12812 29508
rect 12868 29452 12972 29508
rect 13028 29452 13132 29508
rect 13188 29452 13292 29508
rect 13348 29452 13452 29508
rect 13508 29452 13612 29508
rect 13668 29452 13772 29508
rect 13828 29452 13932 29508
rect 13988 29452 14092 29508
rect 14148 29452 14252 29508
rect 14308 29452 14412 29508
rect 14468 29452 14572 29508
rect 14628 29452 14732 29508
rect 14788 29452 14892 29508
rect 14948 29452 15052 29508
rect 15108 29452 15212 29508
rect 15268 29452 15372 29508
rect 15428 29452 15532 29508
rect 15588 29452 15692 29508
rect 15748 29452 15852 29508
rect 15908 29452 16012 29508
rect 16068 29452 16172 29508
rect 16228 29452 16332 29508
rect 16388 29452 16492 29508
rect 16548 29452 16652 29508
rect 16708 29452 16812 29508
rect 16868 29452 16972 29508
rect 17028 29452 17132 29508
rect 17188 29452 17292 29508
rect 17348 29452 17452 29508
rect 17508 29452 17612 29508
rect 17668 29452 17772 29508
rect 17828 29452 17932 29508
rect 17988 29452 18092 29508
rect 18148 29452 18252 29508
rect 18308 29452 18412 29508
rect 18468 29452 18572 29508
rect 18628 29452 18732 29508
rect 18788 29452 18892 29508
rect 18948 29452 22572 29508
rect 22628 29452 22892 29508
rect 22948 29452 23132 29508
rect 23188 29452 23292 29508
rect 23348 29452 23452 29508
rect 23508 29452 23612 29508
rect 23668 29452 23772 29508
rect 23828 29452 23932 29508
rect 23988 29452 24092 29508
rect 24148 29452 24252 29508
rect 24308 29452 24412 29508
rect 24468 29452 24572 29508
rect 24628 29452 24732 29508
rect 24788 29452 24892 29508
rect 24948 29452 25052 29508
rect 25108 29452 25212 29508
rect 25268 29452 25372 29508
rect 25428 29452 25532 29508
rect 25588 29452 25692 29508
rect 25748 29452 25852 29508
rect 25908 29452 26012 29508
rect 26068 29452 26172 29508
rect 26228 29452 26332 29508
rect 26388 29452 26492 29508
rect 26548 29452 26652 29508
rect 26708 29452 26812 29508
rect 26868 29452 26972 29508
rect 27028 29452 27132 29508
rect 27188 29452 27292 29508
rect 27348 29452 27452 29508
rect 27508 29452 27612 29508
rect 27668 29452 27772 29508
rect 27828 29452 27932 29508
rect 27988 29452 28092 29508
rect 28148 29452 28252 29508
rect 28308 29452 28412 29508
rect 28468 29452 28572 29508
rect 28628 29452 28732 29508
rect 28788 29452 28892 29508
rect 28948 29452 29052 29508
rect 29108 29452 29212 29508
rect 29268 29452 29372 29508
rect 29428 29452 29532 29508
rect 29588 29452 29852 29508
rect 29908 29452 33532 29508
rect 33588 29452 33692 29508
rect 33748 29452 33852 29508
rect 33908 29452 34012 29508
rect 34068 29452 34172 29508
rect 34228 29452 34332 29508
rect 34388 29452 34492 29508
rect 34548 29452 34652 29508
rect 34708 29452 34812 29508
rect 34868 29452 34972 29508
rect 35028 29452 35132 29508
rect 35188 29452 35292 29508
rect 35348 29452 35452 29508
rect 35508 29452 35612 29508
rect 35668 29452 35772 29508
rect 35828 29452 35932 29508
rect 35988 29452 36092 29508
rect 36148 29452 36252 29508
rect 36308 29452 36412 29508
rect 36468 29452 36572 29508
rect 36628 29452 36732 29508
rect 36788 29452 36892 29508
rect 36948 29452 37052 29508
rect 37108 29452 37212 29508
rect 37268 29452 37372 29508
rect 37428 29452 37532 29508
rect 37588 29452 37692 29508
rect 37748 29452 37852 29508
rect 37908 29452 38012 29508
rect 38068 29452 38172 29508
rect 38228 29452 38332 29508
rect 38388 29452 38492 29508
rect 38548 29452 38652 29508
rect 38708 29452 38812 29508
rect 38868 29452 38972 29508
rect 39028 29452 39132 29508
rect 39188 29452 39292 29508
rect 39348 29452 39452 29508
rect 39508 29452 39612 29508
rect 39668 29452 39772 29508
rect 39828 29452 39932 29508
rect 39988 29452 40092 29508
rect 40148 29452 40252 29508
rect 40308 29452 40412 29508
rect 40468 29452 40572 29508
rect 40628 29452 40732 29508
rect 40788 29452 40892 29508
rect 40948 29452 41052 29508
rect 41108 29452 41212 29508
rect 41268 29452 41372 29508
rect 41428 29452 41532 29508
rect 41588 29452 41692 29508
rect 41748 29452 41852 29508
rect 41908 29452 41920 29508
rect 0 29440 41920 29452
<< via2 >>
rect 12 37346 68 37348
rect 12 37294 14 37346
rect 14 37294 66 37346
rect 66 37294 68 37346
rect 12 37292 68 37294
rect 172 37346 228 37348
rect 172 37294 174 37346
rect 174 37294 226 37346
rect 226 37294 228 37346
rect 172 37292 228 37294
rect 332 37346 388 37348
rect 332 37294 334 37346
rect 334 37294 386 37346
rect 386 37294 388 37346
rect 332 37292 388 37294
rect 492 37346 548 37348
rect 492 37294 494 37346
rect 494 37294 546 37346
rect 546 37294 548 37346
rect 492 37292 548 37294
rect 652 37346 708 37348
rect 652 37294 654 37346
rect 654 37294 706 37346
rect 706 37294 708 37346
rect 652 37292 708 37294
rect 812 37346 868 37348
rect 812 37294 814 37346
rect 814 37294 866 37346
rect 866 37294 868 37346
rect 812 37292 868 37294
rect 972 37346 1028 37348
rect 972 37294 974 37346
rect 974 37294 1026 37346
rect 1026 37294 1028 37346
rect 972 37292 1028 37294
rect 1132 37346 1188 37348
rect 1132 37294 1134 37346
rect 1134 37294 1186 37346
rect 1186 37294 1188 37346
rect 1132 37292 1188 37294
rect 1292 37346 1348 37348
rect 1292 37294 1294 37346
rect 1294 37294 1346 37346
rect 1346 37294 1348 37346
rect 1292 37292 1348 37294
rect 1452 37346 1508 37348
rect 1452 37294 1454 37346
rect 1454 37294 1506 37346
rect 1506 37294 1508 37346
rect 1452 37292 1508 37294
rect 1612 37346 1668 37348
rect 1612 37294 1614 37346
rect 1614 37294 1666 37346
rect 1666 37294 1668 37346
rect 1612 37292 1668 37294
rect 1772 37346 1828 37348
rect 1772 37294 1774 37346
rect 1774 37294 1826 37346
rect 1826 37294 1828 37346
rect 1772 37292 1828 37294
rect 1932 37346 1988 37348
rect 1932 37294 1934 37346
rect 1934 37294 1986 37346
rect 1986 37294 1988 37346
rect 1932 37292 1988 37294
rect 2092 37346 2148 37348
rect 2092 37294 2094 37346
rect 2094 37294 2146 37346
rect 2146 37294 2148 37346
rect 2092 37292 2148 37294
rect 2252 37346 2308 37348
rect 2252 37294 2254 37346
rect 2254 37294 2306 37346
rect 2306 37294 2308 37346
rect 2252 37292 2308 37294
rect 2412 37346 2468 37348
rect 2412 37294 2414 37346
rect 2414 37294 2466 37346
rect 2466 37294 2468 37346
rect 2412 37292 2468 37294
rect 2572 37346 2628 37348
rect 2572 37294 2574 37346
rect 2574 37294 2626 37346
rect 2626 37294 2628 37346
rect 2572 37292 2628 37294
rect 2732 37346 2788 37348
rect 2732 37294 2734 37346
rect 2734 37294 2786 37346
rect 2786 37294 2788 37346
rect 2732 37292 2788 37294
rect 2892 37346 2948 37348
rect 2892 37294 2894 37346
rect 2894 37294 2946 37346
rect 2946 37294 2948 37346
rect 2892 37292 2948 37294
rect 3052 37346 3108 37348
rect 3052 37294 3054 37346
rect 3054 37294 3106 37346
rect 3106 37294 3108 37346
rect 3052 37292 3108 37294
rect 3212 37346 3268 37348
rect 3212 37294 3214 37346
rect 3214 37294 3266 37346
rect 3266 37294 3268 37346
rect 3212 37292 3268 37294
rect 3372 37346 3428 37348
rect 3372 37294 3374 37346
rect 3374 37294 3426 37346
rect 3426 37294 3428 37346
rect 3372 37292 3428 37294
rect 3532 37346 3588 37348
rect 3532 37294 3534 37346
rect 3534 37294 3586 37346
rect 3586 37294 3588 37346
rect 3532 37292 3588 37294
rect 3692 37346 3748 37348
rect 3692 37294 3694 37346
rect 3694 37294 3746 37346
rect 3746 37294 3748 37346
rect 3692 37292 3748 37294
rect 3852 37346 3908 37348
rect 3852 37294 3854 37346
rect 3854 37294 3906 37346
rect 3906 37294 3908 37346
rect 3852 37292 3908 37294
rect 4012 37346 4068 37348
rect 4012 37294 4014 37346
rect 4014 37294 4066 37346
rect 4066 37294 4068 37346
rect 4012 37292 4068 37294
rect 4172 37346 4228 37348
rect 4172 37294 4174 37346
rect 4174 37294 4226 37346
rect 4226 37294 4228 37346
rect 4172 37292 4228 37294
rect 4332 37346 4388 37348
rect 4332 37294 4334 37346
rect 4334 37294 4386 37346
rect 4386 37294 4388 37346
rect 4332 37292 4388 37294
rect 4492 37346 4548 37348
rect 4492 37294 4494 37346
rect 4494 37294 4546 37346
rect 4546 37294 4548 37346
rect 4492 37292 4548 37294
rect 4652 37346 4708 37348
rect 4652 37294 4654 37346
rect 4654 37294 4706 37346
rect 4706 37294 4708 37346
rect 4652 37292 4708 37294
rect 4812 37346 4868 37348
rect 4812 37294 4814 37346
rect 4814 37294 4866 37346
rect 4866 37294 4868 37346
rect 4812 37292 4868 37294
rect 4972 37346 5028 37348
rect 4972 37294 4974 37346
rect 4974 37294 5026 37346
rect 5026 37294 5028 37346
rect 4972 37292 5028 37294
rect 5132 37346 5188 37348
rect 5132 37294 5134 37346
rect 5134 37294 5186 37346
rect 5186 37294 5188 37346
rect 5132 37292 5188 37294
rect 5292 37346 5348 37348
rect 5292 37294 5294 37346
rect 5294 37294 5346 37346
rect 5346 37294 5348 37346
rect 5292 37292 5348 37294
rect 5452 37346 5508 37348
rect 5452 37294 5454 37346
rect 5454 37294 5506 37346
rect 5506 37294 5508 37346
rect 5452 37292 5508 37294
rect 5612 37346 5668 37348
rect 5612 37294 5614 37346
rect 5614 37294 5666 37346
rect 5666 37294 5668 37346
rect 5612 37292 5668 37294
rect 5772 37346 5828 37348
rect 5772 37294 5774 37346
rect 5774 37294 5826 37346
rect 5826 37294 5828 37346
rect 5772 37292 5828 37294
rect 5932 37346 5988 37348
rect 5932 37294 5934 37346
rect 5934 37294 5986 37346
rect 5986 37294 5988 37346
rect 5932 37292 5988 37294
rect 6092 37346 6148 37348
rect 6092 37294 6094 37346
rect 6094 37294 6146 37346
rect 6146 37294 6148 37346
rect 6092 37292 6148 37294
rect 6252 37346 6308 37348
rect 6252 37294 6254 37346
rect 6254 37294 6306 37346
rect 6306 37294 6308 37346
rect 6252 37292 6308 37294
rect 6412 37346 6468 37348
rect 6412 37294 6414 37346
rect 6414 37294 6466 37346
rect 6466 37294 6468 37346
rect 6412 37292 6468 37294
rect 6572 37346 6628 37348
rect 6572 37294 6574 37346
rect 6574 37294 6626 37346
rect 6626 37294 6628 37346
rect 6572 37292 6628 37294
rect 6732 37346 6788 37348
rect 6732 37294 6734 37346
rect 6734 37294 6786 37346
rect 6786 37294 6788 37346
rect 6732 37292 6788 37294
rect 6892 37346 6948 37348
rect 6892 37294 6894 37346
rect 6894 37294 6946 37346
rect 6946 37294 6948 37346
rect 6892 37292 6948 37294
rect 7052 37346 7108 37348
rect 7052 37294 7054 37346
rect 7054 37294 7106 37346
rect 7106 37294 7108 37346
rect 7052 37292 7108 37294
rect 7212 37346 7268 37348
rect 7212 37294 7214 37346
rect 7214 37294 7266 37346
rect 7266 37294 7268 37346
rect 7212 37292 7268 37294
rect 7372 37346 7428 37348
rect 7372 37294 7374 37346
rect 7374 37294 7426 37346
rect 7426 37294 7428 37346
rect 7372 37292 7428 37294
rect 7532 37346 7588 37348
rect 7532 37294 7534 37346
rect 7534 37294 7586 37346
rect 7586 37294 7588 37346
rect 7532 37292 7588 37294
rect 7692 37346 7748 37348
rect 7692 37294 7694 37346
rect 7694 37294 7746 37346
rect 7746 37294 7748 37346
rect 7692 37292 7748 37294
rect 7852 37346 7908 37348
rect 7852 37294 7854 37346
rect 7854 37294 7906 37346
rect 7906 37294 7908 37346
rect 7852 37292 7908 37294
rect 8012 37346 8068 37348
rect 8012 37294 8014 37346
rect 8014 37294 8066 37346
rect 8066 37294 8068 37346
rect 8012 37292 8068 37294
rect 8172 37346 8228 37348
rect 8172 37294 8174 37346
rect 8174 37294 8226 37346
rect 8226 37294 8228 37346
rect 8172 37292 8228 37294
rect 8332 37346 8388 37348
rect 8332 37294 8334 37346
rect 8334 37294 8386 37346
rect 8386 37294 8388 37346
rect 8332 37292 8388 37294
rect 8492 37292 8548 37348
rect 8812 37292 8868 37348
rect 12492 37346 12548 37348
rect 12492 37294 12494 37346
rect 12494 37294 12546 37346
rect 12546 37294 12548 37346
rect 12492 37292 12548 37294
rect 12652 37346 12708 37348
rect 12652 37294 12654 37346
rect 12654 37294 12706 37346
rect 12706 37294 12708 37346
rect 12652 37292 12708 37294
rect 12812 37346 12868 37348
rect 12812 37294 12814 37346
rect 12814 37294 12866 37346
rect 12866 37294 12868 37346
rect 12812 37292 12868 37294
rect 12972 37346 13028 37348
rect 12972 37294 12974 37346
rect 12974 37294 13026 37346
rect 13026 37294 13028 37346
rect 12972 37292 13028 37294
rect 13132 37346 13188 37348
rect 13132 37294 13134 37346
rect 13134 37294 13186 37346
rect 13186 37294 13188 37346
rect 13132 37292 13188 37294
rect 13292 37346 13348 37348
rect 13292 37294 13294 37346
rect 13294 37294 13346 37346
rect 13346 37294 13348 37346
rect 13292 37292 13348 37294
rect 13452 37346 13508 37348
rect 13452 37294 13454 37346
rect 13454 37294 13506 37346
rect 13506 37294 13508 37346
rect 13452 37292 13508 37294
rect 13612 37346 13668 37348
rect 13612 37294 13614 37346
rect 13614 37294 13666 37346
rect 13666 37294 13668 37346
rect 13612 37292 13668 37294
rect 13772 37346 13828 37348
rect 13772 37294 13774 37346
rect 13774 37294 13826 37346
rect 13826 37294 13828 37346
rect 13772 37292 13828 37294
rect 13932 37346 13988 37348
rect 13932 37294 13934 37346
rect 13934 37294 13986 37346
rect 13986 37294 13988 37346
rect 13932 37292 13988 37294
rect 14092 37346 14148 37348
rect 14092 37294 14094 37346
rect 14094 37294 14146 37346
rect 14146 37294 14148 37346
rect 14092 37292 14148 37294
rect 14252 37346 14308 37348
rect 14252 37294 14254 37346
rect 14254 37294 14306 37346
rect 14306 37294 14308 37346
rect 14252 37292 14308 37294
rect 14412 37346 14468 37348
rect 14412 37294 14414 37346
rect 14414 37294 14466 37346
rect 14466 37294 14468 37346
rect 14412 37292 14468 37294
rect 14572 37346 14628 37348
rect 14572 37294 14574 37346
rect 14574 37294 14626 37346
rect 14626 37294 14628 37346
rect 14572 37292 14628 37294
rect 14732 37346 14788 37348
rect 14732 37294 14734 37346
rect 14734 37294 14786 37346
rect 14786 37294 14788 37346
rect 14732 37292 14788 37294
rect 14892 37346 14948 37348
rect 14892 37294 14894 37346
rect 14894 37294 14946 37346
rect 14946 37294 14948 37346
rect 14892 37292 14948 37294
rect 15052 37346 15108 37348
rect 15052 37294 15054 37346
rect 15054 37294 15106 37346
rect 15106 37294 15108 37346
rect 15052 37292 15108 37294
rect 15212 37346 15268 37348
rect 15212 37294 15214 37346
rect 15214 37294 15266 37346
rect 15266 37294 15268 37346
rect 15212 37292 15268 37294
rect 15372 37346 15428 37348
rect 15372 37294 15374 37346
rect 15374 37294 15426 37346
rect 15426 37294 15428 37346
rect 15372 37292 15428 37294
rect 15532 37346 15588 37348
rect 15532 37294 15534 37346
rect 15534 37294 15586 37346
rect 15586 37294 15588 37346
rect 15532 37292 15588 37294
rect 15692 37346 15748 37348
rect 15692 37294 15694 37346
rect 15694 37294 15746 37346
rect 15746 37294 15748 37346
rect 15692 37292 15748 37294
rect 15852 37346 15908 37348
rect 15852 37294 15854 37346
rect 15854 37294 15906 37346
rect 15906 37294 15908 37346
rect 15852 37292 15908 37294
rect 16012 37346 16068 37348
rect 16012 37294 16014 37346
rect 16014 37294 16066 37346
rect 16066 37294 16068 37346
rect 16012 37292 16068 37294
rect 16172 37346 16228 37348
rect 16172 37294 16174 37346
rect 16174 37294 16226 37346
rect 16226 37294 16228 37346
rect 16172 37292 16228 37294
rect 16332 37346 16388 37348
rect 16332 37294 16334 37346
rect 16334 37294 16386 37346
rect 16386 37294 16388 37346
rect 16332 37292 16388 37294
rect 16492 37346 16548 37348
rect 16492 37294 16494 37346
rect 16494 37294 16546 37346
rect 16546 37294 16548 37346
rect 16492 37292 16548 37294
rect 16652 37346 16708 37348
rect 16652 37294 16654 37346
rect 16654 37294 16706 37346
rect 16706 37294 16708 37346
rect 16652 37292 16708 37294
rect 16812 37346 16868 37348
rect 16812 37294 16814 37346
rect 16814 37294 16866 37346
rect 16866 37294 16868 37346
rect 16812 37292 16868 37294
rect 16972 37346 17028 37348
rect 16972 37294 16974 37346
rect 16974 37294 17026 37346
rect 17026 37294 17028 37346
rect 16972 37292 17028 37294
rect 17132 37346 17188 37348
rect 17132 37294 17134 37346
rect 17134 37294 17186 37346
rect 17186 37294 17188 37346
rect 17132 37292 17188 37294
rect 17292 37346 17348 37348
rect 17292 37294 17294 37346
rect 17294 37294 17346 37346
rect 17346 37294 17348 37346
rect 17292 37292 17348 37294
rect 17452 37346 17508 37348
rect 17452 37294 17454 37346
rect 17454 37294 17506 37346
rect 17506 37294 17508 37346
rect 17452 37292 17508 37294
rect 17612 37346 17668 37348
rect 17612 37294 17614 37346
rect 17614 37294 17666 37346
rect 17666 37294 17668 37346
rect 17612 37292 17668 37294
rect 17772 37346 17828 37348
rect 17772 37294 17774 37346
rect 17774 37294 17826 37346
rect 17826 37294 17828 37346
rect 17772 37292 17828 37294
rect 17932 37346 17988 37348
rect 17932 37294 17934 37346
rect 17934 37294 17986 37346
rect 17986 37294 17988 37346
rect 17932 37292 17988 37294
rect 18092 37346 18148 37348
rect 18092 37294 18094 37346
rect 18094 37294 18146 37346
rect 18146 37294 18148 37346
rect 18092 37292 18148 37294
rect 18252 37346 18308 37348
rect 18252 37294 18254 37346
rect 18254 37294 18306 37346
rect 18306 37294 18308 37346
rect 18252 37292 18308 37294
rect 18412 37346 18468 37348
rect 18412 37294 18414 37346
rect 18414 37294 18466 37346
rect 18466 37294 18468 37346
rect 18412 37292 18468 37294
rect 18572 37346 18628 37348
rect 18572 37294 18574 37346
rect 18574 37294 18626 37346
rect 18626 37294 18628 37346
rect 18572 37292 18628 37294
rect 18732 37346 18788 37348
rect 18732 37294 18734 37346
rect 18734 37294 18786 37346
rect 18786 37294 18788 37346
rect 18732 37292 18788 37294
rect 18892 37346 18948 37348
rect 18892 37294 18894 37346
rect 18894 37294 18946 37346
rect 18946 37294 18948 37346
rect 18892 37292 18948 37294
rect 22572 37292 22628 37348
rect 22892 37292 22948 37348
rect 23132 37346 23188 37348
rect 23132 37294 23134 37346
rect 23134 37294 23186 37346
rect 23186 37294 23188 37346
rect 23132 37292 23188 37294
rect 23292 37346 23348 37348
rect 23292 37294 23294 37346
rect 23294 37294 23346 37346
rect 23346 37294 23348 37346
rect 23292 37292 23348 37294
rect 23452 37346 23508 37348
rect 23452 37294 23454 37346
rect 23454 37294 23506 37346
rect 23506 37294 23508 37346
rect 23452 37292 23508 37294
rect 23612 37346 23668 37348
rect 23612 37294 23614 37346
rect 23614 37294 23666 37346
rect 23666 37294 23668 37346
rect 23612 37292 23668 37294
rect 23772 37346 23828 37348
rect 23772 37294 23774 37346
rect 23774 37294 23826 37346
rect 23826 37294 23828 37346
rect 23772 37292 23828 37294
rect 23932 37346 23988 37348
rect 23932 37294 23934 37346
rect 23934 37294 23986 37346
rect 23986 37294 23988 37346
rect 23932 37292 23988 37294
rect 24092 37346 24148 37348
rect 24092 37294 24094 37346
rect 24094 37294 24146 37346
rect 24146 37294 24148 37346
rect 24092 37292 24148 37294
rect 24252 37346 24308 37348
rect 24252 37294 24254 37346
rect 24254 37294 24306 37346
rect 24306 37294 24308 37346
rect 24252 37292 24308 37294
rect 24412 37346 24468 37348
rect 24412 37294 24414 37346
rect 24414 37294 24466 37346
rect 24466 37294 24468 37346
rect 24412 37292 24468 37294
rect 24572 37346 24628 37348
rect 24572 37294 24574 37346
rect 24574 37294 24626 37346
rect 24626 37294 24628 37346
rect 24572 37292 24628 37294
rect 24732 37346 24788 37348
rect 24732 37294 24734 37346
rect 24734 37294 24786 37346
rect 24786 37294 24788 37346
rect 24732 37292 24788 37294
rect 24892 37346 24948 37348
rect 24892 37294 24894 37346
rect 24894 37294 24946 37346
rect 24946 37294 24948 37346
rect 24892 37292 24948 37294
rect 25052 37346 25108 37348
rect 25052 37294 25054 37346
rect 25054 37294 25106 37346
rect 25106 37294 25108 37346
rect 25052 37292 25108 37294
rect 25212 37346 25268 37348
rect 25212 37294 25214 37346
rect 25214 37294 25266 37346
rect 25266 37294 25268 37346
rect 25212 37292 25268 37294
rect 25372 37346 25428 37348
rect 25372 37294 25374 37346
rect 25374 37294 25426 37346
rect 25426 37294 25428 37346
rect 25372 37292 25428 37294
rect 25532 37346 25588 37348
rect 25532 37294 25534 37346
rect 25534 37294 25586 37346
rect 25586 37294 25588 37346
rect 25532 37292 25588 37294
rect 25692 37346 25748 37348
rect 25692 37294 25694 37346
rect 25694 37294 25746 37346
rect 25746 37294 25748 37346
rect 25692 37292 25748 37294
rect 25852 37346 25908 37348
rect 25852 37294 25854 37346
rect 25854 37294 25906 37346
rect 25906 37294 25908 37346
rect 25852 37292 25908 37294
rect 26012 37346 26068 37348
rect 26012 37294 26014 37346
rect 26014 37294 26066 37346
rect 26066 37294 26068 37346
rect 26012 37292 26068 37294
rect 26172 37346 26228 37348
rect 26172 37294 26174 37346
rect 26174 37294 26226 37346
rect 26226 37294 26228 37346
rect 26172 37292 26228 37294
rect 26332 37346 26388 37348
rect 26332 37294 26334 37346
rect 26334 37294 26386 37346
rect 26386 37294 26388 37346
rect 26332 37292 26388 37294
rect 26492 37346 26548 37348
rect 26492 37294 26494 37346
rect 26494 37294 26546 37346
rect 26546 37294 26548 37346
rect 26492 37292 26548 37294
rect 26652 37346 26708 37348
rect 26652 37294 26654 37346
rect 26654 37294 26706 37346
rect 26706 37294 26708 37346
rect 26652 37292 26708 37294
rect 26812 37346 26868 37348
rect 26812 37294 26814 37346
rect 26814 37294 26866 37346
rect 26866 37294 26868 37346
rect 26812 37292 26868 37294
rect 26972 37346 27028 37348
rect 26972 37294 26974 37346
rect 26974 37294 27026 37346
rect 27026 37294 27028 37346
rect 26972 37292 27028 37294
rect 27132 37346 27188 37348
rect 27132 37294 27134 37346
rect 27134 37294 27186 37346
rect 27186 37294 27188 37346
rect 27132 37292 27188 37294
rect 27292 37346 27348 37348
rect 27292 37294 27294 37346
rect 27294 37294 27346 37346
rect 27346 37294 27348 37346
rect 27292 37292 27348 37294
rect 27452 37346 27508 37348
rect 27452 37294 27454 37346
rect 27454 37294 27506 37346
rect 27506 37294 27508 37346
rect 27452 37292 27508 37294
rect 27612 37346 27668 37348
rect 27612 37294 27614 37346
rect 27614 37294 27666 37346
rect 27666 37294 27668 37346
rect 27612 37292 27668 37294
rect 27772 37346 27828 37348
rect 27772 37294 27774 37346
rect 27774 37294 27826 37346
rect 27826 37294 27828 37346
rect 27772 37292 27828 37294
rect 27932 37346 27988 37348
rect 27932 37294 27934 37346
rect 27934 37294 27986 37346
rect 27986 37294 27988 37346
rect 27932 37292 27988 37294
rect 28092 37346 28148 37348
rect 28092 37294 28094 37346
rect 28094 37294 28146 37346
rect 28146 37294 28148 37346
rect 28092 37292 28148 37294
rect 28252 37346 28308 37348
rect 28252 37294 28254 37346
rect 28254 37294 28306 37346
rect 28306 37294 28308 37346
rect 28252 37292 28308 37294
rect 28412 37346 28468 37348
rect 28412 37294 28414 37346
rect 28414 37294 28466 37346
rect 28466 37294 28468 37346
rect 28412 37292 28468 37294
rect 28572 37346 28628 37348
rect 28572 37294 28574 37346
rect 28574 37294 28626 37346
rect 28626 37294 28628 37346
rect 28572 37292 28628 37294
rect 28732 37346 28788 37348
rect 28732 37294 28734 37346
rect 28734 37294 28786 37346
rect 28786 37294 28788 37346
rect 28732 37292 28788 37294
rect 28892 37346 28948 37348
rect 28892 37294 28894 37346
rect 28894 37294 28946 37346
rect 28946 37294 28948 37346
rect 28892 37292 28948 37294
rect 29052 37346 29108 37348
rect 29052 37294 29054 37346
rect 29054 37294 29106 37346
rect 29106 37294 29108 37346
rect 29052 37292 29108 37294
rect 29212 37346 29268 37348
rect 29212 37294 29214 37346
rect 29214 37294 29266 37346
rect 29266 37294 29268 37346
rect 29212 37292 29268 37294
rect 29372 37346 29428 37348
rect 29372 37294 29374 37346
rect 29374 37294 29426 37346
rect 29426 37294 29428 37346
rect 29372 37292 29428 37294
rect 33052 37292 33108 37348
rect 33372 37292 33428 37348
rect 33532 37346 33588 37348
rect 33532 37294 33534 37346
rect 33534 37294 33586 37346
rect 33586 37294 33588 37346
rect 33532 37292 33588 37294
rect 33692 37346 33748 37348
rect 33692 37294 33694 37346
rect 33694 37294 33746 37346
rect 33746 37294 33748 37346
rect 33692 37292 33748 37294
rect 33852 37346 33908 37348
rect 33852 37294 33854 37346
rect 33854 37294 33906 37346
rect 33906 37294 33908 37346
rect 33852 37292 33908 37294
rect 34012 37346 34068 37348
rect 34012 37294 34014 37346
rect 34014 37294 34066 37346
rect 34066 37294 34068 37346
rect 34012 37292 34068 37294
rect 34172 37346 34228 37348
rect 34172 37294 34174 37346
rect 34174 37294 34226 37346
rect 34226 37294 34228 37346
rect 34172 37292 34228 37294
rect 34332 37346 34388 37348
rect 34332 37294 34334 37346
rect 34334 37294 34386 37346
rect 34386 37294 34388 37346
rect 34332 37292 34388 37294
rect 34492 37346 34548 37348
rect 34492 37294 34494 37346
rect 34494 37294 34546 37346
rect 34546 37294 34548 37346
rect 34492 37292 34548 37294
rect 34652 37346 34708 37348
rect 34652 37294 34654 37346
rect 34654 37294 34706 37346
rect 34706 37294 34708 37346
rect 34652 37292 34708 37294
rect 34812 37346 34868 37348
rect 34812 37294 34814 37346
rect 34814 37294 34866 37346
rect 34866 37294 34868 37346
rect 34812 37292 34868 37294
rect 34972 37346 35028 37348
rect 34972 37294 34974 37346
rect 34974 37294 35026 37346
rect 35026 37294 35028 37346
rect 34972 37292 35028 37294
rect 35132 37346 35188 37348
rect 35132 37294 35134 37346
rect 35134 37294 35186 37346
rect 35186 37294 35188 37346
rect 35132 37292 35188 37294
rect 35292 37346 35348 37348
rect 35292 37294 35294 37346
rect 35294 37294 35346 37346
rect 35346 37294 35348 37346
rect 35292 37292 35348 37294
rect 35452 37346 35508 37348
rect 35452 37294 35454 37346
rect 35454 37294 35506 37346
rect 35506 37294 35508 37346
rect 35452 37292 35508 37294
rect 35612 37346 35668 37348
rect 35612 37294 35614 37346
rect 35614 37294 35666 37346
rect 35666 37294 35668 37346
rect 35612 37292 35668 37294
rect 35772 37346 35828 37348
rect 35772 37294 35774 37346
rect 35774 37294 35826 37346
rect 35826 37294 35828 37346
rect 35772 37292 35828 37294
rect 35932 37346 35988 37348
rect 35932 37294 35934 37346
rect 35934 37294 35986 37346
rect 35986 37294 35988 37346
rect 35932 37292 35988 37294
rect 36092 37346 36148 37348
rect 36092 37294 36094 37346
rect 36094 37294 36146 37346
rect 36146 37294 36148 37346
rect 36092 37292 36148 37294
rect 36252 37346 36308 37348
rect 36252 37294 36254 37346
rect 36254 37294 36306 37346
rect 36306 37294 36308 37346
rect 36252 37292 36308 37294
rect 36412 37346 36468 37348
rect 36412 37294 36414 37346
rect 36414 37294 36466 37346
rect 36466 37294 36468 37346
rect 36412 37292 36468 37294
rect 36572 37346 36628 37348
rect 36572 37294 36574 37346
rect 36574 37294 36626 37346
rect 36626 37294 36628 37346
rect 36572 37292 36628 37294
rect 36732 37346 36788 37348
rect 36732 37294 36734 37346
rect 36734 37294 36786 37346
rect 36786 37294 36788 37346
rect 36732 37292 36788 37294
rect 36892 37346 36948 37348
rect 36892 37294 36894 37346
rect 36894 37294 36946 37346
rect 36946 37294 36948 37346
rect 36892 37292 36948 37294
rect 37052 37346 37108 37348
rect 37052 37294 37054 37346
rect 37054 37294 37106 37346
rect 37106 37294 37108 37346
rect 37052 37292 37108 37294
rect 37212 37346 37268 37348
rect 37212 37294 37214 37346
rect 37214 37294 37266 37346
rect 37266 37294 37268 37346
rect 37212 37292 37268 37294
rect 37372 37346 37428 37348
rect 37372 37294 37374 37346
rect 37374 37294 37426 37346
rect 37426 37294 37428 37346
rect 37372 37292 37428 37294
rect 37532 37346 37588 37348
rect 37532 37294 37534 37346
rect 37534 37294 37586 37346
rect 37586 37294 37588 37346
rect 37532 37292 37588 37294
rect 37692 37346 37748 37348
rect 37692 37294 37694 37346
rect 37694 37294 37746 37346
rect 37746 37294 37748 37346
rect 37692 37292 37748 37294
rect 37852 37346 37908 37348
rect 37852 37294 37854 37346
rect 37854 37294 37906 37346
rect 37906 37294 37908 37346
rect 37852 37292 37908 37294
rect 38012 37346 38068 37348
rect 38012 37294 38014 37346
rect 38014 37294 38066 37346
rect 38066 37294 38068 37346
rect 38012 37292 38068 37294
rect 38172 37346 38228 37348
rect 38172 37294 38174 37346
rect 38174 37294 38226 37346
rect 38226 37294 38228 37346
rect 38172 37292 38228 37294
rect 38332 37346 38388 37348
rect 38332 37294 38334 37346
rect 38334 37294 38386 37346
rect 38386 37294 38388 37346
rect 38332 37292 38388 37294
rect 38492 37346 38548 37348
rect 38492 37294 38494 37346
rect 38494 37294 38546 37346
rect 38546 37294 38548 37346
rect 38492 37292 38548 37294
rect 38652 37346 38708 37348
rect 38652 37294 38654 37346
rect 38654 37294 38706 37346
rect 38706 37294 38708 37346
rect 38652 37292 38708 37294
rect 38812 37346 38868 37348
rect 38812 37294 38814 37346
rect 38814 37294 38866 37346
rect 38866 37294 38868 37346
rect 38812 37292 38868 37294
rect 38972 37346 39028 37348
rect 38972 37294 38974 37346
rect 38974 37294 39026 37346
rect 39026 37294 39028 37346
rect 38972 37292 39028 37294
rect 39132 37346 39188 37348
rect 39132 37294 39134 37346
rect 39134 37294 39186 37346
rect 39186 37294 39188 37346
rect 39132 37292 39188 37294
rect 39292 37346 39348 37348
rect 39292 37294 39294 37346
rect 39294 37294 39346 37346
rect 39346 37294 39348 37346
rect 39292 37292 39348 37294
rect 39452 37346 39508 37348
rect 39452 37294 39454 37346
rect 39454 37294 39506 37346
rect 39506 37294 39508 37346
rect 39452 37292 39508 37294
rect 39612 37346 39668 37348
rect 39612 37294 39614 37346
rect 39614 37294 39666 37346
rect 39666 37294 39668 37346
rect 39612 37292 39668 37294
rect 39772 37346 39828 37348
rect 39772 37294 39774 37346
rect 39774 37294 39826 37346
rect 39826 37294 39828 37346
rect 39772 37292 39828 37294
rect 39932 37346 39988 37348
rect 39932 37294 39934 37346
rect 39934 37294 39986 37346
rect 39986 37294 39988 37346
rect 39932 37292 39988 37294
rect 40092 37346 40148 37348
rect 40092 37294 40094 37346
rect 40094 37294 40146 37346
rect 40146 37294 40148 37346
rect 40092 37292 40148 37294
rect 40252 37346 40308 37348
rect 40252 37294 40254 37346
rect 40254 37294 40306 37346
rect 40306 37294 40308 37346
rect 40252 37292 40308 37294
rect 40412 37346 40468 37348
rect 40412 37294 40414 37346
rect 40414 37294 40466 37346
rect 40466 37294 40468 37346
rect 40412 37292 40468 37294
rect 40572 37346 40628 37348
rect 40572 37294 40574 37346
rect 40574 37294 40626 37346
rect 40626 37294 40628 37346
rect 40572 37292 40628 37294
rect 40732 37346 40788 37348
rect 40732 37294 40734 37346
rect 40734 37294 40786 37346
rect 40786 37294 40788 37346
rect 40732 37292 40788 37294
rect 40892 37346 40948 37348
rect 40892 37294 40894 37346
rect 40894 37294 40946 37346
rect 40946 37294 40948 37346
rect 40892 37292 40948 37294
rect 41052 37346 41108 37348
rect 41052 37294 41054 37346
rect 41054 37294 41106 37346
rect 41106 37294 41108 37346
rect 41052 37292 41108 37294
rect 41212 37346 41268 37348
rect 41212 37294 41214 37346
rect 41214 37294 41266 37346
rect 41266 37294 41268 37346
rect 41212 37292 41268 37294
rect 41372 37346 41428 37348
rect 41372 37294 41374 37346
rect 41374 37294 41426 37346
rect 41426 37294 41428 37346
rect 41372 37292 41428 37294
rect 41532 37346 41588 37348
rect 41532 37294 41534 37346
rect 41534 37294 41586 37346
rect 41586 37294 41588 37346
rect 41532 37292 41588 37294
rect 41692 37346 41748 37348
rect 41692 37294 41694 37346
rect 41694 37294 41746 37346
rect 41746 37294 41748 37346
rect 41692 37292 41748 37294
rect 41852 37346 41908 37348
rect 41852 37294 41854 37346
rect 41854 37294 41906 37346
rect 41906 37294 41908 37346
rect 41852 37292 41908 37294
rect 8652 37132 8708 37188
rect 22732 37132 22788 37188
rect 33212 37132 33268 37188
rect 12 37026 68 37028
rect 12 36974 14 37026
rect 14 36974 66 37026
rect 66 36974 68 37026
rect 12 36972 68 36974
rect 172 37026 228 37028
rect 172 36974 174 37026
rect 174 36974 226 37026
rect 226 36974 228 37026
rect 172 36972 228 36974
rect 332 37026 388 37028
rect 332 36974 334 37026
rect 334 36974 386 37026
rect 386 36974 388 37026
rect 332 36972 388 36974
rect 492 37026 548 37028
rect 492 36974 494 37026
rect 494 36974 546 37026
rect 546 36974 548 37026
rect 492 36972 548 36974
rect 652 37026 708 37028
rect 652 36974 654 37026
rect 654 36974 706 37026
rect 706 36974 708 37026
rect 652 36972 708 36974
rect 812 37026 868 37028
rect 812 36974 814 37026
rect 814 36974 866 37026
rect 866 36974 868 37026
rect 812 36972 868 36974
rect 972 37026 1028 37028
rect 972 36974 974 37026
rect 974 36974 1026 37026
rect 1026 36974 1028 37026
rect 972 36972 1028 36974
rect 1132 37026 1188 37028
rect 1132 36974 1134 37026
rect 1134 36974 1186 37026
rect 1186 36974 1188 37026
rect 1132 36972 1188 36974
rect 1292 37026 1348 37028
rect 1292 36974 1294 37026
rect 1294 36974 1346 37026
rect 1346 36974 1348 37026
rect 1292 36972 1348 36974
rect 1452 37026 1508 37028
rect 1452 36974 1454 37026
rect 1454 36974 1506 37026
rect 1506 36974 1508 37026
rect 1452 36972 1508 36974
rect 1612 37026 1668 37028
rect 1612 36974 1614 37026
rect 1614 36974 1666 37026
rect 1666 36974 1668 37026
rect 1612 36972 1668 36974
rect 1772 37026 1828 37028
rect 1772 36974 1774 37026
rect 1774 36974 1826 37026
rect 1826 36974 1828 37026
rect 1772 36972 1828 36974
rect 1932 37026 1988 37028
rect 1932 36974 1934 37026
rect 1934 36974 1986 37026
rect 1986 36974 1988 37026
rect 1932 36972 1988 36974
rect 2092 37026 2148 37028
rect 2092 36974 2094 37026
rect 2094 36974 2146 37026
rect 2146 36974 2148 37026
rect 2092 36972 2148 36974
rect 2252 37026 2308 37028
rect 2252 36974 2254 37026
rect 2254 36974 2306 37026
rect 2306 36974 2308 37026
rect 2252 36972 2308 36974
rect 2412 37026 2468 37028
rect 2412 36974 2414 37026
rect 2414 36974 2466 37026
rect 2466 36974 2468 37026
rect 2412 36972 2468 36974
rect 2572 37026 2628 37028
rect 2572 36974 2574 37026
rect 2574 36974 2626 37026
rect 2626 36974 2628 37026
rect 2572 36972 2628 36974
rect 2732 37026 2788 37028
rect 2732 36974 2734 37026
rect 2734 36974 2786 37026
rect 2786 36974 2788 37026
rect 2732 36972 2788 36974
rect 2892 37026 2948 37028
rect 2892 36974 2894 37026
rect 2894 36974 2946 37026
rect 2946 36974 2948 37026
rect 2892 36972 2948 36974
rect 3052 37026 3108 37028
rect 3052 36974 3054 37026
rect 3054 36974 3106 37026
rect 3106 36974 3108 37026
rect 3052 36972 3108 36974
rect 3212 37026 3268 37028
rect 3212 36974 3214 37026
rect 3214 36974 3266 37026
rect 3266 36974 3268 37026
rect 3212 36972 3268 36974
rect 3372 37026 3428 37028
rect 3372 36974 3374 37026
rect 3374 36974 3426 37026
rect 3426 36974 3428 37026
rect 3372 36972 3428 36974
rect 3532 37026 3588 37028
rect 3532 36974 3534 37026
rect 3534 36974 3586 37026
rect 3586 36974 3588 37026
rect 3532 36972 3588 36974
rect 3692 37026 3748 37028
rect 3692 36974 3694 37026
rect 3694 36974 3746 37026
rect 3746 36974 3748 37026
rect 3692 36972 3748 36974
rect 3852 37026 3908 37028
rect 3852 36974 3854 37026
rect 3854 36974 3906 37026
rect 3906 36974 3908 37026
rect 3852 36972 3908 36974
rect 4012 37026 4068 37028
rect 4012 36974 4014 37026
rect 4014 36974 4066 37026
rect 4066 36974 4068 37026
rect 4012 36972 4068 36974
rect 4172 37026 4228 37028
rect 4172 36974 4174 37026
rect 4174 36974 4226 37026
rect 4226 36974 4228 37026
rect 4172 36972 4228 36974
rect 4332 37026 4388 37028
rect 4332 36974 4334 37026
rect 4334 36974 4386 37026
rect 4386 36974 4388 37026
rect 4332 36972 4388 36974
rect 4492 37026 4548 37028
rect 4492 36974 4494 37026
rect 4494 36974 4546 37026
rect 4546 36974 4548 37026
rect 4492 36972 4548 36974
rect 4652 37026 4708 37028
rect 4652 36974 4654 37026
rect 4654 36974 4706 37026
rect 4706 36974 4708 37026
rect 4652 36972 4708 36974
rect 4812 37026 4868 37028
rect 4812 36974 4814 37026
rect 4814 36974 4866 37026
rect 4866 36974 4868 37026
rect 4812 36972 4868 36974
rect 4972 37026 5028 37028
rect 4972 36974 4974 37026
rect 4974 36974 5026 37026
rect 5026 36974 5028 37026
rect 4972 36972 5028 36974
rect 5132 37026 5188 37028
rect 5132 36974 5134 37026
rect 5134 36974 5186 37026
rect 5186 36974 5188 37026
rect 5132 36972 5188 36974
rect 5292 37026 5348 37028
rect 5292 36974 5294 37026
rect 5294 36974 5346 37026
rect 5346 36974 5348 37026
rect 5292 36972 5348 36974
rect 5452 37026 5508 37028
rect 5452 36974 5454 37026
rect 5454 36974 5506 37026
rect 5506 36974 5508 37026
rect 5452 36972 5508 36974
rect 5612 37026 5668 37028
rect 5612 36974 5614 37026
rect 5614 36974 5666 37026
rect 5666 36974 5668 37026
rect 5612 36972 5668 36974
rect 5772 37026 5828 37028
rect 5772 36974 5774 37026
rect 5774 36974 5826 37026
rect 5826 36974 5828 37026
rect 5772 36972 5828 36974
rect 5932 37026 5988 37028
rect 5932 36974 5934 37026
rect 5934 36974 5986 37026
rect 5986 36974 5988 37026
rect 5932 36972 5988 36974
rect 6092 37026 6148 37028
rect 6092 36974 6094 37026
rect 6094 36974 6146 37026
rect 6146 36974 6148 37026
rect 6092 36972 6148 36974
rect 6252 37026 6308 37028
rect 6252 36974 6254 37026
rect 6254 36974 6306 37026
rect 6306 36974 6308 37026
rect 6252 36972 6308 36974
rect 6412 37026 6468 37028
rect 6412 36974 6414 37026
rect 6414 36974 6466 37026
rect 6466 36974 6468 37026
rect 6412 36972 6468 36974
rect 6572 37026 6628 37028
rect 6572 36974 6574 37026
rect 6574 36974 6626 37026
rect 6626 36974 6628 37026
rect 6572 36972 6628 36974
rect 6732 37026 6788 37028
rect 6732 36974 6734 37026
rect 6734 36974 6786 37026
rect 6786 36974 6788 37026
rect 6732 36972 6788 36974
rect 6892 37026 6948 37028
rect 6892 36974 6894 37026
rect 6894 36974 6946 37026
rect 6946 36974 6948 37026
rect 6892 36972 6948 36974
rect 7052 37026 7108 37028
rect 7052 36974 7054 37026
rect 7054 36974 7106 37026
rect 7106 36974 7108 37026
rect 7052 36972 7108 36974
rect 7212 37026 7268 37028
rect 7212 36974 7214 37026
rect 7214 36974 7266 37026
rect 7266 36974 7268 37026
rect 7212 36972 7268 36974
rect 7372 37026 7428 37028
rect 7372 36974 7374 37026
rect 7374 36974 7426 37026
rect 7426 36974 7428 37026
rect 7372 36972 7428 36974
rect 7532 37026 7588 37028
rect 7532 36974 7534 37026
rect 7534 36974 7586 37026
rect 7586 36974 7588 37026
rect 7532 36972 7588 36974
rect 7692 37026 7748 37028
rect 7692 36974 7694 37026
rect 7694 36974 7746 37026
rect 7746 36974 7748 37026
rect 7692 36972 7748 36974
rect 7852 37026 7908 37028
rect 7852 36974 7854 37026
rect 7854 36974 7906 37026
rect 7906 36974 7908 37026
rect 7852 36972 7908 36974
rect 8012 37026 8068 37028
rect 8012 36974 8014 37026
rect 8014 36974 8066 37026
rect 8066 36974 8068 37026
rect 8012 36972 8068 36974
rect 8172 37026 8228 37028
rect 8172 36974 8174 37026
rect 8174 36974 8226 37026
rect 8226 36974 8228 37026
rect 8172 36972 8228 36974
rect 8332 37026 8388 37028
rect 8332 36974 8334 37026
rect 8334 36974 8386 37026
rect 8386 36974 8388 37026
rect 8332 36972 8388 36974
rect 8492 36972 8548 37028
rect 8812 36972 8868 37028
rect 12492 37026 12548 37028
rect 12492 36974 12494 37026
rect 12494 36974 12546 37026
rect 12546 36974 12548 37026
rect 12492 36972 12548 36974
rect 12652 37026 12708 37028
rect 12652 36974 12654 37026
rect 12654 36974 12706 37026
rect 12706 36974 12708 37026
rect 12652 36972 12708 36974
rect 12812 37026 12868 37028
rect 12812 36974 12814 37026
rect 12814 36974 12866 37026
rect 12866 36974 12868 37026
rect 12812 36972 12868 36974
rect 12972 37026 13028 37028
rect 12972 36974 12974 37026
rect 12974 36974 13026 37026
rect 13026 36974 13028 37026
rect 12972 36972 13028 36974
rect 13132 37026 13188 37028
rect 13132 36974 13134 37026
rect 13134 36974 13186 37026
rect 13186 36974 13188 37026
rect 13132 36972 13188 36974
rect 13292 37026 13348 37028
rect 13292 36974 13294 37026
rect 13294 36974 13346 37026
rect 13346 36974 13348 37026
rect 13292 36972 13348 36974
rect 13452 37026 13508 37028
rect 13452 36974 13454 37026
rect 13454 36974 13506 37026
rect 13506 36974 13508 37026
rect 13452 36972 13508 36974
rect 13612 37026 13668 37028
rect 13612 36974 13614 37026
rect 13614 36974 13666 37026
rect 13666 36974 13668 37026
rect 13612 36972 13668 36974
rect 13772 37026 13828 37028
rect 13772 36974 13774 37026
rect 13774 36974 13826 37026
rect 13826 36974 13828 37026
rect 13772 36972 13828 36974
rect 13932 37026 13988 37028
rect 13932 36974 13934 37026
rect 13934 36974 13986 37026
rect 13986 36974 13988 37026
rect 13932 36972 13988 36974
rect 14092 37026 14148 37028
rect 14092 36974 14094 37026
rect 14094 36974 14146 37026
rect 14146 36974 14148 37026
rect 14092 36972 14148 36974
rect 14252 37026 14308 37028
rect 14252 36974 14254 37026
rect 14254 36974 14306 37026
rect 14306 36974 14308 37026
rect 14252 36972 14308 36974
rect 14412 37026 14468 37028
rect 14412 36974 14414 37026
rect 14414 36974 14466 37026
rect 14466 36974 14468 37026
rect 14412 36972 14468 36974
rect 14572 37026 14628 37028
rect 14572 36974 14574 37026
rect 14574 36974 14626 37026
rect 14626 36974 14628 37026
rect 14572 36972 14628 36974
rect 14732 37026 14788 37028
rect 14732 36974 14734 37026
rect 14734 36974 14786 37026
rect 14786 36974 14788 37026
rect 14732 36972 14788 36974
rect 14892 37026 14948 37028
rect 14892 36974 14894 37026
rect 14894 36974 14946 37026
rect 14946 36974 14948 37026
rect 14892 36972 14948 36974
rect 15052 37026 15108 37028
rect 15052 36974 15054 37026
rect 15054 36974 15106 37026
rect 15106 36974 15108 37026
rect 15052 36972 15108 36974
rect 15212 37026 15268 37028
rect 15212 36974 15214 37026
rect 15214 36974 15266 37026
rect 15266 36974 15268 37026
rect 15212 36972 15268 36974
rect 15372 37026 15428 37028
rect 15372 36974 15374 37026
rect 15374 36974 15426 37026
rect 15426 36974 15428 37026
rect 15372 36972 15428 36974
rect 15532 37026 15588 37028
rect 15532 36974 15534 37026
rect 15534 36974 15586 37026
rect 15586 36974 15588 37026
rect 15532 36972 15588 36974
rect 15692 37026 15748 37028
rect 15692 36974 15694 37026
rect 15694 36974 15746 37026
rect 15746 36974 15748 37026
rect 15692 36972 15748 36974
rect 15852 37026 15908 37028
rect 15852 36974 15854 37026
rect 15854 36974 15906 37026
rect 15906 36974 15908 37026
rect 15852 36972 15908 36974
rect 16012 37026 16068 37028
rect 16012 36974 16014 37026
rect 16014 36974 16066 37026
rect 16066 36974 16068 37026
rect 16012 36972 16068 36974
rect 16172 37026 16228 37028
rect 16172 36974 16174 37026
rect 16174 36974 16226 37026
rect 16226 36974 16228 37026
rect 16172 36972 16228 36974
rect 16332 37026 16388 37028
rect 16332 36974 16334 37026
rect 16334 36974 16386 37026
rect 16386 36974 16388 37026
rect 16332 36972 16388 36974
rect 16492 37026 16548 37028
rect 16492 36974 16494 37026
rect 16494 36974 16546 37026
rect 16546 36974 16548 37026
rect 16492 36972 16548 36974
rect 16652 37026 16708 37028
rect 16652 36974 16654 37026
rect 16654 36974 16706 37026
rect 16706 36974 16708 37026
rect 16652 36972 16708 36974
rect 16812 37026 16868 37028
rect 16812 36974 16814 37026
rect 16814 36974 16866 37026
rect 16866 36974 16868 37026
rect 16812 36972 16868 36974
rect 16972 37026 17028 37028
rect 16972 36974 16974 37026
rect 16974 36974 17026 37026
rect 17026 36974 17028 37026
rect 16972 36972 17028 36974
rect 17132 37026 17188 37028
rect 17132 36974 17134 37026
rect 17134 36974 17186 37026
rect 17186 36974 17188 37026
rect 17132 36972 17188 36974
rect 17292 37026 17348 37028
rect 17292 36974 17294 37026
rect 17294 36974 17346 37026
rect 17346 36974 17348 37026
rect 17292 36972 17348 36974
rect 17452 37026 17508 37028
rect 17452 36974 17454 37026
rect 17454 36974 17506 37026
rect 17506 36974 17508 37026
rect 17452 36972 17508 36974
rect 17612 37026 17668 37028
rect 17612 36974 17614 37026
rect 17614 36974 17666 37026
rect 17666 36974 17668 37026
rect 17612 36972 17668 36974
rect 17772 37026 17828 37028
rect 17772 36974 17774 37026
rect 17774 36974 17826 37026
rect 17826 36974 17828 37026
rect 17772 36972 17828 36974
rect 17932 37026 17988 37028
rect 17932 36974 17934 37026
rect 17934 36974 17986 37026
rect 17986 36974 17988 37026
rect 17932 36972 17988 36974
rect 18092 37026 18148 37028
rect 18092 36974 18094 37026
rect 18094 36974 18146 37026
rect 18146 36974 18148 37026
rect 18092 36972 18148 36974
rect 18252 37026 18308 37028
rect 18252 36974 18254 37026
rect 18254 36974 18306 37026
rect 18306 36974 18308 37026
rect 18252 36972 18308 36974
rect 18412 37026 18468 37028
rect 18412 36974 18414 37026
rect 18414 36974 18466 37026
rect 18466 36974 18468 37026
rect 18412 36972 18468 36974
rect 18572 37026 18628 37028
rect 18572 36974 18574 37026
rect 18574 36974 18626 37026
rect 18626 36974 18628 37026
rect 18572 36972 18628 36974
rect 18732 37026 18788 37028
rect 18732 36974 18734 37026
rect 18734 36974 18786 37026
rect 18786 36974 18788 37026
rect 18732 36972 18788 36974
rect 18892 37026 18948 37028
rect 18892 36974 18894 37026
rect 18894 36974 18946 37026
rect 18946 36974 18948 37026
rect 18892 36972 18948 36974
rect 22572 36972 22628 37028
rect 22892 36972 22948 37028
rect 23132 37026 23188 37028
rect 23132 36974 23134 37026
rect 23134 36974 23186 37026
rect 23186 36974 23188 37026
rect 23132 36972 23188 36974
rect 23292 37026 23348 37028
rect 23292 36974 23294 37026
rect 23294 36974 23346 37026
rect 23346 36974 23348 37026
rect 23292 36972 23348 36974
rect 23452 37026 23508 37028
rect 23452 36974 23454 37026
rect 23454 36974 23506 37026
rect 23506 36974 23508 37026
rect 23452 36972 23508 36974
rect 23612 37026 23668 37028
rect 23612 36974 23614 37026
rect 23614 36974 23666 37026
rect 23666 36974 23668 37026
rect 23612 36972 23668 36974
rect 23772 37026 23828 37028
rect 23772 36974 23774 37026
rect 23774 36974 23826 37026
rect 23826 36974 23828 37026
rect 23772 36972 23828 36974
rect 23932 37026 23988 37028
rect 23932 36974 23934 37026
rect 23934 36974 23986 37026
rect 23986 36974 23988 37026
rect 23932 36972 23988 36974
rect 24092 37026 24148 37028
rect 24092 36974 24094 37026
rect 24094 36974 24146 37026
rect 24146 36974 24148 37026
rect 24092 36972 24148 36974
rect 24252 37026 24308 37028
rect 24252 36974 24254 37026
rect 24254 36974 24306 37026
rect 24306 36974 24308 37026
rect 24252 36972 24308 36974
rect 24412 37026 24468 37028
rect 24412 36974 24414 37026
rect 24414 36974 24466 37026
rect 24466 36974 24468 37026
rect 24412 36972 24468 36974
rect 24572 37026 24628 37028
rect 24572 36974 24574 37026
rect 24574 36974 24626 37026
rect 24626 36974 24628 37026
rect 24572 36972 24628 36974
rect 24732 37026 24788 37028
rect 24732 36974 24734 37026
rect 24734 36974 24786 37026
rect 24786 36974 24788 37026
rect 24732 36972 24788 36974
rect 24892 37026 24948 37028
rect 24892 36974 24894 37026
rect 24894 36974 24946 37026
rect 24946 36974 24948 37026
rect 24892 36972 24948 36974
rect 25052 37026 25108 37028
rect 25052 36974 25054 37026
rect 25054 36974 25106 37026
rect 25106 36974 25108 37026
rect 25052 36972 25108 36974
rect 25212 37026 25268 37028
rect 25212 36974 25214 37026
rect 25214 36974 25266 37026
rect 25266 36974 25268 37026
rect 25212 36972 25268 36974
rect 25372 37026 25428 37028
rect 25372 36974 25374 37026
rect 25374 36974 25426 37026
rect 25426 36974 25428 37026
rect 25372 36972 25428 36974
rect 25532 37026 25588 37028
rect 25532 36974 25534 37026
rect 25534 36974 25586 37026
rect 25586 36974 25588 37026
rect 25532 36972 25588 36974
rect 25692 37026 25748 37028
rect 25692 36974 25694 37026
rect 25694 36974 25746 37026
rect 25746 36974 25748 37026
rect 25692 36972 25748 36974
rect 25852 37026 25908 37028
rect 25852 36974 25854 37026
rect 25854 36974 25906 37026
rect 25906 36974 25908 37026
rect 25852 36972 25908 36974
rect 26012 37026 26068 37028
rect 26012 36974 26014 37026
rect 26014 36974 26066 37026
rect 26066 36974 26068 37026
rect 26012 36972 26068 36974
rect 26172 37026 26228 37028
rect 26172 36974 26174 37026
rect 26174 36974 26226 37026
rect 26226 36974 26228 37026
rect 26172 36972 26228 36974
rect 26332 37026 26388 37028
rect 26332 36974 26334 37026
rect 26334 36974 26386 37026
rect 26386 36974 26388 37026
rect 26332 36972 26388 36974
rect 26492 37026 26548 37028
rect 26492 36974 26494 37026
rect 26494 36974 26546 37026
rect 26546 36974 26548 37026
rect 26492 36972 26548 36974
rect 26652 37026 26708 37028
rect 26652 36974 26654 37026
rect 26654 36974 26706 37026
rect 26706 36974 26708 37026
rect 26652 36972 26708 36974
rect 26812 37026 26868 37028
rect 26812 36974 26814 37026
rect 26814 36974 26866 37026
rect 26866 36974 26868 37026
rect 26812 36972 26868 36974
rect 26972 37026 27028 37028
rect 26972 36974 26974 37026
rect 26974 36974 27026 37026
rect 27026 36974 27028 37026
rect 26972 36972 27028 36974
rect 27132 37026 27188 37028
rect 27132 36974 27134 37026
rect 27134 36974 27186 37026
rect 27186 36974 27188 37026
rect 27132 36972 27188 36974
rect 27292 37026 27348 37028
rect 27292 36974 27294 37026
rect 27294 36974 27346 37026
rect 27346 36974 27348 37026
rect 27292 36972 27348 36974
rect 27452 37026 27508 37028
rect 27452 36974 27454 37026
rect 27454 36974 27506 37026
rect 27506 36974 27508 37026
rect 27452 36972 27508 36974
rect 27612 37026 27668 37028
rect 27612 36974 27614 37026
rect 27614 36974 27666 37026
rect 27666 36974 27668 37026
rect 27612 36972 27668 36974
rect 27772 37026 27828 37028
rect 27772 36974 27774 37026
rect 27774 36974 27826 37026
rect 27826 36974 27828 37026
rect 27772 36972 27828 36974
rect 27932 37026 27988 37028
rect 27932 36974 27934 37026
rect 27934 36974 27986 37026
rect 27986 36974 27988 37026
rect 27932 36972 27988 36974
rect 28092 37026 28148 37028
rect 28092 36974 28094 37026
rect 28094 36974 28146 37026
rect 28146 36974 28148 37026
rect 28092 36972 28148 36974
rect 28252 37026 28308 37028
rect 28252 36974 28254 37026
rect 28254 36974 28306 37026
rect 28306 36974 28308 37026
rect 28252 36972 28308 36974
rect 28412 37026 28468 37028
rect 28412 36974 28414 37026
rect 28414 36974 28466 37026
rect 28466 36974 28468 37026
rect 28412 36972 28468 36974
rect 28572 37026 28628 37028
rect 28572 36974 28574 37026
rect 28574 36974 28626 37026
rect 28626 36974 28628 37026
rect 28572 36972 28628 36974
rect 28732 37026 28788 37028
rect 28732 36974 28734 37026
rect 28734 36974 28786 37026
rect 28786 36974 28788 37026
rect 28732 36972 28788 36974
rect 28892 37026 28948 37028
rect 28892 36974 28894 37026
rect 28894 36974 28946 37026
rect 28946 36974 28948 37026
rect 28892 36972 28948 36974
rect 29052 37026 29108 37028
rect 29052 36974 29054 37026
rect 29054 36974 29106 37026
rect 29106 36974 29108 37026
rect 29052 36972 29108 36974
rect 29212 37026 29268 37028
rect 29212 36974 29214 37026
rect 29214 36974 29266 37026
rect 29266 36974 29268 37026
rect 29212 36972 29268 36974
rect 29372 37026 29428 37028
rect 29372 36974 29374 37026
rect 29374 36974 29426 37026
rect 29426 36974 29428 37026
rect 29372 36972 29428 36974
rect 33052 36972 33108 37028
rect 33372 36972 33428 37028
rect 33532 37026 33588 37028
rect 33532 36974 33534 37026
rect 33534 36974 33586 37026
rect 33586 36974 33588 37026
rect 33532 36972 33588 36974
rect 33692 37026 33748 37028
rect 33692 36974 33694 37026
rect 33694 36974 33746 37026
rect 33746 36974 33748 37026
rect 33692 36972 33748 36974
rect 33852 37026 33908 37028
rect 33852 36974 33854 37026
rect 33854 36974 33906 37026
rect 33906 36974 33908 37026
rect 33852 36972 33908 36974
rect 34012 37026 34068 37028
rect 34012 36974 34014 37026
rect 34014 36974 34066 37026
rect 34066 36974 34068 37026
rect 34012 36972 34068 36974
rect 34172 37026 34228 37028
rect 34172 36974 34174 37026
rect 34174 36974 34226 37026
rect 34226 36974 34228 37026
rect 34172 36972 34228 36974
rect 34332 37026 34388 37028
rect 34332 36974 34334 37026
rect 34334 36974 34386 37026
rect 34386 36974 34388 37026
rect 34332 36972 34388 36974
rect 34492 37026 34548 37028
rect 34492 36974 34494 37026
rect 34494 36974 34546 37026
rect 34546 36974 34548 37026
rect 34492 36972 34548 36974
rect 34652 37026 34708 37028
rect 34652 36974 34654 37026
rect 34654 36974 34706 37026
rect 34706 36974 34708 37026
rect 34652 36972 34708 36974
rect 34812 37026 34868 37028
rect 34812 36974 34814 37026
rect 34814 36974 34866 37026
rect 34866 36974 34868 37026
rect 34812 36972 34868 36974
rect 34972 37026 35028 37028
rect 34972 36974 34974 37026
rect 34974 36974 35026 37026
rect 35026 36974 35028 37026
rect 34972 36972 35028 36974
rect 35132 37026 35188 37028
rect 35132 36974 35134 37026
rect 35134 36974 35186 37026
rect 35186 36974 35188 37026
rect 35132 36972 35188 36974
rect 35292 37026 35348 37028
rect 35292 36974 35294 37026
rect 35294 36974 35346 37026
rect 35346 36974 35348 37026
rect 35292 36972 35348 36974
rect 35452 37026 35508 37028
rect 35452 36974 35454 37026
rect 35454 36974 35506 37026
rect 35506 36974 35508 37026
rect 35452 36972 35508 36974
rect 35612 37026 35668 37028
rect 35612 36974 35614 37026
rect 35614 36974 35666 37026
rect 35666 36974 35668 37026
rect 35612 36972 35668 36974
rect 35772 37026 35828 37028
rect 35772 36974 35774 37026
rect 35774 36974 35826 37026
rect 35826 36974 35828 37026
rect 35772 36972 35828 36974
rect 35932 37026 35988 37028
rect 35932 36974 35934 37026
rect 35934 36974 35986 37026
rect 35986 36974 35988 37026
rect 35932 36972 35988 36974
rect 36092 37026 36148 37028
rect 36092 36974 36094 37026
rect 36094 36974 36146 37026
rect 36146 36974 36148 37026
rect 36092 36972 36148 36974
rect 36252 37026 36308 37028
rect 36252 36974 36254 37026
rect 36254 36974 36306 37026
rect 36306 36974 36308 37026
rect 36252 36972 36308 36974
rect 36412 37026 36468 37028
rect 36412 36974 36414 37026
rect 36414 36974 36466 37026
rect 36466 36974 36468 37026
rect 36412 36972 36468 36974
rect 36572 37026 36628 37028
rect 36572 36974 36574 37026
rect 36574 36974 36626 37026
rect 36626 36974 36628 37026
rect 36572 36972 36628 36974
rect 36732 37026 36788 37028
rect 36732 36974 36734 37026
rect 36734 36974 36786 37026
rect 36786 36974 36788 37026
rect 36732 36972 36788 36974
rect 36892 37026 36948 37028
rect 36892 36974 36894 37026
rect 36894 36974 36946 37026
rect 36946 36974 36948 37026
rect 36892 36972 36948 36974
rect 37052 37026 37108 37028
rect 37052 36974 37054 37026
rect 37054 36974 37106 37026
rect 37106 36974 37108 37026
rect 37052 36972 37108 36974
rect 37212 37026 37268 37028
rect 37212 36974 37214 37026
rect 37214 36974 37266 37026
rect 37266 36974 37268 37026
rect 37212 36972 37268 36974
rect 37372 37026 37428 37028
rect 37372 36974 37374 37026
rect 37374 36974 37426 37026
rect 37426 36974 37428 37026
rect 37372 36972 37428 36974
rect 37532 37026 37588 37028
rect 37532 36974 37534 37026
rect 37534 36974 37586 37026
rect 37586 36974 37588 37026
rect 37532 36972 37588 36974
rect 37692 37026 37748 37028
rect 37692 36974 37694 37026
rect 37694 36974 37746 37026
rect 37746 36974 37748 37026
rect 37692 36972 37748 36974
rect 37852 37026 37908 37028
rect 37852 36974 37854 37026
rect 37854 36974 37906 37026
rect 37906 36974 37908 37026
rect 37852 36972 37908 36974
rect 38012 37026 38068 37028
rect 38012 36974 38014 37026
rect 38014 36974 38066 37026
rect 38066 36974 38068 37026
rect 38012 36972 38068 36974
rect 38172 37026 38228 37028
rect 38172 36974 38174 37026
rect 38174 36974 38226 37026
rect 38226 36974 38228 37026
rect 38172 36972 38228 36974
rect 38332 37026 38388 37028
rect 38332 36974 38334 37026
rect 38334 36974 38386 37026
rect 38386 36974 38388 37026
rect 38332 36972 38388 36974
rect 38492 37026 38548 37028
rect 38492 36974 38494 37026
rect 38494 36974 38546 37026
rect 38546 36974 38548 37026
rect 38492 36972 38548 36974
rect 38652 37026 38708 37028
rect 38652 36974 38654 37026
rect 38654 36974 38706 37026
rect 38706 36974 38708 37026
rect 38652 36972 38708 36974
rect 38812 37026 38868 37028
rect 38812 36974 38814 37026
rect 38814 36974 38866 37026
rect 38866 36974 38868 37026
rect 38812 36972 38868 36974
rect 38972 37026 39028 37028
rect 38972 36974 38974 37026
rect 38974 36974 39026 37026
rect 39026 36974 39028 37026
rect 38972 36972 39028 36974
rect 39132 37026 39188 37028
rect 39132 36974 39134 37026
rect 39134 36974 39186 37026
rect 39186 36974 39188 37026
rect 39132 36972 39188 36974
rect 39292 37026 39348 37028
rect 39292 36974 39294 37026
rect 39294 36974 39346 37026
rect 39346 36974 39348 37026
rect 39292 36972 39348 36974
rect 39452 37026 39508 37028
rect 39452 36974 39454 37026
rect 39454 36974 39506 37026
rect 39506 36974 39508 37026
rect 39452 36972 39508 36974
rect 39612 37026 39668 37028
rect 39612 36974 39614 37026
rect 39614 36974 39666 37026
rect 39666 36974 39668 37026
rect 39612 36972 39668 36974
rect 39772 37026 39828 37028
rect 39772 36974 39774 37026
rect 39774 36974 39826 37026
rect 39826 36974 39828 37026
rect 39772 36972 39828 36974
rect 39932 37026 39988 37028
rect 39932 36974 39934 37026
rect 39934 36974 39986 37026
rect 39986 36974 39988 37026
rect 39932 36972 39988 36974
rect 40092 37026 40148 37028
rect 40092 36974 40094 37026
rect 40094 36974 40146 37026
rect 40146 36974 40148 37026
rect 40092 36972 40148 36974
rect 40252 37026 40308 37028
rect 40252 36974 40254 37026
rect 40254 36974 40306 37026
rect 40306 36974 40308 37026
rect 40252 36972 40308 36974
rect 40412 37026 40468 37028
rect 40412 36974 40414 37026
rect 40414 36974 40466 37026
rect 40466 36974 40468 37026
rect 40412 36972 40468 36974
rect 40572 37026 40628 37028
rect 40572 36974 40574 37026
rect 40574 36974 40626 37026
rect 40626 36974 40628 37026
rect 40572 36972 40628 36974
rect 40732 37026 40788 37028
rect 40732 36974 40734 37026
rect 40734 36974 40786 37026
rect 40786 36974 40788 37026
rect 40732 36972 40788 36974
rect 40892 37026 40948 37028
rect 40892 36974 40894 37026
rect 40894 36974 40946 37026
rect 40946 36974 40948 37026
rect 40892 36972 40948 36974
rect 41052 37026 41108 37028
rect 41052 36974 41054 37026
rect 41054 36974 41106 37026
rect 41106 36974 41108 37026
rect 41052 36972 41108 36974
rect 41212 37026 41268 37028
rect 41212 36974 41214 37026
rect 41214 36974 41266 37026
rect 41266 36974 41268 37026
rect 41212 36972 41268 36974
rect 41372 37026 41428 37028
rect 41372 36974 41374 37026
rect 41374 36974 41426 37026
rect 41426 36974 41428 37026
rect 41372 36972 41428 36974
rect 41532 37026 41588 37028
rect 41532 36974 41534 37026
rect 41534 36974 41586 37026
rect 41586 36974 41588 37026
rect 41532 36972 41588 36974
rect 41692 37026 41748 37028
rect 41692 36974 41694 37026
rect 41694 36974 41746 37026
rect 41746 36974 41748 37026
rect 41692 36972 41748 36974
rect 41852 37026 41908 37028
rect 41852 36974 41854 37026
rect 41854 36974 41906 37026
rect 41906 36974 41908 37026
rect 41852 36972 41908 36974
rect 12 36866 68 36868
rect 12 36814 14 36866
rect 14 36814 66 36866
rect 66 36814 68 36866
rect 12 36812 68 36814
rect 172 36866 228 36868
rect 172 36814 174 36866
rect 174 36814 226 36866
rect 226 36814 228 36866
rect 172 36812 228 36814
rect 332 36866 388 36868
rect 332 36814 334 36866
rect 334 36814 386 36866
rect 386 36814 388 36866
rect 332 36812 388 36814
rect 492 36866 548 36868
rect 492 36814 494 36866
rect 494 36814 546 36866
rect 546 36814 548 36866
rect 492 36812 548 36814
rect 652 36866 708 36868
rect 652 36814 654 36866
rect 654 36814 706 36866
rect 706 36814 708 36866
rect 652 36812 708 36814
rect 812 36866 868 36868
rect 812 36814 814 36866
rect 814 36814 866 36866
rect 866 36814 868 36866
rect 812 36812 868 36814
rect 972 36866 1028 36868
rect 972 36814 974 36866
rect 974 36814 1026 36866
rect 1026 36814 1028 36866
rect 972 36812 1028 36814
rect 1132 36866 1188 36868
rect 1132 36814 1134 36866
rect 1134 36814 1186 36866
rect 1186 36814 1188 36866
rect 1132 36812 1188 36814
rect 1292 36866 1348 36868
rect 1292 36814 1294 36866
rect 1294 36814 1346 36866
rect 1346 36814 1348 36866
rect 1292 36812 1348 36814
rect 1452 36866 1508 36868
rect 1452 36814 1454 36866
rect 1454 36814 1506 36866
rect 1506 36814 1508 36866
rect 1452 36812 1508 36814
rect 1612 36866 1668 36868
rect 1612 36814 1614 36866
rect 1614 36814 1666 36866
rect 1666 36814 1668 36866
rect 1612 36812 1668 36814
rect 1772 36866 1828 36868
rect 1772 36814 1774 36866
rect 1774 36814 1826 36866
rect 1826 36814 1828 36866
rect 1772 36812 1828 36814
rect 1932 36866 1988 36868
rect 1932 36814 1934 36866
rect 1934 36814 1986 36866
rect 1986 36814 1988 36866
rect 1932 36812 1988 36814
rect 2092 36866 2148 36868
rect 2092 36814 2094 36866
rect 2094 36814 2146 36866
rect 2146 36814 2148 36866
rect 2092 36812 2148 36814
rect 2252 36866 2308 36868
rect 2252 36814 2254 36866
rect 2254 36814 2306 36866
rect 2306 36814 2308 36866
rect 2252 36812 2308 36814
rect 2412 36866 2468 36868
rect 2412 36814 2414 36866
rect 2414 36814 2466 36866
rect 2466 36814 2468 36866
rect 2412 36812 2468 36814
rect 2572 36866 2628 36868
rect 2572 36814 2574 36866
rect 2574 36814 2626 36866
rect 2626 36814 2628 36866
rect 2572 36812 2628 36814
rect 2732 36866 2788 36868
rect 2732 36814 2734 36866
rect 2734 36814 2786 36866
rect 2786 36814 2788 36866
rect 2732 36812 2788 36814
rect 2892 36866 2948 36868
rect 2892 36814 2894 36866
rect 2894 36814 2946 36866
rect 2946 36814 2948 36866
rect 2892 36812 2948 36814
rect 3052 36866 3108 36868
rect 3052 36814 3054 36866
rect 3054 36814 3106 36866
rect 3106 36814 3108 36866
rect 3052 36812 3108 36814
rect 3212 36866 3268 36868
rect 3212 36814 3214 36866
rect 3214 36814 3266 36866
rect 3266 36814 3268 36866
rect 3212 36812 3268 36814
rect 3372 36866 3428 36868
rect 3372 36814 3374 36866
rect 3374 36814 3426 36866
rect 3426 36814 3428 36866
rect 3372 36812 3428 36814
rect 3532 36866 3588 36868
rect 3532 36814 3534 36866
rect 3534 36814 3586 36866
rect 3586 36814 3588 36866
rect 3532 36812 3588 36814
rect 3692 36866 3748 36868
rect 3692 36814 3694 36866
rect 3694 36814 3746 36866
rect 3746 36814 3748 36866
rect 3692 36812 3748 36814
rect 3852 36866 3908 36868
rect 3852 36814 3854 36866
rect 3854 36814 3906 36866
rect 3906 36814 3908 36866
rect 3852 36812 3908 36814
rect 4012 36866 4068 36868
rect 4012 36814 4014 36866
rect 4014 36814 4066 36866
rect 4066 36814 4068 36866
rect 4012 36812 4068 36814
rect 4172 36866 4228 36868
rect 4172 36814 4174 36866
rect 4174 36814 4226 36866
rect 4226 36814 4228 36866
rect 4172 36812 4228 36814
rect 4332 36866 4388 36868
rect 4332 36814 4334 36866
rect 4334 36814 4386 36866
rect 4386 36814 4388 36866
rect 4332 36812 4388 36814
rect 4492 36866 4548 36868
rect 4492 36814 4494 36866
rect 4494 36814 4546 36866
rect 4546 36814 4548 36866
rect 4492 36812 4548 36814
rect 4652 36866 4708 36868
rect 4652 36814 4654 36866
rect 4654 36814 4706 36866
rect 4706 36814 4708 36866
rect 4652 36812 4708 36814
rect 4812 36866 4868 36868
rect 4812 36814 4814 36866
rect 4814 36814 4866 36866
rect 4866 36814 4868 36866
rect 4812 36812 4868 36814
rect 4972 36866 5028 36868
rect 4972 36814 4974 36866
rect 4974 36814 5026 36866
rect 5026 36814 5028 36866
rect 4972 36812 5028 36814
rect 5132 36866 5188 36868
rect 5132 36814 5134 36866
rect 5134 36814 5186 36866
rect 5186 36814 5188 36866
rect 5132 36812 5188 36814
rect 5292 36866 5348 36868
rect 5292 36814 5294 36866
rect 5294 36814 5346 36866
rect 5346 36814 5348 36866
rect 5292 36812 5348 36814
rect 5452 36866 5508 36868
rect 5452 36814 5454 36866
rect 5454 36814 5506 36866
rect 5506 36814 5508 36866
rect 5452 36812 5508 36814
rect 5612 36866 5668 36868
rect 5612 36814 5614 36866
rect 5614 36814 5666 36866
rect 5666 36814 5668 36866
rect 5612 36812 5668 36814
rect 5772 36866 5828 36868
rect 5772 36814 5774 36866
rect 5774 36814 5826 36866
rect 5826 36814 5828 36866
rect 5772 36812 5828 36814
rect 5932 36866 5988 36868
rect 5932 36814 5934 36866
rect 5934 36814 5986 36866
rect 5986 36814 5988 36866
rect 5932 36812 5988 36814
rect 6092 36866 6148 36868
rect 6092 36814 6094 36866
rect 6094 36814 6146 36866
rect 6146 36814 6148 36866
rect 6092 36812 6148 36814
rect 6252 36866 6308 36868
rect 6252 36814 6254 36866
rect 6254 36814 6306 36866
rect 6306 36814 6308 36866
rect 6252 36812 6308 36814
rect 6412 36866 6468 36868
rect 6412 36814 6414 36866
rect 6414 36814 6466 36866
rect 6466 36814 6468 36866
rect 6412 36812 6468 36814
rect 6572 36866 6628 36868
rect 6572 36814 6574 36866
rect 6574 36814 6626 36866
rect 6626 36814 6628 36866
rect 6572 36812 6628 36814
rect 6732 36866 6788 36868
rect 6732 36814 6734 36866
rect 6734 36814 6786 36866
rect 6786 36814 6788 36866
rect 6732 36812 6788 36814
rect 6892 36866 6948 36868
rect 6892 36814 6894 36866
rect 6894 36814 6946 36866
rect 6946 36814 6948 36866
rect 6892 36812 6948 36814
rect 7052 36866 7108 36868
rect 7052 36814 7054 36866
rect 7054 36814 7106 36866
rect 7106 36814 7108 36866
rect 7052 36812 7108 36814
rect 7212 36866 7268 36868
rect 7212 36814 7214 36866
rect 7214 36814 7266 36866
rect 7266 36814 7268 36866
rect 7212 36812 7268 36814
rect 7372 36866 7428 36868
rect 7372 36814 7374 36866
rect 7374 36814 7426 36866
rect 7426 36814 7428 36866
rect 7372 36812 7428 36814
rect 7532 36866 7588 36868
rect 7532 36814 7534 36866
rect 7534 36814 7586 36866
rect 7586 36814 7588 36866
rect 7532 36812 7588 36814
rect 7692 36866 7748 36868
rect 7692 36814 7694 36866
rect 7694 36814 7746 36866
rect 7746 36814 7748 36866
rect 7692 36812 7748 36814
rect 7852 36866 7908 36868
rect 7852 36814 7854 36866
rect 7854 36814 7906 36866
rect 7906 36814 7908 36866
rect 7852 36812 7908 36814
rect 8012 36866 8068 36868
rect 8012 36814 8014 36866
rect 8014 36814 8066 36866
rect 8066 36814 8068 36866
rect 8012 36812 8068 36814
rect 8172 36866 8228 36868
rect 8172 36814 8174 36866
rect 8174 36814 8226 36866
rect 8226 36814 8228 36866
rect 8172 36812 8228 36814
rect 8332 36866 8388 36868
rect 8332 36814 8334 36866
rect 8334 36814 8386 36866
rect 8386 36814 8388 36866
rect 8332 36812 8388 36814
rect 8972 36812 9028 36868
rect 9292 36812 9348 36868
rect 12492 36866 12548 36868
rect 12492 36814 12494 36866
rect 12494 36814 12546 36866
rect 12546 36814 12548 36866
rect 12492 36812 12548 36814
rect 12652 36866 12708 36868
rect 12652 36814 12654 36866
rect 12654 36814 12706 36866
rect 12706 36814 12708 36866
rect 12652 36812 12708 36814
rect 12812 36866 12868 36868
rect 12812 36814 12814 36866
rect 12814 36814 12866 36866
rect 12866 36814 12868 36866
rect 12812 36812 12868 36814
rect 12972 36866 13028 36868
rect 12972 36814 12974 36866
rect 12974 36814 13026 36866
rect 13026 36814 13028 36866
rect 12972 36812 13028 36814
rect 13132 36866 13188 36868
rect 13132 36814 13134 36866
rect 13134 36814 13186 36866
rect 13186 36814 13188 36866
rect 13132 36812 13188 36814
rect 13292 36866 13348 36868
rect 13292 36814 13294 36866
rect 13294 36814 13346 36866
rect 13346 36814 13348 36866
rect 13292 36812 13348 36814
rect 13452 36866 13508 36868
rect 13452 36814 13454 36866
rect 13454 36814 13506 36866
rect 13506 36814 13508 36866
rect 13452 36812 13508 36814
rect 13612 36866 13668 36868
rect 13612 36814 13614 36866
rect 13614 36814 13666 36866
rect 13666 36814 13668 36866
rect 13612 36812 13668 36814
rect 13772 36866 13828 36868
rect 13772 36814 13774 36866
rect 13774 36814 13826 36866
rect 13826 36814 13828 36866
rect 13772 36812 13828 36814
rect 13932 36866 13988 36868
rect 13932 36814 13934 36866
rect 13934 36814 13986 36866
rect 13986 36814 13988 36866
rect 13932 36812 13988 36814
rect 14092 36866 14148 36868
rect 14092 36814 14094 36866
rect 14094 36814 14146 36866
rect 14146 36814 14148 36866
rect 14092 36812 14148 36814
rect 14252 36866 14308 36868
rect 14252 36814 14254 36866
rect 14254 36814 14306 36866
rect 14306 36814 14308 36866
rect 14252 36812 14308 36814
rect 14412 36866 14468 36868
rect 14412 36814 14414 36866
rect 14414 36814 14466 36866
rect 14466 36814 14468 36866
rect 14412 36812 14468 36814
rect 14572 36866 14628 36868
rect 14572 36814 14574 36866
rect 14574 36814 14626 36866
rect 14626 36814 14628 36866
rect 14572 36812 14628 36814
rect 14732 36866 14788 36868
rect 14732 36814 14734 36866
rect 14734 36814 14786 36866
rect 14786 36814 14788 36866
rect 14732 36812 14788 36814
rect 14892 36866 14948 36868
rect 14892 36814 14894 36866
rect 14894 36814 14946 36866
rect 14946 36814 14948 36866
rect 14892 36812 14948 36814
rect 15052 36866 15108 36868
rect 15052 36814 15054 36866
rect 15054 36814 15106 36866
rect 15106 36814 15108 36866
rect 15052 36812 15108 36814
rect 15212 36866 15268 36868
rect 15212 36814 15214 36866
rect 15214 36814 15266 36866
rect 15266 36814 15268 36866
rect 15212 36812 15268 36814
rect 15372 36866 15428 36868
rect 15372 36814 15374 36866
rect 15374 36814 15426 36866
rect 15426 36814 15428 36866
rect 15372 36812 15428 36814
rect 15532 36866 15588 36868
rect 15532 36814 15534 36866
rect 15534 36814 15586 36866
rect 15586 36814 15588 36866
rect 15532 36812 15588 36814
rect 15692 36866 15748 36868
rect 15692 36814 15694 36866
rect 15694 36814 15746 36866
rect 15746 36814 15748 36866
rect 15692 36812 15748 36814
rect 15852 36866 15908 36868
rect 15852 36814 15854 36866
rect 15854 36814 15906 36866
rect 15906 36814 15908 36866
rect 15852 36812 15908 36814
rect 16012 36866 16068 36868
rect 16012 36814 16014 36866
rect 16014 36814 16066 36866
rect 16066 36814 16068 36866
rect 16012 36812 16068 36814
rect 16172 36866 16228 36868
rect 16172 36814 16174 36866
rect 16174 36814 16226 36866
rect 16226 36814 16228 36866
rect 16172 36812 16228 36814
rect 16332 36866 16388 36868
rect 16332 36814 16334 36866
rect 16334 36814 16386 36866
rect 16386 36814 16388 36866
rect 16332 36812 16388 36814
rect 16492 36866 16548 36868
rect 16492 36814 16494 36866
rect 16494 36814 16546 36866
rect 16546 36814 16548 36866
rect 16492 36812 16548 36814
rect 16652 36866 16708 36868
rect 16652 36814 16654 36866
rect 16654 36814 16706 36866
rect 16706 36814 16708 36866
rect 16652 36812 16708 36814
rect 16812 36866 16868 36868
rect 16812 36814 16814 36866
rect 16814 36814 16866 36866
rect 16866 36814 16868 36866
rect 16812 36812 16868 36814
rect 16972 36866 17028 36868
rect 16972 36814 16974 36866
rect 16974 36814 17026 36866
rect 17026 36814 17028 36866
rect 16972 36812 17028 36814
rect 17132 36866 17188 36868
rect 17132 36814 17134 36866
rect 17134 36814 17186 36866
rect 17186 36814 17188 36866
rect 17132 36812 17188 36814
rect 17292 36866 17348 36868
rect 17292 36814 17294 36866
rect 17294 36814 17346 36866
rect 17346 36814 17348 36866
rect 17292 36812 17348 36814
rect 17452 36866 17508 36868
rect 17452 36814 17454 36866
rect 17454 36814 17506 36866
rect 17506 36814 17508 36866
rect 17452 36812 17508 36814
rect 17612 36866 17668 36868
rect 17612 36814 17614 36866
rect 17614 36814 17666 36866
rect 17666 36814 17668 36866
rect 17612 36812 17668 36814
rect 17772 36866 17828 36868
rect 17772 36814 17774 36866
rect 17774 36814 17826 36866
rect 17826 36814 17828 36866
rect 17772 36812 17828 36814
rect 17932 36866 17988 36868
rect 17932 36814 17934 36866
rect 17934 36814 17986 36866
rect 17986 36814 17988 36866
rect 17932 36812 17988 36814
rect 18092 36866 18148 36868
rect 18092 36814 18094 36866
rect 18094 36814 18146 36866
rect 18146 36814 18148 36866
rect 18092 36812 18148 36814
rect 18252 36866 18308 36868
rect 18252 36814 18254 36866
rect 18254 36814 18306 36866
rect 18306 36814 18308 36866
rect 18252 36812 18308 36814
rect 18412 36866 18468 36868
rect 18412 36814 18414 36866
rect 18414 36814 18466 36866
rect 18466 36814 18468 36866
rect 18412 36812 18468 36814
rect 18572 36866 18628 36868
rect 18572 36814 18574 36866
rect 18574 36814 18626 36866
rect 18626 36814 18628 36866
rect 18572 36812 18628 36814
rect 18732 36866 18788 36868
rect 18732 36814 18734 36866
rect 18734 36814 18786 36866
rect 18786 36814 18788 36866
rect 18732 36812 18788 36814
rect 18892 36866 18948 36868
rect 18892 36814 18894 36866
rect 18894 36814 18946 36866
rect 18946 36814 18948 36866
rect 18892 36812 18948 36814
rect 22092 36812 22148 36868
rect 22412 36812 22468 36868
rect 23132 36866 23188 36868
rect 23132 36814 23134 36866
rect 23134 36814 23186 36866
rect 23186 36814 23188 36866
rect 23132 36812 23188 36814
rect 23292 36866 23348 36868
rect 23292 36814 23294 36866
rect 23294 36814 23346 36866
rect 23346 36814 23348 36866
rect 23292 36812 23348 36814
rect 23452 36866 23508 36868
rect 23452 36814 23454 36866
rect 23454 36814 23506 36866
rect 23506 36814 23508 36866
rect 23452 36812 23508 36814
rect 23612 36866 23668 36868
rect 23612 36814 23614 36866
rect 23614 36814 23666 36866
rect 23666 36814 23668 36866
rect 23612 36812 23668 36814
rect 23772 36866 23828 36868
rect 23772 36814 23774 36866
rect 23774 36814 23826 36866
rect 23826 36814 23828 36866
rect 23772 36812 23828 36814
rect 23932 36866 23988 36868
rect 23932 36814 23934 36866
rect 23934 36814 23986 36866
rect 23986 36814 23988 36866
rect 23932 36812 23988 36814
rect 24092 36866 24148 36868
rect 24092 36814 24094 36866
rect 24094 36814 24146 36866
rect 24146 36814 24148 36866
rect 24092 36812 24148 36814
rect 24252 36866 24308 36868
rect 24252 36814 24254 36866
rect 24254 36814 24306 36866
rect 24306 36814 24308 36866
rect 24252 36812 24308 36814
rect 24412 36866 24468 36868
rect 24412 36814 24414 36866
rect 24414 36814 24466 36866
rect 24466 36814 24468 36866
rect 24412 36812 24468 36814
rect 24572 36866 24628 36868
rect 24572 36814 24574 36866
rect 24574 36814 24626 36866
rect 24626 36814 24628 36866
rect 24572 36812 24628 36814
rect 24732 36866 24788 36868
rect 24732 36814 24734 36866
rect 24734 36814 24786 36866
rect 24786 36814 24788 36866
rect 24732 36812 24788 36814
rect 24892 36866 24948 36868
rect 24892 36814 24894 36866
rect 24894 36814 24946 36866
rect 24946 36814 24948 36866
rect 24892 36812 24948 36814
rect 25052 36866 25108 36868
rect 25052 36814 25054 36866
rect 25054 36814 25106 36866
rect 25106 36814 25108 36866
rect 25052 36812 25108 36814
rect 25212 36866 25268 36868
rect 25212 36814 25214 36866
rect 25214 36814 25266 36866
rect 25266 36814 25268 36866
rect 25212 36812 25268 36814
rect 25372 36866 25428 36868
rect 25372 36814 25374 36866
rect 25374 36814 25426 36866
rect 25426 36814 25428 36866
rect 25372 36812 25428 36814
rect 25532 36866 25588 36868
rect 25532 36814 25534 36866
rect 25534 36814 25586 36866
rect 25586 36814 25588 36866
rect 25532 36812 25588 36814
rect 25692 36866 25748 36868
rect 25692 36814 25694 36866
rect 25694 36814 25746 36866
rect 25746 36814 25748 36866
rect 25692 36812 25748 36814
rect 25852 36866 25908 36868
rect 25852 36814 25854 36866
rect 25854 36814 25906 36866
rect 25906 36814 25908 36866
rect 25852 36812 25908 36814
rect 26012 36866 26068 36868
rect 26012 36814 26014 36866
rect 26014 36814 26066 36866
rect 26066 36814 26068 36866
rect 26012 36812 26068 36814
rect 26172 36866 26228 36868
rect 26172 36814 26174 36866
rect 26174 36814 26226 36866
rect 26226 36814 26228 36866
rect 26172 36812 26228 36814
rect 26332 36866 26388 36868
rect 26332 36814 26334 36866
rect 26334 36814 26386 36866
rect 26386 36814 26388 36866
rect 26332 36812 26388 36814
rect 26492 36866 26548 36868
rect 26492 36814 26494 36866
rect 26494 36814 26546 36866
rect 26546 36814 26548 36866
rect 26492 36812 26548 36814
rect 26652 36866 26708 36868
rect 26652 36814 26654 36866
rect 26654 36814 26706 36866
rect 26706 36814 26708 36866
rect 26652 36812 26708 36814
rect 26812 36866 26868 36868
rect 26812 36814 26814 36866
rect 26814 36814 26866 36866
rect 26866 36814 26868 36866
rect 26812 36812 26868 36814
rect 26972 36866 27028 36868
rect 26972 36814 26974 36866
rect 26974 36814 27026 36866
rect 27026 36814 27028 36866
rect 26972 36812 27028 36814
rect 27132 36866 27188 36868
rect 27132 36814 27134 36866
rect 27134 36814 27186 36866
rect 27186 36814 27188 36866
rect 27132 36812 27188 36814
rect 27292 36866 27348 36868
rect 27292 36814 27294 36866
rect 27294 36814 27346 36866
rect 27346 36814 27348 36866
rect 27292 36812 27348 36814
rect 27452 36866 27508 36868
rect 27452 36814 27454 36866
rect 27454 36814 27506 36866
rect 27506 36814 27508 36866
rect 27452 36812 27508 36814
rect 27612 36866 27668 36868
rect 27612 36814 27614 36866
rect 27614 36814 27666 36866
rect 27666 36814 27668 36866
rect 27612 36812 27668 36814
rect 27772 36866 27828 36868
rect 27772 36814 27774 36866
rect 27774 36814 27826 36866
rect 27826 36814 27828 36866
rect 27772 36812 27828 36814
rect 27932 36866 27988 36868
rect 27932 36814 27934 36866
rect 27934 36814 27986 36866
rect 27986 36814 27988 36866
rect 27932 36812 27988 36814
rect 28092 36866 28148 36868
rect 28092 36814 28094 36866
rect 28094 36814 28146 36866
rect 28146 36814 28148 36866
rect 28092 36812 28148 36814
rect 28252 36866 28308 36868
rect 28252 36814 28254 36866
rect 28254 36814 28306 36866
rect 28306 36814 28308 36866
rect 28252 36812 28308 36814
rect 28412 36866 28468 36868
rect 28412 36814 28414 36866
rect 28414 36814 28466 36866
rect 28466 36814 28468 36866
rect 28412 36812 28468 36814
rect 28572 36866 28628 36868
rect 28572 36814 28574 36866
rect 28574 36814 28626 36866
rect 28626 36814 28628 36866
rect 28572 36812 28628 36814
rect 28732 36866 28788 36868
rect 28732 36814 28734 36866
rect 28734 36814 28786 36866
rect 28786 36814 28788 36866
rect 28732 36812 28788 36814
rect 28892 36866 28948 36868
rect 28892 36814 28894 36866
rect 28894 36814 28946 36866
rect 28946 36814 28948 36866
rect 28892 36812 28948 36814
rect 29052 36866 29108 36868
rect 29052 36814 29054 36866
rect 29054 36814 29106 36866
rect 29106 36814 29108 36866
rect 29052 36812 29108 36814
rect 29212 36866 29268 36868
rect 29212 36814 29214 36866
rect 29214 36814 29266 36866
rect 29266 36814 29268 36866
rect 29212 36812 29268 36814
rect 29372 36866 29428 36868
rect 29372 36814 29374 36866
rect 29374 36814 29426 36866
rect 29426 36814 29428 36866
rect 29372 36812 29428 36814
rect 32572 36812 32628 36868
rect 32892 36812 32948 36868
rect 33532 36866 33588 36868
rect 33532 36814 33534 36866
rect 33534 36814 33586 36866
rect 33586 36814 33588 36866
rect 33532 36812 33588 36814
rect 33692 36866 33748 36868
rect 33692 36814 33694 36866
rect 33694 36814 33746 36866
rect 33746 36814 33748 36866
rect 33692 36812 33748 36814
rect 33852 36866 33908 36868
rect 33852 36814 33854 36866
rect 33854 36814 33906 36866
rect 33906 36814 33908 36866
rect 33852 36812 33908 36814
rect 34012 36866 34068 36868
rect 34012 36814 34014 36866
rect 34014 36814 34066 36866
rect 34066 36814 34068 36866
rect 34012 36812 34068 36814
rect 34172 36866 34228 36868
rect 34172 36814 34174 36866
rect 34174 36814 34226 36866
rect 34226 36814 34228 36866
rect 34172 36812 34228 36814
rect 34332 36866 34388 36868
rect 34332 36814 34334 36866
rect 34334 36814 34386 36866
rect 34386 36814 34388 36866
rect 34332 36812 34388 36814
rect 34492 36866 34548 36868
rect 34492 36814 34494 36866
rect 34494 36814 34546 36866
rect 34546 36814 34548 36866
rect 34492 36812 34548 36814
rect 34652 36866 34708 36868
rect 34652 36814 34654 36866
rect 34654 36814 34706 36866
rect 34706 36814 34708 36866
rect 34652 36812 34708 36814
rect 34812 36866 34868 36868
rect 34812 36814 34814 36866
rect 34814 36814 34866 36866
rect 34866 36814 34868 36866
rect 34812 36812 34868 36814
rect 34972 36866 35028 36868
rect 34972 36814 34974 36866
rect 34974 36814 35026 36866
rect 35026 36814 35028 36866
rect 34972 36812 35028 36814
rect 35132 36866 35188 36868
rect 35132 36814 35134 36866
rect 35134 36814 35186 36866
rect 35186 36814 35188 36866
rect 35132 36812 35188 36814
rect 35292 36866 35348 36868
rect 35292 36814 35294 36866
rect 35294 36814 35346 36866
rect 35346 36814 35348 36866
rect 35292 36812 35348 36814
rect 35452 36866 35508 36868
rect 35452 36814 35454 36866
rect 35454 36814 35506 36866
rect 35506 36814 35508 36866
rect 35452 36812 35508 36814
rect 35612 36866 35668 36868
rect 35612 36814 35614 36866
rect 35614 36814 35666 36866
rect 35666 36814 35668 36866
rect 35612 36812 35668 36814
rect 35772 36866 35828 36868
rect 35772 36814 35774 36866
rect 35774 36814 35826 36866
rect 35826 36814 35828 36866
rect 35772 36812 35828 36814
rect 35932 36866 35988 36868
rect 35932 36814 35934 36866
rect 35934 36814 35986 36866
rect 35986 36814 35988 36866
rect 35932 36812 35988 36814
rect 36092 36866 36148 36868
rect 36092 36814 36094 36866
rect 36094 36814 36146 36866
rect 36146 36814 36148 36866
rect 36092 36812 36148 36814
rect 36252 36866 36308 36868
rect 36252 36814 36254 36866
rect 36254 36814 36306 36866
rect 36306 36814 36308 36866
rect 36252 36812 36308 36814
rect 36412 36866 36468 36868
rect 36412 36814 36414 36866
rect 36414 36814 36466 36866
rect 36466 36814 36468 36866
rect 36412 36812 36468 36814
rect 36572 36866 36628 36868
rect 36572 36814 36574 36866
rect 36574 36814 36626 36866
rect 36626 36814 36628 36866
rect 36572 36812 36628 36814
rect 36732 36866 36788 36868
rect 36732 36814 36734 36866
rect 36734 36814 36786 36866
rect 36786 36814 36788 36866
rect 36732 36812 36788 36814
rect 36892 36866 36948 36868
rect 36892 36814 36894 36866
rect 36894 36814 36946 36866
rect 36946 36814 36948 36866
rect 36892 36812 36948 36814
rect 37052 36866 37108 36868
rect 37052 36814 37054 36866
rect 37054 36814 37106 36866
rect 37106 36814 37108 36866
rect 37052 36812 37108 36814
rect 37212 36866 37268 36868
rect 37212 36814 37214 36866
rect 37214 36814 37266 36866
rect 37266 36814 37268 36866
rect 37212 36812 37268 36814
rect 37372 36866 37428 36868
rect 37372 36814 37374 36866
rect 37374 36814 37426 36866
rect 37426 36814 37428 36866
rect 37372 36812 37428 36814
rect 37532 36866 37588 36868
rect 37532 36814 37534 36866
rect 37534 36814 37586 36866
rect 37586 36814 37588 36866
rect 37532 36812 37588 36814
rect 37692 36866 37748 36868
rect 37692 36814 37694 36866
rect 37694 36814 37746 36866
rect 37746 36814 37748 36866
rect 37692 36812 37748 36814
rect 37852 36866 37908 36868
rect 37852 36814 37854 36866
rect 37854 36814 37906 36866
rect 37906 36814 37908 36866
rect 37852 36812 37908 36814
rect 38012 36866 38068 36868
rect 38012 36814 38014 36866
rect 38014 36814 38066 36866
rect 38066 36814 38068 36866
rect 38012 36812 38068 36814
rect 38172 36866 38228 36868
rect 38172 36814 38174 36866
rect 38174 36814 38226 36866
rect 38226 36814 38228 36866
rect 38172 36812 38228 36814
rect 38332 36866 38388 36868
rect 38332 36814 38334 36866
rect 38334 36814 38386 36866
rect 38386 36814 38388 36866
rect 38332 36812 38388 36814
rect 38492 36866 38548 36868
rect 38492 36814 38494 36866
rect 38494 36814 38546 36866
rect 38546 36814 38548 36866
rect 38492 36812 38548 36814
rect 38652 36866 38708 36868
rect 38652 36814 38654 36866
rect 38654 36814 38706 36866
rect 38706 36814 38708 36866
rect 38652 36812 38708 36814
rect 38812 36866 38868 36868
rect 38812 36814 38814 36866
rect 38814 36814 38866 36866
rect 38866 36814 38868 36866
rect 38812 36812 38868 36814
rect 38972 36866 39028 36868
rect 38972 36814 38974 36866
rect 38974 36814 39026 36866
rect 39026 36814 39028 36866
rect 38972 36812 39028 36814
rect 39132 36866 39188 36868
rect 39132 36814 39134 36866
rect 39134 36814 39186 36866
rect 39186 36814 39188 36866
rect 39132 36812 39188 36814
rect 39292 36866 39348 36868
rect 39292 36814 39294 36866
rect 39294 36814 39346 36866
rect 39346 36814 39348 36866
rect 39292 36812 39348 36814
rect 39452 36866 39508 36868
rect 39452 36814 39454 36866
rect 39454 36814 39506 36866
rect 39506 36814 39508 36866
rect 39452 36812 39508 36814
rect 39612 36866 39668 36868
rect 39612 36814 39614 36866
rect 39614 36814 39666 36866
rect 39666 36814 39668 36866
rect 39612 36812 39668 36814
rect 39772 36866 39828 36868
rect 39772 36814 39774 36866
rect 39774 36814 39826 36866
rect 39826 36814 39828 36866
rect 39772 36812 39828 36814
rect 39932 36866 39988 36868
rect 39932 36814 39934 36866
rect 39934 36814 39986 36866
rect 39986 36814 39988 36866
rect 39932 36812 39988 36814
rect 40092 36866 40148 36868
rect 40092 36814 40094 36866
rect 40094 36814 40146 36866
rect 40146 36814 40148 36866
rect 40092 36812 40148 36814
rect 40252 36866 40308 36868
rect 40252 36814 40254 36866
rect 40254 36814 40306 36866
rect 40306 36814 40308 36866
rect 40252 36812 40308 36814
rect 40412 36866 40468 36868
rect 40412 36814 40414 36866
rect 40414 36814 40466 36866
rect 40466 36814 40468 36866
rect 40412 36812 40468 36814
rect 40572 36866 40628 36868
rect 40572 36814 40574 36866
rect 40574 36814 40626 36866
rect 40626 36814 40628 36866
rect 40572 36812 40628 36814
rect 40732 36866 40788 36868
rect 40732 36814 40734 36866
rect 40734 36814 40786 36866
rect 40786 36814 40788 36866
rect 40732 36812 40788 36814
rect 40892 36866 40948 36868
rect 40892 36814 40894 36866
rect 40894 36814 40946 36866
rect 40946 36814 40948 36866
rect 40892 36812 40948 36814
rect 41052 36866 41108 36868
rect 41052 36814 41054 36866
rect 41054 36814 41106 36866
rect 41106 36814 41108 36866
rect 41052 36812 41108 36814
rect 41212 36866 41268 36868
rect 41212 36814 41214 36866
rect 41214 36814 41266 36866
rect 41266 36814 41268 36866
rect 41212 36812 41268 36814
rect 41372 36866 41428 36868
rect 41372 36814 41374 36866
rect 41374 36814 41426 36866
rect 41426 36814 41428 36866
rect 41372 36812 41428 36814
rect 41532 36866 41588 36868
rect 41532 36814 41534 36866
rect 41534 36814 41586 36866
rect 41586 36814 41588 36866
rect 41532 36812 41588 36814
rect 41692 36866 41748 36868
rect 41692 36814 41694 36866
rect 41694 36814 41746 36866
rect 41746 36814 41748 36866
rect 41692 36812 41748 36814
rect 41852 36866 41908 36868
rect 41852 36814 41854 36866
rect 41854 36814 41906 36866
rect 41906 36814 41908 36866
rect 41852 36812 41908 36814
rect 9132 36652 9188 36708
rect 22252 36652 22308 36708
rect 32732 36652 32788 36708
rect 12 36546 68 36548
rect 12 36494 14 36546
rect 14 36494 66 36546
rect 66 36494 68 36546
rect 12 36492 68 36494
rect 172 36546 228 36548
rect 172 36494 174 36546
rect 174 36494 226 36546
rect 226 36494 228 36546
rect 172 36492 228 36494
rect 332 36546 388 36548
rect 332 36494 334 36546
rect 334 36494 386 36546
rect 386 36494 388 36546
rect 332 36492 388 36494
rect 492 36546 548 36548
rect 492 36494 494 36546
rect 494 36494 546 36546
rect 546 36494 548 36546
rect 492 36492 548 36494
rect 652 36546 708 36548
rect 652 36494 654 36546
rect 654 36494 706 36546
rect 706 36494 708 36546
rect 652 36492 708 36494
rect 812 36546 868 36548
rect 812 36494 814 36546
rect 814 36494 866 36546
rect 866 36494 868 36546
rect 812 36492 868 36494
rect 972 36546 1028 36548
rect 972 36494 974 36546
rect 974 36494 1026 36546
rect 1026 36494 1028 36546
rect 972 36492 1028 36494
rect 1132 36546 1188 36548
rect 1132 36494 1134 36546
rect 1134 36494 1186 36546
rect 1186 36494 1188 36546
rect 1132 36492 1188 36494
rect 1292 36546 1348 36548
rect 1292 36494 1294 36546
rect 1294 36494 1346 36546
rect 1346 36494 1348 36546
rect 1292 36492 1348 36494
rect 1452 36546 1508 36548
rect 1452 36494 1454 36546
rect 1454 36494 1506 36546
rect 1506 36494 1508 36546
rect 1452 36492 1508 36494
rect 1612 36546 1668 36548
rect 1612 36494 1614 36546
rect 1614 36494 1666 36546
rect 1666 36494 1668 36546
rect 1612 36492 1668 36494
rect 1772 36546 1828 36548
rect 1772 36494 1774 36546
rect 1774 36494 1826 36546
rect 1826 36494 1828 36546
rect 1772 36492 1828 36494
rect 1932 36546 1988 36548
rect 1932 36494 1934 36546
rect 1934 36494 1986 36546
rect 1986 36494 1988 36546
rect 1932 36492 1988 36494
rect 2092 36546 2148 36548
rect 2092 36494 2094 36546
rect 2094 36494 2146 36546
rect 2146 36494 2148 36546
rect 2092 36492 2148 36494
rect 2252 36546 2308 36548
rect 2252 36494 2254 36546
rect 2254 36494 2306 36546
rect 2306 36494 2308 36546
rect 2252 36492 2308 36494
rect 2412 36546 2468 36548
rect 2412 36494 2414 36546
rect 2414 36494 2466 36546
rect 2466 36494 2468 36546
rect 2412 36492 2468 36494
rect 2572 36546 2628 36548
rect 2572 36494 2574 36546
rect 2574 36494 2626 36546
rect 2626 36494 2628 36546
rect 2572 36492 2628 36494
rect 2732 36546 2788 36548
rect 2732 36494 2734 36546
rect 2734 36494 2786 36546
rect 2786 36494 2788 36546
rect 2732 36492 2788 36494
rect 2892 36546 2948 36548
rect 2892 36494 2894 36546
rect 2894 36494 2946 36546
rect 2946 36494 2948 36546
rect 2892 36492 2948 36494
rect 3052 36546 3108 36548
rect 3052 36494 3054 36546
rect 3054 36494 3106 36546
rect 3106 36494 3108 36546
rect 3052 36492 3108 36494
rect 3212 36546 3268 36548
rect 3212 36494 3214 36546
rect 3214 36494 3266 36546
rect 3266 36494 3268 36546
rect 3212 36492 3268 36494
rect 3372 36546 3428 36548
rect 3372 36494 3374 36546
rect 3374 36494 3426 36546
rect 3426 36494 3428 36546
rect 3372 36492 3428 36494
rect 3532 36546 3588 36548
rect 3532 36494 3534 36546
rect 3534 36494 3586 36546
rect 3586 36494 3588 36546
rect 3532 36492 3588 36494
rect 3692 36546 3748 36548
rect 3692 36494 3694 36546
rect 3694 36494 3746 36546
rect 3746 36494 3748 36546
rect 3692 36492 3748 36494
rect 3852 36546 3908 36548
rect 3852 36494 3854 36546
rect 3854 36494 3906 36546
rect 3906 36494 3908 36546
rect 3852 36492 3908 36494
rect 4012 36546 4068 36548
rect 4012 36494 4014 36546
rect 4014 36494 4066 36546
rect 4066 36494 4068 36546
rect 4012 36492 4068 36494
rect 4172 36546 4228 36548
rect 4172 36494 4174 36546
rect 4174 36494 4226 36546
rect 4226 36494 4228 36546
rect 4172 36492 4228 36494
rect 4332 36546 4388 36548
rect 4332 36494 4334 36546
rect 4334 36494 4386 36546
rect 4386 36494 4388 36546
rect 4332 36492 4388 36494
rect 4492 36546 4548 36548
rect 4492 36494 4494 36546
rect 4494 36494 4546 36546
rect 4546 36494 4548 36546
rect 4492 36492 4548 36494
rect 4652 36546 4708 36548
rect 4652 36494 4654 36546
rect 4654 36494 4706 36546
rect 4706 36494 4708 36546
rect 4652 36492 4708 36494
rect 4812 36546 4868 36548
rect 4812 36494 4814 36546
rect 4814 36494 4866 36546
rect 4866 36494 4868 36546
rect 4812 36492 4868 36494
rect 4972 36546 5028 36548
rect 4972 36494 4974 36546
rect 4974 36494 5026 36546
rect 5026 36494 5028 36546
rect 4972 36492 5028 36494
rect 5132 36546 5188 36548
rect 5132 36494 5134 36546
rect 5134 36494 5186 36546
rect 5186 36494 5188 36546
rect 5132 36492 5188 36494
rect 5292 36546 5348 36548
rect 5292 36494 5294 36546
rect 5294 36494 5346 36546
rect 5346 36494 5348 36546
rect 5292 36492 5348 36494
rect 5452 36546 5508 36548
rect 5452 36494 5454 36546
rect 5454 36494 5506 36546
rect 5506 36494 5508 36546
rect 5452 36492 5508 36494
rect 5612 36546 5668 36548
rect 5612 36494 5614 36546
rect 5614 36494 5666 36546
rect 5666 36494 5668 36546
rect 5612 36492 5668 36494
rect 5772 36546 5828 36548
rect 5772 36494 5774 36546
rect 5774 36494 5826 36546
rect 5826 36494 5828 36546
rect 5772 36492 5828 36494
rect 5932 36546 5988 36548
rect 5932 36494 5934 36546
rect 5934 36494 5986 36546
rect 5986 36494 5988 36546
rect 5932 36492 5988 36494
rect 6092 36546 6148 36548
rect 6092 36494 6094 36546
rect 6094 36494 6146 36546
rect 6146 36494 6148 36546
rect 6092 36492 6148 36494
rect 6252 36546 6308 36548
rect 6252 36494 6254 36546
rect 6254 36494 6306 36546
rect 6306 36494 6308 36546
rect 6252 36492 6308 36494
rect 6412 36546 6468 36548
rect 6412 36494 6414 36546
rect 6414 36494 6466 36546
rect 6466 36494 6468 36546
rect 6412 36492 6468 36494
rect 6572 36546 6628 36548
rect 6572 36494 6574 36546
rect 6574 36494 6626 36546
rect 6626 36494 6628 36546
rect 6572 36492 6628 36494
rect 6732 36546 6788 36548
rect 6732 36494 6734 36546
rect 6734 36494 6786 36546
rect 6786 36494 6788 36546
rect 6732 36492 6788 36494
rect 6892 36546 6948 36548
rect 6892 36494 6894 36546
rect 6894 36494 6946 36546
rect 6946 36494 6948 36546
rect 6892 36492 6948 36494
rect 7052 36546 7108 36548
rect 7052 36494 7054 36546
rect 7054 36494 7106 36546
rect 7106 36494 7108 36546
rect 7052 36492 7108 36494
rect 7212 36546 7268 36548
rect 7212 36494 7214 36546
rect 7214 36494 7266 36546
rect 7266 36494 7268 36546
rect 7212 36492 7268 36494
rect 7372 36546 7428 36548
rect 7372 36494 7374 36546
rect 7374 36494 7426 36546
rect 7426 36494 7428 36546
rect 7372 36492 7428 36494
rect 7532 36546 7588 36548
rect 7532 36494 7534 36546
rect 7534 36494 7586 36546
rect 7586 36494 7588 36546
rect 7532 36492 7588 36494
rect 7692 36546 7748 36548
rect 7692 36494 7694 36546
rect 7694 36494 7746 36546
rect 7746 36494 7748 36546
rect 7692 36492 7748 36494
rect 7852 36546 7908 36548
rect 7852 36494 7854 36546
rect 7854 36494 7906 36546
rect 7906 36494 7908 36546
rect 7852 36492 7908 36494
rect 8012 36546 8068 36548
rect 8012 36494 8014 36546
rect 8014 36494 8066 36546
rect 8066 36494 8068 36546
rect 8012 36492 8068 36494
rect 8172 36546 8228 36548
rect 8172 36494 8174 36546
rect 8174 36494 8226 36546
rect 8226 36494 8228 36546
rect 8172 36492 8228 36494
rect 8332 36546 8388 36548
rect 8332 36494 8334 36546
rect 8334 36494 8386 36546
rect 8386 36494 8388 36546
rect 8332 36492 8388 36494
rect 8972 36492 9028 36548
rect 9292 36492 9348 36548
rect 12492 36546 12548 36548
rect 12492 36494 12494 36546
rect 12494 36494 12546 36546
rect 12546 36494 12548 36546
rect 12492 36492 12548 36494
rect 12652 36546 12708 36548
rect 12652 36494 12654 36546
rect 12654 36494 12706 36546
rect 12706 36494 12708 36546
rect 12652 36492 12708 36494
rect 12812 36546 12868 36548
rect 12812 36494 12814 36546
rect 12814 36494 12866 36546
rect 12866 36494 12868 36546
rect 12812 36492 12868 36494
rect 12972 36546 13028 36548
rect 12972 36494 12974 36546
rect 12974 36494 13026 36546
rect 13026 36494 13028 36546
rect 12972 36492 13028 36494
rect 13132 36546 13188 36548
rect 13132 36494 13134 36546
rect 13134 36494 13186 36546
rect 13186 36494 13188 36546
rect 13132 36492 13188 36494
rect 13292 36546 13348 36548
rect 13292 36494 13294 36546
rect 13294 36494 13346 36546
rect 13346 36494 13348 36546
rect 13292 36492 13348 36494
rect 13452 36546 13508 36548
rect 13452 36494 13454 36546
rect 13454 36494 13506 36546
rect 13506 36494 13508 36546
rect 13452 36492 13508 36494
rect 13612 36546 13668 36548
rect 13612 36494 13614 36546
rect 13614 36494 13666 36546
rect 13666 36494 13668 36546
rect 13612 36492 13668 36494
rect 13772 36546 13828 36548
rect 13772 36494 13774 36546
rect 13774 36494 13826 36546
rect 13826 36494 13828 36546
rect 13772 36492 13828 36494
rect 13932 36546 13988 36548
rect 13932 36494 13934 36546
rect 13934 36494 13986 36546
rect 13986 36494 13988 36546
rect 13932 36492 13988 36494
rect 14092 36546 14148 36548
rect 14092 36494 14094 36546
rect 14094 36494 14146 36546
rect 14146 36494 14148 36546
rect 14092 36492 14148 36494
rect 14252 36546 14308 36548
rect 14252 36494 14254 36546
rect 14254 36494 14306 36546
rect 14306 36494 14308 36546
rect 14252 36492 14308 36494
rect 14412 36546 14468 36548
rect 14412 36494 14414 36546
rect 14414 36494 14466 36546
rect 14466 36494 14468 36546
rect 14412 36492 14468 36494
rect 14572 36546 14628 36548
rect 14572 36494 14574 36546
rect 14574 36494 14626 36546
rect 14626 36494 14628 36546
rect 14572 36492 14628 36494
rect 14732 36546 14788 36548
rect 14732 36494 14734 36546
rect 14734 36494 14786 36546
rect 14786 36494 14788 36546
rect 14732 36492 14788 36494
rect 14892 36546 14948 36548
rect 14892 36494 14894 36546
rect 14894 36494 14946 36546
rect 14946 36494 14948 36546
rect 14892 36492 14948 36494
rect 15052 36546 15108 36548
rect 15052 36494 15054 36546
rect 15054 36494 15106 36546
rect 15106 36494 15108 36546
rect 15052 36492 15108 36494
rect 15212 36546 15268 36548
rect 15212 36494 15214 36546
rect 15214 36494 15266 36546
rect 15266 36494 15268 36546
rect 15212 36492 15268 36494
rect 15372 36546 15428 36548
rect 15372 36494 15374 36546
rect 15374 36494 15426 36546
rect 15426 36494 15428 36546
rect 15372 36492 15428 36494
rect 15532 36546 15588 36548
rect 15532 36494 15534 36546
rect 15534 36494 15586 36546
rect 15586 36494 15588 36546
rect 15532 36492 15588 36494
rect 15692 36546 15748 36548
rect 15692 36494 15694 36546
rect 15694 36494 15746 36546
rect 15746 36494 15748 36546
rect 15692 36492 15748 36494
rect 15852 36546 15908 36548
rect 15852 36494 15854 36546
rect 15854 36494 15906 36546
rect 15906 36494 15908 36546
rect 15852 36492 15908 36494
rect 16012 36546 16068 36548
rect 16012 36494 16014 36546
rect 16014 36494 16066 36546
rect 16066 36494 16068 36546
rect 16012 36492 16068 36494
rect 16172 36546 16228 36548
rect 16172 36494 16174 36546
rect 16174 36494 16226 36546
rect 16226 36494 16228 36546
rect 16172 36492 16228 36494
rect 16332 36546 16388 36548
rect 16332 36494 16334 36546
rect 16334 36494 16386 36546
rect 16386 36494 16388 36546
rect 16332 36492 16388 36494
rect 16492 36546 16548 36548
rect 16492 36494 16494 36546
rect 16494 36494 16546 36546
rect 16546 36494 16548 36546
rect 16492 36492 16548 36494
rect 16652 36546 16708 36548
rect 16652 36494 16654 36546
rect 16654 36494 16706 36546
rect 16706 36494 16708 36546
rect 16652 36492 16708 36494
rect 16812 36546 16868 36548
rect 16812 36494 16814 36546
rect 16814 36494 16866 36546
rect 16866 36494 16868 36546
rect 16812 36492 16868 36494
rect 16972 36546 17028 36548
rect 16972 36494 16974 36546
rect 16974 36494 17026 36546
rect 17026 36494 17028 36546
rect 16972 36492 17028 36494
rect 17132 36546 17188 36548
rect 17132 36494 17134 36546
rect 17134 36494 17186 36546
rect 17186 36494 17188 36546
rect 17132 36492 17188 36494
rect 17292 36546 17348 36548
rect 17292 36494 17294 36546
rect 17294 36494 17346 36546
rect 17346 36494 17348 36546
rect 17292 36492 17348 36494
rect 17452 36546 17508 36548
rect 17452 36494 17454 36546
rect 17454 36494 17506 36546
rect 17506 36494 17508 36546
rect 17452 36492 17508 36494
rect 17612 36546 17668 36548
rect 17612 36494 17614 36546
rect 17614 36494 17666 36546
rect 17666 36494 17668 36546
rect 17612 36492 17668 36494
rect 17772 36546 17828 36548
rect 17772 36494 17774 36546
rect 17774 36494 17826 36546
rect 17826 36494 17828 36546
rect 17772 36492 17828 36494
rect 17932 36546 17988 36548
rect 17932 36494 17934 36546
rect 17934 36494 17986 36546
rect 17986 36494 17988 36546
rect 17932 36492 17988 36494
rect 18092 36546 18148 36548
rect 18092 36494 18094 36546
rect 18094 36494 18146 36546
rect 18146 36494 18148 36546
rect 18092 36492 18148 36494
rect 18252 36546 18308 36548
rect 18252 36494 18254 36546
rect 18254 36494 18306 36546
rect 18306 36494 18308 36546
rect 18252 36492 18308 36494
rect 18412 36546 18468 36548
rect 18412 36494 18414 36546
rect 18414 36494 18466 36546
rect 18466 36494 18468 36546
rect 18412 36492 18468 36494
rect 18572 36546 18628 36548
rect 18572 36494 18574 36546
rect 18574 36494 18626 36546
rect 18626 36494 18628 36546
rect 18572 36492 18628 36494
rect 18732 36546 18788 36548
rect 18732 36494 18734 36546
rect 18734 36494 18786 36546
rect 18786 36494 18788 36546
rect 18732 36492 18788 36494
rect 18892 36546 18948 36548
rect 18892 36494 18894 36546
rect 18894 36494 18946 36546
rect 18946 36494 18948 36546
rect 18892 36492 18948 36494
rect 22092 36492 22148 36548
rect 22412 36492 22468 36548
rect 23132 36546 23188 36548
rect 23132 36494 23134 36546
rect 23134 36494 23186 36546
rect 23186 36494 23188 36546
rect 23132 36492 23188 36494
rect 23292 36546 23348 36548
rect 23292 36494 23294 36546
rect 23294 36494 23346 36546
rect 23346 36494 23348 36546
rect 23292 36492 23348 36494
rect 23452 36546 23508 36548
rect 23452 36494 23454 36546
rect 23454 36494 23506 36546
rect 23506 36494 23508 36546
rect 23452 36492 23508 36494
rect 23612 36546 23668 36548
rect 23612 36494 23614 36546
rect 23614 36494 23666 36546
rect 23666 36494 23668 36546
rect 23612 36492 23668 36494
rect 23772 36546 23828 36548
rect 23772 36494 23774 36546
rect 23774 36494 23826 36546
rect 23826 36494 23828 36546
rect 23772 36492 23828 36494
rect 23932 36546 23988 36548
rect 23932 36494 23934 36546
rect 23934 36494 23986 36546
rect 23986 36494 23988 36546
rect 23932 36492 23988 36494
rect 24092 36546 24148 36548
rect 24092 36494 24094 36546
rect 24094 36494 24146 36546
rect 24146 36494 24148 36546
rect 24092 36492 24148 36494
rect 24252 36546 24308 36548
rect 24252 36494 24254 36546
rect 24254 36494 24306 36546
rect 24306 36494 24308 36546
rect 24252 36492 24308 36494
rect 24412 36546 24468 36548
rect 24412 36494 24414 36546
rect 24414 36494 24466 36546
rect 24466 36494 24468 36546
rect 24412 36492 24468 36494
rect 24572 36546 24628 36548
rect 24572 36494 24574 36546
rect 24574 36494 24626 36546
rect 24626 36494 24628 36546
rect 24572 36492 24628 36494
rect 24732 36546 24788 36548
rect 24732 36494 24734 36546
rect 24734 36494 24786 36546
rect 24786 36494 24788 36546
rect 24732 36492 24788 36494
rect 24892 36546 24948 36548
rect 24892 36494 24894 36546
rect 24894 36494 24946 36546
rect 24946 36494 24948 36546
rect 24892 36492 24948 36494
rect 25052 36546 25108 36548
rect 25052 36494 25054 36546
rect 25054 36494 25106 36546
rect 25106 36494 25108 36546
rect 25052 36492 25108 36494
rect 25212 36546 25268 36548
rect 25212 36494 25214 36546
rect 25214 36494 25266 36546
rect 25266 36494 25268 36546
rect 25212 36492 25268 36494
rect 25372 36546 25428 36548
rect 25372 36494 25374 36546
rect 25374 36494 25426 36546
rect 25426 36494 25428 36546
rect 25372 36492 25428 36494
rect 25532 36546 25588 36548
rect 25532 36494 25534 36546
rect 25534 36494 25586 36546
rect 25586 36494 25588 36546
rect 25532 36492 25588 36494
rect 25692 36546 25748 36548
rect 25692 36494 25694 36546
rect 25694 36494 25746 36546
rect 25746 36494 25748 36546
rect 25692 36492 25748 36494
rect 25852 36546 25908 36548
rect 25852 36494 25854 36546
rect 25854 36494 25906 36546
rect 25906 36494 25908 36546
rect 25852 36492 25908 36494
rect 26012 36546 26068 36548
rect 26012 36494 26014 36546
rect 26014 36494 26066 36546
rect 26066 36494 26068 36546
rect 26012 36492 26068 36494
rect 26172 36546 26228 36548
rect 26172 36494 26174 36546
rect 26174 36494 26226 36546
rect 26226 36494 26228 36546
rect 26172 36492 26228 36494
rect 26332 36546 26388 36548
rect 26332 36494 26334 36546
rect 26334 36494 26386 36546
rect 26386 36494 26388 36546
rect 26332 36492 26388 36494
rect 26492 36546 26548 36548
rect 26492 36494 26494 36546
rect 26494 36494 26546 36546
rect 26546 36494 26548 36546
rect 26492 36492 26548 36494
rect 26652 36546 26708 36548
rect 26652 36494 26654 36546
rect 26654 36494 26706 36546
rect 26706 36494 26708 36546
rect 26652 36492 26708 36494
rect 26812 36546 26868 36548
rect 26812 36494 26814 36546
rect 26814 36494 26866 36546
rect 26866 36494 26868 36546
rect 26812 36492 26868 36494
rect 26972 36546 27028 36548
rect 26972 36494 26974 36546
rect 26974 36494 27026 36546
rect 27026 36494 27028 36546
rect 26972 36492 27028 36494
rect 27132 36546 27188 36548
rect 27132 36494 27134 36546
rect 27134 36494 27186 36546
rect 27186 36494 27188 36546
rect 27132 36492 27188 36494
rect 27292 36546 27348 36548
rect 27292 36494 27294 36546
rect 27294 36494 27346 36546
rect 27346 36494 27348 36546
rect 27292 36492 27348 36494
rect 27452 36546 27508 36548
rect 27452 36494 27454 36546
rect 27454 36494 27506 36546
rect 27506 36494 27508 36546
rect 27452 36492 27508 36494
rect 27612 36546 27668 36548
rect 27612 36494 27614 36546
rect 27614 36494 27666 36546
rect 27666 36494 27668 36546
rect 27612 36492 27668 36494
rect 27772 36546 27828 36548
rect 27772 36494 27774 36546
rect 27774 36494 27826 36546
rect 27826 36494 27828 36546
rect 27772 36492 27828 36494
rect 27932 36546 27988 36548
rect 27932 36494 27934 36546
rect 27934 36494 27986 36546
rect 27986 36494 27988 36546
rect 27932 36492 27988 36494
rect 28092 36546 28148 36548
rect 28092 36494 28094 36546
rect 28094 36494 28146 36546
rect 28146 36494 28148 36546
rect 28092 36492 28148 36494
rect 28252 36546 28308 36548
rect 28252 36494 28254 36546
rect 28254 36494 28306 36546
rect 28306 36494 28308 36546
rect 28252 36492 28308 36494
rect 28412 36546 28468 36548
rect 28412 36494 28414 36546
rect 28414 36494 28466 36546
rect 28466 36494 28468 36546
rect 28412 36492 28468 36494
rect 28572 36546 28628 36548
rect 28572 36494 28574 36546
rect 28574 36494 28626 36546
rect 28626 36494 28628 36546
rect 28572 36492 28628 36494
rect 28732 36546 28788 36548
rect 28732 36494 28734 36546
rect 28734 36494 28786 36546
rect 28786 36494 28788 36546
rect 28732 36492 28788 36494
rect 28892 36546 28948 36548
rect 28892 36494 28894 36546
rect 28894 36494 28946 36546
rect 28946 36494 28948 36546
rect 28892 36492 28948 36494
rect 29052 36546 29108 36548
rect 29052 36494 29054 36546
rect 29054 36494 29106 36546
rect 29106 36494 29108 36546
rect 29052 36492 29108 36494
rect 29212 36546 29268 36548
rect 29212 36494 29214 36546
rect 29214 36494 29266 36546
rect 29266 36494 29268 36546
rect 29212 36492 29268 36494
rect 29372 36546 29428 36548
rect 29372 36494 29374 36546
rect 29374 36494 29426 36546
rect 29426 36494 29428 36546
rect 29372 36492 29428 36494
rect 32572 36492 32628 36548
rect 32892 36492 32948 36548
rect 33532 36546 33588 36548
rect 33532 36494 33534 36546
rect 33534 36494 33586 36546
rect 33586 36494 33588 36546
rect 33532 36492 33588 36494
rect 33692 36546 33748 36548
rect 33692 36494 33694 36546
rect 33694 36494 33746 36546
rect 33746 36494 33748 36546
rect 33692 36492 33748 36494
rect 33852 36546 33908 36548
rect 33852 36494 33854 36546
rect 33854 36494 33906 36546
rect 33906 36494 33908 36546
rect 33852 36492 33908 36494
rect 34012 36546 34068 36548
rect 34012 36494 34014 36546
rect 34014 36494 34066 36546
rect 34066 36494 34068 36546
rect 34012 36492 34068 36494
rect 34172 36546 34228 36548
rect 34172 36494 34174 36546
rect 34174 36494 34226 36546
rect 34226 36494 34228 36546
rect 34172 36492 34228 36494
rect 34332 36546 34388 36548
rect 34332 36494 34334 36546
rect 34334 36494 34386 36546
rect 34386 36494 34388 36546
rect 34332 36492 34388 36494
rect 34492 36546 34548 36548
rect 34492 36494 34494 36546
rect 34494 36494 34546 36546
rect 34546 36494 34548 36546
rect 34492 36492 34548 36494
rect 34652 36546 34708 36548
rect 34652 36494 34654 36546
rect 34654 36494 34706 36546
rect 34706 36494 34708 36546
rect 34652 36492 34708 36494
rect 34812 36546 34868 36548
rect 34812 36494 34814 36546
rect 34814 36494 34866 36546
rect 34866 36494 34868 36546
rect 34812 36492 34868 36494
rect 34972 36546 35028 36548
rect 34972 36494 34974 36546
rect 34974 36494 35026 36546
rect 35026 36494 35028 36546
rect 34972 36492 35028 36494
rect 35132 36546 35188 36548
rect 35132 36494 35134 36546
rect 35134 36494 35186 36546
rect 35186 36494 35188 36546
rect 35132 36492 35188 36494
rect 35292 36546 35348 36548
rect 35292 36494 35294 36546
rect 35294 36494 35346 36546
rect 35346 36494 35348 36546
rect 35292 36492 35348 36494
rect 35452 36546 35508 36548
rect 35452 36494 35454 36546
rect 35454 36494 35506 36546
rect 35506 36494 35508 36546
rect 35452 36492 35508 36494
rect 35612 36546 35668 36548
rect 35612 36494 35614 36546
rect 35614 36494 35666 36546
rect 35666 36494 35668 36546
rect 35612 36492 35668 36494
rect 35772 36546 35828 36548
rect 35772 36494 35774 36546
rect 35774 36494 35826 36546
rect 35826 36494 35828 36546
rect 35772 36492 35828 36494
rect 35932 36546 35988 36548
rect 35932 36494 35934 36546
rect 35934 36494 35986 36546
rect 35986 36494 35988 36546
rect 35932 36492 35988 36494
rect 36092 36546 36148 36548
rect 36092 36494 36094 36546
rect 36094 36494 36146 36546
rect 36146 36494 36148 36546
rect 36092 36492 36148 36494
rect 36252 36546 36308 36548
rect 36252 36494 36254 36546
rect 36254 36494 36306 36546
rect 36306 36494 36308 36546
rect 36252 36492 36308 36494
rect 36412 36546 36468 36548
rect 36412 36494 36414 36546
rect 36414 36494 36466 36546
rect 36466 36494 36468 36546
rect 36412 36492 36468 36494
rect 36572 36546 36628 36548
rect 36572 36494 36574 36546
rect 36574 36494 36626 36546
rect 36626 36494 36628 36546
rect 36572 36492 36628 36494
rect 36732 36546 36788 36548
rect 36732 36494 36734 36546
rect 36734 36494 36786 36546
rect 36786 36494 36788 36546
rect 36732 36492 36788 36494
rect 36892 36546 36948 36548
rect 36892 36494 36894 36546
rect 36894 36494 36946 36546
rect 36946 36494 36948 36546
rect 36892 36492 36948 36494
rect 37052 36546 37108 36548
rect 37052 36494 37054 36546
rect 37054 36494 37106 36546
rect 37106 36494 37108 36546
rect 37052 36492 37108 36494
rect 37212 36546 37268 36548
rect 37212 36494 37214 36546
rect 37214 36494 37266 36546
rect 37266 36494 37268 36546
rect 37212 36492 37268 36494
rect 37372 36546 37428 36548
rect 37372 36494 37374 36546
rect 37374 36494 37426 36546
rect 37426 36494 37428 36546
rect 37372 36492 37428 36494
rect 37532 36546 37588 36548
rect 37532 36494 37534 36546
rect 37534 36494 37586 36546
rect 37586 36494 37588 36546
rect 37532 36492 37588 36494
rect 37692 36546 37748 36548
rect 37692 36494 37694 36546
rect 37694 36494 37746 36546
rect 37746 36494 37748 36546
rect 37692 36492 37748 36494
rect 37852 36546 37908 36548
rect 37852 36494 37854 36546
rect 37854 36494 37906 36546
rect 37906 36494 37908 36546
rect 37852 36492 37908 36494
rect 38012 36546 38068 36548
rect 38012 36494 38014 36546
rect 38014 36494 38066 36546
rect 38066 36494 38068 36546
rect 38012 36492 38068 36494
rect 38172 36546 38228 36548
rect 38172 36494 38174 36546
rect 38174 36494 38226 36546
rect 38226 36494 38228 36546
rect 38172 36492 38228 36494
rect 38332 36546 38388 36548
rect 38332 36494 38334 36546
rect 38334 36494 38386 36546
rect 38386 36494 38388 36546
rect 38332 36492 38388 36494
rect 38492 36546 38548 36548
rect 38492 36494 38494 36546
rect 38494 36494 38546 36546
rect 38546 36494 38548 36546
rect 38492 36492 38548 36494
rect 38652 36546 38708 36548
rect 38652 36494 38654 36546
rect 38654 36494 38706 36546
rect 38706 36494 38708 36546
rect 38652 36492 38708 36494
rect 38812 36546 38868 36548
rect 38812 36494 38814 36546
rect 38814 36494 38866 36546
rect 38866 36494 38868 36546
rect 38812 36492 38868 36494
rect 38972 36546 39028 36548
rect 38972 36494 38974 36546
rect 38974 36494 39026 36546
rect 39026 36494 39028 36546
rect 38972 36492 39028 36494
rect 39132 36546 39188 36548
rect 39132 36494 39134 36546
rect 39134 36494 39186 36546
rect 39186 36494 39188 36546
rect 39132 36492 39188 36494
rect 39292 36546 39348 36548
rect 39292 36494 39294 36546
rect 39294 36494 39346 36546
rect 39346 36494 39348 36546
rect 39292 36492 39348 36494
rect 39452 36546 39508 36548
rect 39452 36494 39454 36546
rect 39454 36494 39506 36546
rect 39506 36494 39508 36546
rect 39452 36492 39508 36494
rect 39612 36546 39668 36548
rect 39612 36494 39614 36546
rect 39614 36494 39666 36546
rect 39666 36494 39668 36546
rect 39612 36492 39668 36494
rect 39772 36546 39828 36548
rect 39772 36494 39774 36546
rect 39774 36494 39826 36546
rect 39826 36494 39828 36546
rect 39772 36492 39828 36494
rect 39932 36546 39988 36548
rect 39932 36494 39934 36546
rect 39934 36494 39986 36546
rect 39986 36494 39988 36546
rect 39932 36492 39988 36494
rect 40092 36546 40148 36548
rect 40092 36494 40094 36546
rect 40094 36494 40146 36546
rect 40146 36494 40148 36546
rect 40092 36492 40148 36494
rect 40252 36546 40308 36548
rect 40252 36494 40254 36546
rect 40254 36494 40306 36546
rect 40306 36494 40308 36546
rect 40252 36492 40308 36494
rect 40412 36546 40468 36548
rect 40412 36494 40414 36546
rect 40414 36494 40466 36546
rect 40466 36494 40468 36546
rect 40412 36492 40468 36494
rect 40572 36546 40628 36548
rect 40572 36494 40574 36546
rect 40574 36494 40626 36546
rect 40626 36494 40628 36546
rect 40572 36492 40628 36494
rect 40732 36546 40788 36548
rect 40732 36494 40734 36546
rect 40734 36494 40786 36546
rect 40786 36494 40788 36546
rect 40732 36492 40788 36494
rect 40892 36546 40948 36548
rect 40892 36494 40894 36546
rect 40894 36494 40946 36546
rect 40946 36494 40948 36546
rect 40892 36492 40948 36494
rect 41052 36546 41108 36548
rect 41052 36494 41054 36546
rect 41054 36494 41106 36546
rect 41106 36494 41108 36546
rect 41052 36492 41108 36494
rect 41212 36546 41268 36548
rect 41212 36494 41214 36546
rect 41214 36494 41266 36546
rect 41266 36494 41268 36546
rect 41212 36492 41268 36494
rect 41372 36546 41428 36548
rect 41372 36494 41374 36546
rect 41374 36494 41426 36546
rect 41426 36494 41428 36546
rect 41372 36492 41428 36494
rect 41532 36546 41588 36548
rect 41532 36494 41534 36546
rect 41534 36494 41586 36546
rect 41586 36494 41588 36546
rect 41532 36492 41588 36494
rect 41692 36546 41748 36548
rect 41692 36494 41694 36546
rect 41694 36494 41746 36546
rect 41746 36494 41748 36546
rect 41692 36492 41748 36494
rect 41852 36546 41908 36548
rect 41852 36494 41854 36546
rect 41854 36494 41906 36546
rect 41906 36494 41908 36546
rect 41852 36492 41908 36494
rect 12 36386 68 36388
rect 12 36334 14 36386
rect 14 36334 66 36386
rect 66 36334 68 36386
rect 12 36332 68 36334
rect 172 36386 228 36388
rect 172 36334 174 36386
rect 174 36334 226 36386
rect 226 36334 228 36386
rect 172 36332 228 36334
rect 332 36386 388 36388
rect 332 36334 334 36386
rect 334 36334 386 36386
rect 386 36334 388 36386
rect 332 36332 388 36334
rect 492 36386 548 36388
rect 492 36334 494 36386
rect 494 36334 546 36386
rect 546 36334 548 36386
rect 492 36332 548 36334
rect 652 36386 708 36388
rect 652 36334 654 36386
rect 654 36334 706 36386
rect 706 36334 708 36386
rect 652 36332 708 36334
rect 812 36386 868 36388
rect 812 36334 814 36386
rect 814 36334 866 36386
rect 866 36334 868 36386
rect 812 36332 868 36334
rect 972 36386 1028 36388
rect 972 36334 974 36386
rect 974 36334 1026 36386
rect 1026 36334 1028 36386
rect 972 36332 1028 36334
rect 1132 36386 1188 36388
rect 1132 36334 1134 36386
rect 1134 36334 1186 36386
rect 1186 36334 1188 36386
rect 1132 36332 1188 36334
rect 1292 36386 1348 36388
rect 1292 36334 1294 36386
rect 1294 36334 1346 36386
rect 1346 36334 1348 36386
rect 1292 36332 1348 36334
rect 1452 36386 1508 36388
rect 1452 36334 1454 36386
rect 1454 36334 1506 36386
rect 1506 36334 1508 36386
rect 1452 36332 1508 36334
rect 1612 36386 1668 36388
rect 1612 36334 1614 36386
rect 1614 36334 1666 36386
rect 1666 36334 1668 36386
rect 1612 36332 1668 36334
rect 1772 36386 1828 36388
rect 1772 36334 1774 36386
rect 1774 36334 1826 36386
rect 1826 36334 1828 36386
rect 1772 36332 1828 36334
rect 1932 36386 1988 36388
rect 1932 36334 1934 36386
rect 1934 36334 1986 36386
rect 1986 36334 1988 36386
rect 1932 36332 1988 36334
rect 2092 36386 2148 36388
rect 2092 36334 2094 36386
rect 2094 36334 2146 36386
rect 2146 36334 2148 36386
rect 2092 36332 2148 36334
rect 2252 36386 2308 36388
rect 2252 36334 2254 36386
rect 2254 36334 2306 36386
rect 2306 36334 2308 36386
rect 2252 36332 2308 36334
rect 2412 36386 2468 36388
rect 2412 36334 2414 36386
rect 2414 36334 2466 36386
rect 2466 36334 2468 36386
rect 2412 36332 2468 36334
rect 2572 36386 2628 36388
rect 2572 36334 2574 36386
rect 2574 36334 2626 36386
rect 2626 36334 2628 36386
rect 2572 36332 2628 36334
rect 2732 36386 2788 36388
rect 2732 36334 2734 36386
rect 2734 36334 2786 36386
rect 2786 36334 2788 36386
rect 2732 36332 2788 36334
rect 2892 36386 2948 36388
rect 2892 36334 2894 36386
rect 2894 36334 2946 36386
rect 2946 36334 2948 36386
rect 2892 36332 2948 36334
rect 3052 36386 3108 36388
rect 3052 36334 3054 36386
rect 3054 36334 3106 36386
rect 3106 36334 3108 36386
rect 3052 36332 3108 36334
rect 3212 36386 3268 36388
rect 3212 36334 3214 36386
rect 3214 36334 3266 36386
rect 3266 36334 3268 36386
rect 3212 36332 3268 36334
rect 3372 36386 3428 36388
rect 3372 36334 3374 36386
rect 3374 36334 3426 36386
rect 3426 36334 3428 36386
rect 3372 36332 3428 36334
rect 3532 36386 3588 36388
rect 3532 36334 3534 36386
rect 3534 36334 3586 36386
rect 3586 36334 3588 36386
rect 3532 36332 3588 36334
rect 3692 36386 3748 36388
rect 3692 36334 3694 36386
rect 3694 36334 3746 36386
rect 3746 36334 3748 36386
rect 3692 36332 3748 36334
rect 3852 36386 3908 36388
rect 3852 36334 3854 36386
rect 3854 36334 3906 36386
rect 3906 36334 3908 36386
rect 3852 36332 3908 36334
rect 4012 36386 4068 36388
rect 4012 36334 4014 36386
rect 4014 36334 4066 36386
rect 4066 36334 4068 36386
rect 4012 36332 4068 36334
rect 4172 36386 4228 36388
rect 4172 36334 4174 36386
rect 4174 36334 4226 36386
rect 4226 36334 4228 36386
rect 4172 36332 4228 36334
rect 4332 36386 4388 36388
rect 4332 36334 4334 36386
rect 4334 36334 4386 36386
rect 4386 36334 4388 36386
rect 4332 36332 4388 36334
rect 4492 36386 4548 36388
rect 4492 36334 4494 36386
rect 4494 36334 4546 36386
rect 4546 36334 4548 36386
rect 4492 36332 4548 36334
rect 4652 36386 4708 36388
rect 4652 36334 4654 36386
rect 4654 36334 4706 36386
rect 4706 36334 4708 36386
rect 4652 36332 4708 36334
rect 4812 36386 4868 36388
rect 4812 36334 4814 36386
rect 4814 36334 4866 36386
rect 4866 36334 4868 36386
rect 4812 36332 4868 36334
rect 4972 36386 5028 36388
rect 4972 36334 4974 36386
rect 4974 36334 5026 36386
rect 5026 36334 5028 36386
rect 4972 36332 5028 36334
rect 5132 36386 5188 36388
rect 5132 36334 5134 36386
rect 5134 36334 5186 36386
rect 5186 36334 5188 36386
rect 5132 36332 5188 36334
rect 5292 36386 5348 36388
rect 5292 36334 5294 36386
rect 5294 36334 5346 36386
rect 5346 36334 5348 36386
rect 5292 36332 5348 36334
rect 5452 36386 5508 36388
rect 5452 36334 5454 36386
rect 5454 36334 5506 36386
rect 5506 36334 5508 36386
rect 5452 36332 5508 36334
rect 5612 36386 5668 36388
rect 5612 36334 5614 36386
rect 5614 36334 5666 36386
rect 5666 36334 5668 36386
rect 5612 36332 5668 36334
rect 5772 36386 5828 36388
rect 5772 36334 5774 36386
rect 5774 36334 5826 36386
rect 5826 36334 5828 36386
rect 5772 36332 5828 36334
rect 5932 36386 5988 36388
rect 5932 36334 5934 36386
rect 5934 36334 5986 36386
rect 5986 36334 5988 36386
rect 5932 36332 5988 36334
rect 6092 36386 6148 36388
rect 6092 36334 6094 36386
rect 6094 36334 6146 36386
rect 6146 36334 6148 36386
rect 6092 36332 6148 36334
rect 6252 36386 6308 36388
rect 6252 36334 6254 36386
rect 6254 36334 6306 36386
rect 6306 36334 6308 36386
rect 6252 36332 6308 36334
rect 6412 36386 6468 36388
rect 6412 36334 6414 36386
rect 6414 36334 6466 36386
rect 6466 36334 6468 36386
rect 6412 36332 6468 36334
rect 6572 36386 6628 36388
rect 6572 36334 6574 36386
rect 6574 36334 6626 36386
rect 6626 36334 6628 36386
rect 6572 36332 6628 36334
rect 6732 36386 6788 36388
rect 6732 36334 6734 36386
rect 6734 36334 6786 36386
rect 6786 36334 6788 36386
rect 6732 36332 6788 36334
rect 6892 36386 6948 36388
rect 6892 36334 6894 36386
rect 6894 36334 6946 36386
rect 6946 36334 6948 36386
rect 6892 36332 6948 36334
rect 7052 36386 7108 36388
rect 7052 36334 7054 36386
rect 7054 36334 7106 36386
rect 7106 36334 7108 36386
rect 7052 36332 7108 36334
rect 7212 36386 7268 36388
rect 7212 36334 7214 36386
rect 7214 36334 7266 36386
rect 7266 36334 7268 36386
rect 7212 36332 7268 36334
rect 7372 36386 7428 36388
rect 7372 36334 7374 36386
rect 7374 36334 7426 36386
rect 7426 36334 7428 36386
rect 7372 36332 7428 36334
rect 7532 36386 7588 36388
rect 7532 36334 7534 36386
rect 7534 36334 7586 36386
rect 7586 36334 7588 36386
rect 7532 36332 7588 36334
rect 7692 36386 7748 36388
rect 7692 36334 7694 36386
rect 7694 36334 7746 36386
rect 7746 36334 7748 36386
rect 7692 36332 7748 36334
rect 7852 36386 7908 36388
rect 7852 36334 7854 36386
rect 7854 36334 7906 36386
rect 7906 36334 7908 36386
rect 7852 36332 7908 36334
rect 8012 36386 8068 36388
rect 8012 36334 8014 36386
rect 8014 36334 8066 36386
rect 8066 36334 8068 36386
rect 8012 36332 8068 36334
rect 8172 36386 8228 36388
rect 8172 36334 8174 36386
rect 8174 36334 8226 36386
rect 8226 36334 8228 36386
rect 8172 36332 8228 36334
rect 8332 36386 8388 36388
rect 8332 36334 8334 36386
rect 8334 36334 8386 36386
rect 8386 36334 8388 36386
rect 8332 36332 8388 36334
rect 9452 36332 9508 36388
rect 9772 36332 9828 36388
rect 10092 36332 10148 36388
rect 10412 36332 10468 36388
rect 10732 36332 10788 36388
rect 11052 36332 11108 36388
rect 11372 36332 11428 36388
rect 12492 36386 12548 36388
rect 12492 36334 12494 36386
rect 12494 36334 12546 36386
rect 12546 36334 12548 36386
rect 12492 36332 12548 36334
rect 12652 36386 12708 36388
rect 12652 36334 12654 36386
rect 12654 36334 12706 36386
rect 12706 36334 12708 36386
rect 12652 36332 12708 36334
rect 12812 36386 12868 36388
rect 12812 36334 12814 36386
rect 12814 36334 12866 36386
rect 12866 36334 12868 36386
rect 12812 36332 12868 36334
rect 12972 36386 13028 36388
rect 12972 36334 12974 36386
rect 12974 36334 13026 36386
rect 13026 36334 13028 36386
rect 12972 36332 13028 36334
rect 13132 36386 13188 36388
rect 13132 36334 13134 36386
rect 13134 36334 13186 36386
rect 13186 36334 13188 36386
rect 13132 36332 13188 36334
rect 13292 36386 13348 36388
rect 13292 36334 13294 36386
rect 13294 36334 13346 36386
rect 13346 36334 13348 36386
rect 13292 36332 13348 36334
rect 13452 36386 13508 36388
rect 13452 36334 13454 36386
rect 13454 36334 13506 36386
rect 13506 36334 13508 36386
rect 13452 36332 13508 36334
rect 13612 36386 13668 36388
rect 13612 36334 13614 36386
rect 13614 36334 13666 36386
rect 13666 36334 13668 36386
rect 13612 36332 13668 36334
rect 13772 36386 13828 36388
rect 13772 36334 13774 36386
rect 13774 36334 13826 36386
rect 13826 36334 13828 36386
rect 13772 36332 13828 36334
rect 13932 36386 13988 36388
rect 13932 36334 13934 36386
rect 13934 36334 13986 36386
rect 13986 36334 13988 36386
rect 13932 36332 13988 36334
rect 14092 36386 14148 36388
rect 14092 36334 14094 36386
rect 14094 36334 14146 36386
rect 14146 36334 14148 36386
rect 14092 36332 14148 36334
rect 14252 36386 14308 36388
rect 14252 36334 14254 36386
rect 14254 36334 14306 36386
rect 14306 36334 14308 36386
rect 14252 36332 14308 36334
rect 14412 36386 14468 36388
rect 14412 36334 14414 36386
rect 14414 36334 14466 36386
rect 14466 36334 14468 36386
rect 14412 36332 14468 36334
rect 14572 36386 14628 36388
rect 14572 36334 14574 36386
rect 14574 36334 14626 36386
rect 14626 36334 14628 36386
rect 14572 36332 14628 36334
rect 14732 36386 14788 36388
rect 14732 36334 14734 36386
rect 14734 36334 14786 36386
rect 14786 36334 14788 36386
rect 14732 36332 14788 36334
rect 14892 36386 14948 36388
rect 14892 36334 14894 36386
rect 14894 36334 14946 36386
rect 14946 36334 14948 36386
rect 14892 36332 14948 36334
rect 15052 36386 15108 36388
rect 15052 36334 15054 36386
rect 15054 36334 15106 36386
rect 15106 36334 15108 36386
rect 15052 36332 15108 36334
rect 15212 36386 15268 36388
rect 15212 36334 15214 36386
rect 15214 36334 15266 36386
rect 15266 36334 15268 36386
rect 15212 36332 15268 36334
rect 15372 36386 15428 36388
rect 15372 36334 15374 36386
rect 15374 36334 15426 36386
rect 15426 36334 15428 36386
rect 15372 36332 15428 36334
rect 15532 36386 15588 36388
rect 15532 36334 15534 36386
rect 15534 36334 15586 36386
rect 15586 36334 15588 36386
rect 15532 36332 15588 36334
rect 15692 36386 15748 36388
rect 15692 36334 15694 36386
rect 15694 36334 15746 36386
rect 15746 36334 15748 36386
rect 15692 36332 15748 36334
rect 15852 36386 15908 36388
rect 15852 36334 15854 36386
rect 15854 36334 15906 36386
rect 15906 36334 15908 36386
rect 15852 36332 15908 36334
rect 16012 36386 16068 36388
rect 16012 36334 16014 36386
rect 16014 36334 16066 36386
rect 16066 36334 16068 36386
rect 16012 36332 16068 36334
rect 16172 36386 16228 36388
rect 16172 36334 16174 36386
rect 16174 36334 16226 36386
rect 16226 36334 16228 36386
rect 16172 36332 16228 36334
rect 16332 36386 16388 36388
rect 16332 36334 16334 36386
rect 16334 36334 16386 36386
rect 16386 36334 16388 36386
rect 16332 36332 16388 36334
rect 16492 36386 16548 36388
rect 16492 36334 16494 36386
rect 16494 36334 16546 36386
rect 16546 36334 16548 36386
rect 16492 36332 16548 36334
rect 16652 36386 16708 36388
rect 16652 36334 16654 36386
rect 16654 36334 16706 36386
rect 16706 36334 16708 36386
rect 16652 36332 16708 36334
rect 16812 36386 16868 36388
rect 16812 36334 16814 36386
rect 16814 36334 16866 36386
rect 16866 36334 16868 36386
rect 16812 36332 16868 36334
rect 16972 36386 17028 36388
rect 16972 36334 16974 36386
rect 16974 36334 17026 36386
rect 17026 36334 17028 36386
rect 16972 36332 17028 36334
rect 17132 36386 17188 36388
rect 17132 36334 17134 36386
rect 17134 36334 17186 36386
rect 17186 36334 17188 36386
rect 17132 36332 17188 36334
rect 17292 36386 17348 36388
rect 17292 36334 17294 36386
rect 17294 36334 17346 36386
rect 17346 36334 17348 36386
rect 17292 36332 17348 36334
rect 17452 36386 17508 36388
rect 17452 36334 17454 36386
rect 17454 36334 17506 36386
rect 17506 36334 17508 36386
rect 17452 36332 17508 36334
rect 17612 36386 17668 36388
rect 17612 36334 17614 36386
rect 17614 36334 17666 36386
rect 17666 36334 17668 36386
rect 17612 36332 17668 36334
rect 17772 36386 17828 36388
rect 17772 36334 17774 36386
rect 17774 36334 17826 36386
rect 17826 36334 17828 36386
rect 17772 36332 17828 36334
rect 17932 36386 17988 36388
rect 17932 36334 17934 36386
rect 17934 36334 17986 36386
rect 17986 36334 17988 36386
rect 17932 36332 17988 36334
rect 18092 36386 18148 36388
rect 18092 36334 18094 36386
rect 18094 36334 18146 36386
rect 18146 36334 18148 36386
rect 18092 36332 18148 36334
rect 18252 36386 18308 36388
rect 18252 36334 18254 36386
rect 18254 36334 18306 36386
rect 18306 36334 18308 36386
rect 18252 36332 18308 36334
rect 18412 36386 18468 36388
rect 18412 36334 18414 36386
rect 18414 36334 18466 36386
rect 18466 36334 18468 36386
rect 18412 36332 18468 36334
rect 18572 36386 18628 36388
rect 18572 36334 18574 36386
rect 18574 36334 18626 36386
rect 18626 36334 18628 36386
rect 18572 36332 18628 36334
rect 18732 36386 18788 36388
rect 18732 36334 18734 36386
rect 18734 36334 18786 36386
rect 18786 36334 18788 36386
rect 18732 36332 18788 36334
rect 18892 36386 18948 36388
rect 18892 36334 18894 36386
rect 18894 36334 18946 36386
rect 18946 36334 18948 36386
rect 18892 36332 18948 36334
rect 20012 36332 20068 36388
rect 20332 36332 20388 36388
rect 20652 36332 20708 36388
rect 20972 36332 21028 36388
rect 21292 36332 21348 36388
rect 21612 36332 21668 36388
rect 21932 36332 21988 36388
rect 23132 36386 23188 36388
rect 23132 36334 23134 36386
rect 23134 36334 23186 36386
rect 23186 36334 23188 36386
rect 23132 36332 23188 36334
rect 23292 36386 23348 36388
rect 23292 36334 23294 36386
rect 23294 36334 23346 36386
rect 23346 36334 23348 36386
rect 23292 36332 23348 36334
rect 23452 36386 23508 36388
rect 23452 36334 23454 36386
rect 23454 36334 23506 36386
rect 23506 36334 23508 36386
rect 23452 36332 23508 36334
rect 23612 36386 23668 36388
rect 23612 36334 23614 36386
rect 23614 36334 23666 36386
rect 23666 36334 23668 36386
rect 23612 36332 23668 36334
rect 23772 36386 23828 36388
rect 23772 36334 23774 36386
rect 23774 36334 23826 36386
rect 23826 36334 23828 36386
rect 23772 36332 23828 36334
rect 23932 36386 23988 36388
rect 23932 36334 23934 36386
rect 23934 36334 23986 36386
rect 23986 36334 23988 36386
rect 23932 36332 23988 36334
rect 24092 36386 24148 36388
rect 24092 36334 24094 36386
rect 24094 36334 24146 36386
rect 24146 36334 24148 36386
rect 24092 36332 24148 36334
rect 24252 36386 24308 36388
rect 24252 36334 24254 36386
rect 24254 36334 24306 36386
rect 24306 36334 24308 36386
rect 24252 36332 24308 36334
rect 24412 36386 24468 36388
rect 24412 36334 24414 36386
rect 24414 36334 24466 36386
rect 24466 36334 24468 36386
rect 24412 36332 24468 36334
rect 24572 36386 24628 36388
rect 24572 36334 24574 36386
rect 24574 36334 24626 36386
rect 24626 36334 24628 36386
rect 24572 36332 24628 36334
rect 24732 36386 24788 36388
rect 24732 36334 24734 36386
rect 24734 36334 24786 36386
rect 24786 36334 24788 36386
rect 24732 36332 24788 36334
rect 24892 36386 24948 36388
rect 24892 36334 24894 36386
rect 24894 36334 24946 36386
rect 24946 36334 24948 36386
rect 24892 36332 24948 36334
rect 25052 36386 25108 36388
rect 25052 36334 25054 36386
rect 25054 36334 25106 36386
rect 25106 36334 25108 36386
rect 25052 36332 25108 36334
rect 25212 36386 25268 36388
rect 25212 36334 25214 36386
rect 25214 36334 25266 36386
rect 25266 36334 25268 36386
rect 25212 36332 25268 36334
rect 25372 36386 25428 36388
rect 25372 36334 25374 36386
rect 25374 36334 25426 36386
rect 25426 36334 25428 36386
rect 25372 36332 25428 36334
rect 25532 36386 25588 36388
rect 25532 36334 25534 36386
rect 25534 36334 25586 36386
rect 25586 36334 25588 36386
rect 25532 36332 25588 36334
rect 25692 36386 25748 36388
rect 25692 36334 25694 36386
rect 25694 36334 25746 36386
rect 25746 36334 25748 36386
rect 25692 36332 25748 36334
rect 25852 36386 25908 36388
rect 25852 36334 25854 36386
rect 25854 36334 25906 36386
rect 25906 36334 25908 36386
rect 25852 36332 25908 36334
rect 26012 36386 26068 36388
rect 26012 36334 26014 36386
rect 26014 36334 26066 36386
rect 26066 36334 26068 36386
rect 26012 36332 26068 36334
rect 26172 36386 26228 36388
rect 26172 36334 26174 36386
rect 26174 36334 26226 36386
rect 26226 36334 26228 36386
rect 26172 36332 26228 36334
rect 26332 36386 26388 36388
rect 26332 36334 26334 36386
rect 26334 36334 26386 36386
rect 26386 36334 26388 36386
rect 26332 36332 26388 36334
rect 26492 36386 26548 36388
rect 26492 36334 26494 36386
rect 26494 36334 26546 36386
rect 26546 36334 26548 36386
rect 26492 36332 26548 36334
rect 26652 36386 26708 36388
rect 26652 36334 26654 36386
rect 26654 36334 26706 36386
rect 26706 36334 26708 36386
rect 26652 36332 26708 36334
rect 26812 36386 26868 36388
rect 26812 36334 26814 36386
rect 26814 36334 26866 36386
rect 26866 36334 26868 36386
rect 26812 36332 26868 36334
rect 26972 36386 27028 36388
rect 26972 36334 26974 36386
rect 26974 36334 27026 36386
rect 27026 36334 27028 36386
rect 26972 36332 27028 36334
rect 27132 36386 27188 36388
rect 27132 36334 27134 36386
rect 27134 36334 27186 36386
rect 27186 36334 27188 36386
rect 27132 36332 27188 36334
rect 27292 36386 27348 36388
rect 27292 36334 27294 36386
rect 27294 36334 27346 36386
rect 27346 36334 27348 36386
rect 27292 36332 27348 36334
rect 27452 36386 27508 36388
rect 27452 36334 27454 36386
rect 27454 36334 27506 36386
rect 27506 36334 27508 36386
rect 27452 36332 27508 36334
rect 27612 36386 27668 36388
rect 27612 36334 27614 36386
rect 27614 36334 27666 36386
rect 27666 36334 27668 36386
rect 27612 36332 27668 36334
rect 27772 36386 27828 36388
rect 27772 36334 27774 36386
rect 27774 36334 27826 36386
rect 27826 36334 27828 36386
rect 27772 36332 27828 36334
rect 27932 36386 27988 36388
rect 27932 36334 27934 36386
rect 27934 36334 27986 36386
rect 27986 36334 27988 36386
rect 27932 36332 27988 36334
rect 28092 36386 28148 36388
rect 28092 36334 28094 36386
rect 28094 36334 28146 36386
rect 28146 36334 28148 36386
rect 28092 36332 28148 36334
rect 28252 36386 28308 36388
rect 28252 36334 28254 36386
rect 28254 36334 28306 36386
rect 28306 36334 28308 36386
rect 28252 36332 28308 36334
rect 28412 36386 28468 36388
rect 28412 36334 28414 36386
rect 28414 36334 28466 36386
rect 28466 36334 28468 36386
rect 28412 36332 28468 36334
rect 28572 36386 28628 36388
rect 28572 36334 28574 36386
rect 28574 36334 28626 36386
rect 28626 36334 28628 36386
rect 28572 36332 28628 36334
rect 28732 36386 28788 36388
rect 28732 36334 28734 36386
rect 28734 36334 28786 36386
rect 28786 36334 28788 36386
rect 28732 36332 28788 36334
rect 28892 36386 28948 36388
rect 28892 36334 28894 36386
rect 28894 36334 28946 36386
rect 28946 36334 28948 36386
rect 28892 36332 28948 36334
rect 29052 36386 29108 36388
rect 29052 36334 29054 36386
rect 29054 36334 29106 36386
rect 29106 36334 29108 36386
rect 29052 36332 29108 36334
rect 29212 36386 29268 36388
rect 29212 36334 29214 36386
rect 29214 36334 29266 36386
rect 29266 36334 29268 36386
rect 29212 36332 29268 36334
rect 29372 36386 29428 36388
rect 29372 36334 29374 36386
rect 29374 36334 29426 36386
rect 29426 36334 29428 36386
rect 29372 36332 29428 36334
rect 30492 36332 30548 36388
rect 30812 36332 30868 36388
rect 31132 36332 31188 36388
rect 31452 36332 31508 36388
rect 31772 36332 31828 36388
rect 32092 36332 32148 36388
rect 32412 36332 32468 36388
rect 33532 36386 33588 36388
rect 33532 36334 33534 36386
rect 33534 36334 33586 36386
rect 33586 36334 33588 36386
rect 33532 36332 33588 36334
rect 33692 36386 33748 36388
rect 33692 36334 33694 36386
rect 33694 36334 33746 36386
rect 33746 36334 33748 36386
rect 33692 36332 33748 36334
rect 33852 36386 33908 36388
rect 33852 36334 33854 36386
rect 33854 36334 33906 36386
rect 33906 36334 33908 36386
rect 33852 36332 33908 36334
rect 34012 36386 34068 36388
rect 34012 36334 34014 36386
rect 34014 36334 34066 36386
rect 34066 36334 34068 36386
rect 34012 36332 34068 36334
rect 34172 36386 34228 36388
rect 34172 36334 34174 36386
rect 34174 36334 34226 36386
rect 34226 36334 34228 36386
rect 34172 36332 34228 36334
rect 34332 36386 34388 36388
rect 34332 36334 34334 36386
rect 34334 36334 34386 36386
rect 34386 36334 34388 36386
rect 34332 36332 34388 36334
rect 34492 36386 34548 36388
rect 34492 36334 34494 36386
rect 34494 36334 34546 36386
rect 34546 36334 34548 36386
rect 34492 36332 34548 36334
rect 34652 36386 34708 36388
rect 34652 36334 34654 36386
rect 34654 36334 34706 36386
rect 34706 36334 34708 36386
rect 34652 36332 34708 36334
rect 34812 36386 34868 36388
rect 34812 36334 34814 36386
rect 34814 36334 34866 36386
rect 34866 36334 34868 36386
rect 34812 36332 34868 36334
rect 34972 36386 35028 36388
rect 34972 36334 34974 36386
rect 34974 36334 35026 36386
rect 35026 36334 35028 36386
rect 34972 36332 35028 36334
rect 35132 36386 35188 36388
rect 35132 36334 35134 36386
rect 35134 36334 35186 36386
rect 35186 36334 35188 36386
rect 35132 36332 35188 36334
rect 35292 36386 35348 36388
rect 35292 36334 35294 36386
rect 35294 36334 35346 36386
rect 35346 36334 35348 36386
rect 35292 36332 35348 36334
rect 35452 36386 35508 36388
rect 35452 36334 35454 36386
rect 35454 36334 35506 36386
rect 35506 36334 35508 36386
rect 35452 36332 35508 36334
rect 35612 36386 35668 36388
rect 35612 36334 35614 36386
rect 35614 36334 35666 36386
rect 35666 36334 35668 36386
rect 35612 36332 35668 36334
rect 35772 36386 35828 36388
rect 35772 36334 35774 36386
rect 35774 36334 35826 36386
rect 35826 36334 35828 36386
rect 35772 36332 35828 36334
rect 35932 36386 35988 36388
rect 35932 36334 35934 36386
rect 35934 36334 35986 36386
rect 35986 36334 35988 36386
rect 35932 36332 35988 36334
rect 36092 36386 36148 36388
rect 36092 36334 36094 36386
rect 36094 36334 36146 36386
rect 36146 36334 36148 36386
rect 36092 36332 36148 36334
rect 36252 36386 36308 36388
rect 36252 36334 36254 36386
rect 36254 36334 36306 36386
rect 36306 36334 36308 36386
rect 36252 36332 36308 36334
rect 36412 36386 36468 36388
rect 36412 36334 36414 36386
rect 36414 36334 36466 36386
rect 36466 36334 36468 36386
rect 36412 36332 36468 36334
rect 36572 36386 36628 36388
rect 36572 36334 36574 36386
rect 36574 36334 36626 36386
rect 36626 36334 36628 36386
rect 36572 36332 36628 36334
rect 36732 36386 36788 36388
rect 36732 36334 36734 36386
rect 36734 36334 36786 36386
rect 36786 36334 36788 36386
rect 36732 36332 36788 36334
rect 36892 36386 36948 36388
rect 36892 36334 36894 36386
rect 36894 36334 36946 36386
rect 36946 36334 36948 36386
rect 36892 36332 36948 36334
rect 37052 36386 37108 36388
rect 37052 36334 37054 36386
rect 37054 36334 37106 36386
rect 37106 36334 37108 36386
rect 37052 36332 37108 36334
rect 37212 36386 37268 36388
rect 37212 36334 37214 36386
rect 37214 36334 37266 36386
rect 37266 36334 37268 36386
rect 37212 36332 37268 36334
rect 37372 36386 37428 36388
rect 37372 36334 37374 36386
rect 37374 36334 37426 36386
rect 37426 36334 37428 36386
rect 37372 36332 37428 36334
rect 37532 36386 37588 36388
rect 37532 36334 37534 36386
rect 37534 36334 37586 36386
rect 37586 36334 37588 36386
rect 37532 36332 37588 36334
rect 37692 36386 37748 36388
rect 37692 36334 37694 36386
rect 37694 36334 37746 36386
rect 37746 36334 37748 36386
rect 37692 36332 37748 36334
rect 37852 36386 37908 36388
rect 37852 36334 37854 36386
rect 37854 36334 37906 36386
rect 37906 36334 37908 36386
rect 37852 36332 37908 36334
rect 38012 36386 38068 36388
rect 38012 36334 38014 36386
rect 38014 36334 38066 36386
rect 38066 36334 38068 36386
rect 38012 36332 38068 36334
rect 38172 36386 38228 36388
rect 38172 36334 38174 36386
rect 38174 36334 38226 36386
rect 38226 36334 38228 36386
rect 38172 36332 38228 36334
rect 38332 36386 38388 36388
rect 38332 36334 38334 36386
rect 38334 36334 38386 36386
rect 38386 36334 38388 36386
rect 38332 36332 38388 36334
rect 38492 36386 38548 36388
rect 38492 36334 38494 36386
rect 38494 36334 38546 36386
rect 38546 36334 38548 36386
rect 38492 36332 38548 36334
rect 38652 36386 38708 36388
rect 38652 36334 38654 36386
rect 38654 36334 38706 36386
rect 38706 36334 38708 36386
rect 38652 36332 38708 36334
rect 38812 36386 38868 36388
rect 38812 36334 38814 36386
rect 38814 36334 38866 36386
rect 38866 36334 38868 36386
rect 38812 36332 38868 36334
rect 38972 36386 39028 36388
rect 38972 36334 38974 36386
rect 38974 36334 39026 36386
rect 39026 36334 39028 36386
rect 38972 36332 39028 36334
rect 39132 36386 39188 36388
rect 39132 36334 39134 36386
rect 39134 36334 39186 36386
rect 39186 36334 39188 36386
rect 39132 36332 39188 36334
rect 39292 36386 39348 36388
rect 39292 36334 39294 36386
rect 39294 36334 39346 36386
rect 39346 36334 39348 36386
rect 39292 36332 39348 36334
rect 39452 36386 39508 36388
rect 39452 36334 39454 36386
rect 39454 36334 39506 36386
rect 39506 36334 39508 36386
rect 39452 36332 39508 36334
rect 39612 36386 39668 36388
rect 39612 36334 39614 36386
rect 39614 36334 39666 36386
rect 39666 36334 39668 36386
rect 39612 36332 39668 36334
rect 39772 36386 39828 36388
rect 39772 36334 39774 36386
rect 39774 36334 39826 36386
rect 39826 36334 39828 36386
rect 39772 36332 39828 36334
rect 39932 36386 39988 36388
rect 39932 36334 39934 36386
rect 39934 36334 39986 36386
rect 39986 36334 39988 36386
rect 39932 36332 39988 36334
rect 40092 36386 40148 36388
rect 40092 36334 40094 36386
rect 40094 36334 40146 36386
rect 40146 36334 40148 36386
rect 40092 36332 40148 36334
rect 40252 36386 40308 36388
rect 40252 36334 40254 36386
rect 40254 36334 40306 36386
rect 40306 36334 40308 36386
rect 40252 36332 40308 36334
rect 40412 36386 40468 36388
rect 40412 36334 40414 36386
rect 40414 36334 40466 36386
rect 40466 36334 40468 36386
rect 40412 36332 40468 36334
rect 40572 36386 40628 36388
rect 40572 36334 40574 36386
rect 40574 36334 40626 36386
rect 40626 36334 40628 36386
rect 40572 36332 40628 36334
rect 40732 36386 40788 36388
rect 40732 36334 40734 36386
rect 40734 36334 40786 36386
rect 40786 36334 40788 36386
rect 40732 36332 40788 36334
rect 40892 36386 40948 36388
rect 40892 36334 40894 36386
rect 40894 36334 40946 36386
rect 40946 36334 40948 36386
rect 40892 36332 40948 36334
rect 41052 36386 41108 36388
rect 41052 36334 41054 36386
rect 41054 36334 41106 36386
rect 41106 36334 41108 36386
rect 41052 36332 41108 36334
rect 41212 36386 41268 36388
rect 41212 36334 41214 36386
rect 41214 36334 41266 36386
rect 41266 36334 41268 36386
rect 41212 36332 41268 36334
rect 41372 36386 41428 36388
rect 41372 36334 41374 36386
rect 41374 36334 41426 36386
rect 41426 36334 41428 36386
rect 41372 36332 41428 36334
rect 41532 36386 41588 36388
rect 41532 36334 41534 36386
rect 41534 36334 41586 36386
rect 41586 36334 41588 36386
rect 41532 36332 41588 36334
rect 41692 36386 41748 36388
rect 41692 36334 41694 36386
rect 41694 36334 41746 36386
rect 41746 36334 41748 36386
rect 41692 36332 41748 36334
rect 41852 36386 41908 36388
rect 41852 36334 41854 36386
rect 41854 36334 41906 36386
rect 41906 36334 41908 36386
rect 41852 36332 41908 36334
rect 9612 36172 9668 36228
rect 21772 36172 21828 36228
rect 32252 36172 32308 36228
rect 12 36066 68 36068
rect 12 36014 14 36066
rect 14 36014 66 36066
rect 66 36014 68 36066
rect 12 36012 68 36014
rect 172 36066 228 36068
rect 172 36014 174 36066
rect 174 36014 226 36066
rect 226 36014 228 36066
rect 172 36012 228 36014
rect 332 36066 388 36068
rect 332 36014 334 36066
rect 334 36014 386 36066
rect 386 36014 388 36066
rect 332 36012 388 36014
rect 492 36066 548 36068
rect 492 36014 494 36066
rect 494 36014 546 36066
rect 546 36014 548 36066
rect 492 36012 548 36014
rect 652 36066 708 36068
rect 652 36014 654 36066
rect 654 36014 706 36066
rect 706 36014 708 36066
rect 652 36012 708 36014
rect 812 36066 868 36068
rect 812 36014 814 36066
rect 814 36014 866 36066
rect 866 36014 868 36066
rect 812 36012 868 36014
rect 972 36066 1028 36068
rect 972 36014 974 36066
rect 974 36014 1026 36066
rect 1026 36014 1028 36066
rect 972 36012 1028 36014
rect 1132 36066 1188 36068
rect 1132 36014 1134 36066
rect 1134 36014 1186 36066
rect 1186 36014 1188 36066
rect 1132 36012 1188 36014
rect 1292 36066 1348 36068
rect 1292 36014 1294 36066
rect 1294 36014 1346 36066
rect 1346 36014 1348 36066
rect 1292 36012 1348 36014
rect 1452 36066 1508 36068
rect 1452 36014 1454 36066
rect 1454 36014 1506 36066
rect 1506 36014 1508 36066
rect 1452 36012 1508 36014
rect 1612 36066 1668 36068
rect 1612 36014 1614 36066
rect 1614 36014 1666 36066
rect 1666 36014 1668 36066
rect 1612 36012 1668 36014
rect 1772 36066 1828 36068
rect 1772 36014 1774 36066
rect 1774 36014 1826 36066
rect 1826 36014 1828 36066
rect 1772 36012 1828 36014
rect 1932 36066 1988 36068
rect 1932 36014 1934 36066
rect 1934 36014 1986 36066
rect 1986 36014 1988 36066
rect 1932 36012 1988 36014
rect 2092 36066 2148 36068
rect 2092 36014 2094 36066
rect 2094 36014 2146 36066
rect 2146 36014 2148 36066
rect 2092 36012 2148 36014
rect 2252 36066 2308 36068
rect 2252 36014 2254 36066
rect 2254 36014 2306 36066
rect 2306 36014 2308 36066
rect 2252 36012 2308 36014
rect 2412 36066 2468 36068
rect 2412 36014 2414 36066
rect 2414 36014 2466 36066
rect 2466 36014 2468 36066
rect 2412 36012 2468 36014
rect 2572 36066 2628 36068
rect 2572 36014 2574 36066
rect 2574 36014 2626 36066
rect 2626 36014 2628 36066
rect 2572 36012 2628 36014
rect 2732 36066 2788 36068
rect 2732 36014 2734 36066
rect 2734 36014 2786 36066
rect 2786 36014 2788 36066
rect 2732 36012 2788 36014
rect 2892 36066 2948 36068
rect 2892 36014 2894 36066
rect 2894 36014 2946 36066
rect 2946 36014 2948 36066
rect 2892 36012 2948 36014
rect 3052 36066 3108 36068
rect 3052 36014 3054 36066
rect 3054 36014 3106 36066
rect 3106 36014 3108 36066
rect 3052 36012 3108 36014
rect 3212 36066 3268 36068
rect 3212 36014 3214 36066
rect 3214 36014 3266 36066
rect 3266 36014 3268 36066
rect 3212 36012 3268 36014
rect 3372 36066 3428 36068
rect 3372 36014 3374 36066
rect 3374 36014 3426 36066
rect 3426 36014 3428 36066
rect 3372 36012 3428 36014
rect 3532 36066 3588 36068
rect 3532 36014 3534 36066
rect 3534 36014 3586 36066
rect 3586 36014 3588 36066
rect 3532 36012 3588 36014
rect 3692 36066 3748 36068
rect 3692 36014 3694 36066
rect 3694 36014 3746 36066
rect 3746 36014 3748 36066
rect 3692 36012 3748 36014
rect 3852 36066 3908 36068
rect 3852 36014 3854 36066
rect 3854 36014 3906 36066
rect 3906 36014 3908 36066
rect 3852 36012 3908 36014
rect 4012 36066 4068 36068
rect 4012 36014 4014 36066
rect 4014 36014 4066 36066
rect 4066 36014 4068 36066
rect 4012 36012 4068 36014
rect 4172 36066 4228 36068
rect 4172 36014 4174 36066
rect 4174 36014 4226 36066
rect 4226 36014 4228 36066
rect 4172 36012 4228 36014
rect 4332 36066 4388 36068
rect 4332 36014 4334 36066
rect 4334 36014 4386 36066
rect 4386 36014 4388 36066
rect 4332 36012 4388 36014
rect 4492 36066 4548 36068
rect 4492 36014 4494 36066
rect 4494 36014 4546 36066
rect 4546 36014 4548 36066
rect 4492 36012 4548 36014
rect 4652 36066 4708 36068
rect 4652 36014 4654 36066
rect 4654 36014 4706 36066
rect 4706 36014 4708 36066
rect 4652 36012 4708 36014
rect 4812 36066 4868 36068
rect 4812 36014 4814 36066
rect 4814 36014 4866 36066
rect 4866 36014 4868 36066
rect 4812 36012 4868 36014
rect 4972 36066 5028 36068
rect 4972 36014 4974 36066
rect 4974 36014 5026 36066
rect 5026 36014 5028 36066
rect 4972 36012 5028 36014
rect 5132 36066 5188 36068
rect 5132 36014 5134 36066
rect 5134 36014 5186 36066
rect 5186 36014 5188 36066
rect 5132 36012 5188 36014
rect 5292 36066 5348 36068
rect 5292 36014 5294 36066
rect 5294 36014 5346 36066
rect 5346 36014 5348 36066
rect 5292 36012 5348 36014
rect 5452 36066 5508 36068
rect 5452 36014 5454 36066
rect 5454 36014 5506 36066
rect 5506 36014 5508 36066
rect 5452 36012 5508 36014
rect 5612 36066 5668 36068
rect 5612 36014 5614 36066
rect 5614 36014 5666 36066
rect 5666 36014 5668 36066
rect 5612 36012 5668 36014
rect 5772 36066 5828 36068
rect 5772 36014 5774 36066
rect 5774 36014 5826 36066
rect 5826 36014 5828 36066
rect 5772 36012 5828 36014
rect 5932 36066 5988 36068
rect 5932 36014 5934 36066
rect 5934 36014 5986 36066
rect 5986 36014 5988 36066
rect 5932 36012 5988 36014
rect 6092 36066 6148 36068
rect 6092 36014 6094 36066
rect 6094 36014 6146 36066
rect 6146 36014 6148 36066
rect 6092 36012 6148 36014
rect 6252 36066 6308 36068
rect 6252 36014 6254 36066
rect 6254 36014 6306 36066
rect 6306 36014 6308 36066
rect 6252 36012 6308 36014
rect 6412 36066 6468 36068
rect 6412 36014 6414 36066
rect 6414 36014 6466 36066
rect 6466 36014 6468 36066
rect 6412 36012 6468 36014
rect 6572 36066 6628 36068
rect 6572 36014 6574 36066
rect 6574 36014 6626 36066
rect 6626 36014 6628 36066
rect 6572 36012 6628 36014
rect 6732 36066 6788 36068
rect 6732 36014 6734 36066
rect 6734 36014 6786 36066
rect 6786 36014 6788 36066
rect 6732 36012 6788 36014
rect 6892 36066 6948 36068
rect 6892 36014 6894 36066
rect 6894 36014 6946 36066
rect 6946 36014 6948 36066
rect 6892 36012 6948 36014
rect 7052 36066 7108 36068
rect 7052 36014 7054 36066
rect 7054 36014 7106 36066
rect 7106 36014 7108 36066
rect 7052 36012 7108 36014
rect 7212 36066 7268 36068
rect 7212 36014 7214 36066
rect 7214 36014 7266 36066
rect 7266 36014 7268 36066
rect 7212 36012 7268 36014
rect 7372 36066 7428 36068
rect 7372 36014 7374 36066
rect 7374 36014 7426 36066
rect 7426 36014 7428 36066
rect 7372 36012 7428 36014
rect 7532 36066 7588 36068
rect 7532 36014 7534 36066
rect 7534 36014 7586 36066
rect 7586 36014 7588 36066
rect 7532 36012 7588 36014
rect 7692 36066 7748 36068
rect 7692 36014 7694 36066
rect 7694 36014 7746 36066
rect 7746 36014 7748 36066
rect 7692 36012 7748 36014
rect 7852 36066 7908 36068
rect 7852 36014 7854 36066
rect 7854 36014 7906 36066
rect 7906 36014 7908 36066
rect 7852 36012 7908 36014
rect 8012 36066 8068 36068
rect 8012 36014 8014 36066
rect 8014 36014 8066 36066
rect 8066 36014 8068 36066
rect 8012 36012 8068 36014
rect 8172 36066 8228 36068
rect 8172 36014 8174 36066
rect 8174 36014 8226 36066
rect 8226 36014 8228 36066
rect 8172 36012 8228 36014
rect 8332 36066 8388 36068
rect 8332 36014 8334 36066
rect 8334 36014 8386 36066
rect 8386 36014 8388 36066
rect 8332 36012 8388 36014
rect 9452 36012 9508 36068
rect 9772 36012 9828 36068
rect 10092 36012 10148 36068
rect 10412 36012 10468 36068
rect 10732 36012 10788 36068
rect 11052 36012 11108 36068
rect 11372 36012 11428 36068
rect 12492 36066 12548 36068
rect 12492 36014 12494 36066
rect 12494 36014 12546 36066
rect 12546 36014 12548 36066
rect 12492 36012 12548 36014
rect 12652 36066 12708 36068
rect 12652 36014 12654 36066
rect 12654 36014 12706 36066
rect 12706 36014 12708 36066
rect 12652 36012 12708 36014
rect 12812 36066 12868 36068
rect 12812 36014 12814 36066
rect 12814 36014 12866 36066
rect 12866 36014 12868 36066
rect 12812 36012 12868 36014
rect 12972 36066 13028 36068
rect 12972 36014 12974 36066
rect 12974 36014 13026 36066
rect 13026 36014 13028 36066
rect 12972 36012 13028 36014
rect 13132 36066 13188 36068
rect 13132 36014 13134 36066
rect 13134 36014 13186 36066
rect 13186 36014 13188 36066
rect 13132 36012 13188 36014
rect 13292 36066 13348 36068
rect 13292 36014 13294 36066
rect 13294 36014 13346 36066
rect 13346 36014 13348 36066
rect 13292 36012 13348 36014
rect 13452 36066 13508 36068
rect 13452 36014 13454 36066
rect 13454 36014 13506 36066
rect 13506 36014 13508 36066
rect 13452 36012 13508 36014
rect 13612 36066 13668 36068
rect 13612 36014 13614 36066
rect 13614 36014 13666 36066
rect 13666 36014 13668 36066
rect 13612 36012 13668 36014
rect 13772 36066 13828 36068
rect 13772 36014 13774 36066
rect 13774 36014 13826 36066
rect 13826 36014 13828 36066
rect 13772 36012 13828 36014
rect 13932 36066 13988 36068
rect 13932 36014 13934 36066
rect 13934 36014 13986 36066
rect 13986 36014 13988 36066
rect 13932 36012 13988 36014
rect 14092 36066 14148 36068
rect 14092 36014 14094 36066
rect 14094 36014 14146 36066
rect 14146 36014 14148 36066
rect 14092 36012 14148 36014
rect 14252 36066 14308 36068
rect 14252 36014 14254 36066
rect 14254 36014 14306 36066
rect 14306 36014 14308 36066
rect 14252 36012 14308 36014
rect 14412 36066 14468 36068
rect 14412 36014 14414 36066
rect 14414 36014 14466 36066
rect 14466 36014 14468 36066
rect 14412 36012 14468 36014
rect 14572 36066 14628 36068
rect 14572 36014 14574 36066
rect 14574 36014 14626 36066
rect 14626 36014 14628 36066
rect 14572 36012 14628 36014
rect 14732 36066 14788 36068
rect 14732 36014 14734 36066
rect 14734 36014 14786 36066
rect 14786 36014 14788 36066
rect 14732 36012 14788 36014
rect 14892 36066 14948 36068
rect 14892 36014 14894 36066
rect 14894 36014 14946 36066
rect 14946 36014 14948 36066
rect 14892 36012 14948 36014
rect 15052 36066 15108 36068
rect 15052 36014 15054 36066
rect 15054 36014 15106 36066
rect 15106 36014 15108 36066
rect 15052 36012 15108 36014
rect 15212 36066 15268 36068
rect 15212 36014 15214 36066
rect 15214 36014 15266 36066
rect 15266 36014 15268 36066
rect 15212 36012 15268 36014
rect 15372 36066 15428 36068
rect 15372 36014 15374 36066
rect 15374 36014 15426 36066
rect 15426 36014 15428 36066
rect 15372 36012 15428 36014
rect 15532 36066 15588 36068
rect 15532 36014 15534 36066
rect 15534 36014 15586 36066
rect 15586 36014 15588 36066
rect 15532 36012 15588 36014
rect 15692 36066 15748 36068
rect 15692 36014 15694 36066
rect 15694 36014 15746 36066
rect 15746 36014 15748 36066
rect 15692 36012 15748 36014
rect 15852 36066 15908 36068
rect 15852 36014 15854 36066
rect 15854 36014 15906 36066
rect 15906 36014 15908 36066
rect 15852 36012 15908 36014
rect 16012 36066 16068 36068
rect 16012 36014 16014 36066
rect 16014 36014 16066 36066
rect 16066 36014 16068 36066
rect 16012 36012 16068 36014
rect 16172 36066 16228 36068
rect 16172 36014 16174 36066
rect 16174 36014 16226 36066
rect 16226 36014 16228 36066
rect 16172 36012 16228 36014
rect 16332 36066 16388 36068
rect 16332 36014 16334 36066
rect 16334 36014 16386 36066
rect 16386 36014 16388 36066
rect 16332 36012 16388 36014
rect 16492 36066 16548 36068
rect 16492 36014 16494 36066
rect 16494 36014 16546 36066
rect 16546 36014 16548 36066
rect 16492 36012 16548 36014
rect 16652 36066 16708 36068
rect 16652 36014 16654 36066
rect 16654 36014 16706 36066
rect 16706 36014 16708 36066
rect 16652 36012 16708 36014
rect 16812 36066 16868 36068
rect 16812 36014 16814 36066
rect 16814 36014 16866 36066
rect 16866 36014 16868 36066
rect 16812 36012 16868 36014
rect 16972 36066 17028 36068
rect 16972 36014 16974 36066
rect 16974 36014 17026 36066
rect 17026 36014 17028 36066
rect 16972 36012 17028 36014
rect 17132 36066 17188 36068
rect 17132 36014 17134 36066
rect 17134 36014 17186 36066
rect 17186 36014 17188 36066
rect 17132 36012 17188 36014
rect 17292 36066 17348 36068
rect 17292 36014 17294 36066
rect 17294 36014 17346 36066
rect 17346 36014 17348 36066
rect 17292 36012 17348 36014
rect 17452 36066 17508 36068
rect 17452 36014 17454 36066
rect 17454 36014 17506 36066
rect 17506 36014 17508 36066
rect 17452 36012 17508 36014
rect 17612 36066 17668 36068
rect 17612 36014 17614 36066
rect 17614 36014 17666 36066
rect 17666 36014 17668 36066
rect 17612 36012 17668 36014
rect 17772 36066 17828 36068
rect 17772 36014 17774 36066
rect 17774 36014 17826 36066
rect 17826 36014 17828 36066
rect 17772 36012 17828 36014
rect 17932 36066 17988 36068
rect 17932 36014 17934 36066
rect 17934 36014 17986 36066
rect 17986 36014 17988 36066
rect 17932 36012 17988 36014
rect 18092 36066 18148 36068
rect 18092 36014 18094 36066
rect 18094 36014 18146 36066
rect 18146 36014 18148 36066
rect 18092 36012 18148 36014
rect 18252 36066 18308 36068
rect 18252 36014 18254 36066
rect 18254 36014 18306 36066
rect 18306 36014 18308 36066
rect 18252 36012 18308 36014
rect 18412 36066 18468 36068
rect 18412 36014 18414 36066
rect 18414 36014 18466 36066
rect 18466 36014 18468 36066
rect 18412 36012 18468 36014
rect 18572 36066 18628 36068
rect 18572 36014 18574 36066
rect 18574 36014 18626 36066
rect 18626 36014 18628 36066
rect 18572 36012 18628 36014
rect 18732 36066 18788 36068
rect 18732 36014 18734 36066
rect 18734 36014 18786 36066
rect 18786 36014 18788 36066
rect 18732 36012 18788 36014
rect 18892 36066 18948 36068
rect 18892 36014 18894 36066
rect 18894 36014 18946 36066
rect 18946 36014 18948 36066
rect 18892 36012 18948 36014
rect 20012 36012 20068 36068
rect 20332 36012 20388 36068
rect 20652 36012 20708 36068
rect 20972 36012 21028 36068
rect 21292 36012 21348 36068
rect 21612 36012 21668 36068
rect 21932 36012 21988 36068
rect 23132 36066 23188 36068
rect 23132 36014 23134 36066
rect 23134 36014 23186 36066
rect 23186 36014 23188 36066
rect 23132 36012 23188 36014
rect 23292 36066 23348 36068
rect 23292 36014 23294 36066
rect 23294 36014 23346 36066
rect 23346 36014 23348 36066
rect 23292 36012 23348 36014
rect 23452 36066 23508 36068
rect 23452 36014 23454 36066
rect 23454 36014 23506 36066
rect 23506 36014 23508 36066
rect 23452 36012 23508 36014
rect 23612 36066 23668 36068
rect 23612 36014 23614 36066
rect 23614 36014 23666 36066
rect 23666 36014 23668 36066
rect 23612 36012 23668 36014
rect 23772 36066 23828 36068
rect 23772 36014 23774 36066
rect 23774 36014 23826 36066
rect 23826 36014 23828 36066
rect 23772 36012 23828 36014
rect 23932 36066 23988 36068
rect 23932 36014 23934 36066
rect 23934 36014 23986 36066
rect 23986 36014 23988 36066
rect 23932 36012 23988 36014
rect 24092 36066 24148 36068
rect 24092 36014 24094 36066
rect 24094 36014 24146 36066
rect 24146 36014 24148 36066
rect 24092 36012 24148 36014
rect 24252 36066 24308 36068
rect 24252 36014 24254 36066
rect 24254 36014 24306 36066
rect 24306 36014 24308 36066
rect 24252 36012 24308 36014
rect 24412 36066 24468 36068
rect 24412 36014 24414 36066
rect 24414 36014 24466 36066
rect 24466 36014 24468 36066
rect 24412 36012 24468 36014
rect 24572 36066 24628 36068
rect 24572 36014 24574 36066
rect 24574 36014 24626 36066
rect 24626 36014 24628 36066
rect 24572 36012 24628 36014
rect 24732 36066 24788 36068
rect 24732 36014 24734 36066
rect 24734 36014 24786 36066
rect 24786 36014 24788 36066
rect 24732 36012 24788 36014
rect 24892 36066 24948 36068
rect 24892 36014 24894 36066
rect 24894 36014 24946 36066
rect 24946 36014 24948 36066
rect 24892 36012 24948 36014
rect 25052 36066 25108 36068
rect 25052 36014 25054 36066
rect 25054 36014 25106 36066
rect 25106 36014 25108 36066
rect 25052 36012 25108 36014
rect 25212 36066 25268 36068
rect 25212 36014 25214 36066
rect 25214 36014 25266 36066
rect 25266 36014 25268 36066
rect 25212 36012 25268 36014
rect 25372 36066 25428 36068
rect 25372 36014 25374 36066
rect 25374 36014 25426 36066
rect 25426 36014 25428 36066
rect 25372 36012 25428 36014
rect 25532 36066 25588 36068
rect 25532 36014 25534 36066
rect 25534 36014 25586 36066
rect 25586 36014 25588 36066
rect 25532 36012 25588 36014
rect 25692 36066 25748 36068
rect 25692 36014 25694 36066
rect 25694 36014 25746 36066
rect 25746 36014 25748 36066
rect 25692 36012 25748 36014
rect 25852 36066 25908 36068
rect 25852 36014 25854 36066
rect 25854 36014 25906 36066
rect 25906 36014 25908 36066
rect 25852 36012 25908 36014
rect 26012 36066 26068 36068
rect 26012 36014 26014 36066
rect 26014 36014 26066 36066
rect 26066 36014 26068 36066
rect 26012 36012 26068 36014
rect 26172 36066 26228 36068
rect 26172 36014 26174 36066
rect 26174 36014 26226 36066
rect 26226 36014 26228 36066
rect 26172 36012 26228 36014
rect 26332 36066 26388 36068
rect 26332 36014 26334 36066
rect 26334 36014 26386 36066
rect 26386 36014 26388 36066
rect 26332 36012 26388 36014
rect 26492 36066 26548 36068
rect 26492 36014 26494 36066
rect 26494 36014 26546 36066
rect 26546 36014 26548 36066
rect 26492 36012 26548 36014
rect 26652 36066 26708 36068
rect 26652 36014 26654 36066
rect 26654 36014 26706 36066
rect 26706 36014 26708 36066
rect 26652 36012 26708 36014
rect 26812 36066 26868 36068
rect 26812 36014 26814 36066
rect 26814 36014 26866 36066
rect 26866 36014 26868 36066
rect 26812 36012 26868 36014
rect 26972 36066 27028 36068
rect 26972 36014 26974 36066
rect 26974 36014 27026 36066
rect 27026 36014 27028 36066
rect 26972 36012 27028 36014
rect 27132 36066 27188 36068
rect 27132 36014 27134 36066
rect 27134 36014 27186 36066
rect 27186 36014 27188 36066
rect 27132 36012 27188 36014
rect 27292 36066 27348 36068
rect 27292 36014 27294 36066
rect 27294 36014 27346 36066
rect 27346 36014 27348 36066
rect 27292 36012 27348 36014
rect 27452 36066 27508 36068
rect 27452 36014 27454 36066
rect 27454 36014 27506 36066
rect 27506 36014 27508 36066
rect 27452 36012 27508 36014
rect 27612 36066 27668 36068
rect 27612 36014 27614 36066
rect 27614 36014 27666 36066
rect 27666 36014 27668 36066
rect 27612 36012 27668 36014
rect 27772 36066 27828 36068
rect 27772 36014 27774 36066
rect 27774 36014 27826 36066
rect 27826 36014 27828 36066
rect 27772 36012 27828 36014
rect 27932 36066 27988 36068
rect 27932 36014 27934 36066
rect 27934 36014 27986 36066
rect 27986 36014 27988 36066
rect 27932 36012 27988 36014
rect 28092 36066 28148 36068
rect 28092 36014 28094 36066
rect 28094 36014 28146 36066
rect 28146 36014 28148 36066
rect 28092 36012 28148 36014
rect 28252 36066 28308 36068
rect 28252 36014 28254 36066
rect 28254 36014 28306 36066
rect 28306 36014 28308 36066
rect 28252 36012 28308 36014
rect 28412 36066 28468 36068
rect 28412 36014 28414 36066
rect 28414 36014 28466 36066
rect 28466 36014 28468 36066
rect 28412 36012 28468 36014
rect 28572 36066 28628 36068
rect 28572 36014 28574 36066
rect 28574 36014 28626 36066
rect 28626 36014 28628 36066
rect 28572 36012 28628 36014
rect 28732 36066 28788 36068
rect 28732 36014 28734 36066
rect 28734 36014 28786 36066
rect 28786 36014 28788 36066
rect 28732 36012 28788 36014
rect 28892 36066 28948 36068
rect 28892 36014 28894 36066
rect 28894 36014 28946 36066
rect 28946 36014 28948 36066
rect 28892 36012 28948 36014
rect 29052 36066 29108 36068
rect 29052 36014 29054 36066
rect 29054 36014 29106 36066
rect 29106 36014 29108 36066
rect 29052 36012 29108 36014
rect 29212 36066 29268 36068
rect 29212 36014 29214 36066
rect 29214 36014 29266 36066
rect 29266 36014 29268 36066
rect 29212 36012 29268 36014
rect 29372 36066 29428 36068
rect 29372 36014 29374 36066
rect 29374 36014 29426 36066
rect 29426 36014 29428 36066
rect 29372 36012 29428 36014
rect 30492 36012 30548 36068
rect 30812 36012 30868 36068
rect 31132 36012 31188 36068
rect 31452 36012 31508 36068
rect 31772 36012 31828 36068
rect 32092 36012 32148 36068
rect 32412 36012 32468 36068
rect 33532 36066 33588 36068
rect 33532 36014 33534 36066
rect 33534 36014 33586 36066
rect 33586 36014 33588 36066
rect 33532 36012 33588 36014
rect 33692 36066 33748 36068
rect 33692 36014 33694 36066
rect 33694 36014 33746 36066
rect 33746 36014 33748 36066
rect 33692 36012 33748 36014
rect 33852 36066 33908 36068
rect 33852 36014 33854 36066
rect 33854 36014 33906 36066
rect 33906 36014 33908 36066
rect 33852 36012 33908 36014
rect 34012 36066 34068 36068
rect 34012 36014 34014 36066
rect 34014 36014 34066 36066
rect 34066 36014 34068 36066
rect 34012 36012 34068 36014
rect 34172 36066 34228 36068
rect 34172 36014 34174 36066
rect 34174 36014 34226 36066
rect 34226 36014 34228 36066
rect 34172 36012 34228 36014
rect 34332 36066 34388 36068
rect 34332 36014 34334 36066
rect 34334 36014 34386 36066
rect 34386 36014 34388 36066
rect 34332 36012 34388 36014
rect 34492 36066 34548 36068
rect 34492 36014 34494 36066
rect 34494 36014 34546 36066
rect 34546 36014 34548 36066
rect 34492 36012 34548 36014
rect 34652 36066 34708 36068
rect 34652 36014 34654 36066
rect 34654 36014 34706 36066
rect 34706 36014 34708 36066
rect 34652 36012 34708 36014
rect 34812 36066 34868 36068
rect 34812 36014 34814 36066
rect 34814 36014 34866 36066
rect 34866 36014 34868 36066
rect 34812 36012 34868 36014
rect 34972 36066 35028 36068
rect 34972 36014 34974 36066
rect 34974 36014 35026 36066
rect 35026 36014 35028 36066
rect 34972 36012 35028 36014
rect 35132 36066 35188 36068
rect 35132 36014 35134 36066
rect 35134 36014 35186 36066
rect 35186 36014 35188 36066
rect 35132 36012 35188 36014
rect 35292 36066 35348 36068
rect 35292 36014 35294 36066
rect 35294 36014 35346 36066
rect 35346 36014 35348 36066
rect 35292 36012 35348 36014
rect 35452 36066 35508 36068
rect 35452 36014 35454 36066
rect 35454 36014 35506 36066
rect 35506 36014 35508 36066
rect 35452 36012 35508 36014
rect 35612 36066 35668 36068
rect 35612 36014 35614 36066
rect 35614 36014 35666 36066
rect 35666 36014 35668 36066
rect 35612 36012 35668 36014
rect 35772 36066 35828 36068
rect 35772 36014 35774 36066
rect 35774 36014 35826 36066
rect 35826 36014 35828 36066
rect 35772 36012 35828 36014
rect 35932 36066 35988 36068
rect 35932 36014 35934 36066
rect 35934 36014 35986 36066
rect 35986 36014 35988 36066
rect 35932 36012 35988 36014
rect 36092 36066 36148 36068
rect 36092 36014 36094 36066
rect 36094 36014 36146 36066
rect 36146 36014 36148 36066
rect 36092 36012 36148 36014
rect 36252 36066 36308 36068
rect 36252 36014 36254 36066
rect 36254 36014 36306 36066
rect 36306 36014 36308 36066
rect 36252 36012 36308 36014
rect 36412 36066 36468 36068
rect 36412 36014 36414 36066
rect 36414 36014 36466 36066
rect 36466 36014 36468 36066
rect 36412 36012 36468 36014
rect 36572 36066 36628 36068
rect 36572 36014 36574 36066
rect 36574 36014 36626 36066
rect 36626 36014 36628 36066
rect 36572 36012 36628 36014
rect 36732 36066 36788 36068
rect 36732 36014 36734 36066
rect 36734 36014 36786 36066
rect 36786 36014 36788 36066
rect 36732 36012 36788 36014
rect 36892 36066 36948 36068
rect 36892 36014 36894 36066
rect 36894 36014 36946 36066
rect 36946 36014 36948 36066
rect 36892 36012 36948 36014
rect 37052 36066 37108 36068
rect 37052 36014 37054 36066
rect 37054 36014 37106 36066
rect 37106 36014 37108 36066
rect 37052 36012 37108 36014
rect 37212 36066 37268 36068
rect 37212 36014 37214 36066
rect 37214 36014 37266 36066
rect 37266 36014 37268 36066
rect 37212 36012 37268 36014
rect 37372 36066 37428 36068
rect 37372 36014 37374 36066
rect 37374 36014 37426 36066
rect 37426 36014 37428 36066
rect 37372 36012 37428 36014
rect 37532 36066 37588 36068
rect 37532 36014 37534 36066
rect 37534 36014 37586 36066
rect 37586 36014 37588 36066
rect 37532 36012 37588 36014
rect 37692 36066 37748 36068
rect 37692 36014 37694 36066
rect 37694 36014 37746 36066
rect 37746 36014 37748 36066
rect 37692 36012 37748 36014
rect 37852 36066 37908 36068
rect 37852 36014 37854 36066
rect 37854 36014 37906 36066
rect 37906 36014 37908 36066
rect 37852 36012 37908 36014
rect 38012 36066 38068 36068
rect 38012 36014 38014 36066
rect 38014 36014 38066 36066
rect 38066 36014 38068 36066
rect 38012 36012 38068 36014
rect 38172 36066 38228 36068
rect 38172 36014 38174 36066
rect 38174 36014 38226 36066
rect 38226 36014 38228 36066
rect 38172 36012 38228 36014
rect 38332 36066 38388 36068
rect 38332 36014 38334 36066
rect 38334 36014 38386 36066
rect 38386 36014 38388 36066
rect 38332 36012 38388 36014
rect 38492 36066 38548 36068
rect 38492 36014 38494 36066
rect 38494 36014 38546 36066
rect 38546 36014 38548 36066
rect 38492 36012 38548 36014
rect 38652 36066 38708 36068
rect 38652 36014 38654 36066
rect 38654 36014 38706 36066
rect 38706 36014 38708 36066
rect 38652 36012 38708 36014
rect 38812 36066 38868 36068
rect 38812 36014 38814 36066
rect 38814 36014 38866 36066
rect 38866 36014 38868 36066
rect 38812 36012 38868 36014
rect 38972 36066 39028 36068
rect 38972 36014 38974 36066
rect 38974 36014 39026 36066
rect 39026 36014 39028 36066
rect 38972 36012 39028 36014
rect 39132 36066 39188 36068
rect 39132 36014 39134 36066
rect 39134 36014 39186 36066
rect 39186 36014 39188 36066
rect 39132 36012 39188 36014
rect 39292 36066 39348 36068
rect 39292 36014 39294 36066
rect 39294 36014 39346 36066
rect 39346 36014 39348 36066
rect 39292 36012 39348 36014
rect 39452 36066 39508 36068
rect 39452 36014 39454 36066
rect 39454 36014 39506 36066
rect 39506 36014 39508 36066
rect 39452 36012 39508 36014
rect 39612 36066 39668 36068
rect 39612 36014 39614 36066
rect 39614 36014 39666 36066
rect 39666 36014 39668 36066
rect 39612 36012 39668 36014
rect 39772 36066 39828 36068
rect 39772 36014 39774 36066
rect 39774 36014 39826 36066
rect 39826 36014 39828 36066
rect 39772 36012 39828 36014
rect 39932 36066 39988 36068
rect 39932 36014 39934 36066
rect 39934 36014 39986 36066
rect 39986 36014 39988 36066
rect 39932 36012 39988 36014
rect 40092 36066 40148 36068
rect 40092 36014 40094 36066
rect 40094 36014 40146 36066
rect 40146 36014 40148 36066
rect 40092 36012 40148 36014
rect 40252 36066 40308 36068
rect 40252 36014 40254 36066
rect 40254 36014 40306 36066
rect 40306 36014 40308 36066
rect 40252 36012 40308 36014
rect 40412 36066 40468 36068
rect 40412 36014 40414 36066
rect 40414 36014 40466 36066
rect 40466 36014 40468 36066
rect 40412 36012 40468 36014
rect 40572 36066 40628 36068
rect 40572 36014 40574 36066
rect 40574 36014 40626 36066
rect 40626 36014 40628 36066
rect 40572 36012 40628 36014
rect 40732 36066 40788 36068
rect 40732 36014 40734 36066
rect 40734 36014 40786 36066
rect 40786 36014 40788 36066
rect 40732 36012 40788 36014
rect 40892 36066 40948 36068
rect 40892 36014 40894 36066
rect 40894 36014 40946 36066
rect 40946 36014 40948 36066
rect 40892 36012 40948 36014
rect 41052 36066 41108 36068
rect 41052 36014 41054 36066
rect 41054 36014 41106 36066
rect 41106 36014 41108 36066
rect 41052 36012 41108 36014
rect 41212 36066 41268 36068
rect 41212 36014 41214 36066
rect 41214 36014 41266 36066
rect 41266 36014 41268 36066
rect 41212 36012 41268 36014
rect 41372 36066 41428 36068
rect 41372 36014 41374 36066
rect 41374 36014 41426 36066
rect 41426 36014 41428 36066
rect 41372 36012 41428 36014
rect 41532 36066 41588 36068
rect 41532 36014 41534 36066
rect 41534 36014 41586 36066
rect 41586 36014 41588 36066
rect 41532 36012 41588 36014
rect 41692 36066 41748 36068
rect 41692 36014 41694 36066
rect 41694 36014 41746 36066
rect 41746 36014 41748 36066
rect 41692 36012 41748 36014
rect 41852 36066 41908 36068
rect 41852 36014 41854 36066
rect 41854 36014 41906 36066
rect 41906 36014 41908 36066
rect 41852 36012 41908 36014
rect 9932 35852 9988 35908
rect 21452 35852 21508 35908
rect 31932 35852 31988 35908
rect 12 35746 68 35748
rect 12 35694 14 35746
rect 14 35694 66 35746
rect 66 35694 68 35746
rect 12 35692 68 35694
rect 172 35746 228 35748
rect 172 35694 174 35746
rect 174 35694 226 35746
rect 226 35694 228 35746
rect 172 35692 228 35694
rect 332 35746 388 35748
rect 332 35694 334 35746
rect 334 35694 386 35746
rect 386 35694 388 35746
rect 332 35692 388 35694
rect 492 35746 548 35748
rect 492 35694 494 35746
rect 494 35694 546 35746
rect 546 35694 548 35746
rect 492 35692 548 35694
rect 652 35746 708 35748
rect 652 35694 654 35746
rect 654 35694 706 35746
rect 706 35694 708 35746
rect 652 35692 708 35694
rect 812 35746 868 35748
rect 812 35694 814 35746
rect 814 35694 866 35746
rect 866 35694 868 35746
rect 812 35692 868 35694
rect 972 35746 1028 35748
rect 972 35694 974 35746
rect 974 35694 1026 35746
rect 1026 35694 1028 35746
rect 972 35692 1028 35694
rect 1132 35746 1188 35748
rect 1132 35694 1134 35746
rect 1134 35694 1186 35746
rect 1186 35694 1188 35746
rect 1132 35692 1188 35694
rect 1292 35746 1348 35748
rect 1292 35694 1294 35746
rect 1294 35694 1346 35746
rect 1346 35694 1348 35746
rect 1292 35692 1348 35694
rect 1452 35746 1508 35748
rect 1452 35694 1454 35746
rect 1454 35694 1506 35746
rect 1506 35694 1508 35746
rect 1452 35692 1508 35694
rect 1612 35746 1668 35748
rect 1612 35694 1614 35746
rect 1614 35694 1666 35746
rect 1666 35694 1668 35746
rect 1612 35692 1668 35694
rect 1772 35746 1828 35748
rect 1772 35694 1774 35746
rect 1774 35694 1826 35746
rect 1826 35694 1828 35746
rect 1772 35692 1828 35694
rect 1932 35746 1988 35748
rect 1932 35694 1934 35746
rect 1934 35694 1986 35746
rect 1986 35694 1988 35746
rect 1932 35692 1988 35694
rect 2092 35746 2148 35748
rect 2092 35694 2094 35746
rect 2094 35694 2146 35746
rect 2146 35694 2148 35746
rect 2092 35692 2148 35694
rect 2252 35746 2308 35748
rect 2252 35694 2254 35746
rect 2254 35694 2306 35746
rect 2306 35694 2308 35746
rect 2252 35692 2308 35694
rect 2412 35746 2468 35748
rect 2412 35694 2414 35746
rect 2414 35694 2466 35746
rect 2466 35694 2468 35746
rect 2412 35692 2468 35694
rect 2572 35746 2628 35748
rect 2572 35694 2574 35746
rect 2574 35694 2626 35746
rect 2626 35694 2628 35746
rect 2572 35692 2628 35694
rect 2732 35746 2788 35748
rect 2732 35694 2734 35746
rect 2734 35694 2786 35746
rect 2786 35694 2788 35746
rect 2732 35692 2788 35694
rect 2892 35746 2948 35748
rect 2892 35694 2894 35746
rect 2894 35694 2946 35746
rect 2946 35694 2948 35746
rect 2892 35692 2948 35694
rect 3052 35746 3108 35748
rect 3052 35694 3054 35746
rect 3054 35694 3106 35746
rect 3106 35694 3108 35746
rect 3052 35692 3108 35694
rect 3212 35746 3268 35748
rect 3212 35694 3214 35746
rect 3214 35694 3266 35746
rect 3266 35694 3268 35746
rect 3212 35692 3268 35694
rect 3372 35746 3428 35748
rect 3372 35694 3374 35746
rect 3374 35694 3426 35746
rect 3426 35694 3428 35746
rect 3372 35692 3428 35694
rect 3532 35746 3588 35748
rect 3532 35694 3534 35746
rect 3534 35694 3586 35746
rect 3586 35694 3588 35746
rect 3532 35692 3588 35694
rect 3692 35746 3748 35748
rect 3692 35694 3694 35746
rect 3694 35694 3746 35746
rect 3746 35694 3748 35746
rect 3692 35692 3748 35694
rect 3852 35746 3908 35748
rect 3852 35694 3854 35746
rect 3854 35694 3906 35746
rect 3906 35694 3908 35746
rect 3852 35692 3908 35694
rect 4012 35746 4068 35748
rect 4012 35694 4014 35746
rect 4014 35694 4066 35746
rect 4066 35694 4068 35746
rect 4012 35692 4068 35694
rect 4172 35746 4228 35748
rect 4172 35694 4174 35746
rect 4174 35694 4226 35746
rect 4226 35694 4228 35746
rect 4172 35692 4228 35694
rect 4332 35746 4388 35748
rect 4332 35694 4334 35746
rect 4334 35694 4386 35746
rect 4386 35694 4388 35746
rect 4332 35692 4388 35694
rect 4492 35746 4548 35748
rect 4492 35694 4494 35746
rect 4494 35694 4546 35746
rect 4546 35694 4548 35746
rect 4492 35692 4548 35694
rect 4652 35746 4708 35748
rect 4652 35694 4654 35746
rect 4654 35694 4706 35746
rect 4706 35694 4708 35746
rect 4652 35692 4708 35694
rect 4812 35746 4868 35748
rect 4812 35694 4814 35746
rect 4814 35694 4866 35746
rect 4866 35694 4868 35746
rect 4812 35692 4868 35694
rect 4972 35746 5028 35748
rect 4972 35694 4974 35746
rect 4974 35694 5026 35746
rect 5026 35694 5028 35746
rect 4972 35692 5028 35694
rect 5132 35746 5188 35748
rect 5132 35694 5134 35746
rect 5134 35694 5186 35746
rect 5186 35694 5188 35746
rect 5132 35692 5188 35694
rect 5292 35746 5348 35748
rect 5292 35694 5294 35746
rect 5294 35694 5346 35746
rect 5346 35694 5348 35746
rect 5292 35692 5348 35694
rect 5452 35746 5508 35748
rect 5452 35694 5454 35746
rect 5454 35694 5506 35746
rect 5506 35694 5508 35746
rect 5452 35692 5508 35694
rect 5612 35746 5668 35748
rect 5612 35694 5614 35746
rect 5614 35694 5666 35746
rect 5666 35694 5668 35746
rect 5612 35692 5668 35694
rect 5772 35746 5828 35748
rect 5772 35694 5774 35746
rect 5774 35694 5826 35746
rect 5826 35694 5828 35746
rect 5772 35692 5828 35694
rect 5932 35746 5988 35748
rect 5932 35694 5934 35746
rect 5934 35694 5986 35746
rect 5986 35694 5988 35746
rect 5932 35692 5988 35694
rect 6092 35746 6148 35748
rect 6092 35694 6094 35746
rect 6094 35694 6146 35746
rect 6146 35694 6148 35746
rect 6092 35692 6148 35694
rect 6252 35746 6308 35748
rect 6252 35694 6254 35746
rect 6254 35694 6306 35746
rect 6306 35694 6308 35746
rect 6252 35692 6308 35694
rect 6412 35746 6468 35748
rect 6412 35694 6414 35746
rect 6414 35694 6466 35746
rect 6466 35694 6468 35746
rect 6412 35692 6468 35694
rect 6572 35746 6628 35748
rect 6572 35694 6574 35746
rect 6574 35694 6626 35746
rect 6626 35694 6628 35746
rect 6572 35692 6628 35694
rect 6732 35746 6788 35748
rect 6732 35694 6734 35746
rect 6734 35694 6786 35746
rect 6786 35694 6788 35746
rect 6732 35692 6788 35694
rect 6892 35746 6948 35748
rect 6892 35694 6894 35746
rect 6894 35694 6946 35746
rect 6946 35694 6948 35746
rect 6892 35692 6948 35694
rect 7052 35746 7108 35748
rect 7052 35694 7054 35746
rect 7054 35694 7106 35746
rect 7106 35694 7108 35746
rect 7052 35692 7108 35694
rect 7212 35746 7268 35748
rect 7212 35694 7214 35746
rect 7214 35694 7266 35746
rect 7266 35694 7268 35746
rect 7212 35692 7268 35694
rect 7372 35746 7428 35748
rect 7372 35694 7374 35746
rect 7374 35694 7426 35746
rect 7426 35694 7428 35746
rect 7372 35692 7428 35694
rect 7532 35746 7588 35748
rect 7532 35694 7534 35746
rect 7534 35694 7586 35746
rect 7586 35694 7588 35746
rect 7532 35692 7588 35694
rect 7692 35746 7748 35748
rect 7692 35694 7694 35746
rect 7694 35694 7746 35746
rect 7746 35694 7748 35746
rect 7692 35692 7748 35694
rect 7852 35746 7908 35748
rect 7852 35694 7854 35746
rect 7854 35694 7906 35746
rect 7906 35694 7908 35746
rect 7852 35692 7908 35694
rect 8012 35746 8068 35748
rect 8012 35694 8014 35746
rect 8014 35694 8066 35746
rect 8066 35694 8068 35746
rect 8012 35692 8068 35694
rect 8172 35746 8228 35748
rect 8172 35694 8174 35746
rect 8174 35694 8226 35746
rect 8226 35694 8228 35746
rect 8172 35692 8228 35694
rect 8332 35746 8388 35748
rect 8332 35694 8334 35746
rect 8334 35694 8386 35746
rect 8386 35694 8388 35746
rect 8332 35692 8388 35694
rect 9452 35692 9508 35748
rect 9772 35692 9828 35748
rect 10092 35692 10148 35748
rect 10412 35692 10468 35748
rect 10732 35692 10788 35748
rect 11052 35692 11108 35748
rect 11372 35692 11428 35748
rect 12492 35746 12548 35748
rect 12492 35694 12494 35746
rect 12494 35694 12546 35746
rect 12546 35694 12548 35746
rect 12492 35692 12548 35694
rect 12652 35746 12708 35748
rect 12652 35694 12654 35746
rect 12654 35694 12706 35746
rect 12706 35694 12708 35746
rect 12652 35692 12708 35694
rect 12812 35746 12868 35748
rect 12812 35694 12814 35746
rect 12814 35694 12866 35746
rect 12866 35694 12868 35746
rect 12812 35692 12868 35694
rect 12972 35746 13028 35748
rect 12972 35694 12974 35746
rect 12974 35694 13026 35746
rect 13026 35694 13028 35746
rect 12972 35692 13028 35694
rect 13132 35746 13188 35748
rect 13132 35694 13134 35746
rect 13134 35694 13186 35746
rect 13186 35694 13188 35746
rect 13132 35692 13188 35694
rect 13292 35746 13348 35748
rect 13292 35694 13294 35746
rect 13294 35694 13346 35746
rect 13346 35694 13348 35746
rect 13292 35692 13348 35694
rect 13452 35746 13508 35748
rect 13452 35694 13454 35746
rect 13454 35694 13506 35746
rect 13506 35694 13508 35746
rect 13452 35692 13508 35694
rect 13612 35746 13668 35748
rect 13612 35694 13614 35746
rect 13614 35694 13666 35746
rect 13666 35694 13668 35746
rect 13612 35692 13668 35694
rect 13772 35746 13828 35748
rect 13772 35694 13774 35746
rect 13774 35694 13826 35746
rect 13826 35694 13828 35746
rect 13772 35692 13828 35694
rect 13932 35746 13988 35748
rect 13932 35694 13934 35746
rect 13934 35694 13986 35746
rect 13986 35694 13988 35746
rect 13932 35692 13988 35694
rect 14092 35746 14148 35748
rect 14092 35694 14094 35746
rect 14094 35694 14146 35746
rect 14146 35694 14148 35746
rect 14092 35692 14148 35694
rect 14252 35746 14308 35748
rect 14252 35694 14254 35746
rect 14254 35694 14306 35746
rect 14306 35694 14308 35746
rect 14252 35692 14308 35694
rect 14412 35746 14468 35748
rect 14412 35694 14414 35746
rect 14414 35694 14466 35746
rect 14466 35694 14468 35746
rect 14412 35692 14468 35694
rect 14572 35746 14628 35748
rect 14572 35694 14574 35746
rect 14574 35694 14626 35746
rect 14626 35694 14628 35746
rect 14572 35692 14628 35694
rect 14732 35746 14788 35748
rect 14732 35694 14734 35746
rect 14734 35694 14786 35746
rect 14786 35694 14788 35746
rect 14732 35692 14788 35694
rect 14892 35746 14948 35748
rect 14892 35694 14894 35746
rect 14894 35694 14946 35746
rect 14946 35694 14948 35746
rect 14892 35692 14948 35694
rect 15052 35746 15108 35748
rect 15052 35694 15054 35746
rect 15054 35694 15106 35746
rect 15106 35694 15108 35746
rect 15052 35692 15108 35694
rect 15212 35746 15268 35748
rect 15212 35694 15214 35746
rect 15214 35694 15266 35746
rect 15266 35694 15268 35746
rect 15212 35692 15268 35694
rect 15372 35746 15428 35748
rect 15372 35694 15374 35746
rect 15374 35694 15426 35746
rect 15426 35694 15428 35746
rect 15372 35692 15428 35694
rect 15532 35746 15588 35748
rect 15532 35694 15534 35746
rect 15534 35694 15586 35746
rect 15586 35694 15588 35746
rect 15532 35692 15588 35694
rect 15692 35746 15748 35748
rect 15692 35694 15694 35746
rect 15694 35694 15746 35746
rect 15746 35694 15748 35746
rect 15692 35692 15748 35694
rect 15852 35746 15908 35748
rect 15852 35694 15854 35746
rect 15854 35694 15906 35746
rect 15906 35694 15908 35746
rect 15852 35692 15908 35694
rect 16012 35746 16068 35748
rect 16012 35694 16014 35746
rect 16014 35694 16066 35746
rect 16066 35694 16068 35746
rect 16012 35692 16068 35694
rect 16172 35746 16228 35748
rect 16172 35694 16174 35746
rect 16174 35694 16226 35746
rect 16226 35694 16228 35746
rect 16172 35692 16228 35694
rect 16332 35746 16388 35748
rect 16332 35694 16334 35746
rect 16334 35694 16386 35746
rect 16386 35694 16388 35746
rect 16332 35692 16388 35694
rect 16492 35746 16548 35748
rect 16492 35694 16494 35746
rect 16494 35694 16546 35746
rect 16546 35694 16548 35746
rect 16492 35692 16548 35694
rect 16652 35746 16708 35748
rect 16652 35694 16654 35746
rect 16654 35694 16706 35746
rect 16706 35694 16708 35746
rect 16652 35692 16708 35694
rect 16812 35746 16868 35748
rect 16812 35694 16814 35746
rect 16814 35694 16866 35746
rect 16866 35694 16868 35746
rect 16812 35692 16868 35694
rect 16972 35746 17028 35748
rect 16972 35694 16974 35746
rect 16974 35694 17026 35746
rect 17026 35694 17028 35746
rect 16972 35692 17028 35694
rect 17132 35746 17188 35748
rect 17132 35694 17134 35746
rect 17134 35694 17186 35746
rect 17186 35694 17188 35746
rect 17132 35692 17188 35694
rect 17292 35746 17348 35748
rect 17292 35694 17294 35746
rect 17294 35694 17346 35746
rect 17346 35694 17348 35746
rect 17292 35692 17348 35694
rect 17452 35746 17508 35748
rect 17452 35694 17454 35746
rect 17454 35694 17506 35746
rect 17506 35694 17508 35746
rect 17452 35692 17508 35694
rect 17612 35746 17668 35748
rect 17612 35694 17614 35746
rect 17614 35694 17666 35746
rect 17666 35694 17668 35746
rect 17612 35692 17668 35694
rect 17772 35746 17828 35748
rect 17772 35694 17774 35746
rect 17774 35694 17826 35746
rect 17826 35694 17828 35746
rect 17772 35692 17828 35694
rect 17932 35746 17988 35748
rect 17932 35694 17934 35746
rect 17934 35694 17986 35746
rect 17986 35694 17988 35746
rect 17932 35692 17988 35694
rect 18092 35746 18148 35748
rect 18092 35694 18094 35746
rect 18094 35694 18146 35746
rect 18146 35694 18148 35746
rect 18092 35692 18148 35694
rect 18252 35746 18308 35748
rect 18252 35694 18254 35746
rect 18254 35694 18306 35746
rect 18306 35694 18308 35746
rect 18252 35692 18308 35694
rect 18412 35746 18468 35748
rect 18412 35694 18414 35746
rect 18414 35694 18466 35746
rect 18466 35694 18468 35746
rect 18412 35692 18468 35694
rect 18572 35746 18628 35748
rect 18572 35694 18574 35746
rect 18574 35694 18626 35746
rect 18626 35694 18628 35746
rect 18572 35692 18628 35694
rect 18732 35746 18788 35748
rect 18732 35694 18734 35746
rect 18734 35694 18786 35746
rect 18786 35694 18788 35746
rect 18732 35692 18788 35694
rect 18892 35746 18948 35748
rect 18892 35694 18894 35746
rect 18894 35694 18946 35746
rect 18946 35694 18948 35746
rect 18892 35692 18948 35694
rect 20012 35692 20068 35748
rect 20332 35692 20388 35748
rect 20652 35692 20708 35748
rect 20972 35692 21028 35748
rect 21292 35692 21348 35748
rect 21612 35692 21668 35748
rect 21932 35692 21988 35748
rect 23132 35746 23188 35748
rect 23132 35694 23134 35746
rect 23134 35694 23186 35746
rect 23186 35694 23188 35746
rect 23132 35692 23188 35694
rect 23292 35746 23348 35748
rect 23292 35694 23294 35746
rect 23294 35694 23346 35746
rect 23346 35694 23348 35746
rect 23292 35692 23348 35694
rect 23452 35746 23508 35748
rect 23452 35694 23454 35746
rect 23454 35694 23506 35746
rect 23506 35694 23508 35746
rect 23452 35692 23508 35694
rect 23612 35746 23668 35748
rect 23612 35694 23614 35746
rect 23614 35694 23666 35746
rect 23666 35694 23668 35746
rect 23612 35692 23668 35694
rect 23772 35746 23828 35748
rect 23772 35694 23774 35746
rect 23774 35694 23826 35746
rect 23826 35694 23828 35746
rect 23772 35692 23828 35694
rect 23932 35746 23988 35748
rect 23932 35694 23934 35746
rect 23934 35694 23986 35746
rect 23986 35694 23988 35746
rect 23932 35692 23988 35694
rect 24092 35746 24148 35748
rect 24092 35694 24094 35746
rect 24094 35694 24146 35746
rect 24146 35694 24148 35746
rect 24092 35692 24148 35694
rect 24252 35746 24308 35748
rect 24252 35694 24254 35746
rect 24254 35694 24306 35746
rect 24306 35694 24308 35746
rect 24252 35692 24308 35694
rect 24412 35746 24468 35748
rect 24412 35694 24414 35746
rect 24414 35694 24466 35746
rect 24466 35694 24468 35746
rect 24412 35692 24468 35694
rect 24572 35746 24628 35748
rect 24572 35694 24574 35746
rect 24574 35694 24626 35746
rect 24626 35694 24628 35746
rect 24572 35692 24628 35694
rect 24732 35746 24788 35748
rect 24732 35694 24734 35746
rect 24734 35694 24786 35746
rect 24786 35694 24788 35746
rect 24732 35692 24788 35694
rect 24892 35746 24948 35748
rect 24892 35694 24894 35746
rect 24894 35694 24946 35746
rect 24946 35694 24948 35746
rect 24892 35692 24948 35694
rect 25052 35746 25108 35748
rect 25052 35694 25054 35746
rect 25054 35694 25106 35746
rect 25106 35694 25108 35746
rect 25052 35692 25108 35694
rect 25212 35746 25268 35748
rect 25212 35694 25214 35746
rect 25214 35694 25266 35746
rect 25266 35694 25268 35746
rect 25212 35692 25268 35694
rect 25372 35746 25428 35748
rect 25372 35694 25374 35746
rect 25374 35694 25426 35746
rect 25426 35694 25428 35746
rect 25372 35692 25428 35694
rect 25532 35746 25588 35748
rect 25532 35694 25534 35746
rect 25534 35694 25586 35746
rect 25586 35694 25588 35746
rect 25532 35692 25588 35694
rect 25692 35746 25748 35748
rect 25692 35694 25694 35746
rect 25694 35694 25746 35746
rect 25746 35694 25748 35746
rect 25692 35692 25748 35694
rect 25852 35746 25908 35748
rect 25852 35694 25854 35746
rect 25854 35694 25906 35746
rect 25906 35694 25908 35746
rect 25852 35692 25908 35694
rect 26012 35746 26068 35748
rect 26012 35694 26014 35746
rect 26014 35694 26066 35746
rect 26066 35694 26068 35746
rect 26012 35692 26068 35694
rect 26172 35746 26228 35748
rect 26172 35694 26174 35746
rect 26174 35694 26226 35746
rect 26226 35694 26228 35746
rect 26172 35692 26228 35694
rect 26332 35746 26388 35748
rect 26332 35694 26334 35746
rect 26334 35694 26386 35746
rect 26386 35694 26388 35746
rect 26332 35692 26388 35694
rect 26492 35746 26548 35748
rect 26492 35694 26494 35746
rect 26494 35694 26546 35746
rect 26546 35694 26548 35746
rect 26492 35692 26548 35694
rect 26652 35746 26708 35748
rect 26652 35694 26654 35746
rect 26654 35694 26706 35746
rect 26706 35694 26708 35746
rect 26652 35692 26708 35694
rect 26812 35746 26868 35748
rect 26812 35694 26814 35746
rect 26814 35694 26866 35746
rect 26866 35694 26868 35746
rect 26812 35692 26868 35694
rect 26972 35746 27028 35748
rect 26972 35694 26974 35746
rect 26974 35694 27026 35746
rect 27026 35694 27028 35746
rect 26972 35692 27028 35694
rect 27132 35746 27188 35748
rect 27132 35694 27134 35746
rect 27134 35694 27186 35746
rect 27186 35694 27188 35746
rect 27132 35692 27188 35694
rect 27292 35746 27348 35748
rect 27292 35694 27294 35746
rect 27294 35694 27346 35746
rect 27346 35694 27348 35746
rect 27292 35692 27348 35694
rect 27452 35746 27508 35748
rect 27452 35694 27454 35746
rect 27454 35694 27506 35746
rect 27506 35694 27508 35746
rect 27452 35692 27508 35694
rect 27612 35746 27668 35748
rect 27612 35694 27614 35746
rect 27614 35694 27666 35746
rect 27666 35694 27668 35746
rect 27612 35692 27668 35694
rect 27772 35746 27828 35748
rect 27772 35694 27774 35746
rect 27774 35694 27826 35746
rect 27826 35694 27828 35746
rect 27772 35692 27828 35694
rect 27932 35746 27988 35748
rect 27932 35694 27934 35746
rect 27934 35694 27986 35746
rect 27986 35694 27988 35746
rect 27932 35692 27988 35694
rect 28092 35746 28148 35748
rect 28092 35694 28094 35746
rect 28094 35694 28146 35746
rect 28146 35694 28148 35746
rect 28092 35692 28148 35694
rect 28252 35746 28308 35748
rect 28252 35694 28254 35746
rect 28254 35694 28306 35746
rect 28306 35694 28308 35746
rect 28252 35692 28308 35694
rect 28412 35746 28468 35748
rect 28412 35694 28414 35746
rect 28414 35694 28466 35746
rect 28466 35694 28468 35746
rect 28412 35692 28468 35694
rect 28572 35746 28628 35748
rect 28572 35694 28574 35746
rect 28574 35694 28626 35746
rect 28626 35694 28628 35746
rect 28572 35692 28628 35694
rect 28732 35746 28788 35748
rect 28732 35694 28734 35746
rect 28734 35694 28786 35746
rect 28786 35694 28788 35746
rect 28732 35692 28788 35694
rect 28892 35746 28948 35748
rect 28892 35694 28894 35746
rect 28894 35694 28946 35746
rect 28946 35694 28948 35746
rect 28892 35692 28948 35694
rect 29052 35746 29108 35748
rect 29052 35694 29054 35746
rect 29054 35694 29106 35746
rect 29106 35694 29108 35746
rect 29052 35692 29108 35694
rect 29212 35746 29268 35748
rect 29212 35694 29214 35746
rect 29214 35694 29266 35746
rect 29266 35694 29268 35746
rect 29212 35692 29268 35694
rect 29372 35746 29428 35748
rect 29372 35694 29374 35746
rect 29374 35694 29426 35746
rect 29426 35694 29428 35746
rect 29372 35692 29428 35694
rect 30492 35692 30548 35748
rect 30812 35692 30868 35748
rect 31132 35692 31188 35748
rect 31452 35692 31508 35748
rect 31772 35692 31828 35748
rect 32092 35692 32148 35748
rect 32412 35692 32468 35748
rect 33532 35746 33588 35748
rect 33532 35694 33534 35746
rect 33534 35694 33586 35746
rect 33586 35694 33588 35746
rect 33532 35692 33588 35694
rect 33692 35746 33748 35748
rect 33692 35694 33694 35746
rect 33694 35694 33746 35746
rect 33746 35694 33748 35746
rect 33692 35692 33748 35694
rect 33852 35746 33908 35748
rect 33852 35694 33854 35746
rect 33854 35694 33906 35746
rect 33906 35694 33908 35746
rect 33852 35692 33908 35694
rect 34012 35746 34068 35748
rect 34012 35694 34014 35746
rect 34014 35694 34066 35746
rect 34066 35694 34068 35746
rect 34012 35692 34068 35694
rect 34172 35746 34228 35748
rect 34172 35694 34174 35746
rect 34174 35694 34226 35746
rect 34226 35694 34228 35746
rect 34172 35692 34228 35694
rect 34332 35746 34388 35748
rect 34332 35694 34334 35746
rect 34334 35694 34386 35746
rect 34386 35694 34388 35746
rect 34332 35692 34388 35694
rect 34492 35746 34548 35748
rect 34492 35694 34494 35746
rect 34494 35694 34546 35746
rect 34546 35694 34548 35746
rect 34492 35692 34548 35694
rect 34652 35746 34708 35748
rect 34652 35694 34654 35746
rect 34654 35694 34706 35746
rect 34706 35694 34708 35746
rect 34652 35692 34708 35694
rect 34812 35746 34868 35748
rect 34812 35694 34814 35746
rect 34814 35694 34866 35746
rect 34866 35694 34868 35746
rect 34812 35692 34868 35694
rect 34972 35746 35028 35748
rect 34972 35694 34974 35746
rect 34974 35694 35026 35746
rect 35026 35694 35028 35746
rect 34972 35692 35028 35694
rect 35132 35746 35188 35748
rect 35132 35694 35134 35746
rect 35134 35694 35186 35746
rect 35186 35694 35188 35746
rect 35132 35692 35188 35694
rect 35292 35746 35348 35748
rect 35292 35694 35294 35746
rect 35294 35694 35346 35746
rect 35346 35694 35348 35746
rect 35292 35692 35348 35694
rect 35452 35746 35508 35748
rect 35452 35694 35454 35746
rect 35454 35694 35506 35746
rect 35506 35694 35508 35746
rect 35452 35692 35508 35694
rect 35612 35746 35668 35748
rect 35612 35694 35614 35746
rect 35614 35694 35666 35746
rect 35666 35694 35668 35746
rect 35612 35692 35668 35694
rect 35772 35746 35828 35748
rect 35772 35694 35774 35746
rect 35774 35694 35826 35746
rect 35826 35694 35828 35746
rect 35772 35692 35828 35694
rect 35932 35746 35988 35748
rect 35932 35694 35934 35746
rect 35934 35694 35986 35746
rect 35986 35694 35988 35746
rect 35932 35692 35988 35694
rect 36092 35746 36148 35748
rect 36092 35694 36094 35746
rect 36094 35694 36146 35746
rect 36146 35694 36148 35746
rect 36092 35692 36148 35694
rect 36252 35746 36308 35748
rect 36252 35694 36254 35746
rect 36254 35694 36306 35746
rect 36306 35694 36308 35746
rect 36252 35692 36308 35694
rect 36412 35746 36468 35748
rect 36412 35694 36414 35746
rect 36414 35694 36466 35746
rect 36466 35694 36468 35746
rect 36412 35692 36468 35694
rect 36572 35746 36628 35748
rect 36572 35694 36574 35746
rect 36574 35694 36626 35746
rect 36626 35694 36628 35746
rect 36572 35692 36628 35694
rect 36732 35746 36788 35748
rect 36732 35694 36734 35746
rect 36734 35694 36786 35746
rect 36786 35694 36788 35746
rect 36732 35692 36788 35694
rect 36892 35746 36948 35748
rect 36892 35694 36894 35746
rect 36894 35694 36946 35746
rect 36946 35694 36948 35746
rect 36892 35692 36948 35694
rect 37052 35746 37108 35748
rect 37052 35694 37054 35746
rect 37054 35694 37106 35746
rect 37106 35694 37108 35746
rect 37052 35692 37108 35694
rect 37212 35746 37268 35748
rect 37212 35694 37214 35746
rect 37214 35694 37266 35746
rect 37266 35694 37268 35746
rect 37212 35692 37268 35694
rect 37372 35746 37428 35748
rect 37372 35694 37374 35746
rect 37374 35694 37426 35746
rect 37426 35694 37428 35746
rect 37372 35692 37428 35694
rect 37532 35746 37588 35748
rect 37532 35694 37534 35746
rect 37534 35694 37586 35746
rect 37586 35694 37588 35746
rect 37532 35692 37588 35694
rect 37692 35746 37748 35748
rect 37692 35694 37694 35746
rect 37694 35694 37746 35746
rect 37746 35694 37748 35746
rect 37692 35692 37748 35694
rect 37852 35746 37908 35748
rect 37852 35694 37854 35746
rect 37854 35694 37906 35746
rect 37906 35694 37908 35746
rect 37852 35692 37908 35694
rect 38012 35746 38068 35748
rect 38012 35694 38014 35746
rect 38014 35694 38066 35746
rect 38066 35694 38068 35746
rect 38012 35692 38068 35694
rect 38172 35746 38228 35748
rect 38172 35694 38174 35746
rect 38174 35694 38226 35746
rect 38226 35694 38228 35746
rect 38172 35692 38228 35694
rect 38332 35746 38388 35748
rect 38332 35694 38334 35746
rect 38334 35694 38386 35746
rect 38386 35694 38388 35746
rect 38332 35692 38388 35694
rect 38492 35746 38548 35748
rect 38492 35694 38494 35746
rect 38494 35694 38546 35746
rect 38546 35694 38548 35746
rect 38492 35692 38548 35694
rect 38652 35746 38708 35748
rect 38652 35694 38654 35746
rect 38654 35694 38706 35746
rect 38706 35694 38708 35746
rect 38652 35692 38708 35694
rect 38812 35746 38868 35748
rect 38812 35694 38814 35746
rect 38814 35694 38866 35746
rect 38866 35694 38868 35746
rect 38812 35692 38868 35694
rect 38972 35746 39028 35748
rect 38972 35694 38974 35746
rect 38974 35694 39026 35746
rect 39026 35694 39028 35746
rect 38972 35692 39028 35694
rect 39132 35746 39188 35748
rect 39132 35694 39134 35746
rect 39134 35694 39186 35746
rect 39186 35694 39188 35746
rect 39132 35692 39188 35694
rect 39292 35746 39348 35748
rect 39292 35694 39294 35746
rect 39294 35694 39346 35746
rect 39346 35694 39348 35746
rect 39292 35692 39348 35694
rect 39452 35746 39508 35748
rect 39452 35694 39454 35746
rect 39454 35694 39506 35746
rect 39506 35694 39508 35746
rect 39452 35692 39508 35694
rect 39612 35746 39668 35748
rect 39612 35694 39614 35746
rect 39614 35694 39666 35746
rect 39666 35694 39668 35746
rect 39612 35692 39668 35694
rect 39772 35746 39828 35748
rect 39772 35694 39774 35746
rect 39774 35694 39826 35746
rect 39826 35694 39828 35746
rect 39772 35692 39828 35694
rect 39932 35746 39988 35748
rect 39932 35694 39934 35746
rect 39934 35694 39986 35746
rect 39986 35694 39988 35746
rect 39932 35692 39988 35694
rect 40092 35746 40148 35748
rect 40092 35694 40094 35746
rect 40094 35694 40146 35746
rect 40146 35694 40148 35746
rect 40092 35692 40148 35694
rect 40252 35746 40308 35748
rect 40252 35694 40254 35746
rect 40254 35694 40306 35746
rect 40306 35694 40308 35746
rect 40252 35692 40308 35694
rect 40412 35746 40468 35748
rect 40412 35694 40414 35746
rect 40414 35694 40466 35746
rect 40466 35694 40468 35746
rect 40412 35692 40468 35694
rect 40572 35746 40628 35748
rect 40572 35694 40574 35746
rect 40574 35694 40626 35746
rect 40626 35694 40628 35746
rect 40572 35692 40628 35694
rect 40732 35746 40788 35748
rect 40732 35694 40734 35746
rect 40734 35694 40786 35746
rect 40786 35694 40788 35746
rect 40732 35692 40788 35694
rect 40892 35746 40948 35748
rect 40892 35694 40894 35746
rect 40894 35694 40946 35746
rect 40946 35694 40948 35746
rect 40892 35692 40948 35694
rect 41052 35746 41108 35748
rect 41052 35694 41054 35746
rect 41054 35694 41106 35746
rect 41106 35694 41108 35746
rect 41052 35692 41108 35694
rect 41212 35746 41268 35748
rect 41212 35694 41214 35746
rect 41214 35694 41266 35746
rect 41266 35694 41268 35746
rect 41212 35692 41268 35694
rect 41372 35746 41428 35748
rect 41372 35694 41374 35746
rect 41374 35694 41426 35746
rect 41426 35694 41428 35746
rect 41372 35692 41428 35694
rect 41532 35746 41588 35748
rect 41532 35694 41534 35746
rect 41534 35694 41586 35746
rect 41586 35694 41588 35746
rect 41532 35692 41588 35694
rect 41692 35746 41748 35748
rect 41692 35694 41694 35746
rect 41694 35694 41746 35746
rect 41746 35694 41748 35746
rect 41692 35692 41748 35694
rect 41852 35746 41908 35748
rect 41852 35694 41854 35746
rect 41854 35694 41906 35746
rect 41906 35694 41908 35746
rect 41852 35692 41908 35694
rect 10252 35532 10308 35588
rect 21132 35532 21188 35588
rect 31612 35532 31668 35588
rect 12 35426 68 35428
rect 12 35374 14 35426
rect 14 35374 66 35426
rect 66 35374 68 35426
rect 12 35372 68 35374
rect 172 35426 228 35428
rect 172 35374 174 35426
rect 174 35374 226 35426
rect 226 35374 228 35426
rect 172 35372 228 35374
rect 332 35426 388 35428
rect 332 35374 334 35426
rect 334 35374 386 35426
rect 386 35374 388 35426
rect 332 35372 388 35374
rect 492 35426 548 35428
rect 492 35374 494 35426
rect 494 35374 546 35426
rect 546 35374 548 35426
rect 492 35372 548 35374
rect 652 35426 708 35428
rect 652 35374 654 35426
rect 654 35374 706 35426
rect 706 35374 708 35426
rect 652 35372 708 35374
rect 812 35426 868 35428
rect 812 35374 814 35426
rect 814 35374 866 35426
rect 866 35374 868 35426
rect 812 35372 868 35374
rect 972 35426 1028 35428
rect 972 35374 974 35426
rect 974 35374 1026 35426
rect 1026 35374 1028 35426
rect 972 35372 1028 35374
rect 1132 35426 1188 35428
rect 1132 35374 1134 35426
rect 1134 35374 1186 35426
rect 1186 35374 1188 35426
rect 1132 35372 1188 35374
rect 1292 35426 1348 35428
rect 1292 35374 1294 35426
rect 1294 35374 1346 35426
rect 1346 35374 1348 35426
rect 1292 35372 1348 35374
rect 1452 35426 1508 35428
rect 1452 35374 1454 35426
rect 1454 35374 1506 35426
rect 1506 35374 1508 35426
rect 1452 35372 1508 35374
rect 1612 35426 1668 35428
rect 1612 35374 1614 35426
rect 1614 35374 1666 35426
rect 1666 35374 1668 35426
rect 1612 35372 1668 35374
rect 1772 35426 1828 35428
rect 1772 35374 1774 35426
rect 1774 35374 1826 35426
rect 1826 35374 1828 35426
rect 1772 35372 1828 35374
rect 1932 35426 1988 35428
rect 1932 35374 1934 35426
rect 1934 35374 1986 35426
rect 1986 35374 1988 35426
rect 1932 35372 1988 35374
rect 2092 35426 2148 35428
rect 2092 35374 2094 35426
rect 2094 35374 2146 35426
rect 2146 35374 2148 35426
rect 2092 35372 2148 35374
rect 2252 35426 2308 35428
rect 2252 35374 2254 35426
rect 2254 35374 2306 35426
rect 2306 35374 2308 35426
rect 2252 35372 2308 35374
rect 2412 35426 2468 35428
rect 2412 35374 2414 35426
rect 2414 35374 2466 35426
rect 2466 35374 2468 35426
rect 2412 35372 2468 35374
rect 2572 35426 2628 35428
rect 2572 35374 2574 35426
rect 2574 35374 2626 35426
rect 2626 35374 2628 35426
rect 2572 35372 2628 35374
rect 2732 35426 2788 35428
rect 2732 35374 2734 35426
rect 2734 35374 2786 35426
rect 2786 35374 2788 35426
rect 2732 35372 2788 35374
rect 2892 35426 2948 35428
rect 2892 35374 2894 35426
rect 2894 35374 2946 35426
rect 2946 35374 2948 35426
rect 2892 35372 2948 35374
rect 3052 35426 3108 35428
rect 3052 35374 3054 35426
rect 3054 35374 3106 35426
rect 3106 35374 3108 35426
rect 3052 35372 3108 35374
rect 3212 35426 3268 35428
rect 3212 35374 3214 35426
rect 3214 35374 3266 35426
rect 3266 35374 3268 35426
rect 3212 35372 3268 35374
rect 3372 35426 3428 35428
rect 3372 35374 3374 35426
rect 3374 35374 3426 35426
rect 3426 35374 3428 35426
rect 3372 35372 3428 35374
rect 3532 35426 3588 35428
rect 3532 35374 3534 35426
rect 3534 35374 3586 35426
rect 3586 35374 3588 35426
rect 3532 35372 3588 35374
rect 3692 35426 3748 35428
rect 3692 35374 3694 35426
rect 3694 35374 3746 35426
rect 3746 35374 3748 35426
rect 3692 35372 3748 35374
rect 3852 35426 3908 35428
rect 3852 35374 3854 35426
rect 3854 35374 3906 35426
rect 3906 35374 3908 35426
rect 3852 35372 3908 35374
rect 4012 35426 4068 35428
rect 4012 35374 4014 35426
rect 4014 35374 4066 35426
rect 4066 35374 4068 35426
rect 4012 35372 4068 35374
rect 4172 35426 4228 35428
rect 4172 35374 4174 35426
rect 4174 35374 4226 35426
rect 4226 35374 4228 35426
rect 4172 35372 4228 35374
rect 4332 35426 4388 35428
rect 4332 35374 4334 35426
rect 4334 35374 4386 35426
rect 4386 35374 4388 35426
rect 4332 35372 4388 35374
rect 4492 35426 4548 35428
rect 4492 35374 4494 35426
rect 4494 35374 4546 35426
rect 4546 35374 4548 35426
rect 4492 35372 4548 35374
rect 4652 35426 4708 35428
rect 4652 35374 4654 35426
rect 4654 35374 4706 35426
rect 4706 35374 4708 35426
rect 4652 35372 4708 35374
rect 4812 35426 4868 35428
rect 4812 35374 4814 35426
rect 4814 35374 4866 35426
rect 4866 35374 4868 35426
rect 4812 35372 4868 35374
rect 4972 35426 5028 35428
rect 4972 35374 4974 35426
rect 4974 35374 5026 35426
rect 5026 35374 5028 35426
rect 4972 35372 5028 35374
rect 5132 35426 5188 35428
rect 5132 35374 5134 35426
rect 5134 35374 5186 35426
rect 5186 35374 5188 35426
rect 5132 35372 5188 35374
rect 5292 35426 5348 35428
rect 5292 35374 5294 35426
rect 5294 35374 5346 35426
rect 5346 35374 5348 35426
rect 5292 35372 5348 35374
rect 5452 35426 5508 35428
rect 5452 35374 5454 35426
rect 5454 35374 5506 35426
rect 5506 35374 5508 35426
rect 5452 35372 5508 35374
rect 5612 35426 5668 35428
rect 5612 35374 5614 35426
rect 5614 35374 5666 35426
rect 5666 35374 5668 35426
rect 5612 35372 5668 35374
rect 5772 35426 5828 35428
rect 5772 35374 5774 35426
rect 5774 35374 5826 35426
rect 5826 35374 5828 35426
rect 5772 35372 5828 35374
rect 5932 35426 5988 35428
rect 5932 35374 5934 35426
rect 5934 35374 5986 35426
rect 5986 35374 5988 35426
rect 5932 35372 5988 35374
rect 6092 35426 6148 35428
rect 6092 35374 6094 35426
rect 6094 35374 6146 35426
rect 6146 35374 6148 35426
rect 6092 35372 6148 35374
rect 6252 35426 6308 35428
rect 6252 35374 6254 35426
rect 6254 35374 6306 35426
rect 6306 35374 6308 35426
rect 6252 35372 6308 35374
rect 6412 35426 6468 35428
rect 6412 35374 6414 35426
rect 6414 35374 6466 35426
rect 6466 35374 6468 35426
rect 6412 35372 6468 35374
rect 6572 35426 6628 35428
rect 6572 35374 6574 35426
rect 6574 35374 6626 35426
rect 6626 35374 6628 35426
rect 6572 35372 6628 35374
rect 6732 35426 6788 35428
rect 6732 35374 6734 35426
rect 6734 35374 6786 35426
rect 6786 35374 6788 35426
rect 6732 35372 6788 35374
rect 6892 35426 6948 35428
rect 6892 35374 6894 35426
rect 6894 35374 6946 35426
rect 6946 35374 6948 35426
rect 6892 35372 6948 35374
rect 7052 35426 7108 35428
rect 7052 35374 7054 35426
rect 7054 35374 7106 35426
rect 7106 35374 7108 35426
rect 7052 35372 7108 35374
rect 7212 35426 7268 35428
rect 7212 35374 7214 35426
rect 7214 35374 7266 35426
rect 7266 35374 7268 35426
rect 7212 35372 7268 35374
rect 7372 35426 7428 35428
rect 7372 35374 7374 35426
rect 7374 35374 7426 35426
rect 7426 35374 7428 35426
rect 7372 35372 7428 35374
rect 7532 35426 7588 35428
rect 7532 35374 7534 35426
rect 7534 35374 7586 35426
rect 7586 35374 7588 35426
rect 7532 35372 7588 35374
rect 7692 35426 7748 35428
rect 7692 35374 7694 35426
rect 7694 35374 7746 35426
rect 7746 35374 7748 35426
rect 7692 35372 7748 35374
rect 7852 35426 7908 35428
rect 7852 35374 7854 35426
rect 7854 35374 7906 35426
rect 7906 35374 7908 35426
rect 7852 35372 7908 35374
rect 8012 35426 8068 35428
rect 8012 35374 8014 35426
rect 8014 35374 8066 35426
rect 8066 35374 8068 35426
rect 8012 35372 8068 35374
rect 8172 35426 8228 35428
rect 8172 35374 8174 35426
rect 8174 35374 8226 35426
rect 8226 35374 8228 35426
rect 8172 35372 8228 35374
rect 8332 35426 8388 35428
rect 8332 35374 8334 35426
rect 8334 35374 8386 35426
rect 8386 35374 8388 35426
rect 8332 35372 8388 35374
rect 9452 35372 9508 35428
rect 9772 35372 9828 35428
rect 10092 35372 10148 35428
rect 10412 35372 10468 35428
rect 10732 35372 10788 35428
rect 11052 35372 11108 35428
rect 11372 35372 11428 35428
rect 12492 35426 12548 35428
rect 12492 35374 12494 35426
rect 12494 35374 12546 35426
rect 12546 35374 12548 35426
rect 12492 35372 12548 35374
rect 12652 35426 12708 35428
rect 12652 35374 12654 35426
rect 12654 35374 12706 35426
rect 12706 35374 12708 35426
rect 12652 35372 12708 35374
rect 12812 35426 12868 35428
rect 12812 35374 12814 35426
rect 12814 35374 12866 35426
rect 12866 35374 12868 35426
rect 12812 35372 12868 35374
rect 12972 35426 13028 35428
rect 12972 35374 12974 35426
rect 12974 35374 13026 35426
rect 13026 35374 13028 35426
rect 12972 35372 13028 35374
rect 13132 35426 13188 35428
rect 13132 35374 13134 35426
rect 13134 35374 13186 35426
rect 13186 35374 13188 35426
rect 13132 35372 13188 35374
rect 13292 35426 13348 35428
rect 13292 35374 13294 35426
rect 13294 35374 13346 35426
rect 13346 35374 13348 35426
rect 13292 35372 13348 35374
rect 13452 35426 13508 35428
rect 13452 35374 13454 35426
rect 13454 35374 13506 35426
rect 13506 35374 13508 35426
rect 13452 35372 13508 35374
rect 13612 35426 13668 35428
rect 13612 35374 13614 35426
rect 13614 35374 13666 35426
rect 13666 35374 13668 35426
rect 13612 35372 13668 35374
rect 13772 35426 13828 35428
rect 13772 35374 13774 35426
rect 13774 35374 13826 35426
rect 13826 35374 13828 35426
rect 13772 35372 13828 35374
rect 13932 35426 13988 35428
rect 13932 35374 13934 35426
rect 13934 35374 13986 35426
rect 13986 35374 13988 35426
rect 13932 35372 13988 35374
rect 14092 35426 14148 35428
rect 14092 35374 14094 35426
rect 14094 35374 14146 35426
rect 14146 35374 14148 35426
rect 14092 35372 14148 35374
rect 14252 35426 14308 35428
rect 14252 35374 14254 35426
rect 14254 35374 14306 35426
rect 14306 35374 14308 35426
rect 14252 35372 14308 35374
rect 14412 35426 14468 35428
rect 14412 35374 14414 35426
rect 14414 35374 14466 35426
rect 14466 35374 14468 35426
rect 14412 35372 14468 35374
rect 14572 35426 14628 35428
rect 14572 35374 14574 35426
rect 14574 35374 14626 35426
rect 14626 35374 14628 35426
rect 14572 35372 14628 35374
rect 14732 35426 14788 35428
rect 14732 35374 14734 35426
rect 14734 35374 14786 35426
rect 14786 35374 14788 35426
rect 14732 35372 14788 35374
rect 14892 35426 14948 35428
rect 14892 35374 14894 35426
rect 14894 35374 14946 35426
rect 14946 35374 14948 35426
rect 14892 35372 14948 35374
rect 15052 35426 15108 35428
rect 15052 35374 15054 35426
rect 15054 35374 15106 35426
rect 15106 35374 15108 35426
rect 15052 35372 15108 35374
rect 15212 35426 15268 35428
rect 15212 35374 15214 35426
rect 15214 35374 15266 35426
rect 15266 35374 15268 35426
rect 15212 35372 15268 35374
rect 15372 35426 15428 35428
rect 15372 35374 15374 35426
rect 15374 35374 15426 35426
rect 15426 35374 15428 35426
rect 15372 35372 15428 35374
rect 15532 35426 15588 35428
rect 15532 35374 15534 35426
rect 15534 35374 15586 35426
rect 15586 35374 15588 35426
rect 15532 35372 15588 35374
rect 15692 35426 15748 35428
rect 15692 35374 15694 35426
rect 15694 35374 15746 35426
rect 15746 35374 15748 35426
rect 15692 35372 15748 35374
rect 15852 35426 15908 35428
rect 15852 35374 15854 35426
rect 15854 35374 15906 35426
rect 15906 35374 15908 35426
rect 15852 35372 15908 35374
rect 16012 35426 16068 35428
rect 16012 35374 16014 35426
rect 16014 35374 16066 35426
rect 16066 35374 16068 35426
rect 16012 35372 16068 35374
rect 16172 35426 16228 35428
rect 16172 35374 16174 35426
rect 16174 35374 16226 35426
rect 16226 35374 16228 35426
rect 16172 35372 16228 35374
rect 16332 35426 16388 35428
rect 16332 35374 16334 35426
rect 16334 35374 16386 35426
rect 16386 35374 16388 35426
rect 16332 35372 16388 35374
rect 16492 35426 16548 35428
rect 16492 35374 16494 35426
rect 16494 35374 16546 35426
rect 16546 35374 16548 35426
rect 16492 35372 16548 35374
rect 16652 35426 16708 35428
rect 16652 35374 16654 35426
rect 16654 35374 16706 35426
rect 16706 35374 16708 35426
rect 16652 35372 16708 35374
rect 16812 35426 16868 35428
rect 16812 35374 16814 35426
rect 16814 35374 16866 35426
rect 16866 35374 16868 35426
rect 16812 35372 16868 35374
rect 16972 35426 17028 35428
rect 16972 35374 16974 35426
rect 16974 35374 17026 35426
rect 17026 35374 17028 35426
rect 16972 35372 17028 35374
rect 17132 35426 17188 35428
rect 17132 35374 17134 35426
rect 17134 35374 17186 35426
rect 17186 35374 17188 35426
rect 17132 35372 17188 35374
rect 17292 35426 17348 35428
rect 17292 35374 17294 35426
rect 17294 35374 17346 35426
rect 17346 35374 17348 35426
rect 17292 35372 17348 35374
rect 17452 35426 17508 35428
rect 17452 35374 17454 35426
rect 17454 35374 17506 35426
rect 17506 35374 17508 35426
rect 17452 35372 17508 35374
rect 17612 35426 17668 35428
rect 17612 35374 17614 35426
rect 17614 35374 17666 35426
rect 17666 35374 17668 35426
rect 17612 35372 17668 35374
rect 17772 35426 17828 35428
rect 17772 35374 17774 35426
rect 17774 35374 17826 35426
rect 17826 35374 17828 35426
rect 17772 35372 17828 35374
rect 17932 35426 17988 35428
rect 17932 35374 17934 35426
rect 17934 35374 17986 35426
rect 17986 35374 17988 35426
rect 17932 35372 17988 35374
rect 18092 35426 18148 35428
rect 18092 35374 18094 35426
rect 18094 35374 18146 35426
rect 18146 35374 18148 35426
rect 18092 35372 18148 35374
rect 18252 35426 18308 35428
rect 18252 35374 18254 35426
rect 18254 35374 18306 35426
rect 18306 35374 18308 35426
rect 18252 35372 18308 35374
rect 18412 35426 18468 35428
rect 18412 35374 18414 35426
rect 18414 35374 18466 35426
rect 18466 35374 18468 35426
rect 18412 35372 18468 35374
rect 18572 35426 18628 35428
rect 18572 35374 18574 35426
rect 18574 35374 18626 35426
rect 18626 35374 18628 35426
rect 18572 35372 18628 35374
rect 18732 35426 18788 35428
rect 18732 35374 18734 35426
rect 18734 35374 18786 35426
rect 18786 35374 18788 35426
rect 18732 35372 18788 35374
rect 18892 35426 18948 35428
rect 18892 35374 18894 35426
rect 18894 35374 18946 35426
rect 18946 35374 18948 35426
rect 18892 35372 18948 35374
rect 20012 35372 20068 35428
rect 20332 35372 20388 35428
rect 20652 35372 20708 35428
rect 20972 35372 21028 35428
rect 21292 35372 21348 35428
rect 21612 35372 21668 35428
rect 21932 35372 21988 35428
rect 23132 35426 23188 35428
rect 23132 35374 23134 35426
rect 23134 35374 23186 35426
rect 23186 35374 23188 35426
rect 23132 35372 23188 35374
rect 23292 35426 23348 35428
rect 23292 35374 23294 35426
rect 23294 35374 23346 35426
rect 23346 35374 23348 35426
rect 23292 35372 23348 35374
rect 23452 35426 23508 35428
rect 23452 35374 23454 35426
rect 23454 35374 23506 35426
rect 23506 35374 23508 35426
rect 23452 35372 23508 35374
rect 23612 35426 23668 35428
rect 23612 35374 23614 35426
rect 23614 35374 23666 35426
rect 23666 35374 23668 35426
rect 23612 35372 23668 35374
rect 23772 35426 23828 35428
rect 23772 35374 23774 35426
rect 23774 35374 23826 35426
rect 23826 35374 23828 35426
rect 23772 35372 23828 35374
rect 23932 35426 23988 35428
rect 23932 35374 23934 35426
rect 23934 35374 23986 35426
rect 23986 35374 23988 35426
rect 23932 35372 23988 35374
rect 24092 35426 24148 35428
rect 24092 35374 24094 35426
rect 24094 35374 24146 35426
rect 24146 35374 24148 35426
rect 24092 35372 24148 35374
rect 24252 35426 24308 35428
rect 24252 35374 24254 35426
rect 24254 35374 24306 35426
rect 24306 35374 24308 35426
rect 24252 35372 24308 35374
rect 24412 35426 24468 35428
rect 24412 35374 24414 35426
rect 24414 35374 24466 35426
rect 24466 35374 24468 35426
rect 24412 35372 24468 35374
rect 24572 35426 24628 35428
rect 24572 35374 24574 35426
rect 24574 35374 24626 35426
rect 24626 35374 24628 35426
rect 24572 35372 24628 35374
rect 24732 35426 24788 35428
rect 24732 35374 24734 35426
rect 24734 35374 24786 35426
rect 24786 35374 24788 35426
rect 24732 35372 24788 35374
rect 24892 35426 24948 35428
rect 24892 35374 24894 35426
rect 24894 35374 24946 35426
rect 24946 35374 24948 35426
rect 24892 35372 24948 35374
rect 25052 35426 25108 35428
rect 25052 35374 25054 35426
rect 25054 35374 25106 35426
rect 25106 35374 25108 35426
rect 25052 35372 25108 35374
rect 25212 35426 25268 35428
rect 25212 35374 25214 35426
rect 25214 35374 25266 35426
rect 25266 35374 25268 35426
rect 25212 35372 25268 35374
rect 25372 35426 25428 35428
rect 25372 35374 25374 35426
rect 25374 35374 25426 35426
rect 25426 35374 25428 35426
rect 25372 35372 25428 35374
rect 25532 35426 25588 35428
rect 25532 35374 25534 35426
rect 25534 35374 25586 35426
rect 25586 35374 25588 35426
rect 25532 35372 25588 35374
rect 25692 35426 25748 35428
rect 25692 35374 25694 35426
rect 25694 35374 25746 35426
rect 25746 35374 25748 35426
rect 25692 35372 25748 35374
rect 25852 35426 25908 35428
rect 25852 35374 25854 35426
rect 25854 35374 25906 35426
rect 25906 35374 25908 35426
rect 25852 35372 25908 35374
rect 26012 35426 26068 35428
rect 26012 35374 26014 35426
rect 26014 35374 26066 35426
rect 26066 35374 26068 35426
rect 26012 35372 26068 35374
rect 26172 35426 26228 35428
rect 26172 35374 26174 35426
rect 26174 35374 26226 35426
rect 26226 35374 26228 35426
rect 26172 35372 26228 35374
rect 26332 35426 26388 35428
rect 26332 35374 26334 35426
rect 26334 35374 26386 35426
rect 26386 35374 26388 35426
rect 26332 35372 26388 35374
rect 26492 35426 26548 35428
rect 26492 35374 26494 35426
rect 26494 35374 26546 35426
rect 26546 35374 26548 35426
rect 26492 35372 26548 35374
rect 26652 35426 26708 35428
rect 26652 35374 26654 35426
rect 26654 35374 26706 35426
rect 26706 35374 26708 35426
rect 26652 35372 26708 35374
rect 26812 35426 26868 35428
rect 26812 35374 26814 35426
rect 26814 35374 26866 35426
rect 26866 35374 26868 35426
rect 26812 35372 26868 35374
rect 26972 35426 27028 35428
rect 26972 35374 26974 35426
rect 26974 35374 27026 35426
rect 27026 35374 27028 35426
rect 26972 35372 27028 35374
rect 27132 35426 27188 35428
rect 27132 35374 27134 35426
rect 27134 35374 27186 35426
rect 27186 35374 27188 35426
rect 27132 35372 27188 35374
rect 27292 35426 27348 35428
rect 27292 35374 27294 35426
rect 27294 35374 27346 35426
rect 27346 35374 27348 35426
rect 27292 35372 27348 35374
rect 27452 35426 27508 35428
rect 27452 35374 27454 35426
rect 27454 35374 27506 35426
rect 27506 35374 27508 35426
rect 27452 35372 27508 35374
rect 27612 35426 27668 35428
rect 27612 35374 27614 35426
rect 27614 35374 27666 35426
rect 27666 35374 27668 35426
rect 27612 35372 27668 35374
rect 27772 35426 27828 35428
rect 27772 35374 27774 35426
rect 27774 35374 27826 35426
rect 27826 35374 27828 35426
rect 27772 35372 27828 35374
rect 27932 35426 27988 35428
rect 27932 35374 27934 35426
rect 27934 35374 27986 35426
rect 27986 35374 27988 35426
rect 27932 35372 27988 35374
rect 28092 35426 28148 35428
rect 28092 35374 28094 35426
rect 28094 35374 28146 35426
rect 28146 35374 28148 35426
rect 28092 35372 28148 35374
rect 28252 35426 28308 35428
rect 28252 35374 28254 35426
rect 28254 35374 28306 35426
rect 28306 35374 28308 35426
rect 28252 35372 28308 35374
rect 28412 35426 28468 35428
rect 28412 35374 28414 35426
rect 28414 35374 28466 35426
rect 28466 35374 28468 35426
rect 28412 35372 28468 35374
rect 28572 35426 28628 35428
rect 28572 35374 28574 35426
rect 28574 35374 28626 35426
rect 28626 35374 28628 35426
rect 28572 35372 28628 35374
rect 28732 35426 28788 35428
rect 28732 35374 28734 35426
rect 28734 35374 28786 35426
rect 28786 35374 28788 35426
rect 28732 35372 28788 35374
rect 28892 35426 28948 35428
rect 28892 35374 28894 35426
rect 28894 35374 28946 35426
rect 28946 35374 28948 35426
rect 28892 35372 28948 35374
rect 29052 35426 29108 35428
rect 29052 35374 29054 35426
rect 29054 35374 29106 35426
rect 29106 35374 29108 35426
rect 29052 35372 29108 35374
rect 29212 35426 29268 35428
rect 29212 35374 29214 35426
rect 29214 35374 29266 35426
rect 29266 35374 29268 35426
rect 29212 35372 29268 35374
rect 29372 35426 29428 35428
rect 29372 35374 29374 35426
rect 29374 35374 29426 35426
rect 29426 35374 29428 35426
rect 29372 35372 29428 35374
rect 30492 35372 30548 35428
rect 30812 35372 30868 35428
rect 31132 35372 31188 35428
rect 31452 35372 31508 35428
rect 31772 35372 31828 35428
rect 32092 35372 32148 35428
rect 32412 35372 32468 35428
rect 33532 35426 33588 35428
rect 33532 35374 33534 35426
rect 33534 35374 33586 35426
rect 33586 35374 33588 35426
rect 33532 35372 33588 35374
rect 33692 35426 33748 35428
rect 33692 35374 33694 35426
rect 33694 35374 33746 35426
rect 33746 35374 33748 35426
rect 33692 35372 33748 35374
rect 33852 35426 33908 35428
rect 33852 35374 33854 35426
rect 33854 35374 33906 35426
rect 33906 35374 33908 35426
rect 33852 35372 33908 35374
rect 34012 35426 34068 35428
rect 34012 35374 34014 35426
rect 34014 35374 34066 35426
rect 34066 35374 34068 35426
rect 34012 35372 34068 35374
rect 34172 35426 34228 35428
rect 34172 35374 34174 35426
rect 34174 35374 34226 35426
rect 34226 35374 34228 35426
rect 34172 35372 34228 35374
rect 34332 35426 34388 35428
rect 34332 35374 34334 35426
rect 34334 35374 34386 35426
rect 34386 35374 34388 35426
rect 34332 35372 34388 35374
rect 34492 35426 34548 35428
rect 34492 35374 34494 35426
rect 34494 35374 34546 35426
rect 34546 35374 34548 35426
rect 34492 35372 34548 35374
rect 34652 35426 34708 35428
rect 34652 35374 34654 35426
rect 34654 35374 34706 35426
rect 34706 35374 34708 35426
rect 34652 35372 34708 35374
rect 34812 35426 34868 35428
rect 34812 35374 34814 35426
rect 34814 35374 34866 35426
rect 34866 35374 34868 35426
rect 34812 35372 34868 35374
rect 34972 35426 35028 35428
rect 34972 35374 34974 35426
rect 34974 35374 35026 35426
rect 35026 35374 35028 35426
rect 34972 35372 35028 35374
rect 35132 35426 35188 35428
rect 35132 35374 35134 35426
rect 35134 35374 35186 35426
rect 35186 35374 35188 35426
rect 35132 35372 35188 35374
rect 35292 35426 35348 35428
rect 35292 35374 35294 35426
rect 35294 35374 35346 35426
rect 35346 35374 35348 35426
rect 35292 35372 35348 35374
rect 35452 35426 35508 35428
rect 35452 35374 35454 35426
rect 35454 35374 35506 35426
rect 35506 35374 35508 35426
rect 35452 35372 35508 35374
rect 35612 35426 35668 35428
rect 35612 35374 35614 35426
rect 35614 35374 35666 35426
rect 35666 35374 35668 35426
rect 35612 35372 35668 35374
rect 35772 35426 35828 35428
rect 35772 35374 35774 35426
rect 35774 35374 35826 35426
rect 35826 35374 35828 35426
rect 35772 35372 35828 35374
rect 35932 35426 35988 35428
rect 35932 35374 35934 35426
rect 35934 35374 35986 35426
rect 35986 35374 35988 35426
rect 35932 35372 35988 35374
rect 36092 35426 36148 35428
rect 36092 35374 36094 35426
rect 36094 35374 36146 35426
rect 36146 35374 36148 35426
rect 36092 35372 36148 35374
rect 36252 35426 36308 35428
rect 36252 35374 36254 35426
rect 36254 35374 36306 35426
rect 36306 35374 36308 35426
rect 36252 35372 36308 35374
rect 36412 35426 36468 35428
rect 36412 35374 36414 35426
rect 36414 35374 36466 35426
rect 36466 35374 36468 35426
rect 36412 35372 36468 35374
rect 36572 35426 36628 35428
rect 36572 35374 36574 35426
rect 36574 35374 36626 35426
rect 36626 35374 36628 35426
rect 36572 35372 36628 35374
rect 36732 35426 36788 35428
rect 36732 35374 36734 35426
rect 36734 35374 36786 35426
rect 36786 35374 36788 35426
rect 36732 35372 36788 35374
rect 36892 35426 36948 35428
rect 36892 35374 36894 35426
rect 36894 35374 36946 35426
rect 36946 35374 36948 35426
rect 36892 35372 36948 35374
rect 37052 35426 37108 35428
rect 37052 35374 37054 35426
rect 37054 35374 37106 35426
rect 37106 35374 37108 35426
rect 37052 35372 37108 35374
rect 37212 35426 37268 35428
rect 37212 35374 37214 35426
rect 37214 35374 37266 35426
rect 37266 35374 37268 35426
rect 37212 35372 37268 35374
rect 37372 35426 37428 35428
rect 37372 35374 37374 35426
rect 37374 35374 37426 35426
rect 37426 35374 37428 35426
rect 37372 35372 37428 35374
rect 37532 35426 37588 35428
rect 37532 35374 37534 35426
rect 37534 35374 37586 35426
rect 37586 35374 37588 35426
rect 37532 35372 37588 35374
rect 37692 35426 37748 35428
rect 37692 35374 37694 35426
rect 37694 35374 37746 35426
rect 37746 35374 37748 35426
rect 37692 35372 37748 35374
rect 37852 35426 37908 35428
rect 37852 35374 37854 35426
rect 37854 35374 37906 35426
rect 37906 35374 37908 35426
rect 37852 35372 37908 35374
rect 38012 35426 38068 35428
rect 38012 35374 38014 35426
rect 38014 35374 38066 35426
rect 38066 35374 38068 35426
rect 38012 35372 38068 35374
rect 38172 35426 38228 35428
rect 38172 35374 38174 35426
rect 38174 35374 38226 35426
rect 38226 35374 38228 35426
rect 38172 35372 38228 35374
rect 38332 35426 38388 35428
rect 38332 35374 38334 35426
rect 38334 35374 38386 35426
rect 38386 35374 38388 35426
rect 38332 35372 38388 35374
rect 38492 35426 38548 35428
rect 38492 35374 38494 35426
rect 38494 35374 38546 35426
rect 38546 35374 38548 35426
rect 38492 35372 38548 35374
rect 38652 35426 38708 35428
rect 38652 35374 38654 35426
rect 38654 35374 38706 35426
rect 38706 35374 38708 35426
rect 38652 35372 38708 35374
rect 38812 35426 38868 35428
rect 38812 35374 38814 35426
rect 38814 35374 38866 35426
rect 38866 35374 38868 35426
rect 38812 35372 38868 35374
rect 38972 35426 39028 35428
rect 38972 35374 38974 35426
rect 38974 35374 39026 35426
rect 39026 35374 39028 35426
rect 38972 35372 39028 35374
rect 39132 35426 39188 35428
rect 39132 35374 39134 35426
rect 39134 35374 39186 35426
rect 39186 35374 39188 35426
rect 39132 35372 39188 35374
rect 39292 35426 39348 35428
rect 39292 35374 39294 35426
rect 39294 35374 39346 35426
rect 39346 35374 39348 35426
rect 39292 35372 39348 35374
rect 39452 35426 39508 35428
rect 39452 35374 39454 35426
rect 39454 35374 39506 35426
rect 39506 35374 39508 35426
rect 39452 35372 39508 35374
rect 39612 35426 39668 35428
rect 39612 35374 39614 35426
rect 39614 35374 39666 35426
rect 39666 35374 39668 35426
rect 39612 35372 39668 35374
rect 39772 35426 39828 35428
rect 39772 35374 39774 35426
rect 39774 35374 39826 35426
rect 39826 35374 39828 35426
rect 39772 35372 39828 35374
rect 39932 35426 39988 35428
rect 39932 35374 39934 35426
rect 39934 35374 39986 35426
rect 39986 35374 39988 35426
rect 39932 35372 39988 35374
rect 40092 35426 40148 35428
rect 40092 35374 40094 35426
rect 40094 35374 40146 35426
rect 40146 35374 40148 35426
rect 40092 35372 40148 35374
rect 40252 35426 40308 35428
rect 40252 35374 40254 35426
rect 40254 35374 40306 35426
rect 40306 35374 40308 35426
rect 40252 35372 40308 35374
rect 40412 35426 40468 35428
rect 40412 35374 40414 35426
rect 40414 35374 40466 35426
rect 40466 35374 40468 35426
rect 40412 35372 40468 35374
rect 40572 35426 40628 35428
rect 40572 35374 40574 35426
rect 40574 35374 40626 35426
rect 40626 35374 40628 35426
rect 40572 35372 40628 35374
rect 40732 35426 40788 35428
rect 40732 35374 40734 35426
rect 40734 35374 40786 35426
rect 40786 35374 40788 35426
rect 40732 35372 40788 35374
rect 40892 35426 40948 35428
rect 40892 35374 40894 35426
rect 40894 35374 40946 35426
rect 40946 35374 40948 35426
rect 40892 35372 40948 35374
rect 41052 35426 41108 35428
rect 41052 35374 41054 35426
rect 41054 35374 41106 35426
rect 41106 35374 41108 35426
rect 41052 35372 41108 35374
rect 41212 35426 41268 35428
rect 41212 35374 41214 35426
rect 41214 35374 41266 35426
rect 41266 35374 41268 35426
rect 41212 35372 41268 35374
rect 41372 35426 41428 35428
rect 41372 35374 41374 35426
rect 41374 35374 41426 35426
rect 41426 35374 41428 35426
rect 41372 35372 41428 35374
rect 41532 35426 41588 35428
rect 41532 35374 41534 35426
rect 41534 35374 41586 35426
rect 41586 35374 41588 35426
rect 41532 35372 41588 35374
rect 41692 35426 41748 35428
rect 41692 35374 41694 35426
rect 41694 35374 41746 35426
rect 41746 35374 41748 35426
rect 41692 35372 41748 35374
rect 41852 35426 41908 35428
rect 41852 35374 41854 35426
rect 41854 35374 41906 35426
rect 41906 35374 41908 35426
rect 41852 35372 41908 35374
rect 10572 35212 10628 35268
rect 20812 35212 20868 35268
rect 31292 35212 31348 35268
rect 12 35106 68 35108
rect 12 35054 14 35106
rect 14 35054 66 35106
rect 66 35054 68 35106
rect 12 35052 68 35054
rect 172 35106 228 35108
rect 172 35054 174 35106
rect 174 35054 226 35106
rect 226 35054 228 35106
rect 172 35052 228 35054
rect 332 35106 388 35108
rect 332 35054 334 35106
rect 334 35054 386 35106
rect 386 35054 388 35106
rect 332 35052 388 35054
rect 492 35106 548 35108
rect 492 35054 494 35106
rect 494 35054 546 35106
rect 546 35054 548 35106
rect 492 35052 548 35054
rect 652 35106 708 35108
rect 652 35054 654 35106
rect 654 35054 706 35106
rect 706 35054 708 35106
rect 652 35052 708 35054
rect 812 35106 868 35108
rect 812 35054 814 35106
rect 814 35054 866 35106
rect 866 35054 868 35106
rect 812 35052 868 35054
rect 972 35106 1028 35108
rect 972 35054 974 35106
rect 974 35054 1026 35106
rect 1026 35054 1028 35106
rect 972 35052 1028 35054
rect 1132 35106 1188 35108
rect 1132 35054 1134 35106
rect 1134 35054 1186 35106
rect 1186 35054 1188 35106
rect 1132 35052 1188 35054
rect 1292 35106 1348 35108
rect 1292 35054 1294 35106
rect 1294 35054 1346 35106
rect 1346 35054 1348 35106
rect 1292 35052 1348 35054
rect 1452 35106 1508 35108
rect 1452 35054 1454 35106
rect 1454 35054 1506 35106
rect 1506 35054 1508 35106
rect 1452 35052 1508 35054
rect 1612 35106 1668 35108
rect 1612 35054 1614 35106
rect 1614 35054 1666 35106
rect 1666 35054 1668 35106
rect 1612 35052 1668 35054
rect 1772 35106 1828 35108
rect 1772 35054 1774 35106
rect 1774 35054 1826 35106
rect 1826 35054 1828 35106
rect 1772 35052 1828 35054
rect 1932 35106 1988 35108
rect 1932 35054 1934 35106
rect 1934 35054 1986 35106
rect 1986 35054 1988 35106
rect 1932 35052 1988 35054
rect 2092 35106 2148 35108
rect 2092 35054 2094 35106
rect 2094 35054 2146 35106
rect 2146 35054 2148 35106
rect 2092 35052 2148 35054
rect 2252 35106 2308 35108
rect 2252 35054 2254 35106
rect 2254 35054 2306 35106
rect 2306 35054 2308 35106
rect 2252 35052 2308 35054
rect 2412 35106 2468 35108
rect 2412 35054 2414 35106
rect 2414 35054 2466 35106
rect 2466 35054 2468 35106
rect 2412 35052 2468 35054
rect 2572 35106 2628 35108
rect 2572 35054 2574 35106
rect 2574 35054 2626 35106
rect 2626 35054 2628 35106
rect 2572 35052 2628 35054
rect 2732 35106 2788 35108
rect 2732 35054 2734 35106
rect 2734 35054 2786 35106
rect 2786 35054 2788 35106
rect 2732 35052 2788 35054
rect 2892 35106 2948 35108
rect 2892 35054 2894 35106
rect 2894 35054 2946 35106
rect 2946 35054 2948 35106
rect 2892 35052 2948 35054
rect 3052 35106 3108 35108
rect 3052 35054 3054 35106
rect 3054 35054 3106 35106
rect 3106 35054 3108 35106
rect 3052 35052 3108 35054
rect 3212 35106 3268 35108
rect 3212 35054 3214 35106
rect 3214 35054 3266 35106
rect 3266 35054 3268 35106
rect 3212 35052 3268 35054
rect 3372 35106 3428 35108
rect 3372 35054 3374 35106
rect 3374 35054 3426 35106
rect 3426 35054 3428 35106
rect 3372 35052 3428 35054
rect 3532 35106 3588 35108
rect 3532 35054 3534 35106
rect 3534 35054 3586 35106
rect 3586 35054 3588 35106
rect 3532 35052 3588 35054
rect 3692 35106 3748 35108
rect 3692 35054 3694 35106
rect 3694 35054 3746 35106
rect 3746 35054 3748 35106
rect 3692 35052 3748 35054
rect 3852 35106 3908 35108
rect 3852 35054 3854 35106
rect 3854 35054 3906 35106
rect 3906 35054 3908 35106
rect 3852 35052 3908 35054
rect 4012 35106 4068 35108
rect 4012 35054 4014 35106
rect 4014 35054 4066 35106
rect 4066 35054 4068 35106
rect 4012 35052 4068 35054
rect 4172 35106 4228 35108
rect 4172 35054 4174 35106
rect 4174 35054 4226 35106
rect 4226 35054 4228 35106
rect 4172 35052 4228 35054
rect 4332 35106 4388 35108
rect 4332 35054 4334 35106
rect 4334 35054 4386 35106
rect 4386 35054 4388 35106
rect 4332 35052 4388 35054
rect 4492 35106 4548 35108
rect 4492 35054 4494 35106
rect 4494 35054 4546 35106
rect 4546 35054 4548 35106
rect 4492 35052 4548 35054
rect 4652 35106 4708 35108
rect 4652 35054 4654 35106
rect 4654 35054 4706 35106
rect 4706 35054 4708 35106
rect 4652 35052 4708 35054
rect 4812 35106 4868 35108
rect 4812 35054 4814 35106
rect 4814 35054 4866 35106
rect 4866 35054 4868 35106
rect 4812 35052 4868 35054
rect 4972 35106 5028 35108
rect 4972 35054 4974 35106
rect 4974 35054 5026 35106
rect 5026 35054 5028 35106
rect 4972 35052 5028 35054
rect 5132 35106 5188 35108
rect 5132 35054 5134 35106
rect 5134 35054 5186 35106
rect 5186 35054 5188 35106
rect 5132 35052 5188 35054
rect 5292 35106 5348 35108
rect 5292 35054 5294 35106
rect 5294 35054 5346 35106
rect 5346 35054 5348 35106
rect 5292 35052 5348 35054
rect 5452 35106 5508 35108
rect 5452 35054 5454 35106
rect 5454 35054 5506 35106
rect 5506 35054 5508 35106
rect 5452 35052 5508 35054
rect 5612 35106 5668 35108
rect 5612 35054 5614 35106
rect 5614 35054 5666 35106
rect 5666 35054 5668 35106
rect 5612 35052 5668 35054
rect 5772 35106 5828 35108
rect 5772 35054 5774 35106
rect 5774 35054 5826 35106
rect 5826 35054 5828 35106
rect 5772 35052 5828 35054
rect 5932 35106 5988 35108
rect 5932 35054 5934 35106
rect 5934 35054 5986 35106
rect 5986 35054 5988 35106
rect 5932 35052 5988 35054
rect 6092 35106 6148 35108
rect 6092 35054 6094 35106
rect 6094 35054 6146 35106
rect 6146 35054 6148 35106
rect 6092 35052 6148 35054
rect 6252 35106 6308 35108
rect 6252 35054 6254 35106
rect 6254 35054 6306 35106
rect 6306 35054 6308 35106
rect 6252 35052 6308 35054
rect 6412 35106 6468 35108
rect 6412 35054 6414 35106
rect 6414 35054 6466 35106
rect 6466 35054 6468 35106
rect 6412 35052 6468 35054
rect 6572 35106 6628 35108
rect 6572 35054 6574 35106
rect 6574 35054 6626 35106
rect 6626 35054 6628 35106
rect 6572 35052 6628 35054
rect 6732 35106 6788 35108
rect 6732 35054 6734 35106
rect 6734 35054 6786 35106
rect 6786 35054 6788 35106
rect 6732 35052 6788 35054
rect 6892 35106 6948 35108
rect 6892 35054 6894 35106
rect 6894 35054 6946 35106
rect 6946 35054 6948 35106
rect 6892 35052 6948 35054
rect 7052 35106 7108 35108
rect 7052 35054 7054 35106
rect 7054 35054 7106 35106
rect 7106 35054 7108 35106
rect 7052 35052 7108 35054
rect 7212 35106 7268 35108
rect 7212 35054 7214 35106
rect 7214 35054 7266 35106
rect 7266 35054 7268 35106
rect 7212 35052 7268 35054
rect 7372 35106 7428 35108
rect 7372 35054 7374 35106
rect 7374 35054 7426 35106
rect 7426 35054 7428 35106
rect 7372 35052 7428 35054
rect 7532 35106 7588 35108
rect 7532 35054 7534 35106
rect 7534 35054 7586 35106
rect 7586 35054 7588 35106
rect 7532 35052 7588 35054
rect 7692 35106 7748 35108
rect 7692 35054 7694 35106
rect 7694 35054 7746 35106
rect 7746 35054 7748 35106
rect 7692 35052 7748 35054
rect 7852 35106 7908 35108
rect 7852 35054 7854 35106
rect 7854 35054 7906 35106
rect 7906 35054 7908 35106
rect 7852 35052 7908 35054
rect 8012 35106 8068 35108
rect 8012 35054 8014 35106
rect 8014 35054 8066 35106
rect 8066 35054 8068 35106
rect 8012 35052 8068 35054
rect 8172 35106 8228 35108
rect 8172 35054 8174 35106
rect 8174 35054 8226 35106
rect 8226 35054 8228 35106
rect 8172 35052 8228 35054
rect 8332 35106 8388 35108
rect 8332 35054 8334 35106
rect 8334 35054 8386 35106
rect 8386 35054 8388 35106
rect 8332 35052 8388 35054
rect 9452 35052 9508 35108
rect 9772 35052 9828 35108
rect 10092 35052 10148 35108
rect 10412 35052 10468 35108
rect 10732 35052 10788 35108
rect 11052 35052 11108 35108
rect 11372 35052 11428 35108
rect 12492 35106 12548 35108
rect 12492 35054 12494 35106
rect 12494 35054 12546 35106
rect 12546 35054 12548 35106
rect 12492 35052 12548 35054
rect 12652 35106 12708 35108
rect 12652 35054 12654 35106
rect 12654 35054 12706 35106
rect 12706 35054 12708 35106
rect 12652 35052 12708 35054
rect 12812 35106 12868 35108
rect 12812 35054 12814 35106
rect 12814 35054 12866 35106
rect 12866 35054 12868 35106
rect 12812 35052 12868 35054
rect 12972 35106 13028 35108
rect 12972 35054 12974 35106
rect 12974 35054 13026 35106
rect 13026 35054 13028 35106
rect 12972 35052 13028 35054
rect 13132 35106 13188 35108
rect 13132 35054 13134 35106
rect 13134 35054 13186 35106
rect 13186 35054 13188 35106
rect 13132 35052 13188 35054
rect 13292 35106 13348 35108
rect 13292 35054 13294 35106
rect 13294 35054 13346 35106
rect 13346 35054 13348 35106
rect 13292 35052 13348 35054
rect 13452 35106 13508 35108
rect 13452 35054 13454 35106
rect 13454 35054 13506 35106
rect 13506 35054 13508 35106
rect 13452 35052 13508 35054
rect 13612 35106 13668 35108
rect 13612 35054 13614 35106
rect 13614 35054 13666 35106
rect 13666 35054 13668 35106
rect 13612 35052 13668 35054
rect 13772 35106 13828 35108
rect 13772 35054 13774 35106
rect 13774 35054 13826 35106
rect 13826 35054 13828 35106
rect 13772 35052 13828 35054
rect 13932 35106 13988 35108
rect 13932 35054 13934 35106
rect 13934 35054 13986 35106
rect 13986 35054 13988 35106
rect 13932 35052 13988 35054
rect 14092 35106 14148 35108
rect 14092 35054 14094 35106
rect 14094 35054 14146 35106
rect 14146 35054 14148 35106
rect 14092 35052 14148 35054
rect 14252 35106 14308 35108
rect 14252 35054 14254 35106
rect 14254 35054 14306 35106
rect 14306 35054 14308 35106
rect 14252 35052 14308 35054
rect 14412 35106 14468 35108
rect 14412 35054 14414 35106
rect 14414 35054 14466 35106
rect 14466 35054 14468 35106
rect 14412 35052 14468 35054
rect 14572 35106 14628 35108
rect 14572 35054 14574 35106
rect 14574 35054 14626 35106
rect 14626 35054 14628 35106
rect 14572 35052 14628 35054
rect 14732 35106 14788 35108
rect 14732 35054 14734 35106
rect 14734 35054 14786 35106
rect 14786 35054 14788 35106
rect 14732 35052 14788 35054
rect 14892 35106 14948 35108
rect 14892 35054 14894 35106
rect 14894 35054 14946 35106
rect 14946 35054 14948 35106
rect 14892 35052 14948 35054
rect 15052 35106 15108 35108
rect 15052 35054 15054 35106
rect 15054 35054 15106 35106
rect 15106 35054 15108 35106
rect 15052 35052 15108 35054
rect 15212 35106 15268 35108
rect 15212 35054 15214 35106
rect 15214 35054 15266 35106
rect 15266 35054 15268 35106
rect 15212 35052 15268 35054
rect 15372 35106 15428 35108
rect 15372 35054 15374 35106
rect 15374 35054 15426 35106
rect 15426 35054 15428 35106
rect 15372 35052 15428 35054
rect 15532 35106 15588 35108
rect 15532 35054 15534 35106
rect 15534 35054 15586 35106
rect 15586 35054 15588 35106
rect 15532 35052 15588 35054
rect 15692 35106 15748 35108
rect 15692 35054 15694 35106
rect 15694 35054 15746 35106
rect 15746 35054 15748 35106
rect 15692 35052 15748 35054
rect 15852 35106 15908 35108
rect 15852 35054 15854 35106
rect 15854 35054 15906 35106
rect 15906 35054 15908 35106
rect 15852 35052 15908 35054
rect 16012 35106 16068 35108
rect 16012 35054 16014 35106
rect 16014 35054 16066 35106
rect 16066 35054 16068 35106
rect 16012 35052 16068 35054
rect 16172 35106 16228 35108
rect 16172 35054 16174 35106
rect 16174 35054 16226 35106
rect 16226 35054 16228 35106
rect 16172 35052 16228 35054
rect 16332 35106 16388 35108
rect 16332 35054 16334 35106
rect 16334 35054 16386 35106
rect 16386 35054 16388 35106
rect 16332 35052 16388 35054
rect 16492 35106 16548 35108
rect 16492 35054 16494 35106
rect 16494 35054 16546 35106
rect 16546 35054 16548 35106
rect 16492 35052 16548 35054
rect 16652 35106 16708 35108
rect 16652 35054 16654 35106
rect 16654 35054 16706 35106
rect 16706 35054 16708 35106
rect 16652 35052 16708 35054
rect 16812 35106 16868 35108
rect 16812 35054 16814 35106
rect 16814 35054 16866 35106
rect 16866 35054 16868 35106
rect 16812 35052 16868 35054
rect 16972 35106 17028 35108
rect 16972 35054 16974 35106
rect 16974 35054 17026 35106
rect 17026 35054 17028 35106
rect 16972 35052 17028 35054
rect 17132 35106 17188 35108
rect 17132 35054 17134 35106
rect 17134 35054 17186 35106
rect 17186 35054 17188 35106
rect 17132 35052 17188 35054
rect 17292 35106 17348 35108
rect 17292 35054 17294 35106
rect 17294 35054 17346 35106
rect 17346 35054 17348 35106
rect 17292 35052 17348 35054
rect 17452 35106 17508 35108
rect 17452 35054 17454 35106
rect 17454 35054 17506 35106
rect 17506 35054 17508 35106
rect 17452 35052 17508 35054
rect 17612 35106 17668 35108
rect 17612 35054 17614 35106
rect 17614 35054 17666 35106
rect 17666 35054 17668 35106
rect 17612 35052 17668 35054
rect 17772 35106 17828 35108
rect 17772 35054 17774 35106
rect 17774 35054 17826 35106
rect 17826 35054 17828 35106
rect 17772 35052 17828 35054
rect 17932 35106 17988 35108
rect 17932 35054 17934 35106
rect 17934 35054 17986 35106
rect 17986 35054 17988 35106
rect 17932 35052 17988 35054
rect 18092 35106 18148 35108
rect 18092 35054 18094 35106
rect 18094 35054 18146 35106
rect 18146 35054 18148 35106
rect 18092 35052 18148 35054
rect 18252 35106 18308 35108
rect 18252 35054 18254 35106
rect 18254 35054 18306 35106
rect 18306 35054 18308 35106
rect 18252 35052 18308 35054
rect 18412 35106 18468 35108
rect 18412 35054 18414 35106
rect 18414 35054 18466 35106
rect 18466 35054 18468 35106
rect 18412 35052 18468 35054
rect 18572 35106 18628 35108
rect 18572 35054 18574 35106
rect 18574 35054 18626 35106
rect 18626 35054 18628 35106
rect 18572 35052 18628 35054
rect 18732 35106 18788 35108
rect 18732 35054 18734 35106
rect 18734 35054 18786 35106
rect 18786 35054 18788 35106
rect 18732 35052 18788 35054
rect 18892 35106 18948 35108
rect 18892 35054 18894 35106
rect 18894 35054 18946 35106
rect 18946 35054 18948 35106
rect 18892 35052 18948 35054
rect 20012 35052 20068 35108
rect 20332 35052 20388 35108
rect 20652 35052 20708 35108
rect 20972 35052 21028 35108
rect 21292 35052 21348 35108
rect 21612 35052 21668 35108
rect 21932 35052 21988 35108
rect 23132 35106 23188 35108
rect 23132 35054 23134 35106
rect 23134 35054 23186 35106
rect 23186 35054 23188 35106
rect 23132 35052 23188 35054
rect 23292 35106 23348 35108
rect 23292 35054 23294 35106
rect 23294 35054 23346 35106
rect 23346 35054 23348 35106
rect 23292 35052 23348 35054
rect 23452 35106 23508 35108
rect 23452 35054 23454 35106
rect 23454 35054 23506 35106
rect 23506 35054 23508 35106
rect 23452 35052 23508 35054
rect 23612 35106 23668 35108
rect 23612 35054 23614 35106
rect 23614 35054 23666 35106
rect 23666 35054 23668 35106
rect 23612 35052 23668 35054
rect 23772 35106 23828 35108
rect 23772 35054 23774 35106
rect 23774 35054 23826 35106
rect 23826 35054 23828 35106
rect 23772 35052 23828 35054
rect 23932 35106 23988 35108
rect 23932 35054 23934 35106
rect 23934 35054 23986 35106
rect 23986 35054 23988 35106
rect 23932 35052 23988 35054
rect 24092 35106 24148 35108
rect 24092 35054 24094 35106
rect 24094 35054 24146 35106
rect 24146 35054 24148 35106
rect 24092 35052 24148 35054
rect 24252 35106 24308 35108
rect 24252 35054 24254 35106
rect 24254 35054 24306 35106
rect 24306 35054 24308 35106
rect 24252 35052 24308 35054
rect 24412 35106 24468 35108
rect 24412 35054 24414 35106
rect 24414 35054 24466 35106
rect 24466 35054 24468 35106
rect 24412 35052 24468 35054
rect 24572 35106 24628 35108
rect 24572 35054 24574 35106
rect 24574 35054 24626 35106
rect 24626 35054 24628 35106
rect 24572 35052 24628 35054
rect 24732 35106 24788 35108
rect 24732 35054 24734 35106
rect 24734 35054 24786 35106
rect 24786 35054 24788 35106
rect 24732 35052 24788 35054
rect 24892 35106 24948 35108
rect 24892 35054 24894 35106
rect 24894 35054 24946 35106
rect 24946 35054 24948 35106
rect 24892 35052 24948 35054
rect 25052 35106 25108 35108
rect 25052 35054 25054 35106
rect 25054 35054 25106 35106
rect 25106 35054 25108 35106
rect 25052 35052 25108 35054
rect 25212 35106 25268 35108
rect 25212 35054 25214 35106
rect 25214 35054 25266 35106
rect 25266 35054 25268 35106
rect 25212 35052 25268 35054
rect 25372 35106 25428 35108
rect 25372 35054 25374 35106
rect 25374 35054 25426 35106
rect 25426 35054 25428 35106
rect 25372 35052 25428 35054
rect 25532 35106 25588 35108
rect 25532 35054 25534 35106
rect 25534 35054 25586 35106
rect 25586 35054 25588 35106
rect 25532 35052 25588 35054
rect 25692 35106 25748 35108
rect 25692 35054 25694 35106
rect 25694 35054 25746 35106
rect 25746 35054 25748 35106
rect 25692 35052 25748 35054
rect 25852 35106 25908 35108
rect 25852 35054 25854 35106
rect 25854 35054 25906 35106
rect 25906 35054 25908 35106
rect 25852 35052 25908 35054
rect 26012 35106 26068 35108
rect 26012 35054 26014 35106
rect 26014 35054 26066 35106
rect 26066 35054 26068 35106
rect 26012 35052 26068 35054
rect 26172 35106 26228 35108
rect 26172 35054 26174 35106
rect 26174 35054 26226 35106
rect 26226 35054 26228 35106
rect 26172 35052 26228 35054
rect 26332 35106 26388 35108
rect 26332 35054 26334 35106
rect 26334 35054 26386 35106
rect 26386 35054 26388 35106
rect 26332 35052 26388 35054
rect 26492 35106 26548 35108
rect 26492 35054 26494 35106
rect 26494 35054 26546 35106
rect 26546 35054 26548 35106
rect 26492 35052 26548 35054
rect 26652 35106 26708 35108
rect 26652 35054 26654 35106
rect 26654 35054 26706 35106
rect 26706 35054 26708 35106
rect 26652 35052 26708 35054
rect 26812 35106 26868 35108
rect 26812 35054 26814 35106
rect 26814 35054 26866 35106
rect 26866 35054 26868 35106
rect 26812 35052 26868 35054
rect 26972 35106 27028 35108
rect 26972 35054 26974 35106
rect 26974 35054 27026 35106
rect 27026 35054 27028 35106
rect 26972 35052 27028 35054
rect 27132 35106 27188 35108
rect 27132 35054 27134 35106
rect 27134 35054 27186 35106
rect 27186 35054 27188 35106
rect 27132 35052 27188 35054
rect 27292 35106 27348 35108
rect 27292 35054 27294 35106
rect 27294 35054 27346 35106
rect 27346 35054 27348 35106
rect 27292 35052 27348 35054
rect 27452 35106 27508 35108
rect 27452 35054 27454 35106
rect 27454 35054 27506 35106
rect 27506 35054 27508 35106
rect 27452 35052 27508 35054
rect 27612 35106 27668 35108
rect 27612 35054 27614 35106
rect 27614 35054 27666 35106
rect 27666 35054 27668 35106
rect 27612 35052 27668 35054
rect 27772 35106 27828 35108
rect 27772 35054 27774 35106
rect 27774 35054 27826 35106
rect 27826 35054 27828 35106
rect 27772 35052 27828 35054
rect 27932 35106 27988 35108
rect 27932 35054 27934 35106
rect 27934 35054 27986 35106
rect 27986 35054 27988 35106
rect 27932 35052 27988 35054
rect 28092 35106 28148 35108
rect 28092 35054 28094 35106
rect 28094 35054 28146 35106
rect 28146 35054 28148 35106
rect 28092 35052 28148 35054
rect 28252 35106 28308 35108
rect 28252 35054 28254 35106
rect 28254 35054 28306 35106
rect 28306 35054 28308 35106
rect 28252 35052 28308 35054
rect 28412 35106 28468 35108
rect 28412 35054 28414 35106
rect 28414 35054 28466 35106
rect 28466 35054 28468 35106
rect 28412 35052 28468 35054
rect 28572 35106 28628 35108
rect 28572 35054 28574 35106
rect 28574 35054 28626 35106
rect 28626 35054 28628 35106
rect 28572 35052 28628 35054
rect 28732 35106 28788 35108
rect 28732 35054 28734 35106
rect 28734 35054 28786 35106
rect 28786 35054 28788 35106
rect 28732 35052 28788 35054
rect 28892 35106 28948 35108
rect 28892 35054 28894 35106
rect 28894 35054 28946 35106
rect 28946 35054 28948 35106
rect 28892 35052 28948 35054
rect 29052 35106 29108 35108
rect 29052 35054 29054 35106
rect 29054 35054 29106 35106
rect 29106 35054 29108 35106
rect 29052 35052 29108 35054
rect 29212 35106 29268 35108
rect 29212 35054 29214 35106
rect 29214 35054 29266 35106
rect 29266 35054 29268 35106
rect 29212 35052 29268 35054
rect 29372 35106 29428 35108
rect 29372 35054 29374 35106
rect 29374 35054 29426 35106
rect 29426 35054 29428 35106
rect 29372 35052 29428 35054
rect 30492 35052 30548 35108
rect 30812 35052 30868 35108
rect 31132 35052 31188 35108
rect 31452 35052 31508 35108
rect 31772 35052 31828 35108
rect 32092 35052 32148 35108
rect 32412 35052 32468 35108
rect 33532 35106 33588 35108
rect 33532 35054 33534 35106
rect 33534 35054 33586 35106
rect 33586 35054 33588 35106
rect 33532 35052 33588 35054
rect 33692 35106 33748 35108
rect 33692 35054 33694 35106
rect 33694 35054 33746 35106
rect 33746 35054 33748 35106
rect 33692 35052 33748 35054
rect 33852 35106 33908 35108
rect 33852 35054 33854 35106
rect 33854 35054 33906 35106
rect 33906 35054 33908 35106
rect 33852 35052 33908 35054
rect 34012 35106 34068 35108
rect 34012 35054 34014 35106
rect 34014 35054 34066 35106
rect 34066 35054 34068 35106
rect 34012 35052 34068 35054
rect 34172 35106 34228 35108
rect 34172 35054 34174 35106
rect 34174 35054 34226 35106
rect 34226 35054 34228 35106
rect 34172 35052 34228 35054
rect 34332 35106 34388 35108
rect 34332 35054 34334 35106
rect 34334 35054 34386 35106
rect 34386 35054 34388 35106
rect 34332 35052 34388 35054
rect 34492 35106 34548 35108
rect 34492 35054 34494 35106
rect 34494 35054 34546 35106
rect 34546 35054 34548 35106
rect 34492 35052 34548 35054
rect 34652 35106 34708 35108
rect 34652 35054 34654 35106
rect 34654 35054 34706 35106
rect 34706 35054 34708 35106
rect 34652 35052 34708 35054
rect 34812 35106 34868 35108
rect 34812 35054 34814 35106
rect 34814 35054 34866 35106
rect 34866 35054 34868 35106
rect 34812 35052 34868 35054
rect 34972 35106 35028 35108
rect 34972 35054 34974 35106
rect 34974 35054 35026 35106
rect 35026 35054 35028 35106
rect 34972 35052 35028 35054
rect 35132 35106 35188 35108
rect 35132 35054 35134 35106
rect 35134 35054 35186 35106
rect 35186 35054 35188 35106
rect 35132 35052 35188 35054
rect 35292 35106 35348 35108
rect 35292 35054 35294 35106
rect 35294 35054 35346 35106
rect 35346 35054 35348 35106
rect 35292 35052 35348 35054
rect 35452 35106 35508 35108
rect 35452 35054 35454 35106
rect 35454 35054 35506 35106
rect 35506 35054 35508 35106
rect 35452 35052 35508 35054
rect 35612 35106 35668 35108
rect 35612 35054 35614 35106
rect 35614 35054 35666 35106
rect 35666 35054 35668 35106
rect 35612 35052 35668 35054
rect 35772 35106 35828 35108
rect 35772 35054 35774 35106
rect 35774 35054 35826 35106
rect 35826 35054 35828 35106
rect 35772 35052 35828 35054
rect 35932 35106 35988 35108
rect 35932 35054 35934 35106
rect 35934 35054 35986 35106
rect 35986 35054 35988 35106
rect 35932 35052 35988 35054
rect 36092 35106 36148 35108
rect 36092 35054 36094 35106
rect 36094 35054 36146 35106
rect 36146 35054 36148 35106
rect 36092 35052 36148 35054
rect 36252 35106 36308 35108
rect 36252 35054 36254 35106
rect 36254 35054 36306 35106
rect 36306 35054 36308 35106
rect 36252 35052 36308 35054
rect 36412 35106 36468 35108
rect 36412 35054 36414 35106
rect 36414 35054 36466 35106
rect 36466 35054 36468 35106
rect 36412 35052 36468 35054
rect 36572 35106 36628 35108
rect 36572 35054 36574 35106
rect 36574 35054 36626 35106
rect 36626 35054 36628 35106
rect 36572 35052 36628 35054
rect 36732 35106 36788 35108
rect 36732 35054 36734 35106
rect 36734 35054 36786 35106
rect 36786 35054 36788 35106
rect 36732 35052 36788 35054
rect 36892 35106 36948 35108
rect 36892 35054 36894 35106
rect 36894 35054 36946 35106
rect 36946 35054 36948 35106
rect 36892 35052 36948 35054
rect 37052 35106 37108 35108
rect 37052 35054 37054 35106
rect 37054 35054 37106 35106
rect 37106 35054 37108 35106
rect 37052 35052 37108 35054
rect 37212 35106 37268 35108
rect 37212 35054 37214 35106
rect 37214 35054 37266 35106
rect 37266 35054 37268 35106
rect 37212 35052 37268 35054
rect 37372 35106 37428 35108
rect 37372 35054 37374 35106
rect 37374 35054 37426 35106
rect 37426 35054 37428 35106
rect 37372 35052 37428 35054
rect 37532 35106 37588 35108
rect 37532 35054 37534 35106
rect 37534 35054 37586 35106
rect 37586 35054 37588 35106
rect 37532 35052 37588 35054
rect 37692 35106 37748 35108
rect 37692 35054 37694 35106
rect 37694 35054 37746 35106
rect 37746 35054 37748 35106
rect 37692 35052 37748 35054
rect 37852 35106 37908 35108
rect 37852 35054 37854 35106
rect 37854 35054 37906 35106
rect 37906 35054 37908 35106
rect 37852 35052 37908 35054
rect 38012 35106 38068 35108
rect 38012 35054 38014 35106
rect 38014 35054 38066 35106
rect 38066 35054 38068 35106
rect 38012 35052 38068 35054
rect 38172 35106 38228 35108
rect 38172 35054 38174 35106
rect 38174 35054 38226 35106
rect 38226 35054 38228 35106
rect 38172 35052 38228 35054
rect 38332 35106 38388 35108
rect 38332 35054 38334 35106
rect 38334 35054 38386 35106
rect 38386 35054 38388 35106
rect 38332 35052 38388 35054
rect 38492 35106 38548 35108
rect 38492 35054 38494 35106
rect 38494 35054 38546 35106
rect 38546 35054 38548 35106
rect 38492 35052 38548 35054
rect 38652 35106 38708 35108
rect 38652 35054 38654 35106
rect 38654 35054 38706 35106
rect 38706 35054 38708 35106
rect 38652 35052 38708 35054
rect 38812 35106 38868 35108
rect 38812 35054 38814 35106
rect 38814 35054 38866 35106
rect 38866 35054 38868 35106
rect 38812 35052 38868 35054
rect 38972 35106 39028 35108
rect 38972 35054 38974 35106
rect 38974 35054 39026 35106
rect 39026 35054 39028 35106
rect 38972 35052 39028 35054
rect 39132 35106 39188 35108
rect 39132 35054 39134 35106
rect 39134 35054 39186 35106
rect 39186 35054 39188 35106
rect 39132 35052 39188 35054
rect 39292 35106 39348 35108
rect 39292 35054 39294 35106
rect 39294 35054 39346 35106
rect 39346 35054 39348 35106
rect 39292 35052 39348 35054
rect 39452 35106 39508 35108
rect 39452 35054 39454 35106
rect 39454 35054 39506 35106
rect 39506 35054 39508 35106
rect 39452 35052 39508 35054
rect 39612 35106 39668 35108
rect 39612 35054 39614 35106
rect 39614 35054 39666 35106
rect 39666 35054 39668 35106
rect 39612 35052 39668 35054
rect 39772 35106 39828 35108
rect 39772 35054 39774 35106
rect 39774 35054 39826 35106
rect 39826 35054 39828 35106
rect 39772 35052 39828 35054
rect 39932 35106 39988 35108
rect 39932 35054 39934 35106
rect 39934 35054 39986 35106
rect 39986 35054 39988 35106
rect 39932 35052 39988 35054
rect 40092 35106 40148 35108
rect 40092 35054 40094 35106
rect 40094 35054 40146 35106
rect 40146 35054 40148 35106
rect 40092 35052 40148 35054
rect 40252 35106 40308 35108
rect 40252 35054 40254 35106
rect 40254 35054 40306 35106
rect 40306 35054 40308 35106
rect 40252 35052 40308 35054
rect 40412 35106 40468 35108
rect 40412 35054 40414 35106
rect 40414 35054 40466 35106
rect 40466 35054 40468 35106
rect 40412 35052 40468 35054
rect 40572 35106 40628 35108
rect 40572 35054 40574 35106
rect 40574 35054 40626 35106
rect 40626 35054 40628 35106
rect 40572 35052 40628 35054
rect 40732 35106 40788 35108
rect 40732 35054 40734 35106
rect 40734 35054 40786 35106
rect 40786 35054 40788 35106
rect 40732 35052 40788 35054
rect 40892 35106 40948 35108
rect 40892 35054 40894 35106
rect 40894 35054 40946 35106
rect 40946 35054 40948 35106
rect 40892 35052 40948 35054
rect 41052 35106 41108 35108
rect 41052 35054 41054 35106
rect 41054 35054 41106 35106
rect 41106 35054 41108 35106
rect 41052 35052 41108 35054
rect 41212 35106 41268 35108
rect 41212 35054 41214 35106
rect 41214 35054 41266 35106
rect 41266 35054 41268 35106
rect 41212 35052 41268 35054
rect 41372 35106 41428 35108
rect 41372 35054 41374 35106
rect 41374 35054 41426 35106
rect 41426 35054 41428 35106
rect 41372 35052 41428 35054
rect 41532 35106 41588 35108
rect 41532 35054 41534 35106
rect 41534 35054 41586 35106
rect 41586 35054 41588 35106
rect 41532 35052 41588 35054
rect 41692 35106 41748 35108
rect 41692 35054 41694 35106
rect 41694 35054 41746 35106
rect 41746 35054 41748 35106
rect 41692 35052 41748 35054
rect 41852 35106 41908 35108
rect 41852 35054 41854 35106
rect 41854 35054 41906 35106
rect 41906 35054 41908 35106
rect 41852 35052 41908 35054
rect 10892 34892 10948 34948
rect 20492 34892 20548 34948
rect 30972 34892 31028 34948
rect 12 34786 68 34788
rect 12 34734 14 34786
rect 14 34734 66 34786
rect 66 34734 68 34786
rect 12 34732 68 34734
rect 172 34786 228 34788
rect 172 34734 174 34786
rect 174 34734 226 34786
rect 226 34734 228 34786
rect 172 34732 228 34734
rect 332 34786 388 34788
rect 332 34734 334 34786
rect 334 34734 386 34786
rect 386 34734 388 34786
rect 332 34732 388 34734
rect 492 34786 548 34788
rect 492 34734 494 34786
rect 494 34734 546 34786
rect 546 34734 548 34786
rect 492 34732 548 34734
rect 652 34786 708 34788
rect 652 34734 654 34786
rect 654 34734 706 34786
rect 706 34734 708 34786
rect 652 34732 708 34734
rect 812 34786 868 34788
rect 812 34734 814 34786
rect 814 34734 866 34786
rect 866 34734 868 34786
rect 812 34732 868 34734
rect 972 34786 1028 34788
rect 972 34734 974 34786
rect 974 34734 1026 34786
rect 1026 34734 1028 34786
rect 972 34732 1028 34734
rect 1132 34786 1188 34788
rect 1132 34734 1134 34786
rect 1134 34734 1186 34786
rect 1186 34734 1188 34786
rect 1132 34732 1188 34734
rect 1292 34786 1348 34788
rect 1292 34734 1294 34786
rect 1294 34734 1346 34786
rect 1346 34734 1348 34786
rect 1292 34732 1348 34734
rect 1452 34786 1508 34788
rect 1452 34734 1454 34786
rect 1454 34734 1506 34786
rect 1506 34734 1508 34786
rect 1452 34732 1508 34734
rect 1612 34786 1668 34788
rect 1612 34734 1614 34786
rect 1614 34734 1666 34786
rect 1666 34734 1668 34786
rect 1612 34732 1668 34734
rect 1772 34786 1828 34788
rect 1772 34734 1774 34786
rect 1774 34734 1826 34786
rect 1826 34734 1828 34786
rect 1772 34732 1828 34734
rect 1932 34786 1988 34788
rect 1932 34734 1934 34786
rect 1934 34734 1986 34786
rect 1986 34734 1988 34786
rect 1932 34732 1988 34734
rect 2092 34786 2148 34788
rect 2092 34734 2094 34786
rect 2094 34734 2146 34786
rect 2146 34734 2148 34786
rect 2092 34732 2148 34734
rect 2252 34786 2308 34788
rect 2252 34734 2254 34786
rect 2254 34734 2306 34786
rect 2306 34734 2308 34786
rect 2252 34732 2308 34734
rect 2412 34786 2468 34788
rect 2412 34734 2414 34786
rect 2414 34734 2466 34786
rect 2466 34734 2468 34786
rect 2412 34732 2468 34734
rect 2572 34786 2628 34788
rect 2572 34734 2574 34786
rect 2574 34734 2626 34786
rect 2626 34734 2628 34786
rect 2572 34732 2628 34734
rect 2732 34786 2788 34788
rect 2732 34734 2734 34786
rect 2734 34734 2786 34786
rect 2786 34734 2788 34786
rect 2732 34732 2788 34734
rect 2892 34786 2948 34788
rect 2892 34734 2894 34786
rect 2894 34734 2946 34786
rect 2946 34734 2948 34786
rect 2892 34732 2948 34734
rect 3052 34786 3108 34788
rect 3052 34734 3054 34786
rect 3054 34734 3106 34786
rect 3106 34734 3108 34786
rect 3052 34732 3108 34734
rect 3212 34786 3268 34788
rect 3212 34734 3214 34786
rect 3214 34734 3266 34786
rect 3266 34734 3268 34786
rect 3212 34732 3268 34734
rect 3372 34786 3428 34788
rect 3372 34734 3374 34786
rect 3374 34734 3426 34786
rect 3426 34734 3428 34786
rect 3372 34732 3428 34734
rect 3532 34786 3588 34788
rect 3532 34734 3534 34786
rect 3534 34734 3586 34786
rect 3586 34734 3588 34786
rect 3532 34732 3588 34734
rect 3692 34786 3748 34788
rect 3692 34734 3694 34786
rect 3694 34734 3746 34786
rect 3746 34734 3748 34786
rect 3692 34732 3748 34734
rect 3852 34786 3908 34788
rect 3852 34734 3854 34786
rect 3854 34734 3906 34786
rect 3906 34734 3908 34786
rect 3852 34732 3908 34734
rect 4012 34786 4068 34788
rect 4012 34734 4014 34786
rect 4014 34734 4066 34786
rect 4066 34734 4068 34786
rect 4012 34732 4068 34734
rect 4172 34786 4228 34788
rect 4172 34734 4174 34786
rect 4174 34734 4226 34786
rect 4226 34734 4228 34786
rect 4172 34732 4228 34734
rect 4332 34786 4388 34788
rect 4332 34734 4334 34786
rect 4334 34734 4386 34786
rect 4386 34734 4388 34786
rect 4332 34732 4388 34734
rect 4492 34786 4548 34788
rect 4492 34734 4494 34786
rect 4494 34734 4546 34786
rect 4546 34734 4548 34786
rect 4492 34732 4548 34734
rect 4652 34786 4708 34788
rect 4652 34734 4654 34786
rect 4654 34734 4706 34786
rect 4706 34734 4708 34786
rect 4652 34732 4708 34734
rect 4812 34786 4868 34788
rect 4812 34734 4814 34786
rect 4814 34734 4866 34786
rect 4866 34734 4868 34786
rect 4812 34732 4868 34734
rect 4972 34786 5028 34788
rect 4972 34734 4974 34786
rect 4974 34734 5026 34786
rect 5026 34734 5028 34786
rect 4972 34732 5028 34734
rect 5132 34786 5188 34788
rect 5132 34734 5134 34786
rect 5134 34734 5186 34786
rect 5186 34734 5188 34786
rect 5132 34732 5188 34734
rect 5292 34786 5348 34788
rect 5292 34734 5294 34786
rect 5294 34734 5346 34786
rect 5346 34734 5348 34786
rect 5292 34732 5348 34734
rect 5452 34786 5508 34788
rect 5452 34734 5454 34786
rect 5454 34734 5506 34786
rect 5506 34734 5508 34786
rect 5452 34732 5508 34734
rect 5612 34786 5668 34788
rect 5612 34734 5614 34786
rect 5614 34734 5666 34786
rect 5666 34734 5668 34786
rect 5612 34732 5668 34734
rect 5772 34786 5828 34788
rect 5772 34734 5774 34786
rect 5774 34734 5826 34786
rect 5826 34734 5828 34786
rect 5772 34732 5828 34734
rect 5932 34786 5988 34788
rect 5932 34734 5934 34786
rect 5934 34734 5986 34786
rect 5986 34734 5988 34786
rect 5932 34732 5988 34734
rect 6092 34786 6148 34788
rect 6092 34734 6094 34786
rect 6094 34734 6146 34786
rect 6146 34734 6148 34786
rect 6092 34732 6148 34734
rect 6252 34786 6308 34788
rect 6252 34734 6254 34786
rect 6254 34734 6306 34786
rect 6306 34734 6308 34786
rect 6252 34732 6308 34734
rect 6412 34786 6468 34788
rect 6412 34734 6414 34786
rect 6414 34734 6466 34786
rect 6466 34734 6468 34786
rect 6412 34732 6468 34734
rect 6572 34786 6628 34788
rect 6572 34734 6574 34786
rect 6574 34734 6626 34786
rect 6626 34734 6628 34786
rect 6572 34732 6628 34734
rect 6732 34786 6788 34788
rect 6732 34734 6734 34786
rect 6734 34734 6786 34786
rect 6786 34734 6788 34786
rect 6732 34732 6788 34734
rect 6892 34786 6948 34788
rect 6892 34734 6894 34786
rect 6894 34734 6946 34786
rect 6946 34734 6948 34786
rect 6892 34732 6948 34734
rect 7052 34786 7108 34788
rect 7052 34734 7054 34786
rect 7054 34734 7106 34786
rect 7106 34734 7108 34786
rect 7052 34732 7108 34734
rect 7212 34786 7268 34788
rect 7212 34734 7214 34786
rect 7214 34734 7266 34786
rect 7266 34734 7268 34786
rect 7212 34732 7268 34734
rect 7372 34786 7428 34788
rect 7372 34734 7374 34786
rect 7374 34734 7426 34786
rect 7426 34734 7428 34786
rect 7372 34732 7428 34734
rect 7532 34786 7588 34788
rect 7532 34734 7534 34786
rect 7534 34734 7586 34786
rect 7586 34734 7588 34786
rect 7532 34732 7588 34734
rect 7692 34786 7748 34788
rect 7692 34734 7694 34786
rect 7694 34734 7746 34786
rect 7746 34734 7748 34786
rect 7692 34732 7748 34734
rect 7852 34786 7908 34788
rect 7852 34734 7854 34786
rect 7854 34734 7906 34786
rect 7906 34734 7908 34786
rect 7852 34732 7908 34734
rect 8012 34786 8068 34788
rect 8012 34734 8014 34786
rect 8014 34734 8066 34786
rect 8066 34734 8068 34786
rect 8012 34732 8068 34734
rect 8172 34786 8228 34788
rect 8172 34734 8174 34786
rect 8174 34734 8226 34786
rect 8226 34734 8228 34786
rect 8172 34732 8228 34734
rect 8332 34786 8388 34788
rect 8332 34734 8334 34786
rect 8334 34734 8386 34786
rect 8386 34734 8388 34786
rect 8332 34732 8388 34734
rect 9452 34732 9508 34788
rect 9772 34732 9828 34788
rect 10092 34732 10148 34788
rect 10412 34732 10468 34788
rect 10732 34732 10788 34788
rect 11052 34732 11108 34788
rect 11372 34732 11428 34788
rect 12492 34786 12548 34788
rect 12492 34734 12494 34786
rect 12494 34734 12546 34786
rect 12546 34734 12548 34786
rect 12492 34732 12548 34734
rect 12652 34786 12708 34788
rect 12652 34734 12654 34786
rect 12654 34734 12706 34786
rect 12706 34734 12708 34786
rect 12652 34732 12708 34734
rect 12812 34786 12868 34788
rect 12812 34734 12814 34786
rect 12814 34734 12866 34786
rect 12866 34734 12868 34786
rect 12812 34732 12868 34734
rect 12972 34786 13028 34788
rect 12972 34734 12974 34786
rect 12974 34734 13026 34786
rect 13026 34734 13028 34786
rect 12972 34732 13028 34734
rect 13132 34786 13188 34788
rect 13132 34734 13134 34786
rect 13134 34734 13186 34786
rect 13186 34734 13188 34786
rect 13132 34732 13188 34734
rect 13292 34786 13348 34788
rect 13292 34734 13294 34786
rect 13294 34734 13346 34786
rect 13346 34734 13348 34786
rect 13292 34732 13348 34734
rect 13452 34786 13508 34788
rect 13452 34734 13454 34786
rect 13454 34734 13506 34786
rect 13506 34734 13508 34786
rect 13452 34732 13508 34734
rect 13612 34786 13668 34788
rect 13612 34734 13614 34786
rect 13614 34734 13666 34786
rect 13666 34734 13668 34786
rect 13612 34732 13668 34734
rect 13772 34786 13828 34788
rect 13772 34734 13774 34786
rect 13774 34734 13826 34786
rect 13826 34734 13828 34786
rect 13772 34732 13828 34734
rect 13932 34786 13988 34788
rect 13932 34734 13934 34786
rect 13934 34734 13986 34786
rect 13986 34734 13988 34786
rect 13932 34732 13988 34734
rect 14092 34786 14148 34788
rect 14092 34734 14094 34786
rect 14094 34734 14146 34786
rect 14146 34734 14148 34786
rect 14092 34732 14148 34734
rect 14252 34786 14308 34788
rect 14252 34734 14254 34786
rect 14254 34734 14306 34786
rect 14306 34734 14308 34786
rect 14252 34732 14308 34734
rect 14412 34786 14468 34788
rect 14412 34734 14414 34786
rect 14414 34734 14466 34786
rect 14466 34734 14468 34786
rect 14412 34732 14468 34734
rect 14572 34786 14628 34788
rect 14572 34734 14574 34786
rect 14574 34734 14626 34786
rect 14626 34734 14628 34786
rect 14572 34732 14628 34734
rect 14732 34786 14788 34788
rect 14732 34734 14734 34786
rect 14734 34734 14786 34786
rect 14786 34734 14788 34786
rect 14732 34732 14788 34734
rect 14892 34786 14948 34788
rect 14892 34734 14894 34786
rect 14894 34734 14946 34786
rect 14946 34734 14948 34786
rect 14892 34732 14948 34734
rect 15052 34786 15108 34788
rect 15052 34734 15054 34786
rect 15054 34734 15106 34786
rect 15106 34734 15108 34786
rect 15052 34732 15108 34734
rect 15212 34786 15268 34788
rect 15212 34734 15214 34786
rect 15214 34734 15266 34786
rect 15266 34734 15268 34786
rect 15212 34732 15268 34734
rect 15372 34786 15428 34788
rect 15372 34734 15374 34786
rect 15374 34734 15426 34786
rect 15426 34734 15428 34786
rect 15372 34732 15428 34734
rect 15532 34786 15588 34788
rect 15532 34734 15534 34786
rect 15534 34734 15586 34786
rect 15586 34734 15588 34786
rect 15532 34732 15588 34734
rect 15692 34786 15748 34788
rect 15692 34734 15694 34786
rect 15694 34734 15746 34786
rect 15746 34734 15748 34786
rect 15692 34732 15748 34734
rect 15852 34786 15908 34788
rect 15852 34734 15854 34786
rect 15854 34734 15906 34786
rect 15906 34734 15908 34786
rect 15852 34732 15908 34734
rect 16012 34786 16068 34788
rect 16012 34734 16014 34786
rect 16014 34734 16066 34786
rect 16066 34734 16068 34786
rect 16012 34732 16068 34734
rect 16172 34786 16228 34788
rect 16172 34734 16174 34786
rect 16174 34734 16226 34786
rect 16226 34734 16228 34786
rect 16172 34732 16228 34734
rect 16332 34786 16388 34788
rect 16332 34734 16334 34786
rect 16334 34734 16386 34786
rect 16386 34734 16388 34786
rect 16332 34732 16388 34734
rect 16492 34786 16548 34788
rect 16492 34734 16494 34786
rect 16494 34734 16546 34786
rect 16546 34734 16548 34786
rect 16492 34732 16548 34734
rect 16652 34786 16708 34788
rect 16652 34734 16654 34786
rect 16654 34734 16706 34786
rect 16706 34734 16708 34786
rect 16652 34732 16708 34734
rect 16812 34786 16868 34788
rect 16812 34734 16814 34786
rect 16814 34734 16866 34786
rect 16866 34734 16868 34786
rect 16812 34732 16868 34734
rect 16972 34786 17028 34788
rect 16972 34734 16974 34786
rect 16974 34734 17026 34786
rect 17026 34734 17028 34786
rect 16972 34732 17028 34734
rect 17132 34786 17188 34788
rect 17132 34734 17134 34786
rect 17134 34734 17186 34786
rect 17186 34734 17188 34786
rect 17132 34732 17188 34734
rect 17292 34786 17348 34788
rect 17292 34734 17294 34786
rect 17294 34734 17346 34786
rect 17346 34734 17348 34786
rect 17292 34732 17348 34734
rect 17452 34786 17508 34788
rect 17452 34734 17454 34786
rect 17454 34734 17506 34786
rect 17506 34734 17508 34786
rect 17452 34732 17508 34734
rect 17612 34786 17668 34788
rect 17612 34734 17614 34786
rect 17614 34734 17666 34786
rect 17666 34734 17668 34786
rect 17612 34732 17668 34734
rect 17772 34786 17828 34788
rect 17772 34734 17774 34786
rect 17774 34734 17826 34786
rect 17826 34734 17828 34786
rect 17772 34732 17828 34734
rect 17932 34786 17988 34788
rect 17932 34734 17934 34786
rect 17934 34734 17986 34786
rect 17986 34734 17988 34786
rect 17932 34732 17988 34734
rect 18092 34786 18148 34788
rect 18092 34734 18094 34786
rect 18094 34734 18146 34786
rect 18146 34734 18148 34786
rect 18092 34732 18148 34734
rect 18252 34786 18308 34788
rect 18252 34734 18254 34786
rect 18254 34734 18306 34786
rect 18306 34734 18308 34786
rect 18252 34732 18308 34734
rect 18412 34786 18468 34788
rect 18412 34734 18414 34786
rect 18414 34734 18466 34786
rect 18466 34734 18468 34786
rect 18412 34732 18468 34734
rect 18572 34786 18628 34788
rect 18572 34734 18574 34786
rect 18574 34734 18626 34786
rect 18626 34734 18628 34786
rect 18572 34732 18628 34734
rect 18732 34786 18788 34788
rect 18732 34734 18734 34786
rect 18734 34734 18786 34786
rect 18786 34734 18788 34786
rect 18732 34732 18788 34734
rect 18892 34786 18948 34788
rect 18892 34734 18894 34786
rect 18894 34734 18946 34786
rect 18946 34734 18948 34786
rect 18892 34732 18948 34734
rect 20012 34732 20068 34788
rect 20332 34732 20388 34788
rect 20652 34732 20708 34788
rect 20972 34732 21028 34788
rect 21292 34732 21348 34788
rect 21612 34732 21668 34788
rect 21932 34732 21988 34788
rect 23132 34786 23188 34788
rect 23132 34734 23134 34786
rect 23134 34734 23186 34786
rect 23186 34734 23188 34786
rect 23132 34732 23188 34734
rect 23292 34786 23348 34788
rect 23292 34734 23294 34786
rect 23294 34734 23346 34786
rect 23346 34734 23348 34786
rect 23292 34732 23348 34734
rect 23452 34786 23508 34788
rect 23452 34734 23454 34786
rect 23454 34734 23506 34786
rect 23506 34734 23508 34786
rect 23452 34732 23508 34734
rect 23612 34786 23668 34788
rect 23612 34734 23614 34786
rect 23614 34734 23666 34786
rect 23666 34734 23668 34786
rect 23612 34732 23668 34734
rect 23772 34786 23828 34788
rect 23772 34734 23774 34786
rect 23774 34734 23826 34786
rect 23826 34734 23828 34786
rect 23772 34732 23828 34734
rect 23932 34786 23988 34788
rect 23932 34734 23934 34786
rect 23934 34734 23986 34786
rect 23986 34734 23988 34786
rect 23932 34732 23988 34734
rect 24092 34786 24148 34788
rect 24092 34734 24094 34786
rect 24094 34734 24146 34786
rect 24146 34734 24148 34786
rect 24092 34732 24148 34734
rect 24252 34786 24308 34788
rect 24252 34734 24254 34786
rect 24254 34734 24306 34786
rect 24306 34734 24308 34786
rect 24252 34732 24308 34734
rect 24412 34786 24468 34788
rect 24412 34734 24414 34786
rect 24414 34734 24466 34786
rect 24466 34734 24468 34786
rect 24412 34732 24468 34734
rect 24572 34786 24628 34788
rect 24572 34734 24574 34786
rect 24574 34734 24626 34786
rect 24626 34734 24628 34786
rect 24572 34732 24628 34734
rect 24732 34786 24788 34788
rect 24732 34734 24734 34786
rect 24734 34734 24786 34786
rect 24786 34734 24788 34786
rect 24732 34732 24788 34734
rect 24892 34786 24948 34788
rect 24892 34734 24894 34786
rect 24894 34734 24946 34786
rect 24946 34734 24948 34786
rect 24892 34732 24948 34734
rect 25052 34786 25108 34788
rect 25052 34734 25054 34786
rect 25054 34734 25106 34786
rect 25106 34734 25108 34786
rect 25052 34732 25108 34734
rect 25212 34786 25268 34788
rect 25212 34734 25214 34786
rect 25214 34734 25266 34786
rect 25266 34734 25268 34786
rect 25212 34732 25268 34734
rect 25372 34786 25428 34788
rect 25372 34734 25374 34786
rect 25374 34734 25426 34786
rect 25426 34734 25428 34786
rect 25372 34732 25428 34734
rect 25532 34786 25588 34788
rect 25532 34734 25534 34786
rect 25534 34734 25586 34786
rect 25586 34734 25588 34786
rect 25532 34732 25588 34734
rect 25692 34786 25748 34788
rect 25692 34734 25694 34786
rect 25694 34734 25746 34786
rect 25746 34734 25748 34786
rect 25692 34732 25748 34734
rect 25852 34786 25908 34788
rect 25852 34734 25854 34786
rect 25854 34734 25906 34786
rect 25906 34734 25908 34786
rect 25852 34732 25908 34734
rect 26012 34786 26068 34788
rect 26012 34734 26014 34786
rect 26014 34734 26066 34786
rect 26066 34734 26068 34786
rect 26012 34732 26068 34734
rect 26172 34786 26228 34788
rect 26172 34734 26174 34786
rect 26174 34734 26226 34786
rect 26226 34734 26228 34786
rect 26172 34732 26228 34734
rect 26332 34786 26388 34788
rect 26332 34734 26334 34786
rect 26334 34734 26386 34786
rect 26386 34734 26388 34786
rect 26332 34732 26388 34734
rect 26492 34786 26548 34788
rect 26492 34734 26494 34786
rect 26494 34734 26546 34786
rect 26546 34734 26548 34786
rect 26492 34732 26548 34734
rect 26652 34786 26708 34788
rect 26652 34734 26654 34786
rect 26654 34734 26706 34786
rect 26706 34734 26708 34786
rect 26652 34732 26708 34734
rect 26812 34786 26868 34788
rect 26812 34734 26814 34786
rect 26814 34734 26866 34786
rect 26866 34734 26868 34786
rect 26812 34732 26868 34734
rect 26972 34786 27028 34788
rect 26972 34734 26974 34786
rect 26974 34734 27026 34786
rect 27026 34734 27028 34786
rect 26972 34732 27028 34734
rect 27132 34786 27188 34788
rect 27132 34734 27134 34786
rect 27134 34734 27186 34786
rect 27186 34734 27188 34786
rect 27132 34732 27188 34734
rect 27292 34786 27348 34788
rect 27292 34734 27294 34786
rect 27294 34734 27346 34786
rect 27346 34734 27348 34786
rect 27292 34732 27348 34734
rect 27452 34786 27508 34788
rect 27452 34734 27454 34786
rect 27454 34734 27506 34786
rect 27506 34734 27508 34786
rect 27452 34732 27508 34734
rect 27612 34786 27668 34788
rect 27612 34734 27614 34786
rect 27614 34734 27666 34786
rect 27666 34734 27668 34786
rect 27612 34732 27668 34734
rect 27772 34786 27828 34788
rect 27772 34734 27774 34786
rect 27774 34734 27826 34786
rect 27826 34734 27828 34786
rect 27772 34732 27828 34734
rect 27932 34786 27988 34788
rect 27932 34734 27934 34786
rect 27934 34734 27986 34786
rect 27986 34734 27988 34786
rect 27932 34732 27988 34734
rect 28092 34786 28148 34788
rect 28092 34734 28094 34786
rect 28094 34734 28146 34786
rect 28146 34734 28148 34786
rect 28092 34732 28148 34734
rect 28252 34786 28308 34788
rect 28252 34734 28254 34786
rect 28254 34734 28306 34786
rect 28306 34734 28308 34786
rect 28252 34732 28308 34734
rect 28412 34786 28468 34788
rect 28412 34734 28414 34786
rect 28414 34734 28466 34786
rect 28466 34734 28468 34786
rect 28412 34732 28468 34734
rect 28572 34786 28628 34788
rect 28572 34734 28574 34786
rect 28574 34734 28626 34786
rect 28626 34734 28628 34786
rect 28572 34732 28628 34734
rect 28732 34786 28788 34788
rect 28732 34734 28734 34786
rect 28734 34734 28786 34786
rect 28786 34734 28788 34786
rect 28732 34732 28788 34734
rect 28892 34786 28948 34788
rect 28892 34734 28894 34786
rect 28894 34734 28946 34786
rect 28946 34734 28948 34786
rect 28892 34732 28948 34734
rect 29052 34786 29108 34788
rect 29052 34734 29054 34786
rect 29054 34734 29106 34786
rect 29106 34734 29108 34786
rect 29052 34732 29108 34734
rect 29212 34786 29268 34788
rect 29212 34734 29214 34786
rect 29214 34734 29266 34786
rect 29266 34734 29268 34786
rect 29212 34732 29268 34734
rect 29372 34786 29428 34788
rect 29372 34734 29374 34786
rect 29374 34734 29426 34786
rect 29426 34734 29428 34786
rect 29372 34732 29428 34734
rect 30492 34732 30548 34788
rect 30812 34732 30868 34788
rect 31132 34732 31188 34788
rect 31452 34732 31508 34788
rect 31772 34732 31828 34788
rect 32092 34732 32148 34788
rect 32412 34732 32468 34788
rect 33532 34786 33588 34788
rect 33532 34734 33534 34786
rect 33534 34734 33586 34786
rect 33586 34734 33588 34786
rect 33532 34732 33588 34734
rect 33692 34786 33748 34788
rect 33692 34734 33694 34786
rect 33694 34734 33746 34786
rect 33746 34734 33748 34786
rect 33692 34732 33748 34734
rect 33852 34786 33908 34788
rect 33852 34734 33854 34786
rect 33854 34734 33906 34786
rect 33906 34734 33908 34786
rect 33852 34732 33908 34734
rect 34012 34786 34068 34788
rect 34012 34734 34014 34786
rect 34014 34734 34066 34786
rect 34066 34734 34068 34786
rect 34012 34732 34068 34734
rect 34172 34786 34228 34788
rect 34172 34734 34174 34786
rect 34174 34734 34226 34786
rect 34226 34734 34228 34786
rect 34172 34732 34228 34734
rect 34332 34786 34388 34788
rect 34332 34734 34334 34786
rect 34334 34734 34386 34786
rect 34386 34734 34388 34786
rect 34332 34732 34388 34734
rect 34492 34786 34548 34788
rect 34492 34734 34494 34786
rect 34494 34734 34546 34786
rect 34546 34734 34548 34786
rect 34492 34732 34548 34734
rect 34652 34786 34708 34788
rect 34652 34734 34654 34786
rect 34654 34734 34706 34786
rect 34706 34734 34708 34786
rect 34652 34732 34708 34734
rect 34812 34786 34868 34788
rect 34812 34734 34814 34786
rect 34814 34734 34866 34786
rect 34866 34734 34868 34786
rect 34812 34732 34868 34734
rect 34972 34786 35028 34788
rect 34972 34734 34974 34786
rect 34974 34734 35026 34786
rect 35026 34734 35028 34786
rect 34972 34732 35028 34734
rect 35132 34786 35188 34788
rect 35132 34734 35134 34786
rect 35134 34734 35186 34786
rect 35186 34734 35188 34786
rect 35132 34732 35188 34734
rect 35292 34786 35348 34788
rect 35292 34734 35294 34786
rect 35294 34734 35346 34786
rect 35346 34734 35348 34786
rect 35292 34732 35348 34734
rect 35452 34786 35508 34788
rect 35452 34734 35454 34786
rect 35454 34734 35506 34786
rect 35506 34734 35508 34786
rect 35452 34732 35508 34734
rect 35612 34786 35668 34788
rect 35612 34734 35614 34786
rect 35614 34734 35666 34786
rect 35666 34734 35668 34786
rect 35612 34732 35668 34734
rect 35772 34786 35828 34788
rect 35772 34734 35774 34786
rect 35774 34734 35826 34786
rect 35826 34734 35828 34786
rect 35772 34732 35828 34734
rect 35932 34786 35988 34788
rect 35932 34734 35934 34786
rect 35934 34734 35986 34786
rect 35986 34734 35988 34786
rect 35932 34732 35988 34734
rect 36092 34786 36148 34788
rect 36092 34734 36094 34786
rect 36094 34734 36146 34786
rect 36146 34734 36148 34786
rect 36092 34732 36148 34734
rect 36252 34786 36308 34788
rect 36252 34734 36254 34786
rect 36254 34734 36306 34786
rect 36306 34734 36308 34786
rect 36252 34732 36308 34734
rect 36412 34786 36468 34788
rect 36412 34734 36414 34786
rect 36414 34734 36466 34786
rect 36466 34734 36468 34786
rect 36412 34732 36468 34734
rect 36572 34786 36628 34788
rect 36572 34734 36574 34786
rect 36574 34734 36626 34786
rect 36626 34734 36628 34786
rect 36572 34732 36628 34734
rect 36732 34786 36788 34788
rect 36732 34734 36734 34786
rect 36734 34734 36786 34786
rect 36786 34734 36788 34786
rect 36732 34732 36788 34734
rect 36892 34786 36948 34788
rect 36892 34734 36894 34786
rect 36894 34734 36946 34786
rect 36946 34734 36948 34786
rect 36892 34732 36948 34734
rect 37052 34786 37108 34788
rect 37052 34734 37054 34786
rect 37054 34734 37106 34786
rect 37106 34734 37108 34786
rect 37052 34732 37108 34734
rect 37212 34786 37268 34788
rect 37212 34734 37214 34786
rect 37214 34734 37266 34786
rect 37266 34734 37268 34786
rect 37212 34732 37268 34734
rect 37372 34786 37428 34788
rect 37372 34734 37374 34786
rect 37374 34734 37426 34786
rect 37426 34734 37428 34786
rect 37372 34732 37428 34734
rect 37532 34786 37588 34788
rect 37532 34734 37534 34786
rect 37534 34734 37586 34786
rect 37586 34734 37588 34786
rect 37532 34732 37588 34734
rect 37692 34786 37748 34788
rect 37692 34734 37694 34786
rect 37694 34734 37746 34786
rect 37746 34734 37748 34786
rect 37692 34732 37748 34734
rect 37852 34786 37908 34788
rect 37852 34734 37854 34786
rect 37854 34734 37906 34786
rect 37906 34734 37908 34786
rect 37852 34732 37908 34734
rect 38012 34786 38068 34788
rect 38012 34734 38014 34786
rect 38014 34734 38066 34786
rect 38066 34734 38068 34786
rect 38012 34732 38068 34734
rect 38172 34786 38228 34788
rect 38172 34734 38174 34786
rect 38174 34734 38226 34786
rect 38226 34734 38228 34786
rect 38172 34732 38228 34734
rect 38332 34786 38388 34788
rect 38332 34734 38334 34786
rect 38334 34734 38386 34786
rect 38386 34734 38388 34786
rect 38332 34732 38388 34734
rect 38492 34786 38548 34788
rect 38492 34734 38494 34786
rect 38494 34734 38546 34786
rect 38546 34734 38548 34786
rect 38492 34732 38548 34734
rect 38652 34786 38708 34788
rect 38652 34734 38654 34786
rect 38654 34734 38706 34786
rect 38706 34734 38708 34786
rect 38652 34732 38708 34734
rect 38812 34786 38868 34788
rect 38812 34734 38814 34786
rect 38814 34734 38866 34786
rect 38866 34734 38868 34786
rect 38812 34732 38868 34734
rect 38972 34786 39028 34788
rect 38972 34734 38974 34786
rect 38974 34734 39026 34786
rect 39026 34734 39028 34786
rect 38972 34732 39028 34734
rect 39132 34786 39188 34788
rect 39132 34734 39134 34786
rect 39134 34734 39186 34786
rect 39186 34734 39188 34786
rect 39132 34732 39188 34734
rect 39292 34786 39348 34788
rect 39292 34734 39294 34786
rect 39294 34734 39346 34786
rect 39346 34734 39348 34786
rect 39292 34732 39348 34734
rect 39452 34786 39508 34788
rect 39452 34734 39454 34786
rect 39454 34734 39506 34786
rect 39506 34734 39508 34786
rect 39452 34732 39508 34734
rect 39612 34786 39668 34788
rect 39612 34734 39614 34786
rect 39614 34734 39666 34786
rect 39666 34734 39668 34786
rect 39612 34732 39668 34734
rect 39772 34786 39828 34788
rect 39772 34734 39774 34786
rect 39774 34734 39826 34786
rect 39826 34734 39828 34786
rect 39772 34732 39828 34734
rect 39932 34786 39988 34788
rect 39932 34734 39934 34786
rect 39934 34734 39986 34786
rect 39986 34734 39988 34786
rect 39932 34732 39988 34734
rect 40092 34786 40148 34788
rect 40092 34734 40094 34786
rect 40094 34734 40146 34786
rect 40146 34734 40148 34786
rect 40092 34732 40148 34734
rect 40252 34786 40308 34788
rect 40252 34734 40254 34786
rect 40254 34734 40306 34786
rect 40306 34734 40308 34786
rect 40252 34732 40308 34734
rect 40412 34786 40468 34788
rect 40412 34734 40414 34786
rect 40414 34734 40466 34786
rect 40466 34734 40468 34786
rect 40412 34732 40468 34734
rect 40572 34786 40628 34788
rect 40572 34734 40574 34786
rect 40574 34734 40626 34786
rect 40626 34734 40628 34786
rect 40572 34732 40628 34734
rect 40732 34786 40788 34788
rect 40732 34734 40734 34786
rect 40734 34734 40786 34786
rect 40786 34734 40788 34786
rect 40732 34732 40788 34734
rect 40892 34786 40948 34788
rect 40892 34734 40894 34786
rect 40894 34734 40946 34786
rect 40946 34734 40948 34786
rect 40892 34732 40948 34734
rect 41052 34786 41108 34788
rect 41052 34734 41054 34786
rect 41054 34734 41106 34786
rect 41106 34734 41108 34786
rect 41052 34732 41108 34734
rect 41212 34786 41268 34788
rect 41212 34734 41214 34786
rect 41214 34734 41266 34786
rect 41266 34734 41268 34786
rect 41212 34732 41268 34734
rect 41372 34786 41428 34788
rect 41372 34734 41374 34786
rect 41374 34734 41426 34786
rect 41426 34734 41428 34786
rect 41372 34732 41428 34734
rect 41532 34786 41588 34788
rect 41532 34734 41534 34786
rect 41534 34734 41586 34786
rect 41586 34734 41588 34786
rect 41532 34732 41588 34734
rect 41692 34786 41748 34788
rect 41692 34734 41694 34786
rect 41694 34734 41746 34786
rect 41746 34734 41748 34786
rect 41692 34732 41748 34734
rect 41852 34786 41908 34788
rect 41852 34734 41854 34786
rect 41854 34734 41906 34786
rect 41906 34734 41908 34786
rect 41852 34732 41908 34734
rect 11212 34572 11268 34628
rect 20172 34572 20228 34628
rect 30652 34572 30708 34628
rect 12 34466 68 34468
rect 12 34414 14 34466
rect 14 34414 66 34466
rect 66 34414 68 34466
rect 12 34412 68 34414
rect 172 34466 228 34468
rect 172 34414 174 34466
rect 174 34414 226 34466
rect 226 34414 228 34466
rect 172 34412 228 34414
rect 332 34466 388 34468
rect 332 34414 334 34466
rect 334 34414 386 34466
rect 386 34414 388 34466
rect 332 34412 388 34414
rect 492 34466 548 34468
rect 492 34414 494 34466
rect 494 34414 546 34466
rect 546 34414 548 34466
rect 492 34412 548 34414
rect 652 34466 708 34468
rect 652 34414 654 34466
rect 654 34414 706 34466
rect 706 34414 708 34466
rect 652 34412 708 34414
rect 812 34466 868 34468
rect 812 34414 814 34466
rect 814 34414 866 34466
rect 866 34414 868 34466
rect 812 34412 868 34414
rect 972 34466 1028 34468
rect 972 34414 974 34466
rect 974 34414 1026 34466
rect 1026 34414 1028 34466
rect 972 34412 1028 34414
rect 1132 34466 1188 34468
rect 1132 34414 1134 34466
rect 1134 34414 1186 34466
rect 1186 34414 1188 34466
rect 1132 34412 1188 34414
rect 1292 34466 1348 34468
rect 1292 34414 1294 34466
rect 1294 34414 1346 34466
rect 1346 34414 1348 34466
rect 1292 34412 1348 34414
rect 1452 34466 1508 34468
rect 1452 34414 1454 34466
rect 1454 34414 1506 34466
rect 1506 34414 1508 34466
rect 1452 34412 1508 34414
rect 1612 34466 1668 34468
rect 1612 34414 1614 34466
rect 1614 34414 1666 34466
rect 1666 34414 1668 34466
rect 1612 34412 1668 34414
rect 1772 34466 1828 34468
rect 1772 34414 1774 34466
rect 1774 34414 1826 34466
rect 1826 34414 1828 34466
rect 1772 34412 1828 34414
rect 1932 34466 1988 34468
rect 1932 34414 1934 34466
rect 1934 34414 1986 34466
rect 1986 34414 1988 34466
rect 1932 34412 1988 34414
rect 2092 34466 2148 34468
rect 2092 34414 2094 34466
rect 2094 34414 2146 34466
rect 2146 34414 2148 34466
rect 2092 34412 2148 34414
rect 2252 34466 2308 34468
rect 2252 34414 2254 34466
rect 2254 34414 2306 34466
rect 2306 34414 2308 34466
rect 2252 34412 2308 34414
rect 2412 34466 2468 34468
rect 2412 34414 2414 34466
rect 2414 34414 2466 34466
rect 2466 34414 2468 34466
rect 2412 34412 2468 34414
rect 2572 34466 2628 34468
rect 2572 34414 2574 34466
rect 2574 34414 2626 34466
rect 2626 34414 2628 34466
rect 2572 34412 2628 34414
rect 2732 34466 2788 34468
rect 2732 34414 2734 34466
rect 2734 34414 2786 34466
rect 2786 34414 2788 34466
rect 2732 34412 2788 34414
rect 2892 34466 2948 34468
rect 2892 34414 2894 34466
rect 2894 34414 2946 34466
rect 2946 34414 2948 34466
rect 2892 34412 2948 34414
rect 3052 34466 3108 34468
rect 3052 34414 3054 34466
rect 3054 34414 3106 34466
rect 3106 34414 3108 34466
rect 3052 34412 3108 34414
rect 3212 34466 3268 34468
rect 3212 34414 3214 34466
rect 3214 34414 3266 34466
rect 3266 34414 3268 34466
rect 3212 34412 3268 34414
rect 3372 34466 3428 34468
rect 3372 34414 3374 34466
rect 3374 34414 3426 34466
rect 3426 34414 3428 34466
rect 3372 34412 3428 34414
rect 3532 34466 3588 34468
rect 3532 34414 3534 34466
rect 3534 34414 3586 34466
rect 3586 34414 3588 34466
rect 3532 34412 3588 34414
rect 3692 34466 3748 34468
rect 3692 34414 3694 34466
rect 3694 34414 3746 34466
rect 3746 34414 3748 34466
rect 3692 34412 3748 34414
rect 3852 34466 3908 34468
rect 3852 34414 3854 34466
rect 3854 34414 3906 34466
rect 3906 34414 3908 34466
rect 3852 34412 3908 34414
rect 4012 34466 4068 34468
rect 4012 34414 4014 34466
rect 4014 34414 4066 34466
rect 4066 34414 4068 34466
rect 4012 34412 4068 34414
rect 4172 34466 4228 34468
rect 4172 34414 4174 34466
rect 4174 34414 4226 34466
rect 4226 34414 4228 34466
rect 4172 34412 4228 34414
rect 4332 34466 4388 34468
rect 4332 34414 4334 34466
rect 4334 34414 4386 34466
rect 4386 34414 4388 34466
rect 4332 34412 4388 34414
rect 4492 34466 4548 34468
rect 4492 34414 4494 34466
rect 4494 34414 4546 34466
rect 4546 34414 4548 34466
rect 4492 34412 4548 34414
rect 4652 34466 4708 34468
rect 4652 34414 4654 34466
rect 4654 34414 4706 34466
rect 4706 34414 4708 34466
rect 4652 34412 4708 34414
rect 4812 34466 4868 34468
rect 4812 34414 4814 34466
rect 4814 34414 4866 34466
rect 4866 34414 4868 34466
rect 4812 34412 4868 34414
rect 4972 34466 5028 34468
rect 4972 34414 4974 34466
rect 4974 34414 5026 34466
rect 5026 34414 5028 34466
rect 4972 34412 5028 34414
rect 5132 34466 5188 34468
rect 5132 34414 5134 34466
rect 5134 34414 5186 34466
rect 5186 34414 5188 34466
rect 5132 34412 5188 34414
rect 5292 34466 5348 34468
rect 5292 34414 5294 34466
rect 5294 34414 5346 34466
rect 5346 34414 5348 34466
rect 5292 34412 5348 34414
rect 5452 34466 5508 34468
rect 5452 34414 5454 34466
rect 5454 34414 5506 34466
rect 5506 34414 5508 34466
rect 5452 34412 5508 34414
rect 5612 34466 5668 34468
rect 5612 34414 5614 34466
rect 5614 34414 5666 34466
rect 5666 34414 5668 34466
rect 5612 34412 5668 34414
rect 5772 34466 5828 34468
rect 5772 34414 5774 34466
rect 5774 34414 5826 34466
rect 5826 34414 5828 34466
rect 5772 34412 5828 34414
rect 5932 34466 5988 34468
rect 5932 34414 5934 34466
rect 5934 34414 5986 34466
rect 5986 34414 5988 34466
rect 5932 34412 5988 34414
rect 6092 34466 6148 34468
rect 6092 34414 6094 34466
rect 6094 34414 6146 34466
rect 6146 34414 6148 34466
rect 6092 34412 6148 34414
rect 6252 34466 6308 34468
rect 6252 34414 6254 34466
rect 6254 34414 6306 34466
rect 6306 34414 6308 34466
rect 6252 34412 6308 34414
rect 6412 34466 6468 34468
rect 6412 34414 6414 34466
rect 6414 34414 6466 34466
rect 6466 34414 6468 34466
rect 6412 34412 6468 34414
rect 6572 34466 6628 34468
rect 6572 34414 6574 34466
rect 6574 34414 6626 34466
rect 6626 34414 6628 34466
rect 6572 34412 6628 34414
rect 6732 34466 6788 34468
rect 6732 34414 6734 34466
rect 6734 34414 6786 34466
rect 6786 34414 6788 34466
rect 6732 34412 6788 34414
rect 6892 34466 6948 34468
rect 6892 34414 6894 34466
rect 6894 34414 6946 34466
rect 6946 34414 6948 34466
rect 6892 34412 6948 34414
rect 7052 34466 7108 34468
rect 7052 34414 7054 34466
rect 7054 34414 7106 34466
rect 7106 34414 7108 34466
rect 7052 34412 7108 34414
rect 7212 34466 7268 34468
rect 7212 34414 7214 34466
rect 7214 34414 7266 34466
rect 7266 34414 7268 34466
rect 7212 34412 7268 34414
rect 7372 34466 7428 34468
rect 7372 34414 7374 34466
rect 7374 34414 7426 34466
rect 7426 34414 7428 34466
rect 7372 34412 7428 34414
rect 7532 34466 7588 34468
rect 7532 34414 7534 34466
rect 7534 34414 7586 34466
rect 7586 34414 7588 34466
rect 7532 34412 7588 34414
rect 7692 34466 7748 34468
rect 7692 34414 7694 34466
rect 7694 34414 7746 34466
rect 7746 34414 7748 34466
rect 7692 34412 7748 34414
rect 7852 34466 7908 34468
rect 7852 34414 7854 34466
rect 7854 34414 7906 34466
rect 7906 34414 7908 34466
rect 7852 34412 7908 34414
rect 8012 34466 8068 34468
rect 8012 34414 8014 34466
rect 8014 34414 8066 34466
rect 8066 34414 8068 34466
rect 8012 34412 8068 34414
rect 8172 34466 8228 34468
rect 8172 34414 8174 34466
rect 8174 34414 8226 34466
rect 8226 34414 8228 34466
rect 8172 34412 8228 34414
rect 8332 34466 8388 34468
rect 8332 34414 8334 34466
rect 8334 34414 8386 34466
rect 8386 34414 8388 34466
rect 8332 34412 8388 34414
rect 9452 34412 9508 34468
rect 9772 34412 9828 34468
rect 10092 34412 10148 34468
rect 10412 34412 10468 34468
rect 10732 34412 10788 34468
rect 11052 34412 11108 34468
rect 11372 34412 11428 34468
rect 12492 34466 12548 34468
rect 12492 34414 12494 34466
rect 12494 34414 12546 34466
rect 12546 34414 12548 34466
rect 12492 34412 12548 34414
rect 12652 34466 12708 34468
rect 12652 34414 12654 34466
rect 12654 34414 12706 34466
rect 12706 34414 12708 34466
rect 12652 34412 12708 34414
rect 12812 34466 12868 34468
rect 12812 34414 12814 34466
rect 12814 34414 12866 34466
rect 12866 34414 12868 34466
rect 12812 34412 12868 34414
rect 12972 34466 13028 34468
rect 12972 34414 12974 34466
rect 12974 34414 13026 34466
rect 13026 34414 13028 34466
rect 12972 34412 13028 34414
rect 13132 34466 13188 34468
rect 13132 34414 13134 34466
rect 13134 34414 13186 34466
rect 13186 34414 13188 34466
rect 13132 34412 13188 34414
rect 13292 34466 13348 34468
rect 13292 34414 13294 34466
rect 13294 34414 13346 34466
rect 13346 34414 13348 34466
rect 13292 34412 13348 34414
rect 13452 34466 13508 34468
rect 13452 34414 13454 34466
rect 13454 34414 13506 34466
rect 13506 34414 13508 34466
rect 13452 34412 13508 34414
rect 13612 34466 13668 34468
rect 13612 34414 13614 34466
rect 13614 34414 13666 34466
rect 13666 34414 13668 34466
rect 13612 34412 13668 34414
rect 13772 34466 13828 34468
rect 13772 34414 13774 34466
rect 13774 34414 13826 34466
rect 13826 34414 13828 34466
rect 13772 34412 13828 34414
rect 13932 34466 13988 34468
rect 13932 34414 13934 34466
rect 13934 34414 13986 34466
rect 13986 34414 13988 34466
rect 13932 34412 13988 34414
rect 14092 34466 14148 34468
rect 14092 34414 14094 34466
rect 14094 34414 14146 34466
rect 14146 34414 14148 34466
rect 14092 34412 14148 34414
rect 14252 34466 14308 34468
rect 14252 34414 14254 34466
rect 14254 34414 14306 34466
rect 14306 34414 14308 34466
rect 14252 34412 14308 34414
rect 14412 34466 14468 34468
rect 14412 34414 14414 34466
rect 14414 34414 14466 34466
rect 14466 34414 14468 34466
rect 14412 34412 14468 34414
rect 14572 34466 14628 34468
rect 14572 34414 14574 34466
rect 14574 34414 14626 34466
rect 14626 34414 14628 34466
rect 14572 34412 14628 34414
rect 14732 34466 14788 34468
rect 14732 34414 14734 34466
rect 14734 34414 14786 34466
rect 14786 34414 14788 34466
rect 14732 34412 14788 34414
rect 14892 34466 14948 34468
rect 14892 34414 14894 34466
rect 14894 34414 14946 34466
rect 14946 34414 14948 34466
rect 14892 34412 14948 34414
rect 15052 34466 15108 34468
rect 15052 34414 15054 34466
rect 15054 34414 15106 34466
rect 15106 34414 15108 34466
rect 15052 34412 15108 34414
rect 15212 34466 15268 34468
rect 15212 34414 15214 34466
rect 15214 34414 15266 34466
rect 15266 34414 15268 34466
rect 15212 34412 15268 34414
rect 15372 34466 15428 34468
rect 15372 34414 15374 34466
rect 15374 34414 15426 34466
rect 15426 34414 15428 34466
rect 15372 34412 15428 34414
rect 15532 34466 15588 34468
rect 15532 34414 15534 34466
rect 15534 34414 15586 34466
rect 15586 34414 15588 34466
rect 15532 34412 15588 34414
rect 15692 34466 15748 34468
rect 15692 34414 15694 34466
rect 15694 34414 15746 34466
rect 15746 34414 15748 34466
rect 15692 34412 15748 34414
rect 15852 34466 15908 34468
rect 15852 34414 15854 34466
rect 15854 34414 15906 34466
rect 15906 34414 15908 34466
rect 15852 34412 15908 34414
rect 16012 34466 16068 34468
rect 16012 34414 16014 34466
rect 16014 34414 16066 34466
rect 16066 34414 16068 34466
rect 16012 34412 16068 34414
rect 16172 34466 16228 34468
rect 16172 34414 16174 34466
rect 16174 34414 16226 34466
rect 16226 34414 16228 34466
rect 16172 34412 16228 34414
rect 16332 34466 16388 34468
rect 16332 34414 16334 34466
rect 16334 34414 16386 34466
rect 16386 34414 16388 34466
rect 16332 34412 16388 34414
rect 16492 34466 16548 34468
rect 16492 34414 16494 34466
rect 16494 34414 16546 34466
rect 16546 34414 16548 34466
rect 16492 34412 16548 34414
rect 16652 34466 16708 34468
rect 16652 34414 16654 34466
rect 16654 34414 16706 34466
rect 16706 34414 16708 34466
rect 16652 34412 16708 34414
rect 16812 34466 16868 34468
rect 16812 34414 16814 34466
rect 16814 34414 16866 34466
rect 16866 34414 16868 34466
rect 16812 34412 16868 34414
rect 16972 34466 17028 34468
rect 16972 34414 16974 34466
rect 16974 34414 17026 34466
rect 17026 34414 17028 34466
rect 16972 34412 17028 34414
rect 17132 34466 17188 34468
rect 17132 34414 17134 34466
rect 17134 34414 17186 34466
rect 17186 34414 17188 34466
rect 17132 34412 17188 34414
rect 17292 34466 17348 34468
rect 17292 34414 17294 34466
rect 17294 34414 17346 34466
rect 17346 34414 17348 34466
rect 17292 34412 17348 34414
rect 17452 34466 17508 34468
rect 17452 34414 17454 34466
rect 17454 34414 17506 34466
rect 17506 34414 17508 34466
rect 17452 34412 17508 34414
rect 17612 34466 17668 34468
rect 17612 34414 17614 34466
rect 17614 34414 17666 34466
rect 17666 34414 17668 34466
rect 17612 34412 17668 34414
rect 17772 34466 17828 34468
rect 17772 34414 17774 34466
rect 17774 34414 17826 34466
rect 17826 34414 17828 34466
rect 17772 34412 17828 34414
rect 17932 34466 17988 34468
rect 17932 34414 17934 34466
rect 17934 34414 17986 34466
rect 17986 34414 17988 34466
rect 17932 34412 17988 34414
rect 18092 34466 18148 34468
rect 18092 34414 18094 34466
rect 18094 34414 18146 34466
rect 18146 34414 18148 34466
rect 18092 34412 18148 34414
rect 18252 34466 18308 34468
rect 18252 34414 18254 34466
rect 18254 34414 18306 34466
rect 18306 34414 18308 34466
rect 18252 34412 18308 34414
rect 18412 34466 18468 34468
rect 18412 34414 18414 34466
rect 18414 34414 18466 34466
rect 18466 34414 18468 34466
rect 18412 34412 18468 34414
rect 18572 34466 18628 34468
rect 18572 34414 18574 34466
rect 18574 34414 18626 34466
rect 18626 34414 18628 34466
rect 18572 34412 18628 34414
rect 18732 34466 18788 34468
rect 18732 34414 18734 34466
rect 18734 34414 18786 34466
rect 18786 34414 18788 34466
rect 18732 34412 18788 34414
rect 18892 34466 18948 34468
rect 18892 34414 18894 34466
rect 18894 34414 18946 34466
rect 18946 34414 18948 34466
rect 18892 34412 18948 34414
rect 20012 34412 20068 34468
rect 20332 34412 20388 34468
rect 20652 34412 20708 34468
rect 20972 34412 21028 34468
rect 21292 34412 21348 34468
rect 21612 34412 21668 34468
rect 21932 34412 21988 34468
rect 23132 34466 23188 34468
rect 23132 34414 23134 34466
rect 23134 34414 23186 34466
rect 23186 34414 23188 34466
rect 23132 34412 23188 34414
rect 23292 34466 23348 34468
rect 23292 34414 23294 34466
rect 23294 34414 23346 34466
rect 23346 34414 23348 34466
rect 23292 34412 23348 34414
rect 23452 34466 23508 34468
rect 23452 34414 23454 34466
rect 23454 34414 23506 34466
rect 23506 34414 23508 34466
rect 23452 34412 23508 34414
rect 23612 34466 23668 34468
rect 23612 34414 23614 34466
rect 23614 34414 23666 34466
rect 23666 34414 23668 34466
rect 23612 34412 23668 34414
rect 23772 34466 23828 34468
rect 23772 34414 23774 34466
rect 23774 34414 23826 34466
rect 23826 34414 23828 34466
rect 23772 34412 23828 34414
rect 23932 34466 23988 34468
rect 23932 34414 23934 34466
rect 23934 34414 23986 34466
rect 23986 34414 23988 34466
rect 23932 34412 23988 34414
rect 24092 34466 24148 34468
rect 24092 34414 24094 34466
rect 24094 34414 24146 34466
rect 24146 34414 24148 34466
rect 24092 34412 24148 34414
rect 24252 34466 24308 34468
rect 24252 34414 24254 34466
rect 24254 34414 24306 34466
rect 24306 34414 24308 34466
rect 24252 34412 24308 34414
rect 24412 34466 24468 34468
rect 24412 34414 24414 34466
rect 24414 34414 24466 34466
rect 24466 34414 24468 34466
rect 24412 34412 24468 34414
rect 24572 34466 24628 34468
rect 24572 34414 24574 34466
rect 24574 34414 24626 34466
rect 24626 34414 24628 34466
rect 24572 34412 24628 34414
rect 24732 34466 24788 34468
rect 24732 34414 24734 34466
rect 24734 34414 24786 34466
rect 24786 34414 24788 34466
rect 24732 34412 24788 34414
rect 24892 34466 24948 34468
rect 24892 34414 24894 34466
rect 24894 34414 24946 34466
rect 24946 34414 24948 34466
rect 24892 34412 24948 34414
rect 25052 34466 25108 34468
rect 25052 34414 25054 34466
rect 25054 34414 25106 34466
rect 25106 34414 25108 34466
rect 25052 34412 25108 34414
rect 25212 34466 25268 34468
rect 25212 34414 25214 34466
rect 25214 34414 25266 34466
rect 25266 34414 25268 34466
rect 25212 34412 25268 34414
rect 25372 34466 25428 34468
rect 25372 34414 25374 34466
rect 25374 34414 25426 34466
rect 25426 34414 25428 34466
rect 25372 34412 25428 34414
rect 25532 34466 25588 34468
rect 25532 34414 25534 34466
rect 25534 34414 25586 34466
rect 25586 34414 25588 34466
rect 25532 34412 25588 34414
rect 25692 34466 25748 34468
rect 25692 34414 25694 34466
rect 25694 34414 25746 34466
rect 25746 34414 25748 34466
rect 25692 34412 25748 34414
rect 25852 34466 25908 34468
rect 25852 34414 25854 34466
rect 25854 34414 25906 34466
rect 25906 34414 25908 34466
rect 25852 34412 25908 34414
rect 26012 34466 26068 34468
rect 26012 34414 26014 34466
rect 26014 34414 26066 34466
rect 26066 34414 26068 34466
rect 26012 34412 26068 34414
rect 26172 34466 26228 34468
rect 26172 34414 26174 34466
rect 26174 34414 26226 34466
rect 26226 34414 26228 34466
rect 26172 34412 26228 34414
rect 26332 34466 26388 34468
rect 26332 34414 26334 34466
rect 26334 34414 26386 34466
rect 26386 34414 26388 34466
rect 26332 34412 26388 34414
rect 26492 34466 26548 34468
rect 26492 34414 26494 34466
rect 26494 34414 26546 34466
rect 26546 34414 26548 34466
rect 26492 34412 26548 34414
rect 26652 34466 26708 34468
rect 26652 34414 26654 34466
rect 26654 34414 26706 34466
rect 26706 34414 26708 34466
rect 26652 34412 26708 34414
rect 26812 34466 26868 34468
rect 26812 34414 26814 34466
rect 26814 34414 26866 34466
rect 26866 34414 26868 34466
rect 26812 34412 26868 34414
rect 26972 34466 27028 34468
rect 26972 34414 26974 34466
rect 26974 34414 27026 34466
rect 27026 34414 27028 34466
rect 26972 34412 27028 34414
rect 27132 34466 27188 34468
rect 27132 34414 27134 34466
rect 27134 34414 27186 34466
rect 27186 34414 27188 34466
rect 27132 34412 27188 34414
rect 27292 34466 27348 34468
rect 27292 34414 27294 34466
rect 27294 34414 27346 34466
rect 27346 34414 27348 34466
rect 27292 34412 27348 34414
rect 27452 34466 27508 34468
rect 27452 34414 27454 34466
rect 27454 34414 27506 34466
rect 27506 34414 27508 34466
rect 27452 34412 27508 34414
rect 27612 34466 27668 34468
rect 27612 34414 27614 34466
rect 27614 34414 27666 34466
rect 27666 34414 27668 34466
rect 27612 34412 27668 34414
rect 27772 34466 27828 34468
rect 27772 34414 27774 34466
rect 27774 34414 27826 34466
rect 27826 34414 27828 34466
rect 27772 34412 27828 34414
rect 27932 34466 27988 34468
rect 27932 34414 27934 34466
rect 27934 34414 27986 34466
rect 27986 34414 27988 34466
rect 27932 34412 27988 34414
rect 28092 34466 28148 34468
rect 28092 34414 28094 34466
rect 28094 34414 28146 34466
rect 28146 34414 28148 34466
rect 28092 34412 28148 34414
rect 28252 34466 28308 34468
rect 28252 34414 28254 34466
rect 28254 34414 28306 34466
rect 28306 34414 28308 34466
rect 28252 34412 28308 34414
rect 28412 34466 28468 34468
rect 28412 34414 28414 34466
rect 28414 34414 28466 34466
rect 28466 34414 28468 34466
rect 28412 34412 28468 34414
rect 28572 34466 28628 34468
rect 28572 34414 28574 34466
rect 28574 34414 28626 34466
rect 28626 34414 28628 34466
rect 28572 34412 28628 34414
rect 28732 34466 28788 34468
rect 28732 34414 28734 34466
rect 28734 34414 28786 34466
rect 28786 34414 28788 34466
rect 28732 34412 28788 34414
rect 28892 34466 28948 34468
rect 28892 34414 28894 34466
rect 28894 34414 28946 34466
rect 28946 34414 28948 34466
rect 28892 34412 28948 34414
rect 29052 34466 29108 34468
rect 29052 34414 29054 34466
rect 29054 34414 29106 34466
rect 29106 34414 29108 34466
rect 29052 34412 29108 34414
rect 29212 34466 29268 34468
rect 29212 34414 29214 34466
rect 29214 34414 29266 34466
rect 29266 34414 29268 34466
rect 29212 34412 29268 34414
rect 29372 34466 29428 34468
rect 29372 34414 29374 34466
rect 29374 34414 29426 34466
rect 29426 34414 29428 34466
rect 29372 34412 29428 34414
rect 30492 34412 30548 34468
rect 30812 34412 30868 34468
rect 31132 34412 31188 34468
rect 31452 34412 31508 34468
rect 31772 34412 31828 34468
rect 32092 34412 32148 34468
rect 32412 34412 32468 34468
rect 33532 34466 33588 34468
rect 33532 34414 33534 34466
rect 33534 34414 33586 34466
rect 33586 34414 33588 34466
rect 33532 34412 33588 34414
rect 33692 34466 33748 34468
rect 33692 34414 33694 34466
rect 33694 34414 33746 34466
rect 33746 34414 33748 34466
rect 33692 34412 33748 34414
rect 33852 34466 33908 34468
rect 33852 34414 33854 34466
rect 33854 34414 33906 34466
rect 33906 34414 33908 34466
rect 33852 34412 33908 34414
rect 34012 34466 34068 34468
rect 34012 34414 34014 34466
rect 34014 34414 34066 34466
rect 34066 34414 34068 34466
rect 34012 34412 34068 34414
rect 34172 34466 34228 34468
rect 34172 34414 34174 34466
rect 34174 34414 34226 34466
rect 34226 34414 34228 34466
rect 34172 34412 34228 34414
rect 34332 34466 34388 34468
rect 34332 34414 34334 34466
rect 34334 34414 34386 34466
rect 34386 34414 34388 34466
rect 34332 34412 34388 34414
rect 34492 34466 34548 34468
rect 34492 34414 34494 34466
rect 34494 34414 34546 34466
rect 34546 34414 34548 34466
rect 34492 34412 34548 34414
rect 34652 34466 34708 34468
rect 34652 34414 34654 34466
rect 34654 34414 34706 34466
rect 34706 34414 34708 34466
rect 34652 34412 34708 34414
rect 34812 34466 34868 34468
rect 34812 34414 34814 34466
rect 34814 34414 34866 34466
rect 34866 34414 34868 34466
rect 34812 34412 34868 34414
rect 34972 34466 35028 34468
rect 34972 34414 34974 34466
rect 34974 34414 35026 34466
rect 35026 34414 35028 34466
rect 34972 34412 35028 34414
rect 35132 34466 35188 34468
rect 35132 34414 35134 34466
rect 35134 34414 35186 34466
rect 35186 34414 35188 34466
rect 35132 34412 35188 34414
rect 35292 34466 35348 34468
rect 35292 34414 35294 34466
rect 35294 34414 35346 34466
rect 35346 34414 35348 34466
rect 35292 34412 35348 34414
rect 35452 34466 35508 34468
rect 35452 34414 35454 34466
rect 35454 34414 35506 34466
rect 35506 34414 35508 34466
rect 35452 34412 35508 34414
rect 35612 34466 35668 34468
rect 35612 34414 35614 34466
rect 35614 34414 35666 34466
rect 35666 34414 35668 34466
rect 35612 34412 35668 34414
rect 35772 34466 35828 34468
rect 35772 34414 35774 34466
rect 35774 34414 35826 34466
rect 35826 34414 35828 34466
rect 35772 34412 35828 34414
rect 35932 34466 35988 34468
rect 35932 34414 35934 34466
rect 35934 34414 35986 34466
rect 35986 34414 35988 34466
rect 35932 34412 35988 34414
rect 36092 34466 36148 34468
rect 36092 34414 36094 34466
rect 36094 34414 36146 34466
rect 36146 34414 36148 34466
rect 36092 34412 36148 34414
rect 36252 34466 36308 34468
rect 36252 34414 36254 34466
rect 36254 34414 36306 34466
rect 36306 34414 36308 34466
rect 36252 34412 36308 34414
rect 36412 34466 36468 34468
rect 36412 34414 36414 34466
rect 36414 34414 36466 34466
rect 36466 34414 36468 34466
rect 36412 34412 36468 34414
rect 36572 34466 36628 34468
rect 36572 34414 36574 34466
rect 36574 34414 36626 34466
rect 36626 34414 36628 34466
rect 36572 34412 36628 34414
rect 36732 34466 36788 34468
rect 36732 34414 36734 34466
rect 36734 34414 36786 34466
rect 36786 34414 36788 34466
rect 36732 34412 36788 34414
rect 36892 34466 36948 34468
rect 36892 34414 36894 34466
rect 36894 34414 36946 34466
rect 36946 34414 36948 34466
rect 36892 34412 36948 34414
rect 37052 34466 37108 34468
rect 37052 34414 37054 34466
rect 37054 34414 37106 34466
rect 37106 34414 37108 34466
rect 37052 34412 37108 34414
rect 37212 34466 37268 34468
rect 37212 34414 37214 34466
rect 37214 34414 37266 34466
rect 37266 34414 37268 34466
rect 37212 34412 37268 34414
rect 37372 34466 37428 34468
rect 37372 34414 37374 34466
rect 37374 34414 37426 34466
rect 37426 34414 37428 34466
rect 37372 34412 37428 34414
rect 37532 34466 37588 34468
rect 37532 34414 37534 34466
rect 37534 34414 37586 34466
rect 37586 34414 37588 34466
rect 37532 34412 37588 34414
rect 37692 34466 37748 34468
rect 37692 34414 37694 34466
rect 37694 34414 37746 34466
rect 37746 34414 37748 34466
rect 37692 34412 37748 34414
rect 37852 34466 37908 34468
rect 37852 34414 37854 34466
rect 37854 34414 37906 34466
rect 37906 34414 37908 34466
rect 37852 34412 37908 34414
rect 38012 34466 38068 34468
rect 38012 34414 38014 34466
rect 38014 34414 38066 34466
rect 38066 34414 38068 34466
rect 38012 34412 38068 34414
rect 38172 34466 38228 34468
rect 38172 34414 38174 34466
rect 38174 34414 38226 34466
rect 38226 34414 38228 34466
rect 38172 34412 38228 34414
rect 38332 34466 38388 34468
rect 38332 34414 38334 34466
rect 38334 34414 38386 34466
rect 38386 34414 38388 34466
rect 38332 34412 38388 34414
rect 38492 34466 38548 34468
rect 38492 34414 38494 34466
rect 38494 34414 38546 34466
rect 38546 34414 38548 34466
rect 38492 34412 38548 34414
rect 38652 34466 38708 34468
rect 38652 34414 38654 34466
rect 38654 34414 38706 34466
rect 38706 34414 38708 34466
rect 38652 34412 38708 34414
rect 38812 34466 38868 34468
rect 38812 34414 38814 34466
rect 38814 34414 38866 34466
rect 38866 34414 38868 34466
rect 38812 34412 38868 34414
rect 38972 34466 39028 34468
rect 38972 34414 38974 34466
rect 38974 34414 39026 34466
rect 39026 34414 39028 34466
rect 38972 34412 39028 34414
rect 39132 34466 39188 34468
rect 39132 34414 39134 34466
rect 39134 34414 39186 34466
rect 39186 34414 39188 34466
rect 39132 34412 39188 34414
rect 39292 34466 39348 34468
rect 39292 34414 39294 34466
rect 39294 34414 39346 34466
rect 39346 34414 39348 34466
rect 39292 34412 39348 34414
rect 39452 34466 39508 34468
rect 39452 34414 39454 34466
rect 39454 34414 39506 34466
rect 39506 34414 39508 34466
rect 39452 34412 39508 34414
rect 39612 34466 39668 34468
rect 39612 34414 39614 34466
rect 39614 34414 39666 34466
rect 39666 34414 39668 34466
rect 39612 34412 39668 34414
rect 39772 34466 39828 34468
rect 39772 34414 39774 34466
rect 39774 34414 39826 34466
rect 39826 34414 39828 34466
rect 39772 34412 39828 34414
rect 39932 34466 39988 34468
rect 39932 34414 39934 34466
rect 39934 34414 39986 34466
rect 39986 34414 39988 34466
rect 39932 34412 39988 34414
rect 40092 34466 40148 34468
rect 40092 34414 40094 34466
rect 40094 34414 40146 34466
rect 40146 34414 40148 34466
rect 40092 34412 40148 34414
rect 40252 34466 40308 34468
rect 40252 34414 40254 34466
rect 40254 34414 40306 34466
rect 40306 34414 40308 34466
rect 40252 34412 40308 34414
rect 40412 34466 40468 34468
rect 40412 34414 40414 34466
rect 40414 34414 40466 34466
rect 40466 34414 40468 34466
rect 40412 34412 40468 34414
rect 40572 34466 40628 34468
rect 40572 34414 40574 34466
rect 40574 34414 40626 34466
rect 40626 34414 40628 34466
rect 40572 34412 40628 34414
rect 40732 34466 40788 34468
rect 40732 34414 40734 34466
rect 40734 34414 40786 34466
rect 40786 34414 40788 34466
rect 40732 34412 40788 34414
rect 40892 34466 40948 34468
rect 40892 34414 40894 34466
rect 40894 34414 40946 34466
rect 40946 34414 40948 34466
rect 40892 34412 40948 34414
rect 41052 34466 41108 34468
rect 41052 34414 41054 34466
rect 41054 34414 41106 34466
rect 41106 34414 41108 34466
rect 41052 34412 41108 34414
rect 41212 34466 41268 34468
rect 41212 34414 41214 34466
rect 41214 34414 41266 34466
rect 41266 34414 41268 34466
rect 41212 34412 41268 34414
rect 41372 34466 41428 34468
rect 41372 34414 41374 34466
rect 41374 34414 41426 34466
rect 41426 34414 41428 34466
rect 41372 34412 41428 34414
rect 41532 34466 41588 34468
rect 41532 34414 41534 34466
rect 41534 34414 41586 34466
rect 41586 34414 41588 34466
rect 41532 34412 41588 34414
rect 41692 34466 41748 34468
rect 41692 34414 41694 34466
rect 41694 34414 41746 34466
rect 41746 34414 41748 34466
rect 41692 34412 41748 34414
rect 41852 34466 41908 34468
rect 41852 34414 41854 34466
rect 41854 34414 41906 34466
rect 41906 34414 41908 34466
rect 41852 34412 41908 34414
rect 12 34306 68 34308
rect 12 34254 14 34306
rect 14 34254 66 34306
rect 66 34254 68 34306
rect 12 34252 68 34254
rect 172 34306 228 34308
rect 172 34254 174 34306
rect 174 34254 226 34306
rect 226 34254 228 34306
rect 172 34252 228 34254
rect 332 34306 388 34308
rect 332 34254 334 34306
rect 334 34254 386 34306
rect 386 34254 388 34306
rect 332 34252 388 34254
rect 492 34306 548 34308
rect 492 34254 494 34306
rect 494 34254 546 34306
rect 546 34254 548 34306
rect 492 34252 548 34254
rect 652 34306 708 34308
rect 652 34254 654 34306
rect 654 34254 706 34306
rect 706 34254 708 34306
rect 652 34252 708 34254
rect 812 34306 868 34308
rect 812 34254 814 34306
rect 814 34254 866 34306
rect 866 34254 868 34306
rect 812 34252 868 34254
rect 972 34306 1028 34308
rect 972 34254 974 34306
rect 974 34254 1026 34306
rect 1026 34254 1028 34306
rect 972 34252 1028 34254
rect 1132 34306 1188 34308
rect 1132 34254 1134 34306
rect 1134 34254 1186 34306
rect 1186 34254 1188 34306
rect 1132 34252 1188 34254
rect 1292 34306 1348 34308
rect 1292 34254 1294 34306
rect 1294 34254 1346 34306
rect 1346 34254 1348 34306
rect 1292 34252 1348 34254
rect 1452 34306 1508 34308
rect 1452 34254 1454 34306
rect 1454 34254 1506 34306
rect 1506 34254 1508 34306
rect 1452 34252 1508 34254
rect 1612 34306 1668 34308
rect 1612 34254 1614 34306
rect 1614 34254 1666 34306
rect 1666 34254 1668 34306
rect 1612 34252 1668 34254
rect 1772 34306 1828 34308
rect 1772 34254 1774 34306
rect 1774 34254 1826 34306
rect 1826 34254 1828 34306
rect 1772 34252 1828 34254
rect 1932 34306 1988 34308
rect 1932 34254 1934 34306
rect 1934 34254 1986 34306
rect 1986 34254 1988 34306
rect 1932 34252 1988 34254
rect 2092 34306 2148 34308
rect 2092 34254 2094 34306
rect 2094 34254 2146 34306
rect 2146 34254 2148 34306
rect 2092 34252 2148 34254
rect 2252 34306 2308 34308
rect 2252 34254 2254 34306
rect 2254 34254 2306 34306
rect 2306 34254 2308 34306
rect 2252 34252 2308 34254
rect 2412 34306 2468 34308
rect 2412 34254 2414 34306
rect 2414 34254 2466 34306
rect 2466 34254 2468 34306
rect 2412 34252 2468 34254
rect 2572 34306 2628 34308
rect 2572 34254 2574 34306
rect 2574 34254 2626 34306
rect 2626 34254 2628 34306
rect 2572 34252 2628 34254
rect 2732 34306 2788 34308
rect 2732 34254 2734 34306
rect 2734 34254 2786 34306
rect 2786 34254 2788 34306
rect 2732 34252 2788 34254
rect 2892 34306 2948 34308
rect 2892 34254 2894 34306
rect 2894 34254 2946 34306
rect 2946 34254 2948 34306
rect 2892 34252 2948 34254
rect 3052 34306 3108 34308
rect 3052 34254 3054 34306
rect 3054 34254 3106 34306
rect 3106 34254 3108 34306
rect 3052 34252 3108 34254
rect 3212 34306 3268 34308
rect 3212 34254 3214 34306
rect 3214 34254 3266 34306
rect 3266 34254 3268 34306
rect 3212 34252 3268 34254
rect 3372 34306 3428 34308
rect 3372 34254 3374 34306
rect 3374 34254 3426 34306
rect 3426 34254 3428 34306
rect 3372 34252 3428 34254
rect 3532 34306 3588 34308
rect 3532 34254 3534 34306
rect 3534 34254 3586 34306
rect 3586 34254 3588 34306
rect 3532 34252 3588 34254
rect 3692 34306 3748 34308
rect 3692 34254 3694 34306
rect 3694 34254 3746 34306
rect 3746 34254 3748 34306
rect 3692 34252 3748 34254
rect 3852 34306 3908 34308
rect 3852 34254 3854 34306
rect 3854 34254 3906 34306
rect 3906 34254 3908 34306
rect 3852 34252 3908 34254
rect 4012 34306 4068 34308
rect 4012 34254 4014 34306
rect 4014 34254 4066 34306
rect 4066 34254 4068 34306
rect 4012 34252 4068 34254
rect 4172 34306 4228 34308
rect 4172 34254 4174 34306
rect 4174 34254 4226 34306
rect 4226 34254 4228 34306
rect 4172 34252 4228 34254
rect 4332 34306 4388 34308
rect 4332 34254 4334 34306
rect 4334 34254 4386 34306
rect 4386 34254 4388 34306
rect 4332 34252 4388 34254
rect 4492 34306 4548 34308
rect 4492 34254 4494 34306
rect 4494 34254 4546 34306
rect 4546 34254 4548 34306
rect 4492 34252 4548 34254
rect 4652 34306 4708 34308
rect 4652 34254 4654 34306
rect 4654 34254 4706 34306
rect 4706 34254 4708 34306
rect 4652 34252 4708 34254
rect 4812 34306 4868 34308
rect 4812 34254 4814 34306
rect 4814 34254 4866 34306
rect 4866 34254 4868 34306
rect 4812 34252 4868 34254
rect 4972 34306 5028 34308
rect 4972 34254 4974 34306
rect 4974 34254 5026 34306
rect 5026 34254 5028 34306
rect 4972 34252 5028 34254
rect 5132 34306 5188 34308
rect 5132 34254 5134 34306
rect 5134 34254 5186 34306
rect 5186 34254 5188 34306
rect 5132 34252 5188 34254
rect 5292 34306 5348 34308
rect 5292 34254 5294 34306
rect 5294 34254 5346 34306
rect 5346 34254 5348 34306
rect 5292 34252 5348 34254
rect 5452 34306 5508 34308
rect 5452 34254 5454 34306
rect 5454 34254 5506 34306
rect 5506 34254 5508 34306
rect 5452 34252 5508 34254
rect 5612 34306 5668 34308
rect 5612 34254 5614 34306
rect 5614 34254 5666 34306
rect 5666 34254 5668 34306
rect 5612 34252 5668 34254
rect 5772 34306 5828 34308
rect 5772 34254 5774 34306
rect 5774 34254 5826 34306
rect 5826 34254 5828 34306
rect 5772 34252 5828 34254
rect 5932 34306 5988 34308
rect 5932 34254 5934 34306
rect 5934 34254 5986 34306
rect 5986 34254 5988 34306
rect 5932 34252 5988 34254
rect 6092 34306 6148 34308
rect 6092 34254 6094 34306
rect 6094 34254 6146 34306
rect 6146 34254 6148 34306
rect 6092 34252 6148 34254
rect 6252 34306 6308 34308
rect 6252 34254 6254 34306
rect 6254 34254 6306 34306
rect 6306 34254 6308 34306
rect 6252 34252 6308 34254
rect 6412 34306 6468 34308
rect 6412 34254 6414 34306
rect 6414 34254 6466 34306
rect 6466 34254 6468 34306
rect 6412 34252 6468 34254
rect 6572 34306 6628 34308
rect 6572 34254 6574 34306
rect 6574 34254 6626 34306
rect 6626 34254 6628 34306
rect 6572 34252 6628 34254
rect 6732 34306 6788 34308
rect 6732 34254 6734 34306
rect 6734 34254 6786 34306
rect 6786 34254 6788 34306
rect 6732 34252 6788 34254
rect 6892 34306 6948 34308
rect 6892 34254 6894 34306
rect 6894 34254 6946 34306
rect 6946 34254 6948 34306
rect 6892 34252 6948 34254
rect 7052 34306 7108 34308
rect 7052 34254 7054 34306
rect 7054 34254 7106 34306
rect 7106 34254 7108 34306
rect 7052 34252 7108 34254
rect 7212 34306 7268 34308
rect 7212 34254 7214 34306
rect 7214 34254 7266 34306
rect 7266 34254 7268 34306
rect 7212 34252 7268 34254
rect 7372 34306 7428 34308
rect 7372 34254 7374 34306
rect 7374 34254 7426 34306
rect 7426 34254 7428 34306
rect 7372 34252 7428 34254
rect 7532 34306 7588 34308
rect 7532 34254 7534 34306
rect 7534 34254 7586 34306
rect 7586 34254 7588 34306
rect 7532 34252 7588 34254
rect 7692 34306 7748 34308
rect 7692 34254 7694 34306
rect 7694 34254 7746 34306
rect 7746 34254 7748 34306
rect 7692 34252 7748 34254
rect 7852 34306 7908 34308
rect 7852 34254 7854 34306
rect 7854 34254 7906 34306
rect 7906 34254 7908 34306
rect 7852 34252 7908 34254
rect 8012 34306 8068 34308
rect 8012 34254 8014 34306
rect 8014 34254 8066 34306
rect 8066 34254 8068 34306
rect 8012 34252 8068 34254
rect 8172 34306 8228 34308
rect 8172 34254 8174 34306
rect 8174 34254 8226 34306
rect 8226 34254 8228 34306
rect 8172 34252 8228 34254
rect 8332 34306 8388 34308
rect 8332 34254 8334 34306
rect 8334 34254 8386 34306
rect 8386 34254 8388 34306
rect 8332 34252 8388 34254
rect 11532 34252 11588 34308
rect 11852 34252 11908 34308
rect 12492 34306 12548 34308
rect 12492 34254 12494 34306
rect 12494 34254 12546 34306
rect 12546 34254 12548 34306
rect 12492 34252 12548 34254
rect 12652 34306 12708 34308
rect 12652 34254 12654 34306
rect 12654 34254 12706 34306
rect 12706 34254 12708 34306
rect 12652 34252 12708 34254
rect 12812 34306 12868 34308
rect 12812 34254 12814 34306
rect 12814 34254 12866 34306
rect 12866 34254 12868 34306
rect 12812 34252 12868 34254
rect 12972 34306 13028 34308
rect 12972 34254 12974 34306
rect 12974 34254 13026 34306
rect 13026 34254 13028 34306
rect 12972 34252 13028 34254
rect 13132 34306 13188 34308
rect 13132 34254 13134 34306
rect 13134 34254 13186 34306
rect 13186 34254 13188 34306
rect 13132 34252 13188 34254
rect 13292 34306 13348 34308
rect 13292 34254 13294 34306
rect 13294 34254 13346 34306
rect 13346 34254 13348 34306
rect 13292 34252 13348 34254
rect 13452 34306 13508 34308
rect 13452 34254 13454 34306
rect 13454 34254 13506 34306
rect 13506 34254 13508 34306
rect 13452 34252 13508 34254
rect 13612 34306 13668 34308
rect 13612 34254 13614 34306
rect 13614 34254 13666 34306
rect 13666 34254 13668 34306
rect 13612 34252 13668 34254
rect 13772 34306 13828 34308
rect 13772 34254 13774 34306
rect 13774 34254 13826 34306
rect 13826 34254 13828 34306
rect 13772 34252 13828 34254
rect 13932 34306 13988 34308
rect 13932 34254 13934 34306
rect 13934 34254 13986 34306
rect 13986 34254 13988 34306
rect 13932 34252 13988 34254
rect 14092 34306 14148 34308
rect 14092 34254 14094 34306
rect 14094 34254 14146 34306
rect 14146 34254 14148 34306
rect 14092 34252 14148 34254
rect 14252 34306 14308 34308
rect 14252 34254 14254 34306
rect 14254 34254 14306 34306
rect 14306 34254 14308 34306
rect 14252 34252 14308 34254
rect 14412 34306 14468 34308
rect 14412 34254 14414 34306
rect 14414 34254 14466 34306
rect 14466 34254 14468 34306
rect 14412 34252 14468 34254
rect 14572 34306 14628 34308
rect 14572 34254 14574 34306
rect 14574 34254 14626 34306
rect 14626 34254 14628 34306
rect 14572 34252 14628 34254
rect 14732 34306 14788 34308
rect 14732 34254 14734 34306
rect 14734 34254 14786 34306
rect 14786 34254 14788 34306
rect 14732 34252 14788 34254
rect 14892 34306 14948 34308
rect 14892 34254 14894 34306
rect 14894 34254 14946 34306
rect 14946 34254 14948 34306
rect 14892 34252 14948 34254
rect 15052 34306 15108 34308
rect 15052 34254 15054 34306
rect 15054 34254 15106 34306
rect 15106 34254 15108 34306
rect 15052 34252 15108 34254
rect 15212 34306 15268 34308
rect 15212 34254 15214 34306
rect 15214 34254 15266 34306
rect 15266 34254 15268 34306
rect 15212 34252 15268 34254
rect 15372 34306 15428 34308
rect 15372 34254 15374 34306
rect 15374 34254 15426 34306
rect 15426 34254 15428 34306
rect 15372 34252 15428 34254
rect 15532 34306 15588 34308
rect 15532 34254 15534 34306
rect 15534 34254 15586 34306
rect 15586 34254 15588 34306
rect 15532 34252 15588 34254
rect 15692 34306 15748 34308
rect 15692 34254 15694 34306
rect 15694 34254 15746 34306
rect 15746 34254 15748 34306
rect 15692 34252 15748 34254
rect 15852 34306 15908 34308
rect 15852 34254 15854 34306
rect 15854 34254 15906 34306
rect 15906 34254 15908 34306
rect 15852 34252 15908 34254
rect 16012 34306 16068 34308
rect 16012 34254 16014 34306
rect 16014 34254 16066 34306
rect 16066 34254 16068 34306
rect 16012 34252 16068 34254
rect 16172 34306 16228 34308
rect 16172 34254 16174 34306
rect 16174 34254 16226 34306
rect 16226 34254 16228 34306
rect 16172 34252 16228 34254
rect 16332 34306 16388 34308
rect 16332 34254 16334 34306
rect 16334 34254 16386 34306
rect 16386 34254 16388 34306
rect 16332 34252 16388 34254
rect 16492 34306 16548 34308
rect 16492 34254 16494 34306
rect 16494 34254 16546 34306
rect 16546 34254 16548 34306
rect 16492 34252 16548 34254
rect 16652 34306 16708 34308
rect 16652 34254 16654 34306
rect 16654 34254 16706 34306
rect 16706 34254 16708 34306
rect 16652 34252 16708 34254
rect 16812 34306 16868 34308
rect 16812 34254 16814 34306
rect 16814 34254 16866 34306
rect 16866 34254 16868 34306
rect 16812 34252 16868 34254
rect 16972 34306 17028 34308
rect 16972 34254 16974 34306
rect 16974 34254 17026 34306
rect 17026 34254 17028 34306
rect 16972 34252 17028 34254
rect 17132 34306 17188 34308
rect 17132 34254 17134 34306
rect 17134 34254 17186 34306
rect 17186 34254 17188 34306
rect 17132 34252 17188 34254
rect 17292 34306 17348 34308
rect 17292 34254 17294 34306
rect 17294 34254 17346 34306
rect 17346 34254 17348 34306
rect 17292 34252 17348 34254
rect 17452 34306 17508 34308
rect 17452 34254 17454 34306
rect 17454 34254 17506 34306
rect 17506 34254 17508 34306
rect 17452 34252 17508 34254
rect 17612 34306 17668 34308
rect 17612 34254 17614 34306
rect 17614 34254 17666 34306
rect 17666 34254 17668 34306
rect 17612 34252 17668 34254
rect 17772 34306 17828 34308
rect 17772 34254 17774 34306
rect 17774 34254 17826 34306
rect 17826 34254 17828 34306
rect 17772 34252 17828 34254
rect 17932 34306 17988 34308
rect 17932 34254 17934 34306
rect 17934 34254 17986 34306
rect 17986 34254 17988 34306
rect 17932 34252 17988 34254
rect 18092 34306 18148 34308
rect 18092 34254 18094 34306
rect 18094 34254 18146 34306
rect 18146 34254 18148 34306
rect 18092 34252 18148 34254
rect 18252 34306 18308 34308
rect 18252 34254 18254 34306
rect 18254 34254 18306 34306
rect 18306 34254 18308 34306
rect 18252 34252 18308 34254
rect 18412 34306 18468 34308
rect 18412 34254 18414 34306
rect 18414 34254 18466 34306
rect 18466 34254 18468 34306
rect 18412 34252 18468 34254
rect 18572 34306 18628 34308
rect 18572 34254 18574 34306
rect 18574 34254 18626 34306
rect 18626 34254 18628 34306
rect 18572 34252 18628 34254
rect 18732 34306 18788 34308
rect 18732 34254 18734 34306
rect 18734 34254 18786 34306
rect 18786 34254 18788 34306
rect 18732 34252 18788 34254
rect 18892 34306 18948 34308
rect 18892 34254 18894 34306
rect 18894 34254 18946 34306
rect 18946 34254 18948 34306
rect 18892 34252 18948 34254
rect 19532 34252 19588 34308
rect 19852 34252 19908 34308
rect 23132 34306 23188 34308
rect 23132 34254 23134 34306
rect 23134 34254 23186 34306
rect 23186 34254 23188 34306
rect 23132 34252 23188 34254
rect 23292 34306 23348 34308
rect 23292 34254 23294 34306
rect 23294 34254 23346 34306
rect 23346 34254 23348 34306
rect 23292 34252 23348 34254
rect 23452 34306 23508 34308
rect 23452 34254 23454 34306
rect 23454 34254 23506 34306
rect 23506 34254 23508 34306
rect 23452 34252 23508 34254
rect 23612 34306 23668 34308
rect 23612 34254 23614 34306
rect 23614 34254 23666 34306
rect 23666 34254 23668 34306
rect 23612 34252 23668 34254
rect 23772 34306 23828 34308
rect 23772 34254 23774 34306
rect 23774 34254 23826 34306
rect 23826 34254 23828 34306
rect 23772 34252 23828 34254
rect 23932 34306 23988 34308
rect 23932 34254 23934 34306
rect 23934 34254 23986 34306
rect 23986 34254 23988 34306
rect 23932 34252 23988 34254
rect 24092 34306 24148 34308
rect 24092 34254 24094 34306
rect 24094 34254 24146 34306
rect 24146 34254 24148 34306
rect 24092 34252 24148 34254
rect 24252 34306 24308 34308
rect 24252 34254 24254 34306
rect 24254 34254 24306 34306
rect 24306 34254 24308 34306
rect 24252 34252 24308 34254
rect 24412 34306 24468 34308
rect 24412 34254 24414 34306
rect 24414 34254 24466 34306
rect 24466 34254 24468 34306
rect 24412 34252 24468 34254
rect 24572 34306 24628 34308
rect 24572 34254 24574 34306
rect 24574 34254 24626 34306
rect 24626 34254 24628 34306
rect 24572 34252 24628 34254
rect 24732 34306 24788 34308
rect 24732 34254 24734 34306
rect 24734 34254 24786 34306
rect 24786 34254 24788 34306
rect 24732 34252 24788 34254
rect 24892 34306 24948 34308
rect 24892 34254 24894 34306
rect 24894 34254 24946 34306
rect 24946 34254 24948 34306
rect 24892 34252 24948 34254
rect 25052 34306 25108 34308
rect 25052 34254 25054 34306
rect 25054 34254 25106 34306
rect 25106 34254 25108 34306
rect 25052 34252 25108 34254
rect 25212 34306 25268 34308
rect 25212 34254 25214 34306
rect 25214 34254 25266 34306
rect 25266 34254 25268 34306
rect 25212 34252 25268 34254
rect 25372 34306 25428 34308
rect 25372 34254 25374 34306
rect 25374 34254 25426 34306
rect 25426 34254 25428 34306
rect 25372 34252 25428 34254
rect 25532 34306 25588 34308
rect 25532 34254 25534 34306
rect 25534 34254 25586 34306
rect 25586 34254 25588 34306
rect 25532 34252 25588 34254
rect 25692 34306 25748 34308
rect 25692 34254 25694 34306
rect 25694 34254 25746 34306
rect 25746 34254 25748 34306
rect 25692 34252 25748 34254
rect 25852 34306 25908 34308
rect 25852 34254 25854 34306
rect 25854 34254 25906 34306
rect 25906 34254 25908 34306
rect 25852 34252 25908 34254
rect 26012 34306 26068 34308
rect 26012 34254 26014 34306
rect 26014 34254 26066 34306
rect 26066 34254 26068 34306
rect 26012 34252 26068 34254
rect 26172 34306 26228 34308
rect 26172 34254 26174 34306
rect 26174 34254 26226 34306
rect 26226 34254 26228 34306
rect 26172 34252 26228 34254
rect 26332 34306 26388 34308
rect 26332 34254 26334 34306
rect 26334 34254 26386 34306
rect 26386 34254 26388 34306
rect 26332 34252 26388 34254
rect 26492 34306 26548 34308
rect 26492 34254 26494 34306
rect 26494 34254 26546 34306
rect 26546 34254 26548 34306
rect 26492 34252 26548 34254
rect 26652 34306 26708 34308
rect 26652 34254 26654 34306
rect 26654 34254 26706 34306
rect 26706 34254 26708 34306
rect 26652 34252 26708 34254
rect 26812 34306 26868 34308
rect 26812 34254 26814 34306
rect 26814 34254 26866 34306
rect 26866 34254 26868 34306
rect 26812 34252 26868 34254
rect 26972 34306 27028 34308
rect 26972 34254 26974 34306
rect 26974 34254 27026 34306
rect 27026 34254 27028 34306
rect 26972 34252 27028 34254
rect 27132 34306 27188 34308
rect 27132 34254 27134 34306
rect 27134 34254 27186 34306
rect 27186 34254 27188 34306
rect 27132 34252 27188 34254
rect 27292 34306 27348 34308
rect 27292 34254 27294 34306
rect 27294 34254 27346 34306
rect 27346 34254 27348 34306
rect 27292 34252 27348 34254
rect 27452 34306 27508 34308
rect 27452 34254 27454 34306
rect 27454 34254 27506 34306
rect 27506 34254 27508 34306
rect 27452 34252 27508 34254
rect 27612 34306 27668 34308
rect 27612 34254 27614 34306
rect 27614 34254 27666 34306
rect 27666 34254 27668 34306
rect 27612 34252 27668 34254
rect 27772 34306 27828 34308
rect 27772 34254 27774 34306
rect 27774 34254 27826 34306
rect 27826 34254 27828 34306
rect 27772 34252 27828 34254
rect 27932 34306 27988 34308
rect 27932 34254 27934 34306
rect 27934 34254 27986 34306
rect 27986 34254 27988 34306
rect 27932 34252 27988 34254
rect 28092 34306 28148 34308
rect 28092 34254 28094 34306
rect 28094 34254 28146 34306
rect 28146 34254 28148 34306
rect 28092 34252 28148 34254
rect 28252 34306 28308 34308
rect 28252 34254 28254 34306
rect 28254 34254 28306 34306
rect 28306 34254 28308 34306
rect 28252 34252 28308 34254
rect 28412 34306 28468 34308
rect 28412 34254 28414 34306
rect 28414 34254 28466 34306
rect 28466 34254 28468 34306
rect 28412 34252 28468 34254
rect 28572 34306 28628 34308
rect 28572 34254 28574 34306
rect 28574 34254 28626 34306
rect 28626 34254 28628 34306
rect 28572 34252 28628 34254
rect 28732 34306 28788 34308
rect 28732 34254 28734 34306
rect 28734 34254 28786 34306
rect 28786 34254 28788 34306
rect 28732 34252 28788 34254
rect 28892 34306 28948 34308
rect 28892 34254 28894 34306
rect 28894 34254 28946 34306
rect 28946 34254 28948 34306
rect 28892 34252 28948 34254
rect 29052 34306 29108 34308
rect 29052 34254 29054 34306
rect 29054 34254 29106 34306
rect 29106 34254 29108 34306
rect 29052 34252 29108 34254
rect 29212 34306 29268 34308
rect 29212 34254 29214 34306
rect 29214 34254 29266 34306
rect 29266 34254 29268 34306
rect 29212 34252 29268 34254
rect 29372 34306 29428 34308
rect 29372 34254 29374 34306
rect 29374 34254 29426 34306
rect 29426 34254 29428 34306
rect 29372 34252 29428 34254
rect 30012 34252 30068 34308
rect 30332 34252 30388 34308
rect 33532 34306 33588 34308
rect 33532 34254 33534 34306
rect 33534 34254 33586 34306
rect 33586 34254 33588 34306
rect 33532 34252 33588 34254
rect 33692 34306 33748 34308
rect 33692 34254 33694 34306
rect 33694 34254 33746 34306
rect 33746 34254 33748 34306
rect 33692 34252 33748 34254
rect 33852 34306 33908 34308
rect 33852 34254 33854 34306
rect 33854 34254 33906 34306
rect 33906 34254 33908 34306
rect 33852 34252 33908 34254
rect 34012 34306 34068 34308
rect 34012 34254 34014 34306
rect 34014 34254 34066 34306
rect 34066 34254 34068 34306
rect 34012 34252 34068 34254
rect 34172 34306 34228 34308
rect 34172 34254 34174 34306
rect 34174 34254 34226 34306
rect 34226 34254 34228 34306
rect 34172 34252 34228 34254
rect 34332 34306 34388 34308
rect 34332 34254 34334 34306
rect 34334 34254 34386 34306
rect 34386 34254 34388 34306
rect 34332 34252 34388 34254
rect 34492 34306 34548 34308
rect 34492 34254 34494 34306
rect 34494 34254 34546 34306
rect 34546 34254 34548 34306
rect 34492 34252 34548 34254
rect 34652 34306 34708 34308
rect 34652 34254 34654 34306
rect 34654 34254 34706 34306
rect 34706 34254 34708 34306
rect 34652 34252 34708 34254
rect 34812 34306 34868 34308
rect 34812 34254 34814 34306
rect 34814 34254 34866 34306
rect 34866 34254 34868 34306
rect 34812 34252 34868 34254
rect 34972 34306 35028 34308
rect 34972 34254 34974 34306
rect 34974 34254 35026 34306
rect 35026 34254 35028 34306
rect 34972 34252 35028 34254
rect 35132 34306 35188 34308
rect 35132 34254 35134 34306
rect 35134 34254 35186 34306
rect 35186 34254 35188 34306
rect 35132 34252 35188 34254
rect 35292 34306 35348 34308
rect 35292 34254 35294 34306
rect 35294 34254 35346 34306
rect 35346 34254 35348 34306
rect 35292 34252 35348 34254
rect 35452 34306 35508 34308
rect 35452 34254 35454 34306
rect 35454 34254 35506 34306
rect 35506 34254 35508 34306
rect 35452 34252 35508 34254
rect 35612 34306 35668 34308
rect 35612 34254 35614 34306
rect 35614 34254 35666 34306
rect 35666 34254 35668 34306
rect 35612 34252 35668 34254
rect 35772 34306 35828 34308
rect 35772 34254 35774 34306
rect 35774 34254 35826 34306
rect 35826 34254 35828 34306
rect 35772 34252 35828 34254
rect 35932 34306 35988 34308
rect 35932 34254 35934 34306
rect 35934 34254 35986 34306
rect 35986 34254 35988 34306
rect 35932 34252 35988 34254
rect 36092 34306 36148 34308
rect 36092 34254 36094 34306
rect 36094 34254 36146 34306
rect 36146 34254 36148 34306
rect 36092 34252 36148 34254
rect 36252 34306 36308 34308
rect 36252 34254 36254 34306
rect 36254 34254 36306 34306
rect 36306 34254 36308 34306
rect 36252 34252 36308 34254
rect 36412 34306 36468 34308
rect 36412 34254 36414 34306
rect 36414 34254 36466 34306
rect 36466 34254 36468 34306
rect 36412 34252 36468 34254
rect 36572 34306 36628 34308
rect 36572 34254 36574 34306
rect 36574 34254 36626 34306
rect 36626 34254 36628 34306
rect 36572 34252 36628 34254
rect 36732 34306 36788 34308
rect 36732 34254 36734 34306
rect 36734 34254 36786 34306
rect 36786 34254 36788 34306
rect 36732 34252 36788 34254
rect 36892 34306 36948 34308
rect 36892 34254 36894 34306
rect 36894 34254 36946 34306
rect 36946 34254 36948 34306
rect 36892 34252 36948 34254
rect 37052 34306 37108 34308
rect 37052 34254 37054 34306
rect 37054 34254 37106 34306
rect 37106 34254 37108 34306
rect 37052 34252 37108 34254
rect 37212 34306 37268 34308
rect 37212 34254 37214 34306
rect 37214 34254 37266 34306
rect 37266 34254 37268 34306
rect 37212 34252 37268 34254
rect 37372 34306 37428 34308
rect 37372 34254 37374 34306
rect 37374 34254 37426 34306
rect 37426 34254 37428 34306
rect 37372 34252 37428 34254
rect 37532 34306 37588 34308
rect 37532 34254 37534 34306
rect 37534 34254 37586 34306
rect 37586 34254 37588 34306
rect 37532 34252 37588 34254
rect 37692 34306 37748 34308
rect 37692 34254 37694 34306
rect 37694 34254 37746 34306
rect 37746 34254 37748 34306
rect 37692 34252 37748 34254
rect 37852 34306 37908 34308
rect 37852 34254 37854 34306
rect 37854 34254 37906 34306
rect 37906 34254 37908 34306
rect 37852 34252 37908 34254
rect 38012 34306 38068 34308
rect 38012 34254 38014 34306
rect 38014 34254 38066 34306
rect 38066 34254 38068 34306
rect 38012 34252 38068 34254
rect 38172 34306 38228 34308
rect 38172 34254 38174 34306
rect 38174 34254 38226 34306
rect 38226 34254 38228 34306
rect 38172 34252 38228 34254
rect 38332 34306 38388 34308
rect 38332 34254 38334 34306
rect 38334 34254 38386 34306
rect 38386 34254 38388 34306
rect 38332 34252 38388 34254
rect 38492 34306 38548 34308
rect 38492 34254 38494 34306
rect 38494 34254 38546 34306
rect 38546 34254 38548 34306
rect 38492 34252 38548 34254
rect 38652 34306 38708 34308
rect 38652 34254 38654 34306
rect 38654 34254 38706 34306
rect 38706 34254 38708 34306
rect 38652 34252 38708 34254
rect 38812 34306 38868 34308
rect 38812 34254 38814 34306
rect 38814 34254 38866 34306
rect 38866 34254 38868 34306
rect 38812 34252 38868 34254
rect 38972 34306 39028 34308
rect 38972 34254 38974 34306
rect 38974 34254 39026 34306
rect 39026 34254 39028 34306
rect 38972 34252 39028 34254
rect 39132 34306 39188 34308
rect 39132 34254 39134 34306
rect 39134 34254 39186 34306
rect 39186 34254 39188 34306
rect 39132 34252 39188 34254
rect 39292 34306 39348 34308
rect 39292 34254 39294 34306
rect 39294 34254 39346 34306
rect 39346 34254 39348 34306
rect 39292 34252 39348 34254
rect 39452 34306 39508 34308
rect 39452 34254 39454 34306
rect 39454 34254 39506 34306
rect 39506 34254 39508 34306
rect 39452 34252 39508 34254
rect 39612 34306 39668 34308
rect 39612 34254 39614 34306
rect 39614 34254 39666 34306
rect 39666 34254 39668 34306
rect 39612 34252 39668 34254
rect 39772 34306 39828 34308
rect 39772 34254 39774 34306
rect 39774 34254 39826 34306
rect 39826 34254 39828 34306
rect 39772 34252 39828 34254
rect 39932 34306 39988 34308
rect 39932 34254 39934 34306
rect 39934 34254 39986 34306
rect 39986 34254 39988 34306
rect 39932 34252 39988 34254
rect 40092 34306 40148 34308
rect 40092 34254 40094 34306
rect 40094 34254 40146 34306
rect 40146 34254 40148 34306
rect 40092 34252 40148 34254
rect 40252 34306 40308 34308
rect 40252 34254 40254 34306
rect 40254 34254 40306 34306
rect 40306 34254 40308 34306
rect 40252 34252 40308 34254
rect 40412 34306 40468 34308
rect 40412 34254 40414 34306
rect 40414 34254 40466 34306
rect 40466 34254 40468 34306
rect 40412 34252 40468 34254
rect 40572 34306 40628 34308
rect 40572 34254 40574 34306
rect 40574 34254 40626 34306
rect 40626 34254 40628 34306
rect 40572 34252 40628 34254
rect 40732 34306 40788 34308
rect 40732 34254 40734 34306
rect 40734 34254 40786 34306
rect 40786 34254 40788 34306
rect 40732 34252 40788 34254
rect 40892 34306 40948 34308
rect 40892 34254 40894 34306
rect 40894 34254 40946 34306
rect 40946 34254 40948 34306
rect 40892 34252 40948 34254
rect 41052 34306 41108 34308
rect 41052 34254 41054 34306
rect 41054 34254 41106 34306
rect 41106 34254 41108 34306
rect 41052 34252 41108 34254
rect 41212 34306 41268 34308
rect 41212 34254 41214 34306
rect 41214 34254 41266 34306
rect 41266 34254 41268 34306
rect 41212 34252 41268 34254
rect 41372 34306 41428 34308
rect 41372 34254 41374 34306
rect 41374 34254 41426 34306
rect 41426 34254 41428 34306
rect 41372 34252 41428 34254
rect 41532 34306 41588 34308
rect 41532 34254 41534 34306
rect 41534 34254 41586 34306
rect 41586 34254 41588 34306
rect 41532 34252 41588 34254
rect 41692 34306 41748 34308
rect 41692 34254 41694 34306
rect 41694 34254 41746 34306
rect 41746 34254 41748 34306
rect 41692 34252 41748 34254
rect 41852 34306 41908 34308
rect 41852 34254 41854 34306
rect 41854 34254 41906 34306
rect 41906 34254 41908 34306
rect 41852 34252 41908 34254
rect 11692 34092 11748 34148
rect 19692 34092 19748 34148
rect 30172 34092 30228 34148
rect 12 33986 68 33988
rect 12 33934 14 33986
rect 14 33934 66 33986
rect 66 33934 68 33986
rect 12 33932 68 33934
rect 172 33986 228 33988
rect 172 33934 174 33986
rect 174 33934 226 33986
rect 226 33934 228 33986
rect 172 33932 228 33934
rect 332 33986 388 33988
rect 332 33934 334 33986
rect 334 33934 386 33986
rect 386 33934 388 33986
rect 332 33932 388 33934
rect 492 33986 548 33988
rect 492 33934 494 33986
rect 494 33934 546 33986
rect 546 33934 548 33986
rect 492 33932 548 33934
rect 652 33986 708 33988
rect 652 33934 654 33986
rect 654 33934 706 33986
rect 706 33934 708 33986
rect 652 33932 708 33934
rect 812 33986 868 33988
rect 812 33934 814 33986
rect 814 33934 866 33986
rect 866 33934 868 33986
rect 812 33932 868 33934
rect 972 33986 1028 33988
rect 972 33934 974 33986
rect 974 33934 1026 33986
rect 1026 33934 1028 33986
rect 972 33932 1028 33934
rect 1132 33986 1188 33988
rect 1132 33934 1134 33986
rect 1134 33934 1186 33986
rect 1186 33934 1188 33986
rect 1132 33932 1188 33934
rect 1292 33986 1348 33988
rect 1292 33934 1294 33986
rect 1294 33934 1346 33986
rect 1346 33934 1348 33986
rect 1292 33932 1348 33934
rect 1452 33986 1508 33988
rect 1452 33934 1454 33986
rect 1454 33934 1506 33986
rect 1506 33934 1508 33986
rect 1452 33932 1508 33934
rect 1612 33986 1668 33988
rect 1612 33934 1614 33986
rect 1614 33934 1666 33986
rect 1666 33934 1668 33986
rect 1612 33932 1668 33934
rect 1772 33986 1828 33988
rect 1772 33934 1774 33986
rect 1774 33934 1826 33986
rect 1826 33934 1828 33986
rect 1772 33932 1828 33934
rect 1932 33986 1988 33988
rect 1932 33934 1934 33986
rect 1934 33934 1986 33986
rect 1986 33934 1988 33986
rect 1932 33932 1988 33934
rect 2092 33986 2148 33988
rect 2092 33934 2094 33986
rect 2094 33934 2146 33986
rect 2146 33934 2148 33986
rect 2092 33932 2148 33934
rect 2252 33986 2308 33988
rect 2252 33934 2254 33986
rect 2254 33934 2306 33986
rect 2306 33934 2308 33986
rect 2252 33932 2308 33934
rect 2412 33986 2468 33988
rect 2412 33934 2414 33986
rect 2414 33934 2466 33986
rect 2466 33934 2468 33986
rect 2412 33932 2468 33934
rect 2572 33986 2628 33988
rect 2572 33934 2574 33986
rect 2574 33934 2626 33986
rect 2626 33934 2628 33986
rect 2572 33932 2628 33934
rect 2732 33986 2788 33988
rect 2732 33934 2734 33986
rect 2734 33934 2786 33986
rect 2786 33934 2788 33986
rect 2732 33932 2788 33934
rect 2892 33986 2948 33988
rect 2892 33934 2894 33986
rect 2894 33934 2946 33986
rect 2946 33934 2948 33986
rect 2892 33932 2948 33934
rect 3052 33986 3108 33988
rect 3052 33934 3054 33986
rect 3054 33934 3106 33986
rect 3106 33934 3108 33986
rect 3052 33932 3108 33934
rect 3212 33986 3268 33988
rect 3212 33934 3214 33986
rect 3214 33934 3266 33986
rect 3266 33934 3268 33986
rect 3212 33932 3268 33934
rect 3372 33986 3428 33988
rect 3372 33934 3374 33986
rect 3374 33934 3426 33986
rect 3426 33934 3428 33986
rect 3372 33932 3428 33934
rect 3532 33986 3588 33988
rect 3532 33934 3534 33986
rect 3534 33934 3586 33986
rect 3586 33934 3588 33986
rect 3532 33932 3588 33934
rect 3692 33986 3748 33988
rect 3692 33934 3694 33986
rect 3694 33934 3746 33986
rect 3746 33934 3748 33986
rect 3692 33932 3748 33934
rect 3852 33986 3908 33988
rect 3852 33934 3854 33986
rect 3854 33934 3906 33986
rect 3906 33934 3908 33986
rect 3852 33932 3908 33934
rect 4012 33986 4068 33988
rect 4012 33934 4014 33986
rect 4014 33934 4066 33986
rect 4066 33934 4068 33986
rect 4012 33932 4068 33934
rect 4172 33986 4228 33988
rect 4172 33934 4174 33986
rect 4174 33934 4226 33986
rect 4226 33934 4228 33986
rect 4172 33932 4228 33934
rect 4332 33986 4388 33988
rect 4332 33934 4334 33986
rect 4334 33934 4386 33986
rect 4386 33934 4388 33986
rect 4332 33932 4388 33934
rect 4492 33986 4548 33988
rect 4492 33934 4494 33986
rect 4494 33934 4546 33986
rect 4546 33934 4548 33986
rect 4492 33932 4548 33934
rect 4652 33986 4708 33988
rect 4652 33934 4654 33986
rect 4654 33934 4706 33986
rect 4706 33934 4708 33986
rect 4652 33932 4708 33934
rect 4812 33986 4868 33988
rect 4812 33934 4814 33986
rect 4814 33934 4866 33986
rect 4866 33934 4868 33986
rect 4812 33932 4868 33934
rect 4972 33986 5028 33988
rect 4972 33934 4974 33986
rect 4974 33934 5026 33986
rect 5026 33934 5028 33986
rect 4972 33932 5028 33934
rect 5132 33986 5188 33988
rect 5132 33934 5134 33986
rect 5134 33934 5186 33986
rect 5186 33934 5188 33986
rect 5132 33932 5188 33934
rect 5292 33986 5348 33988
rect 5292 33934 5294 33986
rect 5294 33934 5346 33986
rect 5346 33934 5348 33986
rect 5292 33932 5348 33934
rect 5452 33986 5508 33988
rect 5452 33934 5454 33986
rect 5454 33934 5506 33986
rect 5506 33934 5508 33986
rect 5452 33932 5508 33934
rect 5612 33986 5668 33988
rect 5612 33934 5614 33986
rect 5614 33934 5666 33986
rect 5666 33934 5668 33986
rect 5612 33932 5668 33934
rect 5772 33986 5828 33988
rect 5772 33934 5774 33986
rect 5774 33934 5826 33986
rect 5826 33934 5828 33986
rect 5772 33932 5828 33934
rect 5932 33986 5988 33988
rect 5932 33934 5934 33986
rect 5934 33934 5986 33986
rect 5986 33934 5988 33986
rect 5932 33932 5988 33934
rect 6092 33986 6148 33988
rect 6092 33934 6094 33986
rect 6094 33934 6146 33986
rect 6146 33934 6148 33986
rect 6092 33932 6148 33934
rect 6252 33986 6308 33988
rect 6252 33934 6254 33986
rect 6254 33934 6306 33986
rect 6306 33934 6308 33986
rect 6252 33932 6308 33934
rect 6412 33986 6468 33988
rect 6412 33934 6414 33986
rect 6414 33934 6466 33986
rect 6466 33934 6468 33986
rect 6412 33932 6468 33934
rect 6572 33986 6628 33988
rect 6572 33934 6574 33986
rect 6574 33934 6626 33986
rect 6626 33934 6628 33986
rect 6572 33932 6628 33934
rect 6732 33986 6788 33988
rect 6732 33934 6734 33986
rect 6734 33934 6786 33986
rect 6786 33934 6788 33986
rect 6732 33932 6788 33934
rect 6892 33986 6948 33988
rect 6892 33934 6894 33986
rect 6894 33934 6946 33986
rect 6946 33934 6948 33986
rect 6892 33932 6948 33934
rect 7052 33986 7108 33988
rect 7052 33934 7054 33986
rect 7054 33934 7106 33986
rect 7106 33934 7108 33986
rect 7052 33932 7108 33934
rect 7212 33986 7268 33988
rect 7212 33934 7214 33986
rect 7214 33934 7266 33986
rect 7266 33934 7268 33986
rect 7212 33932 7268 33934
rect 7372 33986 7428 33988
rect 7372 33934 7374 33986
rect 7374 33934 7426 33986
rect 7426 33934 7428 33986
rect 7372 33932 7428 33934
rect 7532 33986 7588 33988
rect 7532 33934 7534 33986
rect 7534 33934 7586 33986
rect 7586 33934 7588 33986
rect 7532 33932 7588 33934
rect 7692 33986 7748 33988
rect 7692 33934 7694 33986
rect 7694 33934 7746 33986
rect 7746 33934 7748 33986
rect 7692 33932 7748 33934
rect 7852 33986 7908 33988
rect 7852 33934 7854 33986
rect 7854 33934 7906 33986
rect 7906 33934 7908 33986
rect 7852 33932 7908 33934
rect 8012 33986 8068 33988
rect 8012 33934 8014 33986
rect 8014 33934 8066 33986
rect 8066 33934 8068 33986
rect 8012 33932 8068 33934
rect 8172 33986 8228 33988
rect 8172 33934 8174 33986
rect 8174 33934 8226 33986
rect 8226 33934 8228 33986
rect 8172 33932 8228 33934
rect 8332 33986 8388 33988
rect 8332 33934 8334 33986
rect 8334 33934 8386 33986
rect 8386 33934 8388 33986
rect 8332 33932 8388 33934
rect 11532 33932 11588 33988
rect 11852 33932 11908 33988
rect 12492 33986 12548 33988
rect 12492 33934 12494 33986
rect 12494 33934 12546 33986
rect 12546 33934 12548 33986
rect 12492 33932 12548 33934
rect 12652 33986 12708 33988
rect 12652 33934 12654 33986
rect 12654 33934 12706 33986
rect 12706 33934 12708 33986
rect 12652 33932 12708 33934
rect 12812 33986 12868 33988
rect 12812 33934 12814 33986
rect 12814 33934 12866 33986
rect 12866 33934 12868 33986
rect 12812 33932 12868 33934
rect 12972 33986 13028 33988
rect 12972 33934 12974 33986
rect 12974 33934 13026 33986
rect 13026 33934 13028 33986
rect 12972 33932 13028 33934
rect 13132 33986 13188 33988
rect 13132 33934 13134 33986
rect 13134 33934 13186 33986
rect 13186 33934 13188 33986
rect 13132 33932 13188 33934
rect 13292 33986 13348 33988
rect 13292 33934 13294 33986
rect 13294 33934 13346 33986
rect 13346 33934 13348 33986
rect 13292 33932 13348 33934
rect 13452 33986 13508 33988
rect 13452 33934 13454 33986
rect 13454 33934 13506 33986
rect 13506 33934 13508 33986
rect 13452 33932 13508 33934
rect 13612 33986 13668 33988
rect 13612 33934 13614 33986
rect 13614 33934 13666 33986
rect 13666 33934 13668 33986
rect 13612 33932 13668 33934
rect 13772 33986 13828 33988
rect 13772 33934 13774 33986
rect 13774 33934 13826 33986
rect 13826 33934 13828 33986
rect 13772 33932 13828 33934
rect 13932 33986 13988 33988
rect 13932 33934 13934 33986
rect 13934 33934 13986 33986
rect 13986 33934 13988 33986
rect 13932 33932 13988 33934
rect 14092 33986 14148 33988
rect 14092 33934 14094 33986
rect 14094 33934 14146 33986
rect 14146 33934 14148 33986
rect 14092 33932 14148 33934
rect 14252 33986 14308 33988
rect 14252 33934 14254 33986
rect 14254 33934 14306 33986
rect 14306 33934 14308 33986
rect 14252 33932 14308 33934
rect 14412 33986 14468 33988
rect 14412 33934 14414 33986
rect 14414 33934 14466 33986
rect 14466 33934 14468 33986
rect 14412 33932 14468 33934
rect 14572 33986 14628 33988
rect 14572 33934 14574 33986
rect 14574 33934 14626 33986
rect 14626 33934 14628 33986
rect 14572 33932 14628 33934
rect 14732 33986 14788 33988
rect 14732 33934 14734 33986
rect 14734 33934 14786 33986
rect 14786 33934 14788 33986
rect 14732 33932 14788 33934
rect 14892 33986 14948 33988
rect 14892 33934 14894 33986
rect 14894 33934 14946 33986
rect 14946 33934 14948 33986
rect 14892 33932 14948 33934
rect 15052 33986 15108 33988
rect 15052 33934 15054 33986
rect 15054 33934 15106 33986
rect 15106 33934 15108 33986
rect 15052 33932 15108 33934
rect 15212 33986 15268 33988
rect 15212 33934 15214 33986
rect 15214 33934 15266 33986
rect 15266 33934 15268 33986
rect 15212 33932 15268 33934
rect 15372 33986 15428 33988
rect 15372 33934 15374 33986
rect 15374 33934 15426 33986
rect 15426 33934 15428 33986
rect 15372 33932 15428 33934
rect 15532 33986 15588 33988
rect 15532 33934 15534 33986
rect 15534 33934 15586 33986
rect 15586 33934 15588 33986
rect 15532 33932 15588 33934
rect 15692 33986 15748 33988
rect 15692 33934 15694 33986
rect 15694 33934 15746 33986
rect 15746 33934 15748 33986
rect 15692 33932 15748 33934
rect 15852 33986 15908 33988
rect 15852 33934 15854 33986
rect 15854 33934 15906 33986
rect 15906 33934 15908 33986
rect 15852 33932 15908 33934
rect 16012 33986 16068 33988
rect 16012 33934 16014 33986
rect 16014 33934 16066 33986
rect 16066 33934 16068 33986
rect 16012 33932 16068 33934
rect 16172 33986 16228 33988
rect 16172 33934 16174 33986
rect 16174 33934 16226 33986
rect 16226 33934 16228 33986
rect 16172 33932 16228 33934
rect 16332 33986 16388 33988
rect 16332 33934 16334 33986
rect 16334 33934 16386 33986
rect 16386 33934 16388 33986
rect 16332 33932 16388 33934
rect 16492 33986 16548 33988
rect 16492 33934 16494 33986
rect 16494 33934 16546 33986
rect 16546 33934 16548 33986
rect 16492 33932 16548 33934
rect 16652 33986 16708 33988
rect 16652 33934 16654 33986
rect 16654 33934 16706 33986
rect 16706 33934 16708 33986
rect 16652 33932 16708 33934
rect 16812 33986 16868 33988
rect 16812 33934 16814 33986
rect 16814 33934 16866 33986
rect 16866 33934 16868 33986
rect 16812 33932 16868 33934
rect 16972 33986 17028 33988
rect 16972 33934 16974 33986
rect 16974 33934 17026 33986
rect 17026 33934 17028 33986
rect 16972 33932 17028 33934
rect 17132 33986 17188 33988
rect 17132 33934 17134 33986
rect 17134 33934 17186 33986
rect 17186 33934 17188 33986
rect 17132 33932 17188 33934
rect 17292 33986 17348 33988
rect 17292 33934 17294 33986
rect 17294 33934 17346 33986
rect 17346 33934 17348 33986
rect 17292 33932 17348 33934
rect 17452 33986 17508 33988
rect 17452 33934 17454 33986
rect 17454 33934 17506 33986
rect 17506 33934 17508 33986
rect 17452 33932 17508 33934
rect 17612 33986 17668 33988
rect 17612 33934 17614 33986
rect 17614 33934 17666 33986
rect 17666 33934 17668 33986
rect 17612 33932 17668 33934
rect 17772 33986 17828 33988
rect 17772 33934 17774 33986
rect 17774 33934 17826 33986
rect 17826 33934 17828 33986
rect 17772 33932 17828 33934
rect 17932 33986 17988 33988
rect 17932 33934 17934 33986
rect 17934 33934 17986 33986
rect 17986 33934 17988 33986
rect 17932 33932 17988 33934
rect 18092 33986 18148 33988
rect 18092 33934 18094 33986
rect 18094 33934 18146 33986
rect 18146 33934 18148 33986
rect 18092 33932 18148 33934
rect 18252 33986 18308 33988
rect 18252 33934 18254 33986
rect 18254 33934 18306 33986
rect 18306 33934 18308 33986
rect 18252 33932 18308 33934
rect 18412 33986 18468 33988
rect 18412 33934 18414 33986
rect 18414 33934 18466 33986
rect 18466 33934 18468 33986
rect 18412 33932 18468 33934
rect 18572 33986 18628 33988
rect 18572 33934 18574 33986
rect 18574 33934 18626 33986
rect 18626 33934 18628 33986
rect 18572 33932 18628 33934
rect 18732 33986 18788 33988
rect 18732 33934 18734 33986
rect 18734 33934 18786 33986
rect 18786 33934 18788 33986
rect 18732 33932 18788 33934
rect 18892 33986 18948 33988
rect 18892 33934 18894 33986
rect 18894 33934 18946 33986
rect 18946 33934 18948 33986
rect 18892 33932 18948 33934
rect 19532 33932 19588 33988
rect 19852 33932 19908 33988
rect 23132 33986 23188 33988
rect 23132 33934 23134 33986
rect 23134 33934 23186 33986
rect 23186 33934 23188 33986
rect 23132 33932 23188 33934
rect 23292 33986 23348 33988
rect 23292 33934 23294 33986
rect 23294 33934 23346 33986
rect 23346 33934 23348 33986
rect 23292 33932 23348 33934
rect 23452 33986 23508 33988
rect 23452 33934 23454 33986
rect 23454 33934 23506 33986
rect 23506 33934 23508 33986
rect 23452 33932 23508 33934
rect 23612 33986 23668 33988
rect 23612 33934 23614 33986
rect 23614 33934 23666 33986
rect 23666 33934 23668 33986
rect 23612 33932 23668 33934
rect 23772 33986 23828 33988
rect 23772 33934 23774 33986
rect 23774 33934 23826 33986
rect 23826 33934 23828 33986
rect 23772 33932 23828 33934
rect 23932 33986 23988 33988
rect 23932 33934 23934 33986
rect 23934 33934 23986 33986
rect 23986 33934 23988 33986
rect 23932 33932 23988 33934
rect 24092 33986 24148 33988
rect 24092 33934 24094 33986
rect 24094 33934 24146 33986
rect 24146 33934 24148 33986
rect 24092 33932 24148 33934
rect 24252 33986 24308 33988
rect 24252 33934 24254 33986
rect 24254 33934 24306 33986
rect 24306 33934 24308 33986
rect 24252 33932 24308 33934
rect 24412 33986 24468 33988
rect 24412 33934 24414 33986
rect 24414 33934 24466 33986
rect 24466 33934 24468 33986
rect 24412 33932 24468 33934
rect 24572 33986 24628 33988
rect 24572 33934 24574 33986
rect 24574 33934 24626 33986
rect 24626 33934 24628 33986
rect 24572 33932 24628 33934
rect 24732 33986 24788 33988
rect 24732 33934 24734 33986
rect 24734 33934 24786 33986
rect 24786 33934 24788 33986
rect 24732 33932 24788 33934
rect 24892 33986 24948 33988
rect 24892 33934 24894 33986
rect 24894 33934 24946 33986
rect 24946 33934 24948 33986
rect 24892 33932 24948 33934
rect 25052 33986 25108 33988
rect 25052 33934 25054 33986
rect 25054 33934 25106 33986
rect 25106 33934 25108 33986
rect 25052 33932 25108 33934
rect 25212 33986 25268 33988
rect 25212 33934 25214 33986
rect 25214 33934 25266 33986
rect 25266 33934 25268 33986
rect 25212 33932 25268 33934
rect 25372 33986 25428 33988
rect 25372 33934 25374 33986
rect 25374 33934 25426 33986
rect 25426 33934 25428 33986
rect 25372 33932 25428 33934
rect 25532 33986 25588 33988
rect 25532 33934 25534 33986
rect 25534 33934 25586 33986
rect 25586 33934 25588 33986
rect 25532 33932 25588 33934
rect 25692 33986 25748 33988
rect 25692 33934 25694 33986
rect 25694 33934 25746 33986
rect 25746 33934 25748 33986
rect 25692 33932 25748 33934
rect 25852 33986 25908 33988
rect 25852 33934 25854 33986
rect 25854 33934 25906 33986
rect 25906 33934 25908 33986
rect 25852 33932 25908 33934
rect 26012 33986 26068 33988
rect 26012 33934 26014 33986
rect 26014 33934 26066 33986
rect 26066 33934 26068 33986
rect 26012 33932 26068 33934
rect 26172 33986 26228 33988
rect 26172 33934 26174 33986
rect 26174 33934 26226 33986
rect 26226 33934 26228 33986
rect 26172 33932 26228 33934
rect 26332 33986 26388 33988
rect 26332 33934 26334 33986
rect 26334 33934 26386 33986
rect 26386 33934 26388 33986
rect 26332 33932 26388 33934
rect 26492 33986 26548 33988
rect 26492 33934 26494 33986
rect 26494 33934 26546 33986
rect 26546 33934 26548 33986
rect 26492 33932 26548 33934
rect 26652 33986 26708 33988
rect 26652 33934 26654 33986
rect 26654 33934 26706 33986
rect 26706 33934 26708 33986
rect 26652 33932 26708 33934
rect 26812 33986 26868 33988
rect 26812 33934 26814 33986
rect 26814 33934 26866 33986
rect 26866 33934 26868 33986
rect 26812 33932 26868 33934
rect 26972 33986 27028 33988
rect 26972 33934 26974 33986
rect 26974 33934 27026 33986
rect 27026 33934 27028 33986
rect 26972 33932 27028 33934
rect 27132 33986 27188 33988
rect 27132 33934 27134 33986
rect 27134 33934 27186 33986
rect 27186 33934 27188 33986
rect 27132 33932 27188 33934
rect 27292 33986 27348 33988
rect 27292 33934 27294 33986
rect 27294 33934 27346 33986
rect 27346 33934 27348 33986
rect 27292 33932 27348 33934
rect 27452 33986 27508 33988
rect 27452 33934 27454 33986
rect 27454 33934 27506 33986
rect 27506 33934 27508 33986
rect 27452 33932 27508 33934
rect 27612 33986 27668 33988
rect 27612 33934 27614 33986
rect 27614 33934 27666 33986
rect 27666 33934 27668 33986
rect 27612 33932 27668 33934
rect 27772 33986 27828 33988
rect 27772 33934 27774 33986
rect 27774 33934 27826 33986
rect 27826 33934 27828 33986
rect 27772 33932 27828 33934
rect 27932 33986 27988 33988
rect 27932 33934 27934 33986
rect 27934 33934 27986 33986
rect 27986 33934 27988 33986
rect 27932 33932 27988 33934
rect 28092 33986 28148 33988
rect 28092 33934 28094 33986
rect 28094 33934 28146 33986
rect 28146 33934 28148 33986
rect 28092 33932 28148 33934
rect 28252 33986 28308 33988
rect 28252 33934 28254 33986
rect 28254 33934 28306 33986
rect 28306 33934 28308 33986
rect 28252 33932 28308 33934
rect 28412 33986 28468 33988
rect 28412 33934 28414 33986
rect 28414 33934 28466 33986
rect 28466 33934 28468 33986
rect 28412 33932 28468 33934
rect 28572 33986 28628 33988
rect 28572 33934 28574 33986
rect 28574 33934 28626 33986
rect 28626 33934 28628 33986
rect 28572 33932 28628 33934
rect 28732 33986 28788 33988
rect 28732 33934 28734 33986
rect 28734 33934 28786 33986
rect 28786 33934 28788 33986
rect 28732 33932 28788 33934
rect 28892 33986 28948 33988
rect 28892 33934 28894 33986
rect 28894 33934 28946 33986
rect 28946 33934 28948 33986
rect 28892 33932 28948 33934
rect 29052 33986 29108 33988
rect 29052 33934 29054 33986
rect 29054 33934 29106 33986
rect 29106 33934 29108 33986
rect 29052 33932 29108 33934
rect 29212 33986 29268 33988
rect 29212 33934 29214 33986
rect 29214 33934 29266 33986
rect 29266 33934 29268 33986
rect 29212 33932 29268 33934
rect 29372 33986 29428 33988
rect 29372 33934 29374 33986
rect 29374 33934 29426 33986
rect 29426 33934 29428 33986
rect 29372 33932 29428 33934
rect 30012 33932 30068 33988
rect 30332 33932 30388 33988
rect 33532 33986 33588 33988
rect 33532 33934 33534 33986
rect 33534 33934 33586 33986
rect 33586 33934 33588 33986
rect 33532 33932 33588 33934
rect 33692 33986 33748 33988
rect 33692 33934 33694 33986
rect 33694 33934 33746 33986
rect 33746 33934 33748 33986
rect 33692 33932 33748 33934
rect 33852 33986 33908 33988
rect 33852 33934 33854 33986
rect 33854 33934 33906 33986
rect 33906 33934 33908 33986
rect 33852 33932 33908 33934
rect 34012 33986 34068 33988
rect 34012 33934 34014 33986
rect 34014 33934 34066 33986
rect 34066 33934 34068 33986
rect 34012 33932 34068 33934
rect 34172 33986 34228 33988
rect 34172 33934 34174 33986
rect 34174 33934 34226 33986
rect 34226 33934 34228 33986
rect 34172 33932 34228 33934
rect 34332 33986 34388 33988
rect 34332 33934 34334 33986
rect 34334 33934 34386 33986
rect 34386 33934 34388 33986
rect 34332 33932 34388 33934
rect 34492 33986 34548 33988
rect 34492 33934 34494 33986
rect 34494 33934 34546 33986
rect 34546 33934 34548 33986
rect 34492 33932 34548 33934
rect 34652 33986 34708 33988
rect 34652 33934 34654 33986
rect 34654 33934 34706 33986
rect 34706 33934 34708 33986
rect 34652 33932 34708 33934
rect 34812 33986 34868 33988
rect 34812 33934 34814 33986
rect 34814 33934 34866 33986
rect 34866 33934 34868 33986
rect 34812 33932 34868 33934
rect 34972 33986 35028 33988
rect 34972 33934 34974 33986
rect 34974 33934 35026 33986
rect 35026 33934 35028 33986
rect 34972 33932 35028 33934
rect 35132 33986 35188 33988
rect 35132 33934 35134 33986
rect 35134 33934 35186 33986
rect 35186 33934 35188 33986
rect 35132 33932 35188 33934
rect 35292 33986 35348 33988
rect 35292 33934 35294 33986
rect 35294 33934 35346 33986
rect 35346 33934 35348 33986
rect 35292 33932 35348 33934
rect 35452 33986 35508 33988
rect 35452 33934 35454 33986
rect 35454 33934 35506 33986
rect 35506 33934 35508 33986
rect 35452 33932 35508 33934
rect 35612 33986 35668 33988
rect 35612 33934 35614 33986
rect 35614 33934 35666 33986
rect 35666 33934 35668 33986
rect 35612 33932 35668 33934
rect 35772 33986 35828 33988
rect 35772 33934 35774 33986
rect 35774 33934 35826 33986
rect 35826 33934 35828 33986
rect 35772 33932 35828 33934
rect 35932 33986 35988 33988
rect 35932 33934 35934 33986
rect 35934 33934 35986 33986
rect 35986 33934 35988 33986
rect 35932 33932 35988 33934
rect 36092 33986 36148 33988
rect 36092 33934 36094 33986
rect 36094 33934 36146 33986
rect 36146 33934 36148 33986
rect 36092 33932 36148 33934
rect 36252 33986 36308 33988
rect 36252 33934 36254 33986
rect 36254 33934 36306 33986
rect 36306 33934 36308 33986
rect 36252 33932 36308 33934
rect 36412 33986 36468 33988
rect 36412 33934 36414 33986
rect 36414 33934 36466 33986
rect 36466 33934 36468 33986
rect 36412 33932 36468 33934
rect 36572 33986 36628 33988
rect 36572 33934 36574 33986
rect 36574 33934 36626 33986
rect 36626 33934 36628 33986
rect 36572 33932 36628 33934
rect 36732 33986 36788 33988
rect 36732 33934 36734 33986
rect 36734 33934 36786 33986
rect 36786 33934 36788 33986
rect 36732 33932 36788 33934
rect 36892 33986 36948 33988
rect 36892 33934 36894 33986
rect 36894 33934 36946 33986
rect 36946 33934 36948 33986
rect 36892 33932 36948 33934
rect 37052 33986 37108 33988
rect 37052 33934 37054 33986
rect 37054 33934 37106 33986
rect 37106 33934 37108 33986
rect 37052 33932 37108 33934
rect 37212 33986 37268 33988
rect 37212 33934 37214 33986
rect 37214 33934 37266 33986
rect 37266 33934 37268 33986
rect 37212 33932 37268 33934
rect 37372 33986 37428 33988
rect 37372 33934 37374 33986
rect 37374 33934 37426 33986
rect 37426 33934 37428 33986
rect 37372 33932 37428 33934
rect 37532 33986 37588 33988
rect 37532 33934 37534 33986
rect 37534 33934 37586 33986
rect 37586 33934 37588 33986
rect 37532 33932 37588 33934
rect 37692 33986 37748 33988
rect 37692 33934 37694 33986
rect 37694 33934 37746 33986
rect 37746 33934 37748 33986
rect 37692 33932 37748 33934
rect 37852 33986 37908 33988
rect 37852 33934 37854 33986
rect 37854 33934 37906 33986
rect 37906 33934 37908 33986
rect 37852 33932 37908 33934
rect 38012 33986 38068 33988
rect 38012 33934 38014 33986
rect 38014 33934 38066 33986
rect 38066 33934 38068 33986
rect 38012 33932 38068 33934
rect 38172 33986 38228 33988
rect 38172 33934 38174 33986
rect 38174 33934 38226 33986
rect 38226 33934 38228 33986
rect 38172 33932 38228 33934
rect 38332 33986 38388 33988
rect 38332 33934 38334 33986
rect 38334 33934 38386 33986
rect 38386 33934 38388 33986
rect 38332 33932 38388 33934
rect 38492 33986 38548 33988
rect 38492 33934 38494 33986
rect 38494 33934 38546 33986
rect 38546 33934 38548 33986
rect 38492 33932 38548 33934
rect 38652 33986 38708 33988
rect 38652 33934 38654 33986
rect 38654 33934 38706 33986
rect 38706 33934 38708 33986
rect 38652 33932 38708 33934
rect 38812 33986 38868 33988
rect 38812 33934 38814 33986
rect 38814 33934 38866 33986
rect 38866 33934 38868 33986
rect 38812 33932 38868 33934
rect 38972 33986 39028 33988
rect 38972 33934 38974 33986
rect 38974 33934 39026 33986
rect 39026 33934 39028 33986
rect 38972 33932 39028 33934
rect 39132 33986 39188 33988
rect 39132 33934 39134 33986
rect 39134 33934 39186 33986
rect 39186 33934 39188 33986
rect 39132 33932 39188 33934
rect 39292 33986 39348 33988
rect 39292 33934 39294 33986
rect 39294 33934 39346 33986
rect 39346 33934 39348 33986
rect 39292 33932 39348 33934
rect 39452 33986 39508 33988
rect 39452 33934 39454 33986
rect 39454 33934 39506 33986
rect 39506 33934 39508 33986
rect 39452 33932 39508 33934
rect 39612 33986 39668 33988
rect 39612 33934 39614 33986
rect 39614 33934 39666 33986
rect 39666 33934 39668 33986
rect 39612 33932 39668 33934
rect 39772 33986 39828 33988
rect 39772 33934 39774 33986
rect 39774 33934 39826 33986
rect 39826 33934 39828 33986
rect 39772 33932 39828 33934
rect 39932 33986 39988 33988
rect 39932 33934 39934 33986
rect 39934 33934 39986 33986
rect 39986 33934 39988 33986
rect 39932 33932 39988 33934
rect 40092 33986 40148 33988
rect 40092 33934 40094 33986
rect 40094 33934 40146 33986
rect 40146 33934 40148 33986
rect 40092 33932 40148 33934
rect 40252 33986 40308 33988
rect 40252 33934 40254 33986
rect 40254 33934 40306 33986
rect 40306 33934 40308 33986
rect 40252 33932 40308 33934
rect 40412 33986 40468 33988
rect 40412 33934 40414 33986
rect 40414 33934 40466 33986
rect 40466 33934 40468 33986
rect 40412 33932 40468 33934
rect 40572 33986 40628 33988
rect 40572 33934 40574 33986
rect 40574 33934 40626 33986
rect 40626 33934 40628 33986
rect 40572 33932 40628 33934
rect 40732 33986 40788 33988
rect 40732 33934 40734 33986
rect 40734 33934 40786 33986
rect 40786 33934 40788 33986
rect 40732 33932 40788 33934
rect 40892 33986 40948 33988
rect 40892 33934 40894 33986
rect 40894 33934 40946 33986
rect 40946 33934 40948 33986
rect 40892 33932 40948 33934
rect 41052 33986 41108 33988
rect 41052 33934 41054 33986
rect 41054 33934 41106 33986
rect 41106 33934 41108 33986
rect 41052 33932 41108 33934
rect 41212 33986 41268 33988
rect 41212 33934 41214 33986
rect 41214 33934 41266 33986
rect 41266 33934 41268 33986
rect 41212 33932 41268 33934
rect 41372 33986 41428 33988
rect 41372 33934 41374 33986
rect 41374 33934 41426 33986
rect 41426 33934 41428 33986
rect 41372 33932 41428 33934
rect 41532 33986 41588 33988
rect 41532 33934 41534 33986
rect 41534 33934 41586 33986
rect 41586 33934 41588 33986
rect 41532 33932 41588 33934
rect 41692 33986 41748 33988
rect 41692 33934 41694 33986
rect 41694 33934 41746 33986
rect 41746 33934 41748 33986
rect 41692 33932 41748 33934
rect 41852 33986 41908 33988
rect 41852 33934 41854 33986
rect 41854 33934 41906 33986
rect 41906 33934 41908 33986
rect 41852 33932 41908 33934
rect 12 33826 68 33828
rect 12 33774 14 33826
rect 14 33774 66 33826
rect 66 33774 68 33826
rect 12 33772 68 33774
rect 172 33826 228 33828
rect 172 33774 174 33826
rect 174 33774 226 33826
rect 226 33774 228 33826
rect 172 33772 228 33774
rect 332 33826 388 33828
rect 332 33774 334 33826
rect 334 33774 386 33826
rect 386 33774 388 33826
rect 332 33772 388 33774
rect 492 33826 548 33828
rect 492 33774 494 33826
rect 494 33774 546 33826
rect 546 33774 548 33826
rect 492 33772 548 33774
rect 652 33826 708 33828
rect 652 33774 654 33826
rect 654 33774 706 33826
rect 706 33774 708 33826
rect 652 33772 708 33774
rect 812 33826 868 33828
rect 812 33774 814 33826
rect 814 33774 866 33826
rect 866 33774 868 33826
rect 812 33772 868 33774
rect 972 33826 1028 33828
rect 972 33774 974 33826
rect 974 33774 1026 33826
rect 1026 33774 1028 33826
rect 972 33772 1028 33774
rect 1132 33826 1188 33828
rect 1132 33774 1134 33826
rect 1134 33774 1186 33826
rect 1186 33774 1188 33826
rect 1132 33772 1188 33774
rect 1292 33826 1348 33828
rect 1292 33774 1294 33826
rect 1294 33774 1346 33826
rect 1346 33774 1348 33826
rect 1292 33772 1348 33774
rect 1452 33826 1508 33828
rect 1452 33774 1454 33826
rect 1454 33774 1506 33826
rect 1506 33774 1508 33826
rect 1452 33772 1508 33774
rect 1612 33826 1668 33828
rect 1612 33774 1614 33826
rect 1614 33774 1666 33826
rect 1666 33774 1668 33826
rect 1612 33772 1668 33774
rect 1772 33826 1828 33828
rect 1772 33774 1774 33826
rect 1774 33774 1826 33826
rect 1826 33774 1828 33826
rect 1772 33772 1828 33774
rect 1932 33826 1988 33828
rect 1932 33774 1934 33826
rect 1934 33774 1986 33826
rect 1986 33774 1988 33826
rect 1932 33772 1988 33774
rect 2092 33826 2148 33828
rect 2092 33774 2094 33826
rect 2094 33774 2146 33826
rect 2146 33774 2148 33826
rect 2092 33772 2148 33774
rect 2252 33826 2308 33828
rect 2252 33774 2254 33826
rect 2254 33774 2306 33826
rect 2306 33774 2308 33826
rect 2252 33772 2308 33774
rect 2412 33826 2468 33828
rect 2412 33774 2414 33826
rect 2414 33774 2466 33826
rect 2466 33774 2468 33826
rect 2412 33772 2468 33774
rect 2572 33826 2628 33828
rect 2572 33774 2574 33826
rect 2574 33774 2626 33826
rect 2626 33774 2628 33826
rect 2572 33772 2628 33774
rect 2732 33826 2788 33828
rect 2732 33774 2734 33826
rect 2734 33774 2786 33826
rect 2786 33774 2788 33826
rect 2732 33772 2788 33774
rect 2892 33826 2948 33828
rect 2892 33774 2894 33826
rect 2894 33774 2946 33826
rect 2946 33774 2948 33826
rect 2892 33772 2948 33774
rect 3052 33826 3108 33828
rect 3052 33774 3054 33826
rect 3054 33774 3106 33826
rect 3106 33774 3108 33826
rect 3052 33772 3108 33774
rect 3212 33826 3268 33828
rect 3212 33774 3214 33826
rect 3214 33774 3266 33826
rect 3266 33774 3268 33826
rect 3212 33772 3268 33774
rect 3372 33826 3428 33828
rect 3372 33774 3374 33826
rect 3374 33774 3426 33826
rect 3426 33774 3428 33826
rect 3372 33772 3428 33774
rect 3532 33826 3588 33828
rect 3532 33774 3534 33826
rect 3534 33774 3586 33826
rect 3586 33774 3588 33826
rect 3532 33772 3588 33774
rect 3692 33826 3748 33828
rect 3692 33774 3694 33826
rect 3694 33774 3746 33826
rect 3746 33774 3748 33826
rect 3692 33772 3748 33774
rect 3852 33826 3908 33828
rect 3852 33774 3854 33826
rect 3854 33774 3906 33826
rect 3906 33774 3908 33826
rect 3852 33772 3908 33774
rect 4012 33826 4068 33828
rect 4012 33774 4014 33826
rect 4014 33774 4066 33826
rect 4066 33774 4068 33826
rect 4012 33772 4068 33774
rect 4172 33826 4228 33828
rect 4172 33774 4174 33826
rect 4174 33774 4226 33826
rect 4226 33774 4228 33826
rect 4172 33772 4228 33774
rect 4332 33826 4388 33828
rect 4332 33774 4334 33826
rect 4334 33774 4386 33826
rect 4386 33774 4388 33826
rect 4332 33772 4388 33774
rect 4492 33826 4548 33828
rect 4492 33774 4494 33826
rect 4494 33774 4546 33826
rect 4546 33774 4548 33826
rect 4492 33772 4548 33774
rect 4652 33826 4708 33828
rect 4652 33774 4654 33826
rect 4654 33774 4706 33826
rect 4706 33774 4708 33826
rect 4652 33772 4708 33774
rect 4812 33826 4868 33828
rect 4812 33774 4814 33826
rect 4814 33774 4866 33826
rect 4866 33774 4868 33826
rect 4812 33772 4868 33774
rect 4972 33826 5028 33828
rect 4972 33774 4974 33826
rect 4974 33774 5026 33826
rect 5026 33774 5028 33826
rect 4972 33772 5028 33774
rect 5132 33826 5188 33828
rect 5132 33774 5134 33826
rect 5134 33774 5186 33826
rect 5186 33774 5188 33826
rect 5132 33772 5188 33774
rect 5292 33826 5348 33828
rect 5292 33774 5294 33826
rect 5294 33774 5346 33826
rect 5346 33774 5348 33826
rect 5292 33772 5348 33774
rect 5452 33826 5508 33828
rect 5452 33774 5454 33826
rect 5454 33774 5506 33826
rect 5506 33774 5508 33826
rect 5452 33772 5508 33774
rect 5612 33826 5668 33828
rect 5612 33774 5614 33826
rect 5614 33774 5666 33826
rect 5666 33774 5668 33826
rect 5612 33772 5668 33774
rect 5772 33826 5828 33828
rect 5772 33774 5774 33826
rect 5774 33774 5826 33826
rect 5826 33774 5828 33826
rect 5772 33772 5828 33774
rect 5932 33826 5988 33828
rect 5932 33774 5934 33826
rect 5934 33774 5986 33826
rect 5986 33774 5988 33826
rect 5932 33772 5988 33774
rect 6092 33826 6148 33828
rect 6092 33774 6094 33826
rect 6094 33774 6146 33826
rect 6146 33774 6148 33826
rect 6092 33772 6148 33774
rect 6252 33826 6308 33828
rect 6252 33774 6254 33826
rect 6254 33774 6306 33826
rect 6306 33774 6308 33826
rect 6252 33772 6308 33774
rect 6412 33826 6468 33828
rect 6412 33774 6414 33826
rect 6414 33774 6466 33826
rect 6466 33774 6468 33826
rect 6412 33772 6468 33774
rect 6572 33826 6628 33828
rect 6572 33774 6574 33826
rect 6574 33774 6626 33826
rect 6626 33774 6628 33826
rect 6572 33772 6628 33774
rect 6732 33826 6788 33828
rect 6732 33774 6734 33826
rect 6734 33774 6786 33826
rect 6786 33774 6788 33826
rect 6732 33772 6788 33774
rect 6892 33826 6948 33828
rect 6892 33774 6894 33826
rect 6894 33774 6946 33826
rect 6946 33774 6948 33826
rect 6892 33772 6948 33774
rect 7052 33826 7108 33828
rect 7052 33774 7054 33826
rect 7054 33774 7106 33826
rect 7106 33774 7108 33826
rect 7052 33772 7108 33774
rect 7212 33826 7268 33828
rect 7212 33774 7214 33826
rect 7214 33774 7266 33826
rect 7266 33774 7268 33826
rect 7212 33772 7268 33774
rect 7372 33826 7428 33828
rect 7372 33774 7374 33826
rect 7374 33774 7426 33826
rect 7426 33774 7428 33826
rect 7372 33772 7428 33774
rect 7532 33826 7588 33828
rect 7532 33774 7534 33826
rect 7534 33774 7586 33826
rect 7586 33774 7588 33826
rect 7532 33772 7588 33774
rect 7692 33826 7748 33828
rect 7692 33774 7694 33826
rect 7694 33774 7746 33826
rect 7746 33774 7748 33826
rect 7692 33772 7748 33774
rect 7852 33826 7908 33828
rect 7852 33774 7854 33826
rect 7854 33774 7906 33826
rect 7906 33774 7908 33826
rect 7852 33772 7908 33774
rect 8012 33826 8068 33828
rect 8012 33774 8014 33826
rect 8014 33774 8066 33826
rect 8066 33774 8068 33826
rect 8012 33772 8068 33774
rect 8172 33826 8228 33828
rect 8172 33774 8174 33826
rect 8174 33774 8226 33826
rect 8226 33774 8228 33826
rect 8172 33772 8228 33774
rect 8332 33826 8388 33828
rect 8332 33774 8334 33826
rect 8334 33774 8386 33826
rect 8386 33774 8388 33826
rect 8332 33772 8388 33774
rect 12012 33772 12068 33828
rect 12332 33772 12388 33828
rect 12492 33826 12548 33828
rect 12492 33774 12494 33826
rect 12494 33774 12546 33826
rect 12546 33774 12548 33826
rect 12492 33772 12548 33774
rect 12652 33826 12708 33828
rect 12652 33774 12654 33826
rect 12654 33774 12706 33826
rect 12706 33774 12708 33826
rect 12652 33772 12708 33774
rect 12812 33826 12868 33828
rect 12812 33774 12814 33826
rect 12814 33774 12866 33826
rect 12866 33774 12868 33826
rect 12812 33772 12868 33774
rect 12972 33826 13028 33828
rect 12972 33774 12974 33826
rect 12974 33774 13026 33826
rect 13026 33774 13028 33826
rect 12972 33772 13028 33774
rect 13132 33826 13188 33828
rect 13132 33774 13134 33826
rect 13134 33774 13186 33826
rect 13186 33774 13188 33826
rect 13132 33772 13188 33774
rect 13292 33826 13348 33828
rect 13292 33774 13294 33826
rect 13294 33774 13346 33826
rect 13346 33774 13348 33826
rect 13292 33772 13348 33774
rect 13452 33826 13508 33828
rect 13452 33774 13454 33826
rect 13454 33774 13506 33826
rect 13506 33774 13508 33826
rect 13452 33772 13508 33774
rect 13612 33826 13668 33828
rect 13612 33774 13614 33826
rect 13614 33774 13666 33826
rect 13666 33774 13668 33826
rect 13612 33772 13668 33774
rect 13772 33826 13828 33828
rect 13772 33774 13774 33826
rect 13774 33774 13826 33826
rect 13826 33774 13828 33826
rect 13772 33772 13828 33774
rect 13932 33826 13988 33828
rect 13932 33774 13934 33826
rect 13934 33774 13986 33826
rect 13986 33774 13988 33826
rect 13932 33772 13988 33774
rect 14092 33826 14148 33828
rect 14092 33774 14094 33826
rect 14094 33774 14146 33826
rect 14146 33774 14148 33826
rect 14092 33772 14148 33774
rect 14252 33826 14308 33828
rect 14252 33774 14254 33826
rect 14254 33774 14306 33826
rect 14306 33774 14308 33826
rect 14252 33772 14308 33774
rect 14412 33826 14468 33828
rect 14412 33774 14414 33826
rect 14414 33774 14466 33826
rect 14466 33774 14468 33826
rect 14412 33772 14468 33774
rect 14572 33826 14628 33828
rect 14572 33774 14574 33826
rect 14574 33774 14626 33826
rect 14626 33774 14628 33826
rect 14572 33772 14628 33774
rect 14732 33826 14788 33828
rect 14732 33774 14734 33826
rect 14734 33774 14786 33826
rect 14786 33774 14788 33826
rect 14732 33772 14788 33774
rect 14892 33826 14948 33828
rect 14892 33774 14894 33826
rect 14894 33774 14946 33826
rect 14946 33774 14948 33826
rect 14892 33772 14948 33774
rect 15052 33826 15108 33828
rect 15052 33774 15054 33826
rect 15054 33774 15106 33826
rect 15106 33774 15108 33826
rect 15052 33772 15108 33774
rect 15212 33826 15268 33828
rect 15212 33774 15214 33826
rect 15214 33774 15266 33826
rect 15266 33774 15268 33826
rect 15212 33772 15268 33774
rect 15372 33826 15428 33828
rect 15372 33774 15374 33826
rect 15374 33774 15426 33826
rect 15426 33774 15428 33826
rect 15372 33772 15428 33774
rect 15532 33826 15588 33828
rect 15532 33774 15534 33826
rect 15534 33774 15586 33826
rect 15586 33774 15588 33826
rect 15532 33772 15588 33774
rect 15692 33826 15748 33828
rect 15692 33774 15694 33826
rect 15694 33774 15746 33826
rect 15746 33774 15748 33826
rect 15692 33772 15748 33774
rect 15852 33826 15908 33828
rect 15852 33774 15854 33826
rect 15854 33774 15906 33826
rect 15906 33774 15908 33826
rect 15852 33772 15908 33774
rect 16012 33826 16068 33828
rect 16012 33774 16014 33826
rect 16014 33774 16066 33826
rect 16066 33774 16068 33826
rect 16012 33772 16068 33774
rect 16172 33826 16228 33828
rect 16172 33774 16174 33826
rect 16174 33774 16226 33826
rect 16226 33774 16228 33826
rect 16172 33772 16228 33774
rect 16332 33826 16388 33828
rect 16332 33774 16334 33826
rect 16334 33774 16386 33826
rect 16386 33774 16388 33826
rect 16332 33772 16388 33774
rect 16492 33826 16548 33828
rect 16492 33774 16494 33826
rect 16494 33774 16546 33826
rect 16546 33774 16548 33826
rect 16492 33772 16548 33774
rect 16652 33826 16708 33828
rect 16652 33774 16654 33826
rect 16654 33774 16706 33826
rect 16706 33774 16708 33826
rect 16652 33772 16708 33774
rect 16812 33826 16868 33828
rect 16812 33774 16814 33826
rect 16814 33774 16866 33826
rect 16866 33774 16868 33826
rect 16812 33772 16868 33774
rect 16972 33826 17028 33828
rect 16972 33774 16974 33826
rect 16974 33774 17026 33826
rect 17026 33774 17028 33826
rect 16972 33772 17028 33774
rect 17132 33826 17188 33828
rect 17132 33774 17134 33826
rect 17134 33774 17186 33826
rect 17186 33774 17188 33826
rect 17132 33772 17188 33774
rect 17292 33826 17348 33828
rect 17292 33774 17294 33826
rect 17294 33774 17346 33826
rect 17346 33774 17348 33826
rect 17292 33772 17348 33774
rect 17452 33826 17508 33828
rect 17452 33774 17454 33826
rect 17454 33774 17506 33826
rect 17506 33774 17508 33826
rect 17452 33772 17508 33774
rect 17612 33826 17668 33828
rect 17612 33774 17614 33826
rect 17614 33774 17666 33826
rect 17666 33774 17668 33826
rect 17612 33772 17668 33774
rect 17772 33826 17828 33828
rect 17772 33774 17774 33826
rect 17774 33774 17826 33826
rect 17826 33774 17828 33826
rect 17772 33772 17828 33774
rect 17932 33826 17988 33828
rect 17932 33774 17934 33826
rect 17934 33774 17986 33826
rect 17986 33774 17988 33826
rect 17932 33772 17988 33774
rect 18092 33826 18148 33828
rect 18092 33774 18094 33826
rect 18094 33774 18146 33826
rect 18146 33774 18148 33826
rect 18092 33772 18148 33774
rect 18252 33826 18308 33828
rect 18252 33774 18254 33826
rect 18254 33774 18306 33826
rect 18306 33774 18308 33826
rect 18252 33772 18308 33774
rect 18412 33826 18468 33828
rect 18412 33774 18414 33826
rect 18414 33774 18466 33826
rect 18466 33774 18468 33826
rect 18412 33772 18468 33774
rect 18572 33826 18628 33828
rect 18572 33774 18574 33826
rect 18574 33774 18626 33826
rect 18626 33774 18628 33826
rect 18572 33772 18628 33774
rect 18732 33826 18788 33828
rect 18732 33774 18734 33826
rect 18734 33774 18786 33826
rect 18786 33774 18788 33826
rect 18732 33772 18788 33774
rect 18892 33826 18948 33828
rect 18892 33774 18894 33826
rect 18894 33774 18946 33826
rect 18946 33774 18948 33826
rect 18892 33772 18948 33774
rect 19052 33772 19108 33828
rect 19372 33772 19428 33828
rect 23132 33826 23188 33828
rect 23132 33774 23134 33826
rect 23134 33774 23186 33826
rect 23186 33774 23188 33826
rect 23132 33772 23188 33774
rect 23292 33826 23348 33828
rect 23292 33774 23294 33826
rect 23294 33774 23346 33826
rect 23346 33774 23348 33826
rect 23292 33772 23348 33774
rect 23452 33826 23508 33828
rect 23452 33774 23454 33826
rect 23454 33774 23506 33826
rect 23506 33774 23508 33826
rect 23452 33772 23508 33774
rect 23612 33826 23668 33828
rect 23612 33774 23614 33826
rect 23614 33774 23666 33826
rect 23666 33774 23668 33826
rect 23612 33772 23668 33774
rect 23772 33826 23828 33828
rect 23772 33774 23774 33826
rect 23774 33774 23826 33826
rect 23826 33774 23828 33826
rect 23772 33772 23828 33774
rect 23932 33826 23988 33828
rect 23932 33774 23934 33826
rect 23934 33774 23986 33826
rect 23986 33774 23988 33826
rect 23932 33772 23988 33774
rect 24092 33826 24148 33828
rect 24092 33774 24094 33826
rect 24094 33774 24146 33826
rect 24146 33774 24148 33826
rect 24092 33772 24148 33774
rect 24252 33826 24308 33828
rect 24252 33774 24254 33826
rect 24254 33774 24306 33826
rect 24306 33774 24308 33826
rect 24252 33772 24308 33774
rect 24412 33826 24468 33828
rect 24412 33774 24414 33826
rect 24414 33774 24466 33826
rect 24466 33774 24468 33826
rect 24412 33772 24468 33774
rect 24572 33826 24628 33828
rect 24572 33774 24574 33826
rect 24574 33774 24626 33826
rect 24626 33774 24628 33826
rect 24572 33772 24628 33774
rect 24732 33826 24788 33828
rect 24732 33774 24734 33826
rect 24734 33774 24786 33826
rect 24786 33774 24788 33826
rect 24732 33772 24788 33774
rect 24892 33826 24948 33828
rect 24892 33774 24894 33826
rect 24894 33774 24946 33826
rect 24946 33774 24948 33826
rect 24892 33772 24948 33774
rect 25052 33826 25108 33828
rect 25052 33774 25054 33826
rect 25054 33774 25106 33826
rect 25106 33774 25108 33826
rect 25052 33772 25108 33774
rect 25212 33826 25268 33828
rect 25212 33774 25214 33826
rect 25214 33774 25266 33826
rect 25266 33774 25268 33826
rect 25212 33772 25268 33774
rect 25372 33826 25428 33828
rect 25372 33774 25374 33826
rect 25374 33774 25426 33826
rect 25426 33774 25428 33826
rect 25372 33772 25428 33774
rect 25532 33826 25588 33828
rect 25532 33774 25534 33826
rect 25534 33774 25586 33826
rect 25586 33774 25588 33826
rect 25532 33772 25588 33774
rect 25692 33826 25748 33828
rect 25692 33774 25694 33826
rect 25694 33774 25746 33826
rect 25746 33774 25748 33826
rect 25692 33772 25748 33774
rect 25852 33826 25908 33828
rect 25852 33774 25854 33826
rect 25854 33774 25906 33826
rect 25906 33774 25908 33826
rect 25852 33772 25908 33774
rect 26012 33826 26068 33828
rect 26012 33774 26014 33826
rect 26014 33774 26066 33826
rect 26066 33774 26068 33826
rect 26012 33772 26068 33774
rect 26172 33826 26228 33828
rect 26172 33774 26174 33826
rect 26174 33774 26226 33826
rect 26226 33774 26228 33826
rect 26172 33772 26228 33774
rect 26332 33826 26388 33828
rect 26332 33774 26334 33826
rect 26334 33774 26386 33826
rect 26386 33774 26388 33826
rect 26332 33772 26388 33774
rect 26492 33826 26548 33828
rect 26492 33774 26494 33826
rect 26494 33774 26546 33826
rect 26546 33774 26548 33826
rect 26492 33772 26548 33774
rect 26652 33826 26708 33828
rect 26652 33774 26654 33826
rect 26654 33774 26706 33826
rect 26706 33774 26708 33826
rect 26652 33772 26708 33774
rect 26812 33826 26868 33828
rect 26812 33774 26814 33826
rect 26814 33774 26866 33826
rect 26866 33774 26868 33826
rect 26812 33772 26868 33774
rect 26972 33826 27028 33828
rect 26972 33774 26974 33826
rect 26974 33774 27026 33826
rect 27026 33774 27028 33826
rect 26972 33772 27028 33774
rect 27132 33826 27188 33828
rect 27132 33774 27134 33826
rect 27134 33774 27186 33826
rect 27186 33774 27188 33826
rect 27132 33772 27188 33774
rect 27292 33826 27348 33828
rect 27292 33774 27294 33826
rect 27294 33774 27346 33826
rect 27346 33774 27348 33826
rect 27292 33772 27348 33774
rect 27452 33826 27508 33828
rect 27452 33774 27454 33826
rect 27454 33774 27506 33826
rect 27506 33774 27508 33826
rect 27452 33772 27508 33774
rect 27612 33826 27668 33828
rect 27612 33774 27614 33826
rect 27614 33774 27666 33826
rect 27666 33774 27668 33826
rect 27612 33772 27668 33774
rect 27772 33826 27828 33828
rect 27772 33774 27774 33826
rect 27774 33774 27826 33826
rect 27826 33774 27828 33826
rect 27772 33772 27828 33774
rect 27932 33826 27988 33828
rect 27932 33774 27934 33826
rect 27934 33774 27986 33826
rect 27986 33774 27988 33826
rect 27932 33772 27988 33774
rect 28092 33826 28148 33828
rect 28092 33774 28094 33826
rect 28094 33774 28146 33826
rect 28146 33774 28148 33826
rect 28092 33772 28148 33774
rect 28252 33826 28308 33828
rect 28252 33774 28254 33826
rect 28254 33774 28306 33826
rect 28306 33774 28308 33826
rect 28252 33772 28308 33774
rect 28412 33826 28468 33828
rect 28412 33774 28414 33826
rect 28414 33774 28466 33826
rect 28466 33774 28468 33826
rect 28412 33772 28468 33774
rect 28572 33826 28628 33828
rect 28572 33774 28574 33826
rect 28574 33774 28626 33826
rect 28626 33774 28628 33826
rect 28572 33772 28628 33774
rect 28732 33826 28788 33828
rect 28732 33774 28734 33826
rect 28734 33774 28786 33826
rect 28786 33774 28788 33826
rect 28732 33772 28788 33774
rect 28892 33826 28948 33828
rect 28892 33774 28894 33826
rect 28894 33774 28946 33826
rect 28946 33774 28948 33826
rect 28892 33772 28948 33774
rect 29052 33826 29108 33828
rect 29052 33774 29054 33826
rect 29054 33774 29106 33826
rect 29106 33774 29108 33826
rect 29052 33772 29108 33774
rect 29212 33826 29268 33828
rect 29212 33774 29214 33826
rect 29214 33774 29266 33826
rect 29266 33774 29268 33826
rect 29212 33772 29268 33774
rect 29372 33826 29428 33828
rect 29372 33774 29374 33826
rect 29374 33774 29426 33826
rect 29426 33774 29428 33826
rect 29372 33772 29428 33774
rect 29532 33772 29588 33828
rect 29852 33772 29908 33828
rect 33532 33826 33588 33828
rect 33532 33774 33534 33826
rect 33534 33774 33586 33826
rect 33586 33774 33588 33826
rect 33532 33772 33588 33774
rect 33692 33826 33748 33828
rect 33692 33774 33694 33826
rect 33694 33774 33746 33826
rect 33746 33774 33748 33826
rect 33692 33772 33748 33774
rect 33852 33826 33908 33828
rect 33852 33774 33854 33826
rect 33854 33774 33906 33826
rect 33906 33774 33908 33826
rect 33852 33772 33908 33774
rect 34012 33826 34068 33828
rect 34012 33774 34014 33826
rect 34014 33774 34066 33826
rect 34066 33774 34068 33826
rect 34012 33772 34068 33774
rect 34172 33826 34228 33828
rect 34172 33774 34174 33826
rect 34174 33774 34226 33826
rect 34226 33774 34228 33826
rect 34172 33772 34228 33774
rect 34332 33826 34388 33828
rect 34332 33774 34334 33826
rect 34334 33774 34386 33826
rect 34386 33774 34388 33826
rect 34332 33772 34388 33774
rect 34492 33826 34548 33828
rect 34492 33774 34494 33826
rect 34494 33774 34546 33826
rect 34546 33774 34548 33826
rect 34492 33772 34548 33774
rect 34652 33826 34708 33828
rect 34652 33774 34654 33826
rect 34654 33774 34706 33826
rect 34706 33774 34708 33826
rect 34652 33772 34708 33774
rect 34812 33826 34868 33828
rect 34812 33774 34814 33826
rect 34814 33774 34866 33826
rect 34866 33774 34868 33826
rect 34812 33772 34868 33774
rect 34972 33826 35028 33828
rect 34972 33774 34974 33826
rect 34974 33774 35026 33826
rect 35026 33774 35028 33826
rect 34972 33772 35028 33774
rect 35132 33826 35188 33828
rect 35132 33774 35134 33826
rect 35134 33774 35186 33826
rect 35186 33774 35188 33826
rect 35132 33772 35188 33774
rect 35292 33826 35348 33828
rect 35292 33774 35294 33826
rect 35294 33774 35346 33826
rect 35346 33774 35348 33826
rect 35292 33772 35348 33774
rect 35452 33826 35508 33828
rect 35452 33774 35454 33826
rect 35454 33774 35506 33826
rect 35506 33774 35508 33826
rect 35452 33772 35508 33774
rect 35612 33826 35668 33828
rect 35612 33774 35614 33826
rect 35614 33774 35666 33826
rect 35666 33774 35668 33826
rect 35612 33772 35668 33774
rect 35772 33826 35828 33828
rect 35772 33774 35774 33826
rect 35774 33774 35826 33826
rect 35826 33774 35828 33826
rect 35772 33772 35828 33774
rect 35932 33826 35988 33828
rect 35932 33774 35934 33826
rect 35934 33774 35986 33826
rect 35986 33774 35988 33826
rect 35932 33772 35988 33774
rect 36092 33826 36148 33828
rect 36092 33774 36094 33826
rect 36094 33774 36146 33826
rect 36146 33774 36148 33826
rect 36092 33772 36148 33774
rect 36252 33826 36308 33828
rect 36252 33774 36254 33826
rect 36254 33774 36306 33826
rect 36306 33774 36308 33826
rect 36252 33772 36308 33774
rect 36412 33826 36468 33828
rect 36412 33774 36414 33826
rect 36414 33774 36466 33826
rect 36466 33774 36468 33826
rect 36412 33772 36468 33774
rect 36572 33826 36628 33828
rect 36572 33774 36574 33826
rect 36574 33774 36626 33826
rect 36626 33774 36628 33826
rect 36572 33772 36628 33774
rect 36732 33826 36788 33828
rect 36732 33774 36734 33826
rect 36734 33774 36786 33826
rect 36786 33774 36788 33826
rect 36732 33772 36788 33774
rect 36892 33826 36948 33828
rect 36892 33774 36894 33826
rect 36894 33774 36946 33826
rect 36946 33774 36948 33826
rect 36892 33772 36948 33774
rect 37052 33826 37108 33828
rect 37052 33774 37054 33826
rect 37054 33774 37106 33826
rect 37106 33774 37108 33826
rect 37052 33772 37108 33774
rect 37212 33826 37268 33828
rect 37212 33774 37214 33826
rect 37214 33774 37266 33826
rect 37266 33774 37268 33826
rect 37212 33772 37268 33774
rect 37372 33826 37428 33828
rect 37372 33774 37374 33826
rect 37374 33774 37426 33826
rect 37426 33774 37428 33826
rect 37372 33772 37428 33774
rect 37532 33826 37588 33828
rect 37532 33774 37534 33826
rect 37534 33774 37586 33826
rect 37586 33774 37588 33826
rect 37532 33772 37588 33774
rect 37692 33826 37748 33828
rect 37692 33774 37694 33826
rect 37694 33774 37746 33826
rect 37746 33774 37748 33826
rect 37692 33772 37748 33774
rect 37852 33826 37908 33828
rect 37852 33774 37854 33826
rect 37854 33774 37906 33826
rect 37906 33774 37908 33826
rect 37852 33772 37908 33774
rect 38012 33826 38068 33828
rect 38012 33774 38014 33826
rect 38014 33774 38066 33826
rect 38066 33774 38068 33826
rect 38012 33772 38068 33774
rect 38172 33826 38228 33828
rect 38172 33774 38174 33826
rect 38174 33774 38226 33826
rect 38226 33774 38228 33826
rect 38172 33772 38228 33774
rect 38332 33826 38388 33828
rect 38332 33774 38334 33826
rect 38334 33774 38386 33826
rect 38386 33774 38388 33826
rect 38332 33772 38388 33774
rect 38492 33826 38548 33828
rect 38492 33774 38494 33826
rect 38494 33774 38546 33826
rect 38546 33774 38548 33826
rect 38492 33772 38548 33774
rect 38652 33826 38708 33828
rect 38652 33774 38654 33826
rect 38654 33774 38706 33826
rect 38706 33774 38708 33826
rect 38652 33772 38708 33774
rect 38812 33826 38868 33828
rect 38812 33774 38814 33826
rect 38814 33774 38866 33826
rect 38866 33774 38868 33826
rect 38812 33772 38868 33774
rect 38972 33826 39028 33828
rect 38972 33774 38974 33826
rect 38974 33774 39026 33826
rect 39026 33774 39028 33826
rect 38972 33772 39028 33774
rect 39132 33826 39188 33828
rect 39132 33774 39134 33826
rect 39134 33774 39186 33826
rect 39186 33774 39188 33826
rect 39132 33772 39188 33774
rect 39292 33826 39348 33828
rect 39292 33774 39294 33826
rect 39294 33774 39346 33826
rect 39346 33774 39348 33826
rect 39292 33772 39348 33774
rect 39452 33826 39508 33828
rect 39452 33774 39454 33826
rect 39454 33774 39506 33826
rect 39506 33774 39508 33826
rect 39452 33772 39508 33774
rect 39612 33826 39668 33828
rect 39612 33774 39614 33826
rect 39614 33774 39666 33826
rect 39666 33774 39668 33826
rect 39612 33772 39668 33774
rect 39772 33826 39828 33828
rect 39772 33774 39774 33826
rect 39774 33774 39826 33826
rect 39826 33774 39828 33826
rect 39772 33772 39828 33774
rect 39932 33826 39988 33828
rect 39932 33774 39934 33826
rect 39934 33774 39986 33826
rect 39986 33774 39988 33826
rect 39932 33772 39988 33774
rect 40092 33826 40148 33828
rect 40092 33774 40094 33826
rect 40094 33774 40146 33826
rect 40146 33774 40148 33826
rect 40092 33772 40148 33774
rect 40252 33826 40308 33828
rect 40252 33774 40254 33826
rect 40254 33774 40306 33826
rect 40306 33774 40308 33826
rect 40252 33772 40308 33774
rect 40412 33826 40468 33828
rect 40412 33774 40414 33826
rect 40414 33774 40466 33826
rect 40466 33774 40468 33826
rect 40412 33772 40468 33774
rect 40572 33826 40628 33828
rect 40572 33774 40574 33826
rect 40574 33774 40626 33826
rect 40626 33774 40628 33826
rect 40572 33772 40628 33774
rect 40732 33826 40788 33828
rect 40732 33774 40734 33826
rect 40734 33774 40786 33826
rect 40786 33774 40788 33826
rect 40732 33772 40788 33774
rect 40892 33826 40948 33828
rect 40892 33774 40894 33826
rect 40894 33774 40946 33826
rect 40946 33774 40948 33826
rect 40892 33772 40948 33774
rect 41052 33826 41108 33828
rect 41052 33774 41054 33826
rect 41054 33774 41106 33826
rect 41106 33774 41108 33826
rect 41052 33772 41108 33774
rect 41212 33826 41268 33828
rect 41212 33774 41214 33826
rect 41214 33774 41266 33826
rect 41266 33774 41268 33826
rect 41212 33772 41268 33774
rect 41372 33826 41428 33828
rect 41372 33774 41374 33826
rect 41374 33774 41426 33826
rect 41426 33774 41428 33826
rect 41372 33772 41428 33774
rect 41532 33826 41588 33828
rect 41532 33774 41534 33826
rect 41534 33774 41586 33826
rect 41586 33774 41588 33826
rect 41532 33772 41588 33774
rect 41692 33826 41748 33828
rect 41692 33774 41694 33826
rect 41694 33774 41746 33826
rect 41746 33774 41748 33826
rect 41692 33772 41748 33774
rect 41852 33826 41908 33828
rect 41852 33774 41854 33826
rect 41854 33774 41906 33826
rect 41906 33774 41908 33826
rect 41852 33772 41908 33774
rect 12172 33612 12228 33668
rect 19212 33612 19268 33668
rect 29692 33612 29748 33668
rect 12 33506 68 33508
rect 12 33454 14 33506
rect 14 33454 66 33506
rect 66 33454 68 33506
rect 12 33452 68 33454
rect 172 33506 228 33508
rect 172 33454 174 33506
rect 174 33454 226 33506
rect 226 33454 228 33506
rect 172 33452 228 33454
rect 332 33506 388 33508
rect 332 33454 334 33506
rect 334 33454 386 33506
rect 386 33454 388 33506
rect 332 33452 388 33454
rect 492 33506 548 33508
rect 492 33454 494 33506
rect 494 33454 546 33506
rect 546 33454 548 33506
rect 492 33452 548 33454
rect 652 33506 708 33508
rect 652 33454 654 33506
rect 654 33454 706 33506
rect 706 33454 708 33506
rect 652 33452 708 33454
rect 812 33506 868 33508
rect 812 33454 814 33506
rect 814 33454 866 33506
rect 866 33454 868 33506
rect 812 33452 868 33454
rect 972 33506 1028 33508
rect 972 33454 974 33506
rect 974 33454 1026 33506
rect 1026 33454 1028 33506
rect 972 33452 1028 33454
rect 1132 33506 1188 33508
rect 1132 33454 1134 33506
rect 1134 33454 1186 33506
rect 1186 33454 1188 33506
rect 1132 33452 1188 33454
rect 1292 33506 1348 33508
rect 1292 33454 1294 33506
rect 1294 33454 1346 33506
rect 1346 33454 1348 33506
rect 1292 33452 1348 33454
rect 1452 33506 1508 33508
rect 1452 33454 1454 33506
rect 1454 33454 1506 33506
rect 1506 33454 1508 33506
rect 1452 33452 1508 33454
rect 1612 33506 1668 33508
rect 1612 33454 1614 33506
rect 1614 33454 1666 33506
rect 1666 33454 1668 33506
rect 1612 33452 1668 33454
rect 1772 33506 1828 33508
rect 1772 33454 1774 33506
rect 1774 33454 1826 33506
rect 1826 33454 1828 33506
rect 1772 33452 1828 33454
rect 1932 33506 1988 33508
rect 1932 33454 1934 33506
rect 1934 33454 1986 33506
rect 1986 33454 1988 33506
rect 1932 33452 1988 33454
rect 2092 33506 2148 33508
rect 2092 33454 2094 33506
rect 2094 33454 2146 33506
rect 2146 33454 2148 33506
rect 2092 33452 2148 33454
rect 2252 33506 2308 33508
rect 2252 33454 2254 33506
rect 2254 33454 2306 33506
rect 2306 33454 2308 33506
rect 2252 33452 2308 33454
rect 2412 33506 2468 33508
rect 2412 33454 2414 33506
rect 2414 33454 2466 33506
rect 2466 33454 2468 33506
rect 2412 33452 2468 33454
rect 2572 33506 2628 33508
rect 2572 33454 2574 33506
rect 2574 33454 2626 33506
rect 2626 33454 2628 33506
rect 2572 33452 2628 33454
rect 2732 33506 2788 33508
rect 2732 33454 2734 33506
rect 2734 33454 2786 33506
rect 2786 33454 2788 33506
rect 2732 33452 2788 33454
rect 2892 33506 2948 33508
rect 2892 33454 2894 33506
rect 2894 33454 2946 33506
rect 2946 33454 2948 33506
rect 2892 33452 2948 33454
rect 3052 33506 3108 33508
rect 3052 33454 3054 33506
rect 3054 33454 3106 33506
rect 3106 33454 3108 33506
rect 3052 33452 3108 33454
rect 3212 33506 3268 33508
rect 3212 33454 3214 33506
rect 3214 33454 3266 33506
rect 3266 33454 3268 33506
rect 3212 33452 3268 33454
rect 3372 33506 3428 33508
rect 3372 33454 3374 33506
rect 3374 33454 3426 33506
rect 3426 33454 3428 33506
rect 3372 33452 3428 33454
rect 3532 33506 3588 33508
rect 3532 33454 3534 33506
rect 3534 33454 3586 33506
rect 3586 33454 3588 33506
rect 3532 33452 3588 33454
rect 3692 33506 3748 33508
rect 3692 33454 3694 33506
rect 3694 33454 3746 33506
rect 3746 33454 3748 33506
rect 3692 33452 3748 33454
rect 3852 33506 3908 33508
rect 3852 33454 3854 33506
rect 3854 33454 3906 33506
rect 3906 33454 3908 33506
rect 3852 33452 3908 33454
rect 4012 33506 4068 33508
rect 4012 33454 4014 33506
rect 4014 33454 4066 33506
rect 4066 33454 4068 33506
rect 4012 33452 4068 33454
rect 4172 33506 4228 33508
rect 4172 33454 4174 33506
rect 4174 33454 4226 33506
rect 4226 33454 4228 33506
rect 4172 33452 4228 33454
rect 4332 33506 4388 33508
rect 4332 33454 4334 33506
rect 4334 33454 4386 33506
rect 4386 33454 4388 33506
rect 4332 33452 4388 33454
rect 4492 33506 4548 33508
rect 4492 33454 4494 33506
rect 4494 33454 4546 33506
rect 4546 33454 4548 33506
rect 4492 33452 4548 33454
rect 4652 33506 4708 33508
rect 4652 33454 4654 33506
rect 4654 33454 4706 33506
rect 4706 33454 4708 33506
rect 4652 33452 4708 33454
rect 4812 33506 4868 33508
rect 4812 33454 4814 33506
rect 4814 33454 4866 33506
rect 4866 33454 4868 33506
rect 4812 33452 4868 33454
rect 4972 33506 5028 33508
rect 4972 33454 4974 33506
rect 4974 33454 5026 33506
rect 5026 33454 5028 33506
rect 4972 33452 5028 33454
rect 5132 33506 5188 33508
rect 5132 33454 5134 33506
rect 5134 33454 5186 33506
rect 5186 33454 5188 33506
rect 5132 33452 5188 33454
rect 5292 33506 5348 33508
rect 5292 33454 5294 33506
rect 5294 33454 5346 33506
rect 5346 33454 5348 33506
rect 5292 33452 5348 33454
rect 5452 33506 5508 33508
rect 5452 33454 5454 33506
rect 5454 33454 5506 33506
rect 5506 33454 5508 33506
rect 5452 33452 5508 33454
rect 5612 33506 5668 33508
rect 5612 33454 5614 33506
rect 5614 33454 5666 33506
rect 5666 33454 5668 33506
rect 5612 33452 5668 33454
rect 5772 33506 5828 33508
rect 5772 33454 5774 33506
rect 5774 33454 5826 33506
rect 5826 33454 5828 33506
rect 5772 33452 5828 33454
rect 5932 33506 5988 33508
rect 5932 33454 5934 33506
rect 5934 33454 5986 33506
rect 5986 33454 5988 33506
rect 5932 33452 5988 33454
rect 6092 33506 6148 33508
rect 6092 33454 6094 33506
rect 6094 33454 6146 33506
rect 6146 33454 6148 33506
rect 6092 33452 6148 33454
rect 6252 33506 6308 33508
rect 6252 33454 6254 33506
rect 6254 33454 6306 33506
rect 6306 33454 6308 33506
rect 6252 33452 6308 33454
rect 6412 33506 6468 33508
rect 6412 33454 6414 33506
rect 6414 33454 6466 33506
rect 6466 33454 6468 33506
rect 6412 33452 6468 33454
rect 6572 33506 6628 33508
rect 6572 33454 6574 33506
rect 6574 33454 6626 33506
rect 6626 33454 6628 33506
rect 6572 33452 6628 33454
rect 6732 33506 6788 33508
rect 6732 33454 6734 33506
rect 6734 33454 6786 33506
rect 6786 33454 6788 33506
rect 6732 33452 6788 33454
rect 6892 33506 6948 33508
rect 6892 33454 6894 33506
rect 6894 33454 6946 33506
rect 6946 33454 6948 33506
rect 6892 33452 6948 33454
rect 7052 33506 7108 33508
rect 7052 33454 7054 33506
rect 7054 33454 7106 33506
rect 7106 33454 7108 33506
rect 7052 33452 7108 33454
rect 7212 33506 7268 33508
rect 7212 33454 7214 33506
rect 7214 33454 7266 33506
rect 7266 33454 7268 33506
rect 7212 33452 7268 33454
rect 7372 33506 7428 33508
rect 7372 33454 7374 33506
rect 7374 33454 7426 33506
rect 7426 33454 7428 33506
rect 7372 33452 7428 33454
rect 7532 33506 7588 33508
rect 7532 33454 7534 33506
rect 7534 33454 7586 33506
rect 7586 33454 7588 33506
rect 7532 33452 7588 33454
rect 7692 33506 7748 33508
rect 7692 33454 7694 33506
rect 7694 33454 7746 33506
rect 7746 33454 7748 33506
rect 7692 33452 7748 33454
rect 7852 33506 7908 33508
rect 7852 33454 7854 33506
rect 7854 33454 7906 33506
rect 7906 33454 7908 33506
rect 7852 33452 7908 33454
rect 8012 33506 8068 33508
rect 8012 33454 8014 33506
rect 8014 33454 8066 33506
rect 8066 33454 8068 33506
rect 8012 33452 8068 33454
rect 8172 33506 8228 33508
rect 8172 33454 8174 33506
rect 8174 33454 8226 33506
rect 8226 33454 8228 33506
rect 8172 33452 8228 33454
rect 8332 33506 8388 33508
rect 8332 33454 8334 33506
rect 8334 33454 8386 33506
rect 8386 33454 8388 33506
rect 8332 33452 8388 33454
rect 12012 33452 12068 33508
rect 12332 33452 12388 33508
rect 12492 33506 12548 33508
rect 12492 33454 12494 33506
rect 12494 33454 12546 33506
rect 12546 33454 12548 33506
rect 12492 33452 12548 33454
rect 12652 33506 12708 33508
rect 12652 33454 12654 33506
rect 12654 33454 12706 33506
rect 12706 33454 12708 33506
rect 12652 33452 12708 33454
rect 12812 33506 12868 33508
rect 12812 33454 12814 33506
rect 12814 33454 12866 33506
rect 12866 33454 12868 33506
rect 12812 33452 12868 33454
rect 12972 33506 13028 33508
rect 12972 33454 12974 33506
rect 12974 33454 13026 33506
rect 13026 33454 13028 33506
rect 12972 33452 13028 33454
rect 13132 33506 13188 33508
rect 13132 33454 13134 33506
rect 13134 33454 13186 33506
rect 13186 33454 13188 33506
rect 13132 33452 13188 33454
rect 13292 33506 13348 33508
rect 13292 33454 13294 33506
rect 13294 33454 13346 33506
rect 13346 33454 13348 33506
rect 13292 33452 13348 33454
rect 13452 33506 13508 33508
rect 13452 33454 13454 33506
rect 13454 33454 13506 33506
rect 13506 33454 13508 33506
rect 13452 33452 13508 33454
rect 13612 33506 13668 33508
rect 13612 33454 13614 33506
rect 13614 33454 13666 33506
rect 13666 33454 13668 33506
rect 13612 33452 13668 33454
rect 13772 33506 13828 33508
rect 13772 33454 13774 33506
rect 13774 33454 13826 33506
rect 13826 33454 13828 33506
rect 13772 33452 13828 33454
rect 13932 33506 13988 33508
rect 13932 33454 13934 33506
rect 13934 33454 13986 33506
rect 13986 33454 13988 33506
rect 13932 33452 13988 33454
rect 14092 33506 14148 33508
rect 14092 33454 14094 33506
rect 14094 33454 14146 33506
rect 14146 33454 14148 33506
rect 14092 33452 14148 33454
rect 14252 33506 14308 33508
rect 14252 33454 14254 33506
rect 14254 33454 14306 33506
rect 14306 33454 14308 33506
rect 14252 33452 14308 33454
rect 14412 33506 14468 33508
rect 14412 33454 14414 33506
rect 14414 33454 14466 33506
rect 14466 33454 14468 33506
rect 14412 33452 14468 33454
rect 14572 33506 14628 33508
rect 14572 33454 14574 33506
rect 14574 33454 14626 33506
rect 14626 33454 14628 33506
rect 14572 33452 14628 33454
rect 14732 33506 14788 33508
rect 14732 33454 14734 33506
rect 14734 33454 14786 33506
rect 14786 33454 14788 33506
rect 14732 33452 14788 33454
rect 14892 33506 14948 33508
rect 14892 33454 14894 33506
rect 14894 33454 14946 33506
rect 14946 33454 14948 33506
rect 14892 33452 14948 33454
rect 15052 33506 15108 33508
rect 15052 33454 15054 33506
rect 15054 33454 15106 33506
rect 15106 33454 15108 33506
rect 15052 33452 15108 33454
rect 15212 33506 15268 33508
rect 15212 33454 15214 33506
rect 15214 33454 15266 33506
rect 15266 33454 15268 33506
rect 15212 33452 15268 33454
rect 15372 33506 15428 33508
rect 15372 33454 15374 33506
rect 15374 33454 15426 33506
rect 15426 33454 15428 33506
rect 15372 33452 15428 33454
rect 15532 33506 15588 33508
rect 15532 33454 15534 33506
rect 15534 33454 15586 33506
rect 15586 33454 15588 33506
rect 15532 33452 15588 33454
rect 15692 33506 15748 33508
rect 15692 33454 15694 33506
rect 15694 33454 15746 33506
rect 15746 33454 15748 33506
rect 15692 33452 15748 33454
rect 15852 33506 15908 33508
rect 15852 33454 15854 33506
rect 15854 33454 15906 33506
rect 15906 33454 15908 33506
rect 15852 33452 15908 33454
rect 16012 33506 16068 33508
rect 16012 33454 16014 33506
rect 16014 33454 16066 33506
rect 16066 33454 16068 33506
rect 16012 33452 16068 33454
rect 16172 33506 16228 33508
rect 16172 33454 16174 33506
rect 16174 33454 16226 33506
rect 16226 33454 16228 33506
rect 16172 33452 16228 33454
rect 16332 33506 16388 33508
rect 16332 33454 16334 33506
rect 16334 33454 16386 33506
rect 16386 33454 16388 33506
rect 16332 33452 16388 33454
rect 16492 33506 16548 33508
rect 16492 33454 16494 33506
rect 16494 33454 16546 33506
rect 16546 33454 16548 33506
rect 16492 33452 16548 33454
rect 16652 33506 16708 33508
rect 16652 33454 16654 33506
rect 16654 33454 16706 33506
rect 16706 33454 16708 33506
rect 16652 33452 16708 33454
rect 16812 33506 16868 33508
rect 16812 33454 16814 33506
rect 16814 33454 16866 33506
rect 16866 33454 16868 33506
rect 16812 33452 16868 33454
rect 16972 33506 17028 33508
rect 16972 33454 16974 33506
rect 16974 33454 17026 33506
rect 17026 33454 17028 33506
rect 16972 33452 17028 33454
rect 17132 33506 17188 33508
rect 17132 33454 17134 33506
rect 17134 33454 17186 33506
rect 17186 33454 17188 33506
rect 17132 33452 17188 33454
rect 17292 33506 17348 33508
rect 17292 33454 17294 33506
rect 17294 33454 17346 33506
rect 17346 33454 17348 33506
rect 17292 33452 17348 33454
rect 17452 33506 17508 33508
rect 17452 33454 17454 33506
rect 17454 33454 17506 33506
rect 17506 33454 17508 33506
rect 17452 33452 17508 33454
rect 17612 33506 17668 33508
rect 17612 33454 17614 33506
rect 17614 33454 17666 33506
rect 17666 33454 17668 33506
rect 17612 33452 17668 33454
rect 17772 33506 17828 33508
rect 17772 33454 17774 33506
rect 17774 33454 17826 33506
rect 17826 33454 17828 33506
rect 17772 33452 17828 33454
rect 17932 33506 17988 33508
rect 17932 33454 17934 33506
rect 17934 33454 17986 33506
rect 17986 33454 17988 33506
rect 17932 33452 17988 33454
rect 18092 33506 18148 33508
rect 18092 33454 18094 33506
rect 18094 33454 18146 33506
rect 18146 33454 18148 33506
rect 18092 33452 18148 33454
rect 18252 33506 18308 33508
rect 18252 33454 18254 33506
rect 18254 33454 18306 33506
rect 18306 33454 18308 33506
rect 18252 33452 18308 33454
rect 18412 33506 18468 33508
rect 18412 33454 18414 33506
rect 18414 33454 18466 33506
rect 18466 33454 18468 33506
rect 18412 33452 18468 33454
rect 18572 33506 18628 33508
rect 18572 33454 18574 33506
rect 18574 33454 18626 33506
rect 18626 33454 18628 33506
rect 18572 33452 18628 33454
rect 18732 33506 18788 33508
rect 18732 33454 18734 33506
rect 18734 33454 18786 33506
rect 18786 33454 18788 33506
rect 18732 33452 18788 33454
rect 18892 33506 18948 33508
rect 18892 33454 18894 33506
rect 18894 33454 18946 33506
rect 18946 33454 18948 33506
rect 18892 33452 18948 33454
rect 19052 33452 19108 33508
rect 19372 33452 19428 33508
rect 23132 33506 23188 33508
rect 23132 33454 23134 33506
rect 23134 33454 23186 33506
rect 23186 33454 23188 33506
rect 23132 33452 23188 33454
rect 23292 33506 23348 33508
rect 23292 33454 23294 33506
rect 23294 33454 23346 33506
rect 23346 33454 23348 33506
rect 23292 33452 23348 33454
rect 23452 33506 23508 33508
rect 23452 33454 23454 33506
rect 23454 33454 23506 33506
rect 23506 33454 23508 33506
rect 23452 33452 23508 33454
rect 23612 33506 23668 33508
rect 23612 33454 23614 33506
rect 23614 33454 23666 33506
rect 23666 33454 23668 33506
rect 23612 33452 23668 33454
rect 23772 33506 23828 33508
rect 23772 33454 23774 33506
rect 23774 33454 23826 33506
rect 23826 33454 23828 33506
rect 23772 33452 23828 33454
rect 23932 33506 23988 33508
rect 23932 33454 23934 33506
rect 23934 33454 23986 33506
rect 23986 33454 23988 33506
rect 23932 33452 23988 33454
rect 24092 33506 24148 33508
rect 24092 33454 24094 33506
rect 24094 33454 24146 33506
rect 24146 33454 24148 33506
rect 24092 33452 24148 33454
rect 24252 33506 24308 33508
rect 24252 33454 24254 33506
rect 24254 33454 24306 33506
rect 24306 33454 24308 33506
rect 24252 33452 24308 33454
rect 24412 33506 24468 33508
rect 24412 33454 24414 33506
rect 24414 33454 24466 33506
rect 24466 33454 24468 33506
rect 24412 33452 24468 33454
rect 24572 33506 24628 33508
rect 24572 33454 24574 33506
rect 24574 33454 24626 33506
rect 24626 33454 24628 33506
rect 24572 33452 24628 33454
rect 24732 33506 24788 33508
rect 24732 33454 24734 33506
rect 24734 33454 24786 33506
rect 24786 33454 24788 33506
rect 24732 33452 24788 33454
rect 24892 33506 24948 33508
rect 24892 33454 24894 33506
rect 24894 33454 24946 33506
rect 24946 33454 24948 33506
rect 24892 33452 24948 33454
rect 25052 33506 25108 33508
rect 25052 33454 25054 33506
rect 25054 33454 25106 33506
rect 25106 33454 25108 33506
rect 25052 33452 25108 33454
rect 25212 33506 25268 33508
rect 25212 33454 25214 33506
rect 25214 33454 25266 33506
rect 25266 33454 25268 33506
rect 25212 33452 25268 33454
rect 25372 33506 25428 33508
rect 25372 33454 25374 33506
rect 25374 33454 25426 33506
rect 25426 33454 25428 33506
rect 25372 33452 25428 33454
rect 25532 33506 25588 33508
rect 25532 33454 25534 33506
rect 25534 33454 25586 33506
rect 25586 33454 25588 33506
rect 25532 33452 25588 33454
rect 25692 33506 25748 33508
rect 25692 33454 25694 33506
rect 25694 33454 25746 33506
rect 25746 33454 25748 33506
rect 25692 33452 25748 33454
rect 25852 33506 25908 33508
rect 25852 33454 25854 33506
rect 25854 33454 25906 33506
rect 25906 33454 25908 33506
rect 25852 33452 25908 33454
rect 26012 33506 26068 33508
rect 26012 33454 26014 33506
rect 26014 33454 26066 33506
rect 26066 33454 26068 33506
rect 26012 33452 26068 33454
rect 26172 33506 26228 33508
rect 26172 33454 26174 33506
rect 26174 33454 26226 33506
rect 26226 33454 26228 33506
rect 26172 33452 26228 33454
rect 26332 33506 26388 33508
rect 26332 33454 26334 33506
rect 26334 33454 26386 33506
rect 26386 33454 26388 33506
rect 26332 33452 26388 33454
rect 26492 33506 26548 33508
rect 26492 33454 26494 33506
rect 26494 33454 26546 33506
rect 26546 33454 26548 33506
rect 26492 33452 26548 33454
rect 26652 33506 26708 33508
rect 26652 33454 26654 33506
rect 26654 33454 26706 33506
rect 26706 33454 26708 33506
rect 26652 33452 26708 33454
rect 26812 33506 26868 33508
rect 26812 33454 26814 33506
rect 26814 33454 26866 33506
rect 26866 33454 26868 33506
rect 26812 33452 26868 33454
rect 26972 33506 27028 33508
rect 26972 33454 26974 33506
rect 26974 33454 27026 33506
rect 27026 33454 27028 33506
rect 26972 33452 27028 33454
rect 27132 33506 27188 33508
rect 27132 33454 27134 33506
rect 27134 33454 27186 33506
rect 27186 33454 27188 33506
rect 27132 33452 27188 33454
rect 27292 33506 27348 33508
rect 27292 33454 27294 33506
rect 27294 33454 27346 33506
rect 27346 33454 27348 33506
rect 27292 33452 27348 33454
rect 27452 33506 27508 33508
rect 27452 33454 27454 33506
rect 27454 33454 27506 33506
rect 27506 33454 27508 33506
rect 27452 33452 27508 33454
rect 27612 33506 27668 33508
rect 27612 33454 27614 33506
rect 27614 33454 27666 33506
rect 27666 33454 27668 33506
rect 27612 33452 27668 33454
rect 27772 33506 27828 33508
rect 27772 33454 27774 33506
rect 27774 33454 27826 33506
rect 27826 33454 27828 33506
rect 27772 33452 27828 33454
rect 27932 33506 27988 33508
rect 27932 33454 27934 33506
rect 27934 33454 27986 33506
rect 27986 33454 27988 33506
rect 27932 33452 27988 33454
rect 28092 33506 28148 33508
rect 28092 33454 28094 33506
rect 28094 33454 28146 33506
rect 28146 33454 28148 33506
rect 28092 33452 28148 33454
rect 28252 33506 28308 33508
rect 28252 33454 28254 33506
rect 28254 33454 28306 33506
rect 28306 33454 28308 33506
rect 28252 33452 28308 33454
rect 28412 33506 28468 33508
rect 28412 33454 28414 33506
rect 28414 33454 28466 33506
rect 28466 33454 28468 33506
rect 28412 33452 28468 33454
rect 28572 33506 28628 33508
rect 28572 33454 28574 33506
rect 28574 33454 28626 33506
rect 28626 33454 28628 33506
rect 28572 33452 28628 33454
rect 28732 33506 28788 33508
rect 28732 33454 28734 33506
rect 28734 33454 28786 33506
rect 28786 33454 28788 33506
rect 28732 33452 28788 33454
rect 28892 33506 28948 33508
rect 28892 33454 28894 33506
rect 28894 33454 28946 33506
rect 28946 33454 28948 33506
rect 28892 33452 28948 33454
rect 29052 33506 29108 33508
rect 29052 33454 29054 33506
rect 29054 33454 29106 33506
rect 29106 33454 29108 33506
rect 29052 33452 29108 33454
rect 29212 33506 29268 33508
rect 29212 33454 29214 33506
rect 29214 33454 29266 33506
rect 29266 33454 29268 33506
rect 29212 33452 29268 33454
rect 29372 33506 29428 33508
rect 29372 33454 29374 33506
rect 29374 33454 29426 33506
rect 29426 33454 29428 33506
rect 29372 33452 29428 33454
rect 29532 33452 29588 33508
rect 29852 33452 29908 33508
rect 33532 33506 33588 33508
rect 33532 33454 33534 33506
rect 33534 33454 33586 33506
rect 33586 33454 33588 33506
rect 33532 33452 33588 33454
rect 33692 33506 33748 33508
rect 33692 33454 33694 33506
rect 33694 33454 33746 33506
rect 33746 33454 33748 33506
rect 33692 33452 33748 33454
rect 33852 33506 33908 33508
rect 33852 33454 33854 33506
rect 33854 33454 33906 33506
rect 33906 33454 33908 33506
rect 33852 33452 33908 33454
rect 34012 33506 34068 33508
rect 34012 33454 34014 33506
rect 34014 33454 34066 33506
rect 34066 33454 34068 33506
rect 34012 33452 34068 33454
rect 34172 33506 34228 33508
rect 34172 33454 34174 33506
rect 34174 33454 34226 33506
rect 34226 33454 34228 33506
rect 34172 33452 34228 33454
rect 34332 33506 34388 33508
rect 34332 33454 34334 33506
rect 34334 33454 34386 33506
rect 34386 33454 34388 33506
rect 34332 33452 34388 33454
rect 34492 33506 34548 33508
rect 34492 33454 34494 33506
rect 34494 33454 34546 33506
rect 34546 33454 34548 33506
rect 34492 33452 34548 33454
rect 34652 33506 34708 33508
rect 34652 33454 34654 33506
rect 34654 33454 34706 33506
rect 34706 33454 34708 33506
rect 34652 33452 34708 33454
rect 34812 33506 34868 33508
rect 34812 33454 34814 33506
rect 34814 33454 34866 33506
rect 34866 33454 34868 33506
rect 34812 33452 34868 33454
rect 34972 33506 35028 33508
rect 34972 33454 34974 33506
rect 34974 33454 35026 33506
rect 35026 33454 35028 33506
rect 34972 33452 35028 33454
rect 35132 33506 35188 33508
rect 35132 33454 35134 33506
rect 35134 33454 35186 33506
rect 35186 33454 35188 33506
rect 35132 33452 35188 33454
rect 35292 33506 35348 33508
rect 35292 33454 35294 33506
rect 35294 33454 35346 33506
rect 35346 33454 35348 33506
rect 35292 33452 35348 33454
rect 35452 33506 35508 33508
rect 35452 33454 35454 33506
rect 35454 33454 35506 33506
rect 35506 33454 35508 33506
rect 35452 33452 35508 33454
rect 35612 33506 35668 33508
rect 35612 33454 35614 33506
rect 35614 33454 35666 33506
rect 35666 33454 35668 33506
rect 35612 33452 35668 33454
rect 35772 33506 35828 33508
rect 35772 33454 35774 33506
rect 35774 33454 35826 33506
rect 35826 33454 35828 33506
rect 35772 33452 35828 33454
rect 35932 33506 35988 33508
rect 35932 33454 35934 33506
rect 35934 33454 35986 33506
rect 35986 33454 35988 33506
rect 35932 33452 35988 33454
rect 36092 33506 36148 33508
rect 36092 33454 36094 33506
rect 36094 33454 36146 33506
rect 36146 33454 36148 33506
rect 36092 33452 36148 33454
rect 36252 33506 36308 33508
rect 36252 33454 36254 33506
rect 36254 33454 36306 33506
rect 36306 33454 36308 33506
rect 36252 33452 36308 33454
rect 36412 33506 36468 33508
rect 36412 33454 36414 33506
rect 36414 33454 36466 33506
rect 36466 33454 36468 33506
rect 36412 33452 36468 33454
rect 36572 33506 36628 33508
rect 36572 33454 36574 33506
rect 36574 33454 36626 33506
rect 36626 33454 36628 33506
rect 36572 33452 36628 33454
rect 36732 33506 36788 33508
rect 36732 33454 36734 33506
rect 36734 33454 36786 33506
rect 36786 33454 36788 33506
rect 36732 33452 36788 33454
rect 36892 33506 36948 33508
rect 36892 33454 36894 33506
rect 36894 33454 36946 33506
rect 36946 33454 36948 33506
rect 36892 33452 36948 33454
rect 37052 33506 37108 33508
rect 37052 33454 37054 33506
rect 37054 33454 37106 33506
rect 37106 33454 37108 33506
rect 37052 33452 37108 33454
rect 37212 33506 37268 33508
rect 37212 33454 37214 33506
rect 37214 33454 37266 33506
rect 37266 33454 37268 33506
rect 37212 33452 37268 33454
rect 37372 33506 37428 33508
rect 37372 33454 37374 33506
rect 37374 33454 37426 33506
rect 37426 33454 37428 33506
rect 37372 33452 37428 33454
rect 37532 33506 37588 33508
rect 37532 33454 37534 33506
rect 37534 33454 37586 33506
rect 37586 33454 37588 33506
rect 37532 33452 37588 33454
rect 37692 33506 37748 33508
rect 37692 33454 37694 33506
rect 37694 33454 37746 33506
rect 37746 33454 37748 33506
rect 37692 33452 37748 33454
rect 37852 33506 37908 33508
rect 37852 33454 37854 33506
rect 37854 33454 37906 33506
rect 37906 33454 37908 33506
rect 37852 33452 37908 33454
rect 38012 33506 38068 33508
rect 38012 33454 38014 33506
rect 38014 33454 38066 33506
rect 38066 33454 38068 33506
rect 38012 33452 38068 33454
rect 38172 33506 38228 33508
rect 38172 33454 38174 33506
rect 38174 33454 38226 33506
rect 38226 33454 38228 33506
rect 38172 33452 38228 33454
rect 38332 33506 38388 33508
rect 38332 33454 38334 33506
rect 38334 33454 38386 33506
rect 38386 33454 38388 33506
rect 38332 33452 38388 33454
rect 38492 33506 38548 33508
rect 38492 33454 38494 33506
rect 38494 33454 38546 33506
rect 38546 33454 38548 33506
rect 38492 33452 38548 33454
rect 38652 33506 38708 33508
rect 38652 33454 38654 33506
rect 38654 33454 38706 33506
rect 38706 33454 38708 33506
rect 38652 33452 38708 33454
rect 38812 33506 38868 33508
rect 38812 33454 38814 33506
rect 38814 33454 38866 33506
rect 38866 33454 38868 33506
rect 38812 33452 38868 33454
rect 38972 33506 39028 33508
rect 38972 33454 38974 33506
rect 38974 33454 39026 33506
rect 39026 33454 39028 33506
rect 38972 33452 39028 33454
rect 39132 33506 39188 33508
rect 39132 33454 39134 33506
rect 39134 33454 39186 33506
rect 39186 33454 39188 33506
rect 39132 33452 39188 33454
rect 39292 33506 39348 33508
rect 39292 33454 39294 33506
rect 39294 33454 39346 33506
rect 39346 33454 39348 33506
rect 39292 33452 39348 33454
rect 39452 33506 39508 33508
rect 39452 33454 39454 33506
rect 39454 33454 39506 33506
rect 39506 33454 39508 33506
rect 39452 33452 39508 33454
rect 39612 33506 39668 33508
rect 39612 33454 39614 33506
rect 39614 33454 39666 33506
rect 39666 33454 39668 33506
rect 39612 33452 39668 33454
rect 39772 33506 39828 33508
rect 39772 33454 39774 33506
rect 39774 33454 39826 33506
rect 39826 33454 39828 33506
rect 39772 33452 39828 33454
rect 39932 33506 39988 33508
rect 39932 33454 39934 33506
rect 39934 33454 39986 33506
rect 39986 33454 39988 33506
rect 39932 33452 39988 33454
rect 40092 33506 40148 33508
rect 40092 33454 40094 33506
rect 40094 33454 40146 33506
rect 40146 33454 40148 33506
rect 40092 33452 40148 33454
rect 40252 33506 40308 33508
rect 40252 33454 40254 33506
rect 40254 33454 40306 33506
rect 40306 33454 40308 33506
rect 40252 33452 40308 33454
rect 40412 33506 40468 33508
rect 40412 33454 40414 33506
rect 40414 33454 40466 33506
rect 40466 33454 40468 33506
rect 40412 33452 40468 33454
rect 40572 33506 40628 33508
rect 40572 33454 40574 33506
rect 40574 33454 40626 33506
rect 40626 33454 40628 33506
rect 40572 33452 40628 33454
rect 40732 33506 40788 33508
rect 40732 33454 40734 33506
rect 40734 33454 40786 33506
rect 40786 33454 40788 33506
rect 40732 33452 40788 33454
rect 40892 33506 40948 33508
rect 40892 33454 40894 33506
rect 40894 33454 40946 33506
rect 40946 33454 40948 33506
rect 40892 33452 40948 33454
rect 41052 33506 41108 33508
rect 41052 33454 41054 33506
rect 41054 33454 41106 33506
rect 41106 33454 41108 33506
rect 41052 33452 41108 33454
rect 41212 33506 41268 33508
rect 41212 33454 41214 33506
rect 41214 33454 41266 33506
rect 41266 33454 41268 33506
rect 41212 33452 41268 33454
rect 41372 33506 41428 33508
rect 41372 33454 41374 33506
rect 41374 33454 41426 33506
rect 41426 33454 41428 33506
rect 41372 33452 41428 33454
rect 41532 33506 41588 33508
rect 41532 33454 41534 33506
rect 41534 33454 41586 33506
rect 41586 33454 41588 33506
rect 41532 33452 41588 33454
rect 41692 33506 41748 33508
rect 41692 33454 41694 33506
rect 41694 33454 41746 33506
rect 41746 33454 41748 33506
rect 41692 33452 41748 33454
rect 41852 33506 41908 33508
rect 41852 33454 41854 33506
rect 41854 33454 41906 33506
rect 41906 33454 41908 33506
rect 41852 33452 41908 33454
rect 12 33346 68 33348
rect 12 33294 14 33346
rect 14 33294 66 33346
rect 66 33294 68 33346
rect 12 33292 68 33294
rect 172 33346 228 33348
rect 172 33294 174 33346
rect 174 33294 226 33346
rect 226 33294 228 33346
rect 172 33292 228 33294
rect 332 33346 388 33348
rect 332 33294 334 33346
rect 334 33294 386 33346
rect 386 33294 388 33346
rect 332 33292 388 33294
rect 492 33346 548 33348
rect 492 33294 494 33346
rect 494 33294 546 33346
rect 546 33294 548 33346
rect 492 33292 548 33294
rect 652 33346 708 33348
rect 652 33294 654 33346
rect 654 33294 706 33346
rect 706 33294 708 33346
rect 652 33292 708 33294
rect 812 33346 868 33348
rect 812 33294 814 33346
rect 814 33294 866 33346
rect 866 33294 868 33346
rect 812 33292 868 33294
rect 972 33346 1028 33348
rect 972 33294 974 33346
rect 974 33294 1026 33346
rect 1026 33294 1028 33346
rect 972 33292 1028 33294
rect 1132 33346 1188 33348
rect 1132 33294 1134 33346
rect 1134 33294 1186 33346
rect 1186 33294 1188 33346
rect 1132 33292 1188 33294
rect 1292 33346 1348 33348
rect 1292 33294 1294 33346
rect 1294 33294 1346 33346
rect 1346 33294 1348 33346
rect 1292 33292 1348 33294
rect 1452 33346 1508 33348
rect 1452 33294 1454 33346
rect 1454 33294 1506 33346
rect 1506 33294 1508 33346
rect 1452 33292 1508 33294
rect 1612 33346 1668 33348
rect 1612 33294 1614 33346
rect 1614 33294 1666 33346
rect 1666 33294 1668 33346
rect 1612 33292 1668 33294
rect 1772 33346 1828 33348
rect 1772 33294 1774 33346
rect 1774 33294 1826 33346
rect 1826 33294 1828 33346
rect 1772 33292 1828 33294
rect 1932 33346 1988 33348
rect 1932 33294 1934 33346
rect 1934 33294 1986 33346
rect 1986 33294 1988 33346
rect 1932 33292 1988 33294
rect 2092 33346 2148 33348
rect 2092 33294 2094 33346
rect 2094 33294 2146 33346
rect 2146 33294 2148 33346
rect 2092 33292 2148 33294
rect 2252 33346 2308 33348
rect 2252 33294 2254 33346
rect 2254 33294 2306 33346
rect 2306 33294 2308 33346
rect 2252 33292 2308 33294
rect 2412 33346 2468 33348
rect 2412 33294 2414 33346
rect 2414 33294 2466 33346
rect 2466 33294 2468 33346
rect 2412 33292 2468 33294
rect 2572 33346 2628 33348
rect 2572 33294 2574 33346
rect 2574 33294 2626 33346
rect 2626 33294 2628 33346
rect 2572 33292 2628 33294
rect 2732 33346 2788 33348
rect 2732 33294 2734 33346
rect 2734 33294 2786 33346
rect 2786 33294 2788 33346
rect 2732 33292 2788 33294
rect 2892 33346 2948 33348
rect 2892 33294 2894 33346
rect 2894 33294 2946 33346
rect 2946 33294 2948 33346
rect 2892 33292 2948 33294
rect 3052 33346 3108 33348
rect 3052 33294 3054 33346
rect 3054 33294 3106 33346
rect 3106 33294 3108 33346
rect 3052 33292 3108 33294
rect 3212 33346 3268 33348
rect 3212 33294 3214 33346
rect 3214 33294 3266 33346
rect 3266 33294 3268 33346
rect 3212 33292 3268 33294
rect 3372 33346 3428 33348
rect 3372 33294 3374 33346
rect 3374 33294 3426 33346
rect 3426 33294 3428 33346
rect 3372 33292 3428 33294
rect 3532 33346 3588 33348
rect 3532 33294 3534 33346
rect 3534 33294 3586 33346
rect 3586 33294 3588 33346
rect 3532 33292 3588 33294
rect 3692 33346 3748 33348
rect 3692 33294 3694 33346
rect 3694 33294 3746 33346
rect 3746 33294 3748 33346
rect 3692 33292 3748 33294
rect 3852 33346 3908 33348
rect 3852 33294 3854 33346
rect 3854 33294 3906 33346
rect 3906 33294 3908 33346
rect 3852 33292 3908 33294
rect 4012 33346 4068 33348
rect 4012 33294 4014 33346
rect 4014 33294 4066 33346
rect 4066 33294 4068 33346
rect 4012 33292 4068 33294
rect 4172 33346 4228 33348
rect 4172 33294 4174 33346
rect 4174 33294 4226 33346
rect 4226 33294 4228 33346
rect 4172 33292 4228 33294
rect 4332 33346 4388 33348
rect 4332 33294 4334 33346
rect 4334 33294 4386 33346
rect 4386 33294 4388 33346
rect 4332 33292 4388 33294
rect 4492 33346 4548 33348
rect 4492 33294 4494 33346
rect 4494 33294 4546 33346
rect 4546 33294 4548 33346
rect 4492 33292 4548 33294
rect 4652 33346 4708 33348
rect 4652 33294 4654 33346
rect 4654 33294 4706 33346
rect 4706 33294 4708 33346
rect 4652 33292 4708 33294
rect 4812 33346 4868 33348
rect 4812 33294 4814 33346
rect 4814 33294 4866 33346
rect 4866 33294 4868 33346
rect 4812 33292 4868 33294
rect 4972 33346 5028 33348
rect 4972 33294 4974 33346
rect 4974 33294 5026 33346
rect 5026 33294 5028 33346
rect 4972 33292 5028 33294
rect 5132 33346 5188 33348
rect 5132 33294 5134 33346
rect 5134 33294 5186 33346
rect 5186 33294 5188 33346
rect 5132 33292 5188 33294
rect 5292 33346 5348 33348
rect 5292 33294 5294 33346
rect 5294 33294 5346 33346
rect 5346 33294 5348 33346
rect 5292 33292 5348 33294
rect 5452 33346 5508 33348
rect 5452 33294 5454 33346
rect 5454 33294 5506 33346
rect 5506 33294 5508 33346
rect 5452 33292 5508 33294
rect 5612 33346 5668 33348
rect 5612 33294 5614 33346
rect 5614 33294 5666 33346
rect 5666 33294 5668 33346
rect 5612 33292 5668 33294
rect 5772 33346 5828 33348
rect 5772 33294 5774 33346
rect 5774 33294 5826 33346
rect 5826 33294 5828 33346
rect 5772 33292 5828 33294
rect 5932 33346 5988 33348
rect 5932 33294 5934 33346
rect 5934 33294 5986 33346
rect 5986 33294 5988 33346
rect 5932 33292 5988 33294
rect 6092 33346 6148 33348
rect 6092 33294 6094 33346
rect 6094 33294 6146 33346
rect 6146 33294 6148 33346
rect 6092 33292 6148 33294
rect 6252 33346 6308 33348
rect 6252 33294 6254 33346
rect 6254 33294 6306 33346
rect 6306 33294 6308 33346
rect 6252 33292 6308 33294
rect 6412 33346 6468 33348
rect 6412 33294 6414 33346
rect 6414 33294 6466 33346
rect 6466 33294 6468 33346
rect 6412 33292 6468 33294
rect 6572 33346 6628 33348
rect 6572 33294 6574 33346
rect 6574 33294 6626 33346
rect 6626 33294 6628 33346
rect 6572 33292 6628 33294
rect 6732 33346 6788 33348
rect 6732 33294 6734 33346
rect 6734 33294 6786 33346
rect 6786 33294 6788 33346
rect 6732 33292 6788 33294
rect 6892 33346 6948 33348
rect 6892 33294 6894 33346
rect 6894 33294 6946 33346
rect 6946 33294 6948 33346
rect 6892 33292 6948 33294
rect 7052 33346 7108 33348
rect 7052 33294 7054 33346
rect 7054 33294 7106 33346
rect 7106 33294 7108 33346
rect 7052 33292 7108 33294
rect 7212 33346 7268 33348
rect 7212 33294 7214 33346
rect 7214 33294 7266 33346
rect 7266 33294 7268 33346
rect 7212 33292 7268 33294
rect 7372 33346 7428 33348
rect 7372 33294 7374 33346
rect 7374 33294 7426 33346
rect 7426 33294 7428 33346
rect 7372 33292 7428 33294
rect 7532 33346 7588 33348
rect 7532 33294 7534 33346
rect 7534 33294 7586 33346
rect 7586 33294 7588 33346
rect 7532 33292 7588 33294
rect 7692 33346 7748 33348
rect 7692 33294 7694 33346
rect 7694 33294 7746 33346
rect 7746 33294 7748 33346
rect 7692 33292 7748 33294
rect 7852 33346 7908 33348
rect 7852 33294 7854 33346
rect 7854 33294 7906 33346
rect 7906 33294 7908 33346
rect 7852 33292 7908 33294
rect 8012 33346 8068 33348
rect 8012 33294 8014 33346
rect 8014 33294 8066 33346
rect 8066 33294 8068 33346
rect 8012 33292 8068 33294
rect 8172 33346 8228 33348
rect 8172 33294 8174 33346
rect 8174 33294 8226 33346
rect 8226 33294 8228 33346
rect 8172 33292 8228 33294
rect 8332 33346 8388 33348
rect 8332 33294 8334 33346
rect 8334 33294 8386 33346
rect 8386 33294 8388 33346
rect 8332 33292 8388 33294
rect 8492 33292 8548 33348
rect 8812 33292 8868 33348
rect 12492 33346 12548 33348
rect 12492 33294 12494 33346
rect 12494 33294 12546 33346
rect 12546 33294 12548 33346
rect 12492 33292 12548 33294
rect 12652 33346 12708 33348
rect 12652 33294 12654 33346
rect 12654 33294 12706 33346
rect 12706 33294 12708 33346
rect 12652 33292 12708 33294
rect 12812 33346 12868 33348
rect 12812 33294 12814 33346
rect 12814 33294 12866 33346
rect 12866 33294 12868 33346
rect 12812 33292 12868 33294
rect 12972 33346 13028 33348
rect 12972 33294 12974 33346
rect 12974 33294 13026 33346
rect 13026 33294 13028 33346
rect 12972 33292 13028 33294
rect 13132 33346 13188 33348
rect 13132 33294 13134 33346
rect 13134 33294 13186 33346
rect 13186 33294 13188 33346
rect 13132 33292 13188 33294
rect 13292 33346 13348 33348
rect 13292 33294 13294 33346
rect 13294 33294 13346 33346
rect 13346 33294 13348 33346
rect 13292 33292 13348 33294
rect 13452 33346 13508 33348
rect 13452 33294 13454 33346
rect 13454 33294 13506 33346
rect 13506 33294 13508 33346
rect 13452 33292 13508 33294
rect 13612 33346 13668 33348
rect 13612 33294 13614 33346
rect 13614 33294 13666 33346
rect 13666 33294 13668 33346
rect 13612 33292 13668 33294
rect 13772 33346 13828 33348
rect 13772 33294 13774 33346
rect 13774 33294 13826 33346
rect 13826 33294 13828 33346
rect 13772 33292 13828 33294
rect 13932 33346 13988 33348
rect 13932 33294 13934 33346
rect 13934 33294 13986 33346
rect 13986 33294 13988 33346
rect 13932 33292 13988 33294
rect 14092 33346 14148 33348
rect 14092 33294 14094 33346
rect 14094 33294 14146 33346
rect 14146 33294 14148 33346
rect 14092 33292 14148 33294
rect 14252 33346 14308 33348
rect 14252 33294 14254 33346
rect 14254 33294 14306 33346
rect 14306 33294 14308 33346
rect 14252 33292 14308 33294
rect 14412 33346 14468 33348
rect 14412 33294 14414 33346
rect 14414 33294 14466 33346
rect 14466 33294 14468 33346
rect 14412 33292 14468 33294
rect 14572 33346 14628 33348
rect 14572 33294 14574 33346
rect 14574 33294 14626 33346
rect 14626 33294 14628 33346
rect 14572 33292 14628 33294
rect 14732 33346 14788 33348
rect 14732 33294 14734 33346
rect 14734 33294 14786 33346
rect 14786 33294 14788 33346
rect 14732 33292 14788 33294
rect 14892 33346 14948 33348
rect 14892 33294 14894 33346
rect 14894 33294 14946 33346
rect 14946 33294 14948 33346
rect 14892 33292 14948 33294
rect 15052 33346 15108 33348
rect 15052 33294 15054 33346
rect 15054 33294 15106 33346
rect 15106 33294 15108 33346
rect 15052 33292 15108 33294
rect 15212 33346 15268 33348
rect 15212 33294 15214 33346
rect 15214 33294 15266 33346
rect 15266 33294 15268 33346
rect 15212 33292 15268 33294
rect 15372 33346 15428 33348
rect 15372 33294 15374 33346
rect 15374 33294 15426 33346
rect 15426 33294 15428 33346
rect 15372 33292 15428 33294
rect 15532 33346 15588 33348
rect 15532 33294 15534 33346
rect 15534 33294 15586 33346
rect 15586 33294 15588 33346
rect 15532 33292 15588 33294
rect 15692 33346 15748 33348
rect 15692 33294 15694 33346
rect 15694 33294 15746 33346
rect 15746 33294 15748 33346
rect 15692 33292 15748 33294
rect 15852 33346 15908 33348
rect 15852 33294 15854 33346
rect 15854 33294 15906 33346
rect 15906 33294 15908 33346
rect 15852 33292 15908 33294
rect 16012 33346 16068 33348
rect 16012 33294 16014 33346
rect 16014 33294 16066 33346
rect 16066 33294 16068 33346
rect 16012 33292 16068 33294
rect 16172 33346 16228 33348
rect 16172 33294 16174 33346
rect 16174 33294 16226 33346
rect 16226 33294 16228 33346
rect 16172 33292 16228 33294
rect 16332 33346 16388 33348
rect 16332 33294 16334 33346
rect 16334 33294 16386 33346
rect 16386 33294 16388 33346
rect 16332 33292 16388 33294
rect 16492 33346 16548 33348
rect 16492 33294 16494 33346
rect 16494 33294 16546 33346
rect 16546 33294 16548 33346
rect 16492 33292 16548 33294
rect 16652 33346 16708 33348
rect 16652 33294 16654 33346
rect 16654 33294 16706 33346
rect 16706 33294 16708 33346
rect 16652 33292 16708 33294
rect 16812 33346 16868 33348
rect 16812 33294 16814 33346
rect 16814 33294 16866 33346
rect 16866 33294 16868 33346
rect 16812 33292 16868 33294
rect 16972 33346 17028 33348
rect 16972 33294 16974 33346
rect 16974 33294 17026 33346
rect 17026 33294 17028 33346
rect 16972 33292 17028 33294
rect 17132 33346 17188 33348
rect 17132 33294 17134 33346
rect 17134 33294 17186 33346
rect 17186 33294 17188 33346
rect 17132 33292 17188 33294
rect 17292 33346 17348 33348
rect 17292 33294 17294 33346
rect 17294 33294 17346 33346
rect 17346 33294 17348 33346
rect 17292 33292 17348 33294
rect 17452 33346 17508 33348
rect 17452 33294 17454 33346
rect 17454 33294 17506 33346
rect 17506 33294 17508 33346
rect 17452 33292 17508 33294
rect 17612 33346 17668 33348
rect 17612 33294 17614 33346
rect 17614 33294 17666 33346
rect 17666 33294 17668 33346
rect 17612 33292 17668 33294
rect 17772 33346 17828 33348
rect 17772 33294 17774 33346
rect 17774 33294 17826 33346
rect 17826 33294 17828 33346
rect 17772 33292 17828 33294
rect 17932 33346 17988 33348
rect 17932 33294 17934 33346
rect 17934 33294 17986 33346
rect 17986 33294 17988 33346
rect 17932 33292 17988 33294
rect 18092 33346 18148 33348
rect 18092 33294 18094 33346
rect 18094 33294 18146 33346
rect 18146 33294 18148 33346
rect 18092 33292 18148 33294
rect 18252 33346 18308 33348
rect 18252 33294 18254 33346
rect 18254 33294 18306 33346
rect 18306 33294 18308 33346
rect 18252 33292 18308 33294
rect 18412 33346 18468 33348
rect 18412 33294 18414 33346
rect 18414 33294 18466 33346
rect 18466 33294 18468 33346
rect 18412 33292 18468 33294
rect 18572 33346 18628 33348
rect 18572 33294 18574 33346
rect 18574 33294 18626 33346
rect 18626 33294 18628 33346
rect 18572 33292 18628 33294
rect 18732 33346 18788 33348
rect 18732 33294 18734 33346
rect 18734 33294 18786 33346
rect 18786 33294 18788 33346
rect 18732 33292 18788 33294
rect 18892 33346 18948 33348
rect 18892 33294 18894 33346
rect 18894 33294 18946 33346
rect 18946 33294 18948 33346
rect 18892 33292 18948 33294
rect 19052 33292 19108 33348
rect 19372 33292 19428 33348
rect 23132 33346 23188 33348
rect 23132 33294 23134 33346
rect 23134 33294 23186 33346
rect 23186 33294 23188 33346
rect 23132 33292 23188 33294
rect 23292 33346 23348 33348
rect 23292 33294 23294 33346
rect 23294 33294 23346 33346
rect 23346 33294 23348 33346
rect 23292 33292 23348 33294
rect 23452 33346 23508 33348
rect 23452 33294 23454 33346
rect 23454 33294 23506 33346
rect 23506 33294 23508 33346
rect 23452 33292 23508 33294
rect 23612 33346 23668 33348
rect 23612 33294 23614 33346
rect 23614 33294 23666 33346
rect 23666 33294 23668 33346
rect 23612 33292 23668 33294
rect 23772 33346 23828 33348
rect 23772 33294 23774 33346
rect 23774 33294 23826 33346
rect 23826 33294 23828 33346
rect 23772 33292 23828 33294
rect 23932 33346 23988 33348
rect 23932 33294 23934 33346
rect 23934 33294 23986 33346
rect 23986 33294 23988 33346
rect 23932 33292 23988 33294
rect 24092 33346 24148 33348
rect 24092 33294 24094 33346
rect 24094 33294 24146 33346
rect 24146 33294 24148 33346
rect 24092 33292 24148 33294
rect 24252 33346 24308 33348
rect 24252 33294 24254 33346
rect 24254 33294 24306 33346
rect 24306 33294 24308 33346
rect 24252 33292 24308 33294
rect 24412 33346 24468 33348
rect 24412 33294 24414 33346
rect 24414 33294 24466 33346
rect 24466 33294 24468 33346
rect 24412 33292 24468 33294
rect 24572 33346 24628 33348
rect 24572 33294 24574 33346
rect 24574 33294 24626 33346
rect 24626 33294 24628 33346
rect 24572 33292 24628 33294
rect 24732 33346 24788 33348
rect 24732 33294 24734 33346
rect 24734 33294 24786 33346
rect 24786 33294 24788 33346
rect 24732 33292 24788 33294
rect 24892 33346 24948 33348
rect 24892 33294 24894 33346
rect 24894 33294 24946 33346
rect 24946 33294 24948 33346
rect 24892 33292 24948 33294
rect 25052 33346 25108 33348
rect 25052 33294 25054 33346
rect 25054 33294 25106 33346
rect 25106 33294 25108 33346
rect 25052 33292 25108 33294
rect 25212 33346 25268 33348
rect 25212 33294 25214 33346
rect 25214 33294 25266 33346
rect 25266 33294 25268 33346
rect 25212 33292 25268 33294
rect 25372 33346 25428 33348
rect 25372 33294 25374 33346
rect 25374 33294 25426 33346
rect 25426 33294 25428 33346
rect 25372 33292 25428 33294
rect 25532 33346 25588 33348
rect 25532 33294 25534 33346
rect 25534 33294 25586 33346
rect 25586 33294 25588 33346
rect 25532 33292 25588 33294
rect 25692 33346 25748 33348
rect 25692 33294 25694 33346
rect 25694 33294 25746 33346
rect 25746 33294 25748 33346
rect 25692 33292 25748 33294
rect 25852 33346 25908 33348
rect 25852 33294 25854 33346
rect 25854 33294 25906 33346
rect 25906 33294 25908 33346
rect 25852 33292 25908 33294
rect 26012 33346 26068 33348
rect 26012 33294 26014 33346
rect 26014 33294 26066 33346
rect 26066 33294 26068 33346
rect 26012 33292 26068 33294
rect 26172 33346 26228 33348
rect 26172 33294 26174 33346
rect 26174 33294 26226 33346
rect 26226 33294 26228 33346
rect 26172 33292 26228 33294
rect 26332 33346 26388 33348
rect 26332 33294 26334 33346
rect 26334 33294 26386 33346
rect 26386 33294 26388 33346
rect 26332 33292 26388 33294
rect 26492 33346 26548 33348
rect 26492 33294 26494 33346
rect 26494 33294 26546 33346
rect 26546 33294 26548 33346
rect 26492 33292 26548 33294
rect 26652 33346 26708 33348
rect 26652 33294 26654 33346
rect 26654 33294 26706 33346
rect 26706 33294 26708 33346
rect 26652 33292 26708 33294
rect 26812 33346 26868 33348
rect 26812 33294 26814 33346
rect 26814 33294 26866 33346
rect 26866 33294 26868 33346
rect 26812 33292 26868 33294
rect 26972 33346 27028 33348
rect 26972 33294 26974 33346
rect 26974 33294 27026 33346
rect 27026 33294 27028 33346
rect 26972 33292 27028 33294
rect 27132 33346 27188 33348
rect 27132 33294 27134 33346
rect 27134 33294 27186 33346
rect 27186 33294 27188 33346
rect 27132 33292 27188 33294
rect 27292 33346 27348 33348
rect 27292 33294 27294 33346
rect 27294 33294 27346 33346
rect 27346 33294 27348 33346
rect 27292 33292 27348 33294
rect 27452 33346 27508 33348
rect 27452 33294 27454 33346
rect 27454 33294 27506 33346
rect 27506 33294 27508 33346
rect 27452 33292 27508 33294
rect 27612 33346 27668 33348
rect 27612 33294 27614 33346
rect 27614 33294 27666 33346
rect 27666 33294 27668 33346
rect 27612 33292 27668 33294
rect 27772 33346 27828 33348
rect 27772 33294 27774 33346
rect 27774 33294 27826 33346
rect 27826 33294 27828 33346
rect 27772 33292 27828 33294
rect 27932 33346 27988 33348
rect 27932 33294 27934 33346
rect 27934 33294 27986 33346
rect 27986 33294 27988 33346
rect 27932 33292 27988 33294
rect 28092 33346 28148 33348
rect 28092 33294 28094 33346
rect 28094 33294 28146 33346
rect 28146 33294 28148 33346
rect 28092 33292 28148 33294
rect 28252 33346 28308 33348
rect 28252 33294 28254 33346
rect 28254 33294 28306 33346
rect 28306 33294 28308 33346
rect 28252 33292 28308 33294
rect 28412 33346 28468 33348
rect 28412 33294 28414 33346
rect 28414 33294 28466 33346
rect 28466 33294 28468 33346
rect 28412 33292 28468 33294
rect 28572 33346 28628 33348
rect 28572 33294 28574 33346
rect 28574 33294 28626 33346
rect 28626 33294 28628 33346
rect 28572 33292 28628 33294
rect 28732 33346 28788 33348
rect 28732 33294 28734 33346
rect 28734 33294 28786 33346
rect 28786 33294 28788 33346
rect 28732 33292 28788 33294
rect 28892 33346 28948 33348
rect 28892 33294 28894 33346
rect 28894 33294 28946 33346
rect 28946 33294 28948 33346
rect 28892 33292 28948 33294
rect 29052 33346 29108 33348
rect 29052 33294 29054 33346
rect 29054 33294 29106 33346
rect 29106 33294 29108 33346
rect 29052 33292 29108 33294
rect 29212 33346 29268 33348
rect 29212 33294 29214 33346
rect 29214 33294 29266 33346
rect 29266 33294 29268 33346
rect 29212 33292 29268 33294
rect 29372 33346 29428 33348
rect 29372 33294 29374 33346
rect 29374 33294 29426 33346
rect 29426 33294 29428 33346
rect 29372 33292 29428 33294
rect 33052 33292 33108 33348
rect 33372 33292 33428 33348
rect 33532 33346 33588 33348
rect 33532 33294 33534 33346
rect 33534 33294 33586 33346
rect 33586 33294 33588 33346
rect 33532 33292 33588 33294
rect 33692 33346 33748 33348
rect 33692 33294 33694 33346
rect 33694 33294 33746 33346
rect 33746 33294 33748 33346
rect 33692 33292 33748 33294
rect 33852 33346 33908 33348
rect 33852 33294 33854 33346
rect 33854 33294 33906 33346
rect 33906 33294 33908 33346
rect 33852 33292 33908 33294
rect 34012 33346 34068 33348
rect 34012 33294 34014 33346
rect 34014 33294 34066 33346
rect 34066 33294 34068 33346
rect 34012 33292 34068 33294
rect 34172 33346 34228 33348
rect 34172 33294 34174 33346
rect 34174 33294 34226 33346
rect 34226 33294 34228 33346
rect 34172 33292 34228 33294
rect 34332 33346 34388 33348
rect 34332 33294 34334 33346
rect 34334 33294 34386 33346
rect 34386 33294 34388 33346
rect 34332 33292 34388 33294
rect 34492 33346 34548 33348
rect 34492 33294 34494 33346
rect 34494 33294 34546 33346
rect 34546 33294 34548 33346
rect 34492 33292 34548 33294
rect 34652 33346 34708 33348
rect 34652 33294 34654 33346
rect 34654 33294 34706 33346
rect 34706 33294 34708 33346
rect 34652 33292 34708 33294
rect 34812 33346 34868 33348
rect 34812 33294 34814 33346
rect 34814 33294 34866 33346
rect 34866 33294 34868 33346
rect 34812 33292 34868 33294
rect 34972 33346 35028 33348
rect 34972 33294 34974 33346
rect 34974 33294 35026 33346
rect 35026 33294 35028 33346
rect 34972 33292 35028 33294
rect 35132 33346 35188 33348
rect 35132 33294 35134 33346
rect 35134 33294 35186 33346
rect 35186 33294 35188 33346
rect 35132 33292 35188 33294
rect 35292 33346 35348 33348
rect 35292 33294 35294 33346
rect 35294 33294 35346 33346
rect 35346 33294 35348 33346
rect 35292 33292 35348 33294
rect 35452 33346 35508 33348
rect 35452 33294 35454 33346
rect 35454 33294 35506 33346
rect 35506 33294 35508 33346
rect 35452 33292 35508 33294
rect 35612 33346 35668 33348
rect 35612 33294 35614 33346
rect 35614 33294 35666 33346
rect 35666 33294 35668 33346
rect 35612 33292 35668 33294
rect 35772 33346 35828 33348
rect 35772 33294 35774 33346
rect 35774 33294 35826 33346
rect 35826 33294 35828 33346
rect 35772 33292 35828 33294
rect 35932 33346 35988 33348
rect 35932 33294 35934 33346
rect 35934 33294 35986 33346
rect 35986 33294 35988 33346
rect 35932 33292 35988 33294
rect 36092 33346 36148 33348
rect 36092 33294 36094 33346
rect 36094 33294 36146 33346
rect 36146 33294 36148 33346
rect 36092 33292 36148 33294
rect 36252 33346 36308 33348
rect 36252 33294 36254 33346
rect 36254 33294 36306 33346
rect 36306 33294 36308 33346
rect 36252 33292 36308 33294
rect 36412 33346 36468 33348
rect 36412 33294 36414 33346
rect 36414 33294 36466 33346
rect 36466 33294 36468 33346
rect 36412 33292 36468 33294
rect 36572 33346 36628 33348
rect 36572 33294 36574 33346
rect 36574 33294 36626 33346
rect 36626 33294 36628 33346
rect 36572 33292 36628 33294
rect 36732 33346 36788 33348
rect 36732 33294 36734 33346
rect 36734 33294 36786 33346
rect 36786 33294 36788 33346
rect 36732 33292 36788 33294
rect 36892 33346 36948 33348
rect 36892 33294 36894 33346
rect 36894 33294 36946 33346
rect 36946 33294 36948 33346
rect 36892 33292 36948 33294
rect 37052 33346 37108 33348
rect 37052 33294 37054 33346
rect 37054 33294 37106 33346
rect 37106 33294 37108 33346
rect 37052 33292 37108 33294
rect 37212 33346 37268 33348
rect 37212 33294 37214 33346
rect 37214 33294 37266 33346
rect 37266 33294 37268 33346
rect 37212 33292 37268 33294
rect 37372 33346 37428 33348
rect 37372 33294 37374 33346
rect 37374 33294 37426 33346
rect 37426 33294 37428 33346
rect 37372 33292 37428 33294
rect 37532 33346 37588 33348
rect 37532 33294 37534 33346
rect 37534 33294 37586 33346
rect 37586 33294 37588 33346
rect 37532 33292 37588 33294
rect 37692 33346 37748 33348
rect 37692 33294 37694 33346
rect 37694 33294 37746 33346
rect 37746 33294 37748 33346
rect 37692 33292 37748 33294
rect 37852 33346 37908 33348
rect 37852 33294 37854 33346
rect 37854 33294 37906 33346
rect 37906 33294 37908 33346
rect 37852 33292 37908 33294
rect 38012 33346 38068 33348
rect 38012 33294 38014 33346
rect 38014 33294 38066 33346
rect 38066 33294 38068 33346
rect 38012 33292 38068 33294
rect 38172 33346 38228 33348
rect 38172 33294 38174 33346
rect 38174 33294 38226 33346
rect 38226 33294 38228 33346
rect 38172 33292 38228 33294
rect 38332 33346 38388 33348
rect 38332 33294 38334 33346
rect 38334 33294 38386 33346
rect 38386 33294 38388 33346
rect 38332 33292 38388 33294
rect 38492 33346 38548 33348
rect 38492 33294 38494 33346
rect 38494 33294 38546 33346
rect 38546 33294 38548 33346
rect 38492 33292 38548 33294
rect 38652 33346 38708 33348
rect 38652 33294 38654 33346
rect 38654 33294 38706 33346
rect 38706 33294 38708 33346
rect 38652 33292 38708 33294
rect 38812 33346 38868 33348
rect 38812 33294 38814 33346
rect 38814 33294 38866 33346
rect 38866 33294 38868 33346
rect 38812 33292 38868 33294
rect 38972 33346 39028 33348
rect 38972 33294 38974 33346
rect 38974 33294 39026 33346
rect 39026 33294 39028 33346
rect 38972 33292 39028 33294
rect 39132 33346 39188 33348
rect 39132 33294 39134 33346
rect 39134 33294 39186 33346
rect 39186 33294 39188 33346
rect 39132 33292 39188 33294
rect 39292 33346 39348 33348
rect 39292 33294 39294 33346
rect 39294 33294 39346 33346
rect 39346 33294 39348 33346
rect 39292 33292 39348 33294
rect 39452 33346 39508 33348
rect 39452 33294 39454 33346
rect 39454 33294 39506 33346
rect 39506 33294 39508 33346
rect 39452 33292 39508 33294
rect 39612 33346 39668 33348
rect 39612 33294 39614 33346
rect 39614 33294 39666 33346
rect 39666 33294 39668 33346
rect 39612 33292 39668 33294
rect 39772 33346 39828 33348
rect 39772 33294 39774 33346
rect 39774 33294 39826 33346
rect 39826 33294 39828 33346
rect 39772 33292 39828 33294
rect 39932 33346 39988 33348
rect 39932 33294 39934 33346
rect 39934 33294 39986 33346
rect 39986 33294 39988 33346
rect 39932 33292 39988 33294
rect 40092 33346 40148 33348
rect 40092 33294 40094 33346
rect 40094 33294 40146 33346
rect 40146 33294 40148 33346
rect 40092 33292 40148 33294
rect 40252 33346 40308 33348
rect 40252 33294 40254 33346
rect 40254 33294 40306 33346
rect 40306 33294 40308 33346
rect 40252 33292 40308 33294
rect 40412 33346 40468 33348
rect 40412 33294 40414 33346
rect 40414 33294 40466 33346
rect 40466 33294 40468 33346
rect 40412 33292 40468 33294
rect 40572 33346 40628 33348
rect 40572 33294 40574 33346
rect 40574 33294 40626 33346
rect 40626 33294 40628 33346
rect 40572 33292 40628 33294
rect 40732 33346 40788 33348
rect 40732 33294 40734 33346
rect 40734 33294 40786 33346
rect 40786 33294 40788 33346
rect 40732 33292 40788 33294
rect 40892 33346 40948 33348
rect 40892 33294 40894 33346
rect 40894 33294 40946 33346
rect 40946 33294 40948 33346
rect 40892 33292 40948 33294
rect 41052 33346 41108 33348
rect 41052 33294 41054 33346
rect 41054 33294 41106 33346
rect 41106 33294 41108 33346
rect 41052 33292 41108 33294
rect 41212 33346 41268 33348
rect 41212 33294 41214 33346
rect 41214 33294 41266 33346
rect 41266 33294 41268 33346
rect 41212 33292 41268 33294
rect 41372 33346 41428 33348
rect 41372 33294 41374 33346
rect 41374 33294 41426 33346
rect 41426 33294 41428 33346
rect 41372 33292 41428 33294
rect 41532 33346 41588 33348
rect 41532 33294 41534 33346
rect 41534 33294 41586 33346
rect 41586 33294 41588 33346
rect 41532 33292 41588 33294
rect 41692 33346 41748 33348
rect 41692 33294 41694 33346
rect 41694 33294 41746 33346
rect 41746 33294 41748 33346
rect 41692 33292 41748 33294
rect 41852 33346 41908 33348
rect 41852 33294 41854 33346
rect 41854 33294 41906 33346
rect 41906 33294 41908 33346
rect 41852 33292 41908 33294
rect 8652 33132 8708 33188
rect 19212 33132 19268 33188
rect 33212 33132 33268 33188
rect 12 33026 68 33028
rect 12 32974 14 33026
rect 14 32974 66 33026
rect 66 32974 68 33026
rect 12 32972 68 32974
rect 172 33026 228 33028
rect 172 32974 174 33026
rect 174 32974 226 33026
rect 226 32974 228 33026
rect 172 32972 228 32974
rect 332 33026 388 33028
rect 332 32974 334 33026
rect 334 32974 386 33026
rect 386 32974 388 33026
rect 332 32972 388 32974
rect 492 33026 548 33028
rect 492 32974 494 33026
rect 494 32974 546 33026
rect 546 32974 548 33026
rect 492 32972 548 32974
rect 652 33026 708 33028
rect 652 32974 654 33026
rect 654 32974 706 33026
rect 706 32974 708 33026
rect 652 32972 708 32974
rect 812 33026 868 33028
rect 812 32974 814 33026
rect 814 32974 866 33026
rect 866 32974 868 33026
rect 812 32972 868 32974
rect 972 33026 1028 33028
rect 972 32974 974 33026
rect 974 32974 1026 33026
rect 1026 32974 1028 33026
rect 972 32972 1028 32974
rect 1132 33026 1188 33028
rect 1132 32974 1134 33026
rect 1134 32974 1186 33026
rect 1186 32974 1188 33026
rect 1132 32972 1188 32974
rect 1292 33026 1348 33028
rect 1292 32974 1294 33026
rect 1294 32974 1346 33026
rect 1346 32974 1348 33026
rect 1292 32972 1348 32974
rect 1452 33026 1508 33028
rect 1452 32974 1454 33026
rect 1454 32974 1506 33026
rect 1506 32974 1508 33026
rect 1452 32972 1508 32974
rect 1612 33026 1668 33028
rect 1612 32974 1614 33026
rect 1614 32974 1666 33026
rect 1666 32974 1668 33026
rect 1612 32972 1668 32974
rect 1772 33026 1828 33028
rect 1772 32974 1774 33026
rect 1774 32974 1826 33026
rect 1826 32974 1828 33026
rect 1772 32972 1828 32974
rect 1932 33026 1988 33028
rect 1932 32974 1934 33026
rect 1934 32974 1986 33026
rect 1986 32974 1988 33026
rect 1932 32972 1988 32974
rect 2092 33026 2148 33028
rect 2092 32974 2094 33026
rect 2094 32974 2146 33026
rect 2146 32974 2148 33026
rect 2092 32972 2148 32974
rect 2252 33026 2308 33028
rect 2252 32974 2254 33026
rect 2254 32974 2306 33026
rect 2306 32974 2308 33026
rect 2252 32972 2308 32974
rect 2412 33026 2468 33028
rect 2412 32974 2414 33026
rect 2414 32974 2466 33026
rect 2466 32974 2468 33026
rect 2412 32972 2468 32974
rect 2572 33026 2628 33028
rect 2572 32974 2574 33026
rect 2574 32974 2626 33026
rect 2626 32974 2628 33026
rect 2572 32972 2628 32974
rect 2732 33026 2788 33028
rect 2732 32974 2734 33026
rect 2734 32974 2786 33026
rect 2786 32974 2788 33026
rect 2732 32972 2788 32974
rect 2892 33026 2948 33028
rect 2892 32974 2894 33026
rect 2894 32974 2946 33026
rect 2946 32974 2948 33026
rect 2892 32972 2948 32974
rect 3052 33026 3108 33028
rect 3052 32974 3054 33026
rect 3054 32974 3106 33026
rect 3106 32974 3108 33026
rect 3052 32972 3108 32974
rect 3212 33026 3268 33028
rect 3212 32974 3214 33026
rect 3214 32974 3266 33026
rect 3266 32974 3268 33026
rect 3212 32972 3268 32974
rect 3372 33026 3428 33028
rect 3372 32974 3374 33026
rect 3374 32974 3426 33026
rect 3426 32974 3428 33026
rect 3372 32972 3428 32974
rect 3532 33026 3588 33028
rect 3532 32974 3534 33026
rect 3534 32974 3586 33026
rect 3586 32974 3588 33026
rect 3532 32972 3588 32974
rect 3692 33026 3748 33028
rect 3692 32974 3694 33026
rect 3694 32974 3746 33026
rect 3746 32974 3748 33026
rect 3692 32972 3748 32974
rect 3852 33026 3908 33028
rect 3852 32974 3854 33026
rect 3854 32974 3906 33026
rect 3906 32974 3908 33026
rect 3852 32972 3908 32974
rect 4012 33026 4068 33028
rect 4012 32974 4014 33026
rect 4014 32974 4066 33026
rect 4066 32974 4068 33026
rect 4012 32972 4068 32974
rect 4172 33026 4228 33028
rect 4172 32974 4174 33026
rect 4174 32974 4226 33026
rect 4226 32974 4228 33026
rect 4172 32972 4228 32974
rect 4332 33026 4388 33028
rect 4332 32974 4334 33026
rect 4334 32974 4386 33026
rect 4386 32974 4388 33026
rect 4332 32972 4388 32974
rect 4492 33026 4548 33028
rect 4492 32974 4494 33026
rect 4494 32974 4546 33026
rect 4546 32974 4548 33026
rect 4492 32972 4548 32974
rect 4652 33026 4708 33028
rect 4652 32974 4654 33026
rect 4654 32974 4706 33026
rect 4706 32974 4708 33026
rect 4652 32972 4708 32974
rect 4812 33026 4868 33028
rect 4812 32974 4814 33026
rect 4814 32974 4866 33026
rect 4866 32974 4868 33026
rect 4812 32972 4868 32974
rect 4972 33026 5028 33028
rect 4972 32974 4974 33026
rect 4974 32974 5026 33026
rect 5026 32974 5028 33026
rect 4972 32972 5028 32974
rect 5132 33026 5188 33028
rect 5132 32974 5134 33026
rect 5134 32974 5186 33026
rect 5186 32974 5188 33026
rect 5132 32972 5188 32974
rect 5292 33026 5348 33028
rect 5292 32974 5294 33026
rect 5294 32974 5346 33026
rect 5346 32974 5348 33026
rect 5292 32972 5348 32974
rect 5452 33026 5508 33028
rect 5452 32974 5454 33026
rect 5454 32974 5506 33026
rect 5506 32974 5508 33026
rect 5452 32972 5508 32974
rect 5612 33026 5668 33028
rect 5612 32974 5614 33026
rect 5614 32974 5666 33026
rect 5666 32974 5668 33026
rect 5612 32972 5668 32974
rect 5772 33026 5828 33028
rect 5772 32974 5774 33026
rect 5774 32974 5826 33026
rect 5826 32974 5828 33026
rect 5772 32972 5828 32974
rect 5932 33026 5988 33028
rect 5932 32974 5934 33026
rect 5934 32974 5986 33026
rect 5986 32974 5988 33026
rect 5932 32972 5988 32974
rect 6092 33026 6148 33028
rect 6092 32974 6094 33026
rect 6094 32974 6146 33026
rect 6146 32974 6148 33026
rect 6092 32972 6148 32974
rect 6252 33026 6308 33028
rect 6252 32974 6254 33026
rect 6254 32974 6306 33026
rect 6306 32974 6308 33026
rect 6252 32972 6308 32974
rect 6412 33026 6468 33028
rect 6412 32974 6414 33026
rect 6414 32974 6466 33026
rect 6466 32974 6468 33026
rect 6412 32972 6468 32974
rect 6572 33026 6628 33028
rect 6572 32974 6574 33026
rect 6574 32974 6626 33026
rect 6626 32974 6628 33026
rect 6572 32972 6628 32974
rect 6732 33026 6788 33028
rect 6732 32974 6734 33026
rect 6734 32974 6786 33026
rect 6786 32974 6788 33026
rect 6732 32972 6788 32974
rect 6892 33026 6948 33028
rect 6892 32974 6894 33026
rect 6894 32974 6946 33026
rect 6946 32974 6948 33026
rect 6892 32972 6948 32974
rect 7052 33026 7108 33028
rect 7052 32974 7054 33026
rect 7054 32974 7106 33026
rect 7106 32974 7108 33026
rect 7052 32972 7108 32974
rect 7212 33026 7268 33028
rect 7212 32974 7214 33026
rect 7214 32974 7266 33026
rect 7266 32974 7268 33026
rect 7212 32972 7268 32974
rect 7372 33026 7428 33028
rect 7372 32974 7374 33026
rect 7374 32974 7426 33026
rect 7426 32974 7428 33026
rect 7372 32972 7428 32974
rect 7532 33026 7588 33028
rect 7532 32974 7534 33026
rect 7534 32974 7586 33026
rect 7586 32974 7588 33026
rect 7532 32972 7588 32974
rect 7692 33026 7748 33028
rect 7692 32974 7694 33026
rect 7694 32974 7746 33026
rect 7746 32974 7748 33026
rect 7692 32972 7748 32974
rect 7852 33026 7908 33028
rect 7852 32974 7854 33026
rect 7854 32974 7906 33026
rect 7906 32974 7908 33026
rect 7852 32972 7908 32974
rect 8012 33026 8068 33028
rect 8012 32974 8014 33026
rect 8014 32974 8066 33026
rect 8066 32974 8068 33026
rect 8012 32972 8068 32974
rect 8172 33026 8228 33028
rect 8172 32974 8174 33026
rect 8174 32974 8226 33026
rect 8226 32974 8228 33026
rect 8172 32972 8228 32974
rect 8332 33026 8388 33028
rect 8332 32974 8334 33026
rect 8334 32974 8386 33026
rect 8386 32974 8388 33026
rect 8332 32972 8388 32974
rect 8492 32972 8548 33028
rect 8812 32972 8868 33028
rect 12492 33026 12548 33028
rect 12492 32974 12494 33026
rect 12494 32974 12546 33026
rect 12546 32974 12548 33026
rect 12492 32972 12548 32974
rect 12652 33026 12708 33028
rect 12652 32974 12654 33026
rect 12654 32974 12706 33026
rect 12706 32974 12708 33026
rect 12652 32972 12708 32974
rect 12812 33026 12868 33028
rect 12812 32974 12814 33026
rect 12814 32974 12866 33026
rect 12866 32974 12868 33026
rect 12812 32972 12868 32974
rect 12972 33026 13028 33028
rect 12972 32974 12974 33026
rect 12974 32974 13026 33026
rect 13026 32974 13028 33026
rect 12972 32972 13028 32974
rect 13132 33026 13188 33028
rect 13132 32974 13134 33026
rect 13134 32974 13186 33026
rect 13186 32974 13188 33026
rect 13132 32972 13188 32974
rect 13292 33026 13348 33028
rect 13292 32974 13294 33026
rect 13294 32974 13346 33026
rect 13346 32974 13348 33026
rect 13292 32972 13348 32974
rect 13452 33026 13508 33028
rect 13452 32974 13454 33026
rect 13454 32974 13506 33026
rect 13506 32974 13508 33026
rect 13452 32972 13508 32974
rect 13612 33026 13668 33028
rect 13612 32974 13614 33026
rect 13614 32974 13666 33026
rect 13666 32974 13668 33026
rect 13612 32972 13668 32974
rect 13772 33026 13828 33028
rect 13772 32974 13774 33026
rect 13774 32974 13826 33026
rect 13826 32974 13828 33026
rect 13772 32972 13828 32974
rect 13932 33026 13988 33028
rect 13932 32974 13934 33026
rect 13934 32974 13986 33026
rect 13986 32974 13988 33026
rect 13932 32972 13988 32974
rect 14092 33026 14148 33028
rect 14092 32974 14094 33026
rect 14094 32974 14146 33026
rect 14146 32974 14148 33026
rect 14092 32972 14148 32974
rect 14252 33026 14308 33028
rect 14252 32974 14254 33026
rect 14254 32974 14306 33026
rect 14306 32974 14308 33026
rect 14252 32972 14308 32974
rect 14412 33026 14468 33028
rect 14412 32974 14414 33026
rect 14414 32974 14466 33026
rect 14466 32974 14468 33026
rect 14412 32972 14468 32974
rect 14572 33026 14628 33028
rect 14572 32974 14574 33026
rect 14574 32974 14626 33026
rect 14626 32974 14628 33026
rect 14572 32972 14628 32974
rect 14732 33026 14788 33028
rect 14732 32974 14734 33026
rect 14734 32974 14786 33026
rect 14786 32974 14788 33026
rect 14732 32972 14788 32974
rect 14892 33026 14948 33028
rect 14892 32974 14894 33026
rect 14894 32974 14946 33026
rect 14946 32974 14948 33026
rect 14892 32972 14948 32974
rect 15052 33026 15108 33028
rect 15052 32974 15054 33026
rect 15054 32974 15106 33026
rect 15106 32974 15108 33026
rect 15052 32972 15108 32974
rect 15212 33026 15268 33028
rect 15212 32974 15214 33026
rect 15214 32974 15266 33026
rect 15266 32974 15268 33026
rect 15212 32972 15268 32974
rect 15372 33026 15428 33028
rect 15372 32974 15374 33026
rect 15374 32974 15426 33026
rect 15426 32974 15428 33026
rect 15372 32972 15428 32974
rect 15532 33026 15588 33028
rect 15532 32974 15534 33026
rect 15534 32974 15586 33026
rect 15586 32974 15588 33026
rect 15532 32972 15588 32974
rect 15692 33026 15748 33028
rect 15692 32974 15694 33026
rect 15694 32974 15746 33026
rect 15746 32974 15748 33026
rect 15692 32972 15748 32974
rect 15852 33026 15908 33028
rect 15852 32974 15854 33026
rect 15854 32974 15906 33026
rect 15906 32974 15908 33026
rect 15852 32972 15908 32974
rect 16012 33026 16068 33028
rect 16012 32974 16014 33026
rect 16014 32974 16066 33026
rect 16066 32974 16068 33026
rect 16012 32972 16068 32974
rect 16172 33026 16228 33028
rect 16172 32974 16174 33026
rect 16174 32974 16226 33026
rect 16226 32974 16228 33026
rect 16172 32972 16228 32974
rect 16332 33026 16388 33028
rect 16332 32974 16334 33026
rect 16334 32974 16386 33026
rect 16386 32974 16388 33026
rect 16332 32972 16388 32974
rect 16492 33026 16548 33028
rect 16492 32974 16494 33026
rect 16494 32974 16546 33026
rect 16546 32974 16548 33026
rect 16492 32972 16548 32974
rect 16652 33026 16708 33028
rect 16652 32974 16654 33026
rect 16654 32974 16706 33026
rect 16706 32974 16708 33026
rect 16652 32972 16708 32974
rect 16812 33026 16868 33028
rect 16812 32974 16814 33026
rect 16814 32974 16866 33026
rect 16866 32974 16868 33026
rect 16812 32972 16868 32974
rect 16972 33026 17028 33028
rect 16972 32974 16974 33026
rect 16974 32974 17026 33026
rect 17026 32974 17028 33026
rect 16972 32972 17028 32974
rect 17132 33026 17188 33028
rect 17132 32974 17134 33026
rect 17134 32974 17186 33026
rect 17186 32974 17188 33026
rect 17132 32972 17188 32974
rect 17292 33026 17348 33028
rect 17292 32974 17294 33026
rect 17294 32974 17346 33026
rect 17346 32974 17348 33026
rect 17292 32972 17348 32974
rect 17452 33026 17508 33028
rect 17452 32974 17454 33026
rect 17454 32974 17506 33026
rect 17506 32974 17508 33026
rect 17452 32972 17508 32974
rect 17612 33026 17668 33028
rect 17612 32974 17614 33026
rect 17614 32974 17666 33026
rect 17666 32974 17668 33026
rect 17612 32972 17668 32974
rect 17772 33026 17828 33028
rect 17772 32974 17774 33026
rect 17774 32974 17826 33026
rect 17826 32974 17828 33026
rect 17772 32972 17828 32974
rect 17932 33026 17988 33028
rect 17932 32974 17934 33026
rect 17934 32974 17986 33026
rect 17986 32974 17988 33026
rect 17932 32972 17988 32974
rect 18092 33026 18148 33028
rect 18092 32974 18094 33026
rect 18094 32974 18146 33026
rect 18146 32974 18148 33026
rect 18092 32972 18148 32974
rect 18252 33026 18308 33028
rect 18252 32974 18254 33026
rect 18254 32974 18306 33026
rect 18306 32974 18308 33026
rect 18252 32972 18308 32974
rect 18412 33026 18468 33028
rect 18412 32974 18414 33026
rect 18414 32974 18466 33026
rect 18466 32974 18468 33026
rect 18412 32972 18468 32974
rect 18572 33026 18628 33028
rect 18572 32974 18574 33026
rect 18574 32974 18626 33026
rect 18626 32974 18628 33026
rect 18572 32972 18628 32974
rect 18732 33026 18788 33028
rect 18732 32974 18734 33026
rect 18734 32974 18786 33026
rect 18786 32974 18788 33026
rect 18732 32972 18788 32974
rect 18892 33026 18948 33028
rect 18892 32974 18894 33026
rect 18894 32974 18946 33026
rect 18946 32974 18948 33026
rect 18892 32972 18948 32974
rect 19052 32972 19108 33028
rect 19372 32972 19428 33028
rect 23132 33026 23188 33028
rect 23132 32974 23134 33026
rect 23134 32974 23186 33026
rect 23186 32974 23188 33026
rect 23132 32972 23188 32974
rect 23292 33026 23348 33028
rect 23292 32974 23294 33026
rect 23294 32974 23346 33026
rect 23346 32974 23348 33026
rect 23292 32972 23348 32974
rect 23452 33026 23508 33028
rect 23452 32974 23454 33026
rect 23454 32974 23506 33026
rect 23506 32974 23508 33026
rect 23452 32972 23508 32974
rect 23612 33026 23668 33028
rect 23612 32974 23614 33026
rect 23614 32974 23666 33026
rect 23666 32974 23668 33026
rect 23612 32972 23668 32974
rect 23772 33026 23828 33028
rect 23772 32974 23774 33026
rect 23774 32974 23826 33026
rect 23826 32974 23828 33026
rect 23772 32972 23828 32974
rect 23932 33026 23988 33028
rect 23932 32974 23934 33026
rect 23934 32974 23986 33026
rect 23986 32974 23988 33026
rect 23932 32972 23988 32974
rect 24092 33026 24148 33028
rect 24092 32974 24094 33026
rect 24094 32974 24146 33026
rect 24146 32974 24148 33026
rect 24092 32972 24148 32974
rect 24252 33026 24308 33028
rect 24252 32974 24254 33026
rect 24254 32974 24306 33026
rect 24306 32974 24308 33026
rect 24252 32972 24308 32974
rect 24412 33026 24468 33028
rect 24412 32974 24414 33026
rect 24414 32974 24466 33026
rect 24466 32974 24468 33026
rect 24412 32972 24468 32974
rect 24572 33026 24628 33028
rect 24572 32974 24574 33026
rect 24574 32974 24626 33026
rect 24626 32974 24628 33026
rect 24572 32972 24628 32974
rect 24732 33026 24788 33028
rect 24732 32974 24734 33026
rect 24734 32974 24786 33026
rect 24786 32974 24788 33026
rect 24732 32972 24788 32974
rect 24892 33026 24948 33028
rect 24892 32974 24894 33026
rect 24894 32974 24946 33026
rect 24946 32974 24948 33026
rect 24892 32972 24948 32974
rect 25052 33026 25108 33028
rect 25052 32974 25054 33026
rect 25054 32974 25106 33026
rect 25106 32974 25108 33026
rect 25052 32972 25108 32974
rect 25212 33026 25268 33028
rect 25212 32974 25214 33026
rect 25214 32974 25266 33026
rect 25266 32974 25268 33026
rect 25212 32972 25268 32974
rect 25372 33026 25428 33028
rect 25372 32974 25374 33026
rect 25374 32974 25426 33026
rect 25426 32974 25428 33026
rect 25372 32972 25428 32974
rect 25532 33026 25588 33028
rect 25532 32974 25534 33026
rect 25534 32974 25586 33026
rect 25586 32974 25588 33026
rect 25532 32972 25588 32974
rect 25692 33026 25748 33028
rect 25692 32974 25694 33026
rect 25694 32974 25746 33026
rect 25746 32974 25748 33026
rect 25692 32972 25748 32974
rect 25852 33026 25908 33028
rect 25852 32974 25854 33026
rect 25854 32974 25906 33026
rect 25906 32974 25908 33026
rect 25852 32972 25908 32974
rect 26012 33026 26068 33028
rect 26012 32974 26014 33026
rect 26014 32974 26066 33026
rect 26066 32974 26068 33026
rect 26012 32972 26068 32974
rect 26172 33026 26228 33028
rect 26172 32974 26174 33026
rect 26174 32974 26226 33026
rect 26226 32974 26228 33026
rect 26172 32972 26228 32974
rect 26332 33026 26388 33028
rect 26332 32974 26334 33026
rect 26334 32974 26386 33026
rect 26386 32974 26388 33026
rect 26332 32972 26388 32974
rect 26492 33026 26548 33028
rect 26492 32974 26494 33026
rect 26494 32974 26546 33026
rect 26546 32974 26548 33026
rect 26492 32972 26548 32974
rect 26652 33026 26708 33028
rect 26652 32974 26654 33026
rect 26654 32974 26706 33026
rect 26706 32974 26708 33026
rect 26652 32972 26708 32974
rect 26812 33026 26868 33028
rect 26812 32974 26814 33026
rect 26814 32974 26866 33026
rect 26866 32974 26868 33026
rect 26812 32972 26868 32974
rect 26972 33026 27028 33028
rect 26972 32974 26974 33026
rect 26974 32974 27026 33026
rect 27026 32974 27028 33026
rect 26972 32972 27028 32974
rect 27132 33026 27188 33028
rect 27132 32974 27134 33026
rect 27134 32974 27186 33026
rect 27186 32974 27188 33026
rect 27132 32972 27188 32974
rect 27292 33026 27348 33028
rect 27292 32974 27294 33026
rect 27294 32974 27346 33026
rect 27346 32974 27348 33026
rect 27292 32972 27348 32974
rect 27452 33026 27508 33028
rect 27452 32974 27454 33026
rect 27454 32974 27506 33026
rect 27506 32974 27508 33026
rect 27452 32972 27508 32974
rect 27612 33026 27668 33028
rect 27612 32974 27614 33026
rect 27614 32974 27666 33026
rect 27666 32974 27668 33026
rect 27612 32972 27668 32974
rect 27772 33026 27828 33028
rect 27772 32974 27774 33026
rect 27774 32974 27826 33026
rect 27826 32974 27828 33026
rect 27772 32972 27828 32974
rect 27932 33026 27988 33028
rect 27932 32974 27934 33026
rect 27934 32974 27986 33026
rect 27986 32974 27988 33026
rect 27932 32972 27988 32974
rect 28092 33026 28148 33028
rect 28092 32974 28094 33026
rect 28094 32974 28146 33026
rect 28146 32974 28148 33026
rect 28092 32972 28148 32974
rect 28252 33026 28308 33028
rect 28252 32974 28254 33026
rect 28254 32974 28306 33026
rect 28306 32974 28308 33026
rect 28252 32972 28308 32974
rect 28412 33026 28468 33028
rect 28412 32974 28414 33026
rect 28414 32974 28466 33026
rect 28466 32974 28468 33026
rect 28412 32972 28468 32974
rect 28572 33026 28628 33028
rect 28572 32974 28574 33026
rect 28574 32974 28626 33026
rect 28626 32974 28628 33026
rect 28572 32972 28628 32974
rect 28732 33026 28788 33028
rect 28732 32974 28734 33026
rect 28734 32974 28786 33026
rect 28786 32974 28788 33026
rect 28732 32972 28788 32974
rect 28892 33026 28948 33028
rect 28892 32974 28894 33026
rect 28894 32974 28946 33026
rect 28946 32974 28948 33026
rect 28892 32972 28948 32974
rect 29052 33026 29108 33028
rect 29052 32974 29054 33026
rect 29054 32974 29106 33026
rect 29106 32974 29108 33026
rect 29052 32972 29108 32974
rect 29212 33026 29268 33028
rect 29212 32974 29214 33026
rect 29214 32974 29266 33026
rect 29266 32974 29268 33026
rect 29212 32972 29268 32974
rect 29372 33026 29428 33028
rect 29372 32974 29374 33026
rect 29374 32974 29426 33026
rect 29426 32974 29428 33026
rect 29372 32972 29428 32974
rect 33052 32972 33108 33028
rect 33372 32972 33428 33028
rect 33532 33026 33588 33028
rect 33532 32974 33534 33026
rect 33534 32974 33586 33026
rect 33586 32974 33588 33026
rect 33532 32972 33588 32974
rect 33692 33026 33748 33028
rect 33692 32974 33694 33026
rect 33694 32974 33746 33026
rect 33746 32974 33748 33026
rect 33692 32972 33748 32974
rect 33852 33026 33908 33028
rect 33852 32974 33854 33026
rect 33854 32974 33906 33026
rect 33906 32974 33908 33026
rect 33852 32972 33908 32974
rect 34012 33026 34068 33028
rect 34012 32974 34014 33026
rect 34014 32974 34066 33026
rect 34066 32974 34068 33026
rect 34012 32972 34068 32974
rect 34172 33026 34228 33028
rect 34172 32974 34174 33026
rect 34174 32974 34226 33026
rect 34226 32974 34228 33026
rect 34172 32972 34228 32974
rect 34332 33026 34388 33028
rect 34332 32974 34334 33026
rect 34334 32974 34386 33026
rect 34386 32974 34388 33026
rect 34332 32972 34388 32974
rect 34492 33026 34548 33028
rect 34492 32974 34494 33026
rect 34494 32974 34546 33026
rect 34546 32974 34548 33026
rect 34492 32972 34548 32974
rect 34652 33026 34708 33028
rect 34652 32974 34654 33026
rect 34654 32974 34706 33026
rect 34706 32974 34708 33026
rect 34652 32972 34708 32974
rect 34812 33026 34868 33028
rect 34812 32974 34814 33026
rect 34814 32974 34866 33026
rect 34866 32974 34868 33026
rect 34812 32972 34868 32974
rect 34972 33026 35028 33028
rect 34972 32974 34974 33026
rect 34974 32974 35026 33026
rect 35026 32974 35028 33026
rect 34972 32972 35028 32974
rect 35132 33026 35188 33028
rect 35132 32974 35134 33026
rect 35134 32974 35186 33026
rect 35186 32974 35188 33026
rect 35132 32972 35188 32974
rect 35292 33026 35348 33028
rect 35292 32974 35294 33026
rect 35294 32974 35346 33026
rect 35346 32974 35348 33026
rect 35292 32972 35348 32974
rect 35452 33026 35508 33028
rect 35452 32974 35454 33026
rect 35454 32974 35506 33026
rect 35506 32974 35508 33026
rect 35452 32972 35508 32974
rect 35612 33026 35668 33028
rect 35612 32974 35614 33026
rect 35614 32974 35666 33026
rect 35666 32974 35668 33026
rect 35612 32972 35668 32974
rect 35772 33026 35828 33028
rect 35772 32974 35774 33026
rect 35774 32974 35826 33026
rect 35826 32974 35828 33026
rect 35772 32972 35828 32974
rect 35932 33026 35988 33028
rect 35932 32974 35934 33026
rect 35934 32974 35986 33026
rect 35986 32974 35988 33026
rect 35932 32972 35988 32974
rect 36092 33026 36148 33028
rect 36092 32974 36094 33026
rect 36094 32974 36146 33026
rect 36146 32974 36148 33026
rect 36092 32972 36148 32974
rect 36252 33026 36308 33028
rect 36252 32974 36254 33026
rect 36254 32974 36306 33026
rect 36306 32974 36308 33026
rect 36252 32972 36308 32974
rect 36412 33026 36468 33028
rect 36412 32974 36414 33026
rect 36414 32974 36466 33026
rect 36466 32974 36468 33026
rect 36412 32972 36468 32974
rect 36572 33026 36628 33028
rect 36572 32974 36574 33026
rect 36574 32974 36626 33026
rect 36626 32974 36628 33026
rect 36572 32972 36628 32974
rect 36732 33026 36788 33028
rect 36732 32974 36734 33026
rect 36734 32974 36786 33026
rect 36786 32974 36788 33026
rect 36732 32972 36788 32974
rect 36892 33026 36948 33028
rect 36892 32974 36894 33026
rect 36894 32974 36946 33026
rect 36946 32974 36948 33026
rect 36892 32972 36948 32974
rect 37052 33026 37108 33028
rect 37052 32974 37054 33026
rect 37054 32974 37106 33026
rect 37106 32974 37108 33026
rect 37052 32972 37108 32974
rect 37212 33026 37268 33028
rect 37212 32974 37214 33026
rect 37214 32974 37266 33026
rect 37266 32974 37268 33026
rect 37212 32972 37268 32974
rect 37372 33026 37428 33028
rect 37372 32974 37374 33026
rect 37374 32974 37426 33026
rect 37426 32974 37428 33026
rect 37372 32972 37428 32974
rect 37532 33026 37588 33028
rect 37532 32974 37534 33026
rect 37534 32974 37586 33026
rect 37586 32974 37588 33026
rect 37532 32972 37588 32974
rect 37692 33026 37748 33028
rect 37692 32974 37694 33026
rect 37694 32974 37746 33026
rect 37746 32974 37748 33026
rect 37692 32972 37748 32974
rect 37852 33026 37908 33028
rect 37852 32974 37854 33026
rect 37854 32974 37906 33026
rect 37906 32974 37908 33026
rect 37852 32972 37908 32974
rect 38012 33026 38068 33028
rect 38012 32974 38014 33026
rect 38014 32974 38066 33026
rect 38066 32974 38068 33026
rect 38012 32972 38068 32974
rect 38172 33026 38228 33028
rect 38172 32974 38174 33026
rect 38174 32974 38226 33026
rect 38226 32974 38228 33026
rect 38172 32972 38228 32974
rect 38332 33026 38388 33028
rect 38332 32974 38334 33026
rect 38334 32974 38386 33026
rect 38386 32974 38388 33026
rect 38332 32972 38388 32974
rect 38492 33026 38548 33028
rect 38492 32974 38494 33026
rect 38494 32974 38546 33026
rect 38546 32974 38548 33026
rect 38492 32972 38548 32974
rect 38652 33026 38708 33028
rect 38652 32974 38654 33026
rect 38654 32974 38706 33026
rect 38706 32974 38708 33026
rect 38652 32972 38708 32974
rect 38812 33026 38868 33028
rect 38812 32974 38814 33026
rect 38814 32974 38866 33026
rect 38866 32974 38868 33026
rect 38812 32972 38868 32974
rect 38972 33026 39028 33028
rect 38972 32974 38974 33026
rect 38974 32974 39026 33026
rect 39026 32974 39028 33026
rect 38972 32972 39028 32974
rect 39132 33026 39188 33028
rect 39132 32974 39134 33026
rect 39134 32974 39186 33026
rect 39186 32974 39188 33026
rect 39132 32972 39188 32974
rect 39292 33026 39348 33028
rect 39292 32974 39294 33026
rect 39294 32974 39346 33026
rect 39346 32974 39348 33026
rect 39292 32972 39348 32974
rect 39452 33026 39508 33028
rect 39452 32974 39454 33026
rect 39454 32974 39506 33026
rect 39506 32974 39508 33026
rect 39452 32972 39508 32974
rect 39612 33026 39668 33028
rect 39612 32974 39614 33026
rect 39614 32974 39666 33026
rect 39666 32974 39668 33026
rect 39612 32972 39668 32974
rect 39772 33026 39828 33028
rect 39772 32974 39774 33026
rect 39774 32974 39826 33026
rect 39826 32974 39828 33026
rect 39772 32972 39828 32974
rect 39932 33026 39988 33028
rect 39932 32974 39934 33026
rect 39934 32974 39986 33026
rect 39986 32974 39988 33026
rect 39932 32972 39988 32974
rect 40092 33026 40148 33028
rect 40092 32974 40094 33026
rect 40094 32974 40146 33026
rect 40146 32974 40148 33026
rect 40092 32972 40148 32974
rect 40252 33026 40308 33028
rect 40252 32974 40254 33026
rect 40254 32974 40306 33026
rect 40306 32974 40308 33026
rect 40252 32972 40308 32974
rect 40412 33026 40468 33028
rect 40412 32974 40414 33026
rect 40414 32974 40466 33026
rect 40466 32974 40468 33026
rect 40412 32972 40468 32974
rect 40572 33026 40628 33028
rect 40572 32974 40574 33026
rect 40574 32974 40626 33026
rect 40626 32974 40628 33026
rect 40572 32972 40628 32974
rect 40732 33026 40788 33028
rect 40732 32974 40734 33026
rect 40734 32974 40786 33026
rect 40786 32974 40788 33026
rect 40732 32972 40788 32974
rect 40892 33026 40948 33028
rect 40892 32974 40894 33026
rect 40894 32974 40946 33026
rect 40946 32974 40948 33026
rect 40892 32972 40948 32974
rect 41052 33026 41108 33028
rect 41052 32974 41054 33026
rect 41054 32974 41106 33026
rect 41106 32974 41108 33026
rect 41052 32972 41108 32974
rect 41212 33026 41268 33028
rect 41212 32974 41214 33026
rect 41214 32974 41266 33026
rect 41266 32974 41268 33026
rect 41212 32972 41268 32974
rect 41372 33026 41428 33028
rect 41372 32974 41374 33026
rect 41374 32974 41426 33026
rect 41426 32974 41428 33026
rect 41372 32972 41428 32974
rect 41532 33026 41588 33028
rect 41532 32974 41534 33026
rect 41534 32974 41586 33026
rect 41586 32974 41588 33026
rect 41532 32972 41588 32974
rect 41692 33026 41748 33028
rect 41692 32974 41694 33026
rect 41694 32974 41746 33026
rect 41746 32974 41748 33026
rect 41692 32972 41748 32974
rect 41852 33026 41908 33028
rect 41852 32974 41854 33026
rect 41854 32974 41906 33026
rect 41906 32974 41908 33026
rect 41852 32972 41908 32974
rect 12 32866 68 32868
rect 12 32814 14 32866
rect 14 32814 66 32866
rect 66 32814 68 32866
rect 12 32812 68 32814
rect 172 32866 228 32868
rect 172 32814 174 32866
rect 174 32814 226 32866
rect 226 32814 228 32866
rect 172 32812 228 32814
rect 332 32866 388 32868
rect 332 32814 334 32866
rect 334 32814 386 32866
rect 386 32814 388 32866
rect 332 32812 388 32814
rect 492 32866 548 32868
rect 492 32814 494 32866
rect 494 32814 546 32866
rect 546 32814 548 32866
rect 492 32812 548 32814
rect 652 32866 708 32868
rect 652 32814 654 32866
rect 654 32814 706 32866
rect 706 32814 708 32866
rect 652 32812 708 32814
rect 812 32866 868 32868
rect 812 32814 814 32866
rect 814 32814 866 32866
rect 866 32814 868 32866
rect 812 32812 868 32814
rect 972 32866 1028 32868
rect 972 32814 974 32866
rect 974 32814 1026 32866
rect 1026 32814 1028 32866
rect 972 32812 1028 32814
rect 1132 32866 1188 32868
rect 1132 32814 1134 32866
rect 1134 32814 1186 32866
rect 1186 32814 1188 32866
rect 1132 32812 1188 32814
rect 1292 32866 1348 32868
rect 1292 32814 1294 32866
rect 1294 32814 1346 32866
rect 1346 32814 1348 32866
rect 1292 32812 1348 32814
rect 1452 32866 1508 32868
rect 1452 32814 1454 32866
rect 1454 32814 1506 32866
rect 1506 32814 1508 32866
rect 1452 32812 1508 32814
rect 1612 32866 1668 32868
rect 1612 32814 1614 32866
rect 1614 32814 1666 32866
rect 1666 32814 1668 32866
rect 1612 32812 1668 32814
rect 1772 32866 1828 32868
rect 1772 32814 1774 32866
rect 1774 32814 1826 32866
rect 1826 32814 1828 32866
rect 1772 32812 1828 32814
rect 1932 32866 1988 32868
rect 1932 32814 1934 32866
rect 1934 32814 1986 32866
rect 1986 32814 1988 32866
rect 1932 32812 1988 32814
rect 2092 32866 2148 32868
rect 2092 32814 2094 32866
rect 2094 32814 2146 32866
rect 2146 32814 2148 32866
rect 2092 32812 2148 32814
rect 2252 32866 2308 32868
rect 2252 32814 2254 32866
rect 2254 32814 2306 32866
rect 2306 32814 2308 32866
rect 2252 32812 2308 32814
rect 2412 32866 2468 32868
rect 2412 32814 2414 32866
rect 2414 32814 2466 32866
rect 2466 32814 2468 32866
rect 2412 32812 2468 32814
rect 2572 32866 2628 32868
rect 2572 32814 2574 32866
rect 2574 32814 2626 32866
rect 2626 32814 2628 32866
rect 2572 32812 2628 32814
rect 2732 32866 2788 32868
rect 2732 32814 2734 32866
rect 2734 32814 2786 32866
rect 2786 32814 2788 32866
rect 2732 32812 2788 32814
rect 2892 32866 2948 32868
rect 2892 32814 2894 32866
rect 2894 32814 2946 32866
rect 2946 32814 2948 32866
rect 2892 32812 2948 32814
rect 3052 32866 3108 32868
rect 3052 32814 3054 32866
rect 3054 32814 3106 32866
rect 3106 32814 3108 32866
rect 3052 32812 3108 32814
rect 3212 32866 3268 32868
rect 3212 32814 3214 32866
rect 3214 32814 3266 32866
rect 3266 32814 3268 32866
rect 3212 32812 3268 32814
rect 3372 32866 3428 32868
rect 3372 32814 3374 32866
rect 3374 32814 3426 32866
rect 3426 32814 3428 32866
rect 3372 32812 3428 32814
rect 3532 32866 3588 32868
rect 3532 32814 3534 32866
rect 3534 32814 3586 32866
rect 3586 32814 3588 32866
rect 3532 32812 3588 32814
rect 3692 32866 3748 32868
rect 3692 32814 3694 32866
rect 3694 32814 3746 32866
rect 3746 32814 3748 32866
rect 3692 32812 3748 32814
rect 3852 32866 3908 32868
rect 3852 32814 3854 32866
rect 3854 32814 3906 32866
rect 3906 32814 3908 32866
rect 3852 32812 3908 32814
rect 4012 32866 4068 32868
rect 4012 32814 4014 32866
rect 4014 32814 4066 32866
rect 4066 32814 4068 32866
rect 4012 32812 4068 32814
rect 4172 32866 4228 32868
rect 4172 32814 4174 32866
rect 4174 32814 4226 32866
rect 4226 32814 4228 32866
rect 4172 32812 4228 32814
rect 4332 32866 4388 32868
rect 4332 32814 4334 32866
rect 4334 32814 4386 32866
rect 4386 32814 4388 32866
rect 4332 32812 4388 32814
rect 4492 32866 4548 32868
rect 4492 32814 4494 32866
rect 4494 32814 4546 32866
rect 4546 32814 4548 32866
rect 4492 32812 4548 32814
rect 4652 32866 4708 32868
rect 4652 32814 4654 32866
rect 4654 32814 4706 32866
rect 4706 32814 4708 32866
rect 4652 32812 4708 32814
rect 4812 32866 4868 32868
rect 4812 32814 4814 32866
rect 4814 32814 4866 32866
rect 4866 32814 4868 32866
rect 4812 32812 4868 32814
rect 4972 32866 5028 32868
rect 4972 32814 4974 32866
rect 4974 32814 5026 32866
rect 5026 32814 5028 32866
rect 4972 32812 5028 32814
rect 5132 32866 5188 32868
rect 5132 32814 5134 32866
rect 5134 32814 5186 32866
rect 5186 32814 5188 32866
rect 5132 32812 5188 32814
rect 5292 32866 5348 32868
rect 5292 32814 5294 32866
rect 5294 32814 5346 32866
rect 5346 32814 5348 32866
rect 5292 32812 5348 32814
rect 5452 32866 5508 32868
rect 5452 32814 5454 32866
rect 5454 32814 5506 32866
rect 5506 32814 5508 32866
rect 5452 32812 5508 32814
rect 5612 32866 5668 32868
rect 5612 32814 5614 32866
rect 5614 32814 5666 32866
rect 5666 32814 5668 32866
rect 5612 32812 5668 32814
rect 5772 32866 5828 32868
rect 5772 32814 5774 32866
rect 5774 32814 5826 32866
rect 5826 32814 5828 32866
rect 5772 32812 5828 32814
rect 5932 32866 5988 32868
rect 5932 32814 5934 32866
rect 5934 32814 5986 32866
rect 5986 32814 5988 32866
rect 5932 32812 5988 32814
rect 6092 32866 6148 32868
rect 6092 32814 6094 32866
rect 6094 32814 6146 32866
rect 6146 32814 6148 32866
rect 6092 32812 6148 32814
rect 6252 32866 6308 32868
rect 6252 32814 6254 32866
rect 6254 32814 6306 32866
rect 6306 32814 6308 32866
rect 6252 32812 6308 32814
rect 6412 32866 6468 32868
rect 6412 32814 6414 32866
rect 6414 32814 6466 32866
rect 6466 32814 6468 32866
rect 6412 32812 6468 32814
rect 6572 32866 6628 32868
rect 6572 32814 6574 32866
rect 6574 32814 6626 32866
rect 6626 32814 6628 32866
rect 6572 32812 6628 32814
rect 6732 32866 6788 32868
rect 6732 32814 6734 32866
rect 6734 32814 6786 32866
rect 6786 32814 6788 32866
rect 6732 32812 6788 32814
rect 6892 32866 6948 32868
rect 6892 32814 6894 32866
rect 6894 32814 6946 32866
rect 6946 32814 6948 32866
rect 6892 32812 6948 32814
rect 7052 32866 7108 32868
rect 7052 32814 7054 32866
rect 7054 32814 7106 32866
rect 7106 32814 7108 32866
rect 7052 32812 7108 32814
rect 7212 32866 7268 32868
rect 7212 32814 7214 32866
rect 7214 32814 7266 32866
rect 7266 32814 7268 32866
rect 7212 32812 7268 32814
rect 7372 32866 7428 32868
rect 7372 32814 7374 32866
rect 7374 32814 7426 32866
rect 7426 32814 7428 32866
rect 7372 32812 7428 32814
rect 7532 32866 7588 32868
rect 7532 32814 7534 32866
rect 7534 32814 7586 32866
rect 7586 32814 7588 32866
rect 7532 32812 7588 32814
rect 7692 32866 7748 32868
rect 7692 32814 7694 32866
rect 7694 32814 7746 32866
rect 7746 32814 7748 32866
rect 7692 32812 7748 32814
rect 7852 32866 7908 32868
rect 7852 32814 7854 32866
rect 7854 32814 7906 32866
rect 7906 32814 7908 32866
rect 7852 32812 7908 32814
rect 8012 32866 8068 32868
rect 8012 32814 8014 32866
rect 8014 32814 8066 32866
rect 8066 32814 8068 32866
rect 8012 32812 8068 32814
rect 8172 32866 8228 32868
rect 8172 32814 8174 32866
rect 8174 32814 8226 32866
rect 8226 32814 8228 32866
rect 8172 32812 8228 32814
rect 8332 32866 8388 32868
rect 8332 32814 8334 32866
rect 8334 32814 8386 32866
rect 8386 32814 8388 32866
rect 8332 32812 8388 32814
rect 8972 32812 9028 32868
rect 9292 32812 9348 32868
rect 12492 32866 12548 32868
rect 12492 32814 12494 32866
rect 12494 32814 12546 32866
rect 12546 32814 12548 32866
rect 12492 32812 12548 32814
rect 12652 32866 12708 32868
rect 12652 32814 12654 32866
rect 12654 32814 12706 32866
rect 12706 32814 12708 32866
rect 12652 32812 12708 32814
rect 12812 32866 12868 32868
rect 12812 32814 12814 32866
rect 12814 32814 12866 32866
rect 12866 32814 12868 32866
rect 12812 32812 12868 32814
rect 12972 32866 13028 32868
rect 12972 32814 12974 32866
rect 12974 32814 13026 32866
rect 13026 32814 13028 32866
rect 12972 32812 13028 32814
rect 13132 32866 13188 32868
rect 13132 32814 13134 32866
rect 13134 32814 13186 32866
rect 13186 32814 13188 32866
rect 13132 32812 13188 32814
rect 13292 32866 13348 32868
rect 13292 32814 13294 32866
rect 13294 32814 13346 32866
rect 13346 32814 13348 32866
rect 13292 32812 13348 32814
rect 13452 32866 13508 32868
rect 13452 32814 13454 32866
rect 13454 32814 13506 32866
rect 13506 32814 13508 32866
rect 13452 32812 13508 32814
rect 13612 32866 13668 32868
rect 13612 32814 13614 32866
rect 13614 32814 13666 32866
rect 13666 32814 13668 32866
rect 13612 32812 13668 32814
rect 13772 32866 13828 32868
rect 13772 32814 13774 32866
rect 13774 32814 13826 32866
rect 13826 32814 13828 32866
rect 13772 32812 13828 32814
rect 13932 32866 13988 32868
rect 13932 32814 13934 32866
rect 13934 32814 13986 32866
rect 13986 32814 13988 32866
rect 13932 32812 13988 32814
rect 14092 32866 14148 32868
rect 14092 32814 14094 32866
rect 14094 32814 14146 32866
rect 14146 32814 14148 32866
rect 14092 32812 14148 32814
rect 14252 32866 14308 32868
rect 14252 32814 14254 32866
rect 14254 32814 14306 32866
rect 14306 32814 14308 32866
rect 14252 32812 14308 32814
rect 14412 32866 14468 32868
rect 14412 32814 14414 32866
rect 14414 32814 14466 32866
rect 14466 32814 14468 32866
rect 14412 32812 14468 32814
rect 14572 32866 14628 32868
rect 14572 32814 14574 32866
rect 14574 32814 14626 32866
rect 14626 32814 14628 32866
rect 14572 32812 14628 32814
rect 14732 32866 14788 32868
rect 14732 32814 14734 32866
rect 14734 32814 14786 32866
rect 14786 32814 14788 32866
rect 14732 32812 14788 32814
rect 14892 32866 14948 32868
rect 14892 32814 14894 32866
rect 14894 32814 14946 32866
rect 14946 32814 14948 32866
rect 14892 32812 14948 32814
rect 15052 32866 15108 32868
rect 15052 32814 15054 32866
rect 15054 32814 15106 32866
rect 15106 32814 15108 32866
rect 15052 32812 15108 32814
rect 15212 32866 15268 32868
rect 15212 32814 15214 32866
rect 15214 32814 15266 32866
rect 15266 32814 15268 32866
rect 15212 32812 15268 32814
rect 15372 32866 15428 32868
rect 15372 32814 15374 32866
rect 15374 32814 15426 32866
rect 15426 32814 15428 32866
rect 15372 32812 15428 32814
rect 15532 32866 15588 32868
rect 15532 32814 15534 32866
rect 15534 32814 15586 32866
rect 15586 32814 15588 32866
rect 15532 32812 15588 32814
rect 15692 32866 15748 32868
rect 15692 32814 15694 32866
rect 15694 32814 15746 32866
rect 15746 32814 15748 32866
rect 15692 32812 15748 32814
rect 15852 32866 15908 32868
rect 15852 32814 15854 32866
rect 15854 32814 15906 32866
rect 15906 32814 15908 32866
rect 15852 32812 15908 32814
rect 16012 32866 16068 32868
rect 16012 32814 16014 32866
rect 16014 32814 16066 32866
rect 16066 32814 16068 32866
rect 16012 32812 16068 32814
rect 16172 32866 16228 32868
rect 16172 32814 16174 32866
rect 16174 32814 16226 32866
rect 16226 32814 16228 32866
rect 16172 32812 16228 32814
rect 16332 32866 16388 32868
rect 16332 32814 16334 32866
rect 16334 32814 16386 32866
rect 16386 32814 16388 32866
rect 16332 32812 16388 32814
rect 16492 32866 16548 32868
rect 16492 32814 16494 32866
rect 16494 32814 16546 32866
rect 16546 32814 16548 32866
rect 16492 32812 16548 32814
rect 16652 32866 16708 32868
rect 16652 32814 16654 32866
rect 16654 32814 16706 32866
rect 16706 32814 16708 32866
rect 16652 32812 16708 32814
rect 16812 32866 16868 32868
rect 16812 32814 16814 32866
rect 16814 32814 16866 32866
rect 16866 32814 16868 32866
rect 16812 32812 16868 32814
rect 16972 32866 17028 32868
rect 16972 32814 16974 32866
rect 16974 32814 17026 32866
rect 17026 32814 17028 32866
rect 16972 32812 17028 32814
rect 17132 32866 17188 32868
rect 17132 32814 17134 32866
rect 17134 32814 17186 32866
rect 17186 32814 17188 32866
rect 17132 32812 17188 32814
rect 17292 32866 17348 32868
rect 17292 32814 17294 32866
rect 17294 32814 17346 32866
rect 17346 32814 17348 32866
rect 17292 32812 17348 32814
rect 17452 32866 17508 32868
rect 17452 32814 17454 32866
rect 17454 32814 17506 32866
rect 17506 32814 17508 32866
rect 17452 32812 17508 32814
rect 17612 32866 17668 32868
rect 17612 32814 17614 32866
rect 17614 32814 17666 32866
rect 17666 32814 17668 32866
rect 17612 32812 17668 32814
rect 17772 32866 17828 32868
rect 17772 32814 17774 32866
rect 17774 32814 17826 32866
rect 17826 32814 17828 32866
rect 17772 32812 17828 32814
rect 17932 32866 17988 32868
rect 17932 32814 17934 32866
rect 17934 32814 17986 32866
rect 17986 32814 17988 32866
rect 17932 32812 17988 32814
rect 18092 32866 18148 32868
rect 18092 32814 18094 32866
rect 18094 32814 18146 32866
rect 18146 32814 18148 32866
rect 18092 32812 18148 32814
rect 18252 32866 18308 32868
rect 18252 32814 18254 32866
rect 18254 32814 18306 32866
rect 18306 32814 18308 32866
rect 18252 32812 18308 32814
rect 18412 32866 18468 32868
rect 18412 32814 18414 32866
rect 18414 32814 18466 32866
rect 18466 32814 18468 32866
rect 18412 32812 18468 32814
rect 18572 32866 18628 32868
rect 18572 32814 18574 32866
rect 18574 32814 18626 32866
rect 18626 32814 18628 32866
rect 18572 32812 18628 32814
rect 18732 32866 18788 32868
rect 18732 32814 18734 32866
rect 18734 32814 18786 32866
rect 18786 32814 18788 32866
rect 18732 32812 18788 32814
rect 18892 32866 18948 32868
rect 18892 32814 18894 32866
rect 18894 32814 18946 32866
rect 18946 32814 18948 32866
rect 18892 32812 18948 32814
rect 19532 32812 19588 32868
rect 19852 32812 19908 32868
rect 23132 32866 23188 32868
rect 23132 32814 23134 32866
rect 23134 32814 23186 32866
rect 23186 32814 23188 32866
rect 23132 32812 23188 32814
rect 23292 32866 23348 32868
rect 23292 32814 23294 32866
rect 23294 32814 23346 32866
rect 23346 32814 23348 32866
rect 23292 32812 23348 32814
rect 23452 32866 23508 32868
rect 23452 32814 23454 32866
rect 23454 32814 23506 32866
rect 23506 32814 23508 32866
rect 23452 32812 23508 32814
rect 23612 32866 23668 32868
rect 23612 32814 23614 32866
rect 23614 32814 23666 32866
rect 23666 32814 23668 32866
rect 23612 32812 23668 32814
rect 23772 32866 23828 32868
rect 23772 32814 23774 32866
rect 23774 32814 23826 32866
rect 23826 32814 23828 32866
rect 23772 32812 23828 32814
rect 23932 32866 23988 32868
rect 23932 32814 23934 32866
rect 23934 32814 23986 32866
rect 23986 32814 23988 32866
rect 23932 32812 23988 32814
rect 24092 32866 24148 32868
rect 24092 32814 24094 32866
rect 24094 32814 24146 32866
rect 24146 32814 24148 32866
rect 24092 32812 24148 32814
rect 24252 32866 24308 32868
rect 24252 32814 24254 32866
rect 24254 32814 24306 32866
rect 24306 32814 24308 32866
rect 24252 32812 24308 32814
rect 24412 32866 24468 32868
rect 24412 32814 24414 32866
rect 24414 32814 24466 32866
rect 24466 32814 24468 32866
rect 24412 32812 24468 32814
rect 24572 32866 24628 32868
rect 24572 32814 24574 32866
rect 24574 32814 24626 32866
rect 24626 32814 24628 32866
rect 24572 32812 24628 32814
rect 24732 32866 24788 32868
rect 24732 32814 24734 32866
rect 24734 32814 24786 32866
rect 24786 32814 24788 32866
rect 24732 32812 24788 32814
rect 24892 32866 24948 32868
rect 24892 32814 24894 32866
rect 24894 32814 24946 32866
rect 24946 32814 24948 32866
rect 24892 32812 24948 32814
rect 25052 32866 25108 32868
rect 25052 32814 25054 32866
rect 25054 32814 25106 32866
rect 25106 32814 25108 32866
rect 25052 32812 25108 32814
rect 25212 32866 25268 32868
rect 25212 32814 25214 32866
rect 25214 32814 25266 32866
rect 25266 32814 25268 32866
rect 25212 32812 25268 32814
rect 25372 32866 25428 32868
rect 25372 32814 25374 32866
rect 25374 32814 25426 32866
rect 25426 32814 25428 32866
rect 25372 32812 25428 32814
rect 25532 32866 25588 32868
rect 25532 32814 25534 32866
rect 25534 32814 25586 32866
rect 25586 32814 25588 32866
rect 25532 32812 25588 32814
rect 25692 32866 25748 32868
rect 25692 32814 25694 32866
rect 25694 32814 25746 32866
rect 25746 32814 25748 32866
rect 25692 32812 25748 32814
rect 25852 32866 25908 32868
rect 25852 32814 25854 32866
rect 25854 32814 25906 32866
rect 25906 32814 25908 32866
rect 25852 32812 25908 32814
rect 26012 32866 26068 32868
rect 26012 32814 26014 32866
rect 26014 32814 26066 32866
rect 26066 32814 26068 32866
rect 26012 32812 26068 32814
rect 26172 32866 26228 32868
rect 26172 32814 26174 32866
rect 26174 32814 26226 32866
rect 26226 32814 26228 32866
rect 26172 32812 26228 32814
rect 26332 32866 26388 32868
rect 26332 32814 26334 32866
rect 26334 32814 26386 32866
rect 26386 32814 26388 32866
rect 26332 32812 26388 32814
rect 26492 32866 26548 32868
rect 26492 32814 26494 32866
rect 26494 32814 26546 32866
rect 26546 32814 26548 32866
rect 26492 32812 26548 32814
rect 26652 32866 26708 32868
rect 26652 32814 26654 32866
rect 26654 32814 26706 32866
rect 26706 32814 26708 32866
rect 26652 32812 26708 32814
rect 26812 32866 26868 32868
rect 26812 32814 26814 32866
rect 26814 32814 26866 32866
rect 26866 32814 26868 32866
rect 26812 32812 26868 32814
rect 26972 32866 27028 32868
rect 26972 32814 26974 32866
rect 26974 32814 27026 32866
rect 27026 32814 27028 32866
rect 26972 32812 27028 32814
rect 27132 32866 27188 32868
rect 27132 32814 27134 32866
rect 27134 32814 27186 32866
rect 27186 32814 27188 32866
rect 27132 32812 27188 32814
rect 27292 32866 27348 32868
rect 27292 32814 27294 32866
rect 27294 32814 27346 32866
rect 27346 32814 27348 32866
rect 27292 32812 27348 32814
rect 27452 32866 27508 32868
rect 27452 32814 27454 32866
rect 27454 32814 27506 32866
rect 27506 32814 27508 32866
rect 27452 32812 27508 32814
rect 27612 32866 27668 32868
rect 27612 32814 27614 32866
rect 27614 32814 27666 32866
rect 27666 32814 27668 32866
rect 27612 32812 27668 32814
rect 27772 32866 27828 32868
rect 27772 32814 27774 32866
rect 27774 32814 27826 32866
rect 27826 32814 27828 32866
rect 27772 32812 27828 32814
rect 27932 32866 27988 32868
rect 27932 32814 27934 32866
rect 27934 32814 27986 32866
rect 27986 32814 27988 32866
rect 27932 32812 27988 32814
rect 28092 32866 28148 32868
rect 28092 32814 28094 32866
rect 28094 32814 28146 32866
rect 28146 32814 28148 32866
rect 28092 32812 28148 32814
rect 28252 32866 28308 32868
rect 28252 32814 28254 32866
rect 28254 32814 28306 32866
rect 28306 32814 28308 32866
rect 28252 32812 28308 32814
rect 28412 32866 28468 32868
rect 28412 32814 28414 32866
rect 28414 32814 28466 32866
rect 28466 32814 28468 32866
rect 28412 32812 28468 32814
rect 28572 32866 28628 32868
rect 28572 32814 28574 32866
rect 28574 32814 28626 32866
rect 28626 32814 28628 32866
rect 28572 32812 28628 32814
rect 28732 32866 28788 32868
rect 28732 32814 28734 32866
rect 28734 32814 28786 32866
rect 28786 32814 28788 32866
rect 28732 32812 28788 32814
rect 28892 32866 28948 32868
rect 28892 32814 28894 32866
rect 28894 32814 28946 32866
rect 28946 32814 28948 32866
rect 28892 32812 28948 32814
rect 29052 32866 29108 32868
rect 29052 32814 29054 32866
rect 29054 32814 29106 32866
rect 29106 32814 29108 32866
rect 29052 32812 29108 32814
rect 29212 32866 29268 32868
rect 29212 32814 29214 32866
rect 29214 32814 29266 32866
rect 29266 32814 29268 32866
rect 29212 32812 29268 32814
rect 29372 32866 29428 32868
rect 29372 32814 29374 32866
rect 29374 32814 29426 32866
rect 29426 32814 29428 32866
rect 29372 32812 29428 32814
rect 32572 32812 32628 32868
rect 32892 32812 32948 32868
rect 33532 32866 33588 32868
rect 33532 32814 33534 32866
rect 33534 32814 33586 32866
rect 33586 32814 33588 32866
rect 33532 32812 33588 32814
rect 33692 32866 33748 32868
rect 33692 32814 33694 32866
rect 33694 32814 33746 32866
rect 33746 32814 33748 32866
rect 33692 32812 33748 32814
rect 33852 32866 33908 32868
rect 33852 32814 33854 32866
rect 33854 32814 33906 32866
rect 33906 32814 33908 32866
rect 33852 32812 33908 32814
rect 34012 32866 34068 32868
rect 34012 32814 34014 32866
rect 34014 32814 34066 32866
rect 34066 32814 34068 32866
rect 34012 32812 34068 32814
rect 34172 32866 34228 32868
rect 34172 32814 34174 32866
rect 34174 32814 34226 32866
rect 34226 32814 34228 32866
rect 34172 32812 34228 32814
rect 34332 32866 34388 32868
rect 34332 32814 34334 32866
rect 34334 32814 34386 32866
rect 34386 32814 34388 32866
rect 34332 32812 34388 32814
rect 34492 32866 34548 32868
rect 34492 32814 34494 32866
rect 34494 32814 34546 32866
rect 34546 32814 34548 32866
rect 34492 32812 34548 32814
rect 34652 32866 34708 32868
rect 34652 32814 34654 32866
rect 34654 32814 34706 32866
rect 34706 32814 34708 32866
rect 34652 32812 34708 32814
rect 34812 32866 34868 32868
rect 34812 32814 34814 32866
rect 34814 32814 34866 32866
rect 34866 32814 34868 32866
rect 34812 32812 34868 32814
rect 34972 32866 35028 32868
rect 34972 32814 34974 32866
rect 34974 32814 35026 32866
rect 35026 32814 35028 32866
rect 34972 32812 35028 32814
rect 35132 32866 35188 32868
rect 35132 32814 35134 32866
rect 35134 32814 35186 32866
rect 35186 32814 35188 32866
rect 35132 32812 35188 32814
rect 35292 32866 35348 32868
rect 35292 32814 35294 32866
rect 35294 32814 35346 32866
rect 35346 32814 35348 32866
rect 35292 32812 35348 32814
rect 35452 32866 35508 32868
rect 35452 32814 35454 32866
rect 35454 32814 35506 32866
rect 35506 32814 35508 32866
rect 35452 32812 35508 32814
rect 35612 32866 35668 32868
rect 35612 32814 35614 32866
rect 35614 32814 35666 32866
rect 35666 32814 35668 32866
rect 35612 32812 35668 32814
rect 35772 32866 35828 32868
rect 35772 32814 35774 32866
rect 35774 32814 35826 32866
rect 35826 32814 35828 32866
rect 35772 32812 35828 32814
rect 35932 32866 35988 32868
rect 35932 32814 35934 32866
rect 35934 32814 35986 32866
rect 35986 32814 35988 32866
rect 35932 32812 35988 32814
rect 36092 32866 36148 32868
rect 36092 32814 36094 32866
rect 36094 32814 36146 32866
rect 36146 32814 36148 32866
rect 36092 32812 36148 32814
rect 36252 32866 36308 32868
rect 36252 32814 36254 32866
rect 36254 32814 36306 32866
rect 36306 32814 36308 32866
rect 36252 32812 36308 32814
rect 36412 32866 36468 32868
rect 36412 32814 36414 32866
rect 36414 32814 36466 32866
rect 36466 32814 36468 32866
rect 36412 32812 36468 32814
rect 36572 32866 36628 32868
rect 36572 32814 36574 32866
rect 36574 32814 36626 32866
rect 36626 32814 36628 32866
rect 36572 32812 36628 32814
rect 36732 32866 36788 32868
rect 36732 32814 36734 32866
rect 36734 32814 36786 32866
rect 36786 32814 36788 32866
rect 36732 32812 36788 32814
rect 36892 32866 36948 32868
rect 36892 32814 36894 32866
rect 36894 32814 36946 32866
rect 36946 32814 36948 32866
rect 36892 32812 36948 32814
rect 37052 32866 37108 32868
rect 37052 32814 37054 32866
rect 37054 32814 37106 32866
rect 37106 32814 37108 32866
rect 37052 32812 37108 32814
rect 37212 32866 37268 32868
rect 37212 32814 37214 32866
rect 37214 32814 37266 32866
rect 37266 32814 37268 32866
rect 37212 32812 37268 32814
rect 37372 32866 37428 32868
rect 37372 32814 37374 32866
rect 37374 32814 37426 32866
rect 37426 32814 37428 32866
rect 37372 32812 37428 32814
rect 37532 32866 37588 32868
rect 37532 32814 37534 32866
rect 37534 32814 37586 32866
rect 37586 32814 37588 32866
rect 37532 32812 37588 32814
rect 37692 32866 37748 32868
rect 37692 32814 37694 32866
rect 37694 32814 37746 32866
rect 37746 32814 37748 32866
rect 37692 32812 37748 32814
rect 37852 32866 37908 32868
rect 37852 32814 37854 32866
rect 37854 32814 37906 32866
rect 37906 32814 37908 32866
rect 37852 32812 37908 32814
rect 38012 32866 38068 32868
rect 38012 32814 38014 32866
rect 38014 32814 38066 32866
rect 38066 32814 38068 32866
rect 38012 32812 38068 32814
rect 38172 32866 38228 32868
rect 38172 32814 38174 32866
rect 38174 32814 38226 32866
rect 38226 32814 38228 32866
rect 38172 32812 38228 32814
rect 38332 32866 38388 32868
rect 38332 32814 38334 32866
rect 38334 32814 38386 32866
rect 38386 32814 38388 32866
rect 38332 32812 38388 32814
rect 38492 32866 38548 32868
rect 38492 32814 38494 32866
rect 38494 32814 38546 32866
rect 38546 32814 38548 32866
rect 38492 32812 38548 32814
rect 38652 32866 38708 32868
rect 38652 32814 38654 32866
rect 38654 32814 38706 32866
rect 38706 32814 38708 32866
rect 38652 32812 38708 32814
rect 38812 32866 38868 32868
rect 38812 32814 38814 32866
rect 38814 32814 38866 32866
rect 38866 32814 38868 32866
rect 38812 32812 38868 32814
rect 38972 32866 39028 32868
rect 38972 32814 38974 32866
rect 38974 32814 39026 32866
rect 39026 32814 39028 32866
rect 38972 32812 39028 32814
rect 39132 32866 39188 32868
rect 39132 32814 39134 32866
rect 39134 32814 39186 32866
rect 39186 32814 39188 32866
rect 39132 32812 39188 32814
rect 39292 32866 39348 32868
rect 39292 32814 39294 32866
rect 39294 32814 39346 32866
rect 39346 32814 39348 32866
rect 39292 32812 39348 32814
rect 39452 32866 39508 32868
rect 39452 32814 39454 32866
rect 39454 32814 39506 32866
rect 39506 32814 39508 32866
rect 39452 32812 39508 32814
rect 39612 32866 39668 32868
rect 39612 32814 39614 32866
rect 39614 32814 39666 32866
rect 39666 32814 39668 32866
rect 39612 32812 39668 32814
rect 39772 32866 39828 32868
rect 39772 32814 39774 32866
rect 39774 32814 39826 32866
rect 39826 32814 39828 32866
rect 39772 32812 39828 32814
rect 39932 32866 39988 32868
rect 39932 32814 39934 32866
rect 39934 32814 39986 32866
rect 39986 32814 39988 32866
rect 39932 32812 39988 32814
rect 40092 32866 40148 32868
rect 40092 32814 40094 32866
rect 40094 32814 40146 32866
rect 40146 32814 40148 32866
rect 40092 32812 40148 32814
rect 40252 32866 40308 32868
rect 40252 32814 40254 32866
rect 40254 32814 40306 32866
rect 40306 32814 40308 32866
rect 40252 32812 40308 32814
rect 40412 32866 40468 32868
rect 40412 32814 40414 32866
rect 40414 32814 40466 32866
rect 40466 32814 40468 32866
rect 40412 32812 40468 32814
rect 40572 32866 40628 32868
rect 40572 32814 40574 32866
rect 40574 32814 40626 32866
rect 40626 32814 40628 32866
rect 40572 32812 40628 32814
rect 40732 32866 40788 32868
rect 40732 32814 40734 32866
rect 40734 32814 40786 32866
rect 40786 32814 40788 32866
rect 40732 32812 40788 32814
rect 40892 32866 40948 32868
rect 40892 32814 40894 32866
rect 40894 32814 40946 32866
rect 40946 32814 40948 32866
rect 40892 32812 40948 32814
rect 41052 32866 41108 32868
rect 41052 32814 41054 32866
rect 41054 32814 41106 32866
rect 41106 32814 41108 32866
rect 41052 32812 41108 32814
rect 41212 32866 41268 32868
rect 41212 32814 41214 32866
rect 41214 32814 41266 32866
rect 41266 32814 41268 32866
rect 41212 32812 41268 32814
rect 41372 32866 41428 32868
rect 41372 32814 41374 32866
rect 41374 32814 41426 32866
rect 41426 32814 41428 32866
rect 41372 32812 41428 32814
rect 41532 32866 41588 32868
rect 41532 32814 41534 32866
rect 41534 32814 41586 32866
rect 41586 32814 41588 32866
rect 41532 32812 41588 32814
rect 41692 32866 41748 32868
rect 41692 32814 41694 32866
rect 41694 32814 41746 32866
rect 41746 32814 41748 32866
rect 41692 32812 41748 32814
rect 41852 32866 41908 32868
rect 41852 32814 41854 32866
rect 41854 32814 41906 32866
rect 41906 32814 41908 32866
rect 41852 32812 41908 32814
rect 9132 32652 9188 32708
rect 19692 32652 19748 32708
rect 32732 32652 32788 32708
rect 12 32546 68 32548
rect 12 32494 14 32546
rect 14 32494 66 32546
rect 66 32494 68 32546
rect 12 32492 68 32494
rect 172 32546 228 32548
rect 172 32494 174 32546
rect 174 32494 226 32546
rect 226 32494 228 32546
rect 172 32492 228 32494
rect 332 32546 388 32548
rect 332 32494 334 32546
rect 334 32494 386 32546
rect 386 32494 388 32546
rect 332 32492 388 32494
rect 492 32546 548 32548
rect 492 32494 494 32546
rect 494 32494 546 32546
rect 546 32494 548 32546
rect 492 32492 548 32494
rect 652 32546 708 32548
rect 652 32494 654 32546
rect 654 32494 706 32546
rect 706 32494 708 32546
rect 652 32492 708 32494
rect 812 32546 868 32548
rect 812 32494 814 32546
rect 814 32494 866 32546
rect 866 32494 868 32546
rect 812 32492 868 32494
rect 972 32546 1028 32548
rect 972 32494 974 32546
rect 974 32494 1026 32546
rect 1026 32494 1028 32546
rect 972 32492 1028 32494
rect 1132 32546 1188 32548
rect 1132 32494 1134 32546
rect 1134 32494 1186 32546
rect 1186 32494 1188 32546
rect 1132 32492 1188 32494
rect 1292 32546 1348 32548
rect 1292 32494 1294 32546
rect 1294 32494 1346 32546
rect 1346 32494 1348 32546
rect 1292 32492 1348 32494
rect 1452 32546 1508 32548
rect 1452 32494 1454 32546
rect 1454 32494 1506 32546
rect 1506 32494 1508 32546
rect 1452 32492 1508 32494
rect 1612 32546 1668 32548
rect 1612 32494 1614 32546
rect 1614 32494 1666 32546
rect 1666 32494 1668 32546
rect 1612 32492 1668 32494
rect 1772 32546 1828 32548
rect 1772 32494 1774 32546
rect 1774 32494 1826 32546
rect 1826 32494 1828 32546
rect 1772 32492 1828 32494
rect 1932 32546 1988 32548
rect 1932 32494 1934 32546
rect 1934 32494 1986 32546
rect 1986 32494 1988 32546
rect 1932 32492 1988 32494
rect 2092 32546 2148 32548
rect 2092 32494 2094 32546
rect 2094 32494 2146 32546
rect 2146 32494 2148 32546
rect 2092 32492 2148 32494
rect 2252 32546 2308 32548
rect 2252 32494 2254 32546
rect 2254 32494 2306 32546
rect 2306 32494 2308 32546
rect 2252 32492 2308 32494
rect 2412 32546 2468 32548
rect 2412 32494 2414 32546
rect 2414 32494 2466 32546
rect 2466 32494 2468 32546
rect 2412 32492 2468 32494
rect 2572 32546 2628 32548
rect 2572 32494 2574 32546
rect 2574 32494 2626 32546
rect 2626 32494 2628 32546
rect 2572 32492 2628 32494
rect 2732 32546 2788 32548
rect 2732 32494 2734 32546
rect 2734 32494 2786 32546
rect 2786 32494 2788 32546
rect 2732 32492 2788 32494
rect 2892 32546 2948 32548
rect 2892 32494 2894 32546
rect 2894 32494 2946 32546
rect 2946 32494 2948 32546
rect 2892 32492 2948 32494
rect 3052 32546 3108 32548
rect 3052 32494 3054 32546
rect 3054 32494 3106 32546
rect 3106 32494 3108 32546
rect 3052 32492 3108 32494
rect 3212 32546 3268 32548
rect 3212 32494 3214 32546
rect 3214 32494 3266 32546
rect 3266 32494 3268 32546
rect 3212 32492 3268 32494
rect 3372 32546 3428 32548
rect 3372 32494 3374 32546
rect 3374 32494 3426 32546
rect 3426 32494 3428 32546
rect 3372 32492 3428 32494
rect 3532 32546 3588 32548
rect 3532 32494 3534 32546
rect 3534 32494 3586 32546
rect 3586 32494 3588 32546
rect 3532 32492 3588 32494
rect 3692 32546 3748 32548
rect 3692 32494 3694 32546
rect 3694 32494 3746 32546
rect 3746 32494 3748 32546
rect 3692 32492 3748 32494
rect 3852 32546 3908 32548
rect 3852 32494 3854 32546
rect 3854 32494 3906 32546
rect 3906 32494 3908 32546
rect 3852 32492 3908 32494
rect 4012 32546 4068 32548
rect 4012 32494 4014 32546
rect 4014 32494 4066 32546
rect 4066 32494 4068 32546
rect 4012 32492 4068 32494
rect 4172 32546 4228 32548
rect 4172 32494 4174 32546
rect 4174 32494 4226 32546
rect 4226 32494 4228 32546
rect 4172 32492 4228 32494
rect 4332 32546 4388 32548
rect 4332 32494 4334 32546
rect 4334 32494 4386 32546
rect 4386 32494 4388 32546
rect 4332 32492 4388 32494
rect 4492 32546 4548 32548
rect 4492 32494 4494 32546
rect 4494 32494 4546 32546
rect 4546 32494 4548 32546
rect 4492 32492 4548 32494
rect 4652 32546 4708 32548
rect 4652 32494 4654 32546
rect 4654 32494 4706 32546
rect 4706 32494 4708 32546
rect 4652 32492 4708 32494
rect 4812 32546 4868 32548
rect 4812 32494 4814 32546
rect 4814 32494 4866 32546
rect 4866 32494 4868 32546
rect 4812 32492 4868 32494
rect 4972 32546 5028 32548
rect 4972 32494 4974 32546
rect 4974 32494 5026 32546
rect 5026 32494 5028 32546
rect 4972 32492 5028 32494
rect 5132 32546 5188 32548
rect 5132 32494 5134 32546
rect 5134 32494 5186 32546
rect 5186 32494 5188 32546
rect 5132 32492 5188 32494
rect 5292 32546 5348 32548
rect 5292 32494 5294 32546
rect 5294 32494 5346 32546
rect 5346 32494 5348 32546
rect 5292 32492 5348 32494
rect 5452 32546 5508 32548
rect 5452 32494 5454 32546
rect 5454 32494 5506 32546
rect 5506 32494 5508 32546
rect 5452 32492 5508 32494
rect 5612 32546 5668 32548
rect 5612 32494 5614 32546
rect 5614 32494 5666 32546
rect 5666 32494 5668 32546
rect 5612 32492 5668 32494
rect 5772 32546 5828 32548
rect 5772 32494 5774 32546
rect 5774 32494 5826 32546
rect 5826 32494 5828 32546
rect 5772 32492 5828 32494
rect 5932 32546 5988 32548
rect 5932 32494 5934 32546
rect 5934 32494 5986 32546
rect 5986 32494 5988 32546
rect 5932 32492 5988 32494
rect 6092 32546 6148 32548
rect 6092 32494 6094 32546
rect 6094 32494 6146 32546
rect 6146 32494 6148 32546
rect 6092 32492 6148 32494
rect 6252 32546 6308 32548
rect 6252 32494 6254 32546
rect 6254 32494 6306 32546
rect 6306 32494 6308 32546
rect 6252 32492 6308 32494
rect 6412 32546 6468 32548
rect 6412 32494 6414 32546
rect 6414 32494 6466 32546
rect 6466 32494 6468 32546
rect 6412 32492 6468 32494
rect 6572 32546 6628 32548
rect 6572 32494 6574 32546
rect 6574 32494 6626 32546
rect 6626 32494 6628 32546
rect 6572 32492 6628 32494
rect 6732 32546 6788 32548
rect 6732 32494 6734 32546
rect 6734 32494 6786 32546
rect 6786 32494 6788 32546
rect 6732 32492 6788 32494
rect 6892 32546 6948 32548
rect 6892 32494 6894 32546
rect 6894 32494 6946 32546
rect 6946 32494 6948 32546
rect 6892 32492 6948 32494
rect 7052 32546 7108 32548
rect 7052 32494 7054 32546
rect 7054 32494 7106 32546
rect 7106 32494 7108 32546
rect 7052 32492 7108 32494
rect 7212 32546 7268 32548
rect 7212 32494 7214 32546
rect 7214 32494 7266 32546
rect 7266 32494 7268 32546
rect 7212 32492 7268 32494
rect 7372 32546 7428 32548
rect 7372 32494 7374 32546
rect 7374 32494 7426 32546
rect 7426 32494 7428 32546
rect 7372 32492 7428 32494
rect 7532 32546 7588 32548
rect 7532 32494 7534 32546
rect 7534 32494 7586 32546
rect 7586 32494 7588 32546
rect 7532 32492 7588 32494
rect 7692 32546 7748 32548
rect 7692 32494 7694 32546
rect 7694 32494 7746 32546
rect 7746 32494 7748 32546
rect 7692 32492 7748 32494
rect 7852 32546 7908 32548
rect 7852 32494 7854 32546
rect 7854 32494 7906 32546
rect 7906 32494 7908 32546
rect 7852 32492 7908 32494
rect 8012 32546 8068 32548
rect 8012 32494 8014 32546
rect 8014 32494 8066 32546
rect 8066 32494 8068 32546
rect 8012 32492 8068 32494
rect 8172 32546 8228 32548
rect 8172 32494 8174 32546
rect 8174 32494 8226 32546
rect 8226 32494 8228 32546
rect 8172 32492 8228 32494
rect 8332 32546 8388 32548
rect 8332 32494 8334 32546
rect 8334 32494 8386 32546
rect 8386 32494 8388 32546
rect 8332 32492 8388 32494
rect 8972 32492 9028 32548
rect 9292 32492 9348 32548
rect 12492 32546 12548 32548
rect 12492 32494 12494 32546
rect 12494 32494 12546 32546
rect 12546 32494 12548 32546
rect 12492 32492 12548 32494
rect 12652 32546 12708 32548
rect 12652 32494 12654 32546
rect 12654 32494 12706 32546
rect 12706 32494 12708 32546
rect 12652 32492 12708 32494
rect 12812 32546 12868 32548
rect 12812 32494 12814 32546
rect 12814 32494 12866 32546
rect 12866 32494 12868 32546
rect 12812 32492 12868 32494
rect 12972 32546 13028 32548
rect 12972 32494 12974 32546
rect 12974 32494 13026 32546
rect 13026 32494 13028 32546
rect 12972 32492 13028 32494
rect 13132 32546 13188 32548
rect 13132 32494 13134 32546
rect 13134 32494 13186 32546
rect 13186 32494 13188 32546
rect 13132 32492 13188 32494
rect 13292 32546 13348 32548
rect 13292 32494 13294 32546
rect 13294 32494 13346 32546
rect 13346 32494 13348 32546
rect 13292 32492 13348 32494
rect 13452 32546 13508 32548
rect 13452 32494 13454 32546
rect 13454 32494 13506 32546
rect 13506 32494 13508 32546
rect 13452 32492 13508 32494
rect 13612 32546 13668 32548
rect 13612 32494 13614 32546
rect 13614 32494 13666 32546
rect 13666 32494 13668 32546
rect 13612 32492 13668 32494
rect 13772 32546 13828 32548
rect 13772 32494 13774 32546
rect 13774 32494 13826 32546
rect 13826 32494 13828 32546
rect 13772 32492 13828 32494
rect 13932 32546 13988 32548
rect 13932 32494 13934 32546
rect 13934 32494 13986 32546
rect 13986 32494 13988 32546
rect 13932 32492 13988 32494
rect 14092 32546 14148 32548
rect 14092 32494 14094 32546
rect 14094 32494 14146 32546
rect 14146 32494 14148 32546
rect 14092 32492 14148 32494
rect 14252 32546 14308 32548
rect 14252 32494 14254 32546
rect 14254 32494 14306 32546
rect 14306 32494 14308 32546
rect 14252 32492 14308 32494
rect 14412 32546 14468 32548
rect 14412 32494 14414 32546
rect 14414 32494 14466 32546
rect 14466 32494 14468 32546
rect 14412 32492 14468 32494
rect 14572 32546 14628 32548
rect 14572 32494 14574 32546
rect 14574 32494 14626 32546
rect 14626 32494 14628 32546
rect 14572 32492 14628 32494
rect 14732 32546 14788 32548
rect 14732 32494 14734 32546
rect 14734 32494 14786 32546
rect 14786 32494 14788 32546
rect 14732 32492 14788 32494
rect 14892 32546 14948 32548
rect 14892 32494 14894 32546
rect 14894 32494 14946 32546
rect 14946 32494 14948 32546
rect 14892 32492 14948 32494
rect 15052 32546 15108 32548
rect 15052 32494 15054 32546
rect 15054 32494 15106 32546
rect 15106 32494 15108 32546
rect 15052 32492 15108 32494
rect 15212 32546 15268 32548
rect 15212 32494 15214 32546
rect 15214 32494 15266 32546
rect 15266 32494 15268 32546
rect 15212 32492 15268 32494
rect 15372 32546 15428 32548
rect 15372 32494 15374 32546
rect 15374 32494 15426 32546
rect 15426 32494 15428 32546
rect 15372 32492 15428 32494
rect 15532 32546 15588 32548
rect 15532 32494 15534 32546
rect 15534 32494 15586 32546
rect 15586 32494 15588 32546
rect 15532 32492 15588 32494
rect 15692 32546 15748 32548
rect 15692 32494 15694 32546
rect 15694 32494 15746 32546
rect 15746 32494 15748 32546
rect 15692 32492 15748 32494
rect 15852 32546 15908 32548
rect 15852 32494 15854 32546
rect 15854 32494 15906 32546
rect 15906 32494 15908 32546
rect 15852 32492 15908 32494
rect 16012 32546 16068 32548
rect 16012 32494 16014 32546
rect 16014 32494 16066 32546
rect 16066 32494 16068 32546
rect 16012 32492 16068 32494
rect 16172 32546 16228 32548
rect 16172 32494 16174 32546
rect 16174 32494 16226 32546
rect 16226 32494 16228 32546
rect 16172 32492 16228 32494
rect 16332 32546 16388 32548
rect 16332 32494 16334 32546
rect 16334 32494 16386 32546
rect 16386 32494 16388 32546
rect 16332 32492 16388 32494
rect 16492 32546 16548 32548
rect 16492 32494 16494 32546
rect 16494 32494 16546 32546
rect 16546 32494 16548 32546
rect 16492 32492 16548 32494
rect 16652 32546 16708 32548
rect 16652 32494 16654 32546
rect 16654 32494 16706 32546
rect 16706 32494 16708 32546
rect 16652 32492 16708 32494
rect 16812 32546 16868 32548
rect 16812 32494 16814 32546
rect 16814 32494 16866 32546
rect 16866 32494 16868 32546
rect 16812 32492 16868 32494
rect 16972 32546 17028 32548
rect 16972 32494 16974 32546
rect 16974 32494 17026 32546
rect 17026 32494 17028 32546
rect 16972 32492 17028 32494
rect 17132 32546 17188 32548
rect 17132 32494 17134 32546
rect 17134 32494 17186 32546
rect 17186 32494 17188 32546
rect 17132 32492 17188 32494
rect 17292 32546 17348 32548
rect 17292 32494 17294 32546
rect 17294 32494 17346 32546
rect 17346 32494 17348 32546
rect 17292 32492 17348 32494
rect 17452 32546 17508 32548
rect 17452 32494 17454 32546
rect 17454 32494 17506 32546
rect 17506 32494 17508 32546
rect 17452 32492 17508 32494
rect 17612 32546 17668 32548
rect 17612 32494 17614 32546
rect 17614 32494 17666 32546
rect 17666 32494 17668 32546
rect 17612 32492 17668 32494
rect 17772 32546 17828 32548
rect 17772 32494 17774 32546
rect 17774 32494 17826 32546
rect 17826 32494 17828 32546
rect 17772 32492 17828 32494
rect 17932 32546 17988 32548
rect 17932 32494 17934 32546
rect 17934 32494 17986 32546
rect 17986 32494 17988 32546
rect 17932 32492 17988 32494
rect 18092 32546 18148 32548
rect 18092 32494 18094 32546
rect 18094 32494 18146 32546
rect 18146 32494 18148 32546
rect 18092 32492 18148 32494
rect 18252 32546 18308 32548
rect 18252 32494 18254 32546
rect 18254 32494 18306 32546
rect 18306 32494 18308 32546
rect 18252 32492 18308 32494
rect 18412 32546 18468 32548
rect 18412 32494 18414 32546
rect 18414 32494 18466 32546
rect 18466 32494 18468 32546
rect 18412 32492 18468 32494
rect 18572 32546 18628 32548
rect 18572 32494 18574 32546
rect 18574 32494 18626 32546
rect 18626 32494 18628 32546
rect 18572 32492 18628 32494
rect 18732 32546 18788 32548
rect 18732 32494 18734 32546
rect 18734 32494 18786 32546
rect 18786 32494 18788 32546
rect 18732 32492 18788 32494
rect 18892 32546 18948 32548
rect 18892 32494 18894 32546
rect 18894 32494 18946 32546
rect 18946 32494 18948 32546
rect 18892 32492 18948 32494
rect 19532 32492 19588 32548
rect 19852 32492 19908 32548
rect 23132 32546 23188 32548
rect 23132 32494 23134 32546
rect 23134 32494 23186 32546
rect 23186 32494 23188 32546
rect 23132 32492 23188 32494
rect 23292 32546 23348 32548
rect 23292 32494 23294 32546
rect 23294 32494 23346 32546
rect 23346 32494 23348 32546
rect 23292 32492 23348 32494
rect 23452 32546 23508 32548
rect 23452 32494 23454 32546
rect 23454 32494 23506 32546
rect 23506 32494 23508 32546
rect 23452 32492 23508 32494
rect 23612 32546 23668 32548
rect 23612 32494 23614 32546
rect 23614 32494 23666 32546
rect 23666 32494 23668 32546
rect 23612 32492 23668 32494
rect 23772 32546 23828 32548
rect 23772 32494 23774 32546
rect 23774 32494 23826 32546
rect 23826 32494 23828 32546
rect 23772 32492 23828 32494
rect 23932 32546 23988 32548
rect 23932 32494 23934 32546
rect 23934 32494 23986 32546
rect 23986 32494 23988 32546
rect 23932 32492 23988 32494
rect 24092 32546 24148 32548
rect 24092 32494 24094 32546
rect 24094 32494 24146 32546
rect 24146 32494 24148 32546
rect 24092 32492 24148 32494
rect 24252 32546 24308 32548
rect 24252 32494 24254 32546
rect 24254 32494 24306 32546
rect 24306 32494 24308 32546
rect 24252 32492 24308 32494
rect 24412 32546 24468 32548
rect 24412 32494 24414 32546
rect 24414 32494 24466 32546
rect 24466 32494 24468 32546
rect 24412 32492 24468 32494
rect 24572 32546 24628 32548
rect 24572 32494 24574 32546
rect 24574 32494 24626 32546
rect 24626 32494 24628 32546
rect 24572 32492 24628 32494
rect 24732 32546 24788 32548
rect 24732 32494 24734 32546
rect 24734 32494 24786 32546
rect 24786 32494 24788 32546
rect 24732 32492 24788 32494
rect 24892 32546 24948 32548
rect 24892 32494 24894 32546
rect 24894 32494 24946 32546
rect 24946 32494 24948 32546
rect 24892 32492 24948 32494
rect 25052 32546 25108 32548
rect 25052 32494 25054 32546
rect 25054 32494 25106 32546
rect 25106 32494 25108 32546
rect 25052 32492 25108 32494
rect 25212 32546 25268 32548
rect 25212 32494 25214 32546
rect 25214 32494 25266 32546
rect 25266 32494 25268 32546
rect 25212 32492 25268 32494
rect 25372 32546 25428 32548
rect 25372 32494 25374 32546
rect 25374 32494 25426 32546
rect 25426 32494 25428 32546
rect 25372 32492 25428 32494
rect 25532 32546 25588 32548
rect 25532 32494 25534 32546
rect 25534 32494 25586 32546
rect 25586 32494 25588 32546
rect 25532 32492 25588 32494
rect 25692 32546 25748 32548
rect 25692 32494 25694 32546
rect 25694 32494 25746 32546
rect 25746 32494 25748 32546
rect 25692 32492 25748 32494
rect 25852 32546 25908 32548
rect 25852 32494 25854 32546
rect 25854 32494 25906 32546
rect 25906 32494 25908 32546
rect 25852 32492 25908 32494
rect 26012 32546 26068 32548
rect 26012 32494 26014 32546
rect 26014 32494 26066 32546
rect 26066 32494 26068 32546
rect 26012 32492 26068 32494
rect 26172 32546 26228 32548
rect 26172 32494 26174 32546
rect 26174 32494 26226 32546
rect 26226 32494 26228 32546
rect 26172 32492 26228 32494
rect 26332 32546 26388 32548
rect 26332 32494 26334 32546
rect 26334 32494 26386 32546
rect 26386 32494 26388 32546
rect 26332 32492 26388 32494
rect 26492 32546 26548 32548
rect 26492 32494 26494 32546
rect 26494 32494 26546 32546
rect 26546 32494 26548 32546
rect 26492 32492 26548 32494
rect 26652 32546 26708 32548
rect 26652 32494 26654 32546
rect 26654 32494 26706 32546
rect 26706 32494 26708 32546
rect 26652 32492 26708 32494
rect 26812 32546 26868 32548
rect 26812 32494 26814 32546
rect 26814 32494 26866 32546
rect 26866 32494 26868 32546
rect 26812 32492 26868 32494
rect 26972 32546 27028 32548
rect 26972 32494 26974 32546
rect 26974 32494 27026 32546
rect 27026 32494 27028 32546
rect 26972 32492 27028 32494
rect 27132 32546 27188 32548
rect 27132 32494 27134 32546
rect 27134 32494 27186 32546
rect 27186 32494 27188 32546
rect 27132 32492 27188 32494
rect 27292 32546 27348 32548
rect 27292 32494 27294 32546
rect 27294 32494 27346 32546
rect 27346 32494 27348 32546
rect 27292 32492 27348 32494
rect 27452 32546 27508 32548
rect 27452 32494 27454 32546
rect 27454 32494 27506 32546
rect 27506 32494 27508 32546
rect 27452 32492 27508 32494
rect 27612 32546 27668 32548
rect 27612 32494 27614 32546
rect 27614 32494 27666 32546
rect 27666 32494 27668 32546
rect 27612 32492 27668 32494
rect 27772 32546 27828 32548
rect 27772 32494 27774 32546
rect 27774 32494 27826 32546
rect 27826 32494 27828 32546
rect 27772 32492 27828 32494
rect 27932 32546 27988 32548
rect 27932 32494 27934 32546
rect 27934 32494 27986 32546
rect 27986 32494 27988 32546
rect 27932 32492 27988 32494
rect 28092 32546 28148 32548
rect 28092 32494 28094 32546
rect 28094 32494 28146 32546
rect 28146 32494 28148 32546
rect 28092 32492 28148 32494
rect 28252 32546 28308 32548
rect 28252 32494 28254 32546
rect 28254 32494 28306 32546
rect 28306 32494 28308 32546
rect 28252 32492 28308 32494
rect 28412 32546 28468 32548
rect 28412 32494 28414 32546
rect 28414 32494 28466 32546
rect 28466 32494 28468 32546
rect 28412 32492 28468 32494
rect 28572 32546 28628 32548
rect 28572 32494 28574 32546
rect 28574 32494 28626 32546
rect 28626 32494 28628 32546
rect 28572 32492 28628 32494
rect 28732 32546 28788 32548
rect 28732 32494 28734 32546
rect 28734 32494 28786 32546
rect 28786 32494 28788 32546
rect 28732 32492 28788 32494
rect 28892 32546 28948 32548
rect 28892 32494 28894 32546
rect 28894 32494 28946 32546
rect 28946 32494 28948 32546
rect 28892 32492 28948 32494
rect 29052 32546 29108 32548
rect 29052 32494 29054 32546
rect 29054 32494 29106 32546
rect 29106 32494 29108 32546
rect 29052 32492 29108 32494
rect 29212 32546 29268 32548
rect 29212 32494 29214 32546
rect 29214 32494 29266 32546
rect 29266 32494 29268 32546
rect 29212 32492 29268 32494
rect 29372 32546 29428 32548
rect 29372 32494 29374 32546
rect 29374 32494 29426 32546
rect 29426 32494 29428 32546
rect 29372 32492 29428 32494
rect 32572 32492 32628 32548
rect 32892 32492 32948 32548
rect 33532 32546 33588 32548
rect 33532 32494 33534 32546
rect 33534 32494 33586 32546
rect 33586 32494 33588 32546
rect 33532 32492 33588 32494
rect 33692 32546 33748 32548
rect 33692 32494 33694 32546
rect 33694 32494 33746 32546
rect 33746 32494 33748 32546
rect 33692 32492 33748 32494
rect 33852 32546 33908 32548
rect 33852 32494 33854 32546
rect 33854 32494 33906 32546
rect 33906 32494 33908 32546
rect 33852 32492 33908 32494
rect 34012 32546 34068 32548
rect 34012 32494 34014 32546
rect 34014 32494 34066 32546
rect 34066 32494 34068 32546
rect 34012 32492 34068 32494
rect 34172 32546 34228 32548
rect 34172 32494 34174 32546
rect 34174 32494 34226 32546
rect 34226 32494 34228 32546
rect 34172 32492 34228 32494
rect 34332 32546 34388 32548
rect 34332 32494 34334 32546
rect 34334 32494 34386 32546
rect 34386 32494 34388 32546
rect 34332 32492 34388 32494
rect 34492 32546 34548 32548
rect 34492 32494 34494 32546
rect 34494 32494 34546 32546
rect 34546 32494 34548 32546
rect 34492 32492 34548 32494
rect 34652 32546 34708 32548
rect 34652 32494 34654 32546
rect 34654 32494 34706 32546
rect 34706 32494 34708 32546
rect 34652 32492 34708 32494
rect 34812 32546 34868 32548
rect 34812 32494 34814 32546
rect 34814 32494 34866 32546
rect 34866 32494 34868 32546
rect 34812 32492 34868 32494
rect 34972 32546 35028 32548
rect 34972 32494 34974 32546
rect 34974 32494 35026 32546
rect 35026 32494 35028 32546
rect 34972 32492 35028 32494
rect 35132 32546 35188 32548
rect 35132 32494 35134 32546
rect 35134 32494 35186 32546
rect 35186 32494 35188 32546
rect 35132 32492 35188 32494
rect 35292 32546 35348 32548
rect 35292 32494 35294 32546
rect 35294 32494 35346 32546
rect 35346 32494 35348 32546
rect 35292 32492 35348 32494
rect 35452 32546 35508 32548
rect 35452 32494 35454 32546
rect 35454 32494 35506 32546
rect 35506 32494 35508 32546
rect 35452 32492 35508 32494
rect 35612 32546 35668 32548
rect 35612 32494 35614 32546
rect 35614 32494 35666 32546
rect 35666 32494 35668 32546
rect 35612 32492 35668 32494
rect 35772 32546 35828 32548
rect 35772 32494 35774 32546
rect 35774 32494 35826 32546
rect 35826 32494 35828 32546
rect 35772 32492 35828 32494
rect 35932 32546 35988 32548
rect 35932 32494 35934 32546
rect 35934 32494 35986 32546
rect 35986 32494 35988 32546
rect 35932 32492 35988 32494
rect 36092 32546 36148 32548
rect 36092 32494 36094 32546
rect 36094 32494 36146 32546
rect 36146 32494 36148 32546
rect 36092 32492 36148 32494
rect 36252 32546 36308 32548
rect 36252 32494 36254 32546
rect 36254 32494 36306 32546
rect 36306 32494 36308 32546
rect 36252 32492 36308 32494
rect 36412 32546 36468 32548
rect 36412 32494 36414 32546
rect 36414 32494 36466 32546
rect 36466 32494 36468 32546
rect 36412 32492 36468 32494
rect 36572 32546 36628 32548
rect 36572 32494 36574 32546
rect 36574 32494 36626 32546
rect 36626 32494 36628 32546
rect 36572 32492 36628 32494
rect 36732 32546 36788 32548
rect 36732 32494 36734 32546
rect 36734 32494 36786 32546
rect 36786 32494 36788 32546
rect 36732 32492 36788 32494
rect 36892 32546 36948 32548
rect 36892 32494 36894 32546
rect 36894 32494 36946 32546
rect 36946 32494 36948 32546
rect 36892 32492 36948 32494
rect 37052 32546 37108 32548
rect 37052 32494 37054 32546
rect 37054 32494 37106 32546
rect 37106 32494 37108 32546
rect 37052 32492 37108 32494
rect 37212 32546 37268 32548
rect 37212 32494 37214 32546
rect 37214 32494 37266 32546
rect 37266 32494 37268 32546
rect 37212 32492 37268 32494
rect 37372 32546 37428 32548
rect 37372 32494 37374 32546
rect 37374 32494 37426 32546
rect 37426 32494 37428 32546
rect 37372 32492 37428 32494
rect 37532 32546 37588 32548
rect 37532 32494 37534 32546
rect 37534 32494 37586 32546
rect 37586 32494 37588 32546
rect 37532 32492 37588 32494
rect 37692 32546 37748 32548
rect 37692 32494 37694 32546
rect 37694 32494 37746 32546
rect 37746 32494 37748 32546
rect 37692 32492 37748 32494
rect 37852 32546 37908 32548
rect 37852 32494 37854 32546
rect 37854 32494 37906 32546
rect 37906 32494 37908 32546
rect 37852 32492 37908 32494
rect 38012 32546 38068 32548
rect 38012 32494 38014 32546
rect 38014 32494 38066 32546
rect 38066 32494 38068 32546
rect 38012 32492 38068 32494
rect 38172 32546 38228 32548
rect 38172 32494 38174 32546
rect 38174 32494 38226 32546
rect 38226 32494 38228 32546
rect 38172 32492 38228 32494
rect 38332 32546 38388 32548
rect 38332 32494 38334 32546
rect 38334 32494 38386 32546
rect 38386 32494 38388 32546
rect 38332 32492 38388 32494
rect 38492 32546 38548 32548
rect 38492 32494 38494 32546
rect 38494 32494 38546 32546
rect 38546 32494 38548 32546
rect 38492 32492 38548 32494
rect 38652 32546 38708 32548
rect 38652 32494 38654 32546
rect 38654 32494 38706 32546
rect 38706 32494 38708 32546
rect 38652 32492 38708 32494
rect 38812 32546 38868 32548
rect 38812 32494 38814 32546
rect 38814 32494 38866 32546
rect 38866 32494 38868 32546
rect 38812 32492 38868 32494
rect 38972 32546 39028 32548
rect 38972 32494 38974 32546
rect 38974 32494 39026 32546
rect 39026 32494 39028 32546
rect 38972 32492 39028 32494
rect 39132 32546 39188 32548
rect 39132 32494 39134 32546
rect 39134 32494 39186 32546
rect 39186 32494 39188 32546
rect 39132 32492 39188 32494
rect 39292 32546 39348 32548
rect 39292 32494 39294 32546
rect 39294 32494 39346 32546
rect 39346 32494 39348 32546
rect 39292 32492 39348 32494
rect 39452 32546 39508 32548
rect 39452 32494 39454 32546
rect 39454 32494 39506 32546
rect 39506 32494 39508 32546
rect 39452 32492 39508 32494
rect 39612 32546 39668 32548
rect 39612 32494 39614 32546
rect 39614 32494 39666 32546
rect 39666 32494 39668 32546
rect 39612 32492 39668 32494
rect 39772 32546 39828 32548
rect 39772 32494 39774 32546
rect 39774 32494 39826 32546
rect 39826 32494 39828 32546
rect 39772 32492 39828 32494
rect 39932 32546 39988 32548
rect 39932 32494 39934 32546
rect 39934 32494 39986 32546
rect 39986 32494 39988 32546
rect 39932 32492 39988 32494
rect 40092 32546 40148 32548
rect 40092 32494 40094 32546
rect 40094 32494 40146 32546
rect 40146 32494 40148 32546
rect 40092 32492 40148 32494
rect 40252 32546 40308 32548
rect 40252 32494 40254 32546
rect 40254 32494 40306 32546
rect 40306 32494 40308 32546
rect 40252 32492 40308 32494
rect 40412 32546 40468 32548
rect 40412 32494 40414 32546
rect 40414 32494 40466 32546
rect 40466 32494 40468 32546
rect 40412 32492 40468 32494
rect 40572 32546 40628 32548
rect 40572 32494 40574 32546
rect 40574 32494 40626 32546
rect 40626 32494 40628 32546
rect 40572 32492 40628 32494
rect 40732 32546 40788 32548
rect 40732 32494 40734 32546
rect 40734 32494 40786 32546
rect 40786 32494 40788 32546
rect 40732 32492 40788 32494
rect 40892 32546 40948 32548
rect 40892 32494 40894 32546
rect 40894 32494 40946 32546
rect 40946 32494 40948 32546
rect 40892 32492 40948 32494
rect 41052 32546 41108 32548
rect 41052 32494 41054 32546
rect 41054 32494 41106 32546
rect 41106 32494 41108 32546
rect 41052 32492 41108 32494
rect 41212 32546 41268 32548
rect 41212 32494 41214 32546
rect 41214 32494 41266 32546
rect 41266 32494 41268 32546
rect 41212 32492 41268 32494
rect 41372 32546 41428 32548
rect 41372 32494 41374 32546
rect 41374 32494 41426 32546
rect 41426 32494 41428 32546
rect 41372 32492 41428 32494
rect 41532 32546 41588 32548
rect 41532 32494 41534 32546
rect 41534 32494 41586 32546
rect 41586 32494 41588 32546
rect 41532 32492 41588 32494
rect 41692 32546 41748 32548
rect 41692 32494 41694 32546
rect 41694 32494 41746 32546
rect 41746 32494 41748 32546
rect 41692 32492 41748 32494
rect 41852 32546 41908 32548
rect 41852 32494 41854 32546
rect 41854 32494 41906 32546
rect 41906 32494 41908 32546
rect 41852 32492 41908 32494
rect 12 32386 68 32388
rect 12 32334 14 32386
rect 14 32334 66 32386
rect 66 32334 68 32386
rect 12 32332 68 32334
rect 172 32386 228 32388
rect 172 32334 174 32386
rect 174 32334 226 32386
rect 226 32334 228 32386
rect 172 32332 228 32334
rect 332 32386 388 32388
rect 332 32334 334 32386
rect 334 32334 386 32386
rect 386 32334 388 32386
rect 332 32332 388 32334
rect 492 32386 548 32388
rect 492 32334 494 32386
rect 494 32334 546 32386
rect 546 32334 548 32386
rect 492 32332 548 32334
rect 652 32386 708 32388
rect 652 32334 654 32386
rect 654 32334 706 32386
rect 706 32334 708 32386
rect 652 32332 708 32334
rect 812 32386 868 32388
rect 812 32334 814 32386
rect 814 32334 866 32386
rect 866 32334 868 32386
rect 812 32332 868 32334
rect 972 32386 1028 32388
rect 972 32334 974 32386
rect 974 32334 1026 32386
rect 1026 32334 1028 32386
rect 972 32332 1028 32334
rect 1132 32386 1188 32388
rect 1132 32334 1134 32386
rect 1134 32334 1186 32386
rect 1186 32334 1188 32386
rect 1132 32332 1188 32334
rect 1292 32386 1348 32388
rect 1292 32334 1294 32386
rect 1294 32334 1346 32386
rect 1346 32334 1348 32386
rect 1292 32332 1348 32334
rect 1452 32386 1508 32388
rect 1452 32334 1454 32386
rect 1454 32334 1506 32386
rect 1506 32334 1508 32386
rect 1452 32332 1508 32334
rect 1612 32386 1668 32388
rect 1612 32334 1614 32386
rect 1614 32334 1666 32386
rect 1666 32334 1668 32386
rect 1612 32332 1668 32334
rect 1772 32386 1828 32388
rect 1772 32334 1774 32386
rect 1774 32334 1826 32386
rect 1826 32334 1828 32386
rect 1772 32332 1828 32334
rect 1932 32386 1988 32388
rect 1932 32334 1934 32386
rect 1934 32334 1986 32386
rect 1986 32334 1988 32386
rect 1932 32332 1988 32334
rect 2092 32386 2148 32388
rect 2092 32334 2094 32386
rect 2094 32334 2146 32386
rect 2146 32334 2148 32386
rect 2092 32332 2148 32334
rect 2252 32386 2308 32388
rect 2252 32334 2254 32386
rect 2254 32334 2306 32386
rect 2306 32334 2308 32386
rect 2252 32332 2308 32334
rect 2412 32386 2468 32388
rect 2412 32334 2414 32386
rect 2414 32334 2466 32386
rect 2466 32334 2468 32386
rect 2412 32332 2468 32334
rect 2572 32386 2628 32388
rect 2572 32334 2574 32386
rect 2574 32334 2626 32386
rect 2626 32334 2628 32386
rect 2572 32332 2628 32334
rect 2732 32386 2788 32388
rect 2732 32334 2734 32386
rect 2734 32334 2786 32386
rect 2786 32334 2788 32386
rect 2732 32332 2788 32334
rect 2892 32386 2948 32388
rect 2892 32334 2894 32386
rect 2894 32334 2946 32386
rect 2946 32334 2948 32386
rect 2892 32332 2948 32334
rect 3052 32386 3108 32388
rect 3052 32334 3054 32386
rect 3054 32334 3106 32386
rect 3106 32334 3108 32386
rect 3052 32332 3108 32334
rect 3212 32386 3268 32388
rect 3212 32334 3214 32386
rect 3214 32334 3266 32386
rect 3266 32334 3268 32386
rect 3212 32332 3268 32334
rect 3372 32386 3428 32388
rect 3372 32334 3374 32386
rect 3374 32334 3426 32386
rect 3426 32334 3428 32386
rect 3372 32332 3428 32334
rect 3532 32386 3588 32388
rect 3532 32334 3534 32386
rect 3534 32334 3586 32386
rect 3586 32334 3588 32386
rect 3532 32332 3588 32334
rect 3692 32386 3748 32388
rect 3692 32334 3694 32386
rect 3694 32334 3746 32386
rect 3746 32334 3748 32386
rect 3692 32332 3748 32334
rect 3852 32386 3908 32388
rect 3852 32334 3854 32386
rect 3854 32334 3906 32386
rect 3906 32334 3908 32386
rect 3852 32332 3908 32334
rect 4012 32386 4068 32388
rect 4012 32334 4014 32386
rect 4014 32334 4066 32386
rect 4066 32334 4068 32386
rect 4012 32332 4068 32334
rect 4172 32386 4228 32388
rect 4172 32334 4174 32386
rect 4174 32334 4226 32386
rect 4226 32334 4228 32386
rect 4172 32332 4228 32334
rect 4332 32386 4388 32388
rect 4332 32334 4334 32386
rect 4334 32334 4386 32386
rect 4386 32334 4388 32386
rect 4332 32332 4388 32334
rect 4492 32386 4548 32388
rect 4492 32334 4494 32386
rect 4494 32334 4546 32386
rect 4546 32334 4548 32386
rect 4492 32332 4548 32334
rect 4652 32386 4708 32388
rect 4652 32334 4654 32386
rect 4654 32334 4706 32386
rect 4706 32334 4708 32386
rect 4652 32332 4708 32334
rect 4812 32386 4868 32388
rect 4812 32334 4814 32386
rect 4814 32334 4866 32386
rect 4866 32334 4868 32386
rect 4812 32332 4868 32334
rect 4972 32386 5028 32388
rect 4972 32334 4974 32386
rect 4974 32334 5026 32386
rect 5026 32334 5028 32386
rect 4972 32332 5028 32334
rect 5132 32386 5188 32388
rect 5132 32334 5134 32386
rect 5134 32334 5186 32386
rect 5186 32334 5188 32386
rect 5132 32332 5188 32334
rect 5292 32386 5348 32388
rect 5292 32334 5294 32386
rect 5294 32334 5346 32386
rect 5346 32334 5348 32386
rect 5292 32332 5348 32334
rect 5452 32386 5508 32388
rect 5452 32334 5454 32386
rect 5454 32334 5506 32386
rect 5506 32334 5508 32386
rect 5452 32332 5508 32334
rect 5612 32386 5668 32388
rect 5612 32334 5614 32386
rect 5614 32334 5666 32386
rect 5666 32334 5668 32386
rect 5612 32332 5668 32334
rect 5772 32386 5828 32388
rect 5772 32334 5774 32386
rect 5774 32334 5826 32386
rect 5826 32334 5828 32386
rect 5772 32332 5828 32334
rect 5932 32386 5988 32388
rect 5932 32334 5934 32386
rect 5934 32334 5986 32386
rect 5986 32334 5988 32386
rect 5932 32332 5988 32334
rect 6092 32386 6148 32388
rect 6092 32334 6094 32386
rect 6094 32334 6146 32386
rect 6146 32334 6148 32386
rect 6092 32332 6148 32334
rect 6252 32386 6308 32388
rect 6252 32334 6254 32386
rect 6254 32334 6306 32386
rect 6306 32334 6308 32386
rect 6252 32332 6308 32334
rect 6412 32386 6468 32388
rect 6412 32334 6414 32386
rect 6414 32334 6466 32386
rect 6466 32334 6468 32386
rect 6412 32332 6468 32334
rect 6572 32386 6628 32388
rect 6572 32334 6574 32386
rect 6574 32334 6626 32386
rect 6626 32334 6628 32386
rect 6572 32332 6628 32334
rect 6732 32386 6788 32388
rect 6732 32334 6734 32386
rect 6734 32334 6786 32386
rect 6786 32334 6788 32386
rect 6732 32332 6788 32334
rect 6892 32386 6948 32388
rect 6892 32334 6894 32386
rect 6894 32334 6946 32386
rect 6946 32334 6948 32386
rect 6892 32332 6948 32334
rect 7052 32386 7108 32388
rect 7052 32334 7054 32386
rect 7054 32334 7106 32386
rect 7106 32334 7108 32386
rect 7052 32332 7108 32334
rect 7212 32386 7268 32388
rect 7212 32334 7214 32386
rect 7214 32334 7266 32386
rect 7266 32334 7268 32386
rect 7212 32332 7268 32334
rect 7372 32386 7428 32388
rect 7372 32334 7374 32386
rect 7374 32334 7426 32386
rect 7426 32334 7428 32386
rect 7372 32332 7428 32334
rect 7532 32386 7588 32388
rect 7532 32334 7534 32386
rect 7534 32334 7586 32386
rect 7586 32334 7588 32386
rect 7532 32332 7588 32334
rect 7692 32386 7748 32388
rect 7692 32334 7694 32386
rect 7694 32334 7746 32386
rect 7746 32334 7748 32386
rect 7692 32332 7748 32334
rect 7852 32386 7908 32388
rect 7852 32334 7854 32386
rect 7854 32334 7906 32386
rect 7906 32334 7908 32386
rect 7852 32332 7908 32334
rect 8012 32386 8068 32388
rect 8012 32334 8014 32386
rect 8014 32334 8066 32386
rect 8066 32334 8068 32386
rect 8012 32332 8068 32334
rect 8172 32386 8228 32388
rect 8172 32334 8174 32386
rect 8174 32334 8226 32386
rect 8226 32334 8228 32386
rect 8172 32332 8228 32334
rect 8332 32386 8388 32388
rect 8332 32334 8334 32386
rect 8334 32334 8386 32386
rect 8386 32334 8388 32386
rect 8332 32332 8388 32334
rect 9452 32332 9508 32388
rect 9772 32332 9828 32388
rect 10092 32332 10148 32388
rect 10412 32332 10468 32388
rect 10732 32332 10788 32388
rect 11052 32332 11108 32388
rect 11372 32332 11428 32388
rect 12492 32386 12548 32388
rect 12492 32334 12494 32386
rect 12494 32334 12546 32386
rect 12546 32334 12548 32386
rect 12492 32332 12548 32334
rect 12652 32386 12708 32388
rect 12652 32334 12654 32386
rect 12654 32334 12706 32386
rect 12706 32334 12708 32386
rect 12652 32332 12708 32334
rect 12812 32386 12868 32388
rect 12812 32334 12814 32386
rect 12814 32334 12866 32386
rect 12866 32334 12868 32386
rect 12812 32332 12868 32334
rect 12972 32386 13028 32388
rect 12972 32334 12974 32386
rect 12974 32334 13026 32386
rect 13026 32334 13028 32386
rect 12972 32332 13028 32334
rect 13132 32386 13188 32388
rect 13132 32334 13134 32386
rect 13134 32334 13186 32386
rect 13186 32334 13188 32386
rect 13132 32332 13188 32334
rect 13292 32386 13348 32388
rect 13292 32334 13294 32386
rect 13294 32334 13346 32386
rect 13346 32334 13348 32386
rect 13292 32332 13348 32334
rect 13452 32386 13508 32388
rect 13452 32334 13454 32386
rect 13454 32334 13506 32386
rect 13506 32334 13508 32386
rect 13452 32332 13508 32334
rect 13612 32386 13668 32388
rect 13612 32334 13614 32386
rect 13614 32334 13666 32386
rect 13666 32334 13668 32386
rect 13612 32332 13668 32334
rect 13772 32386 13828 32388
rect 13772 32334 13774 32386
rect 13774 32334 13826 32386
rect 13826 32334 13828 32386
rect 13772 32332 13828 32334
rect 13932 32386 13988 32388
rect 13932 32334 13934 32386
rect 13934 32334 13986 32386
rect 13986 32334 13988 32386
rect 13932 32332 13988 32334
rect 14092 32386 14148 32388
rect 14092 32334 14094 32386
rect 14094 32334 14146 32386
rect 14146 32334 14148 32386
rect 14092 32332 14148 32334
rect 14252 32386 14308 32388
rect 14252 32334 14254 32386
rect 14254 32334 14306 32386
rect 14306 32334 14308 32386
rect 14252 32332 14308 32334
rect 14412 32386 14468 32388
rect 14412 32334 14414 32386
rect 14414 32334 14466 32386
rect 14466 32334 14468 32386
rect 14412 32332 14468 32334
rect 14572 32386 14628 32388
rect 14572 32334 14574 32386
rect 14574 32334 14626 32386
rect 14626 32334 14628 32386
rect 14572 32332 14628 32334
rect 14732 32386 14788 32388
rect 14732 32334 14734 32386
rect 14734 32334 14786 32386
rect 14786 32334 14788 32386
rect 14732 32332 14788 32334
rect 14892 32386 14948 32388
rect 14892 32334 14894 32386
rect 14894 32334 14946 32386
rect 14946 32334 14948 32386
rect 14892 32332 14948 32334
rect 15052 32386 15108 32388
rect 15052 32334 15054 32386
rect 15054 32334 15106 32386
rect 15106 32334 15108 32386
rect 15052 32332 15108 32334
rect 15212 32386 15268 32388
rect 15212 32334 15214 32386
rect 15214 32334 15266 32386
rect 15266 32334 15268 32386
rect 15212 32332 15268 32334
rect 15372 32386 15428 32388
rect 15372 32334 15374 32386
rect 15374 32334 15426 32386
rect 15426 32334 15428 32386
rect 15372 32332 15428 32334
rect 15532 32386 15588 32388
rect 15532 32334 15534 32386
rect 15534 32334 15586 32386
rect 15586 32334 15588 32386
rect 15532 32332 15588 32334
rect 15692 32386 15748 32388
rect 15692 32334 15694 32386
rect 15694 32334 15746 32386
rect 15746 32334 15748 32386
rect 15692 32332 15748 32334
rect 15852 32386 15908 32388
rect 15852 32334 15854 32386
rect 15854 32334 15906 32386
rect 15906 32334 15908 32386
rect 15852 32332 15908 32334
rect 16012 32386 16068 32388
rect 16012 32334 16014 32386
rect 16014 32334 16066 32386
rect 16066 32334 16068 32386
rect 16012 32332 16068 32334
rect 16172 32386 16228 32388
rect 16172 32334 16174 32386
rect 16174 32334 16226 32386
rect 16226 32334 16228 32386
rect 16172 32332 16228 32334
rect 16332 32386 16388 32388
rect 16332 32334 16334 32386
rect 16334 32334 16386 32386
rect 16386 32334 16388 32386
rect 16332 32332 16388 32334
rect 16492 32386 16548 32388
rect 16492 32334 16494 32386
rect 16494 32334 16546 32386
rect 16546 32334 16548 32386
rect 16492 32332 16548 32334
rect 16652 32386 16708 32388
rect 16652 32334 16654 32386
rect 16654 32334 16706 32386
rect 16706 32334 16708 32386
rect 16652 32332 16708 32334
rect 16812 32386 16868 32388
rect 16812 32334 16814 32386
rect 16814 32334 16866 32386
rect 16866 32334 16868 32386
rect 16812 32332 16868 32334
rect 16972 32386 17028 32388
rect 16972 32334 16974 32386
rect 16974 32334 17026 32386
rect 17026 32334 17028 32386
rect 16972 32332 17028 32334
rect 17132 32386 17188 32388
rect 17132 32334 17134 32386
rect 17134 32334 17186 32386
rect 17186 32334 17188 32386
rect 17132 32332 17188 32334
rect 17292 32386 17348 32388
rect 17292 32334 17294 32386
rect 17294 32334 17346 32386
rect 17346 32334 17348 32386
rect 17292 32332 17348 32334
rect 17452 32386 17508 32388
rect 17452 32334 17454 32386
rect 17454 32334 17506 32386
rect 17506 32334 17508 32386
rect 17452 32332 17508 32334
rect 17612 32386 17668 32388
rect 17612 32334 17614 32386
rect 17614 32334 17666 32386
rect 17666 32334 17668 32386
rect 17612 32332 17668 32334
rect 17772 32386 17828 32388
rect 17772 32334 17774 32386
rect 17774 32334 17826 32386
rect 17826 32334 17828 32386
rect 17772 32332 17828 32334
rect 17932 32386 17988 32388
rect 17932 32334 17934 32386
rect 17934 32334 17986 32386
rect 17986 32334 17988 32386
rect 17932 32332 17988 32334
rect 18092 32386 18148 32388
rect 18092 32334 18094 32386
rect 18094 32334 18146 32386
rect 18146 32334 18148 32386
rect 18092 32332 18148 32334
rect 18252 32386 18308 32388
rect 18252 32334 18254 32386
rect 18254 32334 18306 32386
rect 18306 32334 18308 32386
rect 18252 32332 18308 32334
rect 18412 32386 18468 32388
rect 18412 32334 18414 32386
rect 18414 32334 18466 32386
rect 18466 32334 18468 32386
rect 18412 32332 18468 32334
rect 18572 32386 18628 32388
rect 18572 32334 18574 32386
rect 18574 32334 18626 32386
rect 18626 32334 18628 32386
rect 18572 32332 18628 32334
rect 18732 32386 18788 32388
rect 18732 32334 18734 32386
rect 18734 32334 18786 32386
rect 18786 32334 18788 32386
rect 18732 32332 18788 32334
rect 18892 32386 18948 32388
rect 18892 32334 18894 32386
rect 18894 32334 18946 32386
rect 18946 32334 18948 32386
rect 18892 32332 18948 32334
rect 20012 32332 20068 32388
rect 20332 32332 20388 32388
rect 20652 32332 20708 32388
rect 20972 32332 21028 32388
rect 21292 32332 21348 32388
rect 21612 32332 21668 32388
rect 21932 32332 21988 32388
rect 23132 32386 23188 32388
rect 23132 32334 23134 32386
rect 23134 32334 23186 32386
rect 23186 32334 23188 32386
rect 23132 32332 23188 32334
rect 23292 32386 23348 32388
rect 23292 32334 23294 32386
rect 23294 32334 23346 32386
rect 23346 32334 23348 32386
rect 23292 32332 23348 32334
rect 23452 32386 23508 32388
rect 23452 32334 23454 32386
rect 23454 32334 23506 32386
rect 23506 32334 23508 32386
rect 23452 32332 23508 32334
rect 23612 32386 23668 32388
rect 23612 32334 23614 32386
rect 23614 32334 23666 32386
rect 23666 32334 23668 32386
rect 23612 32332 23668 32334
rect 23772 32386 23828 32388
rect 23772 32334 23774 32386
rect 23774 32334 23826 32386
rect 23826 32334 23828 32386
rect 23772 32332 23828 32334
rect 23932 32386 23988 32388
rect 23932 32334 23934 32386
rect 23934 32334 23986 32386
rect 23986 32334 23988 32386
rect 23932 32332 23988 32334
rect 24092 32386 24148 32388
rect 24092 32334 24094 32386
rect 24094 32334 24146 32386
rect 24146 32334 24148 32386
rect 24092 32332 24148 32334
rect 24252 32386 24308 32388
rect 24252 32334 24254 32386
rect 24254 32334 24306 32386
rect 24306 32334 24308 32386
rect 24252 32332 24308 32334
rect 24412 32386 24468 32388
rect 24412 32334 24414 32386
rect 24414 32334 24466 32386
rect 24466 32334 24468 32386
rect 24412 32332 24468 32334
rect 24572 32386 24628 32388
rect 24572 32334 24574 32386
rect 24574 32334 24626 32386
rect 24626 32334 24628 32386
rect 24572 32332 24628 32334
rect 24732 32386 24788 32388
rect 24732 32334 24734 32386
rect 24734 32334 24786 32386
rect 24786 32334 24788 32386
rect 24732 32332 24788 32334
rect 24892 32386 24948 32388
rect 24892 32334 24894 32386
rect 24894 32334 24946 32386
rect 24946 32334 24948 32386
rect 24892 32332 24948 32334
rect 25052 32386 25108 32388
rect 25052 32334 25054 32386
rect 25054 32334 25106 32386
rect 25106 32334 25108 32386
rect 25052 32332 25108 32334
rect 25212 32386 25268 32388
rect 25212 32334 25214 32386
rect 25214 32334 25266 32386
rect 25266 32334 25268 32386
rect 25212 32332 25268 32334
rect 25372 32386 25428 32388
rect 25372 32334 25374 32386
rect 25374 32334 25426 32386
rect 25426 32334 25428 32386
rect 25372 32332 25428 32334
rect 25532 32386 25588 32388
rect 25532 32334 25534 32386
rect 25534 32334 25586 32386
rect 25586 32334 25588 32386
rect 25532 32332 25588 32334
rect 25692 32386 25748 32388
rect 25692 32334 25694 32386
rect 25694 32334 25746 32386
rect 25746 32334 25748 32386
rect 25692 32332 25748 32334
rect 25852 32386 25908 32388
rect 25852 32334 25854 32386
rect 25854 32334 25906 32386
rect 25906 32334 25908 32386
rect 25852 32332 25908 32334
rect 26012 32386 26068 32388
rect 26012 32334 26014 32386
rect 26014 32334 26066 32386
rect 26066 32334 26068 32386
rect 26012 32332 26068 32334
rect 26172 32386 26228 32388
rect 26172 32334 26174 32386
rect 26174 32334 26226 32386
rect 26226 32334 26228 32386
rect 26172 32332 26228 32334
rect 26332 32386 26388 32388
rect 26332 32334 26334 32386
rect 26334 32334 26386 32386
rect 26386 32334 26388 32386
rect 26332 32332 26388 32334
rect 26492 32386 26548 32388
rect 26492 32334 26494 32386
rect 26494 32334 26546 32386
rect 26546 32334 26548 32386
rect 26492 32332 26548 32334
rect 26652 32386 26708 32388
rect 26652 32334 26654 32386
rect 26654 32334 26706 32386
rect 26706 32334 26708 32386
rect 26652 32332 26708 32334
rect 26812 32386 26868 32388
rect 26812 32334 26814 32386
rect 26814 32334 26866 32386
rect 26866 32334 26868 32386
rect 26812 32332 26868 32334
rect 26972 32386 27028 32388
rect 26972 32334 26974 32386
rect 26974 32334 27026 32386
rect 27026 32334 27028 32386
rect 26972 32332 27028 32334
rect 27132 32386 27188 32388
rect 27132 32334 27134 32386
rect 27134 32334 27186 32386
rect 27186 32334 27188 32386
rect 27132 32332 27188 32334
rect 27292 32386 27348 32388
rect 27292 32334 27294 32386
rect 27294 32334 27346 32386
rect 27346 32334 27348 32386
rect 27292 32332 27348 32334
rect 27452 32386 27508 32388
rect 27452 32334 27454 32386
rect 27454 32334 27506 32386
rect 27506 32334 27508 32386
rect 27452 32332 27508 32334
rect 27612 32386 27668 32388
rect 27612 32334 27614 32386
rect 27614 32334 27666 32386
rect 27666 32334 27668 32386
rect 27612 32332 27668 32334
rect 27772 32386 27828 32388
rect 27772 32334 27774 32386
rect 27774 32334 27826 32386
rect 27826 32334 27828 32386
rect 27772 32332 27828 32334
rect 27932 32386 27988 32388
rect 27932 32334 27934 32386
rect 27934 32334 27986 32386
rect 27986 32334 27988 32386
rect 27932 32332 27988 32334
rect 28092 32386 28148 32388
rect 28092 32334 28094 32386
rect 28094 32334 28146 32386
rect 28146 32334 28148 32386
rect 28092 32332 28148 32334
rect 28252 32386 28308 32388
rect 28252 32334 28254 32386
rect 28254 32334 28306 32386
rect 28306 32334 28308 32386
rect 28252 32332 28308 32334
rect 28412 32386 28468 32388
rect 28412 32334 28414 32386
rect 28414 32334 28466 32386
rect 28466 32334 28468 32386
rect 28412 32332 28468 32334
rect 28572 32386 28628 32388
rect 28572 32334 28574 32386
rect 28574 32334 28626 32386
rect 28626 32334 28628 32386
rect 28572 32332 28628 32334
rect 28732 32386 28788 32388
rect 28732 32334 28734 32386
rect 28734 32334 28786 32386
rect 28786 32334 28788 32386
rect 28732 32332 28788 32334
rect 28892 32386 28948 32388
rect 28892 32334 28894 32386
rect 28894 32334 28946 32386
rect 28946 32334 28948 32386
rect 28892 32332 28948 32334
rect 29052 32386 29108 32388
rect 29052 32334 29054 32386
rect 29054 32334 29106 32386
rect 29106 32334 29108 32386
rect 29052 32332 29108 32334
rect 29212 32386 29268 32388
rect 29212 32334 29214 32386
rect 29214 32334 29266 32386
rect 29266 32334 29268 32386
rect 29212 32332 29268 32334
rect 29372 32386 29428 32388
rect 29372 32334 29374 32386
rect 29374 32334 29426 32386
rect 29426 32334 29428 32386
rect 29372 32332 29428 32334
rect 30492 32332 30548 32388
rect 30812 32332 30868 32388
rect 31132 32332 31188 32388
rect 31452 32332 31508 32388
rect 31772 32332 31828 32388
rect 32092 32332 32148 32388
rect 32412 32332 32468 32388
rect 33532 32386 33588 32388
rect 33532 32334 33534 32386
rect 33534 32334 33586 32386
rect 33586 32334 33588 32386
rect 33532 32332 33588 32334
rect 33692 32386 33748 32388
rect 33692 32334 33694 32386
rect 33694 32334 33746 32386
rect 33746 32334 33748 32386
rect 33692 32332 33748 32334
rect 33852 32386 33908 32388
rect 33852 32334 33854 32386
rect 33854 32334 33906 32386
rect 33906 32334 33908 32386
rect 33852 32332 33908 32334
rect 34012 32386 34068 32388
rect 34012 32334 34014 32386
rect 34014 32334 34066 32386
rect 34066 32334 34068 32386
rect 34012 32332 34068 32334
rect 34172 32386 34228 32388
rect 34172 32334 34174 32386
rect 34174 32334 34226 32386
rect 34226 32334 34228 32386
rect 34172 32332 34228 32334
rect 34332 32386 34388 32388
rect 34332 32334 34334 32386
rect 34334 32334 34386 32386
rect 34386 32334 34388 32386
rect 34332 32332 34388 32334
rect 34492 32386 34548 32388
rect 34492 32334 34494 32386
rect 34494 32334 34546 32386
rect 34546 32334 34548 32386
rect 34492 32332 34548 32334
rect 34652 32386 34708 32388
rect 34652 32334 34654 32386
rect 34654 32334 34706 32386
rect 34706 32334 34708 32386
rect 34652 32332 34708 32334
rect 34812 32386 34868 32388
rect 34812 32334 34814 32386
rect 34814 32334 34866 32386
rect 34866 32334 34868 32386
rect 34812 32332 34868 32334
rect 34972 32386 35028 32388
rect 34972 32334 34974 32386
rect 34974 32334 35026 32386
rect 35026 32334 35028 32386
rect 34972 32332 35028 32334
rect 35132 32386 35188 32388
rect 35132 32334 35134 32386
rect 35134 32334 35186 32386
rect 35186 32334 35188 32386
rect 35132 32332 35188 32334
rect 35292 32386 35348 32388
rect 35292 32334 35294 32386
rect 35294 32334 35346 32386
rect 35346 32334 35348 32386
rect 35292 32332 35348 32334
rect 35452 32386 35508 32388
rect 35452 32334 35454 32386
rect 35454 32334 35506 32386
rect 35506 32334 35508 32386
rect 35452 32332 35508 32334
rect 35612 32386 35668 32388
rect 35612 32334 35614 32386
rect 35614 32334 35666 32386
rect 35666 32334 35668 32386
rect 35612 32332 35668 32334
rect 35772 32386 35828 32388
rect 35772 32334 35774 32386
rect 35774 32334 35826 32386
rect 35826 32334 35828 32386
rect 35772 32332 35828 32334
rect 35932 32386 35988 32388
rect 35932 32334 35934 32386
rect 35934 32334 35986 32386
rect 35986 32334 35988 32386
rect 35932 32332 35988 32334
rect 36092 32386 36148 32388
rect 36092 32334 36094 32386
rect 36094 32334 36146 32386
rect 36146 32334 36148 32386
rect 36092 32332 36148 32334
rect 36252 32386 36308 32388
rect 36252 32334 36254 32386
rect 36254 32334 36306 32386
rect 36306 32334 36308 32386
rect 36252 32332 36308 32334
rect 36412 32386 36468 32388
rect 36412 32334 36414 32386
rect 36414 32334 36466 32386
rect 36466 32334 36468 32386
rect 36412 32332 36468 32334
rect 36572 32386 36628 32388
rect 36572 32334 36574 32386
rect 36574 32334 36626 32386
rect 36626 32334 36628 32386
rect 36572 32332 36628 32334
rect 36732 32386 36788 32388
rect 36732 32334 36734 32386
rect 36734 32334 36786 32386
rect 36786 32334 36788 32386
rect 36732 32332 36788 32334
rect 36892 32386 36948 32388
rect 36892 32334 36894 32386
rect 36894 32334 36946 32386
rect 36946 32334 36948 32386
rect 36892 32332 36948 32334
rect 37052 32386 37108 32388
rect 37052 32334 37054 32386
rect 37054 32334 37106 32386
rect 37106 32334 37108 32386
rect 37052 32332 37108 32334
rect 37212 32386 37268 32388
rect 37212 32334 37214 32386
rect 37214 32334 37266 32386
rect 37266 32334 37268 32386
rect 37212 32332 37268 32334
rect 37372 32386 37428 32388
rect 37372 32334 37374 32386
rect 37374 32334 37426 32386
rect 37426 32334 37428 32386
rect 37372 32332 37428 32334
rect 37532 32386 37588 32388
rect 37532 32334 37534 32386
rect 37534 32334 37586 32386
rect 37586 32334 37588 32386
rect 37532 32332 37588 32334
rect 37692 32386 37748 32388
rect 37692 32334 37694 32386
rect 37694 32334 37746 32386
rect 37746 32334 37748 32386
rect 37692 32332 37748 32334
rect 37852 32386 37908 32388
rect 37852 32334 37854 32386
rect 37854 32334 37906 32386
rect 37906 32334 37908 32386
rect 37852 32332 37908 32334
rect 38012 32386 38068 32388
rect 38012 32334 38014 32386
rect 38014 32334 38066 32386
rect 38066 32334 38068 32386
rect 38012 32332 38068 32334
rect 38172 32386 38228 32388
rect 38172 32334 38174 32386
rect 38174 32334 38226 32386
rect 38226 32334 38228 32386
rect 38172 32332 38228 32334
rect 38332 32386 38388 32388
rect 38332 32334 38334 32386
rect 38334 32334 38386 32386
rect 38386 32334 38388 32386
rect 38332 32332 38388 32334
rect 38492 32386 38548 32388
rect 38492 32334 38494 32386
rect 38494 32334 38546 32386
rect 38546 32334 38548 32386
rect 38492 32332 38548 32334
rect 38652 32386 38708 32388
rect 38652 32334 38654 32386
rect 38654 32334 38706 32386
rect 38706 32334 38708 32386
rect 38652 32332 38708 32334
rect 38812 32386 38868 32388
rect 38812 32334 38814 32386
rect 38814 32334 38866 32386
rect 38866 32334 38868 32386
rect 38812 32332 38868 32334
rect 38972 32386 39028 32388
rect 38972 32334 38974 32386
rect 38974 32334 39026 32386
rect 39026 32334 39028 32386
rect 38972 32332 39028 32334
rect 39132 32386 39188 32388
rect 39132 32334 39134 32386
rect 39134 32334 39186 32386
rect 39186 32334 39188 32386
rect 39132 32332 39188 32334
rect 39292 32386 39348 32388
rect 39292 32334 39294 32386
rect 39294 32334 39346 32386
rect 39346 32334 39348 32386
rect 39292 32332 39348 32334
rect 39452 32386 39508 32388
rect 39452 32334 39454 32386
rect 39454 32334 39506 32386
rect 39506 32334 39508 32386
rect 39452 32332 39508 32334
rect 39612 32386 39668 32388
rect 39612 32334 39614 32386
rect 39614 32334 39666 32386
rect 39666 32334 39668 32386
rect 39612 32332 39668 32334
rect 39772 32386 39828 32388
rect 39772 32334 39774 32386
rect 39774 32334 39826 32386
rect 39826 32334 39828 32386
rect 39772 32332 39828 32334
rect 39932 32386 39988 32388
rect 39932 32334 39934 32386
rect 39934 32334 39986 32386
rect 39986 32334 39988 32386
rect 39932 32332 39988 32334
rect 40092 32386 40148 32388
rect 40092 32334 40094 32386
rect 40094 32334 40146 32386
rect 40146 32334 40148 32386
rect 40092 32332 40148 32334
rect 40252 32386 40308 32388
rect 40252 32334 40254 32386
rect 40254 32334 40306 32386
rect 40306 32334 40308 32386
rect 40252 32332 40308 32334
rect 40412 32386 40468 32388
rect 40412 32334 40414 32386
rect 40414 32334 40466 32386
rect 40466 32334 40468 32386
rect 40412 32332 40468 32334
rect 40572 32386 40628 32388
rect 40572 32334 40574 32386
rect 40574 32334 40626 32386
rect 40626 32334 40628 32386
rect 40572 32332 40628 32334
rect 40732 32386 40788 32388
rect 40732 32334 40734 32386
rect 40734 32334 40786 32386
rect 40786 32334 40788 32386
rect 40732 32332 40788 32334
rect 40892 32386 40948 32388
rect 40892 32334 40894 32386
rect 40894 32334 40946 32386
rect 40946 32334 40948 32386
rect 40892 32332 40948 32334
rect 41052 32386 41108 32388
rect 41052 32334 41054 32386
rect 41054 32334 41106 32386
rect 41106 32334 41108 32386
rect 41052 32332 41108 32334
rect 41212 32386 41268 32388
rect 41212 32334 41214 32386
rect 41214 32334 41266 32386
rect 41266 32334 41268 32386
rect 41212 32332 41268 32334
rect 41372 32386 41428 32388
rect 41372 32334 41374 32386
rect 41374 32334 41426 32386
rect 41426 32334 41428 32386
rect 41372 32332 41428 32334
rect 41532 32386 41588 32388
rect 41532 32334 41534 32386
rect 41534 32334 41586 32386
rect 41586 32334 41588 32386
rect 41532 32332 41588 32334
rect 41692 32386 41748 32388
rect 41692 32334 41694 32386
rect 41694 32334 41746 32386
rect 41746 32334 41748 32386
rect 41692 32332 41748 32334
rect 41852 32386 41908 32388
rect 41852 32334 41854 32386
rect 41854 32334 41906 32386
rect 41906 32334 41908 32386
rect 41852 32332 41908 32334
rect 9612 32172 9668 32228
rect 20172 32172 20228 32228
rect 32252 32172 32308 32228
rect 12 32066 68 32068
rect 12 32014 14 32066
rect 14 32014 66 32066
rect 66 32014 68 32066
rect 12 32012 68 32014
rect 172 32066 228 32068
rect 172 32014 174 32066
rect 174 32014 226 32066
rect 226 32014 228 32066
rect 172 32012 228 32014
rect 332 32066 388 32068
rect 332 32014 334 32066
rect 334 32014 386 32066
rect 386 32014 388 32066
rect 332 32012 388 32014
rect 492 32066 548 32068
rect 492 32014 494 32066
rect 494 32014 546 32066
rect 546 32014 548 32066
rect 492 32012 548 32014
rect 652 32066 708 32068
rect 652 32014 654 32066
rect 654 32014 706 32066
rect 706 32014 708 32066
rect 652 32012 708 32014
rect 812 32066 868 32068
rect 812 32014 814 32066
rect 814 32014 866 32066
rect 866 32014 868 32066
rect 812 32012 868 32014
rect 972 32066 1028 32068
rect 972 32014 974 32066
rect 974 32014 1026 32066
rect 1026 32014 1028 32066
rect 972 32012 1028 32014
rect 1132 32066 1188 32068
rect 1132 32014 1134 32066
rect 1134 32014 1186 32066
rect 1186 32014 1188 32066
rect 1132 32012 1188 32014
rect 1292 32066 1348 32068
rect 1292 32014 1294 32066
rect 1294 32014 1346 32066
rect 1346 32014 1348 32066
rect 1292 32012 1348 32014
rect 1452 32066 1508 32068
rect 1452 32014 1454 32066
rect 1454 32014 1506 32066
rect 1506 32014 1508 32066
rect 1452 32012 1508 32014
rect 1612 32066 1668 32068
rect 1612 32014 1614 32066
rect 1614 32014 1666 32066
rect 1666 32014 1668 32066
rect 1612 32012 1668 32014
rect 1772 32066 1828 32068
rect 1772 32014 1774 32066
rect 1774 32014 1826 32066
rect 1826 32014 1828 32066
rect 1772 32012 1828 32014
rect 1932 32066 1988 32068
rect 1932 32014 1934 32066
rect 1934 32014 1986 32066
rect 1986 32014 1988 32066
rect 1932 32012 1988 32014
rect 2092 32066 2148 32068
rect 2092 32014 2094 32066
rect 2094 32014 2146 32066
rect 2146 32014 2148 32066
rect 2092 32012 2148 32014
rect 2252 32066 2308 32068
rect 2252 32014 2254 32066
rect 2254 32014 2306 32066
rect 2306 32014 2308 32066
rect 2252 32012 2308 32014
rect 2412 32066 2468 32068
rect 2412 32014 2414 32066
rect 2414 32014 2466 32066
rect 2466 32014 2468 32066
rect 2412 32012 2468 32014
rect 2572 32066 2628 32068
rect 2572 32014 2574 32066
rect 2574 32014 2626 32066
rect 2626 32014 2628 32066
rect 2572 32012 2628 32014
rect 2732 32066 2788 32068
rect 2732 32014 2734 32066
rect 2734 32014 2786 32066
rect 2786 32014 2788 32066
rect 2732 32012 2788 32014
rect 2892 32066 2948 32068
rect 2892 32014 2894 32066
rect 2894 32014 2946 32066
rect 2946 32014 2948 32066
rect 2892 32012 2948 32014
rect 3052 32066 3108 32068
rect 3052 32014 3054 32066
rect 3054 32014 3106 32066
rect 3106 32014 3108 32066
rect 3052 32012 3108 32014
rect 3212 32066 3268 32068
rect 3212 32014 3214 32066
rect 3214 32014 3266 32066
rect 3266 32014 3268 32066
rect 3212 32012 3268 32014
rect 3372 32066 3428 32068
rect 3372 32014 3374 32066
rect 3374 32014 3426 32066
rect 3426 32014 3428 32066
rect 3372 32012 3428 32014
rect 3532 32066 3588 32068
rect 3532 32014 3534 32066
rect 3534 32014 3586 32066
rect 3586 32014 3588 32066
rect 3532 32012 3588 32014
rect 3692 32066 3748 32068
rect 3692 32014 3694 32066
rect 3694 32014 3746 32066
rect 3746 32014 3748 32066
rect 3692 32012 3748 32014
rect 3852 32066 3908 32068
rect 3852 32014 3854 32066
rect 3854 32014 3906 32066
rect 3906 32014 3908 32066
rect 3852 32012 3908 32014
rect 4012 32066 4068 32068
rect 4012 32014 4014 32066
rect 4014 32014 4066 32066
rect 4066 32014 4068 32066
rect 4012 32012 4068 32014
rect 4172 32066 4228 32068
rect 4172 32014 4174 32066
rect 4174 32014 4226 32066
rect 4226 32014 4228 32066
rect 4172 32012 4228 32014
rect 4332 32066 4388 32068
rect 4332 32014 4334 32066
rect 4334 32014 4386 32066
rect 4386 32014 4388 32066
rect 4332 32012 4388 32014
rect 4492 32066 4548 32068
rect 4492 32014 4494 32066
rect 4494 32014 4546 32066
rect 4546 32014 4548 32066
rect 4492 32012 4548 32014
rect 4652 32066 4708 32068
rect 4652 32014 4654 32066
rect 4654 32014 4706 32066
rect 4706 32014 4708 32066
rect 4652 32012 4708 32014
rect 4812 32066 4868 32068
rect 4812 32014 4814 32066
rect 4814 32014 4866 32066
rect 4866 32014 4868 32066
rect 4812 32012 4868 32014
rect 4972 32066 5028 32068
rect 4972 32014 4974 32066
rect 4974 32014 5026 32066
rect 5026 32014 5028 32066
rect 4972 32012 5028 32014
rect 5132 32066 5188 32068
rect 5132 32014 5134 32066
rect 5134 32014 5186 32066
rect 5186 32014 5188 32066
rect 5132 32012 5188 32014
rect 5292 32066 5348 32068
rect 5292 32014 5294 32066
rect 5294 32014 5346 32066
rect 5346 32014 5348 32066
rect 5292 32012 5348 32014
rect 5452 32066 5508 32068
rect 5452 32014 5454 32066
rect 5454 32014 5506 32066
rect 5506 32014 5508 32066
rect 5452 32012 5508 32014
rect 5612 32066 5668 32068
rect 5612 32014 5614 32066
rect 5614 32014 5666 32066
rect 5666 32014 5668 32066
rect 5612 32012 5668 32014
rect 5772 32066 5828 32068
rect 5772 32014 5774 32066
rect 5774 32014 5826 32066
rect 5826 32014 5828 32066
rect 5772 32012 5828 32014
rect 5932 32066 5988 32068
rect 5932 32014 5934 32066
rect 5934 32014 5986 32066
rect 5986 32014 5988 32066
rect 5932 32012 5988 32014
rect 6092 32066 6148 32068
rect 6092 32014 6094 32066
rect 6094 32014 6146 32066
rect 6146 32014 6148 32066
rect 6092 32012 6148 32014
rect 6252 32066 6308 32068
rect 6252 32014 6254 32066
rect 6254 32014 6306 32066
rect 6306 32014 6308 32066
rect 6252 32012 6308 32014
rect 6412 32066 6468 32068
rect 6412 32014 6414 32066
rect 6414 32014 6466 32066
rect 6466 32014 6468 32066
rect 6412 32012 6468 32014
rect 6572 32066 6628 32068
rect 6572 32014 6574 32066
rect 6574 32014 6626 32066
rect 6626 32014 6628 32066
rect 6572 32012 6628 32014
rect 6732 32066 6788 32068
rect 6732 32014 6734 32066
rect 6734 32014 6786 32066
rect 6786 32014 6788 32066
rect 6732 32012 6788 32014
rect 6892 32066 6948 32068
rect 6892 32014 6894 32066
rect 6894 32014 6946 32066
rect 6946 32014 6948 32066
rect 6892 32012 6948 32014
rect 7052 32066 7108 32068
rect 7052 32014 7054 32066
rect 7054 32014 7106 32066
rect 7106 32014 7108 32066
rect 7052 32012 7108 32014
rect 7212 32066 7268 32068
rect 7212 32014 7214 32066
rect 7214 32014 7266 32066
rect 7266 32014 7268 32066
rect 7212 32012 7268 32014
rect 7372 32066 7428 32068
rect 7372 32014 7374 32066
rect 7374 32014 7426 32066
rect 7426 32014 7428 32066
rect 7372 32012 7428 32014
rect 7532 32066 7588 32068
rect 7532 32014 7534 32066
rect 7534 32014 7586 32066
rect 7586 32014 7588 32066
rect 7532 32012 7588 32014
rect 7692 32066 7748 32068
rect 7692 32014 7694 32066
rect 7694 32014 7746 32066
rect 7746 32014 7748 32066
rect 7692 32012 7748 32014
rect 7852 32066 7908 32068
rect 7852 32014 7854 32066
rect 7854 32014 7906 32066
rect 7906 32014 7908 32066
rect 7852 32012 7908 32014
rect 8012 32066 8068 32068
rect 8012 32014 8014 32066
rect 8014 32014 8066 32066
rect 8066 32014 8068 32066
rect 8012 32012 8068 32014
rect 8172 32066 8228 32068
rect 8172 32014 8174 32066
rect 8174 32014 8226 32066
rect 8226 32014 8228 32066
rect 8172 32012 8228 32014
rect 8332 32066 8388 32068
rect 8332 32014 8334 32066
rect 8334 32014 8386 32066
rect 8386 32014 8388 32066
rect 8332 32012 8388 32014
rect 9452 32012 9508 32068
rect 9772 32012 9828 32068
rect 10092 32012 10148 32068
rect 10412 32012 10468 32068
rect 10732 32012 10788 32068
rect 11052 32012 11108 32068
rect 11372 32012 11428 32068
rect 12492 32066 12548 32068
rect 12492 32014 12494 32066
rect 12494 32014 12546 32066
rect 12546 32014 12548 32066
rect 12492 32012 12548 32014
rect 12652 32066 12708 32068
rect 12652 32014 12654 32066
rect 12654 32014 12706 32066
rect 12706 32014 12708 32066
rect 12652 32012 12708 32014
rect 12812 32066 12868 32068
rect 12812 32014 12814 32066
rect 12814 32014 12866 32066
rect 12866 32014 12868 32066
rect 12812 32012 12868 32014
rect 12972 32066 13028 32068
rect 12972 32014 12974 32066
rect 12974 32014 13026 32066
rect 13026 32014 13028 32066
rect 12972 32012 13028 32014
rect 13132 32066 13188 32068
rect 13132 32014 13134 32066
rect 13134 32014 13186 32066
rect 13186 32014 13188 32066
rect 13132 32012 13188 32014
rect 13292 32066 13348 32068
rect 13292 32014 13294 32066
rect 13294 32014 13346 32066
rect 13346 32014 13348 32066
rect 13292 32012 13348 32014
rect 13452 32066 13508 32068
rect 13452 32014 13454 32066
rect 13454 32014 13506 32066
rect 13506 32014 13508 32066
rect 13452 32012 13508 32014
rect 13612 32066 13668 32068
rect 13612 32014 13614 32066
rect 13614 32014 13666 32066
rect 13666 32014 13668 32066
rect 13612 32012 13668 32014
rect 13772 32066 13828 32068
rect 13772 32014 13774 32066
rect 13774 32014 13826 32066
rect 13826 32014 13828 32066
rect 13772 32012 13828 32014
rect 13932 32066 13988 32068
rect 13932 32014 13934 32066
rect 13934 32014 13986 32066
rect 13986 32014 13988 32066
rect 13932 32012 13988 32014
rect 14092 32066 14148 32068
rect 14092 32014 14094 32066
rect 14094 32014 14146 32066
rect 14146 32014 14148 32066
rect 14092 32012 14148 32014
rect 14252 32066 14308 32068
rect 14252 32014 14254 32066
rect 14254 32014 14306 32066
rect 14306 32014 14308 32066
rect 14252 32012 14308 32014
rect 14412 32066 14468 32068
rect 14412 32014 14414 32066
rect 14414 32014 14466 32066
rect 14466 32014 14468 32066
rect 14412 32012 14468 32014
rect 14572 32066 14628 32068
rect 14572 32014 14574 32066
rect 14574 32014 14626 32066
rect 14626 32014 14628 32066
rect 14572 32012 14628 32014
rect 14732 32066 14788 32068
rect 14732 32014 14734 32066
rect 14734 32014 14786 32066
rect 14786 32014 14788 32066
rect 14732 32012 14788 32014
rect 14892 32066 14948 32068
rect 14892 32014 14894 32066
rect 14894 32014 14946 32066
rect 14946 32014 14948 32066
rect 14892 32012 14948 32014
rect 15052 32066 15108 32068
rect 15052 32014 15054 32066
rect 15054 32014 15106 32066
rect 15106 32014 15108 32066
rect 15052 32012 15108 32014
rect 15212 32066 15268 32068
rect 15212 32014 15214 32066
rect 15214 32014 15266 32066
rect 15266 32014 15268 32066
rect 15212 32012 15268 32014
rect 15372 32066 15428 32068
rect 15372 32014 15374 32066
rect 15374 32014 15426 32066
rect 15426 32014 15428 32066
rect 15372 32012 15428 32014
rect 15532 32066 15588 32068
rect 15532 32014 15534 32066
rect 15534 32014 15586 32066
rect 15586 32014 15588 32066
rect 15532 32012 15588 32014
rect 15692 32066 15748 32068
rect 15692 32014 15694 32066
rect 15694 32014 15746 32066
rect 15746 32014 15748 32066
rect 15692 32012 15748 32014
rect 15852 32066 15908 32068
rect 15852 32014 15854 32066
rect 15854 32014 15906 32066
rect 15906 32014 15908 32066
rect 15852 32012 15908 32014
rect 16012 32066 16068 32068
rect 16012 32014 16014 32066
rect 16014 32014 16066 32066
rect 16066 32014 16068 32066
rect 16012 32012 16068 32014
rect 16172 32066 16228 32068
rect 16172 32014 16174 32066
rect 16174 32014 16226 32066
rect 16226 32014 16228 32066
rect 16172 32012 16228 32014
rect 16332 32066 16388 32068
rect 16332 32014 16334 32066
rect 16334 32014 16386 32066
rect 16386 32014 16388 32066
rect 16332 32012 16388 32014
rect 16492 32066 16548 32068
rect 16492 32014 16494 32066
rect 16494 32014 16546 32066
rect 16546 32014 16548 32066
rect 16492 32012 16548 32014
rect 16652 32066 16708 32068
rect 16652 32014 16654 32066
rect 16654 32014 16706 32066
rect 16706 32014 16708 32066
rect 16652 32012 16708 32014
rect 16812 32066 16868 32068
rect 16812 32014 16814 32066
rect 16814 32014 16866 32066
rect 16866 32014 16868 32066
rect 16812 32012 16868 32014
rect 16972 32066 17028 32068
rect 16972 32014 16974 32066
rect 16974 32014 17026 32066
rect 17026 32014 17028 32066
rect 16972 32012 17028 32014
rect 17132 32066 17188 32068
rect 17132 32014 17134 32066
rect 17134 32014 17186 32066
rect 17186 32014 17188 32066
rect 17132 32012 17188 32014
rect 17292 32066 17348 32068
rect 17292 32014 17294 32066
rect 17294 32014 17346 32066
rect 17346 32014 17348 32066
rect 17292 32012 17348 32014
rect 17452 32066 17508 32068
rect 17452 32014 17454 32066
rect 17454 32014 17506 32066
rect 17506 32014 17508 32066
rect 17452 32012 17508 32014
rect 17612 32066 17668 32068
rect 17612 32014 17614 32066
rect 17614 32014 17666 32066
rect 17666 32014 17668 32066
rect 17612 32012 17668 32014
rect 17772 32066 17828 32068
rect 17772 32014 17774 32066
rect 17774 32014 17826 32066
rect 17826 32014 17828 32066
rect 17772 32012 17828 32014
rect 17932 32066 17988 32068
rect 17932 32014 17934 32066
rect 17934 32014 17986 32066
rect 17986 32014 17988 32066
rect 17932 32012 17988 32014
rect 18092 32066 18148 32068
rect 18092 32014 18094 32066
rect 18094 32014 18146 32066
rect 18146 32014 18148 32066
rect 18092 32012 18148 32014
rect 18252 32066 18308 32068
rect 18252 32014 18254 32066
rect 18254 32014 18306 32066
rect 18306 32014 18308 32066
rect 18252 32012 18308 32014
rect 18412 32066 18468 32068
rect 18412 32014 18414 32066
rect 18414 32014 18466 32066
rect 18466 32014 18468 32066
rect 18412 32012 18468 32014
rect 18572 32066 18628 32068
rect 18572 32014 18574 32066
rect 18574 32014 18626 32066
rect 18626 32014 18628 32066
rect 18572 32012 18628 32014
rect 18732 32066 18788 32068
rect 18732 32014 18734 32066
rect 18734 32014 18786 32066
rect 18786 32014 18788 32066
rect 18732 32012 18788 32014
rect 18892 32066 18948 32068
rect 18892 32014 18894 32066
rect 18894 32014 18946 32066
rect 18946 32014 18948 32066
rect 18892 32012 18948 32014
rect 20012 32012 20068 32068
rect 20332 32012 20388 32068
rect 20652 32012 20708 32068
rect 20972 32012 21028 32068
rect 21292 32012 21348 32068
rect 21612 32012 21668 32068
rect 21932 32012 21988 32068
rect 23132 32066 23188 32068
rect 23132 32014 23134 32066
rect 23134 32014 23186 32066
rect 23186 32014 23188 32066
rect 23132 32012 23188 32014
rect 23292 32066 23348 32068
rect 23292 32014 23294 32066
rect 23294 32014 23346 32066
rect 23346 32014 23348 32066
rect 23292 32012 23348 32014
rect 23452 32066 23508 32068
rect 23452 32014 23454 32066
rect 23454 32014 23506 32066
rect 23506 32014 23508 32066
rect 23452 32012 23508 32014
rect 23612 32066 23668 32068
rect 23612 32014 23614 32066
rect 23614 32014 23666 32066
rect 23666 32014 23668 32066
rect 23612 32012 23668 32014
rect 23772 32066 23828 32068
rect 23772 32014 23774 32066
rect 23774 32014 23826 32066
rect 23826 32014 23828 32066
rect 23772 32012 23828 32014
rect 23932 32066 23988 32068
rect 23932 32014 23934 32066
rect 23934 32014 23986 32066
rect 23986 32014 23988 32066
rect 23932 32012 23988 32014
rect 24092 32066 24148 32068
rect 24092 32014 24094 32066
rect 24094 32014 24146 32066
rect 24146 32014 24148 32066
rect 24092 32012 24148 32014
rect 24252 32066 24308 32068
rect 24252 32014 24254 32066
rect 24254 32014 24306 32066
rect 24306 32014 24308 32066
rect 24252 32012 24308 32014
rect 24412 32066 24468 32068
rect 24412 32014 24414 32066
rect 24414 32014 24466 32066
rect 24466 32014 24468 32066
rect 24412 32012 24468 32014
rect 24572 32066 24628 32068
rect 24572 32014 24574 32066
rect 24574 32014 24626 32066
rect 24626 32014 24628 32066
rect 24572 32012 24628 32014
rect 24732 32066 24788 32068
rect 24732 32014 24734 32066
rect 24734 32014 24786 32066
rect 24786 32014 24788 32066
rect 24732 32012 24788 32014
rect 24892 32066 24948 32068
rect 24892 32014 24894 32066
rect 24894 32014 24946 32066
rect 24946 32014 24948 32066
rect 24892 32012 24948 32014
rect 25052 32066 25108 32068
rect 25052 32014 25054 32066
rect 25054 32014 25106 32066
rect 25106 32014 25108 32066
rect 25052 32012 25108 32014
rect 25212 32066 25268 32068
rect 25212 32014 25214 32066
rect 25214 32014 25266 32066
rect 25266 32014 25268 32066
rect 25212 32012 25268 32014
rect 25372 32066 25428 32068
rect 25372 32014 25374 32066
rect 25374 32014 25426 32066
rect 25426 32014 25428 32066
rect 25372 32012 25428 32014
rect 25532 32066 25588 32068
rect 25532 32014 25534 32066
rect 25534 32014 25586 32066
rect 25586 32014 25588 32066
rect 25532 32012 25588 32014
rect 25692 32066 25748 32068
rect 25692 32014 25694 32066
rect 25694 32014 25746 32066
rect 25746 32014 25748 32066
rect 25692 32012 25748 32014
rect 25852 32066 25908 32068
rect 25852 32014 25854 32066
rect 25854 32014 25906 32066
rect 25906 32014 25908 32066
rect 25852 32012 25908 32014
rect 26012 32066 26068 32068
rect 26012 32014 26014 32066
rect 26014 32014 26066 32066
rect 26066 32014 26068 32066
rect 26012 32012 26068 32014
rect 26172 32066 26228 32068
rect 26172 32014 26174 32066
rect 26174 32014 26226 32066
rect 26226 32014 26228 32066
rect 26172 32012 26228 32014
rect 26332 32066 26388 32068
rect 26332 32014 26334 32066
rect 26334 32014 26386 32066
rect 26386 32014 26388 32066
rect 26332 32012 26388 32014
rect 26492 32066 26548 32068
rect 26492 32014 26494 32066
rect 26494 32014 26546 32066
rect 26546 32014 26548 32066
rect 26492 32012 26548 32014
rect 26652 32066 26708 32068
rect 26652 32014 26654 32066
rect 26654 32014 26706 32066
rect 26706 32014 26708 32066
rect 26652 32012 26708 32014
rect 26812 32066 26868 32068
rect 26812 32014 26814 32066
rect 26814 32014 26866 32066
rect 26866 32014 26868 32066
rect 26812 32012 26868 32014
rect 26972 32066 27028 32068
rect 26972 32014 26974 32066
rect 26974 32014 27026 32066
rect 27026 32014 27028 32066
rect 26972 32012 27028 32014
rect 27132 32066 27188 32068
rect 27132 32014 27134 32066
rect 27134 32014 27186 32066
rect 27186 32014 27188 32066
rect 27132 32012 27188 32014
rect 27292 32066 27348 32068
rect 27292 32014 27294 32066
rect 27294 32014 27346 32066
rect 27346 32014 27348 32066
rect 27292 32012 27348 32014
rect 27452 32066 27508 32068
rect 27452 32014 27454 32066
rect 27454 32014 27506 32066
rect 27506 32014 27508 32066
rect 27452 32012 27508 32014
rect 27612 32066 27668 32068
rect 27612 32014 27614 32066
rect 27614 32014 27666 32066
rect 27666 32014 27668 32066
rect 27612 32012 27668 32014
rect 27772 32066 27828 32068
rect 27772 32014 27774 32066
rect 27774 32014 27826 32066
rect 27826 32014 27828 32066
rect 27772 32012 27828 32014
rect 27932 32066 27988 32068
rect 27932 32014 27934 32066
rect 27934 32014 27986 32066
rect 27986 32014 27988 32066
rect 27932 32012 27988 32014
rect 28092 32066 28148 32068
rect 28092 32014 28094 32066
rect 28094 32014 28146 32066
rect 28146 32014 28148 32066
rect 28092 32012 28148 32014
rect 28252 32066 28308 32068
rect 28252 32014 28254 32066
rect 28254 32014 28306 32066
rect 28306 32014 28308 32066
rect 28252 32012 28308 32014
rect 28412 32066 28468 32068
rect 28412 32014 28414 32066
rect 28414 32014 28466 32066
rect 28466 32014 28468 32066
rect 28412 32012 28468 32014
rect 28572 32066 28628 32068
rect 28572 32014 28574 32066
rect 28574 32014 28626 32066
rect 28626 32014 28628 32066
rect 28572 32012 28628 32014
rect 28732 32066 28788 32068
rect 28732 32014 28734 32066
rect 28734 32014 28786 32066
rect 28786 32014 28788 32066
rect 28732 32012 28788 32014
rect 28892 32066 28948 32068
rect 28892 32014 28894 32066
rect 28894 32014 28946 32066
rect 28946 32014 28948 32066
rect 28892 32012 28948 32014
rect 29052 32066 29108 32068
rect 29052 32014 29054 32066
rect 29054 32014 29106 32066
rect 29106 32014 29108 32066
rect 29052 32012 29108 32014
rect 29212 32066 29268 32068
rect 29212 32014 29214 32066
rect 29214 32014 29266 32066
rect 29266 32014 29268 32066
rect 29212 32012 29268 32014
rect 29372 32066 29428 32068
rect 29372 32014 29374 32066
rect 29374 32014 29426 32066
rect 29426 32014 29428 32066
rect 29372 32012 29428 32014
rect 30492 32012 30548 32068
rect 30812 32012 30868 32068
rect 31132 32012 31188 32068
rect 31452 32012 31508 32068
rect 31772 32012 31828 32068
rect 32092 32012 32148 32068
rect 32412 32012 32468 32068
rect 33532 32066 33588 32068
rect 33532 32014 33534 32066
rect 33534 32014 33586 32066
rect 33586 32014 33588 32066
rect 33532 32012 33588 32014
rect 33692 32066 33748 32068
rect 33692 32014 33694 32066
rect 33694 32014 33746 32066
rect 33746 32014 33748 32066
rect 33692 32012 33748 32014
rect 33852 32066 33908 32068
rect 33852 32014 33854 32066
rect 33854 32014 33906 32066
rect 33906 32014 33908 32066
rect 33852 32012 33908 32014
rect 34012 32066 34068 32068
rect 34012 32014 34014 32066
rect 34014 32014 34066 32066
rect 34066 32014 34068 32066
rect 34012 32012 34068 32014
rect 34172 32066 34228 32068
rect 34172 32014 34174 32066
rect 34174 32014 34226 32066
rect 34226 32014 34228 32066
rect 34172 32012 34228 32014
rect 34332 32066 34388 32068
rect 34332 32014 34334 32066
rect 34334 32014 34386 32066
rect 34386 32014 34388 32066
rect 34332 32012 34388 32014
rect 34492 32066 34548 32068
rect 34492 32014 34494 32066
rect 34494 32014 34546 32066
rect 34546 32014 34548 32066
rect 34492 32012 34548 32014
rect 34652 32066 34708 32068
rect 34652 32014 34654 32066
rect 34654 32014 34706 32066
rect 34706 32014 34708 32066
rect 34652 32012 34708 32014
rect 34812 32066 34868 32068
rect 34812 32014 34814 32066
rect 34814 32014 34866 32066
rect 34866 32014 34868 32066
rect 34812 32012 34868 32014
rect 34972 32066 35028 32068
rect 34972 32014 34974 32066
rect 34974 32014 35026 32066
rect 35026 32014 35028 32066
rect 34972 32012 35028 32014
rect 35132 32066 35188 32068
rect 35132 32014 35134 32066
rect 35134 32014 35186 32066
rect 35186 32014 35188 32066
rect 35132 32012 35188 32014
rect 35292 32066 35348 32068
rect 35292 32014 35294 32066
rect 35294 32014 35346 32066
rect 35346 32014 35348 32066
rect 35292 32012 35348 32014
rect 35452 32066 35508 32068
rect 35452 32014 35454 32066
rect 35454 32014 35506 32066
rect 35506 32014 35508 32066
rect 35452 32012 35508 32014
rect 35612 32066 35668 32068
rect 35612 32014 35614 32066
rect 35614 32014 35666 32066
rect 35666 32014 35668 32066
rect 35612 32012 35668 32014
rect 35772 32066 35828 32068
rect 35772 32014 35774 32066
rect 35774 32014 35826 32066
rect 35826 32014 35828 32066
rect 35772 32012 35828 32014
rect 35932 32066 35988 32068
rect 35932 32014 35934 32066
rect 35934 32014 35986 32066
rect 35986 32014 35988 32066
rect 35932 32012 35988 32014
rect 36092 32066 36148 32068
rect 36092 32014 36094 32066
rect 36094 32014 36146 32066
rect 36146 32014 36148 32066
rect 36092 32012 36148 32014
rect 36252 32066 36308 32068
rect 36252 32014 36254 32066
rect 36254 32014 36306 32066
rect 36306 32014 36308 32066
rect 36252 32012 36308 32014
rect 36412 32066 36468 32068
rect 36412 32014 36414 32066
rect 36414 32014 36466 32066
rect 36466 32014 36468 32066
rect 36412 32012 36468 32014
rect 36572 32066 36628 32068
rect 36572 32014 36574 32066
rect 36574 32014 36626 32066
rect 36626 32014 36628 32066
rect 36572 32012 36628 32014
rect 36732 32066 36788 32068
rect 36732 32014 36734 32066
rect 36734 32014 36786 32066
rect 36786 32014 36788 32066
rect 36732 32012 36788 32014
rect 36892 32066 36948 32068
rect 36892 32014 36894 32066
rect 36894 32014 36946 32066
rect 36946 32014 36948 32066
rect 36892 32012 36948 32014
rect 37052 32066 37108 32068
rect 37052 32014 37054 32066
rect 37054 32014 37106 32066
rect 37106 32014 37108 32066
rect 37052 32012 37108 32014
rect 37212 32066 37268 32068
rect 37212 32014 37214 32066
rect 37214 32014 37266 32066
rect 37266 32014 37268 32066
rect 37212 32012 37268 32014
rect 37372 32066 37428 32068
rect 37372 32014 37374 32066
rect 37374 32014 37426 32066
rect 37426 32014 37428 32066
rect 37372 32012 37428 32014
rect 37532 32066 37588 32068
rect 37532 32014 37534 32066
rect 37534 32014 37586 32066
rect 37586 32014 37588 32066
rect 37532 32012 37588 32014
rect 37692 32066 37748 32068
rect 37692 32014 37694 32066
rect 37694 32014 37746 32066
rect 37746 32014 37748 32066
rect 37692 32012 37748 32014
rect 37852 32066 37908 32068
rect 37852 32014 37854 32066
rect 37854 32014 37906 32066
rect 37906 32014 37908 32066
rect 37852 32012 37908 32014
rect 38012 32066 38068 32068
rect 38012 32014 38014 32066
rect 38014 32014 38066 32066
rect 38066 32014 38068 32066
rect 38012 32012 38068 32014
rect 38172 32066 38228 32068
rect 38172 32014 38174 32066
rect 38174 32014 38226 32066
rect 38226 32014 38228 32066
rect 38172 32012 38228 32014
rect 38332 32066 38388 32068
rect 38332 32014 38334 32066
rect 38334 32014 38386 32066
rect 38386 32014 38388 32066
rect 38332 32012 38388 32014
rect 38492 32066 38548 32068
rect 38492 32014 38494 32066
rect 38494 32014 38546 32066
rect 38546 32014 38548 32066
rect 38492 32012 38548 32014
rect 38652 32066 38708 32068
rect 38652 32014 38654 32066
rect 38654 32014 38706 32066
rect 38706 32014 38708 32066
rect 38652 32012 38708 32014
rect 38812 32066 38868 32068
rect 38812 32014 38814 32066
rect 38814 32014 38866 32066
rect 38866 32014 38868 32066
rect 38812 32012 38868 32014
rect 38972 32066 39028 32068
rect 38972 32014 38974 32066
rect 38974 32014 39026 32066
rect 39026 32014 39028 32066
rect 38972 32012 39028 32014
rect 39132 32066 39188 32068
rect 39132 32014 39134 32066
rect 39134 32014 39186 32066
rect 39186 32014 39188 32066
rect 39132 32012 39188 32014
rect 39292 32066 39348 32068
rect 39292 32014 39294 32066
rect 39294 32014 39346 32066
rect 39346 32014 39348 32066
rect 39292 32012 39348 32014
rect 39452 32066 39508 32068
rect 39452 32014 39454 32066
rect 39454 32014 39506 32066
rect 39506 32014 39508 32066
rect 39452 32012 39508 32014
rect 39612 32066 39668 32068
rect 39612 32014 39614 32066
rect 39614 32014 39666 32066
rect 39666 32014 39668 32066
rect 39612 32012 39668 32014
rect 39772 32066 39828 32068
rect 39772 32014 39774 32066
rect 39774 32014 39826 32066
rect 39826 32014 39828 32066
rect 39772 32012 39828 32014
rect 39932 32066 39988 32068
rect 39932 32014 39934 32066
rect 39934 32014 39986 32066
rect 39986 32014 39988 32066
rect 39932 32012 39988 32014
rect 40092 32066 40148 32068
rect 40092 32014 40094 32066
rect 40094 32014 40146 32066
rect 40146 32014 40148 32066
rect 40092 32012 40148 32014
rect 40252 32066 40308 32068
rect 40252 32014 40254 32066
rect 40254 32014 40306 32066
rect 40306 32014 40308 32066
rect 40252 32012 40308 32014
rect 40412 32066 40468 32068
rect 40412 32014 40414 32066
rect 40414 32014 40466 32066
rect 40466 32014 40468 32066
rect 40412 32012 40468 32014
rect 40572 32066 40628 32068
rect 40572 32014 40574 32066
rect 40574 32014 40626 32066
rect 40626 32014 40628 32066
rect 40572 32012 40628 32014
rect 40732 32066 40788 32068
rect 40732 32014 40734 32066
rect 40734 32014 40786 32066
rect 40786 32014 40788 32066
rect 40732 32012 40788 32014
rect 40892 32066 40948 32068
rect 40892 32014 40894 32066
rect 40894 32014 40946 32066
rect 40946 32014 40948 32066
rect 40892 32012 40948 32014
rect 41052 32066 41108 32068
rect 41052 32014 41054 32066
rect 41054 32014 41106 32066
rect 41106 32014 41108 32066
rect 41052 32012 41108 32014
rect 41212 32066 41268 32068
rect 41212 32014 41214 32066
rect 41214 32014 41266 32066
rect 41266 32014 41268 32066
rect 41212 32012 41268 32014
rect 41372 32066 41428 32068
rect 41372 32014 41374 32066
rect 41374 32014 41426 32066
rect 41426 32014 41428 32066
rect 41372 32012 41428 32014
rect 41532 32066 41588 32068
rect 41532 32014 41534 32066
rect 41534 32014 41586 32066
rect 41586 32014 41588 32066
rect 41532 32012 41588 32014
rect 41692 32066 41748 32068
rect 41692 32014 41694 32066
rect 41694 32014 41746 32066
rect 41746 32014 41748 32066
rect 41692 32012 41748 32014
rect 41852 32066 41908 32068
rect 41852 32014 41854 32066
rect 41854 32014 41906 32066
rect 41906 32014 41908 32066
rect 41852 32012 41908 32014
rect 9932 31852 9988 31908
rect 20492 31852 20548 31908
rect 31932 31852 31988 31908
rect 12 31746 68 31748
rect 12 31694 14 31746
rect 14 31694 66 31746
rect 66 31694 68 31746
rect 12 31692 68 31694
rect 172 31746 228 31748
rect 172 31694 174 31746
rect 174 31694 226 31746
rect 226 31694 228 31746
rect 172 31692 228 31694
rect 332 31746 388 31748
rect 332 31694 334 31746
rect 334 31694 386 31746
rect 386 31694 388 31746
rect 332 31692 388 31694
rect 492 31746 548 31748
rect 492 31694 494 31746
rect 494 31694 546 31746
rect 546 31694 548 31746
rect 492 31692 548 31694
rect 652 31746 708 31748
rect 652 31694 654 31746
rect 654 31694 706 31746
rect 706 31694 708 31746
rect 652 31692 708 31694
rect 812 31746 868 31748
rect 812 31694 814 31746
rect 814 31694 866 31746
rect 866 31694 868 31746
rect 812 31692 868 31694
rect 972 31746 1028 31748
rect 972 31694 974 31746
rect 974 31694 1026 31746
rect 1026 31694 1028 31746
rect 972 31692 1028 31694
rect 1132 31746 1188 31748
rect 1132 31694 1134 31746
rect 1134 31694 1186 31746
rect 1186 31694 1188 31746
rect 1132 31692 1188 31694
rect 1292 31746 1348 31748
rect 1292 31694 1294 31746
rect 1294 31694 1346 31746
rect 1346 31694 1348 31746
rect 1292 31692 1348 31694
rect 1452 31746 1508 31748
rect 1452 31694 1454 31746
rect 1454 31694 1506 31746
rect 1506 31694 1508 31746
rect 1452 31692 1508 31694
rect 1612 31746 1668 31748
rect 1612 31694 1614 31746
rect 1614 31694 1666 31746
rect 1666 31694 1668 31746
rect 1612 31692 1668 31694
rect 1772 31746 1828 31748
rect 1772 31694 1774 31746
rect 1774 31694 1826 31746
rect 1826 31694 1828 31746
rect 1772 31692 1828 31694
rect 1932 31746 1988 31748
rect 1932 31694 1934 31746
rect 1934 31694 1986 31746
rect 1986 31694 1988 31746
rect 1932 31692 1988 31694
rect 2092 31746 2148 31748
rect 2092 31694 2094 31746
rect 2094 31694 2146 31746
rect 2146 31694 2148 31746
rect 2092 31692 2148 31694
rect 2252 31746 2308 31748
rect 2252 31694 2254 31746
rect 2254 31694 2306 31746
rect 2306 31694 2308 31746
rect 2252 31692 2308 31694
rect 2412 31746 2468 31748
rect 2412 31694 2414 31746
rect 2414 31694 2466 31746
rect 2466 31694 2468 31746
rect 2412 31692 2468 31694
rect 2572 31746 2628 31748
rect 2572 31694 2574 31746
rect 2574 31694 2626 31746
rect 2626 31694 2628 31746
rect 2572 31692 2628 31694
rect 2732 31746 2788 31748
rect 2732 31694 2734 31746
rect 2734 31694 2786 31746
rect 2786 31694 2788 31746
rect 2732 31692 2788 31694
rect 2892 31746 2948 31748
rect 2892 31694 2894 31746
rect 2894 31694 2946 31746
rect 2946 31694 2948 31746
rect 2892 31692 2948 31694
rect 3052 31746 3108 31748
rect 3052 31694 3054 31746
rect 3054 31694 3106 31746
rect 3106 31694 3108 31746
rect 3052 31692 3108 31694
rect 3212 31746 3268 31748
rect 3212 31694 3214 31746
rect 3214 31694 3266 31746
rect 3266 31694 3268 31746
rect 3212 31692 3268 31694
rect 3372 31746 3428 31748
rect 3372 31694 3374 31746
rect 3374 31694 3426 31746
rect 3426 31694 3428 31746
rect 3372 31692 3428 31694
rect 3532 31746 3588 31748
rect 3532 31694 3534 31746
rect 3534 31694 3586 31746
rect 3586 31694 3588 31746
rect 3532 31692 3588 31694
rect 3692 31746 3748 31748
rect 3692 31694 3694 31746
rect 3694 31694 3746 31746
rect 3746 31694 3748 31746
rect 3692 31692 3748 31694
rect 3852 31746 3908 31748
rect 3852 31694 3854 31746
rect 3854 31694 3906 31746
rect 3906 31694 3908 31746
rect 3852 31692 3908 31694
rect 4012 31746 4068 31748
rect 4012 31694 4014 31746
rect 4014 31694 4066 31746
rect 4066 31694 4068 31746
rect 4012 31692 4068 31694
rect 4172 31746 4228 31748
rect 4172 31694 4174 31746
rect 4174 31694 4226 31746
rect 4226 31694 4228 31746
rect 4172 31692 4228 31694
rect 4332 31746 4388 31748
rect 4332 31694 4334 31746
rect 4334 31694 4386 31746
rect 4386 31694 4388 31746
rect 4332 31692 4388 31694
rect 4492 31746 4548 31748
rect 4492 31694 4494 31746
rect 4494 31694 4546 31746
rect 4546 31694 4548 31746
rect 4492 31692 4548 31694
rect 4652 31746 4708 31748
rect 4652 31694 4654 31746
rect 4654 31694 4706 31746
rect 4706 31694 4708 31746
rect 4652 31692 4708 31694
rect 4812 31746 4868 31748
rect 4812 31694 4814 31746
rect 4814 31694 4866 31746
rect 4866 31694 4868 31746
rect 4812 31692 4868 31694
rect 4972 31746 5028 31748
rect 4972 31694 4974 31746
rect 4974 31694 5026 31746
rect 5026 31694 5028 31746
rect 4972 31692 5028 31694
rect 5132 31746 5188 31748
rect 5132 31694 5134 31746
rect 5134 31694 5186 31746
rect 5186 31694 5188 31746
rect 5132 31692 5188 31694
rect 5292 31746 5348 31748
rect 5292 31694 5294 31746
rect 5294 31694 5346 31746
rect 5346 31694 5348 31746
rect 5292 31692 5348 31694
rect 5452 31746 5508 31748
rect 5452 31694 5454 31746
rect 5454 31694 5506 31746
rect 5506 31694 5508 31746
rect 5452 31692 5508 31694
rect 5612 31746 5668 31748
rect 5612 31694 5614 31746
rect 5614 31694 5666 31746
rect 5666 31694 5668 31746
rect 5612 31692 5668 31694
rect 5772 31746 5828 31748
rect 5772 31694 5774 31746
rect 5774 31694 5826 31746
rect 5826 31694 5828 31746
rect 5772 31692 5828 31694
rect 5932 31746 5988 31748
rect 5932 31694 5934 31746
rect 5934 31694 5986 31746
rect 5986 31694 5988 31746
rect 5932 31692 5988 31694
rect 6092 31746 6148 31748
rect 6092 31694 6094 31746
rect 6094 31694 6146 31746
rect 6146 31694 6148 31746
rect 6092 31692 6148 31694
rect 6252 31746 6308 31748
rect 6252 31694 6254 31746
rect 6254 31694 6306 31746
rect 6306 31694 6308 31746
rect 6252 31692 6308 31694
rect 6412 31746 6468 31748
rect 6412 31694 6414 31746
rect 6414 31694 6466 31746
rect 6466 31694 6468 31746
rect 6412 31692 6468 31694
rect 6572 31746 6628 31748
rect 6572 31694 6574 31746
rect 6574 31694 6626 31746
rect 6626 31694 6628 31746
rect 6572 31692 6628 31694
rect 6732 31746 6788 31748
rect 6732 31694 6734 31746
rect 6734 31694 6786 31746
rect 6786 31694 6788 31746
rect 6732 31692 6788 31694
rect 6892 31746 6948 31748
rect 6892 31694 6894 31746
rect 6894 31694 6946 31746
rect 6946 31694 6948 31746
rect 6892 31692 6948 31694
rect 7052 31746 7108 31748
rect 7052 31694 7054 31746
rect 7054 31694 7106 31746
rect 7106 31694 7108 31746
rect 7052 31692 7108 31694
rect 7212 31746 7268 31748
rect 7212 31694 7214 31746
rect 7214 31694 7266 31746
rect 7266 31694 7268 31746
rect 7212 31692 7268 31694
rect 7372 31746 7428 31748
rect 7372 31694 7374 31746
rect 7374 31694 7426 31746
rect 7426 31694 7428 31746
rect 7372 31692 7428 31694
rect 7532 31746 7588 31748
rect 7532 31694 7534 31746
rect 7534 31694 7586 31746
rect 7586 31694 7588 31746
rect 7532 31692 7588 31694
rect 7692 31746 7748 31748
rect 7692 31694 7694 31746
rect 7694 31694 7746 31746
rect 7746 31694 7748 31746
rect 7692 31692 7748 31694
rect 7852 31746 7908 31748
rect 7852 31694 7854 31746
rect 7854 31694 7906 31746
rect 7906 31694 7908 31746
rect 7852 31692 7908 31694
rect 8012 31746 8068 31748
rect 8012 31694 8014 31746
rect 8014 31694 8066 31746
rect 8066 31694 8068 31746
rect 8012 31692 8068 31694
rect 8172 31746 8228 31748
rect 8172 31694 8174 31746
rect 8174 31694 8226 31746
rect 8226 31694 8228 31746
rect 8172 31692 8228 31694
rect 8332 31746 8388 31748
rect 8332 31694 8334 31746
rect 8334 31694 8386 31746
rect 8386 31694 8388 31746
rect 8332 31692 8388 31694
rect 9452 31692 9508 31748
rect 9772 31692 9828 31748
rect 10092 31692 10148 31748
rect 10412 31692 10468 31748
rect 10732 31692 10788 31748
rect 11052 31692 11108 31748
rect 11372 31692 11428 31748
rect 12492 31746 12548 31748
rect 12492 31694 12494 31746
rect 12494 31694 12546 31746
rect 12546 31694 12548 31746
rect 12492 31692 12548 31694
rect 12652 31746 12708 31748
rect 12652 31694 12654 31746
rect 12654 31694 12706 31746
rect 12706 31694 12708 31746
rect 12652 31692 12708 31694
rect 12812 31746 12868 31748
rect 12812 31694 12814 31746
rect 12814 31694 12866 31746
rect 12866 31694 12868 31746
rect 12812 31692 12868 31694
rect 12972 31746 13028 31748
rect 12972 31694 12974 31746
rect 12974 31694 13026 31746
rect 13026 31694 13028 31746
rect 12972 31692 13028 31694
rect 13132 31746 13188 31748
rect 13132 31694 13134 31746
rect 13134 31694 13186 31746
rect 13186 31694 13188 31746
rect 13132 31692 13188 31694
rect 13292 31746 13348 31748
rect 13292 31694 13294 31746
rect 13294 31694 13346 31746
rect 13346 31694 13348 31746
rect 13292 31692 13348 31694
rect 13452 31746 13508 31748
rect 13452 31694 13454 31746
rect 13454 31694 13506 31746
rect 13506 31694 13508 31746
rect 13452 31692 13508 31694
rect 13612 31746 13668 31748
rect 13612 31694 13614 31746
rect 13614 31694 13666 31746
rect 13666 31694 13668 31746
rect 13612 31692 13668 31694
rect 13772 31746 13828 31748
rect 13772 31694 13774 31746
rect 13774 31694 13826 31746
rect 13826 31694 13828 31746
rect 13772 31692 13828 31694
rect 13932 31746 13988 31748
rect 13932 31694 13934 31746
rect 13934 31694 13986 31746
rect 13986 31694 13988 31746
rect 13932 31692 13988 31694
rect 14092 31746 14148 31748
rect 14092 31694 14094 31746
rect 14094 31694 14146 31746
rect 14146 31694 14148 31746
rect 14092 31692 14148 31694
rect 14252 31746 14308 31748
rect 14252 31694 14254 31746
rect 14254 31694 14306 31746
rect 14306 31694 14308 31746
rect 14252 31692 14308 31694
rect 14412 31746 14468 31748
rect 14412 31694 14414 31746
rect 14414 31694 14466 31746
rect 14466 31694 14468 31746
rect 14412 31692 14468 31694
rect 14572 31746 14628 31748
rect 14572 31694 14574 31746
rect 14574 31694 14626 31746
rect 14626 31694 14628 31746
rect 14572 31692 14628 31694
rect 14732 31746 14788 31748
rect 14732 31694 14734 31746
rect 14734 31694 14786 31746
rect 14786 31694 14788 31746
rect 14732 31692 14788 31694
rect 14892 31746 14948 31748
rect 14892 31694 14894 31746
rect 14894 31694 14946 31746
rect 14946 31694 14948 31746
rect 14892 31692 14948 31694
rect 15052 31746 15108 31748
rect 15052 31694 15054 31746
rect 15054 31694 15106 31746
rect 15106 31694 15108 31746
rect 15052 31692 15108 31694
rect 15212 31746 15268 31748
rect 15212 31694 15214 31746
rect 15214 31694 15266 31746
rect 15266 31694 15268 31746
rect 15212 31692 15268 31694
rect 15372 31746 15428 31748
rect 15372 31694 15374 31746
rect 15374 31694 15426 31746
rect 15426 31694 15428 31746
rect 15372 31692 15428 31694
rect 15532 31746 15588 31748
rect 15532 31694 15534 31746
rect 15534 31694 15586 31746
rect 15586 31694 15588 31746
rect 15532 31692 15588 31694
rect 15692 31746 15748 31748
rect 15692 31694 15694 31746
rect 15694 31694 15746 31746
rect 15746 31694 15748 31746
rect 15692 31692 15748 31694
rect 15852 31746 15908 31748
rect 15852 31694 15854 31746
rect 15854 31694 15906 31746
rect 15906 31694 15908 31746
rect 15852 31692 15908 31694
rect 16012 31746 16068 31748
rect 16012 31694 16014 31746
rect 16014 31694 16066 31746
rect 16066 31694 16068 31746
rect 16012 31692 16068 31694
rect 16172 31746 16228 31748
rect 16172 31694 16174 31746
rect 16174 31694 16226 31746
rect 16226 31694 16228 31746
rect 16172 31692 16228 31694
rect 16332 31746 16388 31748
rect 16332 31694 16334 31746
rect 16334 31694 16386 31746
rect 16386 31694 16388 31746
rect 16332 31692 16388 31694
rect 16492 31746 16548 31748
rect 16492 31694 16494 31746
rect 16494 31694 16546 31746
rect 16546 31694 16548 31746
rect 16492 31692 16548 31694
rect 16652 31746 16708 31748
rect 16652 31694 16654 31746
rect 16654 31694 16706 31746
rect 16706 31694 16708 31746
rect 16652 31692 16708 31694
rect 16812 31746 16868 31748
rect 16812 31694 16814 31746
rect 16814 31694 16866 31746
rect 16866 31694 16868 31746
rect 16812 31692 16868 31694
rect 16972 31746 17028 31748
rect 16972 31694 16974 31746
rect 16974 31694 17026 31746
rect 17026 31694 17028 31746
rect 16972 31692 17028 31694
rect 17132 31746 17188 31748
rect 17132 31694 17134 31746
rect 17134 31694 17186 31746
rect 17186 31694 17188 31746
rect 17132 31692 17188 31694
rect 17292 31746 17348 31748
rect 17292 31694 17294 31746
rect 17294 31694 17346 31746
rect 17346 31694 17348 31746
rect 17292 31692 17348 31694
rect 17452 31746 17508 31748
rect 17452 31694 17454 31746
rect 17454 31694 17506 31746
rect 17506 31694 17508 31746
rect 17452 31692 17508 31694
rect 17612 31746 17668 31748
rect 17612 31694 17614 31746
rect 17614 31694 17666 31746
rect 17666 31694 17668 31746
rect 17612 31692 17668 31694
rect 17772 31746 17828 31748
rect 17772 31694 17774 31746
rect 17774 31694 17826 31746
rect 17826 31694 17828 31746
rect 17772 31692 17828 31694
rect 17932 31746 17988 31748
rect 17932 31694 17934 31746
rect 17934 31694 17986 31746
rect 17986 31694 17988 31746
rect 17932 31692 17988 31694
rect 18092 31746 18148 31748
rect 18092 31694 18094 31746
rect 18094 31694 18146 31746
rect 18146 31694 18148 31746
rect 18092 31692 18148 31694
rect 18252 31746 18308 31748
rect 18252 31694 18254 31746
rect 18254 31694 18306 31746
rect 18306 31694 18308 31746
rect 18252 31692 18308 31694
rect 18412 31746 18468 31748
rect 18412 31694 18414 31746
rect 18414 31694 18466 31746
rect 18466 31694 18468 31746
rect 18412 31692 18468 31694
rect 18572 31746 18628 31748
rect 18572 31694 18574 31746
rect 18574 31694 18626 31746
rect 18626 31694 18628 31746
rect 18572 31692 18628 31694
rect 18732 31746 18788 31748
rect 18732 31694 18734 31746
rect 18734 31694 18786 31746
rect 18786 31694 18788 31746
rect 18732 31692 18788 31694
rect 18892 31746 18948 31748
rect 18892 31694 18894 31746
rect 18894 31694 18946 31746
rect 18946 31694 18948 31746
rect 18892 31692 18948 31694
rect 20012 31692 20068 31748
rect 20332 31692 20388 31748
rect 20652 31692 20708 31748
rect 20972 31692 21028 31748
rect 21292 31692 21348 31748
rect 21612 31692 21668 31748
rect 21932 31692 21988 31748
rect 23132 31746 23188 31748
rect 23132 31694 23134 31746
rect 23134 31694 23186 31746
rect 23186 31694 23188 31746
rect 23132 31692 23188 31694
rect 23292 31746 23348 31748
rect 23292 31694 23294 31746
rect 23294 31694 23346 31746
rect 23346 31694 23348 31746
rect 23292 31692 23348 31694
rect 23452 31746 23508 31748
rect 23452 31694 23454 31746
rect 23454 31694 23506 31746
rect 23506 31694 23508 31746
rect 23452 31692 23508 31694
rect 23612 31746 23668 31748
rect 23612 31694 23614 31746
rect 23614 31694 23666 31746
rect 23666 31694 23668 31746
rect 23612 31692 23668 31694
rect 23772 31746 23828 31748
rect 23772 31694 23774 31746
rect 23774 31694 23826 31746
rect 23826 31694 23828 31746
rect 23772 31692 23828 31694
rect 23932 31746 23988 31748
rect 23932 31694 23934 31746
rect 23934 31694 23986 31746
rect 23986 31694 23988 31746
rect 23932 31692 23988 31694
rect 24092 31746 24148 31748
rect 24092 31694 24094 31746
rect 24094 31694 24146 31746
rect 24146 31694 24148 31746
rect 24092 31692 24148 31694
rect 24252 31746 24308 31748
rect 24252 31694 24254 31746
rect 24254 31694 24306 31746
rect 24306 31694 24308 31746
rect 24252 31692 24308 31694
rect 24412 31746 24468 31748
rect 24412 31694 24414 31746
rect 24414 31694 24466 31746
rect 24466 31694 24468 31746
rect 24412 31692 24468 31694
rect 24572 31746 24628 31748
rect 24572 31694 24574 31746
rect 24574 31694 24626 31746
rect 24626 31694 24628 31746
rect 24572 31692 24628 31694
rect 24732 31746 24788 31748
rect 24732 31694 24734 31746
rect 24734 31694 24786 31746
rect 24786 31694 24788 31746
rect 24732 31692 24788 31694
rect 24892 31746 24948 31748
rect 24892 31694 24894 31746
rect 24894 31694 24946 31746
rect 24946 31694 24948 31746
rect 24892 31692 24948 31694
rect 25052 31746 25108 31748
rect 25052 31694 25054 31746
rect 25054 31694 25106 31746
rect 25106 31694 25108 31746
rect 25052 31692 25108 31694
rect 25212 31746 25268 31748
rect 25212 31694 25214 31746
rect 25214 31694 25266 31746
rect 25266 31694 25268 31746
rect 25212 31692 25268 31694
rect 25372 31746 25428 31748
rect 25372 31694 25374 31746
rect 25374 31694 25426 31746
rect 25426 31694 25428 31746
rect 25372 31692 25428 31694
rect 25532 31746 25588 31748
rect 25532 31694 25534 31746
rect 25534 31694 25586 31746
rect 25586 31694 25588 31746
rect 25532 31692 25588 31694
rect 25692 31746 25748 31748
rect 25692 31694 25694 31746
rect 25694 31694 25746 31746
rect 25746 31694 25748 31746
rect 25692 31692 25748 31694
rect 25852 31746 25908 31748
rect 25852 31694 25854 31746
rect 25854 31694 25906 31746
rect 25906 31694 25908 31746
rect 25852 31692 25908 31694
rect 26012 31746 26068 31748
rect 26012 31694 26014 31746
rect 26014 31694 26066 31746
rect 26066 31694 26068 31746
rect 26012 31692 26068 31694
rect 26172 31746 26228 31748
rect 26172 31694 26174 31746
rect 26174 31694 26226 31746
rect 26226 31694 26228 31746
rect 26172 31692 26228 31694
rect 26332 31746 26388 31748
rect 26332 31694 26334 31746
rect 26334 31694 26386 31746
rect 26386 31694 26388 31746
rect 26332 31692 26388 31694
rect 26492 31746 26548 31748
rect 26492 31694 26494 31746
rect 26494 31694 26546 31746
rect 26546 31694 26548 31746
rect 26492 31692 26548 31694
rect 26652 31746 26708 31748
rect 26652 31694 26654 31746
rect 26654 31694 26706 31746
rect 26706 31694 26708 31746
rect 26652 31692 26708 31694
rect 26812 31746 26868 31748
rect 26812 31694 26814 31746
rect 26814 31694 26866 31746
rect 26866 31694 26868 31746
rect 26812 31692 26868 31694
rect 26972 31746 27028 31748
rect 26972 31694 26974 31746
rect 26974 31694 27026 31746
rect 27026 31694 27028 31746
rect 26972 31692 27028 31694
rect 27132 31746 27188 31748
rect 27132 31694 27134 31746
rect 27134 31694 27186 31746
rect 27186 31694 27188 31746
rect 27132 31692 27188 31694
rect 27292 31746 27348 31748
rect 27292 31694 27294 31746
rect 27294 31694 27346 31746
rect 27346 31694 27348 31746
rect 27292 31692 27348 31694
rect 27452 31746 27508 31748
rect 27452 31694 27454 31746
rect 27454 31694 27506 31746
rect 27506 31694 27508 31746
rect 27452 31692 27508 31694
rect 27612 31746 27668 31748
rect 27612 31694 27614 31746
rect 27614 31694 27666 31746
rect 27666 31694 27668 31746
rect 27612 31692 27668 31694
rect 27772 31746 27828 31748
rect 27772 31694 27774 31746
rect 27774 31694 27826 31746
rect 27826 31694 27828 31746
rect 27772 31692 27828 31694
rect 27932 31746 27988 31748
rect 27932 31694 27934 31746
rect 27934 31694 27986 31746
rect 27986 31694 27988 31746
rect 27932 31692 27988 31694
rect 28092 31746 28148 31748
rect 28092 31694 28094 31746
rect 28094 31694 28146 31746
rect 28146 31694 28148 31746
rect 28092 31692 28148 31694
rect 28252 31746 28308 31748
rect 28252 31694 28254 31746
rect 28254 31694 28306 31746
rect 28306 31694 28308 31746
rect 28252 31692 28308 31694
rect 28412 31746 28468 31748
rect 28412 31694 28414 31746
rect 28414 31694 28466 31746
rect 28466 31694 28468 31746
rect 28412 31692 28468 31694
rect 28572 31746 28628 31748
rect 28572 31694 28574 31746
rect 28574 31694 28626 31746
rect 28626 31694 28628 31746
rect 28572 31692 28628 31694
rect 28732 31746 28788 31748
rect 28732 31694 28734 31746
rect 28734 31694 28786 31746
rect 28786 31694 28788 31746
rect 28732 31692 28788 31694
rect 28892 31746 28948 31748
rect 28892 31694 28894 31746
rect 28894 31694 28946 31746
rect 28946 31694 28948 31746
rect 28892 31692 28948 31694
rect 29052 31746 29108 31748
rect 29052 31694 29054 31746
rect 29054 31694 29106 31746
rect 29106 31694 29108 31746
rect 29052 31692 29108 31694
rect 29212 31746 29268 31748
rect 29212 31694 29214 31746
rect 29214 31694 29266 31746
rect 29266 31694 29268 31746
rect 29212 31692 29268 31694
rect 29372 31746 29428 31748
rect 29372 31694 29374 31746
rect 29374 31694 29426 31746
rect 29426 31694 29428 31746
rect 29372 31692 29428 31694
rect 30492 31692 30548 31748
rect 30812 31692 30868 31748
rect 31132 31692 31188 31748
rect 31452 31692 31508 31748
rect 31772 31692 31828 31748
rect 32092 31692 32148 31748
rect 32412 31692 32468 31748
rect 33532 31746 33588 31748
rect 33532 31694 33534 31746
rect 33534 31694 33586 31746
rect 33586 31694 33588 31746
rect 33532 31692 33588 31694
rect 33692 31746 33748 31748
rect 33692 31694 33694 31746
rect 33694 31694 33746 31746
rect 33746 31694 33748 31746
rect 33692 31692 33748 31694
rect 33852 31746 33908 31748
rect 33852 31694 33854 31746
rect 33854 31694 33906 31746
rect 33906 31694 33908 31746
rect 33852 31692 33908 31694
rect 34012 31746 34068 31748
rect 34012 31694 34014 31746
rect 34014 31694 34066 31746
rect 34066 31694 34068 31746
rect 34012 31692 34068 31694
rect 34172 31746 34228 31748
rect 34172 31694 34174 31746
rect 34174 31694 34226 31746
rect 34226 31694 34228 31746
rect 34172 31692 34228 31694
rect 34332 31746 34388 31748
rect 34332 31694 34334 31746
rect 34334 31694 34386 31746
rect 34386 31694 34388 31746
rect 34332 31692 34388 31694
rect 34492 31746 34548 31748
rect 34492 31694 34494 31746
rect 34494 31694 34546 31746
rect 34546 31694 34548 31746
rect 34492 31692 34548 31694
rect 34652 31746 34708 31748
rect 34652 31694 34654 31746
rect 34654 31694 34706 31746
rect 34706 31694 34708 31746
rect 34652 31692 34708 31694
rect 34812 31746 34868 31748
rect 34812 31694 34814 31746
rect 34814 31694 34866 31746
rect 34866 31694 34868 31746
rect 34812 31692 34868 31694
rect 34972 31746 35028 31748
rect 34972 31694 34974 31746
rect 34974 31694 35026 31746
rect 35026 31694 35028 31746
rect 34972 31692 35028 31694
rect 35132 31746 35188 31748
rect 35132 31694 35134 31746
rect 35134 31694 35186 31746
rect 35186 31694 35188 31746
rect 35132 31692 35188 31694
rect 35292 31746 35348 31748
rect 35292 31694 35294 31746
rect 35294 31694 35346 31746
rect 35346 31694 35348 31746
rect 35292 31692 35348 31694
rect 35452 31746 35508 31748
rect 35452 31694 35454 31746
rect 35454 31694 35506 31746
rect 35506 31694 35508 31746
rect 35452 31692 35508 31694
rect 35612 31746 35668 31748
rect 35612 31694 35614 31746
rect 35614 31694 35666 31746
rect 35666 31694 35668 31746
rect 35612 31692 35668 31694
rect 35772 31746 35828 31748
rect 35772 31694 35774 31746
rect 35774 31694 35826 31746
rect 35826 31694 35828 31746
rect 35772 31692 35828 31694
rect 35932 31746 35988 31748
rect 35932 31694 35934 31746
rect 35934 31694 35986 31746
rect 35986 31694 35988 31746
rect 35932 31692 35988 31694
rect 36092 31746 36148 31748
rect 36092 31694 36094 31746
rect 36094 31694 36146 31746
rect 36146 31694 36148 31746
rect 36092 31692 36148 31694
rect 36252 31746 36308 31748
rect 36252 31694 36254 31746
rect 36254 31694 36306 31746
rect 36306 31694 36308 31746
rect 36252 31692 36308 31694
rect 36412 31746 36468 31748
rect 36412 31694 36414 31746
rect 36414 31694 36466 31746
rect 36466 31694 36468 31746
rect 36412 31692 36468 31694
rect 36572 31746 36628 31748
rect 36572 31694 36574 31746
rect 36574 31694 36626 31746
rect 36626 31694 36628 31746
rect 36572 31692 36628 31694
rect 36732 31746 36788 31748
rect 36732 31694 36734 31746
rect 36734 31694 36786 31746
rect 36786 31694 36788 31746
rect 36732 31692 36788 31694
rect 36892 31746 36948 31748
rect 36892 31694 36894 31746
rect 36894 31694 36946 31746
rect 36946 31694 36948 31746
rect 36892 31692 36948 31694
rect 37052 31746 37108 31748
rect 37052 31694 37054 31746
rect 37054 31694 37106 31746
rect 37106 31694 37108 31746
rect 37052 31692 37108 31694
rect 37212 31746 37268 31748
rect 37212 31694 37214 31746
rect 37214 31694 37266 31746
rect 37266 31694 37268 31746
rect 37212 31692 37268 31694
rect 37372 31746 37428 31748
rect 37372 31694 37374 31746
rect 37374 31694 37426 31746
rect 37426 31694 37428 31746
rect 37372 31692 37428 31694
rect 37532 31746 37588 31748
rect 37532 31694 37534 31746
rect 37534 31694 37586 31746
rect 37586 31694 37588 31746
rect 37532 31692 37588 31694
rect 37692 31746 37748 31748
rect 37692 31694 37694 31746
rect 37694 31694 37746 31746
rect 37746 31694 37748 31746
rect 37692 31692 37748 31694
rect 37852 31746 37908 31748
rect 37852 31694 37854 31746
rect 37854 31694 37906 31746
rect 37906 31694 37908 31746
rect 37852 31692 37908 31694
rect 38012 31746 38068 31748
rect 38012 31694 38014 31746
rect 38014 31694 38066 31746
rect 38066 31694 38068 31746
rect 38012 31692 38068 31694
rect 38172 31746 38228 31748
rect 38172 31694 38174 31746
rect 38174 31694 38226 31746
rect 38226 31694 38228 31746
rect 38172 31692 38228 31694
rect 38332 31746 38388 31748
rect 38332 31694 38334 31746
rect 38334 31694 38386 31746
rect 38386 31694 38388 31746
rect 38332 31692 38388 31694
rect 38492 31746 38548 31748
rect 38492 31694 38494 31746
rect 38494 31694 38546 31746
rect 38546 31694 38548 31746
rect 38492 31692 38548 31694
rect 38652 31746 38708 31748
rect 38652 31694 38654 31746
rect 38654 31694 38706 31746
rect 38706 31694 38708 31746
rect 38652 31692 38708 31694
rect 38812 31746 38868 31748
rect 38812 31694 38814 31746
rect 38814 31694 38866 31746
rect 38866 31694 38868 31746
rect 38812 31692 38868 31694
rect 38972 31746 39028 31748
rect 38972 31694 38974 31746
rect 38974 31694 39026 31746
rect 39026 31694 39028 31746
rect 38972 31692 39028 31694
rect 39132 31746 39188 31748
rect 39132 31694 39134 31746
rect 39134 31694 39186 31746
rect 39186 31694 39188 31746
rect 39132 31692 39188 31694
rect 39292 31746 39348 31748
rect 39292 31694 39294 31746
rect 39294 31694 39346 31746
rect 39346 31694 39348 31746
rect 39292 31692 39348 31694
rect 39452 31746 39508 31748
rect 39452 31694 39454 31746
rect 39454 31694 39506 31746
rect 39506 31694 39508 31746
rect 39452 31692 39508 31694
rect 39612 31746 39668 31748
rect 39612 31694 39614 31746
rect 39614 31694 39666 31746
rect 39666 31694 39668 31746
rect 39612 31692 39668 31694
rect 39772 31746 39828 31748
rect 39772 31694 39774 31746
rect 39774 31694 39826 31746
rect 39826 31694 39828 31746
rect 39772 31692 39828 31694
rect 39932 31746 39988 31748
rect 39932 31694 39934 31746
rect 39934 31694 39986 31746
rect 39986 31694 39988 31746
rect 39932 31692 39988 31694
rect 40092 31746 40148 31748
rect 40092 31694 40094 31746
rect 40094 31694 40146 31746
rect 40146 31694 40148 31746
rect 40092 31692 40148 31694
rect 40252 31746 40308 31748
rect 40252 31694 40254 31746
rect 40254 31694 40306 31746
rect 40306 31694 40308 31746
rect 40252 31692 40308 31694
rect 40412 31746 40468 31748
rect 40412 31694 40414 31746
rect 40414 31694 40466 31746
rect 40466 31694 40468 31746
rect 40412 31692 40468 31694
rect 40572 31746 40628 31748
rect 40572 31694 40574 31746
rect 40574 31694 40626 31746
rect 40626 31694 40628 31746
rect 40572 31692 40628 31694
rect 40732 31746 40788 31748
rect 40732 31694 40734 31746
rect 40734 31694 40786 31746
rect 40786 31694 40788 31746
rect 40732 31692 40788 31694
rect 40892 31746 40948 31748
rect 40892 31694 40894 31746
rect 40894 31694 40946 31746
rect 40946 31694 40948 31746
rect 40892 31692 40948 31694
rect 41052 31746 41108 31748
rect 41052 31694 41054 31746
rect 41054 31694 41106 31746
rect 41106 31694 41108 31746
rect 41052 31692 41108 31694
rect 41212 31746 41268 31748
rect 41212 31694 41214 31746
rect 41214 31694 41266 31746
rect 41266 31694 41268 31746
rect 41212 31692 41268 31694
rect 41372 31746 41428 31748
rect 41372 31694 41374 31746
rect 41374 31694 41426 31746
rect 41426 31694 41428 31746
rect 41372 31692 41428 31694
rect 41532 31746 41588 31748
rect 41532 31694 41534 31746
rect 41534 31694 41586 31746
rect 41586 31694 41588 31746
rect 41532 31692 41588 31694
rect 41692 31746 41748 31748
rect 41692 31694 41694 31746
rect 41694 31694 41746 31746
rect 41746 31694 41748 31746
rect 41692 31692 41748 31694
rect 41852 31746 41908 31748
rect 41852 31694 41854 31746
rect 41854 31694 41906 31746
rect 41906 31694 41908 31746
rect 41852 31692 41908 31694
rect 10252 31532 10308 31588
rect 20812 31532 20868 31588
rect 31612 31532 31668 31588
rect 12 31426 68 31428
rect 12 31374 14 31426
rect 14 31374 66 31426
rect 66 31374 68 31426
rect 12 31372 68 31374
rect 172 31426 228 31428
rect 172 31374 174 31426
rect 174 31374 226 31426
rect 226 31374 228 31426
rect 172 31372 228 31374
rect 332 31426 388 31428
rect 332 31374 334 31426
rect 334 31374 386 31426
rect 386 31374 388 31426
rect 332 31372 388 31374
rect 492 31426 548 31428
rect 492 31374 494 31426
rect 494 31374 546 31426
rect 546 31374 548 31426
rect 492 31372 548 31374
rect 652 31426 708 31428
rect 652 31374 654 31426
rect 654 31374 706 31426
rect 706 31374 708 31426
rect 652 31372 708 31374
rect 812 31426 868 31428
rect 812 31374 814 31426
rect 814 31374 866 31426
rect 866 31374 868 31426
rect 812 31372 868 31374
rect 972 31426 1028 31428
rect 972 31374 974 31426
rect 974 31374 1026 31426
rect 1026 31374 1028 31426
rect 972 31372 1028 31374
rect 1132 31426 1188 31428
rect 1132 31374 1134 31426
rect 1134 31374 1186 31426
rect 1186 31374 1188 31426
rect 1132 31372 1188 31374
rect 1292 31426 1348 31428
rect 1292 31374 1294 31426
rect 1294 31374 1346 31426
rect 1346 31374 1348 31426
rect 1292 31372 1348 31374
rect 1452 31426 1508 31428
rect 1452 31374 1454 31426
rect 1454 31374 1506 31426
rect 1506 31374 1508 31426
rect 1452 31372 1508 31374
rect 1612 31426 1668 31428
rect 1612 31374 1614 31426
rect 1614 31374 1666 31426
rect 1666 31374 1668 31426
rect 1612 31372 1668 31374
rect 1772 31426 1828 31428
rect 1772 31374 1774 31426
rect 1774 31374 1826 31426
rect 1826 31374 1828 31426
rect 1772 31372 1828 31374
rect 1932 31426 1988 31428
rect 1932 31374 1934 31426
rect 1934 31374 1986 31426
rect 1986 31374 1988 31426
rect 1932 31372 1988 31374
rect 2092 31426 2148 31428
rect 2092 31374 2094 31426
rect 2094 31374 2146 31426
rect 2146 31374 2148 31426
rect 2092 31372 2148 31374
rect 2252 31426 2308 31428
rect 2252 31374 2254 31426
rect 2254 31374 2306 31426
rect 2306 31374 2308 31426
rect 2252 31372 2308 31374
rect 2412 31426 2468 31428
rect 2412 31374 2414 31426
rect 2414 31374 2466 31426
rect 2466 31374 2468 31426
rect 2412 31372 2468 31374
rect 2572 31426 2628 31428
rect 2572 31374 2574 31426
rect 2574 31374 2626 31426
rect 2626 31374 2628 31426
rect 2572 31372 2628 31374
rect 2732 31426 2788 31428
rect 2732 31374 2734 31426
rect 2734 31374 2786 31426
rect 2786 31374 2788 31426
rect 2732 31372 2788 31374
rect 2892 31426 2948 31428
rect 2892 31374 2894 31426
rect 2894 31374 2946 31426
rect 2946 31374 2948 31426
rect 2892 31372 2948 31374
rect 3052 31426 3108 31428
rect 3052 31374 3054 31426
rect 3054 31374 3106 31426
rect 3106 31374 3108 31426
rect 3052 31372 3108 31374
rect 3212 31426 3268 31428
rect 3212 31374 3214 31426
rect 3214 31374 3266 31426
rect 3266 31374 3268 31426
rect 3212 31372 3268 31374
rect 3372 31426 3428 31428
rect 3372 31374 3374 31426
rect 3374 31374 3426 31426
rect 3426 31374 3428 31426
rect 3372 31372 3428 31374
rect 3532 31426 3588 31428
rect 3532 31374 3534 31426
rect 3534 31374 3586 31426
rect 3586 31374 3588 31426
rect 3532 31372 3588 31374
rect 3692 31426 3748 31428
rect 3692 31374 3694 31426
rect 3694 31374 3746 31426
rect 3746 31374 3748 31426
rect 3692 31372 3748 31374
rect 3852 31426 3908 31428
rect 3852 31374 3854 31426
rect 3854 31374 3906 31426
rect 3906 31374 3908 31426
rect 3852 31372 3908 31374
rect 4012 31426 4068 31428
rect 4012 31374 4014 31426
rect 4014 31374 4066 31426
rect 4066 31374 4068 31426
rect 4012 31372 4068 31374
rect 4172 31426 4228 31428
rect 4172 31374 4174 31426
rect 4174 31374 4226 31426
rect 4226 31374 4228 31426
rect 4172 31372 4228 31374
rect 4332 31426 4388 31428
rect 4332 31374 4334 31426
rect 4334 31374 4386 31426
rect 4386 31374 4388 31426
rect 4332 31372 4388 31374
rect 4492 31426 4548 31428
rect 4492 31374 4494 31426
rect 4494 31374 4546 31426
rect 4546 31374 4548 31426
rect 4492 31372 4548 31374
rect 4652 31426 4708 31428
rect 4652 31374 4654 31426
rect 4654 31374 4706 31426
rect 4706 31374 4708 31426
rect 4652 31372 4708 31374
rect 4812 31426 4868 31428
rect 4812 31374 4814 31426
rect 4814 31374 4866 31426
rect 4866 31374 4868 31426
rect 4812 31372 4868 31374
rect 4972 31426 5028 31428
rect 4972 31374 4974 31426
rect 4974 31374 5026 31426
rect 5026 31374 5028 31426
rect 4972 31372 5028 31374
rect 5132 31426 5188 31428
rect 5132 31374 5134 31426
rect 5134 31374 5186 31426
rect 5186 31374 5188 31426
rect 5132 31372 5188 31374
rect 5292 31426 5348 31428
rect 5292 31374 5294 31426
rect 5294 31374 5346 31426
rect 5346 31374 5348 31426
rect 5292 31372 5348 31374
rect 5452 31426 5508 31428
rect 5452 31374 5454 31426
rect 5454 31374 5506 31426
rect 5506 31374 5508 31426
rect 5452 31372 5508 31374
rect 5612 31426 5668 31428
rect 5612 31374 5614 31426
rect 5614 31374 5666 31426
rect 5666 31374 5668 31426
rect 5612 31372 5668 31374
rect 5772 31426 5828 31428
rect 5772 31374 5774 31426
rect 5774 31374 5826 31426
rect 5826 31374 5828 31426
rect 5772 31372 5828 31374
rect 5932 31426 5988 31428
rect 5932 31374 5934 31426
rect 5934 31374 5986 31426
rect 5986 31374 5988 31426
rect 5932 31372 5988 31374
rect 6092 31426 6148 31428
rect 6092 31374 6094 31426
rect 6094 31374 6146 31426
rect 6146 31374 6148 31426
rect 6092 31372 6148 31374
rect 6252 31426 6308 31428
rect 6252 31374 6254 31426
rect 6254 31374 6306 31426
rect 6306 31374 6308 31426
rect 6252 31372 6308 31374
rect 6412 31426 6468 31428
rect 6412 31374 6414 31426
rect 6414 31374 6466 31426
rect 6466 31374 6468 31426
rect 6412 31372 6468 31374
rect 6572 31426 6628 31428
rect 6572 31374 6574 31426
rect 6574 31374 6626 31426
rect 6626 31374 6628 31426
rect 6572 31372 6628 31374
rect 6732 31426 6788 31428
rect 6732 31374 6734 31426
rect 6734 31374 6786 31426
rect 6786 31374 6788 31426
rect 6732 31372 6788 31374
rect 6892 31426 6948 31428
rect 6892 31374 6894 31426
rect 6894 31374 6946 31426
rect 6946 31374 6948 31426
rect 6892 31372 6948 31374
rect 7052 31426 7108 31428
rect 7052 31374 7054 31426
rect 7054 31374 7106 31426
rect 7106 31374 7108 31426
rect 7052 31372 7108 31374
rect 7212 31426 7268 31428
rect 7212 31374 7214 31426
rect 7214 31374 7266 31426
rect 7266 31374 7268 31426
rect 7212 31372 7268 31374
rect 7372 31426 7428 31428
rect 7372 31374 7374 31426
rect 7374 31374 7426 31426
rect 7426 31374 7428 31426
rect 7372 31372 7428 31374
rect 7532 31426 7588 31428
rect 7532 31374 7534 31426
rect 7534 31374 7586 31426
rect 7586 31374 7588 31426
rect 7532 31372 7588 31374
rect 7692 31426 7748 31428
rect 7692 31374 7694 31426
rect 7694 31374 7746 31426
rect 7746 31374 7748 31426
rect 7692 31372 7748 31374
rect 7852 31426 7908 31428
rect 7852 31374 7854 31426
rect 7854 31374 7906 31426
rect 7906 31374 7908 31426
rect 7852 31372 7908 31374
rect 8012 31426 8068 31428
rect 8012 31374 8014 31426
rect 8014 31374 8066 31426
rect 8066 31374 8068 31426
rect 8012 31372 8068 31374
rect 8172 31426 8228 31428
rect 8172 31374 8174 31426
rect 8174 31374 8226 31426
rect 8226 31374 8228 31426
rect 8172 31372 8228 31374
rect 8332 31426 8388 31428
rect 8332 31374 8334 31426
rect 8334 31374 8386 31426
rect 8386 31374 8388 31426
rect 8332 31372 8388 31374
rect 9452 31372 9508 31428
rect 9772 31372 9828 31428
rect 10092 31372 10148 31428
rect 10412 31372 10468 31428
rect 10732 31372 10788 31428
rect 11052 31372 11108 31428
rect 11372 31372 11428 31428
rect 12492 31426 12548 31428
rect 12492 31374 12494 31426
rect 12494 31374 12546 31426
rect 12546 31374 12548 31426
rect 12492 31372 12548 31374
rect 12652 31426 12708 31428
rect 12652 31374 12654 31426
rect 12654 31374 12706 31426
rect 12706 31374 12708 31426
rect 12652 31372 12708 31374
rect 12812 31426 12868 31428
rect 12812 31374 12814 31426
rect 12814 31374 12866 31426
rect 12866 31374 12868 31426
rect 12812 31372 12868 31374
rect 12972 31426 13028 31428
rect 12972 31374 12974 31426
rect 12974 31374 13026 31426
rect 13026 31374 13028 31426
rect 12972 31372 13028 31374
rect 13132 31426 13188 31428
rect 13132 31374 13134 31426
rect 13134 31374 13186 31426
rect 13186 31374 13188 31426
rect 13132 31372 13188 31374
rect 13292 31426 13348 31428
rect 13292 31374 13294 31426
rect 13294 31374 13346 31426
rect 13346 31374 13348 31426
rect 13292 31372 13348 31374
rect 13452 31426 13508 31428
rect 13452 31374 13454 31426
rect 13454 31374 13506 31426
rect 13506 31374 13508 31426
rect 13452 31372 13508 31374
rect 13612 31426 13668 31428
rect 13612 31374 13614 31426
rect 13614 31374 13666 31426
rect 13666 31374 13668 31426
rect 13612 31372 13668 31374
rect 13772 31426 13828 31428
rect 13772 31374 13774 31426
rect 13774 31374 13826 31426
rect 13826 31374 13828 31426
rect 13772 31372 13828 31374
rect 13932 31426 13988 31428
rect 13932 31374 13934 31426
rect 13934 31374 13986 31426
rect 13986 31374 13988 31426
rect 13932 31372 13988 31374
rect 14092 31426 14148 31428
rect 14092 31374 14094 31426
rect 14094 31374 14146 31426
rect 14146 31374 14148 31426
rect 14092 31372 14148 31374
rect 14252 31426 14308 31428
rect 14252 31374 14254 31426
rect 14254 31374 14306 31426
rect 14306 31374 14308 31426
rect 14252 31372 14308 31374
rect 14412 31426 14468 31428
rect 14412 31374 14414 31426
rect 14414 31374 14466 31426
rect 14466 31374 14468 31426
rect 14412 31372 14468 31374
rect 14572 31426 14628 31428
rect 14572 31374 14574 31426
rect 14574 31374 14626 31426
rect 14626 31374 14628 31426
rect 14572 31372 14628 31374
rect 14732 31426 14788 31428
rect 14732 31374 14734 31426
rect 14734 31374 14786 31426
rect 14786 31374 14788 31426
rect 14732 31372 14788 31374
rect 14892 31426 14948 31428
rect 14892 31374 14894 31426
rect 14894 31374 14946 31426
rect 14946 31374 14948 31426
rect 14892 31372 14948 31374
rect 15052 31426 15108 31428
rect 15052 31374 15054 31426
rect 15054 31374 15106 31426
rect 15106 31374 15108 31426
rect 15052 31372 15108 31374
rect 15212 31426 15268 31428
rect 15212 31374 15214 31426
rect 15214 31374 15266 31426
rect 15266 31374 15268 31426
rect 15212 31372 15268 31374
rect 15372 31426 15428 31428
rect 15372 31374 15374 31426
rect 15374 31374 15426 31426
rect 15426 31374 15428 31426
rect 15372 31372 15428 31374
rect 15532 31426 15588 31428
rect 15532 31374 15534 31426
rect 15534 31374 15586 31426
rect 15586 31374 15588 31426
rect 15532 31372 15588 31374
rect 15692 31426 15748 31428
rect 15692 31374 15694 31426
rect 15694 31374 15746 31426
rect 15746 31374 15748 31426
rect 15692 31372 15748 31374
rect 15852 31426 15908 31428
rect 15852 31374 15854 31426
rect 15854 31374 15906 31426
rect 15906 31374 15908 31426
rect 15852 31372 15908 31374
rect 16012 31426 16068 31428
rect 16012 31374 16014 31426
rect 16014 31374 16066 31426
rect 16066 31374 16068 31426
rect 16012 31372 16068 31374
rect 16172 31426 16228 31428
rect 16172 31374 16174 31426
rect 16174 31374 16226 31426
rect 16226 31374 16228 31426
rect 16172 31372 16228 31374
rect 16332 31426 16388 31428
rect 16332 31374 16334 31426
rect 16334 31374 16386 31426
rect 16386 31374 16388 31426
rect 16332 31372 16388 31374
rect 16492 31426 16548 31428
rect 16492 31374 16494 31426
rect 16494 31374 16546 31426
rect 16546 31374 16548 31426
rect 16492 31372 16548 31374
rect 16652 31426 16708 31428
rect 16652 31374 16654 31426
rect 16654 31374 16706 31426
rect 16706 31374 16708 31426
rect 16652 31372 16708 31374
rect 16812 31426 16868 31428
rect 16812 31374 16814 31426
rect 16814 31374 16866 31426
rect 16866 31374 16868 31426
rect 16812 31372 16868 31374
rect 16972 31426 17028 31428
rect 16972 31374 16974 31426
rect 16974 31374 17026 31426
rect 17026 31374 17028 31426
rect 16972 31372 17028 31374
rect 17132 31426 17188 31428
rect 17132 31374 17134 31426
rect 17134 31374 17186 31426
rect 17186 31374 17188 31426
rect 17132 31372 17188 31374
rect 17292 31426 17348 31428
rect 17292 31374 17294 31426
rect 17294 31374 17346 31426
rect 17346 31374 17348 31426
rect 17292 31372 17348 31374
rect 17452 31426 17508 31428
rect 17452 31374 17454 31426
rect 17454 31374 17506 31426
rect 17506 31374 17508 31426
rect 17452 31372 17508 31374
rect 17612 31426 17668 31428
rect 17612 31374 17614 31426
rect 17614 31374 17666 31426
rect 17666 31374 17668 31426
rect 17612 31372 17668 31374
rect 17772 31426 17828 31428
rect 17772 31374 17774 31426
rect 17774 31374 17826 31426
rect 17826 31374 17828 31426
rect 17772 31372 17828 31374
rect 17932 31426 17988 31428
rect 17932 31374 17934 31426
rect 17934 31374 17986 31426
rect 17986 31374 17988 31426
rect 17932 31372 17988 31374
rect 18092 31426 18148 31428
rect 18092 31374 18094 31426
rect 18094 31374 18146 31426
rect 18146 31374 18148 31426
rect 18092 31372 18148 31374
rect 18252 31426 18308 31428
rect 18252 31374 18254 31426
rect 18254 31374 18306 31426
rect 18306 31374 18308 31426
rect 18252 31372 18308 31374
rect 18412 31426 18468 31428
rect 18412 31374 18414 31426
rect 18414 31374 18466 31426
rect 18466 31374 18468 31426
rect 18412 31372 18468 31374
rect 18572 31426 18628 31428
rect 18572 31374 18574 31426
rect 18574 31374 18626 31426
rect 18626 31374 18628 31426
rect 18572 31372 18628 31374
rect 18732 31426 18788 31428
rect 18732 31374 18734 31426
rect 18734 31374 18786 31426
rect 18786 31374 18788 31426
rect 18732 31372 18788 31374
rect 18892 31426 18948 31428
rect 18892 31374 18894 31426
rect 18894 31374 18946 31426
rect 18946 31374 18948 31426
rect 18892 31372 18948 31374
rect 20012 31372 20068 31428
rect 20332 31372 20388 31428
rect 20652 31372 20708 31428
rect 20972 31372 21028 31428
rect 21292 31372 21348 31428
rect 21612 31372 21668 31428
rect 21932 31372 21988 31428
rect 23132 31426 23188 31428
rect 23132 31374 23134 31426
rect 23134 31374 23186 31426
rect 23186 31374 23188 31426
rect 23132 31372 23188 31374
rect 23292 31426 23348 31428
rect 23292 31374 23294 31426
rect 23294 31374 23346 31426
rect 23346 31374 23348 31426
rect 23292 31372 23348 31374
rect 23452 31426 23508 31428
rect 23452 31374 23454 31426
rect 23454 31374 23506 31426
rect 23506 31374 23508 31426
rect 23452 31372 23508 31374
rect 23612 31426 23668 31428
rect 23612 31374 23614 31426
rect 23614 31374 23666 31426
rect 23666 31374 23668 31426
rect 23612 31372 23668 31374
rect 23772 31426 23828 31428
rect 23772 31374 23774 31426
rect 23774 31374 23826 31426
rect 23826 31374 23828 31426
rect 23772 31372 23828 31374
rect 23932 31426 23988 31428
rect 23932 31374 23934 31426
rect 23934 31374 23986 31426
rect 23986 31374 23988 31426
rect 23932 31372 23988 31374
rect 24092 31426 24148 31428
rect 24092 31374 24094 31426
rect 24094 31374 24146 31426
rect 24146 31374 24148 31426
rect 24092 31372 24148 31374
rect 24252 31426 24308 31428
rect 24252 31374 24254 31426
rect 24254 31374 24306 31426
rect 24306 31374 24308 31426
rect 24252 31372 24308 31374
rect 24412 31426 24468 31428
rect 24412 31374 24414 31426
rect 24414 31374 24466 31426
rect 24466 31374 24468 31426
rect 24412 31372 24468 31374
rect 24572 31426 24628 31428
rect 24572 31374 24574 31426
rect 24574 31374 24626 31426
rect 24626 31374 24628 31426
rect 24572 31372 24628 31374
rect 24732 31426 24788 31428
rect 24732 31374 24734 31426
rect 24734 31374 24786 31426
rect 24786 31374 24788 31426
rect 24732 31372 24788 31374
rect 24892 31426 24948 31428
rect 24892 31374 24894 31426
rect 24894 31374 24946 31426
rect 24946 31374 24948 31426
rect 24892 31372 24948 31374
rect 25052 31426 25108 31428
rect 25052 31374 25054 31426
rect 25054 31374 25106 31426
rect 25106 31374 25108 31426
rect 25052 31372 25108 31374
rect 25212 31426 25268 31428
rect 25212 31374 25214 31426
rect 25214 31374 25266 31426
rect 25266 31374 25268 31426
rect 25212 31372 25268 31374
rect 25372 31426 25428 31428
rect 25372 31374 25374 31426
rect 25374 31374 25426 31426
rect 25426 31374 25428 31426
rect 25372 31372 25428 31374
rect 25532 31426 25588 31428
rect 25532 31374 25534 31426
rect 25534 31374 25586 31426
rect 25586 31374 25588 31426
rect 25532 31372 25588 31374
rect 25692 31426 25748 31428
rect 25692 31374 25694 31426
rect 25694 31374 25746 31426
rect 25746 31374 25748 31426
rect 25692 31372 25748 31374
rect 25852 31426 25908 31428
rect 25852 31374 25854 31426
rect 25854 31374 25906 31426
rect 25906 31374 25908 31426
rect 25852 31372 25908 31374
rect 26012 31426 26068 31428
rect 26012 31374 26014 31426
rect 26014 31374 26066 31426
rect 26066 31374 26068 31426
rect 26012 31372 26068 31374
rect 26172 31426 26228 31428
rect 26172 31374 26174 31426
rect 26174 31374 26226 31426
rect 26226 31374 26228 31426
rect 26172 31372 26228 31374
rect 26332 31426 26388 31428
rect 26332 31374 26334 31426
rect 26334 31374 26386 31426
rect 26386 31374 26388 31426
rect 26332 31372 26388 31374
rect 26492 31426 26548 31428
rect 26492 31374 26494 31426
rect 26494 31374 26546 31426
rect 26546 31374 26548 31426
rect 26492 31372 26548 31374
rect 26652 31426 26708 31428
rect 26652 31374 26654 31426
rect 26654 31374 26706 31426
rect 26706 31374 26708 31426
rect 26652 31372 26708 31374
rect 26812 31426 26868 31428
rect 26812 31374 26814 31426
rect 26814 31374 26866 31426
rect 26866 31374 26868 31426
rect 26812 31372 26868 31374
rect 26972 31426 27028 31428
rect 26972 31374 26974 31426
rect 26974 31374 27026 31426
rect 27026 31374 27028 31426
rect 26972 31372 27028 31374
rect 27132 31426 27188 31428
rect 27132 31374 27134 31426
rect 27134 31374 27186 31426
rect 27186 31374 27188 31426
rect 27132 31372 27188 31374
rect 27292 31426 27348 31428
rect 27292 31374 27294 31426
rect 27294 31374 27346 31426
rect 27346 31374 27348 31426
rect 27292 31372 27348 31374
rect 27452 31426 27508 31428
rect 27452 31374 27454 31426
rect 27454 31374 27506 31426
rect 27506 31374 27508 31426
rect 27452 31372 27508 31374
rect 27612 31426 27668 31428
rect 27612 31374 27614 31426
rect 27614 31374 27666 31426
rect 27666 31374 27668 31426
rect 27612 31372 27668 31374
rect 27772 31426 27828 31428
rect 27772 31374 27774 31426
rect 27774 31374 27826 31426
rect 27826 31374 27828 31426
rect 27772 31372 27828 31374
rect 27932 31426 27988 31428
rect 27932 31374 27934 31426
rect 27934 31374 27986 31426
rect 27986 31374 27988 31426
rect 27932 31372 27988 31374
rect 28092 31426 28148 31428
rect 28092 31374 28094 31426
rect 28094 31374 28146 31426
rect 28146 31374 28148 31426
rect 28092 31372 28148 31374
rect 28252 31426 28308 31428
rect 28252 31374 28254 31426
rect 28254 31374 28306 31426
rect 28306 31374 28308 31426
rect 28252 31372 28308 31374
rect 28412 31426 28468 31428
rect 28412 31374 28414 31426
rect 28414 31374 28466 31426
rect 28466 31374 28468 31426
rect 28412 31372 28468 31374
rect 28572 31426 28628 31428
rect 28572 31374 28574 31426
rect 28574 31374 28626 31426
rect 28626 31374 28628 31426
rect 28572 31372 28628 31374
rect 28732 31426 28788 31428
rect 28732 31374 28734 31426
rect 28734 31374 28786 31426
rect 28786 31374 28788 31426
rect 28732 31372 28788 31374
rect 28892 31426 28948 31428
rect 28892 31374 28894 31426
rect 28894 31374 28946 31426
rect 28946 31374 28948 31426
rect 28892 31372 28948 31374
rect 29052 31426 29108 31428
rect 29052 31374 29054 31426
rect 29054 31374 29106 31426
rect 29106 31374 29108 31426
rect 29052 31372 29108 31374
rect 29212 31426 29268 31428
rect 29212 31374 29214 31426
rect 29214 31374 29266 31426
rect 29266 31374 29268 31426
rect 29212 31372 29268 31374
rect 29372 31426 29428 31428
rect 29372 31374 29374 31426
rect 29374 31374 29426 31426
rect 29426 31374 29428 31426
rect 29372 31372 29428 31374
rect 30492 31372 30548 31428
rect 30812 31372 30868 31428
rect 31132 31372 31188 31428
rect 31452 31372 31508 31428
rect 31772 31372 31828 31428
rect 32092 31372 32148 31428
rect 32412 31372 32468 31428
rect 33532 31426 33588 31428
rect 33532 31374 33534 31426
rect 33534 31374 33586 31426
rect 33586 31374 33588 31426
rect 33532 31372 33588 31374
rect 33692 31426 33748 31428
rect 33692 31374 33694 31426
rect 33694 31374 33746 31426
rect 33746 31374 33748 31426
rect 33692 31372 33748 31374
rect 33852 31426 33908 31428
rect 33852 31374 33854 31426
rect 33854 31374 33906 31426
rect 33906 31374 33908 31426
rect 33852 31372 33908 31374
rect 34012 31426 34068 31428
rect 34012 31374 34014 31426
rect 34014 31374 34066 31426
rect 34066 31374 34068 31426
rect 34012 31372 34068 31374
rect 34172 31426 34228 31428
rect 34172 31374 34174 31426
rect 34174 31374 34226 31426
rect 34226 31374 34228 31426
rect 34172 31372 34228 31374
rect 34332 31426 34388 31428
rect 34332 31374 34334 31426
rect 34334 31374 34386 31426
rect 34386 31374 34388 31426
rect 34332 31372 34388 31374
rect 34492 31426 34548 31428
rect 34492 31374 34494 31426
rect 34494 31374 34546 31426
rect 34546 31374 34548 31426
rect 34492 31372 34548 31374
rect 34652 31426 34708 31428
rect 34652 31374 34654 31426
rect 34654 31374 34706 31426
rect 34706 31374 34708 31426
rect 34652 31372 34708 31374
rect 34812 31426 34868 31428
rect 34812 31374 34814 31426
rect 34814 31374 34866 31426
rect 34866 31374 34868 31426
rect 34812 31372 34868 31374
rect 34972 31426 35028 31428
rect 34972 31374 34974 31426
rect 34974 31374 35026 31426
rect 35026 31374 35028 31426
rect 34972 31372 35028 31374
rect 35132 31426 35188 31428
rect 35132 31374 35134 31426
rect 35134 31374 35186 31426
rect 35186 31374 35188 31426
rect 35132 31372 35188 31374
rect 35292 31426 35348 31428
rect 35292 31374 35294 31426
rect 35294 31374 35346 31426
rect 35346 31374 35348 31426
rect 35292 31372 35348 31374
rect 35452 31426 35508 31428
rect 35452 31374 35454 31426
rect 35454 31374 35506 31426
rect 35506 31374 35508 31426
rect 35452 31372 35508 31374
rect 35612 31426 35668 31428
rect 35612 31374 35614 31426
rect 35614 31374 35666 31426
rect 35666 31374 35668 31426
rect 35612 31372 35668 31374
rect 35772 31426 35828 31428
rect 35772 31374 35774 31426
rect 35774 31374 35826 31426
rect 35826 31374 35828 31426
rect 35772 31372 35828 31374
rect 35932 31426 35988 31428
rect 35932 31374 35934 31426
rect 35934 31374 35986 31426
rect 35986 31374 35988 31426
rect 35932 31372 35988 31374
rect 36092 31426 36148 31428
rect 36092 31374 36094 31426
rect 36094 31374 36146 31426
rect 36146 31374 36148 31426
rect 36092 31372 36148 31374
rect 36252 31426 36308 31428
rect 36252 31374 36254 31426
rect 36254 31374 36306 31426
rect 36306 31374 36308 31426
rect 36252 31372 36308 31374
rect 36412 31426 36468 31428
rect 36412 31374 36414 31426
rect 36414 31374 36466 31426
rect 36466 31374 36468 31426
rect 36412 31372 36468 31374
rect 36572 31426 36628 31428
rect 36572 31374 36574 31426
rect 36574 31374 36626 31426
rect 36626 31374 36628 31426
rect 36572 31372 36628 31374
rect 36732 31426 36788 31428
rect 36732 31374 36734 31426
rect 36734 31374 36786 31426
rect 36786 31374 36788 31426
rect 36732 31372 36788 31374
rect 36892 31426 36948 31428
rect 36892 31374 36894 31426
rect 36894 31374 36946 31426
rect 36946 31374 36948 31426
rect 36892 31372 36948 31374
rect 37052 31426 37108 31428
rect 37052 31374 37054 31426
rect 37054 31374 37106 31426
rect 37106 31374 37108 31426
rect 37052 31372 37108 31374
rect 37212 31426 37268 31428
rect 37212 31374 37214 31426
rect 37214 31374 37266 31426
rect 37266 31374 37268 31426
rect 37212 31372 37268 31374
rect 37372 31426 37428 31428
rect 37372 31374 37374 31426
rect 37374 31374 37426 31426
rect 37426 31374 37428 31426
rect 37372 31372 37428 31374
rect 37532 31426 37588 31428
rect 37532 31374 37534 31426
rect 37534 31374 37586 31426
rect 37586 31374 37588 31426
rect 37532 31372 37588 31374
rect 37692 31426 37748 31428
rect 37692 31374 37694 31426
rect 37694 31374 37746 31426
rect 37746 31374 37748 31426
rect 37692 31372 37748 31374
rect 37852 31426 37908 31428
rect 37852 31374 37854 31426
rect 37854 31374 37906 31426
rect 37906 31374 37908 31426
rect 37852 31372 37908 31374
rect 38012 31426 38068 31428
rect 38012 31374 38014 31426
rect 38014 31374 38066 31426
rect 38066 31374 38068 31426
rect 38012 31372 38068 31374
rect 38172 31426 38228 31428
rect 38172 31374 38174 31426
rect 38174 31374 38226 31426
rect 38226 31374 38228 31426
rect 38172 31372 38228 31374
rect 38332 31426 38388 31428
rect 38332 31374 38334 31426
rect 38334 31374 38386 31426
rect 38386 31374 38388 31426
rect 38332 31372 38388 31374
rect 38492 31426 38548 31428
rect 38492 31374 38494 31426
rect 38494 31374 38546 31426
rect 38546 31374 38548 31426
rect 38492 31372 38548 31374
rect 38652 31426 38708 31428
rect 38652 31374 38654 31426
rect 38654 31374 38706 31426
rect 38706 31374 38708 31426
rect 38652 31372 38708 31374
rect 38812 31426 38868 31428
rect 38812 31374 38814 31426
rect 38814 31374 38866 31426
rect 38866 31374 38868 31426
rect 38812 31372 38868 31374
rect 38972 31426 39028 31428
rect 38972 31374 38974 31426
rect 38974 31374 39026 31426
rect 39026 31374 39028 31426
rect 38972 31372 39028 31374
rect 39132 31426 39188 31428
rect 39132 31374 39134 31426
rect 39134 31374 39186 31426
rect 39186 31374 39188 31426
rect 39132 31372 39188 31374
rect 39292 31426 39348 31428
rect 39292 31374 39294 31426
rect 39294 31374 39346 31426
rect 39346 31374 39348 31426
rect 39292 31372 39348 31374
rect 39452 31426 39508 31428
rect 39452 31374 39454 31426
rect 39454 31374 39506 31426
rect 39506 31374 39508 31426
rect 39452 31372 39508 31374
rect 39612 31426 39668 31428
rect 39612 31374 39614 31426
rect 39614 31374 39666 31426
rect 39666 31374 39668 31426
rect 39612 31372 39668 31374
rect 39772 31426 39828 31428
rect 39772 31374 39774 31426
rect 39774 31374 39826 31426
rect 39826 31374 39828 31426
rect 39772 31372 39828 31374
rect 39932 31426 39988 31428
rect 39932 31374 39934 31426
rect 39934 31374 39986 31426
rect 39986 31374 39988 31426
rect 39932 31372 39988 31374
rect 40092 31426 40148 31428
rect 40092 31374 40094 31426
rect 40094 31374 40146 31426
rect 40146 31374 40148 31426
rect 40092 31372 40148 31374
rect 40252 31426 40308 31428
rect 40252 31374 40254 31426
rect 40254 31374 40306 31426
rect 40306 31374 40308 31426
rect 40252 31372 40308 31374
rect 40412 31426 40468 31428
rect 40412 31374 40414 31426
rect 40414 31374 40466 31426
rect 40466 31374 40468 31426
rect 40412 31372 40468 31374
rect 40572 31426 40628 31428
rect 40572 31374 40574 31426
rect 40574 31374 40626 31426
rect 40626 31374 40628 31426
rect 40572 31372 40628 31374
rect 40732 31426 40788 31428
rect 40732 31374 40734 31426
rect 40734 31374 40786 31426
rect 40786 31374 40788 31426
rect 40732 31372 40788 31374
rect 40892 31426 40948 31428
rect 40892 31374 40894 31426
rect 40894 31374 40946 31426
rect 40946 31374 40948 31426
rect 40892 31372 40948 31374
rect 41052 31426 41108 31428
rect 41052 31374 41054 31426
rect 41054 31374 41106 31426
rect 41106 31374 41108 31426
rect 41052 31372 41108 31374
rect 41212 31426 41268 31428
rect 41212 31374 41214 31426
rect 41214 31374 41266 31426
rect 41266 31374 41268 31426
rect 41212 31372 41268 31374
rect 41372 31426 41428 31428
rect 41372 31374 41374 31426
rect 41374 31374 41426 31426
rect 41426 31374 41428 31426
rect 41372 31372 41428 31374
rect 41532 31426 41588 31428
rect 41532 31374 41534 31426
rect 41534 31374 41586 31426
rect 41586 31374 41588 31426
rect 41532 31372 41588 31374
rect 41692 31426 41748 31428
rect 41692 31374 41694 31426
rect 41694 31374 41746 31426
rect 41746 31374 41748 31426
rect 41692 31372 41748 31374
rect 41852 31426 41908 31428
rect 41852 31374 41854 31426
rect 41854 31374 41906 31426
rect 41906 31374 41908 31426
rect 41852 31372 41908 31374
rect 10572 31212 10628 31268
rect 21132 31212 21188 31268
rect 31292 31212 31348 31268
rect 12 31106 68 31108
rect 12 31054 14 31106
rect 14 31054 66 31106
rect 66 31054 68 31106
rect 12 31052 68 31054
rect 172 31106 228 31108
rect 172 31054 174 31106
rect 174 31054 226 31106
rect 226 31054 228 31106
rect 172 31052 228 31054
rect 332 31106 388 31108
rect 332 31054 334 31106
rect 334 31054 386 31106
rect 386 31054 388 31106
rect 332 31052 388 31054
rect 492 31106 548 31108
rect 492 31054 494 31106
rect 494 31054 546 31106
rect 546 31054 548 31106
rect 492 31052 548 31054
rect 652 31106 708 31108
rect 652 31054 654 31106
rect 654 31054 706 31106
rect 706 31054 708 31106
rect 652 31052 708 31054
rect 812 31106 868 31108
rect 812 31054 814 31106
rect 814 31054 866 31106
rect 866 31054 868 31106
rect 812 31052 868 31054
rect 972 31106 1028 31108
rect 972 31054 974 31106
rect 974 31054 1026 31106
rect 1026 31054 1028 31106
rect 972 31052 1028 31054
rect 1132 31106 1188 31108
rect 1132 31054 1134 31106
rect 1134 31054 1186 31106
rect 1186 31054 1188 31106
rect 1132 31052 1188 31054
rect 1292 31106 1348 31108
rect 1292 31054 1294 31106
rect 1294 31054 1346 31106
rect 1346 31054 1348 31106
rect 1292 31052 1348 31054
rect 1452 31106 1508 31108
rect 1452 31054 1454 31106
rect 1454 31054 1506 31106
rect 1506 31054 1508 31106
rect 1452 31052 1508 31054
rect 1612 31106 1668 31108
rect 1612 31054 1614 31106
rect 1614 31054 1666 31106
rect 1666 31054 1668 31106
rect 1612 31052 1668 31054
rect 1772 31106 1828 31108
rect 1772 31054 1774 31106
rect 1774 31054 1826 31106
rect 1826 31054 1828 31106
rect 1772 31052 1828 31054
rect 1932 31106 1988 31108
rect 1932 31054 1934 31106
rect 1934 31054 1986 31106
rect 1986 31054 1988 31106
rect 1932 31052 1988 31054
rect 2092 31106 2148 31108
rect 2092 31054 2094 31106
rect 2094 31054 2146 31106
rect 2146 31054 2148 31106
rect 2092 31052 2148 31054
rect 2252 31106 2308 31108
rect 2252 31054 2254 31106
rect 2254 31054 2306 31106
rect 2306 31054 2308 31106
rect 2252 31052 2308 31054
rect 2412 31106 2468 31108
rect 2412 31054 2414 31106
rect 2414 31054 2466 31106
rect 2466 31054 2468 31106
rect 2412 31052 2468 31054
rect 2572 31106 2628 31108
rect 2572 31054 2574 31106
rect 2574 31054 2626 31106
rect 2626 31054 2628 31106
rect 2572 31052 2628 31054
rect 2732 31106 2788 31108
rect 2732 31054 2734 31106
rect 2734 31054 2786 31106
rect 2786 31054 2788 31106
rect 2732 31052 2788 31054
rect 2892 31106 2948 31108
rect 2892 31054 2894 31106
rect 2894 31054 2946 31106
rect 2946 31054 2948 31106
rect 2892 31052 2948 31054
rect 3052 31106 3108 31108
rect 3052 31054 3054 31106
rect 3054 31054 3106 31106
rect 3106 31054 3108 31106
rect 3052 31052 3108 31054
rect 3212 31106 3268 31108
rect 3212 31054 3214 31106
rect 3214 31054 3266 31106
rect 3266 31054 3268 31106
rect 3212 31052 3268 31054
rect 3372 31106 3428 31108
rect 3372 31054 3374 31106
rect 3374 31054 3426 31106
rect 3426 31054 3428 31106
rect 3372 31052 3428 31054
rect 3532 31106 3588 31108
rect 3532 31054 3534 31106
rect 3534 31054 3586 31106
rect 3586 31054 3588 31106
rect 3532 31052 3588 31054
rect 3692 31106 3748 31108
rect 3692 31054 3694 31106
rect 3694 31054 3746 31106
rect 3746 31054 3748 31106
rect 3692 31052 3748 31054
rect 3852 31106 3908 31108
rect 3852 31054 3854 31106
rect 3854 31054 3906 31106
rect 3906 31054 3908 31106
rect 3852 31052 3908 31054
rect 4012 31106 4068 31108
rect 4012 31054 4014 31106
rect 4014 31054 4066 31106
rect 4066 31054 4068 31106
rect 4012 31052 4068 31054
rect 4172 31106 4228 31108
rect 4172 31054 4174 31106
rect 4174 31054 4226 31106
rect 4226 31054 4228 31106
rect 4172 31052 4228 31054
rect 4332 31106 4388 31108
rect 4332 31054 4334 31106
rect 4334 31054 4386 31106
rect 4386 31054 4388 31106
rect 4332 31052 4388 31054
rect 4492 31106 4548 31108
rect 4492 31054 4494 31106
rect 4494 31054 4546 31106
rect 4546 31054 4548 31106
rect 4492 31052 4548 31054
rect 4652 31106 4708 31108
rect 4652 31054 4654 31106
rect 4654 31054 4706 31106
rect 4706 31054 4708 31106
rect 4652 31052 4708 31054
rect 4812 31106 4868 31108
rect 4812 31054 4814 31106
rect 4814 31054 4866 31106
rect 4866 31054 4868 31106
rect 4812 31052 4868 31054
rect 4972 31106 5028 31108
rect 4972 31054 4974 31106
rect 4974 31054 5026 31106
rect 5026 31054 5028 31106
rect 4972 31052 5028 31054
rect 5132 31106 5188 31108
rect 5132 31054 5134 31106
rect 5134 31054 5186 31106
rect 5186 31054 5188 31106
rect 5132 31052 5188 31054
rect 5292 31106 5348 31108
rect 5292 31054 5294 31106
rect 5294 31054 5346 31106
rect 5346 31054 5348 31106
rect 5292 31052 5348 31054
rect 5452 31106 5508 31108
rect 5452 31054 5454 31106
rect 5454 31054 5506 31106
rect 5506 31054 5508 31106
rect 5452 31052 5508 31054
rect 5612 31106 5668 31108
rect 5612 31054 5614 31106
rect 5614 31054 5666 31106
rect 5666 31054 5668 31106
rect 5612 31052 5668 31054
rect 5772 31106 5828 31108
rect 5772 31054 5774 31106
rect 5774 31054 5826 31106
rect 5826 31054 5828 31106
rect 5772 31052 5828 31054
rect 5932 31106 5988 31108
rect 5932 31054 5934 31106
rect 5934 31054 5986 31106
rect 5986 31054 5988 31106
rect 5932 31052 5988 31054
rect 6092 31106 6148 31108
rect 6092 31054 6094 31106
rect 6094 31054 6146 31106
rect 6146 31054 6148 31106
rect 6092 31052 6148 31054
rect 6252 31106 6308 31108
rect 6252 31054 6254 31106
rect 6254 31054 6306 31106
rect 6306 31054 6308 31106
rect 6252 31052 6308 31054
rect 6412 31106 6468 31108
rect 6412 31054 6414 31106
rect 6414 31054 6466 31106
rect 6466 31054 6468 31106
rect 6412 31052 6468 31054
rect 6572 31106 6628 31108
rect 6572 31054 6574 31106
rect 6574 31054 6626 31106
rect 6626 31054 6628 31106
rect 6572 31052 6628 31054
rect 6732 31106 6788 31108
rect 6732 31054 6734 31106
rect 6734 31054 6786 31106
rect 6786 31054 6788 31106
rect 6732 31052 6788 31054
rect 6892 31106 6948 31108
rect 6892 31054 6894 31106
rect 6894 31054 6946 31106
rect 6946 31054 6948 31106
rect 6892 31052 6948 31054
rect 7052 31106 7108 31108
rect 7052 31054 7054 31106
rect 7054 31054 7106 31106
rect 7106 31054 7108 31106
rect 7052 31052 7108 31054
rect 7212 31106 7268 31108
rect 7212 31054 7214 31106
rect 7214 31054 7266 31106
rect 7266 31054 7268 31106
rect 7212 31052 7268 31054
rect 7372 31106 7428 31108
rect 7372 31054 7374 31106
rect 7374 31054 7426 31106
rect 7426 31054 7428 31106
rect 7372 31052 7428 31054
rect 7532 31106 7588 31108
rect 7532 31054 7534 31106
rect 7534 31054 7586 31106
rect 7586 31054 7588 31106
rect 7532 31052 7588 31054
rect 7692 31106 7748 31108
rect 7692 31054 7694 31106
rect 7694 31054 7746 31106
rect 7746 31054 7748 31106
rect 7692 31052 7748 31054
rect 7852 31106 7908 31108
rect 7852 31054 7854 31106
rect 7854 31054 7906 31106
rect 7906 31054 7908 31106
rect 7852 31052 7908 31054
rect 8012 31106 8068 31108
rect 8012 31054 8014 31106
rect 8014 31054 8066 31106
rect 8066 31054 8068 31106
rect 8012 31052 8068 31054
rect 8172 31106 8228 31108
rect 8172 31054 8174 31106
rect 8174 31054 8226 31106
rect 8226 31054 8228 31106
rect 8172 31052 8228 31054
rect 8332 31106 8388 31108
rect 8332 31054 8334 31106
rect 8334 31054 8386 31106
rect 8386 31054 8388 31106
rect 8332 31052 8388 31054
rect 9452 31052 9508 31108
rect 9772 31052 9828 31108
rect 10092 31052 10148 31108
rect 10412 31052 10468 31108
rect 10732 31052 10788 31108
rect 11052 31052 11108 31108
rect 11372 31052 11428 31108
rect 12492 31106 12548 31108
rect 12492 31054 12494 31106
rect 12494 31054 12546 31106
rect 12546 31054 12548 31106
rect 12492 31052 12548 31054
rect 12652 31106 12708 31108
rect 12652 31054 12654 31106
rect 12654 31054 12706 31106
rect 12706 31054 12708 31106
rect 12652 31052 12708 31054
rect 12812 31106 12868 31108
rect 12812 31054 12814 31106
rect 12814 31054 12866 31106
rect 12866 31054 12868 31106
rect 12812 31052 12868 31054
rect 12972 31106 13028 31108
rect 12972 31054 12974 31106
rect 12974 31054 13026 31106
rect 13026 31054 13028 31106
rect 12972 31052 13028 31054
rect 13132 31106 13188 31108
rect 13132 31054 13134 31106
rect 13134 31054 13186 31106
rect 13186 31054 13188 31106
rect 13132 31052 13188 31054
rect 13292 31106 13348 31108
rect 13292 31054 13294 31106
rect 13294 31054 13346 31106
rect 13346 31054 13348 31106
rect 13292 31052 13348 31054
rect 13452 31106 13508 31108
rect 13452 31054 13454 31106
rect 13454 31054 13506 31106
rect 13506 31054 13508 31106
rect 13452 31052 13508 31054
rect 13612 31106 13668 31108
rect 13612 31054 13614 31106
rect 13614 31054 13666 31106
rect 13666 31054 13668 31106
rect 13612 31052 13668 31054
rect 13772 31106 13828 31108
rect 13772 31054 13774 31106
rect 13774 31054 13826 31106
rect 13826 31054 13828 31106
rect 13772 31052 13828 31054
rect 13932 31106 13988 31108
rect 13932 31054 13934 31106
rect 13934 31054 13986 31106
rect 13986 31054 13988 31106
rect 13932 31052 13988 31054
rect 14092 31106 14148 31108
rect 14092 31054 14094 31106
rect 14094 31054 14146 31106
rect 14146 31054 14148 31106
rect 14092 31052 14148 31054
rect 14252 31106 14308 31108
rect 14252 31054 14254 31106
rect 14254 31054 14306 31106
rect 14306 31054 14308 31106
rect 14252 31052 14308 31054
rect 14412 31106 14468 31108
rect 14412 31054 14414 31106
rect 14414 31054 14466 31106
rect 14466 31054 14468 31106
rect 14412 31052 14468 31054
rect 14572 31106 14628 31108
rect 14572 31054 14574 31106
rect 14574 31054 14626 31106
rect 14626 31054 14628 31106
rect 14572 31052 14628 31054
rect 14732 31106 14788 31108
rect 14732 31054 14734 31106
rect 14734 31054 14786 31106
rect 14786 31054 14788 31106
rect 14732 31052 14788 31054
rect 14892 31106 14948 31108
rect 14892 31054 14894 31106
rect 14894 31054 14946 31106
rect 14946 31054 14948 31106
rect 14892 31052 14948 31054
rect 15052 31106 15108 31108
rect 15052 31054 15054 31106
rect 15054 31054 15106 31106
rect 15106 31054 15108 31106
rect 15052 31052 15108 31054
rect 15212 31106 15268 31108
rect 15212 31054 15214 31106
rect 15214 31054 15266 31106
rect 15266 31054 15268 31106
rect 15212 31052 15268 31054
rect 15372 31106 15428 31108
rect 15372 31054 15374 31106
rect 15374 31054 15426 31106
rect 15426 31054 15428 31106
rect 15372 31052 15428 31054
rect 15532 31106 15588 31108
rect 15532 31054 15534 31106
rect 15534 31054 15586 31106
rect 15586 31054 15588 31106
rect 15532 31052 15588 31054
rect 15692 31106 15748 31108
rect 15692 31054 15694 31106
rect 15694 31054 15746 31106
rect 15746 31054 15748 31106
rect 15692 31052 15748 31054
rect 15852 31106 15908 31108
rect 15852 31054 15854 31106
rect 15854 31054 15906 31106
rect 15906 31054 15908 31106
rect 15852 31052 15908 31054
rect 16012 31106 16068 31108
rect 16012 31054 16014 31106
rect 16014 31054 16066 31106
rect 16066 31054 16068 31106
rect 16012 31052 16068 31054
rect 16172 31106 16228 31108
rect 16172 31054 16174 31106
rect 16174 31054 16226 31106
rect 16226 31054 16228 31106
rect 16172 31052 16228 31054
rect 16332 31106 16388 31108
rect 16332 31054 16334 31106
rect 16334 31054 16386 31106
rect 16386 31054 16388 31106
rect 16332 31052 16388 31054
rect 16492 31106 16548 31108
rect 16492 31054 16494 31106
rect 16494 31054 16546 31106
rect 16546 31054 16548 31106
rect 16492 31052 16548 31054
rect 16652 31106 16708 31108
rect 16652 31054 16654 31106
rect 16654 31054 16706 31106
rect 16706 31054 16708 31106
rect 16652 31052 16708 31054
rect 16812 31106 16868 31108
rect 16812 31054 16814 31106
rect 16814 31054 16866 31106
rect 16866 31054 16868 31106
rect 16812 31052 16868 31054
rect 16972 31106 17028 31108
rect 16972 31054 16974 31106
rect 16974 31054 17026 31106
rect 17026 31054 17028 31106
rect 16972 31052 17028 31054
rect 17132 31106 17188 31108
rect 17132 31054 17134 31106
rect 17134 31054 17186 31106
rect 17186 31054 17188 31106
rect 17132 31052 17188 31054
rect 17292 31106 17348 31108
rect 17292 31054 17294 31106
rect 17294 31054 17346 31106
rect 17346 31054 17348 31106
rect 17292 31052 17348 31054
rect 17452 31106 17508 31108
rect 17452 31054 17454 31106
rect 17454 31054 17506 31106
rect 17506 31054 17508 31106
rect 17452 31052 17508 31054
rect 17612 31106 17668 31108
rect 17612 31054 17614 31106
rect 17614 31054 17666 31106
rect 17666 31054 17668 31106
rect 17612 31052 17668 31054
rect 17772 31106 17828 31108
rect 17772 31054 17774 31106
rect 17774 31054 17826 31106
rect 17826 31054 17828 31106
rect 17772 31052 17828 31054
rect 17932 31106 17988 31108
rect 17932 31054 17934 31106
rect 17934 31054 17986 31106
rect 17986 31054 17988 31106
rect 17932 31052 17988 31054
rect 18092 31106 18148 31108
rect 18092 31054 18094 31106
rect 18094 31054 18146 31106
rect 18146 31054 18148 31106
rect 18092 31052 18148 31054
rect 18252 31106 18308 31108
rect 18252 31054 18254 31106
rect 18254 31054 18306 31106
rect 18306 31054 18308 31106
rect 18252 31052 18308 31054
rect 18412 31106 18468 31108
rect 18412 31054 18414 31106
rect 18414 31054 18466 31106
rect 18466 31054 18468 31106
rect 18412 31052 18468 31054
rect 18572 31106 18628 31108
rect 18572 31054 18574 31106
rect 18574 31054 18626 31106
rect 18626 31054 18628 31106
rect 18572 31052 18628 31054
rect 18732 31106 18788 31108
rect 18732 31054 18734 31106
rect 18734 31054 18786 31106
rect 18786 31054 18788 31106
rect 18732 31052 18788 31054
rect 18892 31106 18948 31108
rect 18892 31054 18894 31106
rect 18894 31054 18946 31106
rect 18946 31054 18948 31106
rect 18892 31052 18948 31054
rect 20012 31052 20068 31108
rect 20332 31052 20388 31108
rect 20652 31052 20708 31108
rect 20972 31052 21028 31108
rect 21292 31052 21348 31108
rect 21612 31052 21668 31108
rect 21932 31052 21988 31108
rect 23132 31106 23188 31108
rect 23132 31054 23134 31106
rect 23134 31054 23186 31106
rect 23186 31054 23188 31106
rect 23132 31052 23188 31054
rect 23292 31106 23348 31108
rect 23292 31054 23294 31106
rect 23294 31054 23346 31106
rect 23346 31054 23348 31106
rect 23292 31052 23348 31054
rect 23452 31106 23508 31108
rect 23452 31054 23454 31106
rect 23454 31054 23506 31106
rect 23506 31054 23508 31106
rect 23452 31052 23508 31054
rect 23612 31106 23668 31108
rect 23612 31054 23614 31106
rect 23614 31054 23666 31106
rect 23666 31054 23668 31106
rect 23612 31052 23668 31054
rect 23772 31106 23828 31108
rect 23772 31054 23774 31106
rect 23774 31054 23826 31106
rect 23826 31054 23828 31106
rect 23772 31052 23828 31054
rect 23932 31106 23988 31108
rect 23932 31054 23934 31106
rect 23934 31054 23986 31106
rect 23986 31054 23988 31106
rect 23932 31052 23988 31054
rect 24092 31106 24148 31108
rect 24092 31054 24094 31106
rect 24094 31054 24146 31106
rect 24146 31054 24148 31106
rect 24092 31052 24148 31054
rect 24252 31106 24308 31108
rect 24252 31054 24254 31106
rect 24254 31054 24306 31106
rect 24306 31054 24308 31106
rect 24252 31052 24308 31054
rect 24412 31106 24468 31108
rect 24412 31054 24414 31106
rect 24414 31054 24466 31106
rect 24466 31054 24468 31106
rect 24412 31052 24468 31054
rect 24572 31106 24628 31108
rect 24572 31054 24574 31106
rect 24574 31054 24626 31106
rect 24626 31054 24628 31106
rect 24572 31052 24628 31054
rect 24732 31106 24788 31108
rect 24732 31054 24734 31106
rect 24734 31054 24786 31106
rect 24786 31054 24788 31106
rect 24732 31052 24788 31054
rect 24892 31106 24948 31108
rect 24892 31054 24894 31106
rect 24894 31054 24946 31106
rect 24946 31054 24948 31106
rect 24892 31052 24948 31054
rect 25052 31106 25108 31108
rect 25052 31054 25054 31106
rect 25054 31054 25106 31106
rect 25106 31054 25108 31106
rect 25052 31052 25108 31054
rect 25212 31106 25268 31108
rect 25212 31054 25214 31106
rect 25214 31054 25266 31106
rect 25266 31054 25268 31106
rect 25212 31052 25268 31054
rect 25372 31106 25428 31108
rect 25372 31054 25374 31106
rect 25374 31054 25426 31106
rect 25426 31054 25428 31106
rect 25372 31052 25428 31054
rect 25532 31106 25588 31108
rect 25532 31054 25534 31106
rect 25534 31054 25586 31106
rect 25586 31054 25588 31106
rect 25532 31052 25588 31054
rect 25692 31106 25748 31108
rect 25692 31054 25694 31106
rect 25694 31054 25746 31106
rect 25746 31054 25748 31106
rect 25692 31052 25748 31054
rect 25852 31106 25908 31108
rect 25852 31054 25854 31106
rect 25854 31054 25906 31106
rect 25906 31054 25908 31106
rect 25852 31052 25908 31054
rect 26012 31106 26068 31108
rect 26012 31054 26014 31106
rect 26014 31054 26066 31106
rect 26066 31054 26068 31106
rect 26012 31052 26068 31054
rect 26172 31106 26228 31108
rect 26172 31054 26174 31106
rect 26174 31054 26226 31106
rect 26226 31054 26228 31106
rect 26172 31052 26228 31054
rect 26332 31106 26388 31108
rect 26332 31054 26334 31106
rect 26334 31054 26386 31106
rect 26386 31054 26388 31106
rect 26332 31052 26388 31054
rect 26492 31106 26548 31108
rect 26492 31054 26494 31106
rect 26494 31054 26546 31106
rect 26546 31054 26548 31106
rect 26492 31052 26548 31054
rect 26652 31106 26708 31108
rect 26652 31054 26654 31106
rect 26654 31054 26706 31106
rect 26706 31054 26708 31106
rect 26652 31052 26708 31054
rect 26812 31106 26868 31108
rect 26812 31054 26814 31106
rect 26814 31054 26866 31106
rect 26866 31054 26868 31106
rect 26812 31052 26868 31054
rect 26972 31106 27028 31108
rect 26972 31054 26974 31106
rect 26974 31054 27026 31106
rect 27026 31054 27028 31106
rect 26972 31052 27028 31054
rect 27132 31106 27188 31108
rect 27132 31054 27134 31106
rect 27134 31054 27186 31106
rect 27186 31054 27188 31106
rect 27132 31052 27188 31054
rect 27292 31106 27348 31108
rect 27292 31054 27294 31106
rect 27294 31054 27346 31106
rect 27346 31054 27348 31106
rect 27292 31052 27348 31054
rect 27452 31106 27508 31108
rect 27452 31054 27454 31106
rect 27454 31054 27506 31106
rect 27506 31054 27508 31106
rect 27452 31052 27508 31054
rect 27612 31106 27668 31108
rect 27612 31054 27614 31106
rect 27614 31054 27666 31106
rect 27666 31054 27668 31106
rect 27612 31052 27668 31054
rect 27772 31106 27828 31108
rect 27772 31054 27774 31106
rect 27774 31054 27826 31106
rect 27826 31054 27828 31106
rect 27772 31052 27828 31054
rect 27932 31106 27988 31108
rect 27932 31054 27934 31106
rect 27934 31054 27986 31106
rect 27986 31054 27988 31106
rect 27932 31052 27988 31054
rect 28092 31106 28148 31108
rect 28092 31054 28094 31106
rect 28094 31054 28146 31106
rect 28146 31054 28148 31106
rect 28092 31052 28148 31054
rect 28252 31106 28308 31108
rect 28252 31054 28254 31106
rect 28254 31054 28306 31106
rect 28306 31054 28308 31106
rect 28252 31052 28308 31054
rect 28412 31106 28468 31108
rect 28412 31054 28414 31106
rect 28414 31054 28466 31106
rect 28466 31054 28468 31106
rect 28412 31052 28468 31054
rect 28572 31106 28628 31108
rect 28572 31054 28574 31106
rect 28574 31054 28626 31106
rect 28626 31054 28628 31106
rect 28572 31052 28628 31054
rect 28732 31106 28788 31108
rect 28732 31054 28734 31106
rect 28734 31054 28786 31106
rect 28786 31054 28788 31106
rect 28732 31052 28788 31054
rect 28892 31106 28948 31108
rect 28892 31054 28894 31106
rect 28894 31054 28946 31106
rect 28946 31054 28948 31106
rect 28892 31052 28948 31054
rect 29052 31106 29108 31108
rect 29052 31054 29054 31106
rect 29054 31054 29106 31106
rect 29106 31054 29108 31106
rect 29052 31052 29108 31054
rect 29212 31106 29268 31108
rect 29212 31054 29214 31106
rect 29214 31054 29266 31106
rect 29266 31054 29268 31106
rect 29212 31052 29268 31054
rect 29372 31106 29428 31108
rect 29372 31054 29374 31106
rect 29374 31054 29426 31106
rect 29426 31054 29428 31106
rect 29372 31052 29428 31054
rect 30492 31052 30548 31108
rect 30812 31052 30868 31108
rect 31132 31052 31188 31108
rect 31452 31052 31508 31108
rect 31772 31052 31828 31108
rect 32092 31052 32148 31108
rect 32412 31052 32468 31108
rect 33532 31106 33588 31108
rect 33532 31054 33534 31106
rect 33534 31054 33586 31106
rect 33586 31054 33588 31106
rect 33532 31052 33588 31054
rect 33692 31106 33748 31108
rect 33692 31054 33694 31106
rect 33694 31054 33746 31106
rect 33746 31054 33748 31106
rect 33692 31052 33748 31054
rect 33852 31106 33908 31108
rect 33852 31054 33854 31106
rect 33854 31054 33906 31106
rect 33906 31054 33908 31106
rect 33852 31052 33908 31054
rect 34012 31106 34068 31108
rect 34012 31054 34014 31106
rect 34014 31054 34066 31106
rect 34066 31054 34068 31106
rect 34012 31052 34068 31054
rect 34172 31106 34228 31108
rect 34172 31054 34174 31106
rect 34174 31054 34226 31106
rect 34226 31054 34228 31106
rect 34172 31052 34228 31054
rect 34332 31106 34388 31108
rect 34332 31054 34334 31106
rect 34334 31054 34386 31106
rect 34386 31054 34388 31106
rect 34332 31052 34388 31054
rect 34492 31106 34548 31108
rect 34492 31054 34494 31106
rect 34494 31054 34546 31106
rect 34546 31054 34548 31106
rect 34492 31052 34548 31054
rect 34652 31106 34708 31108
rect 34652 31054 34654 31106
rect 34654 31054 34706 31106
rect 34706 31054 34708 31106
rect 34652 31052 34708 31054
rect 34812 31106 34868 31108
rect 34812 31054 34814 31106
rect 34814 31054 34866 31106
rect 34866 31054 34868 31106
rect 34812 31052 34868 31054
rect 34972 31106 35028 31108
rect 34972 31054 34974 31106
rect 34974 31054 35026 31106
rect 35026 31054 35028 31106
rect 34972 31052 35028 31054
rect 35132 31106 35188 31108
rect 35132 31054 35134 31106
rect 35134 31054 35186 31106
rect 35186 31054 35188 31106
rect 35132 31052 35188 31054
rect 35292 31106 35348 31108
rect 35292 31054 35294 31106
rect 35294 31054 35346 31106
rect 35346 31054 35348 31106
rect 35292 31052 35348 31054
rect 35452 31106 35508 31108
rect 35452 31054 35454 31106
rect 35454 31054 35506 31106
rect 35506 31054 35508 31106
rect 35452 31052 35508 31054
rect 35612 31106 35668 31108
rect 35612 31054 35614 31106
rect 35614 31054 35666 31106
rect 35666 31054 35668 31106
rect 35612 31052 35668 31054
rect 35772 31106 35828 31108
rect 35772 31054 35774 31106
rect 35774 31054 35826 31106
rect 35826 31054 35828 31106
rect 35772 31052 35828 31054
rect 35932 31106 35988 31108
rect 35932 31054 35934 31106
rect 35934 31054 35986 31106
rect 35986 31054 35988 31106
rect 35932 31052 35988 31054
rect 36092 31106 36148 31108
rect 36092 31054 36094 31106
rect 36094 31054 36146 31106
rect 36146 31054 36148 31106
rect 36092 31052 36148 31054
rect 36252 31106 36308 31108
rect 36252 31054 36254 31106
rect 36254 31054 36306 31106
rect 36306 31054 36308 31106
rect 36252 31052 36308 31054
rect 36412 31106 36468 31108
rect 36412 31054 36414 31106
rect 36414 31054 36466 31106
rect 36466 31054 36468 31106
rect 36412 31052 36468 31054
rect 36572 31106 36628 31108
rect 36572 31054 36574 31106
rect 36574 31054 36626 31106
rect 36626 31054 36628 31106
rect 36572 31052 36628 31054
rect 36732 31106 36788 31108
rect 36732 31054 36734 31106
rect 36734 31054 36786 31106
rect 36786 31054 36788 31106
rect 36732 31052 36788 31054
rect 36892 31106 36948 31108
rect 36892 31054 36894 31106
rect 36894 31054 36946 31106
rect 36946 31054 36948 31106
rect 36892 31052 36948 31054
rect 37052 31106 37108 31108
rect 37052 31054 37054 31106
rect 37054 31054 37106 31106
rect 37106 31054 37108 31106
rect 37052 31052 37108 31054
rect 37212 31106 37268 31108
rect 37212 31054 37214 31106
rect 37214 31054 37266 31106
rect 37266 31054 37268 31106
rect 37212 31052 37268 31054
rect 37372 31106 37428 31108
rect 37372 31054 37374 31106
rect 37374 31054 37426 31106
rect 37426 31054 37428 31106
rect 37372 31052 37428 31054
rect 37532 31106 37588 31108
rect 37532 31054 37534 31106
rect 37534 31054 37586 31106
rect 37586 31054 37588 31106
rect 37532 31052 37588 31054
rect 37692 31106 37748 31108
rect 37692 31054 37694 31106
rect 37694 31054 37746 31106
rect 37746 31054 37748 31106
rect 37692 31052 37748 31054
rect 37852 31106 37908 31108
rect 37852 31054 37854 31106
rect 37854 31054 37906 31106
rect 37906 31054 37908 31106
rect 37852 31052 37908 31054
rect 38012 31106 38068 31108
rect 38012 31054 38014 31106
rect 38014 31054 38066 31106
rect 38066 31054 38068 31106
rect 38012 31052 38068 31054
rect 38172 31106 38228 31108
rect 38172 31054 38174 31106
rect 38174 31054 38226 31106
rect 38226 31054 38228 31106
rect 38172 31052 38228 31054
rect 38332 31106 38388 31108
rect 38332 31054 38334 31106
rect 38334 31054 38386 31106
rect 38386 31054 38388 31106
rect 38332 31052 38388 31054
rect 38492 31106 38548 31108
rect 38492 31054 38494 31106
rect 38494 31054 38546 31106
rect 38546 31054 38548 31106
rect 38492 31052 38548 31054
rect 38652 31106 38708 31108
rect 38652 31054 38654 31106
rect 38654 31054 38706 31106
rect 38706 31054 38708 31106
rect 38652 31052 38708 31054
rect 38812 31106 38868 31108
rect 38812 31054 38814 31106
rect 38814 31054 38866 31106
rect 38866 31054 38868 31106
rect 38812 31052 38868 31054
rect 38972 31106 39028 31108
rect 38972 31054 38974 31106
rect 38974 31054 39026 31106
rect 39026 31054 39028 31106
rect 38972 31052 39028 31054
rect 39132 31106 39188 31108
rect 39132 31054 39134 31106
rect 39134 31054 39186 31106
rect 39186 31054 39188 31106
rect 39132 31052 39188 31054
rect 39292 31106 39348 31108
rect 39292 31054 39294 31106
rect 39294 31054 39346 31106
rect 39346 31054 39348 31106
rect 39292 31052 39348 31054
rect 39452 31106 39508 31108
rect 39452 31054 39454 31106
rect 39454 31054 39506 31106
rect 39506 31054 39508 31106
rect 39452 31052 39508 31054
rect 39612 31106 39668 31108
rect 39612 31054 39614 31106
rect 39614 31054 39666 31106
rect 39666 31054 39668 31106
rect 39612 31052 39668 31054
rect 39772 31106 39828 31108
rect 39772 31054 39774 31106
rect 39774 31054 39826 31106
rect 39826 31054 39828 31106
rect 39772 31052 39828 31054
rect 39932 31106 39988 31108
rect 39932 31054 39934 31106
rect 39934 31054 39986 31106
rect 39986 31054 39988 31106
rect 39932 31052 39988 31054
rect 40092 31106 40148 31108
rect 40092 31054 40094 31106
rect 40094 31054 40146 31106
rect 40146 31054 40148 31106
rect 40092 31052 40148 31054
rect 40252 31106 40308 31108
rect 40252 31054 40254 31106
rect 40254 31054 40306 31106
rect 40306 31054 40308 31106
rect 40252 31052 40308 31054
rect 40412 31106 40468 31108
rect 40412 31054 40414 31106
rect 40414 31054 40466 31106
rect 40466 31054 40468 31106
rect 40412 31052 40468 31054
rect 40572 31106 40628 31108
rect 40572 31054 40574 31106
rect 40574 31054 40626 31106
rect 40626 31054 40628 31106
rect 40572 31052 40628 31054
rect 40732 31106 40788 31108
rect 40732 31054 40734 31106
rect 40734 31054 40786 31106
rect 40786 31054 40788 31106
rect 40732 31052 40788 31054
rect 40892 31106 40948 31108
rect 40892 31054 40894 31106
rect 40894 31054 40946 31106
rect 40946 31054 40948 31106
rect 40892 31052 40948 31054
rect 41052 31106 41108 31108
rect 41052 31054 41054 31106
rect 41054 31054 41106 31106
rect 41106 31054 41108 31106
rect 41052 31052 41108 31054
rect 41212 31106 41268 31108
rect 41212 31054 41214 31106
rect 41214 31054 41266 31106
rect 41266 31054 41268 31106
rect 41212 31052 41268 31054
rect 41372 31106 41428 31108
rect 41372 31054 41374 31106
rect 41374 31054 41426 31106
rect 41426 31054 41428 31106
rect 41372 31052 41428 31054
rect 41532 31106 41588 31108
rect 41532 31054 41534 31106
rect 41534 31054 41586 31106
rect 41586 31054 41588 31106
rect 41532 31052 41588 31054
rect 41692 31106 41748 31108
rect 41692 31054 41694 31106
rect 41694 31054 41746 31106
rect 41746 31054 41748 31106
rect 41692 31052 41748 31054
rect 41852 31106 41908 31108
rect 41852 31054 41854 31106
rect 41854 31054 41906 31106
rect 41906 31054 41908 31106
rect 41852 31052 41908 31054
rect 10892 30892 10948 30948
rect 21452 30892 21508 30948
rect 30972 30892 31028 30948
rect 12 30786 68 30788
rect 12 30734 14 30786
rect 14 30734 66 30786
rect 66 30734 68 30786
rect 12 30732 68 30734
rect 172 30786 228 30788
rect 172 30734 174 30786
rect 174 30734 226 30786
rect 226 30734 228 30786
rect 172 30732 228 30734
rect 332 30786 388 30788
rect 332 30734 334 30786
rect 334 30734 386 30786
rect 386 30734 388 30786
rect 332 30732 388 30734
rect 492 30786 548 30788
rect 492 30734 494 30786
rect 494 30734 546 30786
rect 546 30734 548 30786
rect 492 30732 548 30734
rect 652 30786 708 30788
rect 652 30734 654 30786
rect 654 30734 706 30786
rect 706 30734 708 30786
rect 652 30732 708 30734
rect 812 30786 868 30788
rect 812 30734 814 30786
rect 814 30734 866 30786
rect 866 30734 868 30786
rect 812 30732 868 30734
rect 972 30786 1028 30788
rect 972 30734 974 30786
rect 974 30734 1026 30786
rect 1026 30734 1028 30786
rect 972 30732 1028 30734
rect 1132 30786 1188 30788
rect 1132 30734 1134 30786
rect 1134 30734 1186 30786
rect 1186 30734 1188 30786
rect 1132 30732 1188 30734
rect 1292 30786 1348 30788
rect 1292 30734 1294 30786
rect 1294 30734 1346 30786
rect 1346 30734 1348 30786
rect 1292 30732 1348 30734
rect 1452 30786 1508 30788
rect 1452 30734 1454 30786
rect 1454 30734 1506 30786
rect 1506 30734 1508 30786
rect 1452 30732 1508 30734
rect 1612 30786 1668 30788
rect 1612 30734 1614 30786
rect 1614 30734 1666 30786
rect 1666 30734 1668 30786
rect 1612 30732 1668 30734
rect 1772 30786 1828 30788
rect 1772 30734 1774 30786
rect 1774 30734 1826 30786
rect 1826 30734 1828 30786
rect 1772 30732 1828 30734
rect 1932 30786 1988 30788
rect 1932 30734 1934 30786
rect 1934 30734 1986 30786
rect 1986 30734 1988 30786
rect 1932 30732 1988 30734
rect 2092 30786 2148 30788
rect 2092 30734 2094 30786
rect 2094 30734 2146 30786
rect 2146 30734 2148 30786
rect 2092 30732 2148 30734
rect 2252 30786 2308 30788
rect 2252 30734 2254 30786
rect 2254 30734 2306 30786
rect 2306 30734 2308 30786
rect 2252 30732 2308 30734
rect 2412 30786 2468 30788
rect 2412 30734 2414 30786
rect 2414 30734 2466 30786
rect 2466 30734 2468 30786
rect 2412 30732 2468 30734
rect 2572 30786 2628 30788
rect 2572 30734 2574 30786
rect 2574 30734 2626 30786
rect 2626 30734 2628 30786
rect 2572 30732 2628 30734
rect 2732 30786 2788 30788
rect 2732 30734 2734 30786
rect 2734 30734 2786 30786
rect 2786 30734 2788 30786
rect 2732 30732 2788 30734
rect 2892 30786 2948 30788
rect 2892 30734 2894 30786
rect 2894 30734 2946 30786
rect 2946 30734 2948 30786
rect 2892 30732 2948 30734
rect 3052 30786 3108 30788
rect 3052 30734 3054 30786
rect 3054 30734 3106 30786
rect 3106 30734 3108 30786
rect 3052 30732 3108 30734
rect 3212 30786 3268 30788
rect 3212 30734 3214 30786
rect 3214 30734 3266 30786
rect 3266 30734 3268 30786
rect 3212 30732 3268 30734
rect 3372 30786 3428 30788
rect 3372 30734 3374 30786
rect 3374 30734 3426 30786
rect 3426 30734 3428 30786
rect 3372 30732 3428 30734
rect 3532 30786 3588 30788
rect 3532 30734 3534 30786
rect 3534 30734 3586 30786
rect 3586 30734 3588 30786
rect 3532 30732 3588 30734
rect 3692 30786 3748 30788
rect 3692 30734 3694 30786
rect 3694 30734 3746 30786
rect 3746 30734 3748 30786
rect 3692 30732 3748 30734
rect 3852 30786 3908 30788
rect 3852 30734 3854 30786
rect 3854 30734 3906 30786
rect 3906 30734 3908 30786
rect 3852 30732 3908 30734
rect 4012 30786 4068 30788
rect 4012 30734 4014 30786
rect 4014 30734 4066 30786
rect 4066 30734 4068 30786
rect 4012 30732 4068 30734
rect 4172 30786 4228 30788
rect 4172 30734 4174 30786
rect 4174 30734 4226 30786
rect 4226 30734 4228 30786
rect 4172 30732 4228 30734
rect 4332 30786 4388 30788
rect 4332 30734 4334 30786
rect 4334 30734 4386 30786
rect 4386 30734 4388 30786
rect 4332 30732 4388 30734
rect 4492 30786 4548 30788
rect 4492 30734 4494 30786
rect 4494 30734 4546 30786
rect 4546 30734 4548 30786
rect 4492 30732 4548 30734
rect 4652 30786 4708 30788
rect 4652 30734 4654 30786
rect 4654 30734 4706 30786
rect 4706 30734 4708 30786
rect 4652 30732 4708 30734
rect 4812 30786 4868 30788
rect 4812 30734 4814 30786
rect 4814 30734 4866 30786
rect 4866 30734 4868 30786
rect 4812 30732 4868 30734
rect 4972 30786 5028 30788
rect 4972 30734 4974 30786
rect 4974 30734 5026 30786
rect 5026 30734 5028 30786
rect 4972 30732 5028 30734
rect 5132 30786 5188 30788
rect 5132 30734 5134 30786
rect 5134 30734 5186 30786
rect 5186 30734 5188 30786
rect 5132 30732 5188 30734
rect 5292 30786 5348 30788
rect 5292 30734 5294 30786
rect 5294 30734 5346 30786
rect 5346 30734 5348 30786
rect 5292 30732 5348 30734
rect 5452 30786 5508 30788
rect 5452 30734 5454 30786
rect 5454 30734 5506 30786
rect 5506 30734 5508 30786
rect 5452 30732 5508 30734
rect 5612 30786 5668 30788
rect 5612 30734 5614 30786
rect 5614 30734 5666 30786
rect 5666 30734 5668 30786
rect 5612 30732 5668 30734
rect 5772 30786 5828 30788
rect 5772 30734 5774 30786
rect 5774 30734 5826 30786
rect 5826 30734 5828 30786
rect 5772 30732 5828 30734
rect 5932 30786 5988 30788
rect 5932 30734 5934 30786
rect 5934 30734 5986 30786
rect 5986 30734 5988 30786
rect 5932 30732 5988 30734
rect 6092 30786 6148 30788
rect 6092 30734 6094 30786
rect 6094 30734 6146 30786
rect 6146 30734 6148 30786
rect 6092 30732 6148 30734
rect 6252 30786 6308 30788
rect 6252 30734 6254 30786
rect 6254 30734 6306 30786
rect 6306 30734 6308 30786
rect 6252 30732 6308 30734
rect 6412 30786 6468 30788
rect 6412 30734 6414 30786
rect 6414 30734 6466 30786
rect 6466 30734 6468 30786
rect 6412 30732 6468 30734
rect 6572 30786 6628 30788
rect 6572 30734 6574 30786
rect 6574 30734 6626 30786
rect 6626 30734 6628 30786
rect 6572 30732 6628 30734
rect 6732 30786 6788 30788
rect 6732 30734 6734 30786
rect 6734 30734 6786 30786
rect 6786 30734 6788 30786
rect 6732 30732 6788 30734
rect 6892 30786 6948 30788
rect 6892 30734 6894 30786
rect 6894 30734 6946 30786
rect 6946 30734 6948 30786
rect 6892 30732 6948 30734
rect 7052 30786 7108 30788
rect 7052 30734 7054 30786
rect 7054 30734 7106 30786
rect 7106 30734 7108 30786
rect 7052 30732 7108 30734
rect 7212 30786 7268 30788
rect 7212 30734 7214 30786
rect 7214 30734 7266 30786
rect 7266 30734 7268 30786
rect 7212 30732 7268 30734
rect 7372 30786 7428 30788
rect 7372 30734 7374 30786
rect 7374 30734 7426 30786
rect 7426 30734 7428 30786
rect 7372 30732 7428 30734
rect 7532 30786 7588 30788
rect 7532 30734 7534 30786
rect 7534 30734 7586 30786
rect 7586 30734 7588 30786
rect 7532 30732 7588 30734
rect 7692 30786 7748 30788
rect 7692 30734 7694 30786
rect 7694 30734 7746 30786
rect 7746 30734 7748 30786
rect 7692 30732 7748 30734
rect 7852 30786 7908 30788
rect 7852 30734 7854 30786
rect 7854 30734 7906 30786
rect 7906 30734 7908 30786
rect 7852 30732 7908 30734
rect 8012 30786 8068 30788
rect 8012 30734 8014 30786
rect 8014 30734 8066 30786
rect 8066 30734 8068 30786
rect 8012 30732 8068 30734
rect 8172 30786 8228 30788
rect 8172 30734 8174 30786
rect 8174 30734 8226 30786
rect 8226 30734 8228 30786
rect 8172 30732 8228 30734
rect 8332 30786 8388 30788
rect 8332 30734 8334 30786
rect 8334 30734 8386 30786
rect 8386 30734 8388 30786
rect 8332 30732 8388 30734
rect 9452 30732 9508 30788
rect 9772 30732 9828 30788
rect 10092 30732 10148 30788
rect 10412 30732 10468 30788
rect 10732 30732 10788 30788
rect 11052 30732 11108 30788
rect 11372 30732 11428 30788
rect 12492 30786 12548 30788
rect 12492 30734 12494 30786
rect 12494 30734 12546 30786
rect 12546 30734 12548 30786
rect 12492 30732 12548 30734
rect 12652 30786 12708 30788
rect 12652 30734 12654 30786
rect 12654 30734 12706 30786
rect 12706 30734 12708 30786
rect 12652 30732 12708 30734
rect 12812 30786 12868 30788
rect 12812 30734 12814 30786
rect 12814 30734 12866 30786
rect 12866 30734 12868 30786
rect 12812 30732 12868 30734
rect 12972 30786 13028 30788
rect 12972 30734 12974 30786
rect 12974 30734 13026 30786
rect 13026 30734 13028 30786
rect 12972 30732 13028 30734
rect 13132 30786 13188 30788
rect 13132 30734 13134 30786
rect 13134 30734 13186 30786
rect 13186 30734 13188 30786
rect 13132 30732 13188 30734
rect 13292 30786 13348 30788
rect 13292 30734 13294 30786
rect 13294 30734 13346 30786
rect 13346 30734 13348 30786
rect 13292 30732 13348 30734
rect 13452 30786 13508 30788
rect 13452 30734 13454 30786
rect 13454 30734 13506 30786
rect 13506 30734 13508 30786
rect 13452 30732 13508 30734
rect 13612 30786 13668 30788
rect 13612 30734 13614 30786
rect 13614 30734 13666 30786
rect 13666 30734 13668 30786
rect 13612 30732 13668 30734
rect 13772 30786 13828 30788
rect 13772 30734 13774 30786
rect 13774 30734 13826 30786
rect 13826 30734 13828 30786
rect 13772 30732 13828 30734
rect 13932 30786 13988 30788
rect 13932 30734 13934 30786
rect 13934 30734 13986 30786
rect 13986 30734 13988 30786
rect 13932 30732 13988 30734
rect 14092 30786 14148 30788
rect 14092 30734 14094 30786
rect 14094 30734 14146 30786
rect 14146 30734 14148 30786
rect 14092 30732 14148 30734
rect 14252 30786 14308 30788
rect 14252 30734 14254 30786
rect 14254 30734 14306 30786
rect 14306 30734 14308 30786
rect 14252 30732 14308 30734
rect 14412 30786 14468 30788
rect 14412 30734 14414 30786
rect 14414 30734 14466 30786
rect 14466 30734 14468 30786
rect 14412 30732 14468 30734
rect 14572 30786 14628 30788
rect 14572 30734 14574 30786
rect 14574 30734 14626 30786
rect 14626 30734 14628 30786
rect 14572 30732 14628 30734
rect 14732 30786 14788 30788
rect 14732 30734 14734 30786
rect 14734 30734 14786 30786
rect 14786 30734 14788 30786
rect 14732 30732 14788 30734
rect 14892 30786 14948 30788
rect 14892 30734 14894 30786
rect 14894 30734 14946 30786
rect 14946 30734 14948 30786
rect 14892 30732 14948 30734
rect 15052 30786 15108 30788
rect 15052 30734 15054 30786
rect 15054 30734 15106 30786
rect 15106 30734 15108 30786
rect 15052 30732 15108 30734
rect 15212 30786 15268 30788
rect 15212 30734 15214 30786
rect 15214 30734 15266 30786
rect 15266 30734 15268 30786
rect 15212 30732 15268 30734
rect 15372 30786 15428 30788
rect 15372 30734 15374 30786
rect 15374 30734 15426 30786
rect 15426 30734 15428 30786
rect 15372 30732 15428 30734
rect 15532 30786 15588 30788
rect 15532 30734 15534 30786
rect 15534 30734 15586 30786
rect 15586 30734 15588 30786
rect 15532 30732 15588 30734
rect 15692 30786 15748 30788
rect 15692 30734 15694 30786
rect 15694 30734 15746 30786
rect 15746 30734 15748 30786
rect 15692 30732 15748 30734
rect 15852 30786 15908 30788
rect 15852 30734 15854 30786
rect 15854 30734 15906 30786
rect 15906 30734 15908 30786
rect 15852 30732 15908 30734
rect 16012 30786 16068 30788
rect 16012 30734 16014 30786
rect 16014 30734 16066 30786
rect 16066 30734 16068 30786
rect 16012 30732 16068 30734
rect 16172 30786 16228 30788
rect 16172 30734 16174 30786
rect 16174 30734 16226 30786
rect 16226 30734 16228 30786
rect 16172 30732 16228 30734
rect 16332 30786 16388 30788
rect 16332 30734 16334 30786
rect 16334 30734 16386 30786
rect 16386 30734 16388 30786
rect 16332 30732 16388 30734
rect 16492 30786 16548 30788
rect 16492 30734 16494 30786
rect 16494 30734 16546 30786
rect 16546 30734 16548 30786
rect 16492 30732 16548 30734
rect 16652 30786 16708 30788
rect 16652 30734 16654 30786
rect 16654 30734 16706 30786
rect 16706 30734 16708 30786
rect 16652 30732 16708 30734
rect 16812 30786 16868 30788
rect 16812 30734 16814 30786
rect 16814 30734 16866 30786
rect 16866 30734 16868 30786
rect 16812 30732 16868 30734
rect 16972 30786 17028 30788
rect 16972 30734 16974 30786
rect 16974 30734 17026 30786
rect 17026 30734 17028 30786
rect 16972 30732 17028 30734
rect 17132 30786 17188 30788
rect 17132 30734 17134 30786
rect 17134 30734 17186 30786
rect 17186 30734 17188 30786
rect 17132 30732 17188 30734
rect 17292 30786 17348 30788
rect 17292 30734 17294 30786
rect 17294 30734 17346 30786
rect 17346 30734 17348 30786
rect 17292 30732 17348 30734
rect 17452 30786 17508 30788
rect 17452 30734 17454 30786
rect 17454 30734 17506 30786
rect 17506 30734 17508 30786
rect 17452 30732 17508 30734
rect 17612 30786 17668 30788
rect 17612 30734 17614 30786
rect 17614 30734 17666 30786
rect 17666 30734 17668 30786
rect 17612 30732 17668 30734
rect 17772 30786 17828 30788
rect 17772 30734 17774 30786
rect 17774 30734 17826 30786
rect 17826 30734 17828 30786
rect 17772 30732 17828 30734
rect 17932 30786 17988 30788
rect 17932 30734 17934 30786
rect 17934 30734 17986 30786
rect 17986 30734 17988 30786
rect 17932 30732 17988 30734
rect 18092 30786 18148 30788
rect 18092 30734 18094 30786
rect 18094 30734 18146 30786
rect 18146 30734 18148 30786
rect 18092 30732 18148 30734
rect 18252 30786 18308 30788
rect 18252 30734 18254 30786
rect 18254 30734 18306 30786
rect 18306 30734 18308 30786
rect 18252 30732 18308 30734
rect 18412 30786 18468 30788
rect 18412 30734 18414 30786
rect 18414 30734 18466 30786
rect 18466 30734 18468 30786
rect 18412 30732 18468 30734
rect 18572 30786 18628 30788
rect 18572 30734 18574 30786
rect 18574 30734 18626 30786
rect 18626 30734 18628 30786
rect 18572 30732 18628 30734
rect 18732 30786 18788 30788
rect 18732 30734 18734 30786
rect 18734 30734 18786 30786
rect 18786 30734 18788 30786
rect 18732 30732 18788 30734
rect 18892 30786 18948 30788
rect 18892 30734 18894 30786
rect 18894 30734 18946 30786
rect 18946 30734 18948 30786
rect 18892 30732 18948 30734
rect 20012 30732 20068 30788
rect 20332 30732 20388 30788
rect 20652 30732 20708 30788
rect 20972 30732 21028 30788
rect 21292 30732 21348 30788
rect 21612 30732 21668 30788
rect 21932 30732 21988 30788
rect 23132 30786 23188 30788
rect 23132 30734 23134 30786
rect 23134 30734 23186 30786
rect 23186 30734 23188 30786
rect 23132 30732 23188 30734
rect 23292 30786 23348 30788
rect 23292 30734 23294 30786
rect 23294 30734 23346 30786
rect 23346 30734 23348 30786
rect 23292 30732 23348 30734
rect 23452 30786 23508 30788
rect 23452 30734 23454 30786
rect 23454 30734 23506 30786
rect 23506 30734 23508 30786
rect 23452 30732 23508 30734
rect 23612 30786 23668 30788
rect 23612 30734 23614 30786
rect 23614 30734 23666 30786
rect 23666 30734 23668 30786
rect 23612 30732 23668 30734
rect 23772 30786 23828 30788
rect 23772 30734 23774 30786
rect 23774 30734 23826 30786
rect 23826 30734 23828 30786
rect 23772 30732 23828 30734
rect 23932 30786 23988 30788
rect 23932 30734 23934 30786
rect 23934 30734 23986 30786
rect 23986 30734 23988 30786
rect 23932 30732 23988 30734
rect 24092 30786 24148 30788
rect 24092 30734 24094 30786
rect 24094 30734 24146 30786
rect 24146 30734 24148 30786
rect 24092 30732 24148 30734
rect 24252 30786 24308 30788
rect 24252 30734 24254 30786
rect 24254 30734 24306 30786
rect 24306 30734 24308 30786
rect 24252 30732 24308 30734
rect 24412 30786 24468 30788
rect 24412 30734 24414 30786
rect 24414 30734 24466 30786
rect 24466 30734 24468 30786
rect 24412 30732 24468 30734
rect 24572 30786 24628 30788
rect 24572 30734 24574 30786
rect 24574 30734 24626 30786
rect 24626 30734 24628 30786
rect 24572 30732 24628 30734
rect 24732 30786 24788 30788
rect 24732 30734 24734 30786
rect 24734 30734 24786 30786
rect 24786 30734 24788 30786
rect 24732 30732 24788 30734
rect 24892 30786 24948 30788
rect 24892 30734 24894 30786
rect 24894 30734 24946 30786
rect 24946 30734 24948 30786
rect 24892 30732 24948 30734
rect 25052 30786 25108 30788
rect 25052 30734 25054 30786
rect 25054 30734 25106 30786
rect 25106 30734 25108 30786
rect 25052 30732 25108 30734
rect 25212 30786 25268 30788
rect 25212 30734 25214 30786
rect 25214 30734 25266 30786
rect 25266 30734 25268 30786
rect 25212 30732 25268 30734
rect 25372 30786 25428 30788
rect 25372 30734 25374 30786
rect 25374 30734 25426 30786
rect 25426 30734 25428 30786
rect 25372 30732 25428 30734
rect 25532 30786 25588 30788
rect 25532 30734 25534 30786
rect 25534 30734 25586 30786
rect 25586 30734 25588 30786
rect 25532 30732 25588 30734
rect 25692 30786 25748 30788
rect 25692 30734 25694 30786
rect 25694 30734 25746 30786
rect 25746 30734 25748 30786
rect 25692 30732 25748 30734
rect 25852 30786 25908 30788
rect 25852 30734 25854 30786
rect 25854 30734 25906 30786
rect 25906 30734 25908 30786
rect 25852 30732 25908 30734
rect 26012 30786 26068 30788
rect 26012 30734 26014 30786
rect 26014 30734 26066 30786
rect 26066 30734 26068 30786
rect 26012 30732 26068 30734
rect 26172 30786 26228 30788
rect 26172 30734 26174 30786
rect 26174 30734 26226 30786
rect 26226 30734 26228 30786
rect 26172 30732 26228 30734
rect 26332 30786 26388 30788
rect 26332 30734 26334 30786
rect 26334 30734 26386 30786
rect 26386 30734 26388 30786
rect 26332 30732 26388 30734
rect 26492 30786 26548 30788
rect 26492 30734 26494 30786
rect 26494 30734 26546 30786
rect 26546 30734 26548 30786
rect 26492 30732 26548 30734
rect 26652 30786 26708 30788
rect 26652 30734 26654 30786
rect 26654 30734 26706 30786
rect 26706 30734 26708 30786
rect 26652 30732 26708 30734
rect 26812 30786 26868 30788
rect 26812 30734 26814 30786
rect 26814 30734 26866 30786
rect 26866 30734 26868 30786
rect 26812 30732 26868 30734
rect 26972 30786 27028 30788
rect 26972 30734 26974 30786
rect 26974 30734 27026 30786
rect 27026 30734 27028 30786
rect 26972 30732 27028 30734
rect 27132 30786 27188 30788
rect 27132 30734 27134 30786
rect 27134 30734 27186 30786
rect 27186 30734 27188 30786
rect 27132 30732 27188 30734
rect 27292 30786 27348 30788
rect 27292 30734 27294 30786
rect 27294 30734 27346 30786
rect 27346 30734 27348 30786
rect 27292 30732 27348 30734
rect 27452 30786 27508 30788
rect 27452 30734 27454 30786
rect 27454 30734 27506 30786
rect 27506 30734 27508 30786
rect 27452 30732 27508 30734
rect 27612 30786 27668 30788
rect 27612 30734 27614 30786
rect 27614 30734 27666 30786
rect 27666 30734 27668 30786
rect 27612 30732 27668 30734
rect 27772 30786 27828 30788
rect 27772 30734 27774 30786
rect 27774 30734 27826 30786
rect 27826 30734 27828 30786
rect 27772 30732 27828 30734
rect 27932 30786 27988 30788
rect 27932 30734 27934 30786
rect 27934 30734 27986 30786
rect 27986 30734 27988 30786
rect 27932 30732 27988 30734
rect 28092 30786 28148 30788
rect 28092 30734 28094 30786
rect 28094 30734 28146 30786
rect 28146 30734 28148 30786
rect 28092 30732 28148 30734
rect 28252 30786 28308 30788
rect 28252 30734 28254 30786
rect 28254 30734 28306 30786
rect 28306 30734 28308 30786
rect 28252 30732 28308 30734
rect 28412 30786 28468 30788
rect 28412 30734 28414 30786
rect 28414 30734 28466 30786
rect 28466 30734 28468 30786
rect 28412 30732 28468 30734
rect 28572 30786 28628 30788
rect 28572 30734 28574 30786
rect 28574 30734 28626 30786
rect 28626 30734 28628 30786
rect 28572 30732 28628 30734
rect 28732 30786 28788 30788
rect 28732 30734 28734 30786
rect 28734 30734 28786 30786
rect 28786 30734 28788 30786
rect 28732 30732 28788 30734
rect 28892 30786 28948 30788
rect 28892 30734 28894 30786
rect 28894 30734 28946 30786
rect 28946 30734 28948 30786
rect 28892 30732 28948 30734
rect 29052 30786 29108 30788
rect 29052 30734 29054 30786
rect 29054 30734 29106 30786
rect 29106 30734 29108 30786
rect 29052 30732 29108 30734
rect 29212 30786 29268 30788
rect 29212 30734 29214 30786
rect 29214 30734 29266 30786
rect 29266 30734 29268 30786
rect 29212 30732 29268 30734
rect 29372 30786 29428 30788
rect 29372 30734 29374 30786
rect 29374 30734 29426 30786
rect 29426 30734 29428 30786
rect 29372 30732 29428 30734
rect 30492 30732 30548 30788
rect 30812 30732 30868 30788
rect 31132 30732 31188 30788
rect 31452 30732 31508 30788
rect 31772 30732 31828 30788
rect 32092 30732 32148 30788
rect 32412 30732 32468 30788
rect 33532 30786 33588 30788
rect 33532 30734 33534 30786
rect 33534 30734 33586 30786
rect 33586 30734 33588 30786
rect 33532 30732 33588 30734
rect 33692 30786 33748 30788
rect 33692 30734 33694 30786
rect 33694 30734 33746 30786
rect 33746 30734 33748 30786
rect 33692 30732 33748 30734
rect 33852 30786 33908 30788
rect 33852 30734 33854 30786
rect 33854 30734 33906 30786
rect 33906 30734 33908 30786
rect 33852 30732 33908 30734
rect 34012 30786 34068 30788
rect 34012 30734 34014 30786
rect 34014 30734 34066 30786
rect 34066 30734 34068 30786
rect 34012 30732 34068 30734
rect 34172 30786 34228 30788
rect 34172 30734 34174 30786
rect 34174 30734 34226 30786
rect 34226 30734 34228 30786
rect 34172 30732 34228 30734
rect 34332 30786 34388 30788
rect 34332 30734 34334 30786
rect 34334 30734 34386 30786
rect 34386 30734 34388 30786
rect 34332 30732 34388 30734
rect 34492 30786 34548 30788
rect 34492 30734 34494 30786
rect 34494 30734 34546 30786
rect 34546 30734 34548 30786
rect 34492 30732 34548 30734
rect 34652 30786 34708 30788
rect 34652 30734 34654 30786
rect 34654 30734 34706 30786
rect 34706 30734 34708 30786
rect 34652 30732 34708 30734
rect 34812 30786 34868 30788
rect 34812 30734 34814 30786
rect 34814 30734 34866 30786
rect 34866 30734 34868 30786
rect 34812 30732 34868 30734
rect 34972 30786 35028 30788
rect 34972 30734 34974 30786
rect 34974 30734 35026 30786
rect 35026 30734 35028 30786
rect 34972 30732 35028 30734
rect 35132 30786 35188 30788
rect 35132 30734 35134 30786
rect 35134 30734 35186 30786
rect 35186 30734 35188 30786
rect 35132 30732 35188 30734
rect 35292 30786 35348 30788
rect 35292 30734 35294 30786
rect 35294 30734 35346 30786
rect 35346 30734 35348 30786
rect 35292 30732 35348 30734
rect 35452 30786 35508 30788
rect 35452 30734 35454 30786
rect 35454 30734 35506 30786
rect 35506 30734 35508 30786
rect 35452 30732 35508 30734
rect 35612 30786 35668 30788
rect 35612 30734 35614 30786
rect 35614 30734 35666 30786
rect 35666 30734 35668 30786
rect 35612 30732 35668 30734
rect 35772 30786 35828 30788
rect 35772 30734 35774 30786
rect 35774 30734 35826 30786
rect 35826 30734 35828 30786
rect 35772 30732 35828 30734
rect 35932 30786 35988 30788
rect 35932 30734 35934 30786
rect 35934 30734 35986 30786
rect 35986 30734 35988 30786
rect 35932 30732 35988 30734
rect 36092 30786 36148 30788
rect 36092 30734 36094 30786
rect 36094 30734 36146 30786
rect 36146 30734 36148 30786
rect 36092 30732 36148 30734
rect 36252 30786 36308 30788
rect 36252 30734 36254 30786
rect 36254 30734 36306 30786
rect 36306 30734 36308 30786
rect 36252 30732 36308 30734
rect 36412 30786 36468 30788
rect 36412 30734 36414 30786
rect 36414 30734 36466 30786
rect 36466 30734 36468 30786
rect 36412 30732 36468 30734
rect 36572 30786 36628 30788
rect 36572 30734 36574 30786
rect 36574 30734 36626 30786
rect 36626 30734 36628 30786
rect 36572 30732 36628 30734
rect 36732 30786 36788 30788
rect 36732 30734 36734 30786
rect 36734 30734 36786 30786
rect 36786 30734 36788 30786
rect 36732 30732 36788 30734
rect 36892 30786 36948 30788
rect 36892 30734 36894 30786
rect 36894 30734 36946 30786
rect 36946 30734 36948 30786
rect 36892 30732 36948 30734
rect 37052 30786 37108 30788
rect 37052 30734 37054 30786
rect 37054 30734 37106 30786
rect 37106 30734 37108 30786
rect 37052 30732 37108 30734
rect 37212 30786 37268 30788
rect 37212 30734 37214 30786
rect 37214 30734 37266 30786
rect 37266 30734 37268 30786
rect 37212 30732 37268 30734
rect 37372 30786 37428 30788
rect 37372 30734 37374 30786
rect 37374 30734 37426 30786
rect 37426 30734 37428 30786
rect 37372 30732 37428 30734
rect 37532 30786 37588 30788
rect 37532 30734 37534 30786
rect 37534 30734 37586 30786
rect 37586 30734 37588 30786
rect 37532 30732 37588 30734
rect 37692 30786 37748 30788
rect 37692 30734 37694 30786
rect 37694 30734 37746 30786
rect 37746 30734 37748 30786
rect 37692 30732 37748 30734
rect 37852 30786 37908 30788
rect 37852 30734 37854 30786
rect 37854 30734 37906 30786
rect 37906 30734 37908 30786
rect 37852 30732 37908 30734
rect 38012 30786 38068 30788
rect 38012 30734 38014 30786
rect 38014 30734 38066 30786
rect 38066 30734 38068 30786
rect 38012 30732 38068 30734
rect 38172 30786 38228 30788
rect 38172 30734 38174 30786
rect 38174 30734 38226 30786
rect 38226 30734 38228 30786
rect 38172 30732 38228 30734
rect 38332 30786 38388 30788
rect 38332 30734 38334 30786
rect 38334 30734 38386 30786
rect 38386 30734 38388 30786
rect 38332 30732 38388 30734
rect 38492 30786 38548 30788
rect 38492 30734 38494 30786
rect 38494 30734 38546 30786
rect 38546 30734 38548 30786
rect 38492 30732 38548 30734
rect 38652 30786 38708 30788
rect 38652 30734 38654 30786
rect 38654 30734 38706 30786
rect 38706 30734 38708 30786
rect 38652 30732 38708 30734
rect 38812 30786 38868 30788
rect 38812 30734 38814 30786
rect 38814 30734 38866 30786
rect 38866 30734 38868 30786
rect 38812 30732 38868 30734
rect 38972 30786 39028 30788
rect 38972 30734 38974 30786
rect 38974 30734 39026 30786
rect 39026 30734 39028 30786
rect 38972 30732 39028 30734
rect 39132 30786 39188 30788
rect 39132 30734 39134 30786
rect 39134 30734 39186 30786
rect 39186 30734 39188 30786
rect 39132 30732 39188 30734
rect 39292 30786 39348 30788
rect 39292 30734 39294 30786
rect 39294 30734 39346 30786
rect 39346 30734 39348 30786
rect 39292 30732 39348 30734
rect 39452 30786 39508 30788
rect 39452 30734 39454 30786
rect 39454 30734 39506 30786
rect 39506 30734 39508 30786
rect 39452 30732 39508 30734
rect 39612 30786 39668 30788
rect 39612 30734 39614 30786
rect 39614 30734 39666 30786
rect 39666 30734 39668 30786
rect 39612 30732 39668 30734
rect 39772 30786 39828 30788
rect 39772 30734 39774 30786
rect 39774 30734 39826 30786
rect 39826 30734 39828 30786
rect 39772 30732 39828 30734
rect 39932 30786 39988 30788
rect 39932 30734 39934 30786
rect 39934 30734 39986 30786
rect 39986 30734 39988 30786
rect 39932 30732 39988 30734
rect 40092 30786 40148 30788
rect 40092 30734 40094 30786
rect 40094 30734 40146 30786
rect 40146 30734 40148 30786
rect 40092 30732 40148 30734
rect 40252 30786 40308 30788
rect 40252 30734 40254 30786
rect 40254 30734 40306 30786
rect 40306 30734 40308 30786
rect 40252 30732 40308 30734
rect 40412 30786 40468 30788
rect 40412 30734 40414 30786
rect 40414 30734 40466 30786
rect 40466 30734 40468 30786
rect 40412 30732 40468 30734
rect 40572 30786 40628 30788
rect 40572 30734 40574 30786
rect 40574 30734 40626 30786
rect 40626 30734 40628 30786
rect 40572 30732 40628 30734
rect 40732 30786 40788 30788
rect 40732 30734 40734 30786
rect 40734 30734 40786 30786
rect 40786 30734 40788 30786
rect 40732 30732 40788 30734
rect 40892 30786 40948 30788
rect 40892 30734 40894 30786
rect 40894 30734 40946 30786
rect 40946 30734 40948 30786
rect 40892 30732 40948 30734
rect 41052 30786 41108 30788
rect 41052 30734 41054 30786
rect 41054 30734 41106 30786
rect 41106 30734 41108 30786
rect 41052 30732 41108 30734
rect 41212 30786 41268 30788
rect 41212 30734 41214 30786
rect 41214 30734 41266 30786
rect 41266 30734 41268 30786
rect 41212 30732 41268 30734
rect 41372 30786 41428 30788
rect 41372 30734 41374 30786
rect 41374 30734 41426 30786
rect 41426 30734 41428 30786
rect 41372 30732 41428 30734
rect 41532 30786 41588 30788
rect 41532 30734 41534 30786
rect 41534 30734 41586 30786
rect 41586 30734 41588 30786
rect 41532 30732 41588 30734
rect 41692 30786 41748 30788
rect 41692 30734 41694 30786
rect 41694 30734 41746 30786
rect 41746 30734 41748 30786
rect 41692 30732 41748 30734
rect 41852 30786 41908 30788
rect 41852 30734 41854 30786
rect 41854 30734 41906 30786
rect 41906 30734 41908 30786
rect 41852 30732 41908 30734
rect 11212 30572 11268 30628
rect 21772 30572 21828 30628
rect 30652 30572 30708 30628
rect 12 30466 68 30468
rect 12 30414 14 30466
rect 14 30414 66 30466
rect 66 30414 68 30466
rect 12 30412 68 30414
rect 172 30466 228 30468
rect 172 30414 174 30466
rect 174 30414 226 30466
rect 226 30414 228 30466
rect 172 30412 228 30414
rect 332 30466 388 30468
rect 332 30414 334 30466
rect 334 30414 386 30466
rect 386 30414 388 30466
rect 332 30412 388 30414
rect 492 30466 548 30468
rect 492 30414 494 30466
rect 494 30414 546 30466
rect 546 30414 548 30466
rect 492 30412 548 30414
rect 652 30466 708 30468
rect 652 30414 654 30466
rect 654 30414 706 30466
rect 706 30414 708 30466
rect 652 30412 708 30414
rect 812 30466 868 30468
rect 812 30414 814 30466
rect 814 30414 866 30466
rect 866 30414 868 30466
rect 812 30412 868 30414
rect 972 30466 1028 30468
rect 972 30414 974 30466
rect 974 30414 1026 30466
rect 1026 30414 1028 30466
rect 972 30412 1028 30414
rect 1132 30466 1188 30468
rect 1132 30414 1134 30466
rect 1134 30414 1186 30466
rect 1186 30414 1188 30466
rect 1132 30412 1188 30414
rect 1292 30466 1348 30468
rect 1292 30414 1294 30466
rect 1294 30414 1346 30466
rect 1346 30414 1348 30466
rect 1292 30412 1348 30414
rect 1452 30466 1508 30468
rect 1452 30414 1454 30466
rect 1454 30414 1506 30466
rect 1506 30414 1508 30466
rect 1452 30412 1508 30414
rect 1612 30466 1668 30468
rect 1612 30414 1614 30466
rect 1614 30414 1666 30466
rect 1666 30414 1668 30466
rect 1612 30412 1668 30414
rect 1772 30466 1828 30468
rect 1772 30414 1774 30466
rect 1774 30414 1826 30466
rect 1826 30414 1828 30466
rect 1772 30412 1828 30414
rect 1932 30466 1988 30468
rect 1932 30414 1934 30466
rect 1934 30414 1986 30466
rect 1986 30414 1988 30466
rect 1932 30412 1988 30414
rect 2092 30466 2148 30468
rect 2092 30414 2094 30466
rect 2094 30414 2146 30466
rect 2146 30414 2148 30466
rect 2092 30412 2148 30414
rect 2252 30466 2308 30468
rect 2252 30414 2254 30466
rect 2254 30414 2306 30466
rect 2306 30414 2308 30466
rect 2252 30412 2308 30414
rect 2412 30466 2468 30468
rect 2412 30414 2414 30466
rect 2414 30414 2466 30466
rect 2466 30414 2468 30466
rect 2412 30412 2468 30414
rect 2572 30466 2628 30468
rect 2572 30414 2574 30466
rect 2574 30414 2626 30466
rect 2626 30414 2628 30466
rect 2572 30412 2628 30414
rect 2732 30466 2788 30468
rect 2732 30414 2734 30466
rect 2734 30414 2786 30466
rect 2786 30414 2788 30466
rect 2732 30412 2788 30414
rect 2892 30466 2948 30468
rect 2892 30414 2894 30466
rect 2894 30414 2946 30466
rect 2946 30414 2948 30466
rect 2892 30412 2948 30414
rect 3052 30466 3108 30468
rect 3052 30414 3054 30466
rect 3054 30414 3106 30466
rect 3106 30414 3108 30466
rect 3052 30412 3108 30414
rect 3212 30466 3268 30468
rect 3212 30414 3214 30466
rect 3214 30414 3266 30466
rect 3266 30414 3268 30466
rect 3212 30412 3268 30414
rect 3372 30466 3428 30468
rect 3372 30414 3374 30466
rect 3374 30414 3426 30466
rect 3426 30414 3428 30466
rect 3372 30412 3428 30414
rect 3532 30466 3588 30468
rect 3532 30414 3534 30466
rect 3534 30414 3586 30466
rect 3586 30414 3588 30466
rect 3532 30412 3588 30414
rect 3692 30466 3748 30468
rect 3692 30414 3694 30466
rect 3694 30414 3746 30466
rect 3746 30414 3748 30466
rect 3692 30412 3748 30414
rect 3852 30466 3908 30468
rect 3852 30414 3854 30466
rect 3854 30414 3906 30466
rect 3906 30414 3908 30466
rect 3852 30412 3908 30414
rect 4012 30466 4068 30468
rect 4012 30414 4014 30466
rect 4014 30414 4066 30466
rect 4066 30414 4068 30466
rect 4012 30412 4068 30414
rect 4172 30466 4228 30468
rect 4172 30414 4174 30466
rect 4174 30414 4226 30466
rect 4226 30414 4228 30466
rect 4172 30412 4228 30414
rect 4332 30466 4388 30468
rect 4332 30414 4334 30466
rect 4334 30414 4386 30466
rect 4386 30414 4388 30466
rect 4332 30412 4388 30414
rect 4492 30466 4548 30468
rect 4492 30414 4494 30466
rect 4494 30414 4546 30466
rect 4546 30414 4548 30466
rect 4492 30412 4548 30414
rect 4652 30466 4708 30468
rect 4652 30414 4654 30466
rect 4654 30414 4706 30466
rect 4706 30414 4708 30466
rect 4652 30412 4708 30414
rect 4812 30466 4868 30468
rect 4812 30414 4814 30466
rect 4814 30414 4866 30466
rect 4866 30414 4868 30466
rect 4812 30412 4868 30414
rect 4972 30466 5028 30468
rect 4972 30414 4974 30466
rect 4974 30414 5026 30466
rect 5026 30414 5028 30466
rect 4972 30412 5028 30414
rect 5132 30466 5188 30468
rect 5132 30414 5134 30466
rect 5134 30414 5186 30466
rect 5186 30414 5188 30466
rect 5132 30412 5188 30414
rect 5292 30466 5348 30468
rect 5292 30414 5294 30466
rect 5294 30414 5346 30466
rect 5346 30414 5348 30466
rect 5292 30412 5348 30414
rect 5452 30466 5508 30468
rect 5452 30414 5454 30466
rect 5454 30414 5506 30466
rect 5506 30414 5508 30466
rect 5452 30412 5508 30414
rect 5612 30466 5668 30468
rect 5612 30414 5614 30466
rect 5614 30414 5666 30466
rect 5666 30414 5668 30466
rect 5612 30412 5668 30414
rect 5772 30466 5828 30468
rect 5772 30414 5774 30466
rect 5774 30414 5826 30466
rect 5826 30414 5828 30466
rect 5772 30412 5828 30414
rect 5932 30466 5988 30468
rect 5932 30414 5934 30466
rect 5934 30414 5986 30466
rect 5986 30414 5988 30466
rect 5932 30412 5988 30414
rect 6092 30466 6148 30468
rect 6092 30414 6094 30466
rect 6094 30414 6146 30466
rect 6146 30414 6148 30466
rect 6092 30412 6148 30414
rect 6252 30466 6308 30468
rect 6252 30414 6254 30466
rect 6254 30414 6306 30466
rect 6306 30414 6308 30466
rect 6252 30412 6308 30414
rect 6412 30466 6468 30468
rect 6412 30414 6414 30466
rect 6414 30414 6466 30466
rect 6466 30414 6468 30466
rect 6412 30412 6468 30414
rect 6572 30466 6628 30468
rect 6572 30414 6574 30466
rect 6574 30414 6626 30466
rect 6626 30414 6628 30466
rect 6572 30412 6628 30414
rect 6732 30466 6788 30468
rect 6732 30414 6734 30466
rect 6734 30414 6786 30466
rect 6786 30414 6788 30466
rect 6732 30412 6788 30414
rect 6892 30466 6948 30468
rect 6892 30414 6894 30466
rect 6894 30414 6946 30466
rect 6946 30414 6948 30466
rect 6892 30412 6948 30414
rect 7052 30466 7108 30468
rect 7052 30414 7054 30466
rect 7054 30414 7106 30466
rect 7106 30414 7108 30466
rect 7052 30412 7108 30414
rect 7212 30466 7268 30468
rect 7212 30414 7214 30466
rect 7214 30414 7266 30466
rect 7266 30414 7268 30466
rect 7212 30412 7268 30414
rect 7372 30466 7428 30468
rect 7372 30414 7374 30466
rect 7374 30414 7426 30466
rect 7426 30414 7428 30466
rect 7372 30412 7428 30414
rect 7532 30466 7588 30468
rect 7532 30414 7534 30466
rect 7534 30414 7586 30466
rect 7586 30414 7588 30466
rect 7532 30412 7588 30414
rect 7692 30466 7748 30468
rect 7692 30414 7694 30466
rect 7694 30414 7746 30466
rect 7746 30414 7748 30466
rect 7692 30412 7748 30414
rect 7852 30466 7908 30468
rect 7852 30414 7854 30466
rect 7854 30414 7906 30466
rect 7906 30414 7908 30466
rect 7852 30412 7908 30414
rect 8012 30466 8068 30468
rect 8012 30414 8014 30466
rect 8014 30414 8066 30466
rect 8066 30414 8068 30466
rect 8012 30412 8068 30414
rect 8172 30466 8228 30468
rect 8172 30414 8174 30466
rect 8174 30414 8226 30466
rect 8226 30414 8228 30466
rect 8172 30412 8228 30414
rect 8332 30466 8388 30468
rect 8332 30414 8334 30466
rect 8334 30414 8386 30466
rect 8386 30414 8388 30466
rect 8332 30412 8388 30414
rect 9452 30412 9508 30468
rect 9772 30412 9828 30468
rect 10092 30412 10148 30468
rect 10412 30412 10468 30468
rect 10732 30412 10788 30468
rect 11052 30412 11108 30468
rect 11372 30412 11428 30468
rect 12492 30466 12548 30468
rect 12492 30414 12494 30466
rect 12494 30414 12546 30466
rect 12546 30414 12548 30466
rect 12492 30412 12548 30414
rect 12652 30466 12708 30468
rect 12652 30414 12654 30466
rect 12654 30414 12706 30466
rect 12706 30414 12708 30466
rect 12652 30412 12708 30414
rect 12812 30466 12868 30468
rect 12812 30414 12814 30466
rect 12814 30414 12866 30466
rect 12866 30414 12868 30466
rect 12812 30412 12868 30414
rect 12972 30466 13028 30468
rect 12972 30414 12974 30466
rect 12974 30414 13026 30466
rect 13026 30414 13028 30466
rect 12972 30412 13028 30414
rect 13132 30466 13188 30468
rect 13132 30414 13134 30466
rect 13134 30414 13186 30466
rect 13186 30414 13188 30466
rect 13132 30412 13188 30414
rect 13292 30466 13348 30468
rect 13292 30414 13294 30466
rect 13294 30414 13346 30466
rect 13346 30414 13348 30466
rect 13292 30412 13348 30414
rect 13452 30466 13508 30468
rect 13452 30414 13454 30466
rect 13454 30414 13506 30466
rect 13506 30414 13508 30466
rect 13452 30412 13508 30414
rect 13612 30466 13668 30468
rect 13612 30414 13614 30466
rect 13614 30414 13666 30466
rect 13666 30414 13668 30466
rect 13612 30412 13668 30414
rect 13772 30466 13828 30468
rect 13772 30414 13774 30466
rect 13774 30414 13826 30466
rect 13826 30414 13828 30466
rect 13772 30412 13828 30414
rect 13932 30466 13988 30468
rect 13932 30414 13934 30466
rect 13934 30414 13986 30466
rect 13986 30414 13988 30466
rect 13932 30412 13988 30414
rect 14092 30466 14148 30468
rect 14092 30414 14094 30466
rect 14094 30414 14146 30466
rect 14146 30414 14148 30466
rect 14092 30412 14148 30414
rect 14252 30466 14308 30468
rect 14252 30414 14254 30466
rect 14254 30414 14306 30466
rect 14306 30414 14308 30466
rect 14252 30412 14308 30414
rect 14412 30466 14468 30468
rect 14412 30414 14414 30466
rect 14414 30414 14466 30466
rect 14466 30414 14468 30466
rect 14412 30412 14468 30414
rect 14572 30466 14628 30468
rect 14572 30414 14574 30466
rect 14574 30414 14626 30466
rect 14626 30414 14628 30466
rect 14572 30412 14628 30414
rect 14732 30466 14788 30468
rect 14732 30414 14734 30466
rect 14734 30414 14786 30466
rect 14786 30414 14788 30466
rect 14732 30412 14788 30414
rect 14892 30466 14948 30468
rect 14892 30414 14894 30466
rect 14894 30414 14946 30466
rect 14946 30414 14948 30466
rect 14892 30412 14948 30414
rect 15052 30466 15108 30468
rect 15052 30414 15054 30466
rect 15054 30414 15106 30466
rect 15106 30414 15108 30466
rect 15052 30412 15108 30414
rect 15212 30466 15268 30468
rect 15212 30414 15214 30466
rect 15214 30414 15266 30466
rect 15266 30414 15268 30466
rect 15212 30412 15268 30414
rect 15372 30466 15428 30468
rect 15372 30414 15374 30466
rect 15374 30414 15426 30466
rect 15426 30414 15428 30466
rect 15372 30412 15428 30414
rect 15532 30466 15588 30468
rect 15532 30414 15534 30466
rect 15534 30414 15586 30466
rect 15586 30414 15588 30466
rect 15532 30412 15588 30414
rect 15692 30466 15748 30468
rect 15692 30414 15694 30466
rect 15694 30414 15746 30466
rect 15746 30414 15748 30466
rect 15692 30412 15748 30414
rect 15852 30466 15908 30468
rect 15852 30414 15854 30466
rect 15854 30414 15906 30466
rect 15906 30414 15908 30466
rect 15852 30412 15908 30414
rect 16012 30466 16068 30468
rect 16012 30414 16014 30466
rect 16014 30414 16066 30466
rect 16066 30414 16068 30466
rect 16012 30412 16068 30414
rect 16172 30466 16228 30468
rect 16172 30414 16174 30466
rect 16174 30414 16226 30466
rect 16226 30414 16228 30466
rect 16172 30412 16228 30414
rect 16332 30466 16388 30468
rect 16332 30414 16334 30466
rect 16334 30414 16386 30466
rect 16386 30414 16388 30466
rect 16332 30412 16388 30414
rect 16492 30466 16548 30468
rect 16492 30414 16494 30466
rect 16494 30414 16546 30466
rect 16546 30414 16548 30466
rect 16492 30412 16548 30414
rect 16652 30466 16708 30468
rect 16652 30414 16654 30466
rect 16654 30414 16706 30466
rect 16706 30414 16708 30466
rect 16652 30412 16708 30414
rect 16812 30466 16868 30468
rect 16812 30414 16814 30466
rect 16814 30414 16866 30466
rect 16866 30414 16868 30466
rect 16812 30412 16868 30414
rect 16972 30466 17028 30468
rect 16972 30414 16974 30466
rect 16974 30414 17026 30466
rect 17026 30414 17028 30466
rect 16972 30412 17028 30414
rect 17132 30466 17188 30468
rect 17132 30414 17134 30466
rect 17134 30414 17186 30466
rect 17186 30414 17188 30466
rect 17132 30412 17188 30414
rect 17292 30466 17348 30468
rect 17292 30414 17294 30466
rect 17294 30414 17346 30466
rect 17346 30414 17348 30466
rect 17292 30412 17348 30414
rect 17452 30466 17508 30468
rect 17452 30414 17454 30466
rect 17454 30414 17506 30466
rect 17506 30414 17508 30466
rect 17452 30412 17508 30414
rect 17612 30466 17668 30468
rect 17612 30414 17614 30466
rect 17614 30414 17666 30466
rect 17666 30414 17668 30466
rect 17612 30412 17668 30414
rect 17772 30466 17828 30468
rect 17772 30414 17774 30466
rect 17774 30414 17826 30466
rect 17826 30414 17828 30466
rect 17772 30412 17828 30414
rect 17932 30466 17988 30468
rect 17932 30414 17934 30466
rect 17934 30414 17986 30466
rect 17986 30414 17988 30466
rect 17932 30412 17988 30414
rect 18092 30466 18148 30468
rect 18092 30414 18094 30466
rect 18094 30414 18146 30466
rect 18146 30414 18148 30466
rect 18092 30412 18148 30414
rect 18252 30466 18308 30468
rect 18252 30414 18254 30466
rect 18254 30414 18306 30466
rect 18306 30414 18308 30466
rect 18252 30412 18308 30414
rect 18412 30466 18468 30468
rect 18412 30414 18414 30466
rect 18414 30414 18466 30466
rect 18466 30414 18468 30466
rect 18412 30412 18468 30414
rect 18572 30466 18628 30468
rect 18572 30414 18574 30466
rect 18574 30414 18626 30466
rect 18626 30414 18628 30466
rect 18572 30412 18628 30414
rect 18732 30466 18788 30468
rect 18732 30414 18734 30466
rect 18734 30414 18786 30466
rect 18786 30414 18788 30466
rect 18732 30412 18788 30414
rect 18892 30466 18948 30468
rect 18892 30414 18894 30466
rect 18894 30414 18946 30466
rect 18946 30414 18948 30466
rect 18892 30412 18948 30414
rect 20012 30412 20068 30468
rect 20332 30412 20388 30468
rect 20652 30412 20708 30468
rect 20972 30412 21028 30468
rect 21292 30412 21348 30468
rect 21612 30412 21668 30468
rect 21932 30412 21988 30468
rect 23132 30466 23188 30468
rect 23132 30414 23134 30466
rect 23134 30414 23186 30466
rect 23186 30414 23188 30466
rect 23132 30412 23188 30414
rect 23292 30466 23348 30468
rect 23292 30414 23294 30466
rect 23294 30414 23346 30466
rect 23346 30414 23348 30466
rect 23292 30412 23348 30414
rect 23452 30466 23508 30468
rect 23452 30414 23454 30466
rect 23454 30414 23506 30466
rect 23506 30414 23508 30466
rect 23452 30412 23508 30414
rect 23612 30466 23668 30468
rect 23612 30414 23614 30466
rect 23614 30414 23666 30466
rect 23666 30414 23668 30466
rect 23612 30412 23668 30414
rect 23772 30466 23828 30468
rect 23772 30414 23774 30466
rect 23774 30414 23826 30466
rect 23826 30414 23828 30466
rect 23772 30412 23828 30414
rect 23932 30466 23988 30468
rect 23932 30414 23934 30466
rect 23934 30414 23986 30466
rect 23986 30414 23988 30466
rect 23932 30412 23988 30414
rect 24092 30466 24148 30468
rect 24092 30414 24094 30466
rect 24094 30414 24146 30466
rect 24146 30414 24148 30466
rect 24092 30412 24148 30414
rect 24252 30466 24308 30468
rect 24252 30414 24254 30466
rect 24254 30414 24306 30466
rect 24306 30414 24308 30466
rect 24252 30412 24308 30414
rect 24412 30466 24468 30468
rect 24412 30414 24414 30466
rect 24414 30414 24466 30466
rect 24466 30414 24468 30466
rect 24412 30412 24468 30414
rect 24572 30466 24628 30468
rect 24572 30414 24574 30466
rect 24574 30414 24626 30466
rect 24626 30414 24628 30466
rect 24572 30412 24628 30414
rect 24732 30466 24788 30468
rect 24732 30414 24734 30466
rect 24734 30414 24786 30466
rect 24786 30414 24788 30466
rect 24732 30412 24788 30414
rect 24892 30466 24948 30468
rect 24892 30414 24894 30466
rect 24894 30414 24946 30466
rect 24946 30414 24948 30466
rect 24892 30412 24948 30414
rect 25052 30466 25108 30468
rect 25052 30414 25054 30466
rect 25054 30414 25106 30466
rect 25106 30414 25108 30466
rect 25052 30412 25108 30414
rect 25212 30466 25268 30468
rect 25212 30414 25214 30466
rect 25214 30414 25266 30466
rect 25266 30414 25268 30466
rect 25212 30412 25268 30414
rect 25372 30466 25428 30468
rect 25372 30414 25374 30466
rect 25374 30414 25426 30466
rect 25426 30414 25428 30466
rect 25372 30412 25428 30414
rect 25532 30466 25588 30468
rect 25532 30414 25534 30466
rect 25534 30414 25586 30466
rect 25586 30414 25588 30466
rect 25532 30412 25588 30414
rect 25692 30466 25748 30468
rect 25692 30414 25694 30466
rect 25694 30414 25746 30466
rect 25746 30414 25748 30466
rect 25692 30412 25748 30414
rect 25852 30466 25908 30468
rect 25852 30414 25854 30466
rect 25854 30414 25906 30466
rect 25906 30414 25908 30466
rect 25852 30412 25908 30414
rect 26012 30466 26068 30468
rect 26012 30414 26014 30466
rect 26014 30414 26066 30466
rect 26066 30414 26068 30466
rect 26012 30412 26068 30414
rect 26172 30466 26228 30468
rect 26172 30414 26174 30466
rect 26174 30414 26226 30466
rect 26226 30414 26228 30466
rect 26172 30412 26228 30414
rect 26332 30466 26388 30468
rect 26332 30414 26334 30466
rect 26334 30414 26386 30466
rect 26386 30414 26388 30466
rect 26332 30412 26388 30414
rect 26492 30466 26548 30468
rect 26492 30414 26494 30466
rect 26494 30414 26546 30466
rect 26546 30414 26548 30466
rect 26492 30412 26548 30414
rect 26652 30466 26708 30468
rect 26652 30414 26654 30466
rect 26654 30414 26706 30466
rect 26706 30414 26708 30466
rect 26652 30412 26708 30414
rect 26812 30466 26868 30468
rect 26812 30414 26814 30466
rect 26814 30414 26866 30466
rect 26866 30414 26868 30466
rect 26812 30412 26868 30414
rect 26972 30466 27028 30468
rect 26972 30414 26974 30466
rect 26974 30414 27026 30466
rect 27026 30414 27028 30466
rect 26972 30412 27028 30414
rect 27132 30466 27188 30468
rect 27132 30414 27134 30466
rect 27134 30414 27186 30466
rect 27186 30414 27188 30466
rect 27132 30412 27188 30414
rect 27292 30466 27348 30468
rect 27292 30414 27294 30466
rect 27294 30414 27346 30466
rect 27346 30414 27348 30466
rect 27292 30412 27348 30414
rect 27452 30466 27508 30468
rect 27452 30414 27454 30466
rect 27454 30414 27506 30466
rect 27506 30414 27508 30466
rect 27452 30412 27508 30414
rect 27612 30466 27668 30468
rect 27612 30414 27614 30466
rect 27614 30414 27666 30466
rect 27666 30414 27668 30466
rect 27612 30412 27668 30414
rect 27772 30466 27828 30468
rect 27772 30414 27774 30466
rect 27774 30414 27826 30466
rect 27826 30414 27828 30466
rect 27772 30412 27828 30414
rect 27932 30466 27988 30468
rect 27932 30414 27934 30466
rect 27934 30414 27986 30466
rect 27986 30414 27988 30466
rect 27932 30412 27988 30414
rect 28092 30466 28148 30468
rect 28092 30414 28094 30466
rect 28094 30414 28146 30466
rect 28146 30414 28148 30466
rect 28092 30412 28148 30414
rect 28252 30466 28308 30468
rect 28252 30414 28254 30466
rect 28254 30414 28306 30466
rect 28306 30414 28308 30466
rect 28252 30412 28308 30414
rect 28412 30466 28468 30468
rect 28412 30414 28414 30466
rect 28414 30414 28466 30466
rect 28466 30414 28468 30466
rect 28412 30412 28468 30414
rect 28572 30466 28628 30468
rect 28572 30414 28574 30466
rect 28574 30414 28626 30466
rect 28626 30414 28628 30466
rect 28572 30412 28628 30414
rect 28732 30466 28788 30468
rect 28732 30414 28734 30466
rect 28734 30414 28786 30466
rect 28786 30414 28788 30466
rect 28732 30412 28788 30414
rect 28892 30466 28948 30468
rect 28892 30414 28894 30466
rect 28894 30414 28946 30466
rect 28946 30414 28948 30466
rect 28892 30412 28948 30414
rect 29052 30466 29108 30468
rect 29052 30414 29054 30466
rect 29054 30414 29106 30466
rect 29106 30414 29108 30466
rect 29052 30412 29108 30414
rect 29212 30466 29268 30468
rect 29212 30414 29214 30466
rect 29214 30414 29266 30466
rect 29266 30414 29268 30466
rect 29212 30412 29268 30414
rect 29372 30466 29428 30468
rect 29372 30414 29374 30466
rect 29374 30414 29426 30466
rect 29426 30414 29428 30466
rect 29372 30412 29428 30414
rect 30492 30412 30548 30468
rect 30812 30412 30868 30468
rect 31132 30412 31188 30468
rect 31452 30412 31508 30468
rect 31772 30412 31828 30468
rect 32092 30412 32148 30468
rect 32412 30412 32468 30468
rect 33532 30466 33588 30468
rect 33532 30414 33534 30466
rect 33534 30414 33586 30466
rect 33586 30414 33588 30466
rect 33532 30412 33588 30414
rect 33692 30466 33748 30468
rect 33692 30414 33694 30466
rect 33694 30414 33746 30466
rect 33746 30414 33748 30466
rect 33692 30412 33748 30414
rect 33852 30466 33908 30468
rect 33852 30414 33854 30466
rect 33854 30414 33906 30466
rect 33906 30414 33908 30466
rect 33852 30412 33908 30414
rect 34012 30466 34068 30468
rect 34012 30414 34014 30466
rect 34014 30414 34066 30466
rect 34066 30414 34068 30466
rect 34012 30412 34068 30414
rect 34172 30466 34228 30468
rect 34172 30414 34174 30466
rect 34174 30414 34226 30466
rect 34226 30414 34228 30466
rect 34172 30412 34228 30414
rect 34332 30466 34388 30468
rect 34332 30414 34334 30466
rect 34334 30414 34386 30466
rect 34386 30414 34388 30466
rect 34332 30412 34388 30414
rect 34492 30466 34548 30468
rect 34492 30414 34494 30466
rect 34494 30414 34546 30466
rect 34546 30414 34548 30466
rect 34492 30412 34548 30414
rect 34652 30466 34708 30468
rect 34652 30414 34654 30466
rect 34654 30414 34706 30466
rect 34706 30414 34708 30466
rect 34652 30412 34708 30414
rect 34812 30466 34868 30468
rect 34812 30414 34814 30466
rect 34814 30414 34866 30466
rect 34866 30414 34868 30466
rect 34812 30412 34868 30414
rect 34972 30466 35028 30468
rect 34972 30414 34974 30466
rect 34974 30414 35026 30466
rect 35026 30414 35028 30466
rect 34972 30412 35028 30414
rect 35132 30466 35188 30468
rect 35132 30414 35134 30466
rect 35134 30414 35186 30466
rect 35186 30414 35188 30466
rect 35132 30412 35188 30414
rect 35292 30466 35348 30468
rect 35292 30414 35294 30466
rect 35294 30414 35346 30466
rect 35346 30414 35348 30466
rect 35292 30412 35348 30414
rect 35452 30466 35508 30468
rect 35452 30414 35454 30466
rect 35454 30414 35506 30466
rect 35506 30414 35508 30466
rect 35452 30412 35508 30414
rect 35612 30466 35668 30468
rect 35612 30414 35614 30466
rect 35614 30414 35666 30466
rect 35666 30414 35668 30466
rect 35612 30412 35668 30414
rect 35772 30466 35828 30468
rect 35772 30414 35774 30466
rect 35774 30414 35826 30466
rect 35826 30414 35828 30466
rect 35772 30412 35828 30414
rect 35932 30466 35988 30468
rect 35932 30414 35934 30466
rect 35934 30414 35986 30466
rect 35986 30414 35988 30466
rect 35932 30412 35988 30414
rect 36092 30466 36148 30468
rect 36092 30414 36094 30466
rect 36094 30414 36146 30466
rect 36146 30414 36148 30466
rect 36092 30412 36148 30414
rect 36252 30466 36308 30468
rect 36252 30414 36254 30466
rect 36254 30414 36306 30466
rect 36306 30414 36308 30466
rect 36252 30412 36308 30414
rect 36412 30466 36468 30468
rect 36412 30414 36414 30466
rect 36414 30414 36466 30466
rect 36466 30414 36468 30466
rect 36412 30412 36468 30414
rect 36572 30466 36628 30468
rect 36572 30414 36574 30466
rect 36574 30414 36626 30466
rect 36626 30414 36628 30466
rect 36572 30412 36628 30414
rect 36732 30466 36788 30468
rect 36732 30414 36734 30466
rect 36734 30414 36786 30466
rect 36786 30414 36788 30466
rect 36732 30412 36788 30414
rect 36892 30466 36948 30468
rect 36892 30414 36894 30466
rect 36894 30414 36946 30466
rect 36946 30414 36948 30466
rect 36892 30412 36948 30414
rect 37052 30466 37108 30468
rect 37052 30414 37054 30466
rect 37054 30414 37106 30466
rect 37106 30414 37108 30466
rect 37052 30412 37108 30414
rect 37212 30466 37268 30468
rect 37212 30414 37214 30466
rect 37214 30414 37266 30466
rect 37266 30414 37268 30466
rect 37212 30412 37268 30414
rect 37372 30466 37428 30468
rect 37372 30414 37374 30466
rect 37374 30414 37426 30466
rect 37426 30414 37428 30466
rect 37372 30412 37428 30414
rect 37532 30466 37588 30468
rect 37532 30414 37534 30466
rect 37534 30414 37586 30466
rect 37586 30414 37588 30466
rect 37532 30412 37588 30414
rect 37692 30466 37748 30468
rect 37692 30414 37694 30466
rect 37694 30414 37746 30466
rect 37746 30414 37748 30466
rect 37692 30412 37748 30414
rect 37852 30466 37908 30468
rect 37852 30414 37854 30466
rect 37854 30414 37906 30466
rect 37906 30414 37908 30466
rect 37852 30412 37908 30414
rect 38012 30466 38068 30468
rect 38012 30414 38014 30466
rect 38014 30414 38066 30466
rect 38066 30414 38068 30466
rect 38012 30412 38068 30414
rect 38172 30466 38228 30468
rect 38172 30414 38174 30466
rect 38174 30414 38226 30466
rect 38226 30414 38228 30466
rect 38172 30412 38228 30414
rect 38332 30466 38388 30468
rect 38332 30414 38334 30466
rect 38334 30414 38386 30466
rect 38386 30414 38388 30466
rect 38332 30412 38388 30414
rect 38492 30466 38548 30468
rect 38492 30414 38494 30466
rect 38494 30414 38546 30466
rect 38546 30414 38548 30466
rect 38492 30412 38548 30414
rect 38652 30466 38708 30468
rect 38652 30414 38654 30466
rect 38654 30414 38706 30466
rect 38706 30414 38708 30466
rect 38652 30412 38708 30414
rect 38812 30466 38868 30468
rect 38812 30414 38814 30466
rect 38814 30414 38866 30466
rect 38866 30414 38868 30466
rect 38812 30412 38868 30414
rect 38972 30466 39028 30468
rect 38972 30414 38974 30466
rect 38974 30414 39026 30466
rect 39026 30414 39028 30466
rect 38972 30412 39028 30414
rect 39132 30466 39188 30468
rect 39132 30414 39134 30466
rect 39134 30414 39186 30466
rect 39186 30414 39188 30466
rect 39132 30412 39188 30414
rect 39292 30466 39348 30468
rect 39292 30414 39294 30466
rect 39294 30414 39346 30466
rect 39346 30414 39348 30466
rect 39292 30412 39348 30414
rect 39452 30466 39508 30468
rect 39452 30414 39454 30466
rect 39454 30414 39506 30466
rect 39506 30414 39508 30466
rect 39452 30412 39508 30414
rect 39612 30466 39668 30468
rect 39612 30414 39614 30466
rect 39614 30414 39666 30466
rect 39666 30414 39668 30466
rect 39612 30412 39668 30414
rect 39772 30466 39828 30468
rect 39772 30414 39774 30466
rect 39774 30414 39826 30466
rect 39826 30414 39828 30466
rect 39772 30412 39828 30414
rect 39932 30466 39988 30468
rect 39932 30414 39934 30466
rect 39934 30414 39986 30466
rect 39986 30414 39988 30466
rect 39932 30412 39988 30414
rect 40092 30466 40148 30468
rect 40092 30414 40094 30466
rect 40094 30414 40146 30466
rect 40146 30414 40148 30466
rect 40092 30412 40148 30414
rect 40252 30466 40308 30468
rect 40252 30414 40254 30466
rect 40254 30414 40306 30466
rect 40306 30414 40308 30466
rect 40252 30412 40308 30414
rect 40412 30466 40468 30468
rect 40412 30414 40414 30466
rect 40414 30414 40466 30466
rect 40466 30414 40468 30466
rect 40412 30412 40468 30414
rect 40572 30466 40628 30468
rect 40572 30414 40574 30466
rect 40574 30414 40626 30466
rect 40626 30414 40628 30466
rect 40572 30412 40628 30414
rect 40732 30466 40788 30468
rect 40732 30414 40734 30466
rect 40734 30414 40786 30466
rect 40786 30414 40788 30466
rect 40732 30412 40788 30414
rect 40892 30466 40948 30468
rect 40892 30414 40894 30466
rect 40894 30414 40946 30466
rect 40946 30414 40948 30466
rect 40892 30412 40948 30414
rect 41052 30466 41108 30468
rect 41052 30414 41054 30466
rect 41054 30414 41106 30466
rect 41106 30414 41108 30466
rect 41052 30412 41108 30414
rect 41212 30466 41268 30468
rect 41212 30414 41214 30466
rect 41214 30414 41266 30466
rect 41266 30414 41268 30466
rect 41212 30412 41268 30414
rect 41372 30466 41428 30468
rect 41372 30414 41374 30466
rect 41374 30414 41426 30466
rect 41426 30414 41428 30466
rect 41372 30412 41428 30414
rect 41532 30466 41588 30468
rect 41532 30414 41534 30466
rect 41534 30414 41586 30466
rect 41586 30414 41588 30466
rect 41532 30412 41588 30414
rect 41692 30466 41748 30468
rect 41692 30414 41694 30466
rect 41694 30414 41746 30466
rect 41746 30414 41748 30466
rect 41692 30412 41748 30414
rect 41852 30466 41908 30468
rect 41852 30414 41854 30466
rect 41854 30414 41906 30466
rect 41906 30414 41908 30466
rect 41852 30412 41908 30414
rect 12 30306 68 30308
rect 12 30254 14 30306
rect 14 30254 66 30306
rect 66 30254 68 30306
rect 12 30252 68 30254
rect 172 30306 228 30308
rect 172 30254 174 30306
rect 174 30254 226 30306
rect 226 30254 228 30306
rect 172 30252 228 30254
rect 332 30306 388 30308
rect 332 30254 334 30306
rect 334 30254 386 30306
rect 386 30254 388 30306
rect 332 30252 388 30254
rect 492 30306 548 30308
rect 492 30254 494 30306
rect 494 30254 546 30306
rect 546 30254 548 30306
rect 492 30252 548 30254
rect 652 30306 708 30308
rect 652 30254 654 30306
rect 654 30254 706 30306
rect 706 30254 708 30306
rect 652 30252 708 30254
rect 812 30306 868 30308
rect 812 30254 814 30306
rect 814 30254 866 30306
rect 866 30254 868 30306
rect 812 30252 868 30254
rect 972 30306 1028 30308
rect 972 30254 974 30306
rect 974 30254 1026 30306
rect 1026 30254 1028 30306
rect 972 30252 1028 30254
rect 1132 30306 1188 30308
rect 1132 30254 1134 30306
rect 1134 30254 1186 30306
rect 1186 30254 1188 30306
rect 1132 30252 1188 30254
rect 1292 30306 1348 30308
rect 1292 30254 1294 30306
rect 1294 30254 1346 30306
rect 1346 30254 1348 30306
rect 1292 30252 1348 30254
rect 1452 30306 1508 30308
rect 1452 30254 1454 30306
rect 1454 30254 1506 30306
rect 1506 30254 1508 30306
rect 1452 30252 1508 30254
rect 1612 30306 1668 30308
rect 1612 30254 1614 30306
rect 1614 30254 1666 30306
rect 1666 30254 1668 30306
rect 1612 30252 1668 30254
rect 1772 30306 1828 30308
rect 1772 30254 1774 30306
rect 1774 30254 1826 30306
rect 1826 30254 1828 30306
rect 1772 30252 1828 30254
rect 1932 30306 1988 30308
rect 1932 30254 1934 30306
rect 1934 30254 1986 30306
rect 1986 30254 1988 30306
rect 1932 30252 1988 30254
rect 2092 30306 2148 30308
rect 2092 30254 2094 30306
rect 2094 30254 2146 30306
rect 2146 30254 2148 30306
rect 2092 30252 2148 30254
rect 2252 30306 2308 30308
rect 2252 30254 2254 30306
rect 2254 30254 2306 30306
rect 2306 30254 2308 30306
rect 2252 30252 2308 30254
rect 2412 30306 2468 30308
rect 2412 30254 2414 30306
rect 2414 30254 2466 30306
rect 2466 30254 2468 30306
rect 2412 30252 2468 30254
rect 2572 30306 2628 30308
rect 2572 30254 2574 30306
rect 2574 30254 2626 30306
rect 2626 30254 2628 30306
rect 2572 30252 2628 30254
rect 2732 30306 2788 30308
rect 2732 30254 2734 30306
rect 2734 30254 2786 30306
rect 2786 30254 2788 30306
rect 2732 30252 2788 30254
rect 2892 30306 2948 30308
rect 2892 30254 2894 30306
rect 2894 30254 2946 30306
rect 2946 30254 2948 30306
rect 2892 30252 2948 30254
rect 3052 30306 3108 30308
rect 3052 30254 3054 30306
rect 3054 30254 3106 30306
rect 3106 30254 3108 30306
rect 3052 30252 3108 30254
rect 3212 30306 3268 30308
rect 3212 30254 3214 30306
rect 3214 30254 3266 30306
rect 3266 30254 3268 30306
rect 3212 30252 3268 30254
rect 3372 30306 3428 30308
rect 3372 30254 3374 30306
rect 3374 30254 3426 30306
rect 3426 30254 3428 30306
rect 3372 30252 3428 30254
rect 3532 30306 3588 30308
rect 3532 30254 3534 30306
rect 3534 30254 3586 30306
rect 3586 30254 3588 30306
rect 3532 30252 3588 30254
rect 3692 30306 3748 30308
rect 3692 30254 3694 30306
rect 3694 30254 3746 30306
rect 3746 30254 3748 30306
rect 3692 30252 3748 30254
rect 3852 30306 3908 30308
rect 3852 30254 3854 30306
rect 3854 30254 3906 30306
rect 3906 30254 3908 30306
rect 3852 30252 3908 30254
rect 4012 30306 4068 30308
rect 4012 30254 4014 30306
rect 4014 30254 4066 30306
rect 4066 30254 4068 30306
rect 4012 30252 4068 30254
rect 4172 30306 4228 30308
rect 4172 30254 4174 30306
rect 4174 30254 4226 30306
rect 4226 30254 4228 30306
rect 4172 30252 4228 30254
rect 4332 30306 4388 30308
rect 4332 30254 4334 30306
rect 4334 30254 4386 30306
rect 4386 30254 4388 30306
rect 4332 30252 4388 30254
rect 4492 30306 4548 30308
rect 4492 30254 4494 30306
rect 4494 30254 4546 30306
rect 4546 30254 4548 30306
rect 4492 30252 4548 30254
rect 4652 30306 4708 30308
rect 4652 30254 4654 30306
rect 4654 30254 4706 30306
rect 4706 30254 4708 30306
rect 4652 30252 4708 30254
rect 4812 30306 4868 30308
rect 4812 30254 4814 30306
rect 4814 30254 4866 30306
rect 4866 30254 4868 30306
rect 4812 30252 4868 30254
rect 4972 30306 5028 30308
rect 4972 30254 4974 30306
rect 4974 30254 5026 30306
rect 5026 30254 5028 30306
rect 4972 30252 5028 30254
rect 5132 30306 5188 30308
rect 5132 30254 5134 30306
rect 5134 30254 5186 30306
rect 5186 30254 5188 30306
rect 5132 30252 5188 30254
rect 5292 30306 5348 30308
rect 5292 30254 5294 30306
rect 5294 30254 5346 30306
rect 5346 30254 5348 30306
rect 5292 30252 5348 30254
rect 5452 30306 5508 30308
rect 5452 30254 5454 30306
rect 5454 30254 5506 30306
rect 5506 30254 5508 30306
rect 5452 30252 5508 30254
rect 5612 30306 5668 30308
rect 5612 30254 5614 30306
rect 5614 30254 5666 30306
rect 5666 30254 5668 30306
rect 5612 30252 5668 30254
rect 5772 30306 5828 30308
rect 5772 30254 5774 30306
rect 5774 30254 5826 30306
rect 5826 30254 5828 30306
rect 5772 30252 5828 30254
rect 5932 30306 5988 30308
rect 5932 30254 5934 30306
rect 5934 30254 5986 30306
rect 5986 30254 5988 30306
rect 5932 30252 5988 30254
rect 6092 30306 6148 30308
rect 6092 30254 6094 30306
rect 6094 30254 6146 30306
rect 6146 30254 6148 30306
rect 6092 30252 6148 30254
rect 6252 30306 6308 30308
rect 6252 30254 6254 30306
rect 6254 30254 6306 30306
rect 6306 30254 6308 30306
rect 6252 30252 6308 30254
rect 6412 30306 6468 30308
rect 6412 30254 6414 30306
rect 6414 30254 6466 30306
rect 6466 30254 6468 30306
rect 6412 30252 6468 30254
rect 6572 30306 6628 30308
rect 6572 30254 6574 30306
rect 6574 30254 6626 30306
rect 6626 30254 6628 30306
rect 6572 30252 6628 30254
rect 6732 30306 6788 30308
rect 6732 30254 6734 30306
rect 6734 30254 6786 30306
rect 6786 30254 6788 30306
rect 6732 30252 6788 30254
rect 6892 30306 6948 30308
rect 6892 30254 6894 30306
rect 6894 30254 6946 30306
rect 6946 30254 6948 30306
rect 6892 30252 6948 30254
rect 7052 30306 7108 30308
rect 7052 30254 7054 30306
rect 7054 30254 7106 30306
rect 7106 30254 7108 30306
rect 7052 30252 7108 30254
rect 7212 30306 7268 30308
rect 7212 30254 7214 30306
rect 7214 30254 7266 30306
rect 7266 30254 7268 30306
rect 7212 30252 7268 30254
rect 7372 30306 7428 30308
rect 7372 30254 7374 30306
rect 7374 30254 7426 30306
rect 7426 30254 7428 30306
rect 7372 30252 7428 30254
rect 7532 30306 7588 30308
rect 7532 30254 7534 30306
rect 7534 30254 7586 30306
rect 7586 30254 7588 30306
rect 7532 30252 7588 30254
rect 7692 30306 7748 30308
rect 7692 30254 7694 30306
rect 7694 30254 7746 30306
rect 7746 30254 7748 30306
rect 7692 30252 7748 30254
rect 7852 30306 7908 30308
rect 7852 30254 7854 30306
rect 7854 30254 7906 30306
rect 7906 30254 7908 30306
rect 7852 30252 7908 30254
rect 8012 30306 8068 30308
rect 8012 30254 8014 30306
rect 8014 30254 8066 30306
rect 8066 30254 8068 30306
rect 8012 30252 8068 30254
rect 8172 30306 8228 30308
rect 8172 30254 8174 30306
rect 8174 30254 8226 30306
rect 8226 30254 8228 30306
rect 8172 30252 8228 30254
rect 8332 30306 8388 30308
rect 8332 30254 8334 30306
rect 8334 30254 8386 30306
rect 8386 30254 8388 30306
rect 8332 30252 8388 30254
rect 11532 30252 11588 30308
rect 11852 30252 11908 30308
rect 12492 30306 12548 30308
rect 12492 30254 12494 30306
rect 12494 30254 12546 30306
rect 12546 30254 12548 30306
rect 12492 30252 12548 30254
rect 12652 30306 12708 30308
rect 12652 30254 12654 30306
rect 12654 30254 12706 30306
rect 12706 30254 12708 30306
rect 12652 30252 12708 30254
rect 12812 30306 12868 30308
rect 12812 30254 12814 30306
rect 12814 30254 12866 30306
rect 12866 30254 12868 30306
rect 12812 30252 12868 30254
rect 12972 30306 13028 30308
rect 12972 30254 12974 30306
rect 12974 30254 13026 30306
rect 13026 30254 13028 30306
rect 12972 30252 13028 30254
rect 13132 30306 13188 30308
rect 13132 30254 13134 30306
rect 13134 30254 13186 30306
rect 13186 30254 13188 30306
rect 13132 30252 13188 30254
rect 13292 30306 13348 30308
rect 13292 30254 13294 30306
rect 13294 30254 13346 30306
rect 13346 30254 13348 30306
rect 13292 30252 13348 30254
rect 13452 30306 13508 30308
rect 13452 30254 13454 30306
rect 13454 30254 13506 30306
rect 13506 30254 13508 30306
rect 13452 30252 13508 30254
rect 13612 30306 13668 30308
rect 13612 30254 13614 30306
rect 13614 30254 13666 30306
rect 13666 30254 13668 30306
rect 13612 30252 13668 30254
rect 13772 30306 13828 30308
rect 13772 30254 13774 30306
rect 13774 30254 13826 30306
rect 13826 30254 13828 30306
rect 13772 30252 13828 30254
rect 13932 30306 13988 30308
rect 13932 30254 13934 30306
rect 13934 30254 13986 30306
rect 13986 30254 13988 30306
rect 13932 30252 13988 30254
rect 14092 30306 14148 30308
rect 14092 30254 14094 30306
rect 14094 30254 14146 30306
rect 14146 30254 14148 30306
rect 14092 30252 14148 30254
rect 14252 30306 14308 30308
rect 14252 30254 14254 30306
rect 14254 30254 14306 30306
rect 14306 30254 14308 30306
rect 14252 30252 14308 30254
rect 14412 30306 14468 30308
rect 14412 30254 14414 30306
rect 14414 30254 14466 30306
rect 14466 30254 14468 30306
rect 14412 30252 14468 30254
rect 14572 30306 14628 30308
rect 14572 30254 14574 30306
rect 14574 30254 14626 30306
rect 14626 30254 14628 30306
rect 14572 30252 14628 30254
rect 14732 30306 14788 30308
rect 14732 30254 14734 30306
rect 14734 30254 14786 30306
rect 14786 30254 14788 30306
rect 14732 30252 14788 30254
rect 14892 30306 14948 30308
rect 14892 30254 14894 30306
rect 14894 30254 14946 30306
rect 14946 30254 14948 30306
rect 14892 30252 14948 30254
rect 15052 30306 15108 30308
rect 15052 30254 15054 30306
rect 15054 30254 15106 30306
rect 15106 30254 15108 30306
rect 15052 30252 15108 30254
rect 15212 30306 15268 30308
rect 15212 30254 15214 30306
rect 15214 30254 15266 30306
rect 15266 30254 15268 30306
rect 15212 30252 15268 30254
rect 15372 30306 15428 30308
rect 15372 30254 15374 30306
rect 15374 30254 15426 30306
rect 15426 30254 15428 30306
rect 15372 30252 15428 30254
rect 15532 30306 15588 30308
rect 15532 30254 15534 30306
rect 15534 30254 15586 30306
rect 15586 30254 15588 30306
rect 15532 30252 15588 30254
rect 15692 30306 15748 30308
rect 15692 30254 15694 30306
rect 15694 30254 15746 30306
rect 15746 30254 15748 30306
rect 15692 30252 15748 30254
rect 15852 30306 15908 30308
rect 15852 30254 15854 30306
rect 15854 30254 15906 30306
rect 15906 30254 15908 30306
rect 15852 30252 15908 30254
rect 16012 30306 16068 30308
rect 16012 30254 16014 30306
rect 16014 30254 16066 30306
rect 16066 30254 16068 30306
rect 16012 30252 16068 30254
rect 16172 30306 16228 30308
rect 16172 30254 16174 30306
rect 16174 30254 16226 30306
rect 16226 30254 16228 30306
rect 16172 30252 16228 30254
rect 16332 30306 16388 30308
rect 16332 30254 16334 30306
rect 16334 30254 16386 30306
rect 16386 30254 16388 30306
rect 16332 30252 16388 30254
rect 16492 30306 16548 30308
rect 16492 30254 16494 30306
rect 16494 30254 16546 30306
rect 16546 30254 16548 30306
rect 16492 30252 16548 30254
rect 16652 30306 16708 30308
rect 16652 30254 16654 30306
rect 16654 30254 16706 30306
rect 16706 30254 16708 30306
rect 16652 30252 16708 30254
rect 16812 30306 16868 30308
rect 16812 30254 16814 30306
rect 16814 30254 16866 30306
rect 16866 30254 16868 30306
rect 16812 30252 16868 30254
rect 16972 30306 17028 30308
rect 16972 30254 16974 30306
rect 16974 30254 17026 30306
rect 17026 30254 17028 30306
rect 16972 30252 17028 30254
rect 17132 30306 17188 30308
rect 17132 30254 17134 30306
rect 17134 30254 17186 30306
rect 17186 30254 17188 30306
rect 17132 30252 17188 30254
rect 17292 30306 17348 30308
rect 17292 30254 17294 30306
rect 17294 30254 17346 30306
rect 17346 30254 17348 30306
rect 17292 30252 17348 30254
rect 17452 30306 17508 30308
rect 17452 30254 17454 30306
rect 17454 30254 17506 30306
rect 17506 30254 17508 30306
rect 17452 30252 17508 30254
rect 17612 30306 17668 30308
rect 17612 30254 17614 30306
rect 17614 30254 17666 30306
rect 17666 30254 17668 30306
rect 17612 30252 17668 30254
rect 17772 30306 17828 30308
rect 17772 30254 17774 30306
rect 17774 30254 17826 30306
rect 17826 30254 17828 30306
rect 17772 30252 17828 30254
rect 17932 30306 17988 30308
rect 17932 30254 17934 30306
rect 17934 30254 17986 30306
rect 17986 30254 17988 30306
rect 17932 30252 17988 30254
rect 18092 30306 18148 30308
rect 18092 30254 18094 30306
rect 18094 30254 18146 30306
rect 18146 30254 18148 30306
rect 18092 30252 18148 30254
rect 18252 30306 18308 30308
rect 18252 30254 18254 30306
rect 18254 30254 18306 30306
rect 18306 30254 18308 30306
rect 18252 30252 18308 30254
rect 18412 30306 18468 30308
rect 18412 30254 18414 30306
rect 18414 30254 18466 30306
rect 18466 30254 18468 30306
rect 18412 30252 18468 30254
rect 18572 30306 18628 30308
rect 18572 30254 18574 30306
rect 18574 30254 18626 30306
rect 18626 30254 18628 30306
rect 18572 30252 18628 30254
rect 18732 30306 18788 30308
rect 18732 30254 18734 30306
rect 18734 30254 18786 30306
rect 18786 30254 18788 30306
rect 18732 30252 18788 30254
rect 18892 30306 18948 30308
rect 18892 30254 18894 30306
rect 18894 30254 18946 30306
rect 18946 30254 18948 30306
rect 18892 30252 18948 30254
rect 22092 30252 22148 30308
rect 22412 30252 22468 30308
rect 23132 30306 23188 30308
rect 23132 30254 23134 30306
rect 23134 30254 23186 30306
rect 23186 30254 23188 30306
rect 23132 30252 23188 30254
rect 23292 30306 23348 30308
rect 23292 30254 23294 30306
rect 23294 30254 23346 30306
rect 23346 30254 23348 30306
rect 23292 30252 23348 30254
rect 23452 30306 23508 30308
rect 23452 30254 23454 30306
rect 23454 30254 23506 30306
rect 23506 30254 23508 30306
rect 23452 30252 23508 30254
rect 23612 30306 23668 30308
rect 23612 30254 23614 30306
rect 23614 30254 23666 30306
rect 23666 30254 23668 30306
rect 23612 30252 23668 30254
rect 23772 30306 23828 30308
rect 23772 30254 23774 30306
rect 23774 30254 23826 30306
rect 23826 30254 23828 30306
rect 23772 30252 23828 30254
rect 23932 30306 23988 30308
rect 23932 30254 23934 30306
rect 23934 30254 23986 30306
rect 23986 30254 23988 30306
rect 23932 30252 23988 30254
rect 24092 30306 24148 30308
rect 24092 30254 24094 30306
rect 24094 30254 24146 30306
rect 24146 30254 24148 30306
rect 24092 30252 24148 30254
rect 24252 30306 24308 30308
rect 24252 30254 24254 30306
rect 24254 30254 24306 30306
rect 24306 30254 24308 30306
rect 24252 30252 24308 30254
rect 24412 30306 24468 30308
rect 24412 30254 24414 30306
rect 24414 30254 24466 30306
rect 24466 30254 24468 30306
rect 24412 30252 24468 30254
rect 24572 30306 24628 30308
rect 24572 30254 24574 30306
rect 24574 30254 24626 30306
rect 24626 30254 24628 30306
rect 24572 30252 24628 30254
rect 24732 30306 24788 30308
rect 24732 30254 24734 30306
rect 24734 30254 24786 30306
rect 24786 30254 24788 30306
rect 24732 30252 24788 30254
rect 24892 30306 24948 30308
rect 24892 30254 24894 30306
rect 24894 30254 24946 30306
rect 24946 30254 24948 30306
rect 24892 30252 24948 30254
rect 25052 30306 25108 30308
rect 25052 30254 25054 30306
rect 25054 30254 25106 30306
rect 25106 30254 25108 30306
rect 25052 30252 25108 30254
rect 25212 30306 25268 30308
rect 25212 30254 25214 30306
rect 25214 30254 25266 30306
rect 25266 30254 25268 30306
rect 25212 30252 25268 30254
rect 25372 30306 25428 30308
rect 25372 30254 25374 30306
rect 25374 30254 25426 30306
rect 25426 30254 25428 30306
rect 25372 30252 25428 30254
rect 25532 30306 25588 30308
rect 25532 30254 25534 30306
rect 25534 30254 25586 30306
rect 25586 30254 25588 30306
rect 25532 30252 25588 30254
rect 25692 30306 25748 30308
rect 25692 30254 25694 30306
rect 25694 30254 25746 30306
rect 25746 30254 25748 30306
rect 25692 30252 25748 30254
rect 25852 30306 25908 30308
rect 25852 30254 25854 30306
rect 25854 30254 25906 30306
rect 25906 30254 25908 30306
rect 25852 30252 25908 30254
rect 26012 30306 26068 30308
rect 26012 30254 26014 30306
rect 26014 30254 26066 30306
rect 26066 30254 26068 30306
rect 26012 30252 26068 30254
rect 26172 30306 26228 30308
rect 26172 30254 26174 30306
rect 26174 30254 26226 30306
rect 26226 30254 26228 30306
rect 26172 30252 26228 30254
rect 26332 30306 26388 30308
rect 26332 30254 26334 30306
rect 26334 30254 26386 30306
rect 26386 30254 26388 30306
rect 26332 30252 26388 30254
rect 26492 30306 26548 30308
rect 26492 30254 26494 30306
rect 26494 30254 26546 30306
rect 26546 30254 26548 30306
rect 26492 30252 26548 30254
rect 26652 30306 26708 30308
rect 26652 30254 26654 30306
rect 26654 30254 26706 30306
rect 26706 30254 26708 30306
rect 26652 30252 26708 30254
rect 26812 30306 26868 30308
rect 26812 30254 26814 30306
rect 26814 30254 26866 30306
rect 26866 30254 26868 30306
rect 26812 30252 26868 30254
rect 26972 30306 27028 30308
rect 26972 30254 26974 30306
rect 26974 30254 27026 30306
rect 27026 30254 27028 30306
rect 26972 30252 27028 30254
rect 27132 30306 27188 30308
rect 27132 30254 27134 30306
rect 27134 30254 27186 30306
rect 27186 30254 27188 30306
rect 27132 30252 27188 30254
rect 27292 30306 27348 30308
rect 27292 30254 27294 30306
rect 27294 30254 27346 30306
rect 27346 30254 27348 30306
rect 27292 30252 27348 30254
rect 27452 30306 27508 30308
rect 27452 30254 27454 30306
rect 27454 30254 27506 30306
rect 27506 30254 27508 30306
rect 27452 30252 27508 30254
rect 27612 30306 27668 30308
rect 27612 30254 27614 30306
rect 27614 30254 27666 30306
rect 27666 30254 27668 30306
rect 27612 30252 27668 30254
rect 27772 30306 27828 30308
rect 27772 30254 27774 30306
rect 27774 30254 27826 30306
rect 27826 30254 27828 30306
rect 27772 30252 27828 30254
rect 27932 30306 27988 30308
rect 27932 30254 27934 30306
rect 27934 30254 27986 30306
rect 27986 30254 27988 30306
rect 27932 30252 27988 30254
rect 28092 30306 28148 30308
rect 28092 30254 28094 30306
rect 28094 30254 28146 30306
rect 28146 30254 28148 30306
rect 28092 30252 28148 30254
rect 28252 30306 28308 30308
rect 28252 30254 28254 30306
rect 28254 30254 28306 30306
rect 28306 30254 28308 30306
rect 28252 30252 28308 30254
rect 28412 30306 28468 30308
rect 28412 30254 28414 30306
rect 28414 30254 28466 30306
rect 28466 30254 28468 30306
rect 28412 30252 28468 30254
rect 28572 30306 28628 30308
rect 28572 30254 28574 30306
rect 28574 30254 28626 30306
rect 28626 30254 28628 30306
rect 28572 30252 28628 30254
rect 28732 30306 28788 30308
rect 28732 30254 28734 30306
rect 28734 30254 28786 30306
rect 28786 30254 28788 30306
rect 28732 30252 28788 30254
rect 28892 30306 28948 30308
rect 28892 30254 28894 30306
rect 28894 30254 28946 30306
rect 28946 30254 28948 30306
rect 28892 30252 28948 30254
rect 29052 30306 29108 30308
rect 29052 30254 29054 30306
rect 29054 30254 29106 30306
rect 29106 30254 29108 30306
rect 29052 30252 29108 30254
rect 29212 30306 29268 30308
rect 29212 30254 29214 30306
rect 29214 30254 29266 30306
rect 29266 30254 29268 30306
rect 29212 30252 29268 30254
rect 29372 30306 29428 30308
rect 29372 30254 29374 30306
rect 29374 30254 29426 30306
rect 29426 30254 29428 30306
rect 29372 30252 29428 30254
rect 30012 30252 30068 30308
rect 30332 30252 30388 30308
rect 33532 30306 33588 30308
rect 33532 30254 33534 30306
rect 33534 30254 33586 30306
rect 33586 30254 33588 30306
rect 33532 30252 33588 30254
rect 33692 30306 33748 30308
rect 33692 30254 33694 30306
rect 33694 30254 33746 30306
rect 33746 30254 33748 30306
rect 33692 30252 33748 30254
rect 33852 30306 33908 30308
rect 33852 30254 33854 30306
rect 33854 30254 33906 30306
rect 33906 30254 33908 30306
rect 33852 30252 33908 30254
rect 34012 30306 34068 30308
rect 34012 30254 34014 30306
rect 34014 30254 34066 30306
rect 34066 30254 34068 30306
rect 34012 30252 34068 30254
rect 34172 30306 34228 30308
rect 34172 30254 34174 30306
rect 34174 30254 34226 30306
rect 34226 30254 34228 30306
rect 34172 30252 34228 30254
rect 34332 30306 34388 30308
rect 34332 30254 34334 30306
rect 34334 30254 34386 30306
rect 34386 30254 34388 30306
rect 34332 30252 34388 30254
rect 34492 30306 34548 30308
rect 34492 30254 34494 30306
rect 34494 30254 34546 30306
rect 34546 30254 34548 30306
rect 34492 30252 34548 30254
rect 34652 30306 34708 30308
rect 34652 30254 34654 30306
rect 34654 30254 34706 30306
rect 34706 30254 34708 30306
rect 34652 30252 34708 30254
rect 34812 30306 34868 30308
rect 34812 30254 34814 30306
rect 34814 30254 34866 30306
rect 34866 30254 34868 30306
rect 34812 30252 34868 30254
rect 34972 30306 35028 30308
rect 34972 30254 34974 30306
rect 34974 30254 35026 30306
rect 35026 30254 35028 30306
rect 34972 30252 35028 30254
rect 35132 30306 35188 30308
rect 35132 30254 35134 30306
rect 35134 30254 35186 30306
rect 35186 30254 35188 30306
rect 35132 30252 35188 30254
rect 35292 30306 35348 30308
rect 35292 30254 35294 30306
rect 35294 30254 35346 30306
rect 35346 30254 35348 30306
rect 35292 30252 35348 30254
rect 35452 30306 35508 30308
rect 35452 30254 35454 30306
rect 35454 30254 35506 30306
rect 35506 30254 35508 30306
rect 35452 30252 35508 30254
rect 35612 30306 35668 30308
rect 35612 30254 35614 30306
rect 35614 30254 35666 30306
rect 35666 30254 35668 30306
rect 35612 30252 35668 30254
rect 35772 30306 35828 30308
rect 35772 30254 35774 30306
rect 35774 30254 35826 30306
rect 35826 30254 35828 30306
rect 35772 30252 35828 30254
rect 35932 30306 35988 30308
rect 35932 30254 35934 30306
rect 35934 30254 35986 30306
rect 35986 30254 35988 30306
rect 35932 30252 35988 30254
rect 36092 30306 36148 30308
rect 36092 30254 36094 30306
rect 36094 30254 36146 30306
rect 36146 30254 36148 30306
rect 36092 30252 36148 30254
rect 36252 30306 36308 30308
rect 36252 30254 36254 30306
rect 36254 30254 36306 30306
rect 36306 30254 36308 30306
rect 36252 30252 36308 30254
rect 36412 30306 36468 30308
rect 36412 30254 36414 30306
rect 36414 30254 36466 30306
rect 36466 30254 36468 30306
rect 36412 30252 36468 30254
rect 36572 30306 36628 30308
rect 36572 30254 36574 30306
rect 36574 30254 36626 30306
rect 36626 30254 36628 30306
rect 36572 30252 36628 30254
rect 36732 30306 36788 30308
rect 36732 30254 36734 30306
rect 36734 30254 36786 30306
rect 36786 30254 36788 30306
rect 36732 30252 36788 30254
rect 36892 30306 36948 30308
rect 36892 30254 36894 30306
rect 36894 30254 36946 30306
rect 36946 30254 36948 30306
rect 36892 30252 36948 30254
rect 37052 30306 37108 30308
rect 37052 30254 37054 30306
rect 37054 30254 37106 30306
rect 37106 30254 37108 30306
rect 37052 30252 37108 30254
rect 37212 30306 37268 30308
rect 37212 30254 37214 30306
rect 37214 30254 37266 30306
rect 37266 30254 37268 30306
rect 37212 30252 37268 30254
rect 37372 30306 37428 30308
rect 37372 30254 37374 30306
rect 37374 30254 37426 30306
rect 37426 30254 37428 30306
rect 37372 30252 37428 30254
rect 37532 30306 37588 30308
rect 37532 30254 37534 30306
rect 37534 30254 37586 30306
rect 37586 30254 37588 30306
rect 37532 30252 37588 30254
rect 37692 30306 37748 30308
rect 37692 30254 37694 30306
rect 37694 30254 37746 30306
rect 37746 30254 37748 30306
rect 37692 30252 37748 30254
rect 37852 30306 37908 30308
rect 37852 30254 37854 30306
rect 37854 30254 37906 30306
rect 37906 30254 37908 30306
rect 37852 30252 37908 30254
rect 38012 30306 38068 30308
rect 38012 30254 38014 30306
rect 38014 30254 38066 30306
rect 38066 30254 38068 30306
rect 38012 30252 38068 30254
rect 38172 30306 38228 30308
rect 38172 30254 38174 30306
rect 38174 30254 38226 30306
rect 38226 30254 38228 30306
rect 38172 30252 38228 30254
rect 38332 30306 38388 30308
rect 38332 30254 38334 30306
rect 38334 30254 38386 30306
rect 38386 30254 38388 30306
rect 38332 30252 38388 30254
rect 38492 30306 38548 30308
rect 38492 30254 38494 30306
rect 38494 30254 38546 30306
rect 38546 30254 38548 30306
rect 38492 30252 38548 30254
rect 38652 30306 38708 30308
rect 38652 30254 38654 30306
rect 38654 30254 38706 30306
rect 38706 30254 38708 30306
rect 38652 30252 38708 30254
rect 38812 30306 38868 30308
rect 38812 30254 38814 30306
rect 38814 30254 38866 30306
rect 38866 30254 38868 30306
rect 38812 30252 38868 30254
rect 38972 30306 39028 30308
rect 38972 30254 38974 30306
rect 38974 30254 39026 30306
rect 39026 30254 39028 30306
rect 38972 30252 39028 30254
rect 39132 30306 39188 30308
rect 39132 30254 39134 30306
rect 39134 30254 39186 30306
rect 39186 30254 39188 30306
rect 39132 30252 39188 30254
rect 39292 30306 39348 30308
rect 39292 30254 39294 30306
rect 39294 30254 39346 30306
rect 39346 30254 39348 30306
rect 39292 30252 39348 30254
rect 39452 30306 39508 30308
rect 39452 30254 39454 30306
rect 39454 30254 39506 30306
rect 39506 30254 39508 30306
rect 39452 30252 39508 30254
rect 39612 30306 39668 30308
rect 39612 30254 39614 30306
rect 39614 30254 39666 30306
rect 39666 30254 39668 30306
rect 39612 30252 39668 30254
rect 39772 30306 39828 30308
rect 39772 30254 39774 30306
rect 39774 30254 39826 30306
rect 39826 30254 39828 30306
rect 39772 30252 39828 30254
rect 39932 30306 39988 30308
rect 39932 30254 39934 30306
rect 39934 30254 39986 30306
rect 39986 30254 39988 30306
rect 39932 30252 39988 30254
rect 40092 30306 40148 30308
rect 40092 30254 40094 30306
rect 40094 30254 40146 30306
rect 40146 30254 40148 30306
rect 40092 30252 40148 30254
rect 40252 30306 40308 30308
rect 40252 30254 40254 30306
rect 40254 30254 40306 30306
rect 40306 30254 40308 30306
rect 40252 30252 40308 30254
rect 40412 30306 40468 30308
rect 40412 30254 40414 30306
rect 40414 30254 40466 30306
rect 40466 30254 40468 30306
rect 40412 30252 40468 30254
rect 40572 30306 40628 30308
rect 40572 30254 40574 30306
rect 40574 30254 40626 30306
rect 40626 30254 40628 30306
rect 40572 30252 40628 30254
rect 40732 30306 40788 30308
rect 40732 30254 40734 30306
rect 40734 30254 40786 30306
rect 40786 30254 40788 30306
rect 40732 30252 40788 30254
rect 40892 30306 40948 30308
rect 40892 30254 40894 30306
rect 40894 30254 40946 30306
rect 40946 30254 40948 30306
rect 40892 30252 40948 30254
rect 41052 30306 41108 30308
rect 41052 30254 41054 30306
rect 41054 30254 41106 30306
rect 41106 30254 41108 30306
rect 41052 30252 41108 30254
rect 41212 30306 41268 30308
rect 41212 30254 41214 30306
rect 41214 30254 41266 30306
rect 41266 30254 41268 30306
rect 41212 30252 41268 30254
rect 41372 30306 41428 30308
rect 41372 30254 41374 30306
rect 41374 30254 41426 30306
rect 41426 30254 41428 30306
rect 41372 30252 41428 30254
rect 41532 30306 41588 30308
rect 41532 30254 41534 30306
rect 41534 30254 41586 30306
rect 41586 30254 41588 30306
rect 41532 30252 41588 30254
rect 41692 30306 41748 30308
rect 41692 30254 41694 30306
rect 41694 30254 41746 30306
rect 41746 30254 41748 30306
rect 41692 30252 41748 30254
rect 41852 30306 41908 30308
rect 41852 30254 41854 30306
rect 41854 30254 41906 30306
rect 41906 30254 41908 30306
rect 41852 30252 41908 30254
rect 11692 30092 11748 30148
rect 22252 30092 22308 30148
rect 30172 30092 30228 30148
rect 12 29986 68 29988
rect 12 29934 14 29986
rect 14 29934 66 29986
rect 66 29934 68 29986
rect 12 29932 68 29934
rect 172 29986 228 29988
rect 172 29934 174 29986
rect 174 29934 226 29986
rect 226 29934 228 29986
rect 172 29932 228 29934
rect 332 29986 388 29988
rect 332 29934 334 29986
rect 334 29934 386 29986
rect 386 29934 388 29986
rect 332 29932 388 29934
rect 492 29986 548 29988
rect 492 29934 494 29986
rect 494 29934 546 29986
rect 546 29934 548 29986
rect 492 29932 548 29934
rect 652 29986 708 29988
rect 652 29934 654 29986
rect 654 29934 706 29986
rect 706 29934 708 29986
rect 652 29932 708 29934
rect 812 29986 868 29988
rect 812 29934 814 29986
rect 814 29934 866 29986
rect 866 29934 868 29986
rect 812 29932 868 29934
rect 972 29986 1028 29988
rect 972 29934 974 29986
rect 974 29934 1026 29986
rect 1026 29934 1028 29986
rect 972 29932 1028 29934
rect 1132 29986 1188 29988
rect 1132 29934 1134 29986
rect 1134 29934 1186 29986
rect 1186 29934 1188 29986
rect 1132 29932 1188 29934
rect 1292 29986 1348 29988
rect 1292 29934 1294 29986
rect 1294 29934 1346 29986
rect 1346 29934 1348 29986
rect 1292 29932 1348 29934
rect 1452 29986 1508 29988
rect 1452 29934 1454 29986
rect 1454 29934 1506 29986
rect 1506 29934 1508 29986
rect 1452 29932 1508 29934
rect 1612 29986 1668 29988
rect 1612 29934 1614 29986
rect 1614 29934 1666 29986
rect 1666 29934 1668 29986
rect 1612 29932 1668 29934
rect 1772 29986 1828 29988
rect 1772 29934 1774 29986
rect 1774 29934 1826 29986
rect 1826 29934 1828 29986
rect 1772 29932 1828 29934
rect 1932 29986 1988 29988
rect 1932 29934 1934 29986
rect 1934 29934 1986 29986
rect 1986 29934 1988 29986
rect 1932 29932 1988 29934
rect 2092 29986 2148 29988
rect 2092 29934 2094 29986
rect 2094 29934 2146 29986
rect 2146 29934 2148 29986
rect 2092 29932 2148 29934
rect 2252 29986 2308 29988
rect 2252 29934 2254 29986
rect 2254 29934 2306 29986
rect 2306 29934 2308 29986
rect 2252 29932 2308 29934
rect 2412 29986 2468 29988
rect 2412 29934 2414 29986
rect 2414 29934 2466 29986
rect 2466 29934 2468 29986
rect 2412 29932 2468 29934
rect 2572 29986 2628 29988
rect 2572 29934 2574 29986
rect 2574 29934 2626 29986
rect 2626 29934 2628 29986
rect 2572 29932 2628 29934
rect 2732 29986 2788 29988
rect 2732 29934 2734 29986
rect 2734 29934 2786 29986
rect 2786 29934 2788 29986
rect 2732 29932 2788 29934
rect 2892 29986 2948 29988
rect 2892 29934 2894 29986
rect 2894 29934 2946 29986
rect 2946 29934 2948 29986
rect 2892 29932 2948 29934
rect 3052 29986 3108 29988
rect 3052 29934 3054 29986
rect 3054 29934 3106 29986
rect 3106 29934 3108 29986
rect 3052 29932 3108 29934
rect 3212 29986 3268 29988
rect 3212 29934 3214 29986
rect 3214 29934 3266 29986
rect 3266 29934 3268 29986
rect 3212 29932 3268 29934
rect 3372 29986 3428 29988
rect 3372 29934 3374 29986
rect 3374 29934 3426 29986
rect 3426 29934 3428 29986
rect 3372 29932 3428 29934
rect 3532 29986 3588 29988
rect 3532 29934 3534 29986
rect 3534 29934 3586 29986
rect 3586 29934 3588 29986
rect 3532 29932 3588 29934
rect 3692 29986 3748 29988
rect 3692 29934 3694 29986
rect 3694 29934 3746 29986
rect 3746 29934 3748 29986
rect 3692 29932 3748 29934
rect 3852 29986 3908 29988
rect 3852 29934 3854 29986
rect 3854 29934 3906 29986
rect 3906 29934 3908 29986
rect 3852 29932 3908 29934
rect 4012 29986 4068 29988
rect 4012 29934 4014 29986
rect 4014 29934 4066 29986
rect 4066 29934 4068 29986
rect 4012 29932 4068 29934
rect 4172 29986 4228 29988
rect 4172 29934 4174 29986
rect 4174 29934 4226 29986
rect 4226 29934 4228 29986
rect 4172 29932 4228 29934
rect 4332 29986 4388 29988
rect 4332 29934 4334 29986
rect 4334 29934 4386 29986
rect 4386 29934 4388 29986
rect 4332 29932 4388 29934
rect 4492 29986 4548 29988
rect 4492 29934 4494 29986
rect 4494 29934 4546 29986
rect 4546 29934 4548 29986
rect 4492 29932 4548 29934
rect 4652 29986 4708 29988
rect 4652 29934 4654 29986
rect 4654 29934 4706 29986
rect 4706 29934 4708 29986
rect 4652 29932 4708 29934
rect 4812 29986 4868 29988
rect 4812 29934 4814 29986
rect 4814 29934 4866 29986
rect 4866 29934 4868 29986
rect 4812 29932 4868 29934
rect 4972 29986 5028 29988
rect 4972 29934 4974 29986
rect 4974 29934 5026 29986
rect 5026 29934 5028 29986
rect 4972 29932 5028 29934
rect 5132 29986 5188 29988
rect 5132 29934 5134 29986
rect 5134 29934 5186 29986
rect 5186 29934 5188 29986
rect 5132 29932 5188 29934
rect 5292 29986 5348 29988
rect 5292 29934 5294 29986
rect 5294 29934 5346 29986
rect 5346 29934 5348 29986
rect 5292 29932 5348 29934
rect 5452 29986 5508 29988
rect 5452 29934 5454 29986
rect 5454 29934 5506 29986
rect 5506 29934 5508 29986
rect 5452 29932 5508 29934
rect 5612 29986 5668 29988
rect 5612 29934 5614 29986
rect 5614 29934 5666 29986
rect 5666 29934 5668 29986
rect 5612 29932 5668 29934
rect 5772 29986 5828 29988
rect 5772 29934 5774 29986
rect 5774 29934 5826 29986
rect 5826 29934 5828 29986
rect 5772 29932 5828 29934
rect 5932 29986 5988 29988
rect 5932 29934 5934 29986
rect 5934 29934 5986 29986
rect 5986 29934 5988 29986
rect 5932 29932 5988 29934
rect 6092 29986 6148 29988
rect 6092 29934 6094 29986
rect 6094 29934 6146 29986
rect 6146 29934 6148 29986
rect 6092 29932 6148 29934
rect 6252 29986 6308 29988
rect 6252 29934 6254 29986
rect 6254 29934 6306 29986
rect 6306 29934 6308 29986
rect 6252 29932 6308 29934
rect 6412 29986 6468 29988
rect 6412 29934 6414 29986
rect 6414 29934 6466 29986
rect 6466 29934 6468 29986
rect 6412 29932 6468 29934
rect 6572 29986 6628 29988
rect 6572 29934 6574 29986
rect 6574 29934 6626 29986
rect 6626 29934 6628 29986
rect 6572 29932 6628 29934
rect 6732 29986 6788 29988
rect 6732 29934 6734 29986
rect 6734 29934 6786 29986
rect 6786 29934 6788 29986
rect 6732 29932 6788 29934
rect 6892 29986 6948 29988
rect 6892 29934 6894 29986
rect 6894 29934 6946 29986
rect 6946 29934 6948 29986
rect 6892 29932 6948 29934
rect 7052 29986 7108 29988
rect 7052 29934 7054 29986
rect 7054 29934 7106 29986
rect 7106 29934 7108 29986
rect 7052 29932 7108 29934
rect 7212 29986 7268 29988
rect 7212 29934 7214 29986
rect 7214 29934 7266 29986
rect 7266 29934 7268 29986
rect 7212 29932 7268 29934
rect 7372 29986 7428 29988
rect 7372 29934 7374 29986
rect 7374 29934 7426 29986
rect 7426 29934 7428 29986
rect 7372 29932 7428 29934
rect 7532 29986 7588 29988
rect 7532 29934 7534 29986
rect 7534 29934 7586 29986
rect 7586 29934 7588 29986
rect 7532 29932 7588 29934
rect 7692 29986 7748 29988
rect 7692 29934 7694 29986
rect 7694 29934 7746 29986
rect 7746 29934 7748 29986
rect 7692 29932 7748 29934
rect 7852 29986 7908 29988
rect 7852 29934 7854 29986
rect 7854 29934 7906 29986
rect 7906 29934 7908 29986
rect 7852 29932 7908 29934
rect 8012 29986 8068 29988
rect 8012 29934 8014 29986
rect 8014 29934 8066 29986
rect 8066 29934 8068 29986
rect 8012 29932 8068 29934
rect 8172 29986 8228 29988
rect 8172 29934 8174 29986
rect 8174 29934 8226 29986
rect 8226 29934 8228 29986
rect 8172 29932 8228 29934
rect 8332 29986 8388 29988
rect 8332 29934 8334 29986
rect 8334 29934 8386 29986
rect 8386 29934 8388 29986
rect 8332 29932 8388 29934
rect 11532 29932 11588 29988
rect 11852 29932 11908 29988
rect 12492 29986 12548 29988
rect 12492 29934 12494 29986
rect 12494 29934 12546 29986
rect 12546 29934 12548 29986
rect 12492 29932 12548 29934
rect 12652 29986 12708 29988
rect 12652 29934 12654 29986
rect 12654 29934 12706 29986
rect 12706 29934 12708 29986
rect 12652 29932 12708 29934
rect 12812 29986 12868 29988
rect 12812 29934 12814 29986
rect 12814 29934 12866 29986
rect 12866 29934 12868 29986
rect 12812 29932 12868 29934
rect 12972 29986 13028 29988
rect 12972 29934 12974 29986
rect 12974 29934 13026 29986
rect 13026 29934 13028 29986
rect 12972 29932 13028 29934
rect 13132 29986 13188 29988
rect 13132 29934 13134 29986
rect 13134 29934 13186 29986
rect 13186 29934 13188 29986
rect 13132 29932 13188 29934
rect 13292 29986 13348 29988
rect 13292 29934 13294 29986
rect 13294 29934 13346 29986
rect 13346 29934 13348 29986
rect 13292 29932 13348 29934
rect 13452 29986 13508 29988
rect 13452 29934 13454 29986
rect 13454 29934 13506 29986
rect 13506 29934 13508 29986
rect 13452 29932 13508 29934
rect 13612 29986 13668 29988
rect 13612 29934 13614 29986
rect 13614 29934 13666 29986
rect 13666 29934 13668 29986
rect 13612 29932 13668 29934
rect 13772 29986 13828 29988
rect 13772 29934 13774 29986
rect 13774 29934 13826 29986
rect 13826 29934 13828 29986
rect 13772 29932 13828 29934
rect 13932 29986 13988 29988
rect 13932 29934 13934 29986
rect 13934 29934 13986 29986
rect 13986 29934 13988 29986
rect 13932 29932 13988 29934
rect 14092 29986 14148 29988
rect 14092 29934 14094 29986
rect 14094 29934 14146 29986
rect 14146 29934 14148 29986
rect 14092 29932 14148 29934
rect 14252 29986 14308 29988
rect 14252 29934 14254 29986
rect 14254 29934 14306 29986
rect 14306 29934 14308 29986
rect 14252 29932 14308 29934
rect 14412 29986 14468 29988
rect 14412 29934 14414 29986
rect 14414 29934 14466 29986
rect 14466 29934 14468 29986
rect 14412 29932 14468 29934
rect 14572 29986 14628 29988
rect 14572 29934 14574 29986
rect 14574 29934 14626 29986
rect 14626 29934 14628 29986
rect 14572 29932 14628 29934
rect 14732 29986 14788 29988
rect 14732 29934 14734 29986
rect 14734 29934 14786 29986
rect 14786 29934 14788 29986
rect 14732 29932 14788 29934
rect 14892 29986 14948 29988
rect 14892 29934 14894 29986
rect 14894 29934 14946 29986
rect 14946 29934 14948 29986
rect 14892 29932 14948 29934
rect 15052 29986 15108 29988
rect 15052 29934 15054 29986
rect 15054 29934 15106 29986
rect 15106 29934 15108 29986
rect 15052 29932 15108 29934
rect 15212 29986 15268 29988
rect 15212 29934 15214 29986
rect 15214 29934 15266 29986
rect 15266 29934 15268 29986
rect 15212 29932 15268 29934
rect 15372 29986 15428 29988
rect 15372 29934 15374 29986
rect 15374 29934 15426 29986
rect 15426 29934 15428 29986
rect 15372 29932 15428 29934
rect 15532 29986 15588 29988
rect 15532 29934 15534 29986
rect 15534 29934 15586 29986
rect 15586 29934 15588 29986
rect 15532 29932 15588 29934
rect 15692 29986 15748 29988
rect 15692 29934 15694 29986
rect 15694 29934 15746 29986
rect 15746 29934 15748 29986
rect 15692 29932 15748 29934
rect 15852 29986 15908 29988
rect 15852 29934 15854 29986
rect 15854 29934 15906 29986
rect 15906 29934 15908 29986
rect 15852 29932 15908 29934
rect 16012 29986 16068 29988
rect 16012 29934 16014 29986
rect 16014 29934 16066 29986
rect 16066 29934 16068 29986
rect 16012 29932 16068 29934
rect 16172 29986 16228 29988
rect 16172 29934 16174 29986
rect 16174 29934 16226 29986
rect 16226 29934 16228 29986
rect 16172 29932 16228 29934
rect 16332 29986 16388 29988
rect 16332 29934 16334 29986
rect 16334 29934 16386 29986
rect 16386 29934 16388 29986
rect 16332 29932 16388 29934
rect 16492 29986 16548 29988
rect 16492 29934 16494 29986
rect 16494 29934 16546 29986
rect 16546 29934 16548 29986
rect 16492 29932 16548 29934
rect 16652 29986 16708 29988
rect 16652 29934 16654 29986
rect 16654 29934 16706 29986
rect 16706 29934 16708 29986
rect 16652 29932 16708 29934
rect 16812 29986 16868 29988
rect 16812 29934 16814 29986
rect 16814 29934 16866 29986
rect 16866 29934 16868 29986
rect 16812 29932 16868 29934
rect 16972 29986 17028 29988
rect 16972 29934 16974 29986
rect 16974 29934 17026 29986
rect 17026 29934 17028 29986
rect 16972 29932 17028 29934
rect 17132 29986 17188 29988
rect 17132 29934 17134 29986
rect 17134 29934 17186 29986
rect 17186 29934 17188 29986
rect 17132 29932 17188 29934
rect 17292 29986 17348 29988
rect 17292 29934 17294 29986
rect 17294 29934 17346 29986
rect 17346 29934 17348 29986
rect 17292 29932 17348 29934
rect 17452 29986 17508 29988
rect 17452 29934 17454 29986
rect 17454 29934 17506 29986
rect 17506 29934 17508 29986
rect 17452 29932 17508 29934
rect 17612 29986 17668 29988
rect 17612 29934 17614 29986
rect 17614 29934 17666 29986
rect 17666 29934 17668 29986
rect 17612 29932 17668 29934
rect 17772 29986 17828 29988
rect 17772 29934 17774 29986
rect 17774 29934 17826 29986
rect 17826 29934 17828 29986
rect 17772 29932 17828 29934
rect 17932 29986 17988 29988
rect 17932 29934 17934 29986
rect 17934 29934 17986 29986
rect 17986 29934 17988 29986
rect 17932 29932 17988 29934
rect 18092 29986 18148 29988
rect 18092 29934 18094 29986
rect 18094 29934 18146 29986
rect 18146 29934 18148 29986
rect 18092 29932 18148 29934
rect 18252 29986 18308 29988
rect 18252 29934 18254 29986
rect 18254 29934 18306 29986
rect 18306 29934 18308 29986
rect 18252 29932 18308 29934
rect 18412 29986 18468 29988
rect 18412 29934 18414 29986
rect 18414 29934 18466 29986
rect 18466 29934 18468 29986
rect 18412 29932 18468 29934
rect 18572 29986 18628 29988
rect 18572 29934 18574 29986
rect 18574 29934 18626 29986
rect 18626 29934 18628 29986
rect 18572 29932 18628 29934
rect 18732 29986 18788 29988
rect 18732 29934 18734 29986
rect 18734 29934 18786 29986
rect 18786 29934 18788 29986
rect 18732 29932 18788 29934
rect 18892 29986 18948 29988
rect 18892 29934 18894 29986
rect 18894 29934 18946 29986
rect 18946 29934 18948 29986
rect 18892 29932 18948 29934
rect 22092 29932 22148 29988
rect 22412 29932 22468 29988
rect 23132 29986 23188 29988
rect 23132 29934 23134 29986
rect 23134 29934 23186 29986
rect 23186 29934 23188 29986
rect 23132 29932 23188 29934
rect 23292 29986 23348 29988
rect 23292 29934 23294 29986
rect 23294 29934 23346 29986
rect 23346 29934 23348 29986
rect 23292 29932 23348 29934
rect 23452 29986 23508 29988
rect 23452 29934 23454 29986
rect 23454 29934 23506 29986
rect 23506 29934 23508 29986
rect 23452 29932 23508 29934
rect 23612 29986 23668 29988
rect 23612 29934 23614 29986
rect 23614 29934 23666 29986
rect 23666 29934 23668 29986
rect 23612 29932 23668 29934
rect 23772 29986 23828 29988
rect 23772 29934 23774 29986
rect 23774 29934 23826 29986
rect 23826 29934 23828 29986
rect 23772 29932 23828 29934
rect 23932 29986 23988 29988
rect 23932 29934 23934 29986
rect 23934 29934 23986 29986
rect 23986 29934 23988 29986
rect 23932 29932 23988 29934
rect 24092 29986 24148 29988
rect 24092 29934 24094 29986
rect 24094 29934 24146 29986
rect 24146 29934 24148 29986
rect 24092 29932 24148 29934
rect 24252 29986 24308 29988
rect 24252 29934 24254 29986
rect 24254 29934 24306 29986
rect 24306 29934 24308 29986
rect 24252 29932 24308 29934
rect 24412 29986 24468 29988
rect 24412 29934 24414 29986
rect 24414 29934 24466 29986
rect 24466 29934 24468 29986
rect 24412 29932 24468 29934
rect 24572 29986 24628 29988
rect 24572 29934 24574 29986
rect 24574 29934 24626 29986
rect 24626 29934 24628 29986
rect 24572 29932 24628 29934
rect 24732 29986 24788 29988
rect 24732 29934 24734 29986
rect 24734 29934 24786 29986
rect 24786 29934 24788 29986
rect 24732 29932 24788 29934
rect 24892 29986 24948 29988
rect 24892 29934 24894 29986
rect 24894 29934 24946 29986
rect 24946 29934 24948 29986
rect 24892 29932 24948 29934
rect 25052 29986 25108 29988
rect 25052 29934 25054 29986
rect 25054 29934 25106 29986
rect 25106 29934 25108 29986
rect 25052 29932 25108 29934
rect 25212 29986 25268 29988
rect 25212 29934 25214 29986
rect 25214 29934 25266 29986
rect 25266 29934 25268 29986
rect 25212 29932 25268 29934
rect 25372 29986 25428 29988
rect 25372 29934 25374 29986
rect 25374 29934 25426 29986
rect 25426 29934 25428 29986
rect 25372 29932 25428 29934
rect 25532 29986 25588 29988
rect 25532 29934 25534 29986
rect 25534 29934 25586 29986
rect 25586 29934 25588 29986
rect 25532 29932 25588 29934
rect 25692 29986 25748 29988
rect 25692 29934 25694 29986
rect 25694 29934 25746 29986
rect 25746 29934 25748 29986
rect 25692 29932 25748 29934
rect 25852 29986 25908 29988
rect 25852 29934 25854 29986
rect 25854 29934 25906 29986
rect 25906 29934 25908 29986
rect 25852 29932 25908 29934
rect 26012 29986 26068 29988
rect 26012 29934 26014 29986
rect 26014 29934 26066 29986
rect 26066 29934 26068 29986
rect 26012 29932 26068 29934
rect 26172 29986 26228 29988
rect 26172 29934 26174 29986
rect 26174 29934 26226 29986
rect 26226 29934 26228 29986
rect 26172 29932 26228 29934
rect 26332 29986 26388 29988
rect 26332 29934 26334 29986
rect 26334 29934 26386 29986
rect 26386 29934 26388 29986
rect 26332 29932 26388 29934
rect 26492 29986 26548 29988
rect 26492 29934 26494 29986
rect 26494 29934 26546 29986
rect 26546 29934 26548 29986
rect 26492 29932 26548 29934
rect 26652 29986 26708 29988
rect 26652 29934 26654 29986
rect 26654 29934 26706 29986
rect 26706 29934 26708 29986
rect 26652 29932 26708 29934
rect 26812 29986 26868 29988
rect 26812 29934 26814 29986
rect 26814 29934 26866 29986
rect 26866 29934 26868 29986
rect 26812 29932 26868 29934
rect 26972 29986 27028 29988
rect 26972 29934 26974 29986
rect 26974 29934 27026 29986
rect 27026 29934 27028 29986
rect 26972 29932 27028 29934
rect 27132 29986 27188 29988
rect 27132 29934 27134 29986
rect 27134 29934 27186 29986
rect 27186 29934 27188 29986
rect 27132 29932 27188 29934
rect 27292 29986 27348 29988
rect 27292 29934 27294 29986
rect 27294 29934 27346 29986
rect 27346 29934 27348 29986
rect 27292 29932 27348 29934
rect 27452 29986 27508 29988
rect 27452 29934 27454 29986
rect 27454 29934 27506 29986
rect 27506 29934 27508 29986
rect 27452 29932 27508 29934
rect 27612 29986 27668 29988
rect 27612 29934 27614 29986
rect 27614 29934 27666 29986
rect 27666 29934 27668 29986
rect 27612 29932 27668 29934
rect 27772 29986 27828 29988
rect 27772 29934 27774 29986
rect 27774 29934 27826 29986
rect 27826 29934 27828 29986
rect 27772 29932 27828 29934
rect 27932 29986 27988 29988
rect 27932 29934 27934 29986
rect 27934 29934 27986 29986
rect 27986 29934 27988 29986
rect 27932 29932 27988 29934
rect 28092 29986 28148 29988
rect 28092 29934 28094 29986
rect 28094 29934 28146 29986
rect 28146 29934 28148 29986
rect 28092 29932 28148 29934
rect 28252 29986 28308 29988
rect 28252 29934 28254 29986
rect 28254 29934 28306 29986
rect 28306 29934 28308 29986
rect 28252 29932 28308 29934
rect 28412 29986 28468 29988
rect 28412 29934 28414 29986
rect 28414 29934 28466 29986
rect 28466 29934 28468 29986
rect 28412 29932 28468 29934
rect 28572 29986 28628 29988
rect 28572 29934 28574 29986
rect 28574 29934 28626 29986
rect 28626 29934 28628 29986
rect 28572 29932 28628 29934
rect 28732 29986 28788 29988
rect 28732 29934 28734 29986
rect 28734 29934 28786 29986
rect 28786 29934 28788 29986
rect 28732 29932 28788 29934
rect 28892 29986 28948 29988
rect 28892 29934 28894 29986
rect 28894 29934 28946 29986
rect 28946 29934 28948 29986
rect 28892 29932 28948 29934
rect 29052 29986 29108 29988
rect 29052 29934 29054 29986
rect 29054 29934 29106 29986
rect 29106 29934 29108 29986
rect 29052 29932 29108 29934
rect 29212 29986 29268 29988
rect 29212 29934 29214 29986
rect 29214 29934 29266 29986
rect 29266 29934 29268 29986
rect 29212 29932 29268 29934
rect 29372 29986 29428 29988
rect 29372 29934 29374 29986
rect 29374 29934 29426 29986
rect 29426 29934 29428 29986
rect 29372 29932 29428 29934
rect 30012 29932 30068 29988
rect 30332 29932 30388 29988
rect 33532 29986 33588 29988
rect 33532 29934 33534 29986
rect 33534 29934 33586 29986
rect 33586 29934 33588 29986
rect 33532 29932 33588 29934
rect 33692 29986 33748 29988
rect 33692 29934 33694 29986
rect 33694 29934 33746 29986
rect 33746 29934 33748 29986
rect 33692 29932 33748 29934
rect 33852 29986 33908 29988
rect 33852 29934 33854 29986
rect 33854 29934 33906 29986
rect 33906 29934 33908 29986
rect 33852 29932 33908 29934
rect 34012 29986 34068 29988
rect 34012 29934 34014 29986
rect 34014 29934 34066 29986
rect 34066 29934 34068 29986
rect 34012 29932 34068 29934
rect 34172 29986 34228 29988
rect 34172 29934 34174 29986
rect 34174 29934 34226 29986
rect 34226 29934 34228 29986
rect 34172 29932 34228 29934
rect 34332 29986 34388 29988
rect 34332 29934 34334 29986
rect 34334 29934 34386 29986
rect 34386 29934 34388 29986
rect 34332 29932 34388 29934
rect 34492 29986 34548 29988
rect 34492 29934 34494 29986
rect 34494 29934 34546 29986
rect 34546 29934 34548 29986
rect 34492 29932 34548 29934
rect 34652 29986 34708 29988
rect 34652 29934 34654 29986
rect 34654 29934 34706 29986
rect 34706 29934 34708 29986
rect 34652 29932 34708 29934
rect 34812 29986 34868 29988
rect 34812 29934 34814 29986
rect 34814 29934 34866 29986
rect 34866 29934 34868 29986
rect 34812 29932 34868 29934
rect 34972 29986 35028 29988
rect 34972 29934 34974 29986
rect 34974 29934 35026 29986
rect 35026 29934 35028 29986
rect 34972 29932 35028 29934
rect 35132 29986 35188 29988
rect 35132 29934 35134 29986
rect 35134 29934 35186 29986
rect 35186 29934 35188 29986
rect 35132 29932 35188 29934
rect 35292 29986 35348 29988
rect 35292 29934 35294 29986
rect 35294 29934 35346 29986
rect 35346 29934 35348 29986
rect 35292 29932 35348 29934
rect 35452 29986 35508 29988
rect 35452 29934 35454 29986
rect 35454 29934 35506 29986
rect 35506 29934 35508 29986
rect 35452 29932 35508 29934
rect 35612 29986 35668 29988
rect 35612 29934 35614 29986
rect 35614 29934 35666 29986
rect 35666 29934 35668 29986
rect 35612 29932 35668 29934
rect 35772 29986 35828 29988
rect 35772 29934 35774 29986
rect 35774 29934 35826 29986
rect 35826 29934 35828 29986
rect 35772 29932 35828 29934
rect 35932 29986 35988 29988
rect 35932 29934 35934 29986
rect 35934 29934 35986 29986
rect 35986 29934 35988 29986
rect 35932 29932 35988 29934
rect 36092 29986 36148 29988
rect 36092 29934 36094 29986
rect 36094 29934 36146 29986
rect 36146 29934 36148 29986
rect 36092 29932 36148 29934
rect 36252 29986 36308 29988
rect 36252 29934 36254 29986
rect 36254 29934 36306 29986
rect 36306 29934 36308 29986
rect 36252 29932 36308 29934
rect 36412 29986 36468 29988
rect 36412 29934 36414 29986
rect 36414 29934 36466 29986
rect 36466 29934 36468 29986
rect 36412 29932 36468 29934
rect 36572 29986 36628 29988
rect 36572 29934 36574 29986
rect 36574 29934 36626 29986
rect 36626 29934 36628 29986
rect 36572 29932 36628 29934
rect 36732 29986 36788 29988
rect 36732 29934 36734 29986
rect 36734 29934 36786 29986
rect 36786 29934 36788 29986
rect 36732 29932 36788 29934
rect 36892 29986 36948 29988
rect 36892 29934 36894 29986
rect 36894 29934 36946 29986
rect 36946 29934 36948 29986
rect 36892 29932 36948 29934
rect 37052 29986 37108 29988
rect 37052 29934 37054 29986
rect 37054 29934 37106 29986
rect 37106 29934 37108 29986
rect 37052 29932 37108 29934
rect 37212 29986 37268 29988
rect 37212 29934 37214 29986
rect 37214 29934 37266 29986
rect 37266 29934 37268 29986
rect 37212 29932 37268 29934
rect 37372 29986 37428 29988
rect 37372 29934 37374 29986
rect 37374 29934 37426 29986
rect 37426 29934 37428 29986
rect 37372 29932 37428 29934
rect 37532 29986 37588 29988
rect 37532 29934 37534 29986
rect 37534 29934 37586 29986
rect 37586 29934 37588 29986
rect 37532 29932 37588 29934
rect 37692 29986 37748 29988
rect 37692 29934 37694 29986
rect 37694 29934 37746 29986
rect 37746 29934 37748 29986
rect 37692 29932 37748 29934
rect 37852 29986 37908 29988
rect 37852 29934 37854 29986
rect 37854 29934 37906 29986
rect 37906 29934 37908 29986
rect 37852 29932 37908 29934
rect 38012 29986 38068 29988
rect 38012 29934 38014 29986
rect 38014 29934 38066 29986
rect 38066 29934 38068 29986
rect 38012 29932 38068 29934
rect 38172 29986 38228 29988
rect 38172 29934 38174 29986
rect 38174 29934 38226 29986
rect 38226 29934 38228 29986
rect 38172 29932 38228 29934
rect 38332 29986 38388 29988
rect 38332 29934 38334 29986
rect 38334 29934 38386 29986
rect 38386 29934 38388 29986
rect 38332 29932 38388 29934
rect 38492 29986 38548 29988
rect 38492 29934 38494 29986
rect 38494 29934 38546 29986
rect 38546 29934 38548 29986
rect 38492 29932 38548 29934
rect 38652 29986 38708 29988
rect 38652 29934 38654 29986
rect 38654 29934 38706 29986
rect 38706 29934 38708 29986
rect 38652 29932 38708 29934
rect 38812 29986 38868 29988
rect 38812 29934 38814 29986
rect 38814 29934 38866 29986
rect 38866 29934 38868 29986
rect 38812 29932 38868 29934
rect 38972 29986 39028 29988
rect 38972 29934 38974 29986
rect 38974 29934 39026 29986
rect 39026 29934 39028 29986
rect 38972 29932 39028 29934
rect 39132 29986 39188 29988
rect 39132 29934 39134 29986
rect 39134 29934 39186 29986
rect 39186 29934 39188 29986
rect 39132 29932 39188 29934
rect 39292 29986 39348 29988
rect 39292 29934 39294 29986
rect 39294 29934 39346 29986
rect 39346 29934 39348 29986
rect 39292 29932 39348 29934
rect 39452 29986 39508 29988
rect 39452 29934 39454 29986
rect 39454 29934 39506 29986
rect 39506 29934 39508 29986
rect 39452 29932 39508 29934
rect 39612 29986 39668 29988
rect 39612 29934 39614 29986
rect 39614 29934 39666 29986
rect 39666 29934 39668 29986
rect 39612 29932 39668 29934
rect 39772 29986 39828 29988
rect 39772 29934 39774 29986
rect 39774 29934 39826 29986
rect 39826 29934 39828 29986
rect 39772 29932 39828 29934
rect 39932 29986 39988 29988
rect 39932 29934 39934 29986
rect 39934 29934 39986 29986
rect 39986 29934 39988 29986
rect 39932 29932 39988 29934
rect 40092 29986 40148 29988
rect 40092 29934 40094 29986
rect 40094 29934 40146 29986
rect 40146 29934 40148 29986
rect 40092 29932 40148 29934
rect 40252 29986 40308 29988
rect 40252 29934 40254 29986
rect 40254 29934 40306 29986
rect 40306 29934 40308 29986
rect 40252 29932 40308 29934
rect 40412 29986 40468 29988
rect 40412 29934 40414 29986
rect 40414 29934 40466 29986
rect 40466 29934 40468 29986
rect 40412 29932 40468 29934
rect 40572 29986 40628 29988
rect 40572 29934 40574 29986
rect 40574 29934 40626 29986
rect 40626 29934 40628 29986
rect 40572 29932 40628 29934
rect 40732 29986 40788 29988
rect 40732 29934 40734 29986
rect 40734 29934 40786 29986
rect 40786 29934 40788 29986
rect 40732 29932 40788 29934
rect 40892 29986 40948 29988
rect 40892 29934 40894 29986
rect 40894 29934 40946 29986
rect 40946 29934 40948 29986
rect 40892 29932 40948 29934
rect 41052 29986 41108 29988
rect 41052 29934 41054 29986
rect 41054 29934 41106 29986
rect 41106 29934 41108 29986
rect 41052 29932 41108 29934
rect 41212 29986 41268 29988
rect 41212 29934 41214 29986
rect 41214 29934 41266 29986
rect 41266 29934 41268 29986
rect 41212 29932 41268 29934
rect 41372 29986 41428 29988
rect 41372 29934 41374 29986
rect 41374 29934 41426 29986
rect 41426 29934 41428 29986
rect 41372 29932 41428 29934
rect 41532 29986 41588 29988
rect 41532 29934 41534 29986
rect 41534 29934 41586 29986
rect 41586 29934 41588 29986
rect 41532 29932 41588 29934
rect 41692 29986 41748 29988
rect 41692 29934 41694 29986
rect 41694 29934 41746 29986
rect 41746 29934 41748 29986
rect 41692 29932 41748 29934
rect 41852 29986 41908 29988
rect 41852 29934 41854 29986
rect 41854 29934 41906 29986
rect 41906 29934 41908 29986
rect 41852 29932 41908 29934
rect 12 29826 68 29828
rect 12 29774 14 29826
rect 14 29774 66 29826
rect 66 29774 68 29826
rect 12 29772 68 29774
rect 172 29826 228 29828
rect 172 29774 174 29826
rect 174 29774 226 29826
rect 226 29774 228 29826
rect 172 29772 228 29774
rect 332 29826 388 29828
rect 332 29774 334 29826
rect 334 29774 386 29826
rect 386 29774 388 29826
rect 332 29772 388 29774
rect 492 29826 548 29828
rect 492 29774 494 29826
rect 494 29774 546 29826
rect 546 29774 548 29826
rect 492 29772 548 29774
rect 652 29826 708 29828
rect 652 29774 654 29826
rect 654 29774 706 29826
rect 706 29774 708 29826
rect 652 29772 708 29774
rect 812 29826 868 29828
rect 812 29774 814 29826
rect 814 29774 866 29826
rect 866 29774 868 29826
rect 812 29772 868 29774
rect 972 29826 1028 29828
rect 972 29774 974 29826
rect 974 29774 1026 29826
rect 1026 29774 1028 29826
rect 972 29772 1028 29774
rect 1132 29826 1188 29828
rect 1132 29774 1134 29826
rect 1134 29774 1186 29826
rect 1186 29774 1188 29826
rect 1132 29772 1188 29774
rect 1292 29826 1348 29828
rect 1292 29774 1294 29826
rect 1294 29774 1346 29826
rect 1346 29774 1348 29826
rect 1292 29772 1348 29774
rect 1452 29826 1508 29828
rect 1452 29774 1454 29826
rect 1454 29774 1506 29826
rect 1506 29774 1508 29826
rect 1452 29772 1508 29774
rect 1612 29826 1668 29828
rect 1612 29774 1614 29826
rect 1614 29774 1666 29826
rect 1666 29774 1668 29826
rect 1612 29772 1668 29774
rect 1772 29826 1828 29828
rect 1772 29774 1774 29826
rect 1774 29774 1826 29826
rect 1826 29774 1828 29826
rect 1772 29772 1828 29774
rect 1932 29826 1988 29828
rect 1932 29774 1934 29826
rect 1934 29774 1986 29826
rect 1986 29774 1988 29826
rect 1932 29772 1988 29774
rect 2092 29826 2148 29828
rect 2092 29774 2094 29826
rect 2094 29774 2146 29826
rect 2146 29774 2148 29826
rect 2092 29772 2148 29774
rect 2252 29826 2308 29828
rect 2252 29774 2254 29826
rect 2254 29774 2306 29826
rect 2306 29774 2308 29826
rect 2252 29772 2308 29774
rect 2412 29826 2468 29828
rect 2412 29774 2414 29826
rect 2414 29774 2466 29826
rect 2466 29774 2468 29826
rect 2412 29772 2468 29774
rect 2572 29826 2628 29828
rect 2572 29774 2574 29826
rect 2574 29774 2626 29826
rect 2626 29774 2628 29826
rect 2572 29772 2628 29774
rect 2732 29826 2788 29828
rect 2732 29774 2734 29826
rect 2734 29774 2786 29826
rect 2786 29774 2788 29826
rect 2732 29772 2788 29774
rect 2892 29826 2948 29828
rect 2892 29774 2894 29826
rect 2894 29774 2946 29826
rect 2946 29774 2948 29826
rect 2892 29772 2948 29774
rect 3052 29826 3108 29828
rect 3052 29774 3054 29826
rect 3054 29774 3106 29826
rect 3106 29774 3108 29826
rect 3052 29772 3108 29774
rect 3212 29826 3268 29828
rect 3212 29774 3214 29826
rect 3214 29774 3266 29826
rect 3266 29774 3268 29826
rect 3212 29772 3268 29774
rect 3372 29826 3428 29828
rect 3372 29774 3374 29826
rect 3374 29774 3426 29826
rect 3426 29774 3428 29826
rect 3372 29772 3428 29774
rect 3532 29826 3588 29828
rect 3532 29774 3534 29826
rect 3534 29774 3586 29826
rect 3586 29774 3588 29826
rect 3532 29772 3588 29774
rect 3692 29826 3748 29828
rect 3692 29774 3694 29826
rect 3694 29774 3746 29826
rect 3746 29774 3748 29826
rect 3692 29772 3748 29774
rect 3852 29826 3908 29828
rect 3852 29774 3854 29826
rect 3854 29774 3906 29826
rect 3906 29774 3908 29826
rect 3852 29772 3908 29774
rect 4012 29826 4068 29828
rect 4012 29774 4014 29826
rect 4014 29774 4066 29826
rect 4066 29774 4068 29826
rect 4012 29772 4068 29774
rect 4172 29826 4228 29828
rect 4172 29774 4174 29826
rect 4174 29774 4226 29826
rect 4226 29774 4228 29826
rect 4172 29772 4228 29774
rect 4332 29826 4388 29828
rect 4332 29774 4334 29826
rect 4334 29774 4386 29826
rect 4386 29774 4388 29826
rect 4332 29772 4388 29774
rect 4492 29826 4548 29828
rect 4492 29774 4494 29826
rect 4494 29774 4546 29826
rect 4546 29774 4548 29826
rect 4492 29772 4548 29774
rect 4652 29826 4708 29828
rect 4652 29774 4654 29826
rect 4654 29774 4706 29826
rect 4706 29774 4708 29826
rect 4652 29772 4708 29774
rect 4812 29826 4868 29828
rect 4812 29774 4814 29826
rect 4814 29774 4866 29826
rect 4866 29774 4868 29826
rect 4812 29772 4868 29774
rect 4972 29826 5028 29828
rect 4972 29774 4974 29826
rect 4974 29774 5026 29826
rect 5026 29774 5028 29826
rect 4972 29772 5028 29774
rect 5132 29826 5188 29828
rect 5132 29774 5134 29826
rect 5134 29774 5186 29826
rect 5186 29774 5188 29826
rect 5132 29772 5188 29774
rect 5292 29826 5348 29828
rect 5292 29774 5294 29826
rect 5294 29774 5346 29826
rect 5346 29774 5348 29826
rect 5292 29772 5348 29774
rect 5452 29826 5508 29828
rect 5452 29774 5454 29826
rect 5454 29774 5506 29826
rect 5506 29774 5508 29826
rect 5452 29772 5508 29774
rect 5612 29826 5668 29828
rect 5612 29774 5614 29826
rect 5614 29774 5666 29826
rect 5666 29774 5668 29826
rect 5612 29772 5668 29774
rect 5772 29826 5828 29828
rect 5772 29774 5774 29826
rect 5774 29774 5826 29826
rect 5826 29774 5828 29826
rect 5772 29772 5828 29774
rect 5932 29826 5988 29828
rect 5932 29774 5934 29826
rect 5934 29774 5986 29826
rect 5986 29774 5988 29826
rect 5932 29772 5988 29774
rect 6092 29826 6148 29828
rect 6092 29774 6094 29826
rect 6094 29774 6146 29826
rect 6146 29774 6148 29826
rect 6092 29772 6148 29774
rect 6252 29826 6308 29828
rect 6252 29774 6254 29826
rect 6254 29774 6306 29826
rect 6306 29774 6308 29826
rect 6252 29772 6308 29774
rect 6412 29826 6468 29828
rect 6412 29774 6414 29826
rect 6414 29774 6466 29826
rect 6466 29774 6468 29826
rect 6412 29772 6468 29774
rect 6572 29826 6628 29828
rect 6572 29774 6574 29826
rect 6574 29774 6626 29826
rect 6626 29774 6628 29826
rect 6572 29772 6628 29774
rect 6732 29826 6788 29828
rect 6732 29774 6734 29826
rect 6734 29774 6786 29826
rect 6786 29774 6788 29826
rect 6732 29772 6788 29774
rect 6892 29826 6948 29828
rect 6892 29774 6894 29826
rect 6894 29774 6946 29826
rect 6946 29774 6948 29826
rect 6892 29772 6948 29774
rect 7052 29826 7108 29828
rect 7052 29774 7054 29826
rect 7054 29774 7106 29826
rect 7106 29774 7108 29826
rect 7052 29772 7108 29774
rect 7212 29826 7268 29828
rect 7212 29774 7214 29826
rect 7214 29774 7266 29826
rect 7266 29774 7268 29826
rect 7212 29772 7268 29774
rect 7372 29826 7428 29828
rect 7372 29774 7374 29826
rect 7374 29774 7426 29826
rect 7426 29774 7428 29826
rect 7372 29772 7428 29774
rect 7532 29826 7588 29828
rect 7532 29774 7534 29826
rect 7534 29774 7586 29826
rect 7586 29774 7588 29826
rect 7532 29772 7588 29774
rect 7692 29826 7748 29828
rect 7692 29774 7694 29826
rect 7694 29774 7746 29826
rect 7746 29774 7748 29826
rect 7692 29772 7748 29774
rect 7852 29826 7908 29828
rect 7852 29774 7854 29826
rect 7854 29774 7906 29826
rect 7906 29774 7908 29826
rect 7852 29772 7908 29774
rect 8012 29826 8068 29828
rect 8012 29774 8014 29826
rect 8014 29774 8066 29826
rect 8066 29774 8068 29826
rect 8012 29772 8068 29774
rect 8172 29826 8228 29828
rect 8172 29774 8174 29826
rect 8174 29774 8226 29826
rect 8226 29774 8228 29826
rect 8172 29772 8228 29774
rect 8332 29826 8388 29828
rect 8332 29774 8334 29826
rect 8334 29774 8386 29826
rect 8386 29774 8388 29826
rect 8332 29772 8388 29774
rect 12012 29772 12068 29828
rect 12332 29772 12388 29828
rect 12492 29826 12548 29828
rect 12492 29774 12494 29826
rect 12494 29774 12546 29826
rect 12546 29774 12548 29826
rect 12492 29772 12548 29774
rect 12652 29826 12708 29828
rect 12652 29774 12654 29826
rect 12654 29774 12706 29826
rect 12706 29774 12708 29826
rect 12652 29772 12708 29774
rect 12812 29826 12868 29828
rect 12812 29774 12814 29826
rect 12814 29774 12866 29826
rect 12866 29774 12868 29826
rect 12812 29772 12868 29774
rect 12972 29826 13028 29828
rect 12972 29774 12974 29826
rect 12974 29774 13026 29826
rect 13026 29774 13028 29826
rect 12972 29772 13028 29774
rect 13132 29826 13188 29828
rect 13132 29774 13134 29826
rect 13134 29774 13186 29826
rect 13186 29774 13188 29826
rect 13132 29772 13188 29774
rect 13292 29826 13348 29828
rect 13292 29774 13294 29826
rect 13294 29774 13346 29826
rect 13346 29774 13348 29826
rect 13292 29772 13348 29774
rect 13452 29826 13508 29828
rect 13452 29774 13454 29826
rect 13454 29774 13506 29826
rect 13506 29774 13508 29826
rect 13452 29772 13508 29774
rect 13612 29826 13668 29828
rect 13612 29774 13614 29826
rect 13614 29774 13666 29826
rect 13666 29774 13668 29826
rect 13612 29772 13668 29774
rect 13772 29826 13828 29828
rect 13772 29774 13774 29826
rect 13774 29774 13826 29826
rect 13826 29774 13828 29826
rect 13772 29772 13828 29774
rect 13932 29826 13988 29828
rect 13932 29774 13934 29826
rect 13934 29774 13986 29826
rect 13986 29774 13988 29826
rect 13932 29772 13988 29774
rect 14092 29826 14148 29828
rect 14092 29774 14094 29826
rect 14094 29774 14146 29826
rect 14146 29774 14148 29826
rect 14092 29772 14148 29774
rect 14252 29826 14308 29828
rect 14252 29774 14254 29826
rect 14254 29774 14306 29826
rect 14306 29774 14308 29826
rect 14252 29772 14308 29774
rect 14412 29826 14468 29828
rect 14412 29774 14414 29826
rect 14414 29774 14466 29826
rect 14466 29774 14468 29826
rect 14412 29772 14468 29774
rect 14572 29826 14628 29828
rect 14572 29774 14574 29826
rect 14574 29774 14626 29826
rect 14626 29774 14628 29826
rect 14572 29772 14628 29774
rect 14732 29826 14788 29828
rect 14732 29774 14734 29826
rect 14734 29774 14786 29826
rect 14786 29774 14788 29826
rect 14732 29772 14788 29774
rect 14892 29826 14948 29828
rect 14892 29774 14894 29826
rect 14894 29774 14946 29826
rect 14946 29774 14948 29826
rect 14892 29772 14948 29774
rect 15052 29826 15108 29828
rect 15052 29774 15054 29826
rect 15054 29774 15106 29826
rect 15106 29774 15108 29826
rect 15052 29772 15108 29774
rect 15212 29826 15268 29828
rect 15212 29774 15214 29826
rect 15214 29774 15266 29826
rect 15266 29774 15268 29826
rect 15212 29772 15268 29774
rect 15372 29826 15428 29828
rect 15372 29774 15374 29826
rect 15374 29774 15426 29826
rect 15426 29774 15428 29826
rect 15372 29772 15428 29774
rect 15532 29826 15588 29828
rect 15532 29774 15534 29826
rect 15534 29774 15586 29826
rect 15586 29774 15588 29826
rect 15532 29772 15588 29774
rect 15692 29826 15748 29828
rect 15692 29774 15694 29826
rect 15694 29774 15746 29826
rect 15746 29774 15748 29826
rect 15692 29772 15748 29774
rect 15852 29826 15908 29828
rect 15852 29774 15854 29826
rect 15854 29774 15906 29826
rect 15906 29774 15908 29826
rect 15852 29772 15908 29774
rect 16012 29826 16068 29828
rect 16012 29774 16014 29826
rect 16014 29774 16066 29826
rect 16066 29774 16068 29826
rect 16012 29772 16068 29774
rect 16172 29826 16228 29828
rect 16172 29774 16174 29826
rect 16174 29774 16226 29826
rect 16226 29774 16228 29826
rect 16172 29772 16228 29774
rect 16332 29826 16388 29828
rect 16332 29774 16334 29826
rect 16334 29774 16386 29826
rect 16386 29774 16388 29826
rect 16332 29772 16388 29774
rect 16492 29826 16548 29828
rect 16492 29774 16494 29826
rect 16494 29774 16546 29826
rect 16546 29774 16548 29826
rect 16492 29772 16548 29774
rect 16652 29826 16708 29828
rect 16652 29774 16654 29826
rect 16654 29774 16706 29826
rect 16706 29774 16708 29826
rect 16652 29772 16708 29774
rect 16812 29826 16868 29828
rect 16812 29774 16814 29826
rect 16814 29774 16866 29826
rect 16866 29774 16868 29826
rect 16812 29772 16868 29774
rect 16972 29826 17028 29828
rect 16972 29774 16974 29826
rect 16974 29774 17026 29826
rect 17026 29774 17028 29826
rect 16972 29772 17028 29774
rect 17132 29826 17188 29828
rect 17132 29774 17134 29826
rect 17134 29774 17186 29826
rect 17186 29774 17188 29826
rect 17132 29772 17188 29774
rect 17292 29826 17348 29828
rect 17292 29774 17294 29826
rect 17294 29774 17346 29826
rect 17346 29774 17348 29826
rect 17292 29772 17348 29774
rect 17452 29826 17508 29828
rect 17452 29774 17454 29826
rect 17454 29774 17506 29826
rect 17506 29774 17508 29826
rect 17452 29772 17508 29774
rect 17612 29826 17668 29828
rect 17612 29774 17614 29826
rect 17614 29774 17666 29826
rect 17666 29774 17668 29826
rect 17612 29772 17668 29774
rect 17772 29826 17828 29828
rect 17772 29774 17774 29826
rect 17774 29774 17826 29826
rect 17826 29774 17828 29826
rect 17772 29772 17828 29774
rect 17932 29826 17988 29828
rect 17932 29774 17934 29826
rect 17934 29774 17986 29826
rect 17986 29774 17988 29826
rect 17932 29772 17988 29774
rect 18092 29826 18148 29828
rect 18092 29774 18094 29826
rect 18094 29774 18146 29826
rect 18146 29774 18148 29826
rect 18092 29772 18148 29774
rect 18252 29826 18308 29828
rect 18252 29774 18254 29826
rect 18254 29774 18306 29826
rect 18306 29774 18308 29826
rect 18252 29772 18308 29774
rect 18412 29826 18468 29828
rect 18412 29774 18414 29826
rect 18414 29774 18466 29826
rect 18466 29774 18468 29826
rect 18412 29772 18468 29774
rect 18572 29826 18628 29828
rect 18572 29774 18574 29826
rect 18574 29774 18626 29826
rect 18626 29774 18628 29826
rect 18572 29772 18628 29774
rect 18732 29826 18788 29828
rect 18732 29774 18734 29826
rect 18734 29774 18786 29826
rect 18786 29774 18788 29826
rect 18732 29772 18788 29774
rect 18892 29826 18948 29828
rect 18892 29774 18894 29826
rect 18894 29774 18946 29826
rect 18946 29774 18948 29826
rect 18892 29772 18948 29774
rect 22572 29772 22628 29828
rect 22892 29772 22948 29828
rect 23132 29826 23188 29828
rect 23132 29774 23134 29826
rect 23134 29774 23186 29826
rect 23186 29774 23188 29826
rect 23132 29772 23188 29774
rect 23292 29826 23348 29828
rect 23292 29774 23294 29826
rect 23294 29774 23346 29826
rect 23346 29774 23348 29826
rect 23292 29772 23348 29774
rect 23452 29826 23508 29828
rect 23452 29774 23454 29826
rect 23454 29774 23506 29826
rect 23506 29774 23508 29826
rect 23452 29772 23508 29774
rect 23612 29826 23668 29828
rect 23612 29774 23614 29826
rect 23614 29774 23666 29826
rect 23666 29774 23668 29826
rect 23612 29772 23668 29774
rect 23772 29826 23828 29828
rect 23772 29774 23774 29826
rect 23774 29774 23826 29826
rect 23826 29774 23828 29826
rect 23772 29772 23828 29774
rect 23932 29826 23988 29828
rect 23932 29774 23934 29826
rect 23934 29774 23986 29826
rect 23986 29774 23988 29826
rect 23932 29772 23988 29774
rect 24092 29826 24148 29828
rect 24092 29774 24094 29826
rect 24094 29774 24146 29826
rect 24146 29774 24148 29826
rect 24092 29772 24148 29774
rect 24252 29826 24308 29828
rect 24252 29774 24254 29826
rect 24254 29774 24306 29826
rect 24306 29774 24308 29826
rect 24252 29772 24308 29774
rect 24412 29826 24468 29828
rect 24412 29774 24414 29826
rect 24414 29774 24466 29826
rect 24466 29774 24468 29826
rect 24412 29772 24468 29774
rect 24572 29826 24628 29828
rect 24572 29774 24574 29826
rect 24574 29774 24626 29826
rect 24626 29774 24628 29826
rect 24572 29772 24628 29774
rect 24732 29826 24788 29828
rect 24732 29774 24734 29826
rect 24734 29774 24786 29826
rect 24786 29774 24788 29826
rect 24732 29772 24788 29774
rect 24892 29826 24948 29828
rect 24892 29774 24894 29826
rect 24894 29774 24946 29826
rect 24946 29774 24948 29826
rect 24892 29772 24948 29774
rect 25052 29826 25108 29828
rect 25052 29774 25054 29826
rect 25054 29774 25106 29826
rect 25106 29774 25108 29826
rect 25052 29772 25108 29774
rect 25212 29826 25268 29828
rect 25212 29774 25214 29826
rect 25214 29774 25266 29826
rect 25266 29774 25268 29826
rect 25212 29772 25268 29774
rect 25372 29826 25428 29828
rect 25372 29774 25374 29826
rect 25374 29774 25426 29826
rect 25426 29774 25428 29826
rect 25372 29772 25428 29774
rect 25532 29826 25588 29828
rect 25532 29774 25534 29826
rect 25534 29774 25586 29826
rect 25586 29774 25588 29826
rect 25532 29772 25588 29774
rect 25692 29826 25748 29828
rect 25692 29774 25694 29826
rect 25694 29774 25746 29826
rect 25746 29774 25748 29826
rect 25692 29772 25748 29774
rect 25852 29826 25908 29828
rect 25852 29774 25854 29826
rect 25854 29774 25906 29826
rect 25906 29774 25908 29826
rect 25852 29772 25908 29774
rect 26012 29826 26068 29828
rect 26012 29774 26014 29826
rect 26014 29774 26066 29826
rect 26066 29774 26068 29826
rect 26012 29772 26068 29774
rect 26172 29826 26228 29828
rect 26172 29774 26174 29826
rect 26174 29774 26226 29826
rect 26226 29774 26228 29826
rect 26172 29772 26228 29774
rect 26332 29826 26388 29828
rect 26332 29774 26334 29826
rect 26334 29774 26386 29826
rect 26386 29774 26388 29826
rect 26332 29772 26388 29774
rect 26492 29826 26548 29828
rect 26492 29774 26494 29826
rect 26494 29774 26546 29826
rect 26546 29774 26548 29826
rect 26492 29772 26548 29774
rect 26652 29826 26708 29828
rect 26652 29774 26654 29826
rect 26654 29774 26706 29826
rect 26706 29774 26708 29826
rect 26652 29772 26708 29774
rect 26812 29826 26868 29828
rect 26812 29774 26814 29826
rect 26814 29774 26866 29826
rect 26866 29774 26868 29826
rect 26812 29772 26868 29774
rect 26972 29826 27028 29828
rect 26972 29774 26974 29826
rect 26974 29774 27026 29826
rect 27026 29774 27028 29826
rect 26972 29772 27028 29774
rect 27132 29826 27188 29828
rect 27132 29774 27134 29826
rect 27134 29774 27186 29826
rect 27186 29774 27188 29826
rect 27132 29772 27188 29774
rect 27292 29826 27348 29828
rect 27292 29774 27294 29826
rect 27294 29774 27346 29826
rect 27346 29774 27348 29826
rect 27292 29772 27348 29774
rect 27452 29826 27508 29828
rect 27452 29774 27454 29826
rect 27454 29774 27506 29826
rect 27506 29774 27508 29826
rect 27452 29772 27508 29774
rect 27612 29826 27668 29828
rect 27612 29774 27614 29826
rect 27614 29774 27666 29826
rect 27666 29774 27668 29826
rect 27612 29772 27668 29774
rect 27772 29826 27828 29828
rect 27772 29774 27774 29826
rect 27774 29774 27826 29826
rect 27826 29774 27828 29826
rect 27772 29772 27828 29774
rect 27932 29826 27988 29828
rect 27932 29774 27934 29826
rect 27934 29774 27986 29826
rect 27986 29774 27988 29826
rect 27932 29772 27988 29774
rect 28092 29826 28148 29828
rect 28092 29774 28094 29826
rect 28094 29774 28146 29826
rect 28146 29774 28148 29826
rect 28092 29772 28148 29774
rect 28252 29826 28308 29828
rect 28252 29774 28254 29826
rect 28254 29774 28306 29826
rect 28306 29774 28308 29826
rect 28252 29772 28308 29774
rect 28412 29826 28468 29828
rect 28412 29774 28414 29826
rect 28414 29774 28466 29826
rect 28466 29774 28468 29826
rect 28412 29772 28468 29774
rect 28572 29826 28628 29828
rect 28572 29774 28574 29826
rect 28574 29774 28626 29826
rect 28626 29774 28628 29826
rect 28572 29772 28628 29774
rect 28732 29826 28788 29828
rect 28732 29774 28734 29826
rect 28734 29774 28786 29826
rect 28786 29774 28788 29826
rect 28732 29772 28788 29774
rect 28892 29826 28948 29828
rect 28892 29774 28894 29826
rect 28894 29774 28946 29826
rect 28946 29774 28948 29826
rect 28892 29772 28948 29774
rect 29052 29826 29108 29828
rect 29052 29774 29054 29826
rect 29054 29774 29106 29826
rect 29106 29774 29108 29826
rect 29052 29772 29108 29774
rect 29212 29826 29268 29828
rect 29212 29774 29214 29826
rect 29214 29774 29266 29826
rect 29266 29774 29268 29826
rect 29212 29772 29268 29774
rect 29372 29826 29428 29828
rect 29372 29774 29374 29826
rect 29374 29774 29426 29826
rect 29426 29774 29428 29826
rect 29372 29772 29428 29774
rect 29532 29772 29588 29828
rect 29852 29772 29908 29828
rect 33532 29826 33588 29828
rect 33532 29774 33534 29826
rect 33534 29774 33586 29826
rect 33586 29774 33588 29826
rect 33532 29772 33588 29774
rect 33692 29826 33748 29828
rect 33692 29774 33694 29826
rect 33694 29774 33746 29826
rect 33746 29774 33748 29826
rect 33692 29772 33748 29774
rect 33852 29826 33908 29828
rect 33852 29774 33854 29826
rect 33854 29774 33906 29826
rect 33906 29774 33908 29826
rect 33852 29772 33908 29774
rect 34012 29826 34068 29828
rect 34012 29774 34014 29826
rect 34014 29774 34066 29826
rect 34066 29774 34068 29826
rect 34012 29772 34068 29774
rect 34172 29826 34228 29828
rect 34172 29774 34174 29826
rect 34174 29774 34226 29826
rect 34226 29774 34228 29826
rect 34172 29772 34228 29774
rect 34332 29826 34388 29828
rect 34332 29774 34334 29826
rect 34334 29774 34386 29826
rect 34386 29774 34388 29826
rect 34332 29772 34388 29774
rect 34492 29826 34548 29828
rect 34492 29774 34494 29826
rect 34494 29774 34546 29826
rect 34546 29774 34548 29826
rect 34492 29772 34548 29774
rect 34652 29826 34708 29828
rect 34652 29774 34654 29826
rect 34654 29774 34706 29826
rect 34706 29774 34708 29826
rect 34652 29772 34708 29774
rect 34812 29826 34868 29828
rect 34812 29774 34814 29826
rect 34814 29774 34866 29826
rect 34866 29774 34868 29826
rect 34812 29772 34868 29774
rect 34972 29826 35028 29828
rect 34972 29774 34974 29826
rect 34974 29774 35026 29826
rect 35026 29774 35028 29826
rect 34972 29772 35028 29774
rect 35132 29826 35188 29828
rect 35132 29774 35134 29826
rect 35134 29774 35186 29826
rect 35186 29774 35188 29826
rect 35132 29772 35188 29774
rect 35292 29826 35348 29828
rect 35292 29774 35294 29826
rect 35294 29774 35346 29826
rect 35346 29774 35348 29826
rect 35292 29772 35348 29774
rect 35452 29826 35508 29828
rect 35452 29774 35454 29826
rect 35454 29774 35506 29826
rect 35506 29774 35508 29826
rect 35452 29772 35508 29774
rect 35612 29826 35668 29828
rect 35612 29774 35614 29826
rect 35614 29774 35666 29826
rect 35666 29774 35668 29826
rect 35612 29772 35668 29774
rect 35772 29826 35828 29828
rect 35772 29774 35774 29826
rect 35774 29774 35826 29826
rect 35826 29774 35828 29826
rect 35772 29772 35828 29774
rect 35932 29826 35988 29828
rect 35932 29774 35934 29826
rect 35934 29774 35986 29826
rect 35986 29774 35988 29826
rect 35932 29772 35988 29774
rect 36092 29826 36148 29828
rect 36092 29774 36094 29826
rect 36094 29774 36146 29826
rect 36146 29774 36148 29826
rect 36092 29772 36148 29774
rect 36252 29826 36308 29828
rect 36252 29774 36254 29826
rect 36254 29774 36306 29826
rect 36306 29774 36308 29826
rect 36252 29772 36308 29774
rect 36412 29826 36468 29828
rect 36412 29774 36414 29826
rect 36414 29774 36466 29826
rect 36466 29774 36468 29826
rect 36412 29772 36468 29774
rect 36572 29826 36628 29828
rect 36572 29774 36574 29826
rect 36574 29774 36626 29826
rect 36626 29774 36628 29826
rect 36572 29772 36628 29774
rect 36732 29826 36788 29828
rect 36732 29774 36734 29826
rect 36734 29774 36786 29826
rect 36786 29774 36788 29826
rect 36732 29772 36788 29774
rect 36892 29826 36948 29828
rect 36892 29774 36894 29826
rect 36894 29774 36946 29826
rect 36946 29774 36948 29826
rect 36892 29772 36948 29774
rect 37052 29826 37108 29828
rect 37052 29774 37054 29826
rect 37054 29774 37106 29826
rect 37106 29774 37108 29826
rect 37052 29772 37108 29774
rect 37212 29826 37268 29828
rect 37212 29774 37214 29826
rect 37214 29774 37266 29826
rect 37266 29774 37268 29826
rect 37212 29772 37268 29774
rect 37372 29826 37428 29828
rect 37372 29774 37374 29826
rect 37374 29774 37426 29826
rect 37426 29774 37428 29826
rect 37372 29772 37428 29774
rect 37532 29826 37588 29828
rect 37532 29774 37534 29826
rect 37534 29774 37586 29826
rect 37586 29774 37588 29826
rect 37532 29772 37588 29774
rect 37692 29826 37748 29828
rect 37692 29774 37694 29826
rect 37694 29774 37746 29826
rect 37746 29774 37748 29826
rect 37692 29772 37748 29774
rect 37852 29826 37908 29828
rect 37852 29774 37854 29826
rect 37854 29774 37906 29826
rect 37906 29774 37908 29826
rect 37852 29772 37908 29774
rect 38012 29826 38068 29828
rect 38012 29774 38014 29826
rect 38014 29774 38066 29826
rect 38066 29774 38068 29826
rect 38012 29772 38068 29774
rect 38172 29826 38228 29828
rect 38172 29774 38174 29826
rect 38174 29774 38226 29826
rect 38226 29774 38228 29826
rect 38172 29772 38228 29774
rect 38332 29826 38388 29828
rect 38332 29774 38334 29826
rect 38334 29774 38386 29826
rect 38386 29774 38388 29826
rect 38332 29772 38388 29774
rect 38492 29826 38548 29828
rect 38492 29774 38494 29826
rect 38494 29774 38546 29826
rect 38546 29774 38548 29826
rect 38492 29772 38548 29774
rect 38652 29826 38708 29828
rect 38652 29774 38654 29826
rect 38654 29774 38706 29826
rect 38706 29774 38708 29826
rect 38652 29772 38708 29774
rect 38812 29826 38868 29828
rect 38812 29774 38814 29826
rect 38814 29774 38866 29826
rect 38866 29774 38868 29826
rect 38812 29772 38868 29774
rect 38972 29826 39028 29828
rect 38972 29774 38974 29826
rect 38974 29774 39026 29826
rect 39026 29774 39028 29826
rect 38972 29772 39028 29774
rect 39132 29826 39188 29828
rect 39132 29774 39134 29826
rect 39134 29774 39186 29826
rect 39186 29774 39188 29826
rect 39132 29772 39188 29774
rect 39292 29826 39348 29828
rect 39292 29774 39294 29826
rect 39294 29774 39346 29826
rect 39346 29774 39348 29826
rect 39292 29772 39348 29774
rect 39452 29826 39508 29828
rect 39452 29774 39454 29826
rect 39454 29774 39506 29826
rect 39506 29774 39508 29826
rect 39452 29772 39508 29774
rect 39612 29826 39668 29828
rect 39612 29774 39614 29826
rect 39614 29774 39666 29826
rect 39666 29774 39668 29826
rect 39612 29772 39668 29774
rect 39772 29826 39828 29828
rect 39772 29774 39774 29826
rect 39774 29774 39826 29826
rect 39826 29774 39828 29826
rect 39772 29772 39828 29774
rect 39932 29826 39988 29828
rect 39932 29774 39934 29826
rect 39934 29774 39986 29826
rect 39986 29774 39988 29826
rect 39932 29772 39988 29774
rect 40092 29826 40148 29828
rect 40092 29774 40094 29826
rect 40094 29774 40146 29826
rect 40146 29774 40148 29826
rect 40092 29772 40148 29774
rect 40252 29826 40308 29828
rect 40252 29774 40254 29826
rect 40254 29774 40306 29826
rect 40306 29774 40308 29826
rect 40252 29772 40308 29774
rect 40412 29826 40468 29828
rect 40412 29774 40414 29826
rect 40414 29774 40466 29826
rect 40466 29774 40468 29826
rect 40412 29772 40468 29774
rect 40572 29826 40628 29828
rect 40572 29774 40574 29826
rect 40574 29774 40626 29826
rect 40626 29774 40628 29826
rect 40572 29772 40628 29774
rect 40732 29826 40788 29828
rect 40732 29774 40734 29826
rect 40734 29774 40786 29826
rect 40786 29774 40788 29826
rect 40732 29772 40788 29774
rect 40892 29826 40948 29828
rect 40892 29774 40894 29826
rect 40894 29774 40946 29826
rect 40946 29774 40948 29826
rect 40892 29772 40948 29774
rect 41052 29826 41108 29828
rect 41052 29774 41054 29826
rect 41054 29774 41106 29826
rect 41106 29774 41108 29826
rect 41052 29772 41108 29774
rect 41212 29826 41268 29828
rect 41212 29774 41214 29826
rect 41214 29774 41266 29826
rect 41266 29774 41268 29826
rect 41212 29772 41268 29774
rect 41372 29826 41428 29828
rect 41372 29774 41374 29826
rect 41374 29774 41426 29826
rect 41426 29774 41428 29826
rect 41372 29772 41428 29774
rect 41532 29826 41588 29828
rect 41532 29774 41534 29826
rect 41534 29774 41586 29826
rect 41586 29774 41588 29826
rect 41532 29772 41588 29774
rect 41692 29826 41748 29828
rect 41692 29774 41694 29826
rect 41694 29774 41746 29826
rect 41746 29774 41748 29826
rect 41692 29772 41748 29774
rect 41852 29826 41908 29828
rect 41852 29774 41854 29826
rect 41854 29774 41906 29826
rect 41906 29774 41908 29826
rect 41852 29772 41908 29774
rect 12172 29612 12228 29668
rect 22732 29612 22788 29668
rect 29692 29612 29748 29668
rect 12 29506 68 29508
rect 12 29454 14 29506
rect 14 29454 66 29506
rect 66 29454 68 29506
rect 12 29452 68 29454
rect 172 29506 228 29508
rect 172 29454 174 29506
rect 174 29454 226 29506
rect 226 29454 228 29506
rect 172 29452 228 29454
rect 332 29506 388 29508
rect 332 29454 334 29506
rect 334 29454 386 29506
rect 386 29454 388 29506
rect 332 29452 388 29454
rect 492 29506 548 29508
rect 492 29454 494 29506
rect 494 29454 546 29506
rect 546 29454 548 29506
rect 492 29452 548 29454
rect 652 29506 708 29508
rect 652 29454 654 29506
rect 654 29454 706 29506
rect 706 29454 708 29506
rect 652 29452 708 29454
rect 812 29506 868 29508
rect 812 29454 814 29506
rect 814 29454 866 29506
rect 866 29454 868 29506
rect 812 29452 868 29454
rect 972 29506 1028 29508
rect 972 29454 974 29506
rect 974 29454 1026 29506
rect 1026 29454 1028 29506
rect 972 29452 1028 29454
rect 1132 29506 1188 29508
rect 1132 29454 1134 29506
rect 1134 29454 1186 29506
rect 1186 29454 1188 29506
rect 1132 29452 1188 29454
rect 1292 29506 1348 29508
rect 1292 29454 1294 29506
rect 1294 29454 1346 29506
rect 1346 29454 1348 29506
rect 1292 29452 1348 29454
rect 1452 29506 1508 29508
rect 1452 29454 1454 29506
rect 1454 29454 1506 29506
rect 1506 29454 1508 29506
rect 1452 29452 1508 29454
rect 1612 29506 1668 29508
rect 1612 29454 1614 29506
rect 1614 29454 1666 29506
rect 1666 29454 1668 29506
rect 1612 29452 1668 29454
rect 1772 29506 1828 29508
rect 1772 29454 1774 29506
rect 1774 29454 1826 29506
rect 1826 29454 1828 29506
rect 1772 29452 1828 29454
rect 1932 29506 1988 29508
rect 1932 29454 1934 29506
rect 1934 29454 1986 29506
rect 1986 29454 1988 29506
rect 1932 29452 1988 29454
rect 2092 29506 2148 29508
rect 2092 29454 2094 29506
rect 2094 29454 2146 29506
rect 2146 29454 2148 29506
rect 2092 29452 2148 29454
rect 2252 29506 2308 29508
rect 2252 29454 2254 29506
rect 2254 29454 2306 29506
rect 2306 29454 2308 29506
rect 2252 29452 2308 29454
rect 2412 29506 2468 29508
rect 2412 29454 2414 29506
rect 2414 29454 2466 29506
rect 2466 29454 2468 29506
rect 2412 29452 2468 29454
rect 2572 29506 2628 29508
rect 2572 29454 2574 29506
rect 2574 29454 2626 29506
rect 2626 29454 2628 29506
rect 2572 29452 2628 29454
rect 2732 29506 2788 29508
rect 2732 29454 2734 29506
rect 2734 29454 2786 29506
rect 2786 29454 2788 29506
rect 2732 29452 2788 29454
rect 2892 29506 2948 29508
rect 2892 29454 2894 29506
rect 2894 29454 2946 29506
rect 2946 29454 2948 29506
rect 2892 29452 2948 29454
rect 3052 29506 3108 29508
rect 3052 29454 3054 29506
rect 3054 29454 3106 29506
rect 3106 29454 3108 29506
rect 3052 29452 3108 29454
rect 3212 29506 3268 29508
rect 3212 29454 3214 29506
rect 3214 29454 3266 29506
rect 3266 29454 3268 29506
rect 3212 29452 3268 29454
rect 3372 29506 3428 29508
rect 3372 29454 3374 29506
rect 3374 29454 3426 29506
rect 3426 29454 3428 29506
rect 3372 29452 3428 29454
rect 3532 29506 3588 29508
rect 3532 29454 3534 29506
rect 3534 29454 3586 29506
rect 3586 29454 3588 29506
rect 3532 29452 3588 29454
rect 3692 29506 3748 29508
rect 3692 29454 3694 29506
rect 3694 29454 3746 29506
rect 3746 29454 3748 29506
rect 3692 29452 3748 29454
rect 3852 29506 3908 29508
rect 3852 29454 3854 29506
rect 3854 29454 3906 29506
rect 3906 29454 3908 29506
rect 3852 29452 3908 29454
rect 4012 29506 4068 29508
rect 4012 29454 4014 29506
rect 4014 29454 4066 29506
rect 4066 29454 4068 29506
rect 4012 29452 4068 29454
rect 4172 29506 4228 29508
rect 4172 29454 4174 29506
rect 4174 29454 4226 29506
rect 4226 29454 4228 29506
rect 4172 29452 4228 29454
rect 4332 29506 4388 29508
rect 4332 29454 4334 29506
rect 4334 29454 4386 29506
rect 4386 29454 4388 29506
rect 4332 29452 4388 29454
rect 4492 29506 4548 29508
rect 4492 29454 4494 29506
rect 4494 29454 4546 29506
rect 4546 29454 4548 29506
rect 4492 29452 4548 29454
rect 4652 29506 4708 29508
rect 4652 29454 4654 29506
rect 4654 29454 4706 29506
rect 4706 29454 4708 29506
rect 4652 29452 4708 29454
rect 4812 29506 4868 29508
rect 4812 29454 4814 29506
rect 4814 29454 4866 29506
rect 4866 29454 4868 29506
rect 4812 29452 4868 29454
rect 4972 29506 5028 29508
rect 4972 29454 4974 29506
rect 4974 29454 5026 29506
rect 5026 29454 5028 29506
rect 4972 29452 5028 29454
rect 5132 29506 5188 29508
rect 5132 29454 5134 29506
rect 5134 29454 5186 29506
rect 5186 29454 5188 29506
rect 5132 29452 5188 29454
rect 5292 29506 5348 29508
rect 5292 29454 5294 29506
rect 5294 29454 5346 29506
rect 5346 29454 5348 29506
rect 5292 29452 5348 29454
rect 5452 29506 5508 29508
rect 5452 29454 5454 29506
rect 5454 29454 5506 29506
rect 5506 29454 5508 29506
rect 5452 29452 5508 29454
rect 5612 29506 5668 29508
rect 5612 29454 5614 29506
rect 5614 29454 5666 29506
rect 5666 29454 5668 29506
rect 5612 29452 5668 29454
rect 5772 29506 5828 29508
rect 5772 29454 5774 29506
rect 5774 29454 5826 29506
rect 5826 29454 5828 29506
rect 5772 29452 5828 29454
rect 5932 29506 5988 29508
rect 5932 29454 5934 29506
rect 5934 29454 5986 29506
rect 5986 29454 5988 29506
rect 5932 29452 5988 29454
rect 6092 29506 6148 29508
rect 6092 29454 6094 29506
rect 6094 29454 6146 29506
rect 6146 29454 6148 29506
rect 6092 29452 6148 29454
rect 6252 29506 6308 29508
rect 6252 29454 6254 29506
rect 6254 29454 6306 29506
rect 6306 29454 6308 29506
rect 6252 29452 6308 29454
rect 6412 29506 6468 29508
rect 6412 29454 6414 29506
rect 6414 29454 6466 29506
rect 6466 29454 6468 29506
rect 6412 29452 6468 29454
rect 6572 29506 6628 29508
rect 6572 29454 6574 29506
rect 6574 29454 6626 29506
rect 6626 29454 6628 29506
rect 6572 29452 6628 29454
rect 6732 29506 6788 29508
rect 6732 29454 6734 29506
rect 6734 29454 6786 29506
rect 6786 29454 6788 29506
rect 6732 29452 6788 29454
rect 6892 29506 6948 29508
rect 6892 29454 6894 29506
rect 6894 29454 6946 29506
rect 6946 29454 6948 29506
rect 6892 29452 6948 29454
rect 7052 29506 7108 29508
rect 7052 29454 7054 29506
rect 7054 29454 7106 29506
rect 7106 29454 7108 29506
rect 7052 29452 7108 29454
rect 7212 29506 7268 29508
rect 7212 29454 7214 29506
rect 7214 29454 7266 29506
rect 7266 29454 7268 29506
rect 7212 29452 7268 29454
rect 7372 29506 7428 29508
rect 7372 29454 7374 29506
rect 7374 29454 7426 29506
rect 7426 29454 7428 29506
rect 7372 29452 7428 29454
rect 7532 29506 7588 29508
rect 7532 29454 7534 29506
rect 7534 29454 7586 29506
rect 7586 29454 7588 29506
rect 7532 29452 7588 29454
rect 7692 29506 7748 29508
rect 7692 29454 7694 29506
rect 7694 29454 7746 29506
rect 7746 29454 7748 29506
rect 7692 29452 7748 29454
rect 7852 29506 7908 29508
rect 7852 29454 7854 29506
rect 7854 29454 7906 29506
rect 7906 29454 7908 29506
rect 7852 29452 7908 29454
rect 8012 29506 8068 29508
rect 8012 29454 8014 29506
rect 8014 29454 8066 29506
rect 8066 29454 8068 29506
rect 8012 29452 8068 29454
rect 8172 29506 8228 29508
rect 8172 29454 8174 29506
rect 8174 29454 8226 29506
rect 8226 29454 8228 29506
rect 8172 29452 8228 29454
rect 8332 29506 8388 29508
rect 8332 29454 8334 29506
rect 8334 29454 8386 29506
rect 8386 29454 8388 29506
rect 8332 29452 8388 29454
rect 12012 29452 12068 29508
rect 12332 29452 12388 29508
rect 12492 29506 12548 29508
rect 12492 29454 12494 29506
rect 12494 29454 12546 29506
rect 12546 29454 12548 29506
rect 12492 29452 12548 29454
rect 12652 29506 12708 29508
rect 12652 29454 12654 29506
rect 12654 29454 12706 29506
rect 12706 29454 12708 29506
rect 12652 29452 12708 29454
rect 12812 29506 12868 29508
rect 12812 29454 12814 29506
rect 12814 29454 12866 29506
rect 12866 29454 12868 29506
rect 12812 29452 12868 29454
rect 12972 29506 13028 29508
rect 12972 29454 12974 29506
rect 12974 29454 13026 29506
rect 13026 29454 13028 29506
rect 12972 29452 13028 29454
rect 13132 29506 13188 29508
rect 13132 29454 13134 29506
rect 13134 29454 13186 29506
rect 13186 29454 13188 29506
rect 13132 29452 13188 29454
rect 13292 29506 13348 29508
rect 13292 29454 13294 29506
rect 13294 29454 13346 29506
rect 13346 29454 13348 29506
rect 13292 29452 13348 29454
rect 13452 29506 13508 29508
rect 13452 29454 13454 29506
rect 13454 29454 13506 29506
rect 13506 29454 13508 29506
rect 13452 29452 13508 29454
rect 13612 29506 13668 29508
rect 13612 29454 13614 29506
rect 13614 29454 13666 29506
rect 13666 29454 13668 29506
rect 13612 29452 13668 29454
rect 13772 29506 13828 29508
rect 13772 29454 13774 29506
rect 13774 29454 13826 29506
rect 13826 29454 13828 29506
rect 13772 29452 13828 29454
rect 13932 29506 13988 29508
rect 13932 29454 13934 29506
rect 13934 29454 13986 29506
rect 13986 29454 13988 29506
rect 13932 29452 13988 29454
rect 14092 29506 14148 29508
rect 14092 29454 14094 29506
rect 14094 29454 14146 29506
rect 14146 29454 14148 29506
rect 14092 29452 14148 29454
rect 14252 29506 14308 29508
rect 14252 29454 14254 29506
rect 14254 29454 14306 29506
rect 14306 29454 14308 29506
rect 14252 29452 14308 29454
rect 14412 29506 14468 29508
rect 14412 29454 14414 29506
rect 14414 29454 14466 29506
rect 14466 29454 14468 29506
rect 14412 29452 14468 29454
rect 14572 29506 14628 29508
rect 14572 29454 14574 29506
rect 14574 29454 14626 29506
rect 14626 29454 14628 29506
rect 14572 29452 14628 29454
rect 14732 29506 14788 29508
rect 14732 29454 14734 29506
rect 14734 29454 14786 29506
rect 14786 29454 14788 29506
rect 14732 29452 14788 29454
rect 14892 29506 14948 29508
rect 14892 29454 14894 29506
rect 14894 29454 14946 29506
rect 14946 29454 14948 29506
rect 14892 29452 14948 29454
rect 15052 29506 15108 29508
rect 15052 29454 15054 29506
rect 15054 29454 15106 29506
rect 15106 29454 15108 29506
rect 15052 29452 15108 29454
rect 15212 29506 15268 29508
rect 15212 29454 15214 29506
rect 15214 29454 15266 29506
rect 15266 29454 15268 29506
rect 15212 29452 15268 29454
rect 15372 29506 15428 29508
rect 15372 29454 15374 29506
rect 15374 29454 15426 29506
rect 15426 29454 15428 29506
rect 15372 29452 15428 29454
rect 15532 29506 15588 29508
rect 15532 29454 15534 29506
rect 15534 29454 15586 29506
rect 15586 29454 15588 29506
rect 15532 29452 15588 29454
rect 15692 29506 15748 29508
rect 15692 29454 15694 29506
rect 15694 29454 15746 29506
rect 15746 29454 15748 29506
rect 15692 29452 15748 29454
rect 15852 29506 15908 29508
rect 15852 29454 15854 29506
rect 15854 29454 15906 29506
rect 15906 29454 15908 29506
rect 15852 29452 15908 29454
rect 16012 29506 16068 29508
rect 16012 29454 16014 29506
rect 16014 29454 16066 29506
rect 16066 29454 16068 29506
rect 16012 29452 16068 29454
rect 16172 29506 16228 29508
rect 16172 29454 16174 29506
rect 16174 29454 16226 29506
rect 16226 29454 16228 29506
rect 16172 29452 16228 29454
rect 16332 29506 16388 29508
rect 16332 29454 16334 29506
rect 16334 29454 16386 29506
rect 16386 29454 16388 29506
rect 16332 29452 16388 29454
rect 16492 29506 16548 29508
rect 16492 29454 16494 29506
rect 16494 29454 16546 29506
rect 16546 29454 16548 29506
rect 16492 29452 16548 29454
rect 16652 29506 16708 29508
rect 16652 29454 16654 29506
rect 16654 29454 16706 29506
rect 16706 29454 16708 29506
rect 16652 29452 16708 29454
rect 16812 29506 16868 29508
rect 16812 29454 16814 29506
rect 16814 29454 16866 29506
rect 16866 29454 16868 29506
rect 16812 29452 16868 29454
rect 16972 29506 17028 29508
rect 16972 29454 16974 29506
rect 16974 29454 17026 29506
rect 17026 29454 17028 29506
rect 16972 29452 17028 29454
rect 17132 29506 17188 29508
rect 17132 29454 17134 29506
rect 17134 29454 17186 29506
rect 17186 29454 17188 29506
rect 17132 29452 17188 29454
rect 17292 29506 17348 29508
rect 17292 29454 17294 29506
rect 17294 29454 17346 29506
rect 17346 29454 17348 29506
rect 17292 29452 17348 29454
rect 17452 29506 17508 29508
rect 17452 29454 17454 29506
rect 17454 29454 17506 29506
rect 17506 29454 17508 29506
rect 17452 29452 17508 29454
rect 17612 29506 17668 29508
rect 17612 29454 17614 29506
rect 17614 29454 17666 29506
rect 17666 29454 17668 29506
rect 17612 29452 17668 29454
rect 17772 29506 17828 29508
rect 17772 29454 17774 29506
rect 17774 29454 17826 29506
rect 17826 29454 17828 29506
rect 17772 29452 17828 29454
rect 17932 29506 17988 29508
rect 17932 29454 17934 29506
rect 17934 29454 17986 29506
rect 17986 29454 17988 29506
rect 17932 29452 17988 29454
rect 18092 29506 18148 29508
rect 18092 29454 18094 29506
rect 18094 29454 18146 29506
rect 18146 29454 18148 29506
rect 18092 29452 18148 29454
rect 18252 29506 18308 29508
rect 18252 29454 18254 29506
rect 18254 29454 18306 29506
rect 18306 29454 18308 29506
rect 18252 29452 18308 29454
rect 18412 29506 18468 29508
rect 18412 29454 18414 29506
rect 18414 29454 18466 29506
rect 18466 29454 18468 29506
rect 18412 29452 18468 29454
rect 18572 29506 18628 29508
rect 18572 29454 18574 29506
rect 18574 29454 18626 29506
rect 18626 29454 18628 29506
rect 18572 29452 18628 29454
rect 18732 29506 18788 29508
rect 18732 29454 18734 29506
rect 18734 29454 18786 29506
rect 18786 29454 18788 29506
rect 18732 29452 18788 29454
rect 18892 29506 18948 29508
rect 18892 29454 18894 29506
rect 18894 29454 18946 29506
rect 18946 29454 18948 29506
rect 18892 29452 18948 29454
rect 22572 29452 22628 29508
rect 22892 29452 22948 29508
rect 23132 29506 23188 29508
rect 23132 29454 23134 29506
rect 23134 29454 23186 29506
rect 23186 29454 23188 29506
rect 23132 29452 23188 29454
rect 23292 29506 23348 29508
rect 23292 29454 23294 29506
rect 23294 29454 23346 29506
rect 23346 29454 23348 29506
rect 23292 29452 23348 29454
rect 23452 29506 23508 29508
rect 23452 29454 23454 29506
rect 23454 29454 23506 29506
rect 23506 29454 23508 29506
rect 23452 29452 23508 29454
rect 23612 29506 23668 29508
rect 23612 29454 23614 29506
rect 23614 29454 23666 29506
rect 23666 29454 23668 29506
rect 23612 29452 23668 29454
rect 23772 29506 23828 29508
rect 23772 29454 23774 29506
rect 23774 29454 23826 29506
rect 23826 29454 23828 29506
rect 23772 29452 23828 29454
rect 23932 29506 23988 29508
rect 23932 29454 23934 29506
rect 23934 29454 23986 29506
rect 23986 29454 23988 29506
rect 23932 29452 23988 29454
rect 24092 29506 24148 29508
rect 24092 29454 24094 29506
rect 24094 29454 24146 29506
rect 24146 29454 24148 29506
rect 24092 29452 24148 29454
rect 24252 29506 24308 29508
rect 24252 29454 24254 29506
rect 24254 29454 24306 29506
rect 24306 29454 24308 29506
rect 24252 29452 24308 29454
rect 24412 29506 24468 29508
rect 24412 29454 24414 29506
rect 24414 29454 24466 29506
rect 24466 29454 24468 29506
rect 24412 29452 24468 29454
rect 24572 29506 24628 29508
rect 24572 29454 24574 29506
rect 24574 29454 24626 29506
rect 24626 29454 24628 29506
rect 24572 29452 24628 29454
rect 24732 29506 24788 29508
rect 24732 29454 24734 29506
rect 24734 29454 24786 29506
rect 24786 29454 24788 29506
rect 24732 29452 24788 29454
rect 24892 29506 24948 29508
rect 24892 29454 24894 29506
rect 24894 29454 24946 29506
rect 24946 29454 24948 29506
rect 24892 29452 24948 29454
rect 25052 29506 25108 29508
rect 25052 29454 25054 29506
rect 25054 29454 25106 29506
rect 25106 29454 25108 29506
rect 25052 29452 25108 29454
rect 25212 29506 25268 29508
rect 25212 29454 25214 29506
rect 25214 29454 25266 29506
rect 25266 29454 25268 29506
rect 25212 29452 25268 29454
rect 25372 29506 25428 29508
rect 25372 29454 25374 29506
rect 25374 29454 25426 29506
rect 25426 29454 25428 29506
rect 25372 29452 25428 29454
rect 25532 29506 25588 29508
rect 25532 29454 25534 29506
rect 25534 29454 25586 29506
rect 25586 29454 25588 29506
rect 25532 29452 25588 29454
rect 25692 29506 25748 29508
rect 25692 29454 25694 29506
rect 25694 29454 25746 29506
rect 25746 29454 25748 29506
rect 25692 29452 25748 29454
rect 25852 29506 25908 29508
rect 25852 29454 25854 29506
rect 25854 29454 25906 29506
rect 25906 29454 25908 29506
rect 25852 29452 25908 29454
rect 26012 29506 26068 29508
rect 26012 29454 26014 29506
rect 26014 29454 26066 29506
rect 26066 29454 26068 29506
rect 26012 29452 26068 29454
rect 26172 29506 26228 29508
rect 26172 29454 26174 29506
rect 26174 29454 26226 29506
rect 26226 29454 26228 29506
rect 26172 29452 26228 29454
rect 26332 29506 26388 29508
rect 26332 29454 26334 29506
rect 26334 29454 26386 29506
rect 26386 29454 26388 29506
rect 26332 29452 26388 29454
rect 26492 29506 26548 29508
rect 26492 29454 26494 29506
rect 26494 29454 26546 29506
rect 26546 29454 26548 29506
rect 26492 29452 26548 29454
rect 26652 29506 26708 29508
rect 26652 29454 26654 29506
rect 26654 29454 26706 29506
rect 26706 29454 26708 29506
rect 26652 29452 26708 29454
rect 26812 29506 26868 29508
rect 26812 29454 26814 29506
rect 26814 29454 26866 29506
rect 26866 29454 26868 29506
rect 26812 29452 26868 29454
rect 26972 29506 27028 29508
rect 26972 29454 26974 29506
rect 26974 29454 27026 29506
rect 27026 29454 27028 29506
rect 26972 29452 27028 29454
rect 27132 29506 27188 29508
rect 27132 29454 27134 29506
rect 27134 29454 27186 29506
rect 27186 29454 27188 29506
rect 27132 29452 27188 29454
rect 27292 29506 27348 29508
rect 27292 29454 27294 29506
rect 27294 29454 27346 29506
rect 27346 29454 27348 29506
rect 27292 29452 27348 29454
rect 27452 29506 27508 29508
rect 27452 29454 27454 29506
rect 27454 29454 27506 29506
rect 27506 29454 27508 29506
rect 27452 29452 27508 29454
rect 27612 29506 27668 29508
rect 27612 29454 27614 29506
rect 27614 29454 27666 29506
rect 27666 29454 27668 29506
rect 27612 29452 27668 29454
rect 27772 29506 27828 29508
rect 27772 29454 27774 29506
rect 27774 29454 27826 29506
rect 27826 29454 27828 29506
rect 27772 29452 27828 29454
rect 27932 29506 27988 29508
rect 27932 29454 27934 29506
rect 27934 29454 27986 29506
rect 27986 29454 27988 29506
rect 27932 29452 27988 29454
rect 28092 29506 28148 29508
rect 28092 29454 28094 29506
rect 28094 29454 28146 29506
rect 28146 29454 28148 29506
rect 28092 29452 28148 29454
rect 28252 29506 28308 29508
rect 28252 29454 28254 29506
rect 28254 29454 28306 29506
rect 28306 29454 28308 29506
rect 28252 29452 28308 29454
rect 28412 29506 28468 29508
rect 28412 29454 28414 29506
rect 28414 29454 28466 29506
rect 28466 29454 28468 29506
rect 28412 29452 28468 29454
rect 28572 29506 28628 29508
rect 28572 29454 28574 29506
rect 28574 29454 28626 29506
rect 28626 29454 28628 29506
rect 28572 29452 28628 29454
rect 28732 29506 28788 29508
rect 28732 29454 28734 29506
rect 28734 29454 28786 29506
rect 28786 29454 28788 29506
rect 28732 29452 28788 29454
rect 28892 29506 28948 29508
rect 28892 29454 28894 29506
rect 28894 29454 28946 29506
rect 28946 29454 28948 29506
rect 28892 29452 28948 29454
rect 29052 29506 29108 29508
rect 29052 29454 29054 29506
rect 29054 29454 29106 29506
rect 29106 29454 29108 29506
rect 29052 29452 29108 29454
rect 29212 29506 29268 29508
rect 29212 29454 29214 29506
rect 29214 29454 29266 29506
rect 29266 29454 29268 29506
rect 29212 29452 29268 29454
rect 29372 29506 29428 29508
rect 29372 29454 29374 29506
rect 29374 29454 29426 29506
rect 29426 29454 29428 29506
rect 29372 29452 29428 29454
rect 29532 29452 29588 29508
rect 29852 29452 29908 29508
rect 33532 29506 33588 29508
rect 33532 29454 33534 29506
rect 33534 29454 33586 29506
rect 33586 29454 33588 29506
rect 33532 29452 33588 29454
rect 33692 29506 33748 29508
rect 33692 29454 33694 29506
rect 33694 29454 33746 29506
rect 33746 29454 33748 29506
rect 33692 29452 33748 29454
rect 33852 29506 33908 29508
rect 33852 29454 33854 29506
rect 33854 29454 33906 29506
rect 33906 29454 33908 29506
rect 33852 29452 33908 29454
rect 34012 29506 34068 29508
rect 34012 29454 34014 29506
rect 34014 29454 34066 29506
rect 34066 29454 34068 29506
rect 34012 29452 34068 29454
rect 34172 29506 34228 29508
rect 34172 29454 34174 29506
rect 34174 29454 34226 29506
rect 34226 29454 34228 29506
rect 34172 29452 34228 29454
rect 34332 29506 34388 29508
rect 34332 29454 34334 29506
rect 34334 29454 34386 29506
rect 34386 29454 34388 29506
rect 34332 29452 34388 29454
rect 34492 29506 34548 29508
rect 34492 29454 34494 29506
rect 34494 29454 34546 29506
rect 34546 29454 34548 29506
rect 34492 29452 34548 29454
rect 34652 29506 34708 29508
rect 34652 29454 34654 29506
rect 34654 29454 34706 29506
rect 34706 29454 34708 29506
rect 34652 29452 34708 29454
rect 34812 29506 34868 29508
rect 34812 29454 34814 29506
rect 34814 29454 34866 29506
rect 34866 29454 34868 29506
rect 34812 29452 34868 29454
rect 34972 29506 35028 29508
rect 34972 29454 34974 29506
rect 34974 29454 35026 29506
rect 35026 29454 35028 29506
rect 34972 29452 35028 29454
rect 35132 29506 35188 29508
rect 35132 29454 35134 29506
rect 35134 29454 35186 29506
rect 35186 29454 35188 29506
rect 35132 29452 35188 29454
rect 35292 29506 35348 29508
rect 35292 29454 35294 29506
rect 35294 29454 35346 29506
rect 35346 29454 35348 29506
rect 35292 29452 35348 29454
rect 35452 29506 35508 29508
rect 35452 29454 35454 29506
rect 35454 29454 35506 29506
rect 35506 29454 35508 29506
rect 35452 29452 35508 29454
rect 35612 29506 35668 29508
rect 35612 29454 35614 29506
rect 35614 29454 35666 29506
rect 35666 29454 35668 29506
rect 35612 29452 35668 29454
rect 35772 29506 35828 29508
rect 35772 29454 35774 29506
rect 35774 29454 35826 29506
rect 35826 29454 35828 29506
rect 35772 29452 35828 29454
rect 35932 29506 35988 29508
rect 35932 29454 35934 29506
rect 35934 29454 35986 29506
rect 35986 29454 35988 29506
rect 35932 29452 35988 29454
rect 36092 29506 36148 29508
rect 36092 29454 36094 29506
rect 36094 29454 36146 29506
rect 36146 29454 36148 29506
rect 36092 29452 36148 29454
rect 36252 29506 36308 29508
rect 36252 29454 36254 29506
rect 36254 29454 36306 29506
rect 36306 29454 36308 29506
rect 36252 29452 36308 29454
rect 36412 29506 36468 29508
rect 36412 29454 36414 29506
rect 36414 29454 36466 29506
rect 36466 29454 36468 29506
rect 36412 29452 36468 29454
rect 36572 29506 36628 29508
rect 36572 29454 36574 29506
rect 36574 29454 36626 29506
rect 36626 29454 36628 29506
rect 36572 29452 36628 29454
rect 36732 29506 36788 29508
rect 36732 29454 36734 29506
rect 36734 29454 36786 29506
rect 36786 29454 36788 29506
rect 36732 29452 36788 29454
rect 36892 29506 36948 29508
rect 36892 29454 36894 29506
rect 36894 29454 36946 29506
rect 36946 29454 36948 29506
rect 36892 29452 36948 29454
rect 37052 29506 37108 29508
rect 37052 29454 37054 29506
rect 37054 29454 37106 29506
rect 37106 29454 37108 29506
rect 37052 29452 37108 29454
rect 37212 29506 37268 29508
rect 37212 29454 37214 29506
rect 37214 29454 37266 29506
rect 37266 29454 37268 29506
rect 37212 29452 37268 29454
rect 37372 29506 37428 29508
rect 37372 29454 37374 29506
rect 37374 29454 37426 29506
rect 37426 29454 37428 29506
rect 37372 29452 37428 29454
rect 37532 29506 37588 29508
rect 37532 29454 37534 29506
rect 37534 29454 37586 29506
rect 37586 29454 37588 29506
rect 37532 29452 37588 29454
rect 37692 29506 37748 29508
rect 37692 29454 37694 29506
rect 37694 29454 37746 29506
rect 37746 29454 37748 29506
rect 37692 29452 37748 29454
rect 37852 29506 37908 29508
rect 37852 29454 37854 29506
rect 37854 29454 37906 29506
rect 37906 29454 37908 29506
rect 37852 29452 37908 29454
rect 38012 29506 38068 29508
rect 38012 29454 38014 29506
rect 38014 29454 38066 29506
rect 38066 29454 38068 29506
rect 38012 29452 38068 29454
rect 38172 29506 38228 29508
rect 38172 29454 38174 29506
rect 38174 29454 38226 29506
rect 38226 29454 38228 29506
rect 38172 29452 38228 29454
rect 38332 29506 38388 29508
rect 38332 29454 38334 29506
rect 38334 29454 38386 29506
rect 38386 29454 38388 29506
rect 38332 29452 38388 29454
rect 38492 29506 38548 29508
rect 38492 29454 38494 29506
rect 38494 29454 38546 29506
rect 38546 29454 38548 29506
rect 38492 29452 38548 29454
rect 38652 29506 38708 29508
rect 38652 29454 38654 29506
rect 38654 29454 38706 29506
rect 38706 29454 38708 29506
rect 38652 29452 38708 29454
rect 38812 29506 38868 29508
rect 38812 29454 38814 29506
rect 38814 29454 38866 29506
rect 38866 29454 38868 29506
rect 38812 29452 38868 29454
rect 38972 29506 39028 29508
rect 38972 29454 38974 29506
rect 38974 29454 39026 29506
rect 39026 29454 39028 29506
rect 38972 29452 39028 29454
rect 39132 29506 39188 29508
rect 39132 29454 39134 29506
rect 39134 29454 39186 29506
rect 39186 29454 39188 29506
rect 39132 29452 39188 29454
rect 39292 29506 39348 29508
rect 39292 29454 39294 29506
rect 39294 29454 39346 29506
rect 39346 29454 39348 29506
rect 39292 29452 39348 29454
rect 39452 29506 39508 29508
rect 39452 29454 39454 29506
rect 39454 29454 39506 29506
rect 39506 29454 39508 29506
rect 39452 29452 39508 29454
rect 39612 29506 39668 29508
rect 39612 29454 39614 29506
rect 39614 29454 39666 29506
rect 39666 29454 39668 29506
rect 39612 29452 39668 29454
rect 39772 29506 39828 29508
rect 39772 29454 39774 29506
rect 39774 29454 39826 29506
rect 39826 29454 39828 29506
rect 39772 29452 39828 29454
rect 39932 29506 39988 29508
rect 39932 29454 39934 29506
rect 39934 29454 39986 29506
rect 39986 29454 39988 29506
rect 39932 29452 39988 29454
rect 40092 29506 40148 29508
rect 40092 29454 40094 29506
rect 40094 29454 40146 29506
rect 40146 29454 40148 29506
rect 40092 29452 40148 29454
rect 40252 29506 40308 29508
rect 40252 29454 40254 29506
rect 40254 29454 40306 29506
rect 40306 29454 40308 29506
rect 40252 29452 40308 29454
rect 40412 29506 40468 29508
rect 40412 29454 40414 29506
rect 40414 29454 40466 29506
rect 40466 29454 40468 29506
rect 40412 29452 40468 29454
rect 40572 29506 40628 29508
rect 40572 29454 40574 29506
rect 40574 29454 40626 29506
rect 40626 29454 40628 29506
rect 40572 29452 40628 29454
rect 40732 29506 40788 29508
rect 40732 29454 40734 29506
rect 40734 29454 40786 29506
rect 40786 29454 40788 29506
rect 40732 29452 40788 29454
rect 40892 29506 40948 29508
rect 40892 29454 40894 29506
rect 40894 29454 40946 29506
rect 40946 29454 40948 29506
rect 40892 29452 40948 29454
rect 41052 29506 41108 29508
rect 41052 29454 41054 29506
rect 41054 29454 41106 29506
rect 41106 29454 41108 29506
rect 41052 29452 41108 29454
rect 41212 29506 41268 29508
rect 41212 29454 41214 29506
rect 41214 29454 41266 29506
rect 41266 29454 41268 29506
rect 41212 29452 41268 29454
rect 41372 29506 41428 29508
rect 41372 29454 41374 29506
rect 41374 29454 41426 29506
rect 41426 29454 41428 29506
rect 41372 29452 41428 29454
rect 41532 29506 41588 29508
rect 41532 29454 41534 29506
rect 41534 29454 41586 29506
rect 41586 29454 41588 29506
rect 41532 29452 41588 29454
rect 41692 29506 41748 29508
rect 41692 29454 41694 29506
rect 41694 29454 41746 29506
rect 41746 29454 41748 29506
rect 41692 29452 41748 29454
rect 41852 29506 41908 29508
rect 41852 29454 41854 29506
rect 41854 29454 41906 29506
rect 41906 29454 41908 29506
rect 41852 29452 41908 29454
<< metal3 >>
rect 0 37348 80 37360
rect 0 37292 12 37348
rect 68 37292 80 37348
rect 0 37028 80 37292
rect 0 36972 12 37028
rect 68 36972 80 37028
rect 0 36960 80 36972
rect 160 37348 240 37360
rect 160 37292 172 37348
rect 228 37292 240 37348
rect 160 37028 240 37292
rect 160 36972 172 37028
rect 228 36972 240 37028
rect 160 36960 240 36972
rect 320 37348 400 37360
rect 320 37292 332 37348
rect 388 37292 400 37348
rect 320 37028 400 37292
rect 320 36972 332 37028
rect 388 36972 400 37028
rect 320 36960 400 36972
rect 480 37348 560 37360
rect 480 37292 492 37348
rect 548 37292 560 37348
rect 480 37028 560 37292
rect 480 36972 492 37028
rect 548 36972 560 37028
rect 480 36960 560 36972
rect 640 37348 720 37360
rect 640 37292 652 37348
rect 708 37292 720 37348
rect 640 37028 720 37292
rect 640 36972 652 37028
rect 708 36972 720 37028
rect 640 36960 720 36972
rect 800 37348 880 37360
rect 800 37292 812 37348
rect 868 37292 880 37348
rect 800 37028 880 37292
rect 800 36972 812 37028
rect 868 36972 880 37028
rect 800 36960 880 36972
rect 960 37348 1040 37360
rect 960 37292 972 37348
rect 1028 37292 1040 37348
rect 960 37028 1040 37292
rect 960 36972 972 37028
rect 1028 36972 1040 37028
rect 960 36960 1040 36972
rect 1120 37348 1200 37360
rect 1120 37292 1132 37348
rect 1188 37292 1200 37348
rect 1120 37028 1200 37292
rect 1120 36972 1132 37028
rect 1188 36972 1200 37028
rect 1120 36960 1200 36972
rect 1280 37348 1360 37360
rect 1280 37292 1292 37348
rect 1348 37292 1360 37348
rect 1280 37028 1360 37292
rect 1280 36972 1292 37028
rect 1348 36972 1360 37028
rect 1280 36960 1360 36972
rect 1440 37348 1520 37360
rect 1440 37292 1452 37348
rect 1508 37292 1520 37348
rect 1440 37028 1520 37292
rect 1440 36972 1452 37028
rect 1508 36972 1520 37028
rect 1440 36960 1520 36972
rect 1600 37348 1680 37360
rect 1600 37292 1612 37348
rect 1668 37292 1680 37348
rect 1600 37028 1680 37292
rect 1600 36972 1612 37028
rect 1668 36972 1680 37028
rect 1600 36960 1680 36972
rect 1760 37348 1840 37360
rect 1760 37292 1772 37348
rect 1828 37292 1840 37348
rect 1760 37028 1840 37292
rect 1760 36972 1772 37028
rect 1828 36972 1840 37028
rect 1760 36960 1840 36972
rect 1920 37348 2000 37360
rect 1920 37292 1932 37348
rect 1988 37292 2000 37348
rect 1920 37028 2000 37292
rect 1920 36972 1932 37028
rect 1988 36972 2000 37028
rect 1920 36960 2000 36972
rect 2080 37348 2160 37360
rect 2080 37292 2092 37348
rect 2148 37292 2160 37348
rect 2080 37028 2160 37292
rect 2080 36972 2092 37028
rect 2148 36972 2160 37028
rect 2080 36960 2160 36972
rect 2240 37348 2320 37360
rect 2240 37292 2252 37348
rect 2308 37292 2320 37348
rect 2240 37028 2320 37292
rect 2240 36972 2252 37028
rect 2308 36972 2320 37028
rect 2240 36960 2320 36972
rect 2400 37348 2480 37360
rect 2400 37292 2412 37348
rect 2468 37292 2480 37348
rect 2400 37028 2480 37292
rect 2400 36972 2412 37028
rect 2468 36972 2480 37028
rect 2400 36960 2480 36972
rect 2560 37348 2640 37360
rect 2560 37292 2572 37348
rect 2628 37292 2640 37348
rect 2560 37028 2640 37292
rect 2560 36972 2572 37028
rect 2628 36972 2640 37028
rect 2560 36960 2640 36972
rect 2720 37348 2800 37360
rect 2720 37292 2732 37348
rect 2788 37292 2800 37348
rect 2720 37028 2800 37292
rect 2720 36972 2732 37028
rect 2788 36972 2800 37028
rect 2720 36960 2800 36972
rect 2880 37348 2960 37360
rect 2880 37292 2892 37348
rect 2948 37292 2960 37348
rect 2880 37028 2960 37292
rect 2880 36972 2892 37028
rect 2948 36972 2960 37028
rect 2880 36960 2960 36972
rect 3040 37348 3120 37360
rect 3040 37292 3052 37348
rect 3108 37292 3120 37348
rect 3040 37028 3120 37292
rect 3040 36972 3052 37028
rect 3108 36972 3120 37028
rect 3040 36960 3120 36972
rect 3200 37348 3280 37360
rect 3200 37292 3212 37348
rect 3268 37292 3280 37348
rect 3200 37028 3280 37292
rect 3200 36972 3212 37028
rect 3268 36972 3280 37028
rect 3200 36960 3280 36972
rect 3360 37348 3440 37360
rect 3360 37292 3372 37348
rect 3428 37292 3440 37348
rect 3360 37028 3440 37292
rect 3360 36972 3372 37028
rect 3428 36972 3440 37028
rect 3360 36960 3440 36972
rect 3520 37348 3600 37360
rect 3520 37292 3532 37348
rect 3588 37292 3600 37348
rect 3520 37028 3600 37292
rect 3520 36972 3532 37028
rect 3588 36972 3600 37028
rect 3520 36960 3600 36972
rect 3680 37348 3760 37360
rect 3680 37292 3692 37348
rect 3748 37292 3760 37348
rect 3680 37028 3760 37292
rect 3680 36972 3692 37028
rect 3748 36972 3760 37028
rect 3680 36960 3760 36972
rect 3840 37348 3920 37360
rect 3840 37292 3852 37348
rect 3908 37292 3920 37348
rect 3840 37028 3920 37292
rect 3840 36972 3852 37028
rect 3908 36972 3920 37028
rect 3840 36960 3920 36972
rect 4000 37348 4080 37360
rect 4000 37292 4012 37348
rect 4068 37292 4080 37348
rect 4000 37028 4080 37292
rect 4000 36972 4012 37028
rect 4068 36972 4080 37028
rect 4000 36960 4080 36972
rect 4160 37348 4240 37360
rect 4160 37292 4172 37348
rect 4228 37292 4240 37348
rect 4160 37028 4240 37292
rect 4160 36972 4172 37028
rect 4228 36972 4240 37028
rect 4160 36960 4240 36972
rect 4320 37348 4400 37360
rect 4320 37292 4332 37348
rect 4388 37292 4400 37348
rect 4320 37028 4400 37292
rect 4320 36972 4332 37028
rect 4388 36972 4400 37028
rect 4320 36960 4400 36972
rect 4480 37348 4560 37360
rect 4480 37292 4492 37348
rect 4548 37292 4560 37348
rect 4480 37028 4560 37292
rect 4480 36972 4492 37028
rect 4548 36972 4560 37028
rect 4480 36960 4560 36972
rect 4640 37348 4720 37360
rect 4640 37292 4652 37348
rect 4708 37292 4720 37348
rect 4640 37028 4720 37292
rect 4640 36972 4652 37028
rect 4708 36972 4720 37028
rect 4640 36960 4720 36972
rect 4800 37348 4880 37360
rect 4800 37292 4812 37348
rect 4868 37292 4880 37348
rect 4800 37028 4880 37292
rect 4800 36972 4812 37028
rect 4868 36972 4880 37028
rect 4800 36960 4880 36972
rect 4960 37348 5040 37360
rect 4960 37292 4972 37348
rect 5028 37292 5040 37348
rect 4960 37028 5040 37292
rect 4960 36972 4972 37028
rect 5028 36972 5040 37028
rect 4960 36960 5040 36972
rect 5120 37348 5200 37360
rect 5120 37292 5132 37348
rect 5188 37292 5200 37348
rect 5120 37028 5200 37292
rect 5120 36972 5132 37028
rect 5188 36972 5200 37028
rect 5120 36960 5200 36972
rect 5280 37348 5360 37360
rect 5280 37292 5292 37348
rect 5348 37292 5360 37348
rect 5280 37028 5360 37292
rect 5280 36972 5292 37028
rect 5348 36972 5360 37028
rect 5280 36960 5360 36972
rect 5440 37348 5520 37360
rect 5440 37292 5452 37348
rect 5508 37292 5520 37348
rect 5440 37028 5520 37292
rect 5440 36972 5452 37028
rect 5508 36972 5520 37028
rect 5440 36960 5520 36972
rect 5600 37348 5680 37360
rect 5600 37292 5612 37348
rect 5668 37292 5680 37348
rect 5600 37028 5680 37292
rect 5600 36972 5612 37028
rect 5668 36972 5680 37028
rect 5600 36960 5680 36972
rect 5760 37348 5840 37360
rect 5760 37292 5772 37348
rect 5828 37292 5840 37348
rect 5760 37028 5840 37292
rect 5760 36972 5772 37028
rect 5828 36972 5840 37028
rect 5760 36960 5840 36972
rect 5920 37348 6000 37360
rect 5920 37292 5932 37348
rect 5988 37292 6000 37348
rect 5920 37028 6000 37292
rect 5920 36972 5932 37028
rect 5988 36972 6000 37028
rect 5920 36960 6000 36972
rect 6080 37348 6160 37360
rect 6080 37292 6092 37348
rect 6148 37292 6160 37348
rect 6080 37028 6160 37292
rect 6080 36972 6092 37028
rect 6148 36972 6160 37028
rect 6080 36960 6160 36972
rect 6240 37348 6320 37360
rect 6240 37292 6252 37348
rect 6308 37292 6320 37348
rect 6240 37028 6320 37292
rect 6240 36972 6252 37028
rect 6308 36972 6320 37028
rect 6240 36960 6320 36972
rect 6400 37348 6480 37360
rect 6400 37292 6412 37348
rect 6468 37292 6480 37348
rect 6400 37028 6480 37292
rect 6400 36972 6412 37028
rect 6468 36972 6480 37028
rect 6400 36960 6480 36972
rect 6560 37348 6640 37360
rect 6560 37292 6572 37348
rect 6628 37292 6640 37348
rect 6560 37028 6640 37292
rect 6560 36972 6572 37028
rect 6628 36972 6640 37028
rect 6560 36960 6640 36972
rect 6720 37348 6800 37360
rect 6720 37292 6732 37348
rect 6788 37292 6800 37348
rect 6720 37028 6800 37292
rect 6720 36972 6732 37028
rect 6788 36972 6800 37028
rect 6720 36960 6800 36972
rect 6880 37348 6960 37360
rect 6880 37292 6892 37348
rect 6948 37292 6960 37348
rect 6880 37028 6960 37292
rect 6880 36972 6892 37028
rect 6948 36972 6960 37028
rect 6880 36960 6960 36972
rect 7040 37348 7120 37360
rect 7040 37292 7052 37348
rect 7108 37292 7120 37348
rect 7040 37028 7120 37292
rect 7040 36972 7052 37028
rect 7108 36972 7120 37028
rect 7040 36960 7120 36972
rect 7200 37348 7280 37360
rect 7200 37292 7212 37348
rect 7268 37292 7280 37348
rect 7200 37028 7280 37292
rect 7200 36972 7212 37028
rect 7268 36972 7280 37028
rect 7200 36960 7280 36972
rect 7360 37348 7440 37360
rect 7360 37292 7372 37348
rect 7428 37292 7440 37348
rect 7360 37028 7440 37292
rect 7360 36972 7372 37028
rect 7428 36972 7440 37028
rect 7360 36960 7440 36972
rect 7520 37348 7600 37360
rect 7520 37292 7532 37348
rect 7588 37292 7600 37348
rect 7520 37028 7600 37292
rect 7520 36972 7532 37028
rect 7588 36972 7600 37028
rect 7520 36960 7600 36972
rect 7680 37348 7760 37360
rect 7680 37292 7692 37348
rect 7748 37292 7760 37348
rect 7680 37028 7760 37292
rect 7680 36972 7692 37028
rect 7748 36972 7760 37028
rect 7680 36960 7760 36972
rect 7840 37348 7920 37360
rect 7840 37292 7852 37348
rect 7908 37292 7920 37348
rect 7840 37028 7920 37292
rect 7840 36972 7852 37028
rect 7908 36972 7920 37028
rect 7840 36960 7920 36972
rect 8000 37348 8080 37360
rect 8000 37292 8012 37348
rect 8068 37292 8080 37348
rect 8000 37028 8080 37292
rect 8000 36972 8012 37028
rect 8068 36972 8080 37028
rect 8000 36960 8080 36972
rect 8160 37348 8240 37360
rect 8160 37292 8172 37348
rect 8228 37292 8240 37348
rect 8160 37028 8240 37292
rect 8160 36972 8172 37028
rect 8228 36972 8240 37028
rect 8160 36960 8240 36972
rect 8320 37348 8400 37360
rect 8320 37292 8332 37348
rect 8388 37292 8400 37348
rect 8320 37028 8400 37292
rect 8320 36972 8332 37028
rect 8388 36972 8400 37028
rect 8320 36960 8400 36972
rect 8480 37348 8560 37440
rect 8480 37292 8492 37348
rect 8548 37292 8560 37348
rect 8480 37028 8560 37292
rect 8480 36972 8492 37028
rect 8548 36972 8560 37028
rect 0 36868 80 36880
rect 0 36812 12 36868
rect 68 36812 80 36868
rect 0 36548 80 36812
rect 0 36492 12 36548
rect 68 36492 80 36548
rect 0 36480 80 36492
rect 160 36868 240 36880
rect 160 36812 172 36868
rect 228 36812 240 36868
rect 160 36548 240 36812
rect 160 36492 172 36548
rect 228 36492 240 36548
rect 160 36480 240 36492
rect 320 36868 400 36880
rect 320 36812 332 36868
rect 388 36812 400 36868
rect 320 36548 400 36812
rect 320 36492 332 36548
rect 388 36492 400 36548
rect 320 36480 400 36492
rect 480 36868 560 36880
rect 480 36812 492 36868
rect 548 36812 560 36868
rect 480 36548 560 36812
rect 480 36492 492 36548
rect 548 36492 560 36548
rect 480 36480 560 36492
rect 640 36868 720 36880
rect 640 36812 652 36868
rect 708 36812 720 36868
rect 640 36548 720 36812
rect 640 36492 652 36548
rect 708 36492 720 36548
rect 640 36480 720 36492
rect 800 36868 880 36880
rect 800 36812 812 36868
rect 868 36812 880 36868
rect 800 36548 880 36812
rect 800 36492 812 36548
rect 868 36492 880 36548
rect 800 36480 880 36492
rect 960 36868 1040 36880
rect 960 36812 972 36868
rect 1028 36812 1040 36868
rect 960 36548 1040 36812
rect 960 36492 972 36548
rect 1028 36492 1040 36548
rect 960 36480 1040 36492
rect 1120 36868 1200 36880
rect 1120 36812 1132 36868
rect 1188 36812 1200 36868
rect 1120 36548 1200 36812
rect 1120 36492 1132 36548
rect 1188 36492 1200 36548
rect 1120 36480 1200 36492
rect 1280 36868 1360 36880
rect 1280 36812 1292 36868
rect 1348 36812 1360 36868
rect 1280 36548 1360 36812
rect 1280 36492 1292 36548
rect 1348 36492 1360 36548
rect 1280 36480 1360 36492
rect 1440 36868 1520 36880
rect 1440 36812 1452 36868
rect 1508 36812 1520 36868
rect 1440 36548 1520 36812
rect 1440 36492 1452 36548
rect 1508 36492 1520 36548
rect 1440 36480 1520 36492
rect 1600 36868 1680 36880
rect 1600 36812 1612 36868
rect 1668 36812 1680 36868
rect 1600 36548 1680 36812
rect 1600 36492 1612 36548
rect 1668 36492 1680 36548
rect 1600 36480 1680 36492
rect 1760 36868 1840 36880
rect 1760 36812 1772 36868
rect 1828 36812 1840 36868
rect 1760 36548 1840 36812
rect 1760 36492 1772 36548
rect 1828 36492 1840 36548
rect 1760 36480 1840 36492
rect 1920 36868 2000 36880
rect 1920 36812 1932 36868
rect 1988 36812 2000 36868
rect 1920 36548 2000 36812
rect 1920 36492 1932 36548
rect 1988 36492 2000 36548
rect 1920 36480 2000 36492
rect 2080 36868 2160 36880
rect 2080 36812 2092 36868
rect 2148 36812 2160 36868
rect 2080 36548 2160 36812
rect 2080 36492 2092 36548
rect 2148 36492 2160 36548
rect 2080 36480 2160 36492
rect 2240 36868 2320 36880
rect 2240 36812 2252 36868
rect 2308 36812 2320 36868
rect 2240 36548 2320 36812
rect 2240 36492 2252 36548
rect 2308 36492 2320 36548
rect 2240 36480 2320 36492
rect 2400 36868 2480 36880
rect 2400 36812 2412 36868
rect 2468 36812 2480 36868
rect 2400 36548 2480 36812
rect 2400 36492 2412 36548
rect 2468 36492 2480 36548
rect 2400 36480 2480 36492
rect 2560 36868 2640 36880
rect 2560 36812 2572 36868
rect 2628 36812 2640 36868
rect 2560 36548 2640 36812
rect 2560 36492 2572 36548
rect 2628 36492 2640 36548
rect 2560 36480 2640 36492
rect 2720 36868 2800 36880
rect 2720 36812 2732 36868
rect 2788 36812 2800 36868
rect 2720 36548 2800 36812
rect 2720 36492 2732 36548
rect 2788 36492 2800 36548
rect 2720 36480 2800 36492
rect 2880 36868 2960 36880
rect 2880 36812 2892 36868
rect 2948 36812 2960 36868
rect 2880 36548 2960 36812
rect 2880 36492 2892 36548
rect 2948 36492 2960 36548
rect 2880 36480 2960 36492
rect 3040 36868 3120 36880
rect 3040 36812 3052 36868
rect 3108 36812 3120 36868
rect 3040 36548 3120 36812
rect 3040 36492 3052 36548
rect 3108 36492 3120 36548
rect 3040 36480 3120 36492
rect 3200 36868 3280 36880
rect 3200 36812 3212 36868
rect 3268 36812 3280 36868
rect 3200 36548 3280 36812
rect 3200 36492 3212 36548
rect 3268 36492 3280 36548
rect 3200 36480 3280 36492
rect 3360 36868 3440 36880
rect 3360 36812 3372 36868
rect 3428 36812 3440 36868
rect 3360 36548 3440 36812
rect 3360 36492 3372 36548
rect 3428 36492 3440 36548
rect 3360 36480 3440 36492
rect 3520 36868 3600 36880
rect 3520 36812 3532 36868
rect 3588 36812 3600 36868
rect 3520 36548 3600 36812
rect 3520 36492 3532 36548
rect 3588 36492 3600 36548
rect 3520 36480 3600 36492
rect 3680 36868 3760 36880
rect 3680 36812 3692 36868
rect 3748 36812 3760 36868
rect 3680 36548 3760 36812
rect 3680 36492 3692 36548
rect 3748 36492 3760 36548
rect 3680 36480 3760 36492
rect 3840 36868 3920 36880
rect 3840 36812 3852 36868
rect 3908 36812 3920 36868
rect 3840 36548 3920 36812
rect 3840 36492 3852 36548
rect 3908 36492 3920 36548
rect 3840 36480 3920 36492
rect 4000 36868 4080 36880
rect 4000 36812 4012 36868
rect 4068 36812 4080 36868
rect 4000 36548 4080 36812
rect 4000 36492 4012 36548
rect 4068 36492 4080 36548
rect 4000 36480 4080 36492
rect 4160 36868 4240 36880
rect 4160 36812 4172 36868
rect 4228 36812 4240 36868
rect 4160 36548 4240 36812
rect 4160 36492 4172 36548
rect 4228 36492 4240 36548
rect 4160 36480 4240 36492
rect 4320 36868 4400 36880
rect 4320 36812 4332 36868
rect 4388 36812 4400 36868
rect 4320 36548 4400 36812
rect 4320 36492 4332 36548
rect 4388 36492 4400 36548
rect 4320 36480 4400 36492
rect 4480 36868 4560 36880
rect 4480 36812 4492 36868
rect 4548 36812 4560 36868
rect 4480 36548 4560 36812
rect 4480 36492 4492 36548
rect 4548 36492 4560 36548
rect 4480 36480 4560 36492
rect 4640 36868 4720 36880
rect 4640 36812 4652 36868
rect 4708 36812 4720 36868
rect 4640 36548 4720 36812
rect 4640 36492 4652 36548
rect 4708 36492 4720 36548
rect 4640 36480 4720 36492
rect 4800 36868 4880 36880
rect 4800 36812 4812 36868
rect 4868 36812 4880 36868
rect 4800 36548 4880 36812
rect 4800 36492 4812 36548
rect 4868 36492 4880 36548
rect 4800 36480 4880 36492
rect 4960 36868 5040 36880
rect 4960 36812 4972 36868
rect 5028 36812 5040 36868
rect 4960 36548 5040 36812
rect 4960 36492 4972 36548
rect 5028 36492 5040 36548
rect 4960 36480 5040 36492
rect 5120 36868 5200 36880
rect 5120 36812 5132 36868
rect 5188 36812 5200 36868
rect 5120 36548 5200 36812
rect 5120 36492 5132 36548
rect 5188 36492 5200 36548
rect 5120 36480 5200 36492
rect 5280 36868 5360 36880
rect 5280 36812 5292 36868
rect 5348 36812 5360 36868
rect 5280 36548 5360 36812
rect 5280 36492 5292 36548
rect 5348 36492 5360 36548
rect 5280 36480 5360 36492
rect 5440 36868 5520 36880
rect 5440 36812 5452 36868
rect 5508 36812 5520 36868
rect 5440 36548 5520 36812
rect 5440 36492 5452 36548
rect 5508 36492 5520 36548
rect 5440 36480 5520 36492
rect 5600 36868 5680 36880
rect 5600 36812 5612 36868
rect 5668 36812 5680 36868
rect 5600 36548 5680 36812
rect 5600 36492 5612 36548
rect 5668 36492 5680 36548
rect 5600 36480 5680 36492
rect 5760 36868 5840 36880
rect 5760 36812 5772 36868
rect 5828 36812 5840 36868
rect 5760 36548 5840 36812
rect 5760 36492 5772 36548
rect 5828 36492 5840 36548
rect 5760 36480 5840 36492
rect 5920 36868 6000 36880
rect 5920 36812 5932 36868
rect 5988 36812 6000 36868
rect 5920 36548 6000 36812
rect 5920 36492 5932 36548
rect 5988 36492 6000 36548
rect 5920 36480 6000 36492
rect 6080 36868 6160 36880
rect 6080 36812 6092 36868
rect 6148 36812 6160 36868
rect 6080 36548 6160 36812
rect 6080 36492 6092 36548
rect 6148 36492 6160 36548
rect 6080 36480 6160 36492
rect 6240 36868 6320 36880
rect 6240 36812 6252 36868
rect 6308 36812 6320 36868
rect 6240 36548 6320 36812
rect 6240 36492 6252 36548
rect 6308 36492 6320 36548
rect 6240 36480 6320 36492
rect 6400 36868 6480 36880
rect 6400 36812 6412 36868
rect 6468 36812 6480 36868
rect 6400 36548 6480 36812
rect 6400 36492 6412 36548
rect 6468 36492 6480 36548
rect 6400 36480 6480 36492
rect 6560 36868 6640 36880
rect 6560 36812 6572 36868
rect 6628 36812 6640 36868
rect 6560 36548 6640 36812
rect 6560 36492 6572 36548
rect 6628 36492 6640 36548
rect 6560 36480 6640 36492
rect 6720 36868 6800 36880
rect 6720 36812 6732 36868
rect 6788 36812 6800 36868
rect 6720 36548 6800 36812
rect 6720 36492 6732 36548
rect 6788 36492 6800 36548
rect 6720 36480 6800 36492
rect 6880 36868 6960 36880
rect 6880 36812 6892 36868
rect 6948 36812 6960 36868
rect 6880 36548 6960 36812
rect 6880 36492 6892 36548
rect 6948 36492 6960 36548
rect 6880 36480 6960 36492
rect 7040 36868 7120 36880
rect 7040 36812 7052 36868
rect 7108 36812 7120 36868
rect 7040 36548 7120 36812
rect 7040 36492 7052 36548
rect 7108 36492 7120 36548
rect 7040 36480 7120 36492
rect 7200 36868 7280 36880
rect 7200 36812 7212 36868
rect 7268 36812 7280 36868
rect 7200 36548 7280 36812
rect 7200 36492 7212 36548
rect 7268 36492 7280 36548
rect 7200 36480 7280 36492
rect 7360 36868 7440 36880
rect 7360 36812 7372 36868
rect 7428 36812 7440 36868
rect 7360 36548 7440 36812
rect 7360 36492 7372 36548
rect 7428 36492 7440 36548
rect 7360 36480 7440 36492
rect 7520 36868 7600 36880
rect 7520 36812 7532 36868
rect 7588 36812 7600 36868
rect 7520 36548 7600 36812
rect 7520 36492 7532 36548
rect 7588 36492 7600 36548
rect 7520 36480 7600 36492
rect 7680 36868 7760 36880
rect 7680 36812 7692 36868
rect 7748 36812 7760 36868
rect 7680 36548 7760 36812
rect 7680 36492 7692 36548
rect 7748 36492 7760 36548
rect 7680 36480 7760 36492
rect 7840 36868 7920 36880
rect 7840 36812 7852 36868
rect 7908 36812 7920 36868
rect 7840 36548 7920 36812
rect 7840 36492 7852 36548
rect 7908 36492 7920 36548
rect 7840 36480 7920 36492
rect 8000 36868 8080 36880
rect 8000 36812 8012 36868
rect 8068 36812 8080 36868
rect 8000 36548 8080 36812
rect 8000 36492 8012 36548
rect 8068 36492 8080 36548
rect 8000 36480 8080 36492
rect 8160 36868 8240 36880
rect 8160 36812 8172 36868
rect 8228 36812 8240 36868
rect 8160 36548 8240 36812
rect 8160 36492 8172 36548
rect 8228 36492 8240 36548
rect 8160 36480 8240 36492
rect 8320 36868 8400 36880
rect 8320 36812 8332 36868
rect 8388 36812 8400 36868
rect 8320 36548 8400 36812
rect 8320 36492 8332 36548
rect 8388 36492 8400 36548
rect 8320 36480 8400 36492
rect 0 36388 80 36400
rect 0 36332 12 36388
rect 68 36332 80 36388
rect 0 36068 80 36332
rect 0 36012 12 36068
rect 68 36012 80 36068
rect 0 35748 80 36012
rect 0 35692 12 35748
rect 68 35692 80 35748
rect 0 35428 80 35692
rect 0 35372 12 35428
rect 68 35372 80 35428
rect 0 35108 80 35372
rect 0 35052 12 35108
rect 68 35052 80 35108
rect 0 34788 80 35052
rect 0 34732 12 34788
rect 68 34732 80 34788
rect 0 34468 80 34732
rect 0 34412 12 34468
rect 68 34412 80 34468
rect 0 34400 80 34412
rect 160 36388 240 36400
rect 160 36332 172 36388
rect 228 36332 240 36388
rect 160 36068 240 36332
rect 160 36012 172 36068
rect 228 36012 240 36068
rect 160 35748 240 36012
rect 160 35692 172 35748
rect 228 35692 240 35748
rect 160 35428 240 35692
rect 160 35372 172 35428
rect 228 35372 240 35428
rect 160 35108 240 35372
rect 160 35052 172 35108
rect 228 35052 240 35108
rect 160 34788 240 35052
rect 160 34732 172 34788
rect 228 34732 240 34788
rect 160 34468 240 34732
rect 160 34412 172 34468
rect 228 34412 240 34468
rect 160 34400 240 34412
rect 320 36388 400 36400
rect 320 36332 332 36388
rect 388 36332 400 36388
rect 320 36068 400 36332
rect 320 36012 332 36068
rect 388 36012 400 36068
rect 320 35748 400 36012
rect 320 35692 332 35748
rect 388 35692 400 35748
rect 320 35428 400 35692
rect 320 35372 332 35428
rect 388 35372 400 35428
rect 320 35108 400 35372
rect 320 35052 332 35108
rect 388 35052 400 35108
rect 320 34788 400 35052
rect 320 34732 332 34788
rect 388 34732 400 34788
rect 320 34468 400 34732
rect 320 34412 332 34468
rect 388 34412 400 34468
rect 320 34400 400 34412
rect 480 36388 560 36400
rect 480 36332 492 36388
rect 548 36332 560 36388
rect 480 36068 560 36332
rect 480 36012 492 36068
rect 548 36012 560 36068
rect 480 35748 560 36012
rect 480 35692 492 35748
rect 548 35692 560 35748
rect 480 35428 560 35692
rect 480 35372 492 35428
rect 548 35372 560 35428
rect 480 35108 560 35372
rect 480 35052 492 35108
rect 548 35052 560 35108
rect 480 34788 560 35052
rect 480 34732 492 34788
rect 548 34732 560 34788
rect 480 34468 560 34732
rect 480 34412 492 34468
rect 548 34412 560 34468
rect 480 34400 560 34412
rect 640 36388 720 36400
rect 640 36332 652 36388
rect 708 36332 720 36388
rect 640 36068 720 36332
rect 640 36012 652 36068
rect 708 36012 720 36068
rect 640 35748 720 36012
rect 640 35692 652 35748
rect 708 35692 720 35748
rect 640 35428 720 35692
rect 640 35372 652 35428
rect 708 35372 720 35428
rect 640 35108 720 35372
rect 640 35052 652 35108
rect 708 35052 720 35108
rect 640 34788 720 35052
rect 640 34732 652 34788
rect 708 34732 720 34788
rect 640 34468 720 34732
rect 640 34412 652 34468
rect 708 34412 720 34468
rect 640 34400 720 34412
rect 800 36388 880 36400
rect 800 36332 812 36388
rect 868 36332 880 36388
rect 800 36068 880 36332
rect 800 36012 812 36068
rect 868 36012 880 36068
rect 800 35748 880 36012
rect 800 35692 812 35748
rect 868 35692 880 35748
rect 800 35428 880 35692
rect 800 35372 812 35428
rect 868 35372 880 35428
rect 800 35108 880 35372
rect 800 35052 812 35108
rect 868 35052 880 35108
rect 800 34788 880 35052
rect 800 34732 812 34788
rect 868 34732 880 34788
rect 800 34468 880 34732
rect 800 34412 812 34468
rect 868 34412 880 34468
rect 800 34400 880 34412
rect 960 36388 1040 36400
rect 960 36332 972 36388
rect 1028 36332 1040 36388
rect 960 36068 1040 36332
rect 960 36012 972 36068
rect 1028 36012 1040 36068
rect 960 35748 1040 36012
rect 960 35692 972 35748
rect 1028 35692 1040 35748
rect 960 35428 1040 35692
rect 960 35372 972 35428
rect 1028 35372 1040 35428
rect 960 35108 1040 35372
rect 960 35052 972 35108
rect 1028 35052 1040 35108
rect 960 34788 1040 35052
rect 960 34732 972 34788
rect 1028 34732 1040 34788
rect 960 34468 1040 34732
rect 960 34412 972 34468
rect 1028 34412 1040 34468
rect 960 34400 1040 34412
rect 1120 36388 1200 36400
rect 1120 36332 1132 36388
rect 1188 36332 1200 36388
rect 1120 36068 1200 36332
rect 1120 36012 1132 36068
rect 1188 36012 1200 36068
rect 1120 35748 1200 36012
rect 1120 35692 1132 35748
rect 1188 35692 1200 35748
rect 1120 35428 1200 35692
rect 1120 35372 1132 35428
rect 1188 35372 1200 35428
rect 1120 35108 1200 35372
rect 1120 35052 1132 35108
rect 1188 35052 1200 35108
rect 1120 34788 1200 35052
rect 1120 34732 1132 34788
rect 1188 34732 1200 34788
rect 1120 34468 1200 34732
rect 1120 34412 1132 34468
rect 1188 34412 1200 34468
rect 1120 34400 1200 34412
rect 1280 36388 1360 36400
rect 1280 36332 1292 36388
rect 1348 36332 1360 36388
rect 1280 36068 1360 36332
rect 1280 36012 1292 36068
rect 1348 36012 1360 36068
rect 1280 35748 1360 36012
rect 1280 35692 1292 35748
rect 1348 35692 1360 35748
rect 1280 35428 1360 35692
rect 1280 35372 1292 35428
rect 1348 35372 1360 35428
rect 1280 35108 1360 35372
rect 1280 35052 1292 35108
rect 1348 35052 1360 35108
rect 1280 34788 1360 35052
rect 1280 34732 1292 34788
rect 1348 34732 1360 34788
rect 1280 34468 1360 34732
rect 1280 34412 1292 34468
rect 1348 34412 1360 34468
rect 1280 34400 1360 34412
rect 1440 36388 1520 36400
rect 1440 36332 1452 36388
rect 1508 36332 1520 36388
rect 1440 36068 1520 36332
rect 1440 36012 1452 36068
rect 1508 36012 1520 36068
rect 1440 35748 1520 36012
rect 1440 35692 1452 35748
rect 1508 35692 1520 35748
rect 1440 35428 1520 35692
rect 1440 35372 1452 35428
rect 1508 35372 1520 35428
rect 1440 35108 1520 35372
rect 1440 35052 1452 35108
rect 1508 35052 1520 35108
rect 1440 34788 1520 35052
rect 1440 34732 1452 34788
rect 1508 34732 1520 34788
rect 1440 34468 1520 34732
rect 1440 34412 1452 34468
rect 1508 34412 1520 34468
rect 1440 34400 1520 34412
rect 1600 36388 1680 36400
rect 1600 36332 1612 36388
rect 1668 36332 1680 36388
rect 1600 36068 1680 36332
rect 1600 36012 1612 36068
rect 1668 36012 1680 36068
rect 1600 35748 1680 36012
rect 1600 35692 1612 35748
rect 1668 35692 1680 35748
rect 1600 35428 1680 35692
rect 1600 35372 1612 35428
rect 1668 35372 1680 35428
rect 1600 35108 1680 35372
rect 1600 35052 1612 35108
rect 1668 35052 1680 35108
rect 1600 34788 1680 35052
rect 1600 34732 1612 34788
rect 1668 34732 1680 34788
rect 1600 34468 1680 34732
rect 1600 34412 1612 34468
rect 1668 34412 1680 34468
rect 1600 34400 1680 34412
rect 1760 36388 1840 36400
rect 1760 36332 1772 36388
rect 1828 36332 1840 36388
rect 1760 36068 1840 36332
rect 1760 36012 1772 36068
rect 1828 36012 1840 36068
rect 1760 35748 1840 36012
rect 1760 35692 1772 35748
rect 1828 35692 1840 35748
rect 1760 35428 1840 35692
rect 1760 35372 1772 35428
rect 1828 35372 1840 35428
rect 1760 35108 1840 35372
rect 1760 35052 1772 35108
rect 1828 35052 1840 35108
rect 1760 34788 1840 35052
rect 1760 34732 1772 34788
rect 1828 34732 1840 34788
rect 1760 34468 1840 34732
rect 1760 34412 1772 34468
rect 1828 34412 1840 34468
rect 1760 34400 1840 34412
rect 1920 36388 2000 36400
rect 1920 36332 1932 36388
rect 1988 36332 2000 36388
rect 1920 36068 2000 36332
rect 1920 36012 1932 36068
rect 1988 36012 2000 36068
rect 1920 35748 2000 36012
rect 1920 35692 1932 35748
rect 1988 35692 2000 35748
rect 1920 35428 2000 35692
rect 1920 35372 1932 35428
rect 1988 35372 2000 35428
rect 1920 35108 2000 35372
rect 1920 35052 1932 35108
rect 1988 35052 2000 35108
rect 1920 34788 2000 35052
rect 1920 34732 1932 34788
rect 1988 34732 2000 34788
rect 1920 34468 2000 34732
rect 1920 34412 1932 34468
rect 1988 34412 2000 34468
rect 1920 34400 2000 34412
rect 2080 36388 2160 36400
rect 2080 36332 2092 36388
rect 2148 36332 2160 36388
rect 2080 36068 2160 36332
rect 2080 36012 2092 36068
rect 2148 36012 2160 36068
rect 2080 35748 2160 36012
rect 2080 35692 2092 35748
rect 2148 35692 2160 35748
rect 2080 35428 2160 35692
rect 2080 35372 2092 35428
rect 2148 35372 2160 35428
rect 2080 35108 2160 35372
rect 2080 35052 2092 35108
rect 2148 35052 2160 35108
rect 2080 34788 2160 35052
rect 2080 34732 2092 34788
rect 2148 34732 2160 34788
rect 2080 34468 2160 34732
rect 2080 34412 2092 34468
rect 2148 34412 2160 34468
rect 2080 34400 2160 34412
rect 2240 36388 2320 36400
rect 2240 36332 2252 36388
rect 2308 36332 2320 36388
rect 2240 36068 2320 36332
rect 2240 36012 2252 36068
rect 2308 36012 2320 36068
rect 2240 35748 2320 36012
rect 2240 35692 2252 35748
rect 2308 35692 2320 35748
rect 2240 35428 2320 35692
rect 2240 35372 2252 35428
rect 2308 35372 2320 35428
rect 2240 35108 2320 35372
rect 2240 35052 2252 35108
rect 2308 35052 2320 35108
rect 2240 34788 2320 35052
rect 2240 34732 2252 34788
rect 2308 34732 2320 34788
rect 2240 34468 2320 34732
rect 2240 34412 2252 34468
rect 2308 34412 2320 34468
rect 2240 34400 2320 34412
rect 2400 36388 2480 36400
rect 2400 36332 2412 36388
rect 2468 36332 2480 36388
rect 2400 36068 2480 36332
rect 2400 36012 2412 36068
rect 2468 36012 2480 36068
rect 2400 35748 2480 36012
rect 2400 35692 2412 35748
rect 2468 35692 2480 35748
rect 2400 35428 2480 35692
rect 2400 35372 2412 35428
rect 2468 35372 2480 35428
rect 2400 35108 2480 35372
rect 2400 35052 2412 35108
rect 2468 35052 2480 35108
rect 2400 34788 2480 35052
rect 2400 34732 2412 34788
rect 2468 34732 2480 34788
rect 2400 34468 2480 34732
rect 2400 34412 2412 34468
rect 2468 34412 2480 34468
rect 2400 34400 2480 34412
rect 2560 36388 2640 36400
rect 2560 36332 2572 36388
rect 2628 36332 2640 36388
rect 2560 36068 2640 36332
rect 2560 36012 2572 36068
rect 2628 36012 2640 36068
rect 2560 35748 2640 36012
rect 2560 35692 2572 35748
rect 2628 35692 2640 35748
rect 2560 35428 2640 35692
rect 2560 35372 2572 35428
rect 2628 35372 2640 35428
rect 2560 35108 2640 35372
rect 2560 35052 2572 35108
rect 2628 35052 2640 35108
rect 2560 34788 2640 35052
rect 2560 34732 2572 34788
rect 2628 34732 2640 34788
rect 2560 34468 2640 34732
rect 2560 34412 2572 34468
rect 2628 34412 2640 34468
rect 2560 34400 2640 34412
rect 2720 36388 2800 36400
rect 2720 36332 2732 36388
rect 2788 36332 2800 36388
rect 2720 36068 2800 36332
rect 2720 36012 2732 36068
rect 2788 36012 2800 36068
rect 2720 35748 2800 36012
rect 2720 35692 2732 35748
rect 2788 35692 2800 35748
rect 2720 35428 2800 35692
rect 2720 35372 2732 35428
rect 2788 35372 2800 35428
rect 2720 35108 2800 35372
rect 2720 35052 2732 35108
rect 2788 35052 2800 35108
rect 2720 34788 2800 35052
rect 2720 34732 2732 34788
rect 2788 34732 2800 34788
rect 2720 34468 2800 34732
rect 2720 34412 2732 34468
rect 2788 34412 2800 34468
rect 2720 34400 2800 34412
rect 2880 36388 2960 36400
rect 2880 36332 2892 36388
rect 2948 36332 2960 36388
rect 2880 36068 2960 36332
rect 2880 36012 2892 36068
rect 2948 36012 2960 36068
rect 2880 35748 2960 36012
rect 2880 35692 2892 35748
rect 2948 35692 2960 35748
rect 2880 35428 2960 35692
rect 2880 35372 2892 35428
rect 2948 35372 2960 35428
rect 2880 35108 2960 35372
rect 2880 35052 2892 35108
rect 2948 35052 2960 35108
rect 2880 34788 2960 35052
rect 2880 34732 2892 34788
rect 2948 34732 2960 34788
rect 2880 34468 2960 34732
rect 2880 34412 2892 34468
rect 2948 34412 2960 34468
rect 2880 34400 2960 34412
rect 3040 36388 3120 36400
rect 3040 36332 3052 36388
rect 3108 36332 3120 36388
rect 3040 36068 3120 36332
rect 3040 36012 3052 36068
rect 3108 36012 3120 36068
rect 3040 35748 3120 36012
rect 3040 35692 3052 35748
rect 3108 35692 3120 35748
rect 3040 35428 3120 35692
rect 3040 35372 3052 35428
rect 3108 35372 3120 35428
rect 3040 35108 3120 35372
rect 3040 35052 3052 35108
rect 3108 35052 3120 35108
rect 3040 34788 3120 35052
rect 3040 34732 3052 34788
rect 3108 34732 3120 34788
rect 3040 34468 3120 34732
rect 3040 34412 3052 34468
rect 3108 34412 3120 34468
rect 3040 34400 3120 34412
rect 3200 36388 3280 36400
rect 3200 36332 3212 36388
rect 3268 36332 3280 36388
rect 3200 36068 3280 36332
rect 3200 36012 3212 36068
rect 3268 36012 3280 36068
rect 3200 35748 3280 36012
rect 3200 35692 3212 35748
rect 3268 35692 3280 35748
rect 3200 35428 3280 35692
rect 3200 35372 3212 35428
rect 3268 35372 3280 35428
rect 3200 35108 3280 35372
rect 3200 35052 3212 35108
rect 3268 35052 3280 35108
rect 3200 34788 3280 35052
rect 3200 34732 3212 34788
rect 3268 34732 3280 34788
rect 3200 34468 3280 34732
rect 3200 34412 3212 34468
rect 3268 34412 3280 34468
rect 3200 34400 3280 34412
rect 3360 36388 3440 36400
rect 3360 36332 3372 36388
rect 3428 36332 3440 36388
rect 3360 36068 3440 36332
rect 3360 36012 3372 36068
rect 3428 36012 3440 36068
rect 3360 35748 3440 36012
rect 3360 35692 3372 35748
rect 3428 35692 3440 35748
rect 3360 35428 3440 35692
rect 3360 35372 3372 35428
rect 3428 35372 3440 35428
rect 3360 35108 3440 35372
rect 3360 35052 3372 35108
rect 3428 35052 3440 35108
rect 3360 34788 3440 35052
rect 3360 34732 3372 34788
rect 3428 34732 3440 34788
rect 3360 34468 3440 34732
rect 3360 34412 3372 34468
rect 3428 34412 3440 34468
rect 3360 34400 3440 34412
rect 3520 36388 3600 36400
rect 3520 36332 3532 36388
rect 3588 36332 3600 36388
rect 3520 36068 3600 36332
rect 3520 36012 3532 36068
rect 3588 36012 3600 36068
rect 3520 35748 3600 36012
rect 3520 35692 3532 35748
rect 3588 35692 3600 35748
rect 3520 35428 3600 35692
rect 3520 35372 3532 35428
rect 3588 35372 3600 35428
rect 3520 35108 3600 35372
rect 3520 35052 3532 35108
rect 3588 35052 3600 35108
rect 3520 34788 3600 35052
rect 3520 34732 3532 34788
rect 3588 34732 3600 34788
rect 3520 34468 3600 34732
rect 3520 34412 3532 34468
rect 3588 34412 3600 34468
rect 3520 34400 3600 34412
rect 3680 36388 3760 36400
rect 3680 36332 3692 36388
rect 3748 36332 3760 36388
rect 3680 36068 3760 36332
rect 3680 36012 3692 36068
rect 3748 36012 3760 36068
rect 3680 35748 3760 36012
rect 3680 35692 3692 35748
rect 3748 35692 3760 35748
rect 3680 35428 3760 35692
rect 3680 35372 3692 35428
rect 3748 35372 3760 35428
rect 3680 35108 3760 35372
rect 3680 35052 3692 35108
rect 3748 35052 3760 35108
rect 3680 34788 3760 35052
rect 3680 34732 3692 34788
rect 3748 34732 3760 34788
rect 3680 34468 3760 34732
rect 3680 34412 3692 34468
rect 3748 34412 3760 34468
rect 3680 34400 3760 34412
rect 3840 36388 3920 36400
rect 3840 36332 3852 36388
rect 3908 36332 3920 36388
rect 3840 36068 3920 36332
rect 3840 36012 3852 36068
rect 3908 36012 3920 36068
rect 3840 35748 3920 36012
rect 3840 35692 3852 35748
rect 3908 35692 3920 35748
rect 3840 35428 3920 35692
rect 3840 35372 3852 35428
rect 3908 35372 3920 35428
rect 3840 35108 3920 35372
rect 3840 35052 3852 35108
rect 3908 35052 3920 35108
rect 3840 34788 3920 35052
rect 3840 34732 3852 34788
rect 3908 34732 3920 34788
rect 3840 34468 3920 34732
rect 3840 34412 3852 34468
rect 3908 34412 3920 34468
rect 3840 34400 3920 34412
rect 4000 36388 4080 36400
rect 4000 36332 4012 36388
rect 4068 36332 4080 36388
rect 4000 36068 4080 36332
rect 4000 36012 4012 36068
rect 4068 36012 4080 36068
rect 4000 35748 4080 36012
rect 4000 35692 4012 35748
rect 4068 35692 4080 35748
rect 4000 35428 4080 35692
rect 4000 35372 4012 35428
rect 4068 35372 4080 35428
rect 4000 35108 4080 35372
rect 4000 35052 4012 35108
rect 4068 35052 4080 35108
rect 4000 34788 4080 35052
rect 4000 34732 4012 34788
rect 4068 34732 4080 34788
rect 4000 34468 4080 34732
rect 4000 34412 4012 34468
rect 4068 34412 4080 34468
rect 4000 34400 4080 34412
rect 4160 36388 4240 36400
rect 4160 36332 4172 36388
rect 4228 36332 4240 36388
rect 4160 36068 4240 36332
rect 4160 36012 4172 36068
rect 4228 36012 4240 36068
rect 4160 35748 4240 36012
rect 4160 35692 4172 35748
rect 4228 35692 4240 35748
rect 4160 35428 4240 35692
rect 4160 35372 4172 35428
rect 4228 35372 4240 35428
rect 4160 35108 4240 35372
rect 4160 35052 4172 35108
rect 4228 35052 4240 35108
rect 4160 34788 4240 35052
rect 4160 34732 4172 34788
rect 4228 34732 4240 34788
rect 4160 34468 4240 34732
rect 4160 34412 4172 34468
rect 4228 34412 4240 34468
rect 4160 34400 4240 34412
rect 4320 36388 4400 36400
rect 4320 36332 4332 36388
rect 4388 36332 4400 36388
rect 4320 36068 4400 36332
rect 4320 36012 4332 36068
rect 4388 36012 4400 36068
rect 4320 35748 4400 36012
rect 4320 35692 4332 35748
rect 4388 35692 4400 35748
rect 4320 35428 4400 35692
rect 4320 35372 4332 35428
rect 4388 35372 4400 35428
rect 4320 35108 4400 35372
rect 4320 35052 4332 35108
rect 4388 35052 4400 35108
rect 4320 34788 4400 35052
rect 4320 34732 4332 34788
rect 4388 34732 4400 34788
rect 4320 34468 4400 34732
rect 4320 34412 4332 34468
rect 4388 34412 4400 34468
rect 4320 34400 4400 34412
rect 4480 36388 4560 36400
rect 4480 36332 4492 36388
rect 4548 36332 4560 36388
rect 4480 36068 4560 36332
rect 4480 36012 4492 36068
rect 4548 36012 4560 36068
rect 4480 35748 4560 36012
rect 4480 35692 4492 35748
rect 4548 35692 4560 35748
rect 4480 35428 4560 35692
rect 4480 35372 4492 35428
rect 4548 35372 4560 35428
rect 4480 35108 4560 35372
rect 4480 35052 4492 35108
rect 4548 35052 4560 35108
rect 4480 34788 4560 35052
rect 4480 34732 4492 34788
rect 4548 34732 4560 34788
rect 4480 34468 4560 34732
rect 4480 34412 4492 34468
rect 4548 34412 4560 34468
rect 4480 34400 4560 34412
rect 4640 36388 4720 36400
rect 4640 36332 4652 36388
rect 4708 36332 4720 36388
rect 4640 36068 4720 36332
rect 4640 36012 4652 36068
rect 4708 36012 4720 36068
rect 4640 35748 4720 36012
rect 4640 35692 4652 35748
rect 4708 35692 4720 35748
rect 4640 35428 4720 35692
rect 4640 35372 4652 35428
rect 4708 35372 4720 35428
rect 4640 35108 4720 35372
rect 4640 35052 4652 35108
rect 4708 35052 4720 35108
rect 4640 34788 4720 35052
rect 4640 34732 4652 34788
rect 4708 34732 4720 34788
rect 4640 34468 4720 34732
rect 4640 34412 4652 34468
rect 4708 34412 4720 34468
rect 4640 34400 4720 34412
rect 4800 36388 4880 36400
rect 4800 36332 4812 36388
rect 4868 36332 4880 36388
rect 4800 36068 4880 36332
rect 4800 36012 4812 36068
rect 4868 36012 4880 36068
rect 4800 35748 4880 36012
rect 4800 35692 4812 35748
rect 4868 35692 4880 35748
rect 4800 35428 4880 35692
rect 4800 35372 4812 35428
rect 4868 35372 4880 35428
rect 4800 35108 4880 35372
rect 4800 35052 4812 35108
rect 4868 35052 4880 35108
rect 4800 34788 4880 35052
rect 4800 34732 4812 34788
rect 4868 34732 4880 34788
rect 4800 34468 4880 34732
rect 4800 34412 4812 34468
rect 4868 34412 4880 34468
rect 4800 34400 4880 34412
rect 4960 36388 5040 36400
rect 4960 36332 4972 36388
rect 5028 36332 5040 36388
rect 4960 36068 5040 36332
rect 4960 36012 4972 36068
rect 5028 36012 5040 36068
rect 4960 35748 5040 36012
rect 4960 35692 4972 35748
rect 5028 35692 5040 35748
rect 4960 35428 5040 35692
rect 4960 35372 4972 35428
rect 5028 35372 5040 35428
rect 4960 35108 5040 35372
rect 4960 35052 4972 35108
rect 5028 35052 5040 35108
rect 4960 34788 5040 35052
rect 4960 34732 4972 34788
rect 5028 34732 5040 34788
rect 4960 34468 5040 34732
rect 4960 34412 4972 34468
rect 5028 34412 5040 34468
rect 4960 34400 5040 34412
rect 5120 36388 5200 36400
rect 5120 36332 5132 36388
rect 5188 36332 5200 36388
rect 5120 36068 5200 36332
rect 5120 36012 5132 36068
rect 5188 36012 5200 36068
rect 5120 35748 5200 36012
rect 5120 35692 5132 35748
rect 5188 35692 5200 35748
rect 5120 35428 5200 35692
rect 5120 35372 5132 35428
rect 5188 35372 5200 35428
rect 5120 35108 5200 35372
rect 5120 35052 5132 35108
rect 5188 35052 5200 35108
rect 5120 34788 5200 35052
rect 5120 34732 5132 34788
rect 5188 34732 5200 34788
rect 5120 34468 5200 34732
rect 5120 34412 5132 34468
rect 5188 34412 5200 34468
rect 5120 34400 5200 34412
rect 5280 36388 5360 36400
rect 5280 36332 5292 36388
rect 5348 36332 5360 36388
rect 5280 36068 5360 36332
rect 5280 36012 5292 36068
rect 5348 36012 5360 36068
rect 5280 35748 5360 36012
rect 5280 35692 5292 35748
rect 5348 35692 5360 35748
rect 5280 35428 5360 35692
rect 5280 35372 5292 35428
rect 5348 35372 5360 35428
rect 5280 35108 5360 35372
rect 5280 35052 5292 35108
rect 5348 35052 5360 35108
rect 5280 34788 5360 35052
rect 5280 34732 5292 34788
rect 5348 34732 5360 34788
rect 5280 34468 5360 34732
rect 5280 34412 5292 34468
rect 5348 34412 5360 34468
rect 5280 34400 5360 34412
rect 5440 36388 5520 36400
rect 5440 36332 5452 36388
rect 5508 36332 5520 36388
rect 5440 36068 5520 36332
rect 5440 36012 5452 36068
rect 5508 36012 5520 36068
rect 5440 35748 5520 36012
rect 5440 35692 5452 35748
rect 5508 35692 5520 35748
rect 5440 35428 5520 35692
rect 5440 35372 5452 35428
rect 5508 35372 5520 35428
rect 5440 35108 5520 35372
rect 5440 35052 5452 35108
rect 5508 35052 5520 35108
rect 5440 34788 5520 35052
rect 5440 34732 5452 34788
rect 5508 34732 5520 34788
rect 5440 34468 5520 34732
rect 5440 34412 5452 34468
rect 5508 34412 5520 34468
rect 5440 34400 5520 34412
rect 5600 36388 5680 36400
rect 5600 36332 5612 36388
rect 5668 36332 5680 36388
rect 5600 36068 5680 36332
rect 5600 36012 5612 36068
rect 5668 36012 5680 36068
rect 5600 35748 5680 36012
rect 5600 35692 5612 35748
rect 5668 35692 5680 35748
rect 5600 35428 5680 35692
rect 5600 35372 5612 35428
rect 5668 35372 5680 35428
rect 5600 35108 5680 35372
rect 5600 35052 5612 35108
rect 5668 35052 5680 35108
rect 5600 34788 5680 35052
rect 5600 34732 5612 34788
rect 5668 34732 5680 34788
rect 5600 34468 5680 34732
rect 5600 34412 5612 34468
rect 5668 34412 5680 34468
rect 5600 34400 5680 34412
rect 5760 36388 5840 36400
rect 5760 36332 5772 36388
rect 5828 36332 5840 36388
rect 5760 36068 5840 36332
rect 5760 36012 5772 36068
rect 5828 36012 5840 36068
rect 5760 35748 5840 36012
rect 5760 35692 5772 35748
rect 5828 35692 5840 35748
rect 5760 35428 5840 35692
rect 5760 35372 5772 35428
rect 5828 35372 5840 35428
rect 5760 35108 5840 35372
rect 5760 35052 5772 35108
rect 5828 35052 5840 35108
rect 5760 34788 5840 35052
rect 5760 34732 5772 34788
rect 5828 34732 5840 34788
rect 5760 34468 5840 34732
rect 5760 34412 5772 34468
rect 5828 34412 5840 34468
rect 5760 34400 5840 34412
rect 5920 36388 6000 36400
rect 5920 36332 5932 36388
rect 5988 36332 6000 36388
rect 5920 36068 6000 36332
rect 5920 36012 5932 36068
rect 5988 36012 6000 36068
rect 5920 35748 6000 36012
rect 5920 35692 5932 35748
rect 5988 35692 6000 35748
rect 5920 35428 6000 35692
rect 5920 35372 5932 35428
rect 5988 35372 6000 35428
rect 5920 35108 6000 35372
rect 5920 35052 5932 35108
rect 5988 35052 6000 35108
rect 5920 34788 6000 35052
rect 5920 34732 5932 34788
rect 5988 34732 6000 34788
rect 5920 34468 6000 34732
rect 5920 34412 5932 34468
rect 5988 34412 6000 34468
rect 5920 34400 6000 34412
rect 6080 36388 6160 36400
rect 6080 36332 6092 36388
rect 6148 36332 6160 36388
rect 6080 36068 6160 36332
rect 6080 36012 6092 36068
rect 6148 36012 6160 36068
rect 6080 35748 6160 36012
rect 6080 35692 6092 35748
rect 6148 35692 6160 35748
rect 6080 35428 6160 35692
rect 6080 35372 6092 35428
rect 6148 35372 6160 35428
rect 6080 35108 6160 35372
rect 6080 35052 6092 35108
rect 6148 35052 6160 35108
rect 6080 34788 6160 35052
rect 6080 34732 6092 34788
rect 6148 34732 6160 34788
rect 6080 34468 6160 34732
rect 6080 34412 6092 34468
rect 6148 34412 6160 34468
rect 6080 34400 6160 34412
rect 6240 36388 6320 36400
rect 6240 36332 6252 36388
rect 6308 36332 6320 36388
rect 6240 36068 6320 36332
rect 6240 36012 6252 36068
rect 6308 36012 6320 36068
rect 6240 35748 6320 36012
rect 6240 35692 6252 35748
rect 6308 35692 6320 35748
rect 6240 35428 6320 35692
rect 6240 35372 6252 35428
rect 6308 35372 6320 35428
rect 6240 35108 6320 35372
rect 6240 35052 6252 35108
rect 6308 35052 6320 35108
rect 6240 34788 6320 35052
rect 6240 34732 6252 34788
rect 6308 34732 6320 34788
rect 6240 34468 6320 34732
rect 6240 34412 6252 34468
rect 6308 34412 6320 34468
rect 6240 34400 6320 34412
rect 6400 36388 6480 36400
rect 6400 36332 6412 36388
rect 6468 36332 6480 36388
rect 6400 36068 6480 36332
rect 6400 36012 6412 36068
rect 6468 36012 6480 36068
rect 6400 35748 6480 36012
rect 6400 35692 6412 35748
rect 6468 35692 6480 35748
rect 6400 35428 6480 35692
rect 6400 35372 6412 35428
rect 6468 35372 6480 35428
rect 6400 35108 6480 35372
rect 6400 35052 6412 35108
rect 6468 35052 6480 35108
rect 6400 34788 6480 35052
rect 6400 34732 6412 34788
rect 6468 34732 6480 34788
rect 6400 34468 6480 34732
rect 6400 34412 6412 34468
rect 6468 34412 6480 34468
rect 6400 34400 6480 34412
rect 6560 36388 6640 36400
rect 6560 36332 6572 36388
rect 6628 36332 6640 36388
rect 6560 36068 6640 36332
rect 6560 36012 6572 36068
rect 6628 36012 6640 36068
rect 6560 35748 6640 36012
rect 6560 35692 6572 35748
rect 6628 35692 6640 35748
rect 6560 35428 6640 35692
rect 6560 35372 6572 35428
rect 6628 35372 6640 35428
rect 6560 35108 6640 35372
rect 6560 35052 6572 35108
rect 6628 35052 6640 35108
rect 6560 34788 6640 35052
rect 6560 34732 6572 34788
rect 6628 34732 6640 34788
rect 6560 34468 6640 34732
rect 6560 34412 6572 34468
rect 6628 34412 6640 34468
rect 6560 34400 6640 34412
rect 6720 36388 6800 36400
rect 6720 36332 6732 36388
rect 6788 36332 6800 36388
rect 6720 36068 6800 36332
rect 6720 36012 6732 36068
rect 6788 36012 6800 36068
rect 6720 35748 6800 36012
rect 6720 35692 6732 35748
rect 6788 35692 6800 35748
rect 6720 35428 6800 35692
rect 6720 35372 6732 35428
rect 6788 35372 6800 35428
rect 6720 35108 6800 35372
rect 6720 35052 6732 35108
rect 6788 35052 6800 35108
rect 6720 34788 6800 35052
rect 6720 34732 6732 34788
rect 6788 34732 6800 34788
rect 6720 34468 6800 34732
rect 6720 34412 6732 34468
rect 6788 34412 6800 34468
rect 6720 34400 6800 34412
rect 6880 36388 6960 36400
rect 6880 36332 6892 36388
rect 6948 36332 6960 36388
rect 6880 36068 6960 36332
rect 6880 36012 6892 36068
rect 6948 36012 6960 36068
rect 6880 35748 6960 36012
rect 6880 35692 6892 35748
rect 6948 35692 6960 35748
rect 6880 35428 6960 35692
rect 6880 35372 6892 35428
rect 6948 35372 6960 35428
rect 6880 35108 6960 35372
rect 6880 35052 6892 35108
rect 6948 35052 6960 35108
rect 6880 34788 6960 35052
rect 6880 34732 6892 34788
rect 6948 34732 6960 34788
rect 6880 34468 6960 34732
rect 6880 34412 6892 34468
rect 6948 34412 6960 34468
rect 6880 34400 6960 34412
rect 7040 36388 7120 36400
rect 7040 36332 7052 36388
rect 7108 36332 7120 36388
rect 7040 36068 7120 36332
rect 7040 36012 7052 36068
rect 7108 36012 7120 36068
rect 7040 35748 7120 36012
rect 7040 35692 7052 35748
rect 7108 35692 7120 35748
rect 7040 35428 7120 35692
rect 7040 35372 7052 35428
rect 7108 35372 7120 35428
rect 7040 35108 7120 35372
rect 7040 35052 7052 35108
rect 7108 35052 7120 35108
rect 7040 34788 7120 35052
rect 7040 34732 7052 34788
rect 7108 34732 7120 34788
rect 7040 34468 7120 34732
rect 7040 34412 7052 34468
rect 7108 34412 7120 34468
rect 7040 34400 7120 34412
rect 7200 36388 7280 36400
rect 7200 36332 7212 36388
rect 7268 36332 7280 36388
rect 7200 36068 7280 36332
rect 7200 36012 7212 36068
rect 7268 36012 7280 36068
rect 7200 35748 7280 36012
rect 7200 35692 7212 35748
rect 7268 35692 7280 35748
rect 7200 35428 7280 35692
rect 7200 35372 7212 35428
rect 7268 35372 7280 35428
rect 7200 35108 7280 35372
rect 7200 35052 7212 35108
rect 7268 35052 7280 35108
rect 7200 34788 7280 35052
rect 7200 34732 7212 34788
rect 7268 34732 7280 34788
rect 7200 34468 7280 34732
rect 7200 34412 7212 34468
rect 7268 34412 7280 34468
rect 7200 34400 7280 34412
rect 7360 36388 7440 36400
rect 7360 36332 7372 36388
rect 7428 36332 7440 36388
rect 7360 36068 7440 36332
rect 7360 36012 7372 36068
rect 7428 36012 7440 36068
rect 7360 35748 7440 36012
rect 7360 35692 7372 35748
rect 7428 35692 7440 35748
rect 7360 35428 7440 35692
rect 7360 35372 7372 35428
rect 7428 35372 7440 35428
rect 7360 35108 7440 35372
rect 7360 35052 7372 35108
rect 7428 35052 7440 35108
rect 7360 34788 7440 35052
rect 7360 34732 7372 34788
rect 7428 34732 7440 34788
rect 7360 34468 7440 34732
rect 7360 34412 7372 34468
rect 7428 34412 7440 34468
rect 7360 34400 7440 34412
rect 7520 36388 7600 36400
rect 7520 36332 7532 36388
rect 7588 36332 7600 36388
rect 7520 36068 7600 36332
rect 7520 36012 7532 36068
rect 7588 36012 7600 36068
rect 7520 35748 7600 36012
rect 7520 35692 7532 35748
rect 7588 35692 7600 35748
rect 7520 35428 7600 35692
rect 7520 35372 7532 35428
rect 7588 35372 7600 35428
rect 7520 35108 7600 35372
rect 7520 35052 7532 35108
rect 7588 35052 7600 35108
rect 7520 34788 7600 35052
rect 7520 34732 7532 34788
rect 7588 34732 7600 34788
rect 7520 34468 7600 34732
rect 7520 34412 7532 34468
rect 7588 34412 7600 34468
rect 7520 34400 7600 34412
rect 7680 36388 7760 36400
rect 7680 36332 7692 36388
rect 7748 36332 7760 36388
rect 7680 36068 7760 36332
rect 7680 36012 7692 36068
rect 7748 36012 7760 36068
rect 7680 35748 7760 36012
rect 7680 35692 7692 35748
rect 7748 35692 7760 35748
rect 7680 35428 7760 35692
rect 7680 35372 7692 35428
rect 7748 35372 7760 35428
rect 7680 35108 7760 35372
rect 7680 35052 7692 35108
rect 7748 35052 7760 35108
rect 7680 34788 7760 35052
rect 7680 34732 7692 34788
rect 7748 34732 7760 34788
rect 7680 34468 7760 34732
rect 7680 34412 7692 34468
rect 7748 34412 7760 34468
rect 7680 34400 7760 34412
rect 7840 36388 7920 36400
rect 7840 36332 7852 36388
rect 7908 36332 7920 36388
rect 7840 36068 7920 36332
rect 7840 36012 7852 36068
rect 7908 36012 7920 36068
rect 7840 35748 7920 36012
rect 7840 35692 7852 35748
rect 7908 35692 7920 35748
rect 7840 35428 7920 35692
rect 7840 35372 7852 35428
rect 7908 35372 7920 35428
rect 7840 35108 7920 35372
rect 7840 35052 7852 35108
rect 7908 35052 7920 35108
rect 7840 34788 7920 35052
rect 7840 34732 7852 34788
rect 7908 34732 7920 34788
rect 7840 34468 7920 34732
rect 7840 34412 7852 34468
rect 7908 34412 7920 34468
rect 7840 34400 7920 34412
rect 8000 36388 8080 36400
rect 8000 36332 8012 36388
rect 8068 36332 8080 36388
rect 8000 36068 8080 36332
rect 8000 36012 8012 36068
rect 8068 36012 8080 36068
rect 8000 35748 8080 36012
rect 8000 35692 8012 35748
rect 8068 35692 8080 35748
rect 8000 35428 8080 35692
rect 8000 35372 8012 35428
rect 8068 35372 8080 35428
rect 8000 35108 8080 35372
rect 8000 35052 8012 35108
rect 8068 35052 8080 35108
rect 8000 34788 8080 35052
rect 8000 34732 8012 34788
rect 8068 34732 8080 34788
rect 8000 34468 8080 34732
rect 8000 34412 8012 34468
rect 8068 34412 8080 34468
rect 8000 34400 8080 34412
rect 8160 36388 8240 36400
rect 8160 36332 8172 36388
rect 8228 36332 8240 36388
rect 8160 36068 8240 36332
rect 8160 36012 8172 36068
rect 8228 36012 8240 36068
rect 8160 35748 8240 36012
rect 8160 35692 8172 35748
rect 8228 35692 8240 35748
rect 8160 35428 8240 35692
rect 8160 35372 8172 35428
rect 8228 35372 8240 35428
rect 8160 35108 8240 35372
rect 8160 35052 8172 35108
rect 8228 35052 8240 35108
rect 8160 34788 8240 35052
rect 8160 34732 8172 34788
rect 8228 34732 8240 34788
rect 8160 34468 8240 34732
rect 8160 34412 8172 34468
rect 8228 34412 8240 34468
rect 8160 34400 8240 34412
rect 8320 36388 8400 36400
rect 8320 36332 8332 36388
rect 8388 36332 8400 36388
rect 8320 36068 8400 36332
rect 8320 36012 8332 36068
rect 8388 36012 8400 36068
rect 8320 35748 8400 36012
rect 8320 35692 8332 35748
rect 8388 35692 8400 35748
rect 8320 35428 8400 35692
rect 8320 35372 8332 35428
rect 8388 35372 8400 35428
rect 8320 35108 8400 35372
rect 8320 35052 8332 35108
rect 8388 35052 8400 35108
rect 8320 34788 8400 35052
rect 8320 34732 8332 34788
rect 8388 34732 8400 34788
rect 8320 34468 8400 34732
rect 8320 34412 8332 34468
rect 8388 34412 8400 34468
rect 8320 34400 8400 34412
rect 0 34308 80 34320
rect 0 34252 12 34308
rect 68 34252 80 34308
rect 0 33988 80 34252
rect 0 33932 12 33988
rect 68 33932 80 33988
rect 0 33920 80 33932
rect 160 34308 240 34320
rect 160 34252 172 34308
rect 228 34252 240 34308
rect 160 33988 240 34252
rect 160 33932 172 33988
rect 228 33932 240 33988
rect 160 33920 240 33932
rect 320 34308 400 34320
rect 320 34252 332 34308
rect 388 34252 400 34308
rect 320 33988 400 34252
rect 320 33932 332 33988
rect 388 33932 400 33988
rect 320 33920 400 33932
rect 480 34308 560 34320
rect 480 34252 492 34308
rect 548 34252 560 34308
rect 480 33988 560 34252
rect 480 33932 492 33988
rect 548 33932 560 33988
rect 480 33920 560 33932
rect 640 34308 720 34320
rect 640 34252 652 34308
rect 708 34252 720 34308
rect 640 33988 720 34252
rect 640 33932 652 33988
rect 708 33932 720 33988
rect 640 33920 720 33932
rect 800 34308 880 34320
rect 800 34252 812 34308
rect 868 34252 880 34308
rect 800 33988 880 34252
rect 800 33932 812 33988
rect 868 33932 880 33988
rect 800 33920 880 33932
rect 960 34308 1040 34320
rect 960 34252 972 34308
rect 1028 34252 1040 34308
rect 960 33988 1040 34252
rect 960 33932 972 33988
rect 1028 33932 1040 33988
rect 960 33920 1040 33932
rect 1120 34308 1200 34320
rect 1120 34252 1132 34308
rect 1188 34252 1200 34308
rect 1120 33988 1200 34252
rect 1120 33932 1132 33988
rect 1188 33932 1200 33988
rect 1120 33920 1200 33932
rect 1280 34308 1360 34320
rect 1280 34252 1292 34308
rect 1348 34252 1360 34308
rect 1280 33988 1360 34252
rect 1280 33932 1292 33988
rect 1348 33932 1360 33988
rect 1280 33920 1360 33932
rect 1440 34308 1520 34320
rect 1440 34252 1452 34308
rect 1508 34252 1520 34308
rect 1440 33988 1520 34252
rect 1440 33932 1452 33988
rect 1508 33932 1520 33988
rect 1440 33920 1520 33932
rect 1600 34308 1680 34320
rect 1600 34252 1612 34308
rect 1668 34252 1680 34308
rect 1600 33988 1680 34252
rect 1600 33932 1612 33988
rect 1668 33932 1680 33988
rect 1600 33920 1680 33932
rect 1760 34308 1840 34320
rect 1760 34252 1772 34308
rect 1828 34252 1840 34308
rect 1760 33988 1840 34252
rect 1760 33932 1772 33988
rect 1828 33932 1840 33988
rect 1760 33920 1840 33932
rect 1920 34308 2000 34320
rect 1920 34252 1932 34308
rect 1988 34252 2000 34308
rect 1920 33988 2000 34252
rect 1920 33932 1932 33988
rect 1988 33932 2000 33988
rect 1920 33920 2000 33932
rect 2080 34308 2160 34320
rect 2080 34252 2092 34308
rect 2148 34252 2160 34308
rect 2080 33988 2160 34252
rect 2080 33932 2092 33988
rect 2148 33932 2160 33988
rect 2080 33920 2160 33932
rect 2240 34308 2320 34320
rect 2240 34252 2252 34308
rect 2308 34252 2320 34308
rect 2240 33988 2320 34252
rect 2240 33932 2252 33988
rect 2308 33932 2320 33988
rect 2240 33920 2320 33932
rect 2400 34308 2480 34320
rect 2400 34252 2412 34308
rect 2468 34252 2480 34308
rect 2400 33988 2480 34252
rect 2400 33932 2412 33988
rect 2468 33932 2480 33988
rect 2400 33920 2480 33932
rect 2560 34308 2640 34320
rect 2560 34252 2572 34308
rect 2628 34252 2640 34308
rect 2560 33988 2640 34252
rect 2560 33932 2572 33988
rect 2628 33932 2640 33988
rect 2560 33920 2640 33932
rect 2720 34308 2800 34320
rect 2720 34252 2732 34308
rect 2788 34252 2800 34308
rect 2720 33988 2800 34252
rect 2720 33932 2732 33988
rect 2788 33932 2800 33988
rect 2720 33920 2800 33932
rect 2880 34308 2960 34320
rect 2880 34252 2892 34308
rect 2948 34252 2960 34308
rect 2880 33988 2960 34252
rect 2880 33932 2892 33988
rect 2948 33932 2960 33988
rect 2880 33920 2960 33932
rect 3040 34308 3120 34320
rect 3040 34252 3052 34308
rect 3108 34252 3120 34308
rect 3040 33988 3120 34252
rect 3040 33932 3052 33988
rect 3108 33932 3120 33988
rect 3040 33920 3120 33932
rect 3200 34308 3280 34320
rect 3200 34252 3212 34308
rect 3268 34252 3280 34308
rect 3200 33988 3280 34252
rect 3200 33932 3212 33988
rect 3268 33932 3280 33988
rect 3200 33920 3280 33932
rect 3360 34308 3440 34320
rect 3360 34252 3372 34308
rect 3428 34252 3440 34308
rect 3360 33988 3440 34252
rect 3360 33932 3372 33988
rect 3428 33932 3440 33988
rect 3360 33920 3440 33932
rect 3520 34308 3600 34320
rect 3520 34252 3532 34308
rect 3588 34252 3600 34308
rect 3520 33988 3600 34252
rect 3520 33932 3532 33988
rect 3588 33932 3600 33988
rect 3520 33920 3600 33932
rect 3680 34308 3760 34320
rect 3680 34252 3692 34308
rect 3748 34252 3760 34308
rect 3680 33988 3760 34252
rect 3680 33932 3692 33988
rect 3748 33932 3760 33988
rect 3680 33920 3760 33932
rect 3840 34308 3920 34320
rect 3840 34252 3852 34308
rect 3908 34252 3920 34308
rect 3840 33988 3920 34252
rect 3840 33932 3852 33988
rect 3908 33932 3920 33988
rect 3840 33920 3920 33932
rect 4000 34308 4080 34320
rect 4000 34252 4012 34308
rect 4068 34252 4080 34308
rect 4000 33988 4080 34252
rect 4000 33932 4012 33988
rect 4068 33932 4080 33988
rect 4000 33920 4080 33932
rect 4160 34308 4240 34320
rect 4160 34252 4172 34308
rect 4228 34252 4240 34308
rect 4160 33988 4240 34252
rect 4160 33932 4172 33988
rect 4228 33932 4240 33988
rect 4160 33920 4240 33932
rect 4320 34308 4400 34320
rect 4320 34252 4332 34308
rect 4388 34252 4400 34308
rect 4320 33988 4400 34252
rect 4320 33932 4332 33988
rect 4388 33932 4400 33988
rect 4320 33920 4400 33932
rect 4480 34308 4560 34320
rect 4480 34252 4492 34308
rect 4548 34252 4560 34308
rect 4480 33988 4560 34252
rect 4480 33932 4492 33988
rect 4548 33932 4560 33988
rect 4480 33920 4560 33932
rect 4640 34308 4720 34320
rect 4640 34252 4652 34308
rect 4708 34252 4720 34308
rect 4640 33988 4720 34252
rect 4640 33932 4652 33988
rect 4708 33932 4720 33988
rect 4640 33920 4720 33932
rect 4800 34308 4880 34320
rect 4800 34252 4812 34308
rect 4868 34252 4880 34308
rect 4800 33988 4880 34252
rect 4800 33932 4812 33988
rect 4868 33932 4880 33988
rect 4800 33920 4880 33932
rect 4960 34308 5040 34320
rect 4960 34252 4972 34308
rect 5028 34252 5040 34308
rect 4960 33988 5040 34252
rect 4960 33932 4972 33988
rect 5028 33932 5040 33988
rect 4960 33920 5040 33932
rect 5120 34308 5200 34320
rect 5120 34252 5132 34308
rect 5188 34252 5200 34308
rect 5120 33988 5200 34252
rect 5120 33932 5132 33988
rect 5188 33932 5200 33988
rect 5120 33920 5200 33932
rect 5280 34308 5360 34320
rect 5280 34252 5292 34308
rect 5348 34252 5360 34308
rect 5280 33988 5360 34252
rect 5280 33932 5292 33988
rect 5348 33932 5360 33988
rect 5280 33920 5360 33932
rect 5440 34308 5520 34320
rect 5440 34252 5452 34308
rect 5508 34252 5520 34308
rect 5440 33988 5520 34252
rect 5440 33932 5452 33988
rect 5508 33932 5520 33988
rect 5440 33920 5520 33932
rect 5600 34308 5680 34320
rect 5600 34252 5612 34308
rect 5668 34252 5680 34308
rect 5600 33988 5680 34252
rect 5600 33932 5612 33988
rect 5668 33932 5680 33988
rect 5600 33920 5680 33932
rect 5760 34308 5840 34320
rect 5760 34252 5772 34308
rect 5828 34252 5840 34308
rect 5760 33988 5840 34252
rect 5760 33932 5772 33988
rect 5828 33932 5840 33988
rect 5760 33920 5840 33932
rect 5920 34308 6000 34320
rect 5920 34252 5932 34308
rect 5988 34252 6000 34308
rect 5920 33988 6000 34252
rect 5920 33932 5932 33988
rect 5988 33932 6000 33988
rect 5920 33920 6000 33932
rect 6080 34308 6160 34320
rect 6080 34252 6092 34308
rect 6148 34252 6160 34308
rect 6080 33988 6160 34252
rect 6080 33932 6092 33988
rect 6148 33932 6160 33988
rect 6080 33920 6160 33932
rect 6240 34308 6320 34320
rect 6240 34252 6252 34308
rect 6308 34252 6320 34308
rect 6240 33988 6320 34252
rect 6240 33932 6252 33988
rect 6308 33932 6320 33988
rect 6240 33920 6320 33932
rect 6400 34308 6480 34320
rect 6400 34252 6412 34308
rect 6468 34252 6480 34308
rect 6400 33988 6480 34252
rect 6400 33932 6412 33988
rect 6468 33932 6480 33988
rect 6400 33920 6480 33932
rect 6560 34308 6640 34320
rect 6560 34252 6572 34308
rect 6628 34252 6640 34308
rect 6560 33988 6640 34252
rect 6560 33932 6572 33988
rect 6628 33932 6640 33988
rect 6560 33920 6640 33932
rect 6720 34308 6800 34320
rect 6720 34252 6732 34308
rect 6788 34252 6800 34308
rect 6720 33988 6800 34252
rect 6720 33932 6732 33988
rect 6788 33932 6800 33988
rect 6720 33920 6800 33932
rect 6880 34308 6960 34320
rect 6880 34252 6892 34308
rect 6948 34252 6960 34308
rect 6880 33988 6960 34252
rect 6880 33932 6892 33988
rect 6948 33932 6960 33988
rect 6880 33920 6960 33932
rect 7040 34308 7120 34320
rect 7040 34252 7052 34308
rect 7108 34252 7120 34308
rect 7040 33988 7120 34252
rect 7040 33932 7052 33988
rect 7108 33932 7120 33988
rect 7040 33920 7120 33932
rect 7200 34308 7280 34320
rect 7200 34252 7212 34308
rect 7268 34252 7280 34308
rect 7200 33988 7280 34252
rect 7200 33932 7212 33988
rect 7268 33932 7280 33988
rect 7200 33920 7280 33932
rect 7360 34308 7440 34320
rect 7360 34252 7372 34308
rect 7428 34252 7440 34308
rect 7360 33988 7440 34252
rect 7360 33932 7372 33988
rect 7428 33932 7440 33988
rect 7360 33920 7440 33932
rect 7520 34308 7600 34320
rect 7520 34252 7532 34308
rect 7588 34252 7600 34308
rect 7520 33988 7600 34252
rect 7520 33932 7532 33988
rect 7588 33932 7600 33988
rect 7520 33920 7600 33932
rect 7680 34308 7760 34320
rect 7680 34252 7692 34308
rect 7748 34252 7760 34308
rect 7680 33988 7760 34252
rect 7680 33932 7692 33988
rect 7748 33932 7760 33988
rect 7680 33920 7760 33932
rect 7840 34308 7920 34320
rect 7840 34252 7852 34308
rect 7908 34252 7920 34308
rect 7840 33988 7920 34252
rect 7840 33932 7852 33988
rect 7908 33932 7920 33988
rect 7840 33920 7920 33932
rect 8000 34308 8080 34320
rect 8000 34252 8012 34308
rect 8068 34252 8080 34308
rect 8000 33988 8080 34252
rect 8000 33932 8012 33988
rect 8068 33932 8080 33988
rect 8000 33920 8080 33932
rect 8160 34308 8240 34320
rect 8160 34252 8172 34308
rect 8228 34252 8240 34308
rect 8160 33988 8240 34252
rect 8160 33932 8172 33988
rect 8228 33932 8240 33988
rect 8160 33920 8240 33932
rect 8320 34308 8400 34320
rect 8320 34252 8332 34308
rect 8388 34252 8400 34308
rect 8320 33988 8400 34252
rect 8320 33932 8332 33988
rect 8388 33932 8400 33988
rect 8320 33920 8400 33932
rect 0 33828 80 33840
rect 0 33772 12 33828
rect 68 33772 80 33828
rect 0 33508 80 33772
rect 0 33452 12 33508
rect 68 33452 80 33508
rect 0 33440 80 33452
rect 160 33828 240 33840
rect 160 33772 172 33828
rect 228 33772 240 33828
rect 160 33508 240 33772
rect 160 33452 172 33508
rect 228 33452 240 33508
rect 160 33440 240 33452
rect 320 33828 400 33840
rect 320 33772 332 33828
rect 388 33772 400 33828
rect 320 33508 400 33772
rect 320 33452 332 33508
rect 388 33452 400 33508
rect 320 33440 400 33452
rect 480 33828 560 33840
rect 480 33772 492 33828
rect 548 33772 560 33828
rect 480 33508 560 33772
rect 480 33452 492 33508
rect 548 33452 560 33508
rect 480 33440 560 33452
rect 640 33828 720 33840
rect 640 33772 652 33828
rect 708 33772 720 33828
rect 640 33508 720 33772
rect 640 33452 652 33508
rect 708 33452 720 33508
rect 640 33440 720 33452
rect 800 33828 880 33840
rect 800 33772 812 33828
rect 868 33772 880 33828
rect 800 33508 880 33772
rect 800 33452 812 33508
rect 868 33452 880 33508
rect 800 33440 880 33452
rect 960 33828 1040 33840
rect 960 33772 972 33828
rect 1028 33772 1040 33828
rect 960 33508 1040 33772
rect 960 33452 972 33508
rect 1028 33452 1040 33508
rect 960 33440 1040 33452
rect 1120 33828 1200 33840
rect 1120 33772 1132 33828
rect 1188 33772 1200 33828
rect 1120 33508 1200 33772
rect 1120 33452 1132 33508
rect 1188 33452 1200 33508
rect 1120 33440 1200 33452
rect 1280 33828 1360 33840
rect 1280 33772 1292 33828
rect 1348 33772 1360 33828
rect 1280 33508 1360 33772
rect 1280 33452 1292 33508
rect 1348 33452 1360 33508
rect 1280 33440 1360 33452
rect 1440 33828 1520 33840
rect 1440 33772 1452 33828
rect 1508 33772 1520 33828
rect 1440 33508 1520 33772
rect 1440 33452 1452 33508
rect 1508 33452 1520 33508
rect 1440 33440 1520 33452
rect 1600 33828 1680 33840
rect 1600 33772 1612 33828
rect 1668 33772 1680 33828
rect 1600 33508 1680 33772
rect 1600 33452 1612 33508
rect 1668 33452 1680 33508
rect 1600 33440 1680 33452
rect 1760 33828 1840 33840
rect 1760 33772 1772 33828
rect 1828 33772 1840 33828
rect 1760 33508 1840 33772
rect 1760 33452 1772 33508
rect 1828 33452 1840 33508
rect 1760 33440 1840 33452
rect 1920 33828 2000 33840
rect 1920 33772 1932 33828
rect 1988 33772 2000 33828
rect 1920 33508 2000 33772
rect 1920 33452 1932 33508
rect 1988 33452 2000 33508
rect 1920 33440 2000 33452
rect 2080 33828 2160 33840
rect 2080 33772 2092 33828
rect 2148 33772 2160 33828
rect 2080 33508 2160 33772
rect 2080 33452 2092 33508
rect 2148 33452 2160 33508
rect 2080 33440 2160 33452
rect 2240 33828 2320 33840
rect 2240 33772 2252 33828
rect 2308 33772 2320 33828
rect 2240 33508 2320 33772
rect 2240 33452 2252 33508
rect 2308 33452 2320 33508
rect 2240 33440 2320 33452
rect 2400 33828 2480 33840
rect 2400 33772 2412 33828
rect 2468 33772 2480 33828
rect 2400 33508 2480 33772
rect 2400 33452 2412 33508
rect 2468 33452 2480 33508
rect 2400 33440 2480 33452
rect 2560 33828 2640 33840
rect 2560 33772 2572 33828
rect 2628 33772 2640 33828
rect 2560 33508 2640 33772
rect 2560 33452 2572 33508
rect 2628 33452 2640 33508
rect 2560 33440 2640 33452
rect 2720 33828 2800 33840
rect 2720 33772 2732 33828
rect 2788 33772 2800 33828
rect 2720 33508 2800 33772
rect 2720 33452 2732 33508
rect 2788 33452 2800 33508
rect 2720 33440 2800 33452
rect 2880 33828 2960 33840
rect 2880 33772 2892 33828
rect 2948 33772 2960 33828
rect 2880 33508 2960 33772
rect 2880 33452 2892 33508
rect 2948 33452 2960 33508
rect 2880 33440 2960 33452
rect 3040 33828 3120 33840
rect 3040 33772 3052 33828
rect 3108 33772 3120 33828
rect 3040 33508 3120 33772
rect 3040 33452 3052 33508
rect 3108 33452 3120 33508
rect 3040 33440 3120 33452
rect 3200 33828 3280 33840
rect 3200 33772 3212 33828
rect 3268 33772 3280 33828
rect 3200 33508 3280 33772
rect 3200 33452 3212 33508
rect 3268 33452 3280 33508
rect 3200 33440 3280 33452
rect 3360 33828 3440 33840
rect 3360 33772 3372 33828
rect 3428 33772 3440 33828
rect 3360 33508 3440 33772
rect 3360 33452 3372 33508
rect 3428 33452 3440 33508
rect 3360 33440 3440 33452
rect 3520 33828 3600 33840
rect 3520 33772 3532 33828
rect 3588 33772 3600 33828
rect 3520 33508 3600 33772
rect 3520 33452 3532 33508
rect 3588 33452 3600 33508
rect 3520 33440 3600 33452
rect 3680 33828 3760 33840
rect 3680 33772 3692 33828
rect 3748 33772 3760 33828
rect 3680 33508 3760 33772
rect 3680 33452 3692 33508
rect 3748 33452 3760 33508
rect 3680 33440 3760 33452
rect 3840 33828 3920 33840
rect 3840 33772 3852 33828
rect 3908 33772 3920 33828
rect 3840 33508 3920 33772
rect 3840 33452 3852 33508
rect 3908 33452 3920 33508
rect 3840 33440 3920 33452
rect 4000 33828 4080 33840
rect 4000 33772 4012 33828
rect 4068 33772 4080 33828
rect 4000 33508 4080 33772
rect 4000 33452 4012 33508
rect 4068 33452 4080 33508
rect 4000 33440 4080 33452
rect 4160 33828 4240 33840
rect 4160 33772 4172 33828
rect 4228 33772 4240 33828
rect 4160 33508 4240 33772
rect 4160 33452 4172 33508
rect 4228 33452 4240 33508
rect 4160 33440 4240 33452
rect 4320 33828 4400 33840
rect 4320 33772 4332 33828
rect 4388 33772 4400 33828
rect 4320 33508 4400 33772
rect 4320 33452 4332 33508
rect 4388 33452 4400 33508
rect 4320 33440 4400 33452
rect 4480 33828 4560 33840
rect 4480 33772 4492 33828
rect 4548 33772 4560 33828
rect 4480 33508 4560 33772
rect 4480 33452 4492 33508
rect 4548 33452 4560 33508
rect 4480 33440 4560 33452
rect 4640 33828 4720 33840
rect 4640 33772 4652 33828
rect 4708 33772 4720 33828
rect 4640 33508 4720 33772
rect 4640 33452 4652 33508
rect 4708 33452 4720 33508
rect 4640 33440 4720 33452
rect 4800 33828 4880 33840
rect 4800 33772 4812 33828
rect 4868 33772 4880 33828
rect 4800 33508 4880 33772
rect 4800 33452 4812 33508
rect 4868 33452 4880 33508
rect 4800 33440 4880 33452
rect 4960 33828 5040 33840
rect 4960 33772 4972 33828
rect 5028 33772 5040 33828
rect 4960 33508 5040 33772
rect 4960 33452 4972 33508
rect 5028 33452 5040 33508
rect 4960 33440 5040 33452
rect 5120 33828 5200 33840
rect 5120 33772 5132 33828
rect 5188 33772 5200 33828
rect 5120 33508 5200 33772
rect 5120 33452 5132 33508
rect 5188 33452 5200 33508
rect 5120 33440 5200 33452
rect 5280 33828 5360 33840
rect 5280 33772 5292 33828
rect 5348 33772 5360 33828
rect 5280 33508 5360 33772
rect 5280 33452 5292 33508
rect 5348 33452 5360 33508
rect 5280 33440 5360 33452
rect 5440 33828 5520 33840
rect 5440 33772 5452 33828
rect 5508 33772 5520 33828
rect 5440 33508 5520 33772
rect 5440 33452 5452 33508
rect 5508 33452 5520 33508
rect 5440 33440 5520 33452
rect 5600 33828 5680 33840
rect 5600 33772 5612 33828
rect 5668 33772 5680 33828
rect 5600 33508 5680 33772
rect 5600 33452 5612 33508
rect 5668 33452 5680 33508
rect 5600 33440 5680 33452
rect 5760 33828 5840 33840
rect 5760 33772 5772 33828
rect 5828 33772 5840 33828
rect 5760 33508 5840 33772
rect 5760 33452 5772 33508
rect 5828 33452 5840 33508
rect 5760 33440 5840 33452
rect 5920 33828 6000 33840
rect 5920 33772 5932 33828
rect 5988 33772 6000 33828
rect 5920 33508 6000 33772
rect 5920 33452 5932 33508
rect 5988 33452 6000 33508
rect 5920 33440 6000 33452
rect 6080 33828 6160 33840
rect 6080 33772 6092 33828
rect 6148 33772 6160 33828
rect 6080 33508 6160 33772
rect 6080 33452 6092 33508
rect 6148 33452 6160 33508
rect 6080 33440 6160 33452
rect 6240 33828 6320 33840
rect 6240 33772 6252 33828
rect 6308 33772 6320 33828
rect 6240 33508 6320 33772
rect 6240 33452 6252 33508
rect 6308 33452 6320 33508
rect 6240 33440 6320 33452
rect 6400 33828 6480 33840
rect 6400 33772 6412 33828
rect 6468 33772 6480 33828
rect 6400 33508 6480 33772
rect 6400 33452 6412 33508
rect 6468 33452 6480 33508
rect 6400 33440 6480 33452
rect 6560 33828 6640 33840
rect 6560 33772 6572 33828
rect 6628 33772 6640 33828
rect 6560 33508 6640 33772
rect 6560 33452 6572 33508
rect 6628 33452 6640 33508
rect 6560 33440 6640 33452
rect 6720 33828 6800 33840
rect 6720 33772 6732 33828
rect 6788 33772 6800 33828
rect 6720 33508 6800 33772
rect 6720 33452 6732 33508
rect 6788 33452 6800 33508
rect 6720 33440 6800 33452
rect 6880 33828 6960 33840
rect 6880 33772 6892 33828
rect 6948 33772 6960 33828
rect 6880 33508 6960 33772
rect 6880 33452 6892 33508
rect 6948 33452 6960 33508
rect 6880 33440 6960 33452
rect 7040 33828 7120 33840
rect 7040 33772 7052 33828
rect 7108 33772 7120 33828
rect 7040 33508 7120 33772
rect 7040 33452 7052 33508
rect 7108 33452 7120 33508
rect 7040 33440 7120 33452
rect 7200 33828 7280 33840
rect 7200 33772 7212 33828
rect 7268 33772 7280 33828
rect 7200 33508 7280 33772
rect 7200 33452 7212 33508
rect 7268 33452 7280 33508
rect 7200 33440 7280 33452
rect 7360 33828 7440 33840
rect 7360 33772 7372 33828
rect 7428 33772 7440 33828
rect 7360 33508 7440 33772
rect 7360 33452 7372 33508
rect 7428 33452 7440 33508
rect 7360 33440 7440 33452
rect 7520 33828 7600 33840
rect 7520 33772 7532 33828
rect 7588 33772 7600 33828
rect 7520 33508 7600 33772
rect 7520 33452 7532 33508
rect 7588 33452 7600 33508
rect 7520 33440 7600 33452
rect 7680 33828 7760 33840
rect 7680 33772 7692 33828
rect 7748 33772 7760 33828
rect 7680 33508 7760 33772
rect 7680 33452 7692 33508
rect 7748 33452 7760 33508
rect 7680 33440 7760 33452
rect 7840 33828 7920 33840
rect 7840 33772 7852 33828
rect 7908 33772 7920 33828
rect 7840 33508 7920 33772
rect 7840 33452 7852 33508
rect 7908 33452 7920 33508
rect 7840 33440 7920 33452
rect 8000 33828 8080 33840
rect 8000 33772 8012 33828
rect 8068 33772 8080 33828
rect 8000 33508 8080 33772
rect 8000 33452 8012 33508
rect 8068 33452 8080 33508
rect 8000 33440 8080 33452
rect 8160 33828 8240 33840
rect 8160 33772 8172 33828
rect 8228 33772 8240 33828
rect 8160 33508 8240 33772
rect 8160 33452 8172 33508
rect 8228 33452 8240 33508
rect 8160 33440 8240 33452
rect 8320 33828 8400 33840
rect 8320 33772 8332 33828
rect 8388 33772 8400 33828
rect 8320 33508 8400 33772
rect 8320 33452 8332 33508
rect 8388 33452 8400 33508
rect 8320 33440 8400 33452
rect 8480 33440 8560 36972
rect 8640 37188 8720 37440
rect 8640 37132 8652 37188
rect 8708 37132 8720 37188
rect 8640 33440 8720 37132
rect 8800 37348 8880 37440
rect 8800 37292 8812 37348
rect 8868 37292 8880 37348
rect 8800 37028 8880 37292
rect 8800 36972 8812 37028
rect 8868 36972 8880 37028
rect 8800 33440 8880 36972
rect 8960 36868 9040 37440
rect 8960 36812 8972 36868
rect 9028 36812 9040 36868
rect 8960 36548 9040 36812
rect 8960 36492 8972 36548
rect 9028 36492 9040 36548
rect 8960 33440 9040 36492
rect 9120 36708 9200 37440
rect 9120 36652 9132 36708
rect 9188 36652 9200 36708
rect 9120 33440 9200 36652
rect 9280 36868 9360 37440
rect 9280 36812 9292 36868
rect 9348 36812 9360 36868
rect 9280 36548 9360 36812
rect 9280 36492 9292 36548
rect 9348 36492 9360 36548
rect 9280 33440 9360 36492
rect 9440 36388 9520 37440
rect 9440 36332 9452 36388
rect 9508 36332 9520 36388
rect 9440 36068 9520 36332
rect 9440 36012 9452 36068
rect 9508 36012 9520 36068
rect 9440 35748 9520 36012
rect 9440 35692 9452 35748
rect 9508 35692 9520 35748
rect 9440 35428 9520 35692
rect 9440 35372 9452 35428
rect 9508 35372 9520 35428
rect 9440 35108 9520 35372
rect 9440 35052 9452 35108
rect 9508 35052 9520 35108
rect 9440 34788 9520 35052
rect 9440 34732 9452 34788
rect 9508 34732 9520 34788
rect 9440 34468 9520 34732
rect 9440 34412 9452 34468
rect 9508 34412 9520 34468
rect 9440 33440 9520 34412
rect 9600 36228 9680 37440
rect 9600 36172 9612 36228
rect 9668 36172 9680 36228
rect 9600 33440 9680 36172
rect 9760 36388 9840 37440
rect 9760 36332 9772 36388
rect 9828 36332 9840 36388
rect 9760 36068 9840 36332
rect 9760 36012 9772 36068
rect 9828 36012 9840 36068
rect 9760 35748 9840 36012
rect 9760 35692 9772 35748
rect 9828 35692 9840 35748
rect 9760 35428 9840 35692
rect 9760 35372 9772 35428
rect 9828 35372 9840 35428
rect 9760 35108 9840 35372
rect 9760 35052 9772 35108
rect 9828 35052 9840 35108
rect 9760 34788 9840 35052
rect 9760 34732 9772 34788
rect 9828 34732 9840 34788
rect 9760 34468 9840 34732
rect 9760 34412 9772 34468
rect 9828 34412 9840 34468
rect 9760 33440 9840 34412
rect 9920 35908 10000 37440
rect 9920 35852 9932 35908
rect 9988 35852 10000 35908
rect 9920 33440 10000 35852
rect 10080 36388 10160 37440
rect 10080 36332 10092 36388
rect 10148 36332 10160 36388
rect 10080 36068 10160 36332
rect 10080 36012 10092 36068
rect 10148 36012 10160 36068
rect 10080 35748 10160 36012
rect 10080 35692 10092 35748
rect 10148 35692 10160 35748
rect 10080 35428 10160 35692
rect 10080 35372 10092 35428
rect 10148 35372 10160 35428
rect 10080 35108 10160 35372
rect 10080 35052 10092 35108
rect 10148 35052 10160 35108
rect 10080 34788 10160 35052
rect 10080 34732 10092 34788
rect 10148 34732 10160 34788
rect 10080 34468 10160 34732
rect 10080 34412 10092 34468
rect 10148 34412 10160 34468
rect 10080 33440 10160 34412
rect 10240 35588 10320 37440
rect 10240 35532 10252 35588
rect 10308 35532 10320 35588
rect 10240 33440 10320 35532
rect 10400 36388 10480 37440
rect 10400 36332 10412 36388
rect 10468 36332 10480 36388
rect 10400 36068 10480 36332
rect 10400 36012 10412 36068
rect 10468 36012 10480 36068
rect 10400 35748 10480 36012
rect 10400 35692 10412 35748
rect 10468 35692 10480 35748
rect 10400 35428 10480 35692
rect 10400 35372 10412 35428
rect 10468 35372 10480 35428
rect 10400 35108 10480 35372
rect 10400 35052 10412 35108
rect 10468 35052 10480 35108
rect 10400 34788 10480 35052
rect 10400 34732 10412 34788
rect 10468 34732 10480 34788
rect 10400 34468 10480 34732
rect 10400 34412 10412 34468
rect 10468 34412 10480 34468
rect 10400 33440 10480 34412
rect 10560 35268 10640 37440
rect 10560 35212 10572 35268
rect 10628 35212 10640 35268
rect 10560 33440 10640 35212
rect 10720 36388 10800 37440
rect 10720 36332 10732 36388
rect 10788 36332 10800 36388
rect 10720 36068 10800 36332
rect 10720 36012 10732 36068
rect 10788 36012 10800 36068
rect 10720 35748 10800 36012
rect 10720 35692 10732 35748
rect 10788 35692 10800 35748
rect 10720 35428 10800 35692
rect 10720 35372 10732 35428
rect 10788 35372 10800 35428
rect 10720 35108 10800 35372
rect 10720 35052 10732 35108
rect 10788 35052 10800 35108
rect 10720 34788 10800 35052
rect 10720 34732 10732 34788
rect 10788 34732 10800 34788
rect 10720 34468 10800 34732
rect 10720 34412 10732 34468
rect 10788 34412 10800 34468
rect 10720 33440 10800 34412
rect 10880 34948 10960 37440
rect 10880 34892 10892 34948
rect 10948 34892 10960 34948
rect 10880 33440 10960 34892
rect 11040 36388 11120 37440
rect 11040 36332 11052 36388
rect 11108 36332 11120 36388
rect 11040 36068 11120 36332
rect 11040 36012 11052 36068
rect 11108 36012 11120 36068
rect 11040 35748 11120 36012
rect 11040 35692 11052 35748
rect 11108 35692 11120 35748
rect 11040 35428 11120 35692
rect 11040 35372 11052 35428
rect 11108 35372 11120 35428
rect 11040 35108 11120 35372
rect 11040 35052 11052 35108
rect 11108 35052 11120 35108
rect 11040 34788 11120 35052
rect 11040 34732 11052 34788
rect 11108 34732 11120 34788
rect 11040 34468 11120 34732
rect 11040 34412 11052 34468
rect 11108 34412 11120 34468
rect 11040 33440 11120 34412
rect 11200 34628 11280 37440
rect 11200 34572 11212 34628
rect 11268 34572 11280 34628
rect 11200 33440 11280 34572
rect 11360 36388 11440 37440
rect 11360 36332 11372 36388
rect 11428 36332 11440 36388
rect 11360 36068 11440 36332
rect 11360 36012 11372 36068
rect 11428 36012 11440 36068
rect 11360 35748 11440 36012
rect 11360 35692 11372 35748
rect 11428 35692 11440 35748
rect 11360 35428 11440 35692
rect 11360 35372 11372 35428
rect 11428 35372 11440 35428
rect 11360 35108 11440 35372
rect 11360 35052 11372 35108
rect 11428 35052 11440 35108
rect 11360 34788 11440 35052
rect 11360 34732 11372 34788
rect 11428 34732 11440 34788
rect 11360 34468 11440 34732
rect 11360 34412 11372 34468
rect 11428 34412 11440 34468
rect 11360 33440 11440 34412
rect 11520 34308 11600 37440
rect 11520 34252 11532 34308
rect 11588 34252 11600 34308
rect 11520 33988 11600 34252
rect 11520 33932 11532 33988
rect 11588 33932 11600 33988
rect 11520 33440 11600 33932
rect 11680 34148 11760 37440
rect 11680 34092 11692 34148
rect 11748 34092 11760 34148
rect 11680 33440 11760 34092
rect 11840 34308 11920 37440
rect 11840 34252 11852 34308
rect 11908 34252 11920 34308
rect 11840 33988 11920 34252
rect 11840 33932 11852 33988
rect 11908 33932 11920 33988
rect 11840 33440 11920 33932
rect 12000 33828 12080 37440
rect 12000 33772 12012 33828
rect 12068 33772 12080 33828
rect 12000 33508 12080 33772
rect 12000 33452 12012 33508
rect 12068 33452 12080 33508
rect 12000 33440 12080 33452
rect 12160 33668 12240 37440
rect 12160 33612 12172 33668
rect 12228 33612 12240 33668
rect 12160 33440 12240 33612
rect 12320 33828 12400 37440
rect 12480 37348 12560 37360
rect 12480 37292 12492 37348
rect 12548 37292 12560 37348
rect 12480 37028 12560 37292
rect 12480 36972 12492 37028
rect 12548 36972 12560 37028
rect 12480 36960 12560 36972
rect 12640 37348 12720 37360
rect 12640 37292 12652 37348
rect 12708 37292 12720 37348
rect 12640 37028 12720 37292
rect 12640 36972 12652 37028
rect 12708 36972 12720 37028
rect 12640 36960 12720 36972
rect 12800 37348 12880 37360
rect 12800 37292 12812 37348
rect 12868 37292 12880 37348
rect 12800 37028 12880 37292
rect 12800 36972 12812 37028
rect 12868 36972 12880 37028
rect 12800 36960 12880 36972
rect 12960 37348 13040 37360
rect 12960 37292 12972 37348
rect 13028 37292 13040 37348
rect 12960 37028 13040 37292
rect 12960 36972 12972 37028
rect 13028 36972 13040 37028
rect 12960 36960 13040 36972
rect 13120 37348 13200 37360
rect 13120 37292 13132 37348
rect 13188 37292 13200 37348
rect 13120 37028 13200 37292
rect 13120 36972 13132 37028
rect 13188 36972 13200 37028
rect 13120 36960 13200 36972
rect 13280 37348 13360 37360
rect 13280 37292 13292 37348
rect 13348 37292 13360 37348
rect 13280 37028 13360 37292
rect 13280 36972 13292 37028
rect 13348 36972 13360 37028
rect 13280 36960 13360 36972
rect 13440 37348 13520 37360
rect 13440 37292 13452 37348
rect 13508 37292 13520 37348
rect 13440 37028 13520 37292
rect 13440 36972 13452 37028
rect 13508 36972 13520 37028
rect 13440 36960 13520 36972
rect 13600 37348 13680 37360
rect 13600 37292 13612 37348
rect 13668 37292 13680 37348
rect 13600 37028 13680 37292
rect 13600 36972 13612 37028
rect 13668 36972 13680 37028
rect 13600 36960 13680 36972
rect 13760 37348 13840 37360
rect 13760 37292 13772 37348
rect 13828 37292 13840 37348
rect 13760 37028 13840 37292
rect 13760 36972 13772 37028
rect 13828 36972 13840 37028
rect 13760 36960 13840 36972
rect 13920 37348 14000 37360
rect 13920 37292 13932 37348
rect 13988 37292 14000 37348
rect 13920 37028 14000 37292
rect 13920 36972 13932 37028
rect 13988 36972 14000 37028
rect 13920 36960 14000 36972
rect 14080 37348 14160 37360
rect 14080 37292 14092 37348
rect 14148 37292 14160 37348
rect 14080 37028 14160 37292
rect 14080 36972 14092 37028
rect 14148 36972 14160 37028
rect 14080 36960 14160 36972
rect 14240 37348 14320 37360
rect 14240 37292 14252 37348
rect 14308 37292 14320 37348
rect 14240 37028 14320 37292
rect 14240 36972 14252 37028
rect 14308 36972 14320 37028
rect 14240 36960 14320 36972
rect 14400 37348 14480 37360
rect 14400 37292 14412 37348
rect 14468 37292 14480 37348
rect 14400 37028 14480 37292
rect 14400 36972 14412 37028
rect 14468 36972 14480 37028
rect 14400 36960 14480 36972
rect 14560 37348 14640 37360
rect 14560 37292 14572 37348
rect 14628 37292 14640 37348
rect 14560 37028 14640 37292
rect 14560 36972 14572 37028
rect 14628 36972 14640 37028
rect 14560 36960 14640 36972
rect 14720 37348 14800 37360
rect 14720 37292 14732 37348
rect 14788 37292 14800 37348
rect 14720 37028 14800 37292
rect 14720 36972 14732 37028
rect 14788 36972 14800 37028
rect 14720 36960 14800 36972
rect 14880 37348 14960 37360
rect 14880 37292 14892 37348
rect 14948 37292 14960 37348
rect 14880 37028 14960 37292
rect 14880 36972 14892 37028
rect 14948 36972 14960 37028
rect 14880 36960 14960 36972
rect 15040 37348 15120 37360
rect 15040 37292 15052 37348
rect 15108 37292 15120 37348
rect 15040 37028 15120 37292
rect 15040 36972 15052 37028
rect 15108 36972 15120 37028
rect 15040 36960 15120 36972
rect 15200 37348 15280 37360
rect 15200 37292 15212 37348
rect 15268 37292 15280 37348
rect 15200 37028 15280 37292
rect 15200 36972 15212 37028
rect 15268 36972 15280 37028
rect 15200 36960 15280 36972
rect 15360 37348 15440 37360
rect 15360 37292 15372 37348
rect 15428 37292 15440 37348
rect 15360 37028 15440 37292
rect 15360 36972 15372 37028
rect 15428 36972 15440 37028
rect 15360 36960 15440 36972
rect 15520 37348 15600 37360
rect 15520 37292 15532 37348
rect 15588 37292 15600 37348
rect 15520 37028 15600 37292
rect 15520 36972 15532 37028
rect 15588 36972 15600 37028
rect 15520 36960 15600 36972
rect 15680 37348 15760 37360
rect 15680 37292 15692 37348
rect 15748 37292 15760 37348
rect 15680 37028 15760 37292
rect 15680 36972 15692 37028
rect 15748 36972 15760 37028
rect 15680 36960 15760 36972
rect 15840 37348 15920 37360
rect 15840 37292 15852 37348
rect 15908 37292 15920 37348
rect 15840 37028 15920 37292
rect 15840 36972 15852 37028
rect 15908 36972 15920 37028
rect 15840 36960 15920 36972
rect 16000 37348 16080 37360
rect 16000 37292 16012 37348
rect 16068 37292 16080 37348
rect 16000 37028 16080 37292
rect 16000 36972 16012 37028
rect 16068 36972 16080 37028
rect 16000 36960 16080 36972
rect 16160 37348 16240 37360
rect 16160 37292 16172 37348
rect 16228 37292 16240 37348
rect 16160 37028 16240 37292
rect 16160 36972 16172 37028
rect 16228 36972 16240 37028
rect 16160 36960 16240 36972
rect 16320 37348 16400 37360
rect 16320 37292 16332 37348
rect 16388 37292 16400 37348
rect 16320 37028 16400 37292
rect 16320 36972 16332 37028
rect 16388 36972 16400 37028
rect 16320 36960 16400 36972
rect 16480 37348 16560 37360
rect 16480 37292 16492 37348
rect 16548 37292 16560 37348
rect 16480 37028 16560 37292
rect 16480 36972 16492 37028
rect 16548 36972 16560 37028
rect 16480 36960 16560 36972
rect 16640 37348 16720 37360
rect 16640 37292 16652 37348
rect 16708 37292 16720 37348
rect 16640 37028 16720 37292
rect 16640 36972 16652 37028
rect 16708 36972 16720 37028
rect 16640 36960 16720 36972
rect 16800 37348 16880 37360
rect 16800 37292 16812 37348
rect 16868 37292 16880 37348
rect 16800 37028 16880 37292
rect 16800 36972 16812 37028
rect 16868 36972 16880 37028
rect 16800 36960 16880 36972
rect 16960 37348 17040 37360
rect 16960 37292 16972 37348
rect 17028 37292 17040 37348
rect 16960 37028 17040 37292
rect 16960 36972 16972 37028
rect 17028 36972 17040 37028
rect 16960 36960 17040 36972
rect 17120 37348 17200 37360
rect 17120 37292 17132 37348
rect 17188 37292 17200 37348
rect 17120 37028 17200 37292
rect 17120 36972 17132 37028
rect 17188 36972 17200 37028
rect 17120 36960 17200 36972
rect 17280 37348 17360 37360
rect 17280 37292 17292 37348
rect 17348 37292 17360 37348
rect 17280 37028 17360 37292
rect 17280 36972 17292 37028
rect 17348 36972 17360 37028
rect 17280 36960 17360 36972
rect 17440 37348 17520 37360
rect 17440 37292 17452 37348
rect 17508 37292 17520 37348
rect 17440 37028 17520 37292
rect 17440 36972 17452 37028
rect 17508 36972 17520 37028
rect 17440 36960 17520 36972
rect 17600 37348 17680 37360
rect 17600 37292 17612 37348
rect 17668 37292 17680 37348
rect 17600 37028 17680 37292
rect 17600 36972 17612 37028
rect 17668 36972 17680 37028
rect 17600 36960 17680 36972
rect 17760 37348 17840 37360
rect 17760 37292 17772 37348
rect 17828 37292 17840 37348
rect 17760 37028 17840 37292
rect 17760 36972 17772 37028
rect 17828 36972 17840 37028
rect 17760 36960 17840 36972
rect 17920 37348 18000 37360
rect 17920 37292 17932 37348
rect 17988 37292 18000 37348
rect 17920 37028 18000 37292
rect 17920 36972 17932 37028
rect 17988 36972 18000 37028
rect 17920 36960 18000 36972
rect 18080 37348 18160 37360
rect 18080 37292 18092 37348
rect 18148 37292 18160 37348
rect 18080 37028 18160 37292
rect 18080 36972 18092 37028
rect 18148 36972 18160 37028
rect 18080 36960 18160 36972
rect 18240 37348 18320 37360
rect 18240 37292 18252 37348
rect 18308 37292 18320 37348
rect 18240 37028 18320 37292
rect 18240 36972 18252 37028
rect 18308 36972 18320 37028
rect 18240 36960 18320 36972
rect 18400 37348 18480 37360
rect 18400 37292 18412 37348
rect 18468 37292 18480 37348
rect 18400 37028 18480 37292
rect 18400 36972 18412 37028
rect 18468 36972 18480 37028
rect 18400 36960 18480 36972
rect 18560 37348 18640 37360
rect 18560 37292 18572 37348
rect 18628 37292 18640 37348
rect 18560 37028 18640 37292
rect 18560 36972 18572 37028
rect 18628 36972 18640 37028
rect 18560 36960 18640 36972
rect 18720 37348 18800 37360
rect 18720 37292 18732 37348
rect 18788 37292 18800 37348
rect 18720 37028 18800 37292
rect 18720 36972 18732 37028
rect 18788 36972 18800 37028
rect 18720 36960 18800 36972
rect 18880 37348 18960 37360
rect 18880 37292 18892 37348
rect 18948 37292 18960 37348
rect 18880 37028 18960 37292
rect 18880 36972 18892 37028
rect 18948 36972 18960 37028
rect 18880 36960 18960 36972
rect 12480 36868 12560 36880
rect 12480 36812 12492 36868
rect 12548 36812 12560 36868
rect 12480 36548 12560 36812
rect 12480 36492 12492 36548
rect 12548 36492 12560 36548
rect 12480 36480 12560 36492
rect 12640 36868 12720 36880
rect 12640 36812 12652 36868
rect 12708 36812 12720 36868
rect 12640 36548 12720 36812
rect 12640 36492 12652 36548
rect 12708 36492 12720 36548
rect 12640 36480 12720 36492
rect 12800 36868 12880 36880
rect 12800 36812 12812 36868
rect 12868 36812 12880 36868
rect 12800 36548 12880 36812
rect 12800 36492 12812 36548
rect 12868 36492 12880 36548
rect 12800 36480 12880 36492
rect 12960 36868 13040 36880
rect 12960 36812 12972 36868
rect 13028 36812 13040 36868
rect 12960 36548 13040 36812
rect 12960 36492 12972 36548
rect 13028 36492 13040 36548
rect 12960 36480 13040 36492
rect 13120 36868 13200 36880
rect 13120 36812 13132 36868
rect 13188 36812 13200 36868
rect 13120 36548 13200 36812
rect 13120 36492 13132 36548
rect 13188 36492 13200 36548
rect 13120 36480 13200 36492
rect 13280 36868 13360 36880
rect 13280 36812 13292 36868
rect 13348 36812 13360 36868
rect 13280 36548 13360 36812
rect 13280 36492 13292 36548
rect 13348 36492 13360 36548
rect 13280 36480 13360 36492
rect 13440 36868 13520 36880
rect 13440 36812 13452 36868
rect 13508 36812 13520 36868
rect 13440 36548 13520 36812
rect 13440 36492 13452 36548
rect 13508 36492 13520 36548
rect 13440 36480 13520 36492
rect 13600 36868 13680 36880
rect 13600 36812 13612 36868
rect 13668 36812 13680 36868
rect 13600 36548 13680 36812
rect 13600 36492 13612 36548
rect 13668 36492 13680 36548
rect 13600 36480 13680 36492
rect 13760 36868 13840 36880
rect 13760 36812 13772 36868
rect 13828 36812 13840 36868
rect 13760 36548 13840 36812
rect 13760 36492 13772 36548
rect 13828 36492 13840 36548
rect 13760 36480 13840 36492
rect 13920 36868 14000 36880
rect 13920 36812 13932 36868
rect 13988 36812 14000 36868
rect 13920 36548 14000 36812
rect 13920 36492 13932 36548
rect 13988 36492 14000 36548
rect 13920 36480 14000 36492
rect 14080 36868 14160 36880
rect 14080 36812 14092 36868
rect 14148 36812 14160 36868
rect 14080 36548 14160 36812
rect 14080 36492 14092 36548
rect 14148 36492 14160 36548
rect 14080 36480 14160 36492
rect 14240 36868 14320 36880
rect 14240 36812 14252 36868
rect 14308 36812 14320 36868
rect 14240 36548 14320 36812
rect 14240 36492 14252 36548
rect 14308 36492 14320 36548
rect 14240 36480 14320 36492
rect 14400 36868 14480 36880
rect 14400 36812 14412 36868
rect 14468 36812 14480 36868
rect 14400 36548 14480 36812
rect 14400 36492 14412 36548
rect 14468 36492 14480 36548
rect 14400 36480 14480 36492
rect 14560 36868 14640 36880
rect 14560 36812 14572 36868
rect 14628 36812 14640 36868
rect 14560 36548 14640 36812
rect 14560 36492 14572 36548
rect 14628 36492 14640 36548
rect 14560 36480 14640 36492
rect 14720 36868 14800 36880
rect 14720 36812 14732 36868
rect 14788 36812 14800 36868
rect 14720 36548 14800 36812
rect 14720 36492 14732 36548
rect 14788 36492 14800 36548
rect 14720 36480 14800 36492
rect 14880 36868 14960 36880
rect 14880 36812 14892 36868
rect 14948 36812 14960 36868
rect 14880 36548 14960 36812
rect 14880 36492 14892 36548
rect 14948 36492 14960 36548
rect 14880 36480 14960 36492
rect 15040 36868 15120 36880
rect 15040 36812 15052 36868
rect 15108 36812 15120 36868
rect 15040 36548 15120 36812
rect 15040 36492 15052 36548
rect 15108 36492 15120 36548
rect 15040 36480 15120 36492
rect 15200 36868 15280 36880
rect 15200 36812 15212 36868
rect 15268 36812 15280 36868
rect 15200 36548 15280 36812
rect 15200 36492 15212 36548
rect 15268 36492 15280 36548
rect 15200 36480 15280 36492
rect 15360 36868 15440 36880
rect 15360 36812 15372 36868
rect 15428 36812 15440 36868
rect 15360 36548 15440 36812
rect 15360 36492 15372 36548
rect 15428 36492 15440 36548
rect 15360 36480 15440 36492
rect 15520 36868 15600 36880
rect 15520 36812 15532 36868
rect 15588 36812 15600 36868
rect 15520 36548 15600 36812
rect 15520 36492 15532 36548
rect 15588 36492 15600 36548
rect 15520 36480 15600 36492
rect 15680 36868 15760 36880
rect 15680 36812 15692 36868
rect 15748 36812 15760 36868
rect 15680 36548 15760 36812
rect 15680 36492 15692 36548
rect 15748 36492 15760 36548
rect 15680 36480 15760 36492
rect 15840 36868 15920 36880
rect 15840 36812 15852 36868
rect 15908 36812 15920 36868
rect 15840 36548 15920 36812
rect 15840 36492 15852 36548
rect 15908 36492 15920 36548
rect 15840 36480 15920 36492
rect 16000 36868 16080 36880
rect 16000 36812 16012 36868
rect 16068 36812 16080 36868
rect 16000 36548 16080 36812
rect 16000 36492 16012 36548
rect 16068 36492 16080 36548
rect 16000 36480 16080 36492
rect 16160 36868 16240 36880
rect 16160 36812 16172 36868
rect 16228 36812 16240 36868
rect 16160 36548 16240 36812
rect 16160 36492 16172 36548
rect 16228 36492 16240 36548
rect 16160 36480 16240 36492
rect 16320 36868 16400 36880
rect 16320 36812 16332 36868
rect 16388 36812 16400 36868
rect 16320 36548 16400 36812
rect 16320 36492 16332 36548
rect 16388 36492 16400 36548
rect 16320 36480 16400 36492
rect 16480 36868 16560 36880
rect 16480 36812 16492 36868
rect 16548 36812 16560 36868
rect 16480 36548 16560 36812
rect 16480 36492 16492 36548
rect 16548 36492 16560 36548
rect 16480 36480 16560 36492
rect 16640 36868 16720 36880
rect 16640 36812 16652 36868
rect 16708 36812 16720 36868
rect 16640 36548 16720 36812
rect 16640 36492 16652 36548
rect 16708 36492 16720 36548
rect 16640 36480 16720 36492
rect 16800 36868 16880 36880
rect 16800 36812 16812 36868
rect 16868 36812 16880 36868
rect 16800 36548 16880 36812
rect 16800 36492 16812 36548
rect 16868 36492 16880 36548
rect 16800 36480 16880 36492
rect 16960 36868 17040 36880
rect 16960 36812 16972 36868
rect 17028 36812 17040 36868
rect 16960 36548 17040 36812
rect 16960 36492 16972 36548
rect 17028 36492 17040 36548
rect 16960 36480 17040 36492
rect 17120 36868 17200 36880
rect 17120 36812 17132 36868
rect 17188 36812 17200 36868
rect 17120 36548 17200 36812
rect 17120 36492 17132 36548
rect 17188 36492 17200 36548
rect 17120 36480 17200 36492
rect 17280 36868 17360 36880
rect 17280 36812 17292 36868
rect 17348 36812 17360 36868
rect 17280 36548 17360 36812
rect 17280 36492 17292 36548
rect 17348 36492 17360 36548
rect 17280 36480 17360 36492
rect 17440 36868 17520 36880
rect 17440 36812 17452 36868
rect 17508 36812 17520 36868
rect 17440 36548 17520 36812
rect 17440 36492 17452 36548
rect 17508 36492 17520 36548
rect 17440 36480 17520 36492
rect 17600 36868 17680 36880
rect 17600 36812 17612 36868
rect 17668 36812 17680 36868
rect 17600 36548 17680 36812
rect 17600 36492 17612 36548
rect 17668 36492 17680 36548
rect 17600 36480 17680 36492
rect 17760 36868 17840 36880
rect 17760 36812 17772 36868
rect 17828 36812 17840 36868
rect 17760 36548 17840 36812
rect 17760 36492 17772 36548
rect 17828 36492 17840 36548
rect 17760 36480 17840 36492
rect 17920 36868 18000 36880
rect 17920 36812 17932 36868
rect 17988 36812 18000 36868
rect 17920 36548 18000 36812
rect 17920 36492 17932 36548
rect 17988 36492 18000 36548
rect 17920 36480 18000 36492
rect 18080 36868 18160 36880
rect 18080 36812 18092 36868
rect 18148 36812 18160 36868
rect 18080 36548 18160 36812
rect 18080 36492 18092 36548
rect 18148 36492 18160 36548
rect 18080 36480 18160 36492
rect 18240 36868 18320 36880
rect 18240 36812 18252 36868
rect 18308 36812 18320 36868
rect 18240 36548 18320 36812
rect 18240 36492 18252 36548
rect 18308 36492 18320 36548
rect 18240 36480 18320 36492
rect 18400 36868 18480 36880
rect 18400 36812 18412 36868
rect 18468 36812 18480 36868
rect 18400 36548 18480 36812
rect 18400 36492 18412 36548
rect 18468 36492 18480 36548
rect 18400 36480 18480 36492
rect 18560 36868 18640 36880
rect 18560 36812 18572 36868
rect 18628 36812 18640 36868
rect 18560 36548 18640 36812
rect 18560 36492 18572 36548
rect 18628 36492 18640 36548
rect 18560 36480 18640 36492
rect 18720 36868 18800 36880
rect 18720 36812 18732 36868
rect 18788 36812 18800 36868
rect 18720 36548 18800 36812
rect 18720 36492 18732 36548
rect 18788 36492 18800 36548
rect 18720 36480 18800 36492
rect 18880 36868 18960 36880
rect 18880 36812 18892 36868
rect 18948 36812 18960 36868
rect 18880 36548 18960 36812
rect 18880 36492 18892 36548
rect 18948 36492 18960 36548
rect 18880 36480 18960 36492
rect 12480 36388 12560 36400
rect 12480 36332 12492 36388
rect 12548 36332 12560 36388
rect 12480 36068 12560 36332
rect 12480 36012 12492 36068
rect 12548 36012 12560 36068
rect 12480 35748 12560 36012
rect 12480 35692 12492 35748
rect 12548 35692 12560 35748
rect 12480 35428 12560 35692
rect 12480 35372 12492 35428
rect 12548 35372 12560 35428
rect 12480 35108 12560 35372
rect 12480 35052 12492 35108
rect 12548 35052 12560 35108
rect 12480 34788 12560 35052
rect 12480 34732 12492 34788
rect 12548 34732 12560 34788
rect 12480 34468 12560 34732
rect 12480 34412 12492 34468
rect 12548 34412 12560 34468
rect 12480 34400 12560 34412
rect 12640 36388 12720 36400
rect 12640 36332 12652 36388
rect 12708 36332 12720 36388
rect 12640 36068 12720 36332
rect 12640 36012 12652 36068
rect 12708 36012 12720 36068
rect 12640 35748 12720 36012
rect 12640 35692 12652 35748
rect 12708 35692 12720 35748
rect 12640 35428 12720 35692
rect 12640 35372 12652 35428
rect 12708 35372 12720 35428
rect 12640 35108 12720 35372
rect 12640 35052 12652 35108
rect 12708 35052 12720 35108
rect 12640 34788 12720 35052
rect 12640 34732 12652 34788
rect 12708 34732 12720 34788
rect 12640 34468 12720 34732
rect 12640 34412 12652 34468
rect 12708 34412 12720 34468
rect 12640 34400 12720 34412
rect 12800 36388 12880 36400
rect 12800 36332 12812 36388
rect 12868 36332 12880 36388
rect 12800 36068 12880 36332
rect 12800 36012 12812 36068
rect 12868 36012 12880 36068
rect 12800 35748 12880 36012
rect 12800 35692 12812 35748
rect 12868 35692 12880 35748
rect 12800 35428 12880 35692
rect 12800 35372 12812 35428
rect 12868 35372 12880 35428
rect 12800 35108 12880 35372
rect 12800 35052 12812 35108
rect 12868 35052 12880 35108
rect 12800 34788 12880 35052
rect 12800 34732 12812 34788
rect 12868 34732 12880 34788
rect 12800 34468 12880 34732
rect 12800 34412 12812 34468
rect 12868 34412 12880 34468
rect 12800 34400 12880 34412
rect 12960 36388 13040 36400
rect 12960 36332 12972 36388
rect 13028 36332 13040 36388
rect 12960 36068 13040 36332
rect 12960 36012 12972 36068
rect 13028 36012 13040 36068
rect 12960 35748 13040 36012
rect 12960 35692 12972 35748
rect 13028 35692 13040 35748
rect 12960 35428 13040 35692
rect 12960 35372 12972 35428
rect 13028 35372 13040 35428
rect 12960 35108 13040 35372
rect 12960 35052 12972 35108
rect 13028 35052 13040 35108
rect 12960 34788 13040 35052
rect 12960 34732 12972 34788
rect 13028 34732 13040 34788
rect 12960 34468 13040 34732
rect 12960 34412 12972 34468
rect 13028 34412 13040 34468
rect 12960 34400 13040 34412
rect 13120 36388 13200 36400
rect 13120 36332 13132 36388
rect 13188 36332 13200 36388
rect 13120 36068 13200 36332
rect 13120 36012 13132 36068
rect 13188 36012 13200 36068
rect 13120 35748 13200 36012
rect 13120 35692 13132 35748
rect 13188 35692 13200 35748
rect 13120 35428 13200 35692
rect 13120 35372 13132 35428
rect 13188 35372 13200 35428
rect 13120 35108 13200 35372
rect 13120 35052 13132 35108
rect 13188 35052 13200 35108
rect 13120 34788 13200 35052
rect 13120 34732 13132 34788
rect 13188 34732 13200 34788
rect 13120 34468 13200 34732
rect 13120 34412 13132 34468
rect 13188 34412 13200 34468
rect 13120 34400 13200 34412
rect 13280 36388 13360 36400
rect 13280 36332 13292 36388
rect 13348 36332 13360 36388
rect 13280 36068 13360 36332
rect 13280 36012 13292 36068
rect 13348 36012 13360 36068
rect 13280 35748 13360 36012
rect 13280 35692 13292 35748
rect 13348 35692 13360 35748
rect 13280 35428 13360 35692
rect 13280 35372 13292 35428
rect 13348 35372 13360 35428
rect 13280 35108 13360 35372
rect 13280 35052 13292 35108
rect 13348 35052 13360 35108
rect 13280 34788 13360 35052
rect 13280 34732 13292 34788
rect 13348 34732 13360 34788
rect 13280 34468 13360 34732
rect 13280 34412 13292 34468
rect 13348 34412 13360 34468
rect 13280 34400 13360 34412
rect 13440 36388 13520 36400
rect 13440 36332 13452 36388
rect 13508 36332 13520 36388
rect 13440 36068 13520 36332
rect 13440 36012 13452 36068
rect 13508 36012 13520 36068
rect 13440 35748 13520 36012
rect 13440 35692 13452 35748
rect 13508 35692 13520 35748
rect 13440 35428 13520 35692
rect 13440 35372 13452 35428
rect 13508 35372 13520 35428
rect 13440 35108 13520 35372
rect 13440 35052 13452 35108
rect 13508 35052 13520 35108
rect 13440 34788 13520 35052
rect 13440 34732 13452 34788
rect 13508 34732 13520 34788
rect 13440 34468 13520 34732
rect 13440 34412 13452 34468
rect 13508 34412 13520 34468
rect 13440 34400 13520 34412
rect 13600 36388 13680 36400
rect 13600 36332 13612 36388
rect 13668 36332 13680 36388
rect 13600 36068 13680 36332
rect 13600 36012 13612 36068
rect 13668 36012 13680 36068
rect 13600 35748 13680 36012
rect 13600 35692 13612 35748
rect 13668 35692 13680 35748
rect 13600 35428 13680 35692
rect 13600 35372 13612 35428
rect 13668 35372 13680 35428
rect 13600 35108 13680 35372
rect 13600 35052 13612 35108
rect 13668 35052 13680 35108
rect 13600 34788 13680 35052
rect 13600 34732 13612 34788
rect 13668 34732 13680 34788
rect 13600 34468 13680 34732
rect 13600 34412 13612 34468
rect 13668 34412 13680 34468
rect 13600 34400 13680 34412
rect 13760 36388 13840 36400
rect 13760 36332 13772 36388
rect 13828 36332 13840 36388
rect 13760 36068 13840 36332
rect 13760 36012 13772 36068
rect 13828 36012 13840 36068
rect 13760 35748 13840 36012
rect 13760 35692 13772 35748
rect 13828 35692 13840 35748
rect 13760 35428 13840 35692
rect 13760 35372 13772 35428
rect 13828 35372 13840 35428
rect 13760 35108 13840 35372
rect 13760 35052 13772 35108
rect 13828 35052 13840 35108
rect 13760 34788 13840 35052
rect 13760 34732 13772 34788
rect 13828 34732 13840 34788
rect 13760 34468 13840 34732
rect 13760 34412 13772 34468
rect 13828 34412 13840 34468
rect 13760 34400 13840 34412
rect 13920 36388 14000 36400
rect 13920 36332 13932 36388
rect 13988 36332 14000 36388
rect 13920 36068 14000 36332
rect 13920 36012 13932 36068
rect 13988 36012 14000 36068
rect 13920 35748 14000 36012
rect 13920 35692 13932 35748
rect 13988 35692 14000 35748
rect 13920 35428 14000 35692
rect 13920 35372 13932 35428
rect 13988 35372 14000 35428
rect 13920 35108 14000 35372
rect 13920 35052 13932 35108
rect 13988 35052 14000 35108
rect 13920 34788 14000 35052
rect 13920 34732 13932 34788
rect 13988 34732 14000 34788
rect 13920 34468 14000 34732
rect 13920 34412 13932 34468
rect 13988 34412 14000 34468
rect 13920 34400 14000 34412
rect 14080 36388 14160 36400
rect 14080 36332 14092 36388
rect 14148 36332 14160 36388
rect 14080 36068 14160 36332
rect 14080 36012 14092 36068
rect 14148 36012 14160 36068
rect 14080 35748 14160 36012
rect 14080 35692 14092 35748
rect 14148 35692 14160 35748
rect 14080 35428 14160 35692
rect 14080 35372 14092 35428
rect 14148 35372 14160 35428
rect 14080 35108 14160 35372
rect 14080 35052 14092 35108
rect 14148 35052 14160 35108
rect 14080 34788 14160 35052
rect 14080 34732 14092 34788
rect 14148 34732 14160 34788
rect 14080 34468 14160 34732
rect 14080 34412 14092 34468
rect 14148 34412 14160 34468
rect 14080 34400 14160 34412
rect 14240 36388 14320 36400
rect 14240 36332 14252 36388
rect 14308 36332 14320 36388
rect 14240 36068 14320 36332
rect 14240 36012 14252 36068
rect 14308 36012 14320 36068
rect 14240 35748 14320 36012
rect 14240 35692 14252 35748
rect 14308 35692 14320 35748
rect 14240 35428 14320 35692
rect 14240 35372 14252 35428
rect 14308 35372 14320 35428
rect 14240 35108 14320 35372
rect 14240 35052 14252 35108
rect 14308 35052 14320 35108
rect 14240 34788 14320 35052
rect 14240 34732 14252 34788
rect 14308 34732 14320 34788
rect 14240 34468 14320 34732
rect 14240 34412 14252 34468
rect 14308 34412 14320 34468
rect 14240 34400 14320 34412
rect 14400 36388 14480 36400
rect 14400 36332 14412 36388
rect 14468 36332 14480 36388
rect 14400 36068 14480 36332
rect 14400 36012 14412 36068
rect 14468 36012 14480 36068
rect 14400 35748 14480 36012
rect 14400 35692 14412 35748
rect 14468 35692 14480 35748
rect 14400 35428 14480 35692
rect 14400 35372 14412 35428
rect 14468 35372 14480 35428
rect 14400 35108 14480 35372
rect 14400 35052 14412 35108
rect 14468 35052 14480 35108
rect 14400 34788 14480 35052
rect 14400 34732 14412 34788
rect 14468 34732 14480 34788
rect 14400 34468 14480 34732
rect 14400 34412 14412 34468
rect 14468 34412 14480 34468
rect 14400 34400 14480 34412
rect 14560 36388 14640 36400
rect 14560 36332 14572 36388
rect 14628 36332 14640 36388
rect 14560 36068 14640 36332
rect 14560 36012 14572 36068
rect 14628 36012 14640 36068
rect 14560 35748 14640 36012
rect 14560 35692 14572 35748
rect 14628 35692 14640 35748
rect 14560 35428 14640 35692
rect 14560 35372 14572 35428
rect 14628 35372 14640 35428
rect 14560 35108 14640 35372
rect 14560 35052 14572 35108
rect 14628 35052 14640 35108
rect 14560 34788 14640 35052
rect 14560 34732 14572 34788
rect 14628 34732 14640 34788
rect 14560 34468 14640 34732
rect 14560 34412 14572 34468
rect 14628 34412 14640 34468
rect 14560 34400 14640 34412
rect 14720 36388 14800 36400
rect 14720 36332 14732 36388
rect 14788 36332 14800 36388
rect 14720 36068 14800 36332
rect 14720 36012 14732 36068
rect 14788 36012 14800 36068
rect 14720 35748 14800 36012
rect 14720 35692 14732 35748
rect 14788 35692 14800 35748
rect 14720 35428 14800 35692
rect 14720 35372 14732 35428
rect 14788 35372 14800 35428
rect 14720 35108 14800 35372
rect 14720 35052 14732 35108
rect 14788 35052 14800 35108
rect 14720 34788 14800 35052
rect 14720 34732 14732 34788
rect 14788 34732 14800 34788
rect 14720 34468 14800 34732
rect 14720 34412 14732 34468
rect 14788 34412 14800 34468
rect 14720 34400 14800 34412
rect 14880 36388 14960 36400
rect 14880 36332 14892 36388
rect 14948 36332 14960 36388
rect 14880 36068 14960 36332
rect 14880 36012 14892 36068
rect 14948 36012 14960 36068
rect 14880 35748 14960 36012
rect 14880 35692 14892 35748
rect 14948 35692 14960 35748
rect 14880 35428 14960 35692
rect 14880 35372 14892 35428
rect 14948 35372 14960 35428
rect 14880 35108 14960 35372
rect 14880 35052 14892 35108
rect 14948 35052 14960 35108
rect 14880 34788 14960 35052
rect 14880 34732 14892 34788
rect 14948 34732 14960 34788
rect 14880 34468 14960 34732
rect 14880 34412 14892 34468
rect 14948 34412 14960 34468
rect 14880 34400 14960 34412
rect 15040 36388 15120 36400
rect 15040 36332 15052 36388
rect 15108 36332 15120 36388
rect 15040 36068 15120 36332
rect 15040 36012 15052 36068
rect 15108 36012 15120 36068
rect 15040 35748 15120 36012
rect 15040 35692 15052 35748
rect 15108 35692 15120 35748
rect 15040 35428 15120 35692
rect 15040 35372 15052 35428
rect 15108 35372 15120 35428
rect 15040 35108 15120 35372
rect 15040 35052 15052 35108
rect 15108 35052 15120 35108
rect 15040 34788 15120 35052
rect 15040 34732 15052 34788
rect 15108 34732 15120 34788
rect 15040 34468 15120 34732
rect 15040 34412 15052 34468
rect 15108 34412 15120 34468
rect 15040 34400 15120 34412
rect 15200 36388 15280 36400
rect 15200 36332 15212 36388
rect 15268 36332 15280 36388
rect 15200 36068 15280 36332
rect 15200 36012 15212 36068
rect 15268 36012 15280 36068
rect 15200 35748 15280 36012
rect 15200 35692 15212 35748
rect 15268 35692 15280 35748
rect 15200 35428 15280 35692
rect 15200 35372 15212 35428
rect 15268 35372 15280 35428
rect 15200 35108 15280 35372
rect 15200 35052 15212 35108
rect 15268 35052 15280 35108
rect 15200 34788 15280 35052
rect 15200 34732 15212 34788
rect 15268 34732 15280 34788
rect 15200 34468 15280 34732
rect 15200 34412 15212 34468
rect 15268 34412 15280 34468
rect 15200 34400 15280 34412
rect 15360 36388 15440 36400
rect 15360 36332 15372 36388
rect 15428 36332 15440 36388
rect 15360 36068 15440 36332
rect 15360 36012 15372 36068
rect 15428 36012 15440 36068
rect 15360 35748 15440 36012
rect 15360 35692 15372 35748
rect 15428 35692 15440 35748
rect 15360 35428 15440 35692
rect 15360 35372 15372 35428
rect 15428 35372 15440 35428
rect 15360 35108 15440 35372
rect 15360 35052 15372 35108
rect 15428 35052 15440 35108
rect 15360 34788 15440 35052
rect 15360 34732 15372 34788
rect 15428 34732 15440 34788
rect 15360 34468 15440 34732
rect 15360 34412 15372 34468
rect 15428 34412 15440 34468
rect 15360 34400 15440 34412
rect 15520 36388 15600 36400
rect 15520 36332 15532 36388
rect 15588 36332 15600 36388
rect 15520 36068 15600 36332
rect 15520 36012 15532 36068
rect 15588 36012 15600 36068
rect 15520 35748 15600 36012
rect 15520 35692 15532 35748
rect 15588 35692 15600 35748
rect 15520 35428 15600 35692
rect 15520 35372 15532 35428
rect 15588 35372 15600 35428
rect 15520 35108 15600 35372
rect 15520 35052 15532 35108
rect 15588 35052 15600 35108
rect 15520 34788 15600 35052
rect 15520 34732 15532 34788
rect 15588 34732 15600 34788
rect 15520 34468 15600 34732
rect 15520 34412 15532 34468
rect 15588 34412 15600 34468
rect 15520 34400 15600 34412
rect 15680 36388 15760 36400
rect 15680 36332 15692 36388
rect 15748 36332 15760 36388
rect 15680 36068 15760 36332
rect 15680 36012 15692 36068
rect 15748 36012 15760 36068
rect 15680 35748 15760 36012
rect 15680 35692 15692 35748
rect 15748 35692 15760 35748
rect 15680 35428 15760 35692
rect 15680 35372 15692 35428
rect 15748 35372 15760 35428
rect 15680 35108 15760 35372
rect 15680 35052 15692 35108
rect 15748 35052 15760 35108
rect 15680 34788 15760 35052
rect 15680 34732 15692 34788
rect 15748 34732 15760 34788
rect 15680 34468 15760 34732
rect 15680 34412 15692 34468
rect 15748 34412 15760 34468
rect 15680 34400 15760 34412
rect 15840 36388 15920 36400
rect 15840 36332 15852 36388
rect 15908 36332 15920 36388
rect 15840 36068 15920 36332
rect 15840 36012 15852 36068
rect 15908 36012 15920 36068
rect 15840 35748 15920 36012
rect 15840 35692 15852 35748
rect 15908 35692 15920 35748
rect 15840 35428 15920 35692
rect 15840 35372 15852 35428
rect 15908 35372 15920 35428
rect 15840 35108 15920 35372
rect 15840 35052 15852 35108
rect 15908 35052 15920 35108
rect 15840 34788 15920 35052
rect 15840 34732 15852 34788
rect 15908 34732 15920 34788
rect 15840 34468 15920 34732
rect 15840 34412 15852 34468
rect 15908 34412 15920 34468
rect 15840 34400 15920 34412
rect 16000 36388 16080 36400
rect 16000 36332 16012 36388
rect 16068 36332 16080 36388
rect 16000 36068 16080 36332
rect 16000 36012 16012 36068
rect 16068 36012 16080 36068
rect 16000 35748 16080 36012
rect 16000 35692 16012 35748
rect 16068 35692 16080 35748
rect 16000 35428 16080 35692
rect 16000 35372 16012 35428
rect 16068 35372 16080 35428
rect 16000 35108 16080 35372
rect 16000 35052 16012 35108
rect 16068 35052 16080 35108
rect 16000 34788 16080 35052
rect 16000 34732 16012 34788
rect 16068 34732 16080 34788
rect 16000 34468 16080 34732
rect 16000 34412 16012 34468
rect 16068 34412 16080 34468
rect 16000 34400 16080 34412
rect 16160 36388 16240 36400
rect 16160 36332 16172 36388
rect 16228 36332 16240 36388
rect 16160 36068 16240 36332
rect 16160 36012 16172 36068
rect 16228 36012 16240 36068
rect 16160 35748 16240 36012
rect 16160 35692 16172 35748
rect 16228 35692 16240 35748
rect 16160 35428 16240 35692
rect 16160 35372 16172 35428
rect 16228 35372 16240 35428
rect 16160 35108 16240 35372
rect 16160 35052 16172 35108
rect 16228 35052 16240 35108
rect 16160 34788 16240 35052
rect 16160 34732 16172 34788
rect 16228 34732 16240 34788
rect 16160 34468 16240 34732
rect 16160 34412 16172 34468
rect 16228 34412 16240 34468
rect 16160 34400 16240 34412
rect 16320 36388 16400 36400
rect 16320 36332 16332 36388
rect 16388 36332 16400 36388
rect 16320 36068 16400 36332
rect 16320 36012 16332 36068
rect 16388 36012 16400 36068
rect 16320 35748 16400 36012
rect 16320 35692 16332 35748
rect 16388 35692 16400 35748
rect 16320 35428 16400 35692
rect 16320 35372 16332 35428
rect 16388 35372 16400 35428
rect 16320 35108 16400 35372
rect 16320 35052 16332 35108
rect 16388 35052 16400 35108
rect 16320 34788 16400 35052
rect 16320 34732 16332 34788
rect 16388 34732 16400 34788
rect 16320 34468 16400 34732
rect 16320 34412 16332 34468
rect 16388 34412 16400 34468
rect 16320 34400 16400 34412
rect 16480 36388 16560 36400
rect 16480 36332 16492 36388
rect 16548 36332 16560 36388
rect 16480 36068 16560 36332
rect 16480 36012 16492 36068
rect 16548 36012 16560 36068
rect 16480 35748 16560 36012
rect 16480 35692 16492 35748
rect 16548 35692 16560 35748
rect 16480 35428 16560 35692
rect 16480 35372 16492 35428
rect 16548 35372 16560 35428
rect 16480 35108 16560 35372
rect 16480 35052 16492 35108
rect 16548 35052 16560 35108
rect 16480 34788 16560 35052
rect 16480 34732 16492 34788
rect 16548 34732 16560 34788
rect 16480 34468 16560 34732
rect 16480 34412 16492 34468
rect 16548 34412 16560 34468
rect 16480 34400 16560 34412
rect 16640 36388 16720 36400
rect 16640 36332 16652 36388
rect 16708 36332 16720 36388
rect 16640 36068 16720 36332
rect 16640 36012 16652 36068
rect 16708 36012 16720 36068
rect 16640 35748 16720 36012
rect 16640 35692 16652 35748
rect 16708 35692 16720 35748
rect 16640 35428 16720 35692
rect 16640 35372 16652 35428
rect 16708 35372 16720 35428
rect 16640 35108 16720 35372
rect 16640 35052 16652 35108
rect 16708 35052 16720 35108
rect 16640 34788 16720 35052
rect 16640 34732 16652 34788
rect 16708 34732 16720 34788
rect 16640 34468 16720 34732
rect 16640 34412 16652 34468
rect 16708 34412 16720 34468
rect 16640 34400 16720 34412
rect 16800 36388 16880 36400
rect 16800 36332 16812 36388
rect 16868 36332 16880 36388
rect 16800 36068 16880 36332
rect 16800 36012 16812 36068
rect 16868 36012 16880 36068
rect 16800 35748 16880 36012
rect 16800 35692 16812 35748
rect 16868 35692 16880 35748
rect 16800 35428 16880 35692
rect 16800 35372 16812 35428
rect 16868 35372 16880 35428
rect 16800 35108 16880 35372
rect 16800 35052 16812 35108
rect 16868 35052 16880 35108
rect 16800 34788 16880 35052
rect 16800 34732 16812 34788
rect 16868 34732 16880 34788
rect 16800 34468 16880 34732
rect 16800 34412 16812 34468
rect 16868 34412 16880 34468
rect 16800 34400 16880 34412
rect 16960 36388 17040 36400
rect 16960 36332 16972 36388
rect 17028 36332 17040 36388
rect 16960 36068 17040 36332
rect 16960 36012 16972 36068
rect 17028 36012 17040 36068
rect 16960 35748 17040 36012
rect 16960 35692 16972 35748
rect 17028 35692 17040 35748
rect 16960 35428 17040 35692
rect 16960 35372 16972 35428
rect 17028 35372 17040 35428
rect 16960 35108 17040 35372
rect 16960 35052 16972 35108
rect 17028 35052 17040 35108
rect 16960 34788 17040 35052
rect 16960 34732 16972 34788
rect 17028 34732 17040 34788
rect 16960 34468 17040 34732
rect 16960 34412 16972 34468
rect 17028 34412 17040 34468
rect 16960 34400 17040 34412
rect 17120 36388 17200 36400
rect 17120 36332 17132 36388
rect 17188 36332 17200 36388
rect 17120 36068 17200 36332
rect 17120 36012 17132 36068
rect 17188 36012 17200 36068
rect 17120 35748 17200 36012
rect 17120 35692 17132 35748
rect 17188 35692 17200 35748
rect 17120 35428 17200 35692
rect 17120 35372 17132 35428
rect 17188 35372 17200 35428
rect 17120 35108 17200 35372
rect 17120 35052 17132 35108
rect 17188 35052 17200 35108
rect 17120 34788 17200 35052
rect 17120 34732 17132 34788
rect 17188 34732 17200 34788
rect 17120 34468 17200 34732
rect 17120 34412 17132 34468
rect 17188 34412 17200 34468
rect 17120 34400 17200 34412
rect 17280 36388 17360 36400
rect 17280 36332 17292 36388
rect 17348 36332 17360 36388
rect 17280 36068 17360 36332
rect 17280 36012 17292 36068
rect 17348 36012 17360 36068
rect 17280 35748 17360 36012
rect 17280 35692 17292 35748
rect 17348 35692 17360 35748
rect 17280 35428 17360 35692
rect 17280 35372 17292 35428
rect 17348 35372 17360 35428
rect 17280 35108 17360 35372
rect 17280 35052 17292 35108
rect 17348 35052 17360 35108
rect 17280 34788 17360 35052
rect 17280 34732 17292 34788
rect 17348 34732 17360 34788
rect 17280 34468 17360 34732
rect 17280 34412 17292 34468
rect 17348 34412 17360 34468
rect 17280 34400 17360 34412
rect 17440 36388 17520 36400
rect 17440 36332 17452 36388
rect 17508 36332 17520 36388
rect 17440 36068 17520 36332
rect 17440 36012 17452 36068
rect 17508 36012 17520 36068
rect 17440 35748 17520 36012
rect 17440 35692 17452 35748
rect 17508 35692 17520 35748
rect 17440 35428 17520 35692
rect 17440 35372 17452 35428
rect 17508 35372 17520 35428
rect 17440 35108 17520 35372
rect 17440 35052 17452 35108
rect 17508 35052 17520 35108
rect 17440 34788 17520 35052
rect 17440 34732 17452 34788
rect 17508 34732 17520 34788
rect 17440 34468 17520 34732
rect 17440 34412 17452 34468
rect 17508 34412 17520 34468
rect 17440 34400 17520 34412
rect 17600 36388 17680 36400
rect 17600 36332 17612 36388
rect 17668 36332 17680 36388
rect 17600 36068 17680 36332
rect 17600 36012 17612 36068
rect 17668 36012 17680 36068
rect 17600 35748 17680 36012
rect 17600 35692 17612 35748
rect 17668 35692 17680 35748
rect 17600 35428 17680 35692
rect 17600 35372 17612 35428
rect 17668 35372 17680 35428
rect 17600 35108 17680 35372
rect 17600 35052 17612 35108
rect 17668 35052 17680 35108
rect 17600 34788 17680 35052
rect 17600 34732 17612 34788
rect 17668 34732 17680 34788
rect 17600 34468 17680 34732
rect 17600 34412 17612 34468
rect 17668 34412 17680 34468
rect 17600 34400 17680 34412
rect 17760 36388 17840 36400
rect 17760 36332 17772 36388
rect 17828 36332 17840 36388
rect 17760 36068 17840 36332
rect 17760 36012 17772 36068
rect 17828 36012 17840 36068
rect 17760 35748 17840 36012
rect 17760 35692 17772 35748
rect 17828 35692 17840 35748
rect 17760 35428 17840 35692
rect 17760 35372 17772 35428
rect 17828 35372 17840 35428
rect 17760 35108 17840 35372
rect 17760 35052 17772 35108
rect 17828 35052 17840 35108
rect 17760 34788 17840 35052
rect 17760 34732 17772 34788
rect 17828 34732 17840 34788
rect 17760 34468 17840 34732
rect 17760 34412 17772 34468
rect 17828 34412 17840 34468
rect 17760 34400 17840 34412
rect 17920 36388 18000 36400
rect 17920 36332 17932 36388
rect 17988 36332 18000 36388
rect 17920 36068 18000 36332
rect 17920 36012 17932 36068
rect 17988 36012 18000 36068
rect 17920 35748 18000 36012
rect 17920 35692 17932 35748
rect 17988 35692 18000 35748
rect 17920 35428 18000 35692
rect 17920 35372 17932 35428
rect 17988 35372 18000 35428
rect 17920 35108 18000 35372
rect 17920 35052 17932 35108
rect 17988 35052 18000 35108
rect 17920 34788 18000 35052
rect 17920 34732 17932 34788
rect 17988 34732 18000 34788
rect 17920 34468 18000 34732
rect 17920 34412 17932 34468
rect 17988 34412 18000 34468
rect 17920 34400 18000 34412
rect 18080 36388 18160 36400
rect 18080 36332 18092 36388
rect 18148 36332 18160 36388
rect 18080 36068 18160 36332
rect 18080 36012 18092 36068
rect 18148 36012 18160 36068
rect 18080 35748 18160 36012
rect 18080 35692 18092 35748
rect 18148 35692 18160 35748
rect 18080 35428 18160 35692
rect 18080 35372 18092 35428
rect 18148 35372 18160 35428
rect 18080 35108 18160 35372
rect 18080 35052 18092 35108
rect 18148 35052 18160 35108
rect 18080 34788 18160 35052
rect 18080 34732 18092 34788
rect 18148 34732 18160 34788
rect 18080 34468 18160 34732
rect 18080 34412 18092 34468
rect 18148 34412 18160 34468
rect 18080 34400 18160 34412
rect 18240 36388 18320 36400
rect 18240 36332 18252 36388
rect 18308 36332 18320 36388
rect 18240 36068 18320 36332
rect 18240 36012 18252 36068
rect 18308 36012 18320 36068
rect 18240 35748 18320 36012
rect 18240 35692 18252 35748
rect 18308 35692 18320 35748
rect 18240 35428 18320 35692
rect 18240 35372 18252 35428
rect 18308 35372 18320 35428
rect 18240 35108 18320 35372
rect 18240 35052 18252 35108
rect 18308 35052 18320 35108
rect 18240 34788 18320 35052
rect 18240 34732 18252 34788
rect 18308 34732 18320 34788
rect 18240 34468 18320 34732
rect 18240 34412 18252 34468
rect 18308 34412 18320 34468
rect 18240 34400 18320 34412
rect 18400 36388 18480 36400
rect 18400 36332 18412 36388
rect 18468 36332 18480 36388
rect 18400 36068 18480 36332
rect 18400 36012 18412 36068
rect 18468 36012 18480 36068
rect 18400 35748 18480 36012
rect 18400 35692 18412 35748
rect 18468 35692 18480 35748
rect 18400 35428 18480 35692
rect 18400 35372 18412 35428
rect 18468 35372 18480 35428
rect 18400 35108 18480 35372
rect 18400 35052 18412 35108
rect 18468 35052 18480 35108
rect 18400 34788 18480 35052
rect 18400 34732 18412 34788
rect 18468 34732 18480 34788
rect 18400 34468 18480 34732
rect 18400 34412 18412 34468
rect 18468 34412 18480 34468
rect 18400 34400 18480 34412
rect 18560 36388 18640 36400
rect 18560 36332 18572 36388
rect 18628 36332 18640 36388
rect 18560 36068 18640 36332
rect 18560 36012 18572 36068
rect 18628 36012 18640 36068
rect 18560 35748 18640 36012
rect 18560 35692 18572 35748
rect 18628 35692 18640 35748
rect 18560 35428 18640 35692
rect 18560 35372 18572 35428
rect 18628 35372 18640 35428
rect 18560 35108 18640 35372
rect 18560 35052 18572 35108
rect 18628 35052 18640 35108
rect 18560 34788 18640 35052
rect 18560 34732 18572 34788
rect 18628 34732 18640 34788
rect 18560 34468 18640 34732
rect 18560 34412 18572 34468
rect 18628 34412 18640 34468
rect 18560 34400 18640 34412
rect 18720 36388 18800 36400
rect 18720 36332 18732 36388
rect 18788 36332 18800 36388
rect 18720 36068 18800 36332
rect 18720 36012 18732 36068
rect 18788 36012 18800 36068
rect 18720 35748 18800 36012
rect 18720 35692 18732 35748
rect 18788 35692 18800 35748
rect 18720 35428 18800 35692
rect 18720 35372 18732 35428
rect 18788 35372 18800 35428
rect 18720 35108 18800 35372
rect 18720 35052 18732 35108
rect 18788 35052 18800 35108
rect 18720 34788 18800 35052
rect 18720 34732 18732 34788
rect 18788 34732 18800 34788
rect 18720 34468 18800 34732
rect 18720 34412 18732 34468
rect 18788 34412 18800 34468
rect 18720 34400 18800 34412
rect 18880 36388 18960 36400
rect 18880 36332 18892 36388
rect 18948 36332 18960 36388
rect 18880 36068 18960 36332
rect 18880 36012 18892 36068
rect 18948 36012 18960 36068
rect 18880 35748 18960 36012
rect 18880 35692 18892 35748
rect 18948 35692 18960 35748
rect 18880 35428 18960 35692
rect 18880 35372 18892 35428
rect 18948 35372 18960 35428
rect 18880 35108 18960 35372
rect 18880 35052 18892 35108
rect 18948 35052 18960 35108
rect 18880 34788 18960 35052
rect 18880 34732 18892 34788
rect 18948 34732 18960 34788
rect 18880 34468 18960 34732
rect 18880 34412 18892 34468
rect 18948 34412 18960 34468
rect 18880 34400 18960 34412
rect 12480 34308 12560 34320
rect 12480 34252 12492 34308
rect 12548 34252 12560 34308
rect 12480 33988 12560 34252
rect 12480 33932 12492 33988
rect 12548 33932 12560 33988
rect 12480 33920 12560 33932
rect 12640 34308 12720 34320
rect 12640 34252 12652 34308
rect 12708 34252 12720 34308
rect 12640 33988 12720 34252
rect 12640 33932 12652 33988
rect 12708 33932 12720 33988
rect 12640 33920 12720 33932
rect 12800 34308 12880 34320
rect 12800 34252 12812 34308
rect 12868 34252 12880 34308
rect 12800 33988 12880 34252
rect 12800 33932 12812 33988
rect 12868 33932 12880 33988
rect 12800 33920 12880 33932
rect 12960 34308 13040 34320
rect 12960 34252 12972 34308
rect 13028 34252 13040 34308
rect 12960 33988 13040 34252
rect 12960 33932 12972 33988
rect 13028 33932 13040 33988
rect 12960 33920 13040 33932
rect 13120 34308 13200 34320
rect 13120 34252 13132 34308
rect 13188 34252 13200 34308
rect 13120 33988 13200 34252
rect 13120 33932 13132 33988
rect 13188 33932 13200 33988
rect 13120 33920 13200 33932
rect 13280 34308 13360 34320
rect 13280 34252 13292 34308
rect 13348 34252 13360 34308
rect 13280 33988 13360 34252
rect 13280 33932 13292 33988
rect 13348 33932 13360 33988
rect 13280 33920 13360 33932
rect 13440 34308 13520 34320
rect 13440 34252 13452 34308
rect 13508 34252 13520 34308
rect 13440 33988 13520 34252
rect 13440 33932 13452 33988
rect 13508 33932 13520 33988
rect 13440 33920 13520 33932
rect 13600 34308 13680 34320
rect 13600 34252 13612 34308
rect 13668 34252 13680 34308
rect 13600 33988 13680 34252
rect 13600 33932 13612 33988
rect 13668 33932 13680 33988
rect 13600 33920 13680 33932
rect 13760 34308 13840 34320
rect 13760 34252 13772 34308
rect 13828 34252 13840 34308
rect 13760 33988 13840 34252
rect 13760 33932 13772 33988
rect 13828 33932 13840 33988
rect 13760 33920 13840 33932
rect 13920 34308 14000 34320
rect 13920 34252 13932 34308
rect 13988 34252 14000 34308
rect 13920 33988 14000 34252
rect 13920 33932 13932 33988
rect 13988 33932 14000 33988
rect 13920 33920 14000 33932
rect 14080 34308 14160 34320
rect 14080 34252 14092 34308
rect 14148 34252 14160 34308
rect 14080 33988 14160 34252
rect 14080 33932 14092 33988
rect 14148 33932 14160 33988
rect 14080 33920 14160 33932
rect 14240 34308 14320 34320
rect 14240 34252 14252 34308
rect 14308 34252 14320 34308
rect 14240 33988 14320 34252
rect 14240 33932 14252 33988
rect 14308 33932 14320 33988
rect 14240 33920 14320 33932
rect 14400 34308 14480 34320
rect 14400 34252 14412 34308
rect 14468 34252 14480 34308
rect 14400 33988 14480 34252
rect 14400 33932 14412 33988
rect 14468 33932 14480 33988
rect 14400 33920 14480 33932
rect 14560 34308 14640 34320
rect 14560 34252 14572 34308
rect 14628 34252 14640 34308
rect 14560 33988 14640 34252
rect 14560 33932 14572 33988
rect 14628 33932 14640 33988
rect 14560 33920 14640 33932
rect 14720 34308 14800 34320
rect 14720 34252 14732 34308
rect 14788 34252 14800 34308
rect 14720 33988 14800 34252
rect 14720 33932 14732 33988
rect 14788 33932 14800 33988
rect 14720 33920 14800 33932
rect 14880 34308 14960 34320
rect 14880 34252 14892 34308
rect 14948 34252 14960 34308
rect 14880 33988 14960 34252
rect 14880 33932 14892 33988
rect 14948 33932 14960 33988
rect 14880 33920 14960 33932
rect 15040 34308 15120 34320
rect 15040 34252 15052 34308
rect 15108 34252 15120 34308
rect 15040 33988 15120 34252
rect 15040 33932 15052 33988
rect 15108 33932 15120 33988
rect 15040 33920 15120 33932
rect 15200 34308 15280 34320
rect 15200 34252 15212 34308
rect 15268 34252 15280 34308
rect 15200 33988 15280 34252
rect 15200 33932 15212 33988
rect 15268 33932 15280 33988
rect 15200 33920 15280 33932
rect 15360 34308 15440 34320
rect 15360 34252 15372 34308
rect 15428 34252 15440 34308
rect 15360 33988 15440 34252
rect 15360 33932 15372 33988
rect 15428 33932 15440 33988
rect 15360 33920 15440 33932
rect 15520 34308 15600 34320
rect 15520 34252 15532 34308
rect 15588 34252 15600 34308
rect 15520 33988 15600 34252
rect 15520 33932 15532 33988
rect 15588 33932 15600 33988
rect 15520 33920 15600 33932
rect 15680 34308 15760 34320
rect 15680 34252 15692 34308
rect 15748 34252 15760 34308
rect 15680 33988 15760 34252
rect 15680 33932 15692 33988
rect 15748 33932 15760 33988
rect 15680 33920 15760 33932
rect 15840 34308 15920 34320
rect 15840 34252 15852 34308
rect 15908 34252 15920 34308
rect 15840 33988 15920 34252
rect 15840 33932 15852 33988
rect 15908 33932 15920 33988
rect 15840 33920 15920 33932
rect 16000 34308 16080 34320
rect 16000 34252 16012 34308
rect 16068 34252 16080 34308
rect 16000 33988 16080 34252
rect 16000 33932 16012 33988
rect 16068 33932 16080 33988
rect 16000 33920 16080 33932
rect 16160 34308 16240 34320
rect 16160 34252 16172 34308
rect 16228 34252 16240 34308
rect 16160 33988 16240 34252
rect 16160 33932 16172 33988
rect 16228 33932 16240 33988
rect 16160 33920 16240 33932
rect 16320 34308 16400 34320
rect 16320 34252 16332 34308
rect 16388 34252 16400 34308
rect 16320 33988 16400 34252
rect 16320 33932 16332 33988
rect 16388 33932 16400 33988
rect 16320 33920 16400 33932
rect 16480 34308 16560 34320
rect 16480 34252 16492 34308
rect 16548 34252 16560 34308
rect 16480 33988 16560 34252
rect 16480 33932 16492 33988
rect 16548 33932 16560 33988
rect 16480 33920 16560 33932
rect 16640 34308 16720 34320
rect 16640 34252 16652 34308
rect 16708 34252 16720 34308
rect 16640 33988 16720 34252
rect 16640 33932 16652 33988
rect 16708 33932 16720 33988
rect 16640 33920 16720 33932
rect 16800 34308 16880 34320
rect 16800 34252 16812 34308
rect 16868 34252 16880 34308
rect 16800 33988 16880 34252
rect 16800 33932 16812 33988
rect 16868 33932 16880 33988
rect 16800 33920 16880 33932
rect 16960 34308 17040 34320
rect 16960 34252 16972 34308
rect 17028 34252 17040 34308
rect 16960 33988 17040 34252
rect 16960 33932 16972 33988
rect 17028 33932 17040 33988
rect 16960 33920 17040 33932
rect 17120 34308 17200 34320
rect 17120 34252 17132 34308
rect 17188 34252 17200 34308
rect 17120 33988 17200 34252
rect 17120 33932 17132 33988
rect 17188 33932 17200 33988
rect 17120 33920 17200 33932
rect 17280 34308 17360 34320
rect 17280 34252 17292 34308
rect 17348 34252 17360 34308
rect 17280 33988 17360 34252
rect 17280 33932 17292 33988
rect 17348 33932 17360 33988
rect 17280 33920 17360 33932
rect 17440 34308 17520 34320
rect 17440 34252 17452 34308
rect 17508 34252 17520 34308
rect 17440 33988 17520 34252
rect 17440 33932 17452 33988
rect 17508 33932 17520 33988
rect 17440 33920 17520 33932
rect 17600 34308 17680 34320
rect 17600 34252 17612 34308
rect 17668 34252 17680 34308
rect 17600 33988 17680 34252
rect 17600 33932 17612 33988
rect 17668 33932 17680 33988
rect 17600 33920 17680 33932
rect 17760 34308 17840 34320
rect 17760 34252 17772 34308
rect 17828 34252 17840 34308
rect 17760 33988 17840 34252
rect 17760 33932 17772 33988
rect 17828 33932 17840 33988
rect 17760 33920 17840 33932
rect 17920 34308 18000 34320
rect 17920 34252 17932 34308
rect 17988 34252 18000 34308
rect 17920 33988 18000 34252
rect 17920 33932 17932 33988
rect 17988 33932 18000 33988
rect 17920 33920 18000 33932
rect 18080 34308 18160 34320
rect 18080 34252 18092 34308
rect 18148 34252 18160 34308
rect 18080 33988 18160 34252
rect 18080 33932 18092 33988
rect 18148 33932 18160 33988
rect 18080 33920 18160 33932
rect 18240 34308 18320 34320
rect 18240 34252 18252 34308
rect 18308 34252 18320 34308
rect 18240 33988 18320 34252
rect 18240 33932 18252 33988
rect 18308 33932 18320 33988
rect 18240 33920 18320 33932
rect 18400 34308 18480 34320
rect 18400 34252 18412 34308
rect 18468 34252 18480 34308
rect 18400 33988 18480 34252
rect 18400 33932 18412 33988
rect 18468 33932 18480 33988
rect 18400 33920 18480 33932
rect 18560 34308 18640 34320
rect 18560 34252 18572 34308
rect 18628 34252 18640 34308
rect 18560 33988 18640 34252
rect 18560 33932 18572 33988
rect 18628 33932 18640 33988
rect 18560 33920 18640 33932
rect 18720 34308 18800 34320
rect 18720 34252 18732 34308
rect 18788 34252 18800 34308
rect 18720 33988 18800 34252
rect 18720 33932 18732 33988
rect 18788 33932 18800 33988
rect 18720 33920 18800 33932
rect 18880 34308 18960 34320
rect 18880 34252 18892 34308
rect 18948 34252 18960 34308
rect 18880 33988 18960 34252
rect 18880 33932 18892 33988
rect 18948 33932 18960 33988
rect 18880 33920 18960 33932
rect 12320 33772 12332 33828
rect 12388 33772 12400 33828
rect 12320 33508 12400 33772
rect 12320 33452 12332 33508
rect 12388 33452 12400 33508
rect 12320 33440 12400 33452
rect 12480 33828 12560 33840
rect 12480 33772 12492 33828
rect 12548 33772 12560 33828
rect 12480 33508 12560 33772
rect 12480 33452 12492 33508
rect 12548 33452 12560 33508
rect 12480 33440 12560 33452
rect 12640 33828 12720 33840
rect 12640 33772 12652 33828
rect 12708 33772 12720 33828
rect 12640 33508 12720 33772
rect 12640 33452 12652 33508
rect 12708 33452 12720 33508
rect 12640 33440 12720 33452
rect 12800 33828 12880 33840
rect 12800 33772 12812 33828
rect 12868 33772 12880 33828
rect 12800 33508 12880 33772
rect 12800 33452 12812 33508
rect 12868 33452 12880 33508
rect 12800 33440 12880 33452
rect 12960 33828 13040 33840
rect 12960 33772 12972 33828
rect 13028 33772 13040 33828
rect 12960 33508 13040 33772
rect 12960 33452 12972 33508
rect 13028 33452 13040 33508
rect 12960 33440 13040 33452
rect 13120 33828 13200 33840
rect 13120 33772 13132 33828
rect 13188 33772 13200 33828
rect 13120 33508 13200 33772
rect 13120 33452 13132 33508
rect 13188 33452 13200 33508
rect 13120 33440 13200 33452
rect 13280 33828 13360 33840
rect 13280 33772 13292 33828
rect 13348 33772 13360 33828
rect 13280 33508 13360 33772
rect 13280 33452 13292 33508
rect 13348 33452 13360 33508
rect 13280 33440 13360 33452
rect 13440 33828 13520 33840
rect 13440 33772 13452 33828
rect 13508 33772 13520 33828
rect 13440 33508 13520 33772
rect 13440 33452 13452 33508
rect 13508 33452 13520 33508
rect 13440 33440 13520 33452
rect 13600 33828 13680 33840
rect 13600 33772 13612 33828
rect 13668 33772 13680 33828
rect 13600 33508 13680 33772
rect 13600 33452 13612 33508
rect 13668 33452 13680 33508
rect 13600 33440 13680 33452
rect 13760 33828 13840 33840
rect 13760 33772 13772 33828
rect 13828 33772 13840 33828
rect 13760 33508 13840 33772
rect 13760 33452 13772 33508
rect 13828 33452 13840 33508
rect 13760 33440 13840 33452
rect 13920 33828 14000 33840
rect 13920 33772 13932 33828
rect 13988 33772 14000 33828
rect 13920 33508 14000 33772
rect 13920 33452 13932 33508
rect 13988 33452 14000 33508
rect 13920 33440 14000 33452
rect 14080 33828 14160 33840
rect 14080 33772 14092 33828
rect 14148 33772 14160 33828
rect 14080 33508 14160 33772
rect 14080 33452 14092 33508
rect 14148 33452 14160 33508
rect 14080 33440 14160 33452
rect 14240 33828 14320 33840
rect 14240 33772 14252 33828
rect 14308 33772 14320 33828
rect 14240 33508 14320 33772
rect 14240 33452 14252 33508
rect 14308 33452 14320 33508
rect 14240 33440 14320 33452
rect 14400 33828 14480 33840
rect 14400 33772 14412 33828
rect 14468 33772 14480 33828
rect 14400 33508 14480 33772
rect 14400 33452 14412 33508
rect 14468 33452 14480 33508
rect 14400 33440 14480 33452
rect 14560 33828 14640 33840
rect 14560 33772 14572 33828
rect 14628 33772 14640 33828
rect 14560 33508 14640 33772
rect 14560 33452 14572 33508
rect 14628 33452 14640 33508
rect 14560 33440 14640 33452
rect 14720 33828 14800 33840
rect 14720 33772 14732 33828
rect 14788 33772 14800 33828
rect 14720 33508 14800 33772
rect 14720 33452 14732 33508
rect 14788 33452 14800 33508
rect 14720 33440 14800 33452
rect 14880 33828 14960 33840
rect 14880 33772 14892 33828
rect 14948 33772 14960 33828
rect 14880 33508 14960 33772
rect 14880 33452 14892 33508
rect 14948 33452 14960 33508
rect 14880 33440 14960 33452
rect 15040 33828 15120 33840
rect 15040 33772 15052 33828
rect 15108 33772 15120 33828
rect 15040 33508 15120 33772
rect 15040 33452 15052 33508
rect 15108 33452 15120 33508
rect 15040 33440 15120 33452
rect 15200 33828 15280 33840
rect 15200 33772 15212 33828
rect 15268 33772 15280 33828
rect 15200 33508 15280 33772
rect 15200 33452 15212 33508
rect 15268 33452 15280 33508
rect 15200 33440 15280 33452
rect 15360 33828 15440 33840
rect 15360 33772 15372 33828
rect 15428 33772 15440 33828
rect 15360 33508 15440 33772
rect 15360 33452 15372 33508
rect 15428 33452 15440 33508
rect 15360 33440 15440 33452
rect 15520 33828 15600 33840
rect 15520 33772 15532 33828
rect 15588 33772 15600 33828
rect 15520 33508 15600 33772
rect 15520 33452 15532 33508
rect 15588 33452 15600 33508
rect 15520 33440 15600 33452
rect 15680 33828 15760 33840
rect 15680 33772 15692 33828
rect 15748 33772 15760 33828
rect 15680 33508 15760 33772
rect 15680 33452 15692 33508
rect 15748 33452 15760 33508
rect 15680 33440 15760 33452
rect 15840 33828 15920 33840
rect 15840 33772 15852 33828
rect 15908 33772 15920 33828
rect 15840 33508 15920 33772
rect 15840 33452 15852 33508
rect 15908 33452 15920 33508
rect 15840 33440 15920 33452
rect 16000 33828 16080 33840
rect 16000 33772 16012 33828
rect 16068 33772 16080 33828
rect 16000 33508 16080 33772
rect 16000 33452 16012 33508
rect 16068 33452 16080 33508
rect 16000 33440 16080 33452
rect 16160 33828 16240 33840
rect 16160 33772 16172 33828
rect 16228 33772 16240 33828
rect 16160 33508 16240 33772
rect 16160 33452 16172 33508
rect 16228 33452 16240 33508
rect 16160 33440 16240 33452
rect 16320 33828 16400 33840
rect 16320 33772 16332 33828
rect 16388 33772 16400 33828
rect 16320 33508 16400 33772
rect 16320 33452 16332 33508
rect 16388 33452 16400 33508
rect 16320 33440 16400 33452
rect 16480 33828 16560 33840
rect 16480 33772 16492 33828
rect 16548 33772 16560 33828
rect 16480 33508 16560 33772
rect 16480 33452 16492 33508
rect 16548 33452 16560 33508
rect 16480 33440 16560 33452
rect 16640 33828 16720 33840
rect 16640 33772 16652 33828
rect 16708 33772 16720 33828
rect 16640 33508 16720 33772
rect 16640 33452 16652 33508
rect 16708 33452 16720 33508
rect 16640 33440 16720 33452
rect 16800 33828 16880 33840
rect 16800 33772 16812 33828
rect 16868 33772 16880 33828
rect 16800 33508 16880 33772
rect 16800 33452 16812 33508
rect 16868 33452 16880 33508
rect 16800 33440 16880 33452
rect 16960 33828 17040 33840
rect 16960 33772 16972 33828
rect 17028 33772 17040 33828
rect 16960 33508 17040 33772
rect 16960 33452 16972 33508
rect 17028 33452 17040 33508
rect 16960 33440 17040 33452
rect 17120 33828 17200 33840
rect 17120 33772 17132 33828
rect 17188 33772 17200 33828
rect 17120 33508 17200 33772
rect 17120 33452 17132 33508
rect 17188 33452 17200 33508
rect 17120 33440 17200 33452
rect 17280 33828 17360 33840
rect 17280 33772 17292 33828
rect 17348 33772 17360 33828
rect 17280 33508 17360 33772
rect 17280 33452 17292 33508
rect 17348 33452 17360 33508
rect 17280 33440 17360 33452
rect 17440 33828 17520 33840
rect 17440 33772 17452 33828
rect 17508 33772 17520 33828
rect 17440 33508 17520 33772
rect 17440 33452 17452 33508
rect 17508 33452 17520 33508
rect 17440 33440 17520 33452
rect 17600 33828 17680 33840
rect 17600 33772 17612 33828
rect 17668 33772 17680 33828
rect 17600 33508 17680 33772
rect 17600 33452 17612 33508
rect 17668 33452 17680 33508
rect 17600 33440 17680 33452
rect 17760 33828 17840 33840
rect 17760 33772 17772 33828
rect 17828 33772 17840 33828
rect 17760 33508 17840 33772
rect 17760 33452 17772 33508
rect 17828 33452 17840 33508
rect 17760 33440 17840 33452
rect 17920 33828 18000 33840
rect 17920 33772 17932 33828
rect 17988 33772 18000 33828
rect 17920 33508 18000 33772
rect 17920 33452 17932 33508
rect 17988 33452 18000 33508
rect 17920 33440 18000 33452
rect 18080 33828 18160 33840
rect 18080 33772 18092 33828
rect 18148 33772 18160 33828
rect 18080 33508 18160 33772
rect 18080 33452 18092 33508
rect 18148 33452 18160 33508
rect 18080 33440 18160 33452
rect 18240 33828 18320 33840
rect 18240 33772 18252 33828
rect 18308 33772 18320 33828
rect 18240 33508 18320 33772
rect 18240 33452 18252 33508
rect 18308 33452 18320 33508
rect 18240 33440 18320 33452
rect 18400 33828 18480 33840
rect 18400 33772 18412 33828
rect 18468 33772 18480 33828
rect 18400 33508 18480 33772
rect 18400 33452 18412 33508
rect 18468 33452 18480 33508
rect 18400 33440 18480 33452
rect 18560 33828 18640 33840
rect 18560 33772 18572 33828
rect 18628 33772 18640 33828
rect 18560 33508 18640 33772
rect 18560 33452 18572 33508
rect 18628 33452 18640 33508
rect 18560 33440 18640 33452
rect 18720 33828 18800 33840
rect 18720 33772 18732 33828
rect 18788 33772 18800 33828
rect 18720 33508 18800 33772
rect 18720 33452 18732 33508
rect 18788 33452 18800 33508
rect 18720 33440 18800 33452
rect 18880 33828 18960 33840
rect 18880 33772 18892 33828
rect 18948 33772 18960 33828
rect 18880 33508 18960 33772
rect 18880 33452 18892 33508
rect 18948 33452 18960 33508
rect 18880 33440 18960 33452
rect 19040 33828 19120 37360
rect 19040 33772 19052 33828
rect 19108 33772 19120 33828
rect 19040 33508 19120 33772
rect 19040 33452 19052 33508
rect 19108 33452 19120 33508
rect 0 33348 80 33360
rect 0 33292 12 33348
rect 68 33292 80 33348
rect 0 33028 80 33292
rect 0 32972 12 33028
rect 68 32972 80 33028
rect 0 32960 80 32972
rect 160 33348 240 33360
rect 160 33292 172 33348
rect 228 33292 240 33348
rect 160 33028 240 33292
rect 160 32972 172 33028
rect 228 32972 240 33028
rect 160 32960 240 32972
rect 320 33348 400 33360
rect 320 33292 332 33348
rect 388 33292 400 33348
rect 320 33028 400 33292
rect 320 32972 332 33028
rect 388 32972 400 33028
rect 320 32960 400 32972
rect 480 33348 560 33360
rect 480 33292 492 33348
rect 548 33292 560 33348
rect 480 33028 560 33292
rect 480 32972 492 33028
rect 548 32972 560 33028
rect 480 32960 560 32972
rect 640 33348 720 33360
rect 640 33292 652 33348
rect 708 33292 720 33348
rect 640 33028 720 33292
rect 640 32972 652 33028
rect 708 32972 720 33028
rect 640 32960 720 32972
rect 800 33348 880 33360
rect 800 33292 812 33348
rect 868 33292 880 33348
rect 800 33028 880 33292
rect 800 32972 812 33028
rect 868 32972 880 33028
rect 800 32960 880 32972
rect 960 33348 1040 33360
rect 960 33292 972 33348
rect 1028 33292 1040 33348
rect 960 33028 1040 33292
rect 960 32972 972 33028
rect 1028 32972 1040 33028
rect 960 32960 1040 32972
rect 1120 33348 1200 33360
rect 1120 33292 1132 33348
rect 1188 33292 1200 33348
rect 1120 33028 1200 33292
rect 1120 32972 1132 33028
rect 1188 32972 1200 33028
rect 1120 32960 1200 32972
rect 1280 33348 1360 33360
rect 1280 33292 1292 33348
rect 1348 33292 1360 33348
rect 1280 33028 1360 33292
rect 1280 32972 1292 33028
rect 1348 32972 1360 33028
rect 1280 32960 1360 32972
rect 1440 33348 1520 33360
rect 1440 33292 1452 33348
rect 1508 33292 1520 33348
rect 1440 33028 1520 33292
rect 1440 32972 1452 33028
rect 1508 32972 1520 33028
rect 1440 32960 1520 32972
rect 1600 33348 1680 33360
rect 1600 33292 1612 33348
rect 1668 33292 1680 33348
rect 1600 33028 1680 33292
rect 1600 32972 1612 33028
rect 1668 32972 1680 33028
rect 1600 32960 1680 32972
rect 1760 33348 1840 33360
rect 1760 33292 1772 33348
rect 1828 33292 1840 33348
rect 1760 33028 1840 33292
rect 1760 32972 1772 33028
rect 1828 32972 1840 33028
rect 1760 32960 1840 32972
rect 1920 33348 2000 33360
rect 1920 33292 1932 33348
rect 1988 33292 2000 33348
rect 1920 33028 2000 33292
rect 1920 32972 1932 33028
rect 1988 32972 2000 33028
rect 1920 32960 2000 32972
rect 2080 33348 2160 33360
rect 2080 33292 2092 33348
rect 2148 33292 2160 33348
rect 2080 33028 2160 33292
rect 2080 32972 2092 33028
rect 2148 32972 2160 33028
rect 2080 32960 2160 32972
rect 2240 33348 2320 33360
rect 2240 33292 2252 33348
rect 2308 33292 2320 33348
rect 2240 33028 2320 33292
rect 2240 32972 2252 33028
rect 2308 32972 2320 33028
rect 2240 32960 2320 32972
rect 2400 33348 2480 33360
rect 2400 33292 2412 33348
rect 2468 33292 2480 33348
rect 2400 33028 2480 33292
rect 2400 32972 2412 33028
rect 2468 32972 2480 33028
rect 2400 32960 2480 32972
rect 2560 33348 2640 33360
rect 2560 33292 2572 33348
rect 2628 33292 2640 33348
rect 2560 33028 2640 33292
rect 2560 32972 2572 33028
rect 2628 32972 2640 33028
rect 2560 32960 2640 32972
rect 2720 33348 2800 33360
rect 2720 33292 2732 33348
rect 2788 33292 2800 33348
rect 2720 33028 2800 33292
rect 2720 32972 2732 33028
rect 2788 32972 2800 33028
rect 2720 32960 2800 32972
rect 2880 33348 2960 33360
rect 2880 33292 2892 33348
rect 2948 33292 2960 33348
rect 2880 33028 2960 33292
rect 2880 32972 2892 33028
rect 2948 32972 2960 33028
rect 2880 32960 2960 32972
rect 3040 33348 3120 33360
rect 3040 33292 3052 33348
rect 3108 33292 3120 33348
rect 3040 33028 3120 33292
rect 3040 32972 3052 33028
rect 3108 32972 3120 33028
rect 3040 32960 3120 32972
rect 3200 33348 3280 33360
rect 3200 33292 3212 33348
rect 3268 33292 3280 33348
rect 3200 33028 3280 33292
rect 3200 32972 3212 33028
rect 3268 32972 3280 33028
rect 3200 32960 3280 32972
rect 3360 33348 3440 33360
rect 3360 33292 3372 33348
rect 3428 33292 3440 33348
rect 3360 33028 3440 33292
rect 3360 32972 3372 33028
rect 3428 32972 3440 33028
rect 3360 32960 3440 32972
rect 3520 33348 3600 33360
rect 3520 33292 3532 33348
rect 3588 33292 3600 33348
rect 3520 33028 3600 33292
rect 3520 32972 3532 33028
rect 3588 32972 3600 33028
rect 3520 32960 3600 32972
rect 3680 33348 3760 33360
rect 3680 33292 3692 33348
rect 3748 33292 3760 33348
rect 3680 33028 3760 33292
rect 3680 32972 3692 33028
rect 3748 32972 3760 33028
rect 3680 32960 3760 32972
rect 3840 33348 3920 33360
rect 3840 33292 3852 33348
rect 3908 33292 3920 33348
rect 3840 33028 3920 33292
rect 3840 32972 3852 33028
rect 3908 32972 3920 33028
rect 3840 32960 3920 32972
rect 4000 33348 4080 33360
rect 4000 33292 4012 33348
rect 4068 33292 4080 33348
rect 4000 33028 4080 33292
rect 4000 32972 4012 33028
rect 4068 32972 4080 33028
rect 4000 32960 4080 32972
rect 4160 33348 4240 33360
rect 4160 33292 4172 33348
rect 4228 33292 4240 33348
rect 4160 33028 4240 33292
rect 4160 32972 4172 33028
rect 4228 32972 4240 33028
rect 4160 32960 4240 32972
rect 4320 33348 4400 33360
rect 4320 33292 4332 33348
rect 4388 33292 4400 33348
rect 4320 33028 4400 33292
rect 4320 32972 4332 33028
rect 4388 32972 4400 33028
rect 4320 32960 4400 32972
rect 4480 33348 4560 33360
rect 4480 33292 4492 33348
rect 4548 33292 4560 33348
rect 4480 33028 4560 33292
rect 4480 32972 4492 33028
rect 4548 32972 4560 33028
rect 4480 32960 4560 32972
rect 4640 33348 4720 33360
rect 4640 33292 4652 33348
rect 4708 33292 4720 33348
rect 4640 33028 4720 33292
rect 4640 32972 4652 33028
rect 4708 32972 4720 33028
rect 4640 32960 4720 32972
rect 4800 33348 4880 33360
rect 4800 33292 4812 33348
rect 4868 33292 4880 33348
rect 4800 33028 4880 33292
rect 4800 32972 4812 33028
rect 4868 32972 4880 33028
rect 4800 32960 4880 32972
rect 4960 33348 5040 33360
rect 4960 33292 4972 33348
rect 5028 33292 5040 33348
rect 4960 33028 5040 33292
rect 4960 32972 4972 33028
rect 5028 32972 5040 33028
rect 4960 32960 5040 32972
rect 5120 33348 5200 33360
rect 5120 33292 5132 33348
rect 5188 33292 5200 33348
rect 5120 33028 5200 33292
rect 5120 32972 5132 33028
rect 5188 32972 5200 33028
rect 5120 32960 5200 32972
rect 5280 33348 5360 33360
rect 5280 33292 5292 33348
rect 5348 33292 5360 33348
rect 5280 33028 5360 33292
rect 5280 32972 5292 33028
rect 5348 32972 5360 33028
rect 5280 32960 5360 32972
rect 5440 33348 5520 33360
rect 5440 33292 5452 33348
rect 5508 33292 5520 33348
rect 5440 33028 5520 33292
rect 5440 32972 5452 33028
rect 5508 32972 5520 33028
rect 5440 32960 5520 32972
rect 5600 33348 5680 33360
rect 5600 33292 5612 33348
rect 5668 33292 5680 33348
rect 5600 33028 5680 33292
rect 5600 32972 5612 33028
rect 5668 32972 5680 33028
rect 5600 32960 5680 32972
rect 5760 33348 5840 33360
rect 5760 33292 5772 33348
rect 5828 33292 5840 33348
rect 5760 33028 5840 33292
rect 5760 32972 5772 33028
rect 5828 32972 5840 33028
rect 5760 32960 5840 32972
rect 5920 33348 6000 33360
rect 5920 33292 5932 33348
rect 5988 33292 6000 33348
rect 5920 33028 6000 33292
rect 5920 32972 5932 33028
rect 5988 32972 6000 33028
rect 5920 32960 6000 32972
rect 6080 33348 6160 33360
rect 6080 33292 6092 33348
rect 6148 33292 6160 33348
rect 6080 33028 6160 33292
rect 6080 32972 6092 33028
rect 6148 32972 6160 33028
rect 6080 32960 6160 32972
rect 6240 33348 6320 33360
rect 6240 33292 6252 33348
rect 6308 33292 6320 33348
rect 6240 33028 6320 33292
rect 6240 32972 6252 33028
rect 6308 32972 6320 33028
rect 6240 32960 6320 32972
rect 6400 33348 6480 33360
rect 6400 33292 6412 33348
rect 6468 33292 6480 33348
rect 6400 33028 6480 33292
rect 6400 32972 6412 33028
rect 6468 32972 6480 33028
rect 6400 32960 6480 32972
rect 6560 33348 6640 33360
rect 6560 33292 6572 33348
rect 6628 33292 6640 33348
rect 6560 33028 6640 33292
rect 6560 32972 6572 33028
rect 6628 32972 6640 33028
rect 6560 32960 6640 32972
rect 6720 33348 6800 33360
rect 6720 33292 6732 33348
rect 6788 33292 6800 33348
rect 6720 33028 6800 33292
rect 6720 32972 6732 33028
rect 6788 32972 6800 33028
rect 6720 32960 6800 32972
rect 6880 33348 6960 33360
rect 6880 33292 6892 33348
rect 6948 33292 6960 33348
rect 6880 33028 6960 33292
rect 6880 32972 6892 33028
rect 6948 32972 6960 33028
rect 6880 32960 6960 32972
rect 7040 33348 7120 33360
rect 7040 33292 7052 33348
rect 7108 33292 7120 33348
rect 7040 33028 7120 33292
rect 7040 32972 7052 33028
rect 7108 32972 7120 33028
rect 7040 32960 7120 32972
rect 7200 33348 7280 33360
rect 7200 33292 7212 33348
rect 7268 33292 7280 33348
rect 7200 33028 7280 33292
rect 7200 32972 7212 33028
rect 7268 32972 7280 33028
rect 7200 32960 7280 32972
rect 7360 33348 7440 33360
rect 7360 33292 7372 33348
rect 7428 33292 7440 33348
rect 7360 33028 7440 33292
rect 7360 32972 7372 33028
rect 7428 32972 7440 33028
rect 7360 32960 7440 32972
rect 7520 33348 7600 33360
rect 7520 33292 7532 33348
rect 7588 33292 7600 33348
rect 7520 33028 7600 33292
rect 7520 32972 7532 33028
rect 7588 32972 7600 33028
rect 7520 32960 7600 32972
rect 7680 33348 7760 33360
rect 7680 33292 7692 33348
rect 7748 33292 7760 33348
rect 7680 33028 7760 33292
rect 7680 32972 7692 33028
rect 7748 32972 7760 33028
rect 7680 32960 7760 32972
rect 7840 33348 7920 33360
rect 7840 33292 7852 33348
rect 7908 33292 7920 33348
rect 7840 33028 7920 33292
rect 7840 32972 7852 33028
rect 7908 32972 7920 33028
rect 7840 32960 7920 32972
rect 8000 33348 8080 33360
rect 8000 33292 8012 33348
rect 8068 33292 8080 33348
rect 8000 33028 8080 33292
rect 8000 32972 8012 33028
rect 8068 32972 8080 33028
rect 8000 32960 8080 32972
rect 8160 33348 8240 33360
rect 8160 33292 8172 33348
rect 8228 33292 8240 33348
rect 8160 33028 8240 33292
rect 8160 32972 8172 33028
rect 8228 32972 8240 33028
rect 8160 32960 8240 32972
rect 8320 33348 8400 33360
rect 8320 33292 8332 33348
rect 8388 33292 8400 33348
rect 8320 33028 8400 33292
rect 8320 32972 8332 33028
rect 8388 32972 8400 33028
rect 8320 32960 8400 32972
rect 8480 33348 8560 33360
rect 8480 33292 8492 33348
rect 8548 33292 8560 33348
rect 8480 33028 8560 33292
rect 8480 32972 8492 33028
rect 8548 32972 8560 33028
rect 0 32868 80 32880
rect 0 32812 12 32868
rect 68 32812 80 32868
rect 0 32548 80 32812
rect 0 32492 12 32548
rect 68 32492 80 32548
rect 0 32480 80 32492
rect 160 32868 240 32880
rect 160 32812 172 32868
rect 228 32812 240 32868
rect 160 32548 240 32812
rect 160 32492 172 32548
rect 228 32492 240 32548
rect 160 32480 240 32492
rect 320 32868 400 32880
rect 320 32812 332 32868
rect 388 32812 400 32868
rect 320 32548 400 32812
rect 320 32492 332 32548
rect 388 32492 400 32548
rect 320 32480 400 32492
rect 480 32868 560 32880
rect 480 32812 492 32868
rect 548 32812 560 32868
rect 480 32548 560 32812
rect 480 32492 492 32548
rect 548 32492 560 32548
rect 480 32480 560 32492
rect 640 32868 720 32880
rect 640 32812 652 32868
rect 708 32812 720 32868
rect 640 32548 720 32812
rect 640 32492 652 32548
rect 708 32492 720 32548
rect 640 32480 720 32492
rect 800 32868 880 32880
rect 800 32812 812 32868
rect 868 32812 880 32868
rect 800 32548 880 32812
rect 800 32492 812 32548
rect 868 32492 880 32548
rect 800 32480 880 32492
rect 960 32868 1040 32880
rect 960 32812 972 32868
rect 1028 32812 1040 32868
rect 960 32548 1040 32812
rect 960 32492 972 32548
rect 1028 32492 1040 32548
rect 960 32480 1040 32492
rect 1120 32868 1200 32880
rect 1120 32812 1132 32868
rect 1188 32812 1200 32868
rect 1120 32548 1200 32812
rect 1120 32492 1132 32548
rect 1188 32492 1200 32548
rect 1120 32480 1200 32492
rect 1280 32868 1360 32880
rect 1280 32812 1292 32868
rect 1348 32812 1360 32868
rect 1280 32548 1360 32812
rect 1280 32492 1292 32548
rect 1348 32492 1360 32548
rect 1280 32480 1360 32492
rect 1440 32868 1520 32880
rect 1440 32812 1452 32868
rect 1508 32812 1520 32868
rect 1440 32548 1520 32812
rect 1440 32492 1452 32548
rect 1508 32492 1520 32548
rect 1440 32480 1520 32492
rect 1600 32868 1680 32880
rect 1600 32812 1612 32868
rect 1668 32812 1680 32868
rect 1600 32548 1680 32812
rect 1600 32492 1612 32548
rect 1668 32492 1680 32548
rect 1600 32480 1680 32492
rect 1760 32868 1840 32880
rect 1760 32812 1772 32868
rect 1828 32812 1840 32868
rect 1760 32548 1840 32812
rect 1760 32492 1772 32548
rect 1828 32492 1840 32548
rect 1760 32480 1840 32492
rect 1920 32868 2000 32880
rect 1920 32812 1932 32868
rect 1988 32812 2000 32868
rect 1920 32548 2000 32812
rect 1920 32492 1932 32548
rect 1988 32492 2000 32548
rect 1920 32480 2000 32492
rect 2080 32868 2160 32880
rect 2080 32812 2092 32868
rect 2148 32812 2160 32868
rect 2080 32548 2160 32812
rect 2080 32492 2092 32548
rect 2148 32492 2160 32548
rect 2080 32480 2160 32492
rect 2240 32868 2320 32880
rect 2240 32812 2252 32868
rect 2308 32812 2320 32868
rect 2240 32548 2320 32812
rect 2240 32492 2252 32548
rect 2308 32492 2320 32548
rect 2240 32480 2320 32492
rect 2400 32868 2480 32880
rect 2400 32812 2412 32868
rect 2468 32812 2480 32868
rect 2400 32548 2480 32812
rect 2400 32492 2412 32548
rect 2468 32492 2480 32548
rect 2400 32480 2480 32492
rect 2560 32868 2640 32880
rect 2560 32812 2572 32868
rect 2628 32812 2640 32868
rect 2560 32548 2640 32812
rect 2560 32492 2572 32548
rect 2628 32492 2640 32548
rect 2560 32480 2640 32492
rect 2720 32868 2800 32880
rect 2720 32812 2732 32868
rect 2788 32812 2800 32868
rect 2720 32548 2800 32812
rect 2720 32492 2732 32548
rect 2788 32492 2800 32548
rect 2720 32480 2800 32492
rect 2880 32868 2960 32880
rect 2880 32812 2892 32868
rect 2948 32812 2960 32868
rect 2880 32548 2960 32812
rect 2880 32492 2892 32548
rect 2948 32492 2960 32548
rect 2880 32480 2960 32492
rect 3040 32868 3120 32880
rect 3040 32812 3052 32868
rect 3108 32812 3120 32868
rect 3040 32548 3120 32812
rect 3040 32492 3052 32548
rect 3108 32492 3120 32548
rect 3040 32480 3120 32492
rect 3200 32868 3280 32880
rect 3200 32812 3212 32868
rect 3268 32812 3280 32868
rect 3200 32548 3280 32812
rect 3200 32492 3212 32548
rect 3268 32492 3280 32548
rect 3200 32480 3280 32492
rect 3360 32868 3440 32880
rect 3360 32812 3372 32868
rect 3428 32812 3440 32868
rect 3360 32548 3440 32812
rect 3360 32492 3372 32548
rect 3428 32492 3440 32548
rect 3360 32480 3440 32492
rect 3520 32868 3600 32880
rect 3520 32812 3532 32868
rect 3588 32812 3600 32868
rect 3520 32548 3600 32812
rect 3520 32492 3532 32548
rect 3588 32492 3600 32548
rect 3520 32480 3600 32492
rect 3680 32868 3760 32880
rect 3680 32812 3692 32868
rect 3748 32812 3760 32868
rect 3680 32548 3760 32812
rect 3680 32492 3692 32548
rect 3748 32492 3760 32548
rect 3680 32480 3760 32492
rect 3840 32868 3920 32880
rect 3840 32812 3852 32868
rect 3908 32812 3920 32868
rect 3840 32548 3920 32812
rect 3840 32492 3852 32548
rect 3908 32492 3920 32548
rect 3840 32480 3920 32492
rect 4000 32868 4080 32880
rect 4000 32812 4012 32868
rect 4068 32812 4080 32868
rect 4000 32548 4080 32812
rect 4000 32492 4012 32548
rect 4068 32492 4080 32548
rect 4000 32480 4080 32492
rect 4160 32868 4240 32880
rect 4160 32812 4172 32868
rect 4228 32812 4240 32868
rect 4160 32548 4240 32812
rect 4160 32492 4172 32548
rect 4228 32492 4240 32548
rect 4160 32480 4240 32492
rect 4320 32868 4400 32880
rect 4320 32812 4332 32868
rect 4388 32812 4400 32868
rect 4320 32548 4400 32812
rect 4320 32492 4332 32548
rect 4388 32492 4400 32548
rect 4320 32480 4400 32492
rect 4480 32868 4560 32880
rect 4480 32812 4492 32868
rect 4548 32812 4560 32868
rect 4480 32548 4560 32812
rect 4480 32492 4492 32548
rect 4548 32492 4560 32548
rect 4480 32480 4560 32492
rect 4640 32868 4720 32880
rect 4640 32812 4652 32868
rect 4708 32812 4720 32868
rect 4640 32548 4720 32812
rect 4640 32492 4652 32548
rect 4708 32492 4720 32548
rect 4640 32480 4720 32492
rect 4800 32868 4880 32880
rect 4800 32812 4812 32868
rect 4868 32812 4880 32868
rect 4800 32548 4880 32812
rect 4800 32492 4812 32548
rect 4868 32492 4880 32548
rect 4800 32480 4880 32492
rect 4960 32868 5040 32880
rect 4960 32812 4972 32868
rect 5028 32812 5040 32868
rect 4960 32548 5040 32812
rect 4960 32492 4972 32548
rect 5028 32492 5040 32548
rect 4960 32480 5040 32492
rect 5120 32868 5200 32880
rect 5120 32812 5132 32868
rect 5188 32812 5200 32868
rect 5120 32548 5200 32812
rect 5120 32492 5132 32548
rect 5188 32492 5200 32548
rect 5120 32480 5200 32492
rect 5280 32868 5360 32880
rect 5280 32812 5292 32868
rect 5348 32812 5360 32868
rect 5280 32548 5360 32812
rect 5280 32492 5292 32548
rect 5348 32492 5360 32548
rect 5280 32480 5360 32492
rect 5440 32868 5520 32880
rect 5440 32812 5452 32868
rect 5508 32812 5520 32868
rect 5440 32548 5520 32812
rect 5440 32492 5452 32548
rect 5508 32492 5520 32548
rect 5440 32480 5520 32492
rect 5600 32868 5680 32880
rect 5600 32812 5612 32868
rect 5668 32812 5680 32868
rect 5600 32548 5680 32812
rect 5600 32492 5612 32548
rect 5668 32492 5680 32548
rect 5600 32480 5680 32492
rect 5760 32868 5840 32880
rect 5760 32812 5772 32868
rect 5828 32812 5840 32868
rect 5760 32548 5840 32812
rect 5760 32492 5772 32548
rect 5828 32492 5840 32548
rect 5760 32480 5840 32492
rect 5920 32868 6000 32880
rect 5920 32812 5932 32868
rect 5988 32812 6000 32868
rect 5920 32548 6000 32812
rect 5920 32492 5932 32548
rect 5988 32492 6000 32548
rect 5920 32480 6000 32492
rect 6080 32868 6160 32880
rect 6080 32812 6092 32868
rect 6148 32812 6160 32868
rect 6080 32548 6160 32812
rect 6080 32492 6092 32548
rect 6148 32492 6160 32548
rect 6080 32480 6160 32492
rect 6240 32868 6320 32880
rect 6240 32812 6252 32868
rect 6308 32812 6320 32868
rect 6240 32548 6320 32812
rect 6240 32492 6252 32548
rect 6308 32492 6320 32548
rect 6240 32480 6320 32492
rect 6400 32868 6480 32880
rect 6400 32812 6412 32868
rect 6468 32812 6480 32868
rect 6400 32548 6480 32812
rect 6400 32492 6412 32548
rect 6468 32492 6480 32548
rect 6400 32480 6480 32492
rect 6560 32868 6640 32880
rect 6560 32812 6572 32868
rect 6628 32812 6640 32868
rect 6560 32548 6640 32812
rect 6560 32492 6572 32548
rect 6628 32492 6640 32548
rect 6560 32480 6640 32492
rect 6720 32868 6800 32880
rect 6720 32812 6732 32868
rect 6788 32812 6800 32868
rect 6720 32548 6800 32812
rect 6720 32492 6732 32548
rect 6788 32492 6800 32548
rect 6720 32480 6800 32492
rect 6880 32868 6960 32880
rect 6880 32812 6892 32868
rect 6948 32812 6960 32868
rect 6880 32548 6960 32812
rect 6880 32492 6892 32548
rect 6948 32492 6960 32548
rect 6880 32480 6960 32492
rect 7040 32868 7120 32880
rect 7040 32812 7052 32868
rect 7108 32812 7120 32868
rect 7040 32548 7120 32812
rect 7040 32492 7052 32548
rect 7108 32492 7120 32548
rect 7040 32480 7120 32492
rect 7200 32868 7280 32880
rect 7200 32812 7212 32868
rect 7268 32812 7280 32868
rect 7200 32548 7280 32812
rect 7200 32492 7212 32548
rect 7268 32492 7280 32548
rect 7200 32480 7280 32492
rect 7360 32868 7440 32880
rect 7360 32812 7372 32868
rect 7428 32812 7440 32868
rect 7360 32548 7440 32812
rect 7360 32492 7372 32548
rect 7428 32492 7440 32548
rect 7360 32480 7440 32492
rect 7520 32868 7600 32880
rect 7520 32812 7532 32868
rect 7588 32812 7600 32868
rect 7520 32548 7600 32812
rect 7520 32492 7532 32548
rect 7588 32492 7600 32548
rect 7520 32480 7600 32492
rect 7680 32868 7760 32880
rect 7680 32812 7692 32868
rect 7748 32812 7760 32868
rect 7680 32548 7760 32812
rect 7680 32492 7692 32548
rect 7748 32492 7760 32548
rect 7680 32480 7760 32492
rect 7840 32868 7920 32880
rect 7840 32812 7852 32868
rect 7908 32812 7920 32868
rect 7840 32548 7920 32812
rect 7840 32492 7852 32548
rect 7908 32492 7920 32548
rect 7840 32480 7920 32492
rect 8000 32868 8080 32880
rect 8000 32812 8012 32868
rect 8068 32812 8080 32868
rect 8000 32548 8080 32812
rect 8000 32492 8012 32548
rect 8068 32492 8080 32548
rect 8000 32480 8080 32492
rect 8160 32868 8240 32880
rect 8160 32812 8172 32868
rect 8228 32812 8240 32868
rect 8160 32548 8240 32812
rect 8160 32492 8172 32548
rect 8228 32492 8240 32548
rect 8160 32480 8240 32492
rect 8320 32868 8400 32880
rect 8320 32812 8332 32868
rect 8388 32812 8400 32868
rect 8320 32548 8400 32812
rect 8320 32492 8332 32548
rect 8388 32492 8400 32548
rect 8320 32480 8400 32492
rect 0 32388 80 32400
rect 0 32332 12 32388
rect 68 32332 80 32388
rect 0 32068 80 32332
rect 0 32012 12 32068
rect 68 32012 80 32068
rect 0 31748 80 32012
rect 0 31692 12 31748
rect 68 31692 80 31748
rect 0 31428 80 31692
rect 0 31372 12 31428
rect 68 31372 80 31428
rect 0 31108 80 31372
rect 0 31052 12 31108
rect 68 31052 80 31108
rect 0 30788 80 31052
rect 0 30732 12 30788
rect 68 30732 80 30788
rect 0 30468 80 30732
rect 0 30412 12 30468
rect 68 30412 80 30468
rect 0 30400 80 30412
rect 160 32388 240 32400
rect 160 32332 172 32388
rect 228 32332 240 32388
rect 160 32068 240 32332
rect 160 32012 172 32068
rect 228 32012 240 32068
rect 160 31748 240 32012
rect 160 31692 172 31748
rect 228 31692 240 31748
rect 160 31428 240 31692
rect 160 31372 172 31428
rect 228 31372 240 31428
rect 160 31108 240 31372
rect 160 31052 172 31108
rect 228 31052 240 31108
rect 160 30788 240 31052
rect 160 30732 172 30788
rect 228 30732 240 30788
rect 160 30468 240 30732
rect 160 30412 172 30468
rect 228 30412 240 30468
rect 160 30400 240 30412
rect 320 32388 400 32400
rect 320 32332 332 32388
rect 388 32332 400 32388
rect 320 32068 400 32332
rect 320 32012 332 32068
rect 388 32012 400 32068
rect 320 31748 400 32012
rect 320 31692 332 31748
rect 388 31692 400 31748
rect 320 31428 400 31692
rect 320 31372 332 31428
rect 388 31372 400 31428
rect 320 31108 400 31372
rect 320 31052 332 31108
rect 388 31052 400 31108
rect 320 30788 400 31052
rect 320 30732 332 30788
rect 388 30732 400 30788
rect 320 30468 400 30732
rect 320 30412 332 30468
rect 388 30412 400 30468
rect 320 30400 400 30412
rect 480 32388 560 32400
rect 480 32332 492 32388
rect 548 32332 560 32388
rect 480 32068 560 32332
rect 480 32012 492 32068
rect 548 32012 560 32068
rect 480 31748 560 32012
rect 480 31692 492 31748
rect 548 31692 560 31748
rect 480 31428 560 31692
rect 480 31372 492 31428
rect 548 31372 560 31428
rect 480 31108 560 31372
rect 480 31052 492 31108
rect 548 31052 560 31108
rect 480 30788 560 31052
rect 480 30732 492 30788
rect 548 30732 560 30788
rect 480 30468 560 30732
rect 480 30412 492 30468
rect 548 30412 560 30468
rect 480 30400 560 30412
rect 640 32388 720 32400
rect 640 32332 652 32388
rect 708 32332 720 32388
rect 640 32068 720 32332
rect 640 32012 652 32068
rect 708 32012 720 32068
rect 640 31748 720 32012
rect 640 31692 652 31748
rect 708 31692 720 31748
rect 640 31428 720 31692
rect 640 31372 652 31428
rect 708 31372 720 31428
rect 640 31108 720 31372
rect 640 31052 652 31108
rect 708 31052 720 31108
rect 640 30788 720 31052
rect 640 30732 652 30788
rect 708 30732 720 30788
rect 640 30468 720 30732
rect 640 30412 652 30468
rect 708 30412 720 30468
rect 640 30400 720 30412
rect 800 32388 880 32400
rect 800 32332 812 32388
rect 868 32332 880 32388
rect 800 32068 880 32332
rect 800 32012 812 32068
rect 868 32012 880 32068
rect 800 31748 880 32012
rect 800 31692 812 31748
rect 868 31692 880 31748
rect 800 31428 880 31692
rect 800 31372 812 31428
rect 868 31372 880 31428
rect 800 31108 880 31372
rect 800 31052 812 31108
rect 868 31052 880 31108
rect 800 30788 880 31052
rect 800 30732 812 30788
rect 868 30732 880 30788
rect 800 30468 880 30732
rect 800 30412 812 30468
rect 868 30412 880 30468
rect 800 30400 880 30412
rect 960 32388 1040 32400
rect 960 32332 972 32388
rect 1028 32332 1040 32388
rect 960 32068 1040 32332
rect 960 32012 972 32068
rect 1028 32012 1040 32068
rect 960 31748 1040 32012
rect 960 31692 972 31748
rect 1028 31692 1040 31748
rect 960 31428 1040 31692
rect 960 31372 972 31428
rect 1028 31372 1040 31428
rect 960 31108 1040 31372
rect 960 31052 972 31108
rect 1028 31052 1040 31108
rect 960 30788 1040 31052
rect 960 30732 972 30788
rect 1028 30732 1040 30788
rect 960 30468 1040 30732
rect 960 30412 972 30468
rect 1028 30412 1040 30468
rect 960 30400 1040 30412
rect 1120 32388 1200 32400
rect 1120 32332 1132 32388
rect 1188 32332 1200 32388
rect 1120 32068 1200 32332
rect 1120 32012 1132 32068
rect 1188 32012 1200 32068
rect 1120 31748 1200 32012
rect 1120 31692 1132 31748
rect 1188 31692 1200 31748
rect 1120 31428 1200 31692
rect 1120 31372 1132 31428
rect 1188 31372 1200 31428
rect 1120 31108 1200 31372
rect 1120 31052 1132 31108
rect 1188 31052 1200 31108
rect 1120 30788 1200 31052
rect 1120 30732 1132 30788
rect 1188 30732 1200 30788
rect 1120 30468 1200 30732
rect 1120 30412 1132 30468
rect 1188 30412 1200 30468
rect 1120 30400 1200 30412
rect 1280 32388 1360 32400
rect 1280 32332 1292 32388
rect 1348 32332 1360 32388
rect 1280 32068 1360 32332
rect 1280 32012 1292 32068
rect 1348 32012 1360 32068
rect 1280 31748 1360 32012
rect 1280 31692 1292 31748
rect 1348 31692 1360 31748
rect 1280 31428 1360 31692
rect 1280 31372 1292 31428
rect 1348 31372 1360 31428
rect 1280 31108 1360 31372
rect 1280 31052 1292 31108
rect 1348 31052 1360 31108
rect 1280 30788 1360 31052
rect 1280 30732 1292 30788
rect 1348 30732 1360 30788
rect 1280 30468 1360 30732
rect 1280 30412 1292 30468
rect 1348 30412 1360 30468
rect 1280 30400 1360 30412
rect 1440 32388 1520 32400
rect 1440 32332 1452 32388
rect 1508 32332 1520 32388
rect 1440 32068 1520 32332
rect 1440 32012 1452 32068
rect 1508 32012 1520 32068
rect 1440 31748 1520 32012
rect 1440 31692 1452 31748
rect 1508 31692 1520 31748
rect 1440 31428 1520 31692
rect 1440 31372 1452 31428
rect 1508 31372 1520 31428
rect 1440 31108 1520 31372
rect 1440 31052 1452 31108
rect 1508 31052 1520 31108
rect 1440 30788 1520 31052
rect 1440 30732 1452 30788
rect 1508 30732 1520 30788
rect 1440 30468 1520 30732
rect 1440 30412 1452 30468
rect 1508 30412 1520 30468
rect 1440 30400 1520 30412
rect 1600 32388 1680 32400
rect 1600 32332 1612 32388
rect 1668 32332 1680 32388
rect 1600 32068 1680 32332
rect 1600 32012 1612 32068
rect 1668 32012 1680 32068
rect 1600 31748 1680 32012
rect 1600 31692 1612 31748
rect 1668 31692 1680 31748
rect 1600 31428 1680 31692
rect 1600 31372 1612 31428
rect 1668 31372 1680 31428
rect 1600 31108 1680 31372
rect 1600 31052 1612 31108
rect 1668 31052 1680 31108
rect 1600 30788 1680 31052
rect 1600 30732 1612 30788
rect 1668 30732 1680 30788
rect 1600 30468 1680 30732
rect 1600 30412 1612 30468
rect 1668 30412 1680 30468
rect 1600 30400 1680 30412
rect 1760 32388 1840 32400
rect 1760 32332 1772 32388
rect 1828 32332 1840 32388
rect 1760 32068 1840 32332
rect 1760 32012 1772 32068
rect 1828 32012 1840 32068
rect 1760 31748 1840 32012
rect 1760 31692 1772 31748
rect 1828 31692 1840 31748
rect 1760 31428 1840 31692
rect 1760 31372 1772 31428
rect 1828 31372 1840 31428
rect 1760 31108 1840 31372
rect 1760 31052 1772 31108
rect 1828 31052 1840 31108
rect 1760 30788 1840 31052
rect 1760 30732 1772 30788
rect 1828 30732 1840 30788
rect 1760 30468 1840 30732
rect 1760 30412 1772 30468
rect 1828 30412 1840 30468
rect 1760 30400 1840 30412
rect 1920 32388 2000 32400
rect 1920 32332 1932 32388
rect 1988 32332 2000 32388
rect 1920 32068 2000 32332
rect 1920 32012 1932 32068
rect 1988 32012 2000 32068
rect 1920 31748 2000 32012
rect 1920 31692 1932 31748
rect 1988 31692 2000 31748
rect 1920 31428 2000 31692
rect 1920 31372 1932 31428
rect 1988 31372 2000 31428
rect 1920 31108 2000 31372
rect 1920 31052 1932 31108
rect 1988 31052 2000 31108
rect 1920 30788 2000 31052
rect 1920 30732 1932 30788
rect 1988 30732 2000 30788
rect 1920 30468 2000 30732
rect 1920 30412 1932 30468
rect 1988 30412 2000 30468
rect 1920 30400 2000 30412
rect 2080 32388 2160 32400
rect 2080 32332 2092 32388
rect 2148 32332 2160 32388
rect 2080 32068 2160 32332
rect 2080 32012 2092 32068
rect 2148 32012 2160 32068
rect 2080 31748 2160 32012
rect 2080 31692 2092 31748
rect 2148 31692 2160 31748
rect 2080 31428 2160 31692
rect 2080 31372 2092 31428
rect 2148 31372 2160 31428
rect 2080 31108 2160 31372
rect 2080 31052 2092 31108
rect 2148 31052 2160 31108
rect 2080 30788 2160 31052
rect 2080 30732 2092 30788
rect 2148 30732 2160 30788
rect 2080 30468 2160 30732
rect 2080 30412 2092 30468
rect 2148 30412 2160 30468
rect 2080 30400 2160 30412
rect 2240 32388 2320 32400
rect 2240 32332 2252 32388
rect 2308 32332 2320 32388
rect 2240 32068 2320 32332
rect 2240 32012 2252 32068
rect 2308 32012 2320 32068
rect 2240 31748 2320 32012
rect 2240 31692 2252 31748
rect 2308 31692 2320 31748
rect 2240 31428 2320 31692
rect 2240 31372 2252 31428
rect 2308 31372 2320 31428
rect 2240 31108 2320 31372
rect 2240 31052 2252 31108
rect 2308 31052 2320 31108
rect 2240 30788 2320 31052
rect 2240 30732 2252 30788
rect 2308 30732 2320 30788
rect 2240 30468 2320 30732
rect 2240 30412 2252 30468
rect 2308 30412 2320 30468
rect 2240 30400 2320 30412
rect 2400 32388 2480 32400
rect 2400 32332 2412 32388
rect 2468 32332 2480 32388
rect 2400 32068 2480 32332
rect 2400 32012 2412 32068
rect 2468 32012 2480 32068
rect 2400 31748 2480 32012
rect 2400 31692 2412 31748
rect 2468 31692 2480 31748
rect 2400 31428 2480 31692
rect 2400 31372 2412 31428
rect 2468 31372 2480 31428
rect 2400 31108 2480 31372
rect 2400 31052 2412 31108
rect 2468 31052 2480 31108
rect 2400 30788 2480 31052
rect 2400 30732 2412 30788
rect 2468 30732 2480 30788
rect 2400 30468 2480 30732
rect 2400 30412 2412 30468
rect 2468 30412 2480 30468
rect 2400 30400 2480 30412
rect 2560 32388 2640 32400
rect 2560 32332 2572 32388
rect 2628 32332 2640 32388
rect 2560 32068 2640 32332
rect 2560 32012 2572 32068
rect 2628 32012 2640 32068
rect 2560 31748 2640 32012
rect 2560 31692 2572 31748
rect 2628 31692 2640 31748
rect 2560 31428 2640 31692
rect 2560 31372 2572 31428
rect 2628 31372 2640 31428
rect 2560 31108 2640 31372
rect 2560 31052 2572 31108
rect 2628 31052 2640 31108
rect 2560 30788 2640 31052
rect 2560 30732 2572 30788
rect 2628 30732 2640 30788
rect 2560 30468 2640 30732
rect 2560 30412 2572 30468
rect 2628 30412 2640 30468
rect 2560 30400 2640 30412
rect 2720 32388 2800 32400
rect 2720 32332 2732 32388
rect 2788 32332 2800 32388
rect 2720 32068 2800 32332
rect 2720 32012 2732 32068
rect 2788 32012 2800 32068
rect 2720 31748 2800 32012
rect 2720 31692 2732 31748
rect 2788 31692 2800 31748
rect 2720 31428 2800 31692
rect 2720 31372 2732 31428
rect 2788 31372 2800 31428
rect 2720 31108 2800 31372
rect 2720 31052 2732 31108
rect 2788 31052 2800 31108
rect 2720 30788 2800 31052
rect 2720 30732 2732 30788
rect 2788 30732 2800 30788
rect 2720 30468 2800 30732
rect 2720 30412 2732 30468
rect 2788 30412 2800 30468
rect 2720 30400 2800 30412
rect 2880 32388 2960 32400
rect 2880 32332 2892 32388
rect 2948 32332 2960 32388
rect 2880 32068 2960 32332
rect 2880 32012 2892 32068
rect 2948 32012 2960 32068
rect 2880 31748 2960 32012
rect 2880 31692 2892 31748
rect 2948 31692 2960 31748
rect 2880 31428 2960 31692
rect 2880 31372 2892 31428
rect 2948 31372 2960 31428
rect 2880 31108 2960 31372
rect 2880 31052 2892 31108
rect 2948 31052 2960 31108
rect 2880 30788 2960 31052
rect 2880 30732 2892 30788
rect 2948 30732 2960 30788
rect 2880 30468 2960 30732
rect 2880 30412 2892 30468
rect 2948 30412 2960 30468
rect 2880 30400 2960 30412
rect 3040 32388 3120 32400
rect 3040 32332 3052 32388
rect 3108 32332 3120 32388
rect 3040 32068 3120 32332
rect 3040 32012 3052 32068
rect 3108 32012 3120 32068
rect 3040 31748 3120 32012
rect 3040 31692 3052 31748
rect 3108 31692 3120 31748
rect 3040 31428 3120 31692
rect 3040 31372 3052 31428
rect 3108 31372 3120 31428
rect 3040 31108 3120 31372
rect 3040 31052 3052 31108
rect 3108 31052 3120 31108
rect 3040 30788 3120 31052
rect 3040 30732 3052 30788
rect 3108 30732 3120 30788
rect 3040 30468 3120 30732
rect 3040 30412 3052 30468
rect 3108 30412 3120 30468
rect 3040 30400 3120 30412
rect 3200 32388 3280 32400
rect 3200 32332 3212 32388
rect 3268 32332 3280 32388
rect 3200 32068 3280 32332
rect 3200 32012 3212 32068
rect 3268 32012 3280 32068
rect 3200 31748 3280 32012
rect 3200 31692 3212 31748
rect 3268 31692 3280 31748
rect 3200 31428 3280 31692
rect 3200 31372 3212 31428
rect 3268 31372 3280 31428
rect 3200 31108 3280 31372
rect 3200 31052 3212 31108
rect 3268 31052 3280 31108
rect 3200 30788 3280 31052
rect 3200 30732 3212 30788
rect 3268 30732 3280 30788
rect 3200 30468 3280 30732
rect 3200 30412 3212 30468
rect 3268 30412 3280 30468
rect 3200 30400 3280 30412
rect 3360 32388 3440 32400
rect 3360 32332 3372 32388
rect 3428 32332 3440 32388
rect 3360 32068 3440 32332
rect 3360 32012 3372 32068
rect 3428 32012 3440 32068
rect 3360 31748 3440 32012
rect 3360 31692 3372 31748
rect 3428 31692 3440 31748
rect 3360 31428 3440 31692
rect 3360 31372 3372 31428
rect 3428 31372 3440 31428
rect 3360 31108 3440 31372
rect 3360 31052 3372 31108
rect 3428 31052 3440 31108
rect 3360 30788 3440 31052
rect 3360 30732 3372 30788
rect 3428 30732 3440 30788
rect 3360 30468 3440 30732
rect 3360 30412 3372 30468
rect 3428 30412 3440 30468
rect 3360 30400 3440 30412
rect 3520 32388 3600 32400
rect 3520 32332 3532 32388
rect 3588 32332 3600 32388
rect 3520 32068 3600 32332
rect 3520 32012 3532 32068
rect 3588 32012 3600 32068
rect 3520 31748 3600 32012
rect 3520 31692 3532 31748
rect 3588 31692 3600 31748
rect 3520 31428 3600 31692
rect 3520 31372 3532 31428
rect 3588 31372 3600 31428
rect 3520 31108 3600 31372
rect 3520 31052 3532 31108
rect 3588 31052 3600 31108
rect 3520 30788 3600 31052
rect 3520 30732 3532 30788
rect 3588 30732 3600 30788
rect 3520 30468 3600 30732
rect 3520 30412 3532 30468
rect 3588 30412 3600 30468
rect 3520 30400 3600 30412
rect 3680 32388 3760 32400
rect 3680 32332 3692 32388
rect 3748 32332 3760 32388
rect 3680 32068 3760 32332
rect 3680 32012 3692 32068
rect 3748 32012 3760 32068
rect 3680 31748 3760 32012
rect 3680 31692 3692 31748
rect 3748 31692 3760 31748
rect 3680 31428 3760 31692
rect 3680 31372 3692 31428
rect 3748 31372 3760 31428
rect 3680 31108 3760 31372
rect 3680 31052 3692 31108
rect 3748 31052 3760 31108
rect 3680 30788 3760 31052
rect 3680 30732 3692 30788
rect 3748 30732 3760 30788
rect 3680 30468 3760 30732
rect 3680 30412 3692 30468
rect 3748 30412 3760 30468
rect 3680 30400 3760 30412
rect 3840 32388 3920 32400
rect 3840 32332 3852 32388
rect 3908 32332 3920 32388
rect 3840 32068 3920 32332
rect 3840 32012 3852 32068
rect 3908 32012 3920 32068
rect 3840 31748 3920 32012
rect 3840 31692 3852 31748
rect 3908 31692 3920 31748
rect 3840 31428 3920 31692
rect 3840 31372 3852 31428
rect 3908 31372 3920 31428
rect 3840 31108 3920 31372
rect 3840 31052 3852 31108
rect 3908 31052 3920 31108
rect 3840 30788 3920 31052
rect 3840 30732 3852 30788
rect 3908 30732 3920 30788
rect 3840 30468 3920 30732
rect 3840 30412 3852 30468
rect 3908 30412 3920 30468
rect 3840 30400 3920 30412
rect 4000 32388 4080 32400
rect 4000 32332 4012 32388
rect 4068 32332 4080 32388
rect 4000 32068 4080 32332
rect 4000 32012 4012 32068
rect 4068 32012 4080 32068
rect 4000 31748 4080 32012
rect 4000 31692 4012 31748
rect 4068 31692 4080 31748
rect 4000 31428 4080 31692
rect 4000 31372 4012 31428
rect 4068 31372 4080 31428
rect 4000 31108 4080 31372
rect 4000 31052 4012 31108
rect 4068 31052 4080 31108
rect 4000 30788 4080 31052
rect 4000 30732 4012 30788
rect 4068 30732 4080 30788
rect 4000 30468 4080 30732
rect 4000 30412 4012 30468
rect 4068 30412 4080 30468
rect 4000 30400 4080 30412
rect 4160 32388 4240 32400
rect 4160 32332 4172 32388
rect 4228 32332 4240 32388
rect 4160 32068 4240 32332
rect 4160 32012 4172 32068
rect 4228 32012 4240 32068
rect 4160 31748 4240 32012
rect 4160 31692 4172 31748
rect 4228 31692 4240 31748
rect 4160 31428 4240 31692
rect 4160 31372 4172 31428
rect 4228 31372 4240 31428
rect 4160 31108 4240 31372
rect 4160 31052 4172 31108
rect 4228 31052 4240 31108
rect 4160 30788 4240 31052
rect 4160 30732 4172 30788
rect 4228 30732 4240 30788
rect 4160 30468 4240 30732
rect 4160 30412 4172 30468
rect 4228 30412 4240 30468
rect 4160 30400 4240 30412
rect 4320 32388 4400 32400
rect 4320 32332 4332 32388
rect 4388 32332 4400 32388
rect 4320 32068 4400 32332
rect 4320 32012 4332 32068
rect 4388 32012 4400 32068
rect 4320 31748 4400 32012
rect 4320 31692 4332 31748
rect 4388 31692 4400 31748
rect 4320 31428 4400 31692
rect 4320 31372 4332 31428
rect 4388 31372 4400 31428
rect 4320 31108 4400 31372
rect 4320 31052 4332 31108
rect 4388 31052 4400 31108
rect 4320 30788 4400 31052
rect 4320 30732 4332 30788
rect 4388 30732 4400 30788
rect 4320 30468 4400 30732
rect 4320 30412 4332 30468
rect 4388 30412 4400 30468
rect 4320 30400 4400 30412
rect 4480 32388 4560 32400
rect 4480 32332 4492 32388
rect 4548 32332 4560 32388
rect 4480 32068 4560 32332
rect 4480 32012 4492 32068
rect 4548 32012 4560 32068
rect 4480 31748 4560 32012
rect 4480 31692 4492 31748
rect 4548 31692 4560 31748
rect 4480 31428 4560 31692
rect 4480 31372 4492 31428
rect 4548 31372 4560 31428
rect 4480 31108 4560 31372
rect 4480 31052 4492 31108
rect 4548 31052 4560 31108
rect 4480 30788 4560 31052
rect 4480 30732 4492 30788
rect 4548 30732 4560 30788
rect 4480 30468 4560 30732
rect 4480 30412 4492 30468
rect 4548 30412 4560 30468
rect 4480 30400 4560 30412
rect 4640 32388 4720 32400
rect 4640 32332 4652 32388
rect 4708 32332 4720 32388
rect 4640 32068 4720 32332
rect 4640 32012 4652 32068
rect 4708 32012 4720 32068
rect 4640 31748 4720 32012
rect 4640 31692 4652 31748
rect 4708 31692 4720 31748
rect 4640 31428 4720 31692
rect 4640 31372 4652 31428
rect 4708 31372 4720 31428
rect 4640 31108 4720 31372
rect 4640 31052 4652 31108
rect 4708 31052 4720 31108
rect 4640 30788 4720 31052
rect 4640 30732 4652 30788
rect 4708 30732 4720 30788
rect 4640 30468 4720 30732
rect 4640 30412 4652 30468
rect 4708 30412 4720 30468
rect 4640 30400 4720 30412
rect 4800 32388 4880 32400
rect 4800 32332 4812 32388
rect 4868 32332 4880 32388
rect 4800 32068 4880 32332
rect 4800 32012 4812 32068
rect 4868 32012 4880 32068
rect 4800 31748 4880 32012
rect 4800 31692 4812 31748
rect 4868 31692 4880 31748
rect 4800 31428 4880 31692
rect 4800 31372 4812 31428
rect 4868 31372 4880 31428
rect 4800 31108 4880 31372
rect 4800 31052 4812 31108
rect 4868 31052 4880 31108
rect 4800 30788 4880 31052
rect 4800 30732 4812 30788
rect 4868 30732 4880 30788
rect 4800 30468 4880 30732
rect 4800 30412 4812 30468
rect 4868 30412 4880 30468
rect 4800 30400 4880 30412
rect 4960 32388 5040 32400
rect 4960 32332 4972 32388
rect 5028 32332 5040 32388
rect 4960 32068 5040 32332
rect 4960 32012 4972 32068
rect 5028 32012 5040 32068
rect 4960 31748 5040 32012
rect 4960 31692 4972 31748
rect 5028 31692 5040 31748
rect 4960 31428 5040 31692
rect 4960 31372 4972 31428
rect 5028 31372 5040 31428
rect 4960 31108 5040 31372
rect 4960 31052 4972 31108
rect 5028 31052 5040 31108
rect 4960 30788 5040 31052
rect 4960 30732 4972 30788
rect 5028 30732 5040 30788
rect 4960 30468 5040 30732
rect 4960 30412 4972 30468
rect 5028 30412 5040 30468
rect 4960 30400 5040 30412
rect 5120 32388 5200 32400
rect 5120 32332 5132 32388
rect 5188 32332 5200 32388
rect 5120 32068 5200 32332
rect 5120 32012 5132 32068
rect 5188 32012 5200 32068
rect 5120 31748 5200 32012
rect 5120 31692 5132 31748
rect 5188 31692 5200 31748
rect 5120 31428 5200 31692
rect 5120 31372 5132 31428
rect 5188 31372 5200 31428
rect 5120 31108 5200 31372
rect 5120 31052 5132 31108
rect 5188 31052 5200 31108
rect 5120 30788 5200 31052
rect 5120 30732 5132 30788
rect 5188 30732 5200 30788
rect 5120 30468 5200 30732
rect 5120 30412 5132 30468
rect 5188 30412 5200 30468
rect 5120 30400 5200 30412
rect 5280 32388 5360 32400
rect 5280 32332 5292 32388
rect 5348 32332 5360 32388
rect 5280 32068 5360 32332
rect 5280 32012 5292 32068
rect 5348 32012 5360 32068
rect 5280 31748 5360 32012
rect 5280 31692 5292 31748
rect 5348 31692 5360 31748
rect 5280 31428 5360 31692
rect 5280 31372 5292 31428
rect 5348 31372 5360 31428
rect 5280 31108 5360 31372
rect 5280 31052 5292 31108
rect 5348 31052 5360 31108
rect 5280 30788 5360 31052
rect 5280 30732 5292 30788
rect 5348 30732 5360 30788
rect 5280 30468 5360 30732
rect 5280 30412 5292 30468
rect 5348 30412 5360 30468
rect 5280 30400 5360 30412
rect 5440 32388 5520 32400
rect 5440 32332 5452 32388
rect 5508 32332 5520 32388
rect 5440 32068 5520 32332
rect 5440 32012 5452 32068
rect 5508 32012 5520 32068
rect 5440 31748 5520 32012
rect 5440 31692 5452 31748
rect 5508 31692 5520 31748
rect 5440 31428 5520 31692
rect 5440 31372 5452 31428
rect 5508 31372 5520 31428
rect 5440 31108 5520 31372
rect 5440 31052 5452 31108
rect 5508 31052 5520 31108
rect 5440 30788 5520 31052
rect 5440 30732 5452 30788
rect 5508 30732 5520 30788
rect 5440 30468 5520 30732
rect 5440 30412 5452 30468
rect 5508 30412 5520 30468
rect 5440 30400 5520 30412
rect 5600 32388 5680 32400
rect 5600 32332 5612 32388
rect 5668 32332 5680 32388
rect 5600 32068 5680 32332
rect 5600 32012 5612 32068
rect 5668 32012 5680 32068
rect 5600 31748 5680 32012
rect 5600 31692 5612 31748
rect 5668 31692 5680 31748
rect 5600 31428 5680 31692
rect 5600 31372 5612 31428
rect 5668 31372 5680 31428
rect 5600 31108 5680 31372
rect 5600 31052 5612 31108
rect 5668 31052 5680 31108
rect 5600 30788 5680 31052
rect 5600 30732 5612 30788
rect 5668 30732 5680 30788
rect 5600 30468 5680 30732
rect 5600 30412 5612 30468
rect 5668 30412 5680 30468
rect 5600 30400 5680 30412
rect 5760 32388 5840 32400
rect 5760 32332 5772 32388
rect 5828 32332 5840 32388
rect 5760 32068 5840 32332
rect 5760 32012 5772 32068
rect 5828 32012 5840 32068
rect 5760 31748 5840 32012
rect 5760 31692 5772 31748
rect 5828 31692 5840 31748
rect 5760 31428 5840 31692
rect 5760 31372 5772 31428
rect 5828 31372 5840 31428
rect 5760 31108 5840 31372
rect 5760 31052 5772 31108
rect 5828 31052 5840 31108
rect 5760 30788 5840 31052
rect 5760 30732 5772 30788
rect 5828 30732 5840 30788
rect 5760 30468 5840 30732
rect 5760 30412 5772 30468
rect 5828 30412 5840 30468
rect 5760 30400 5840 30412
rect 5920 32388 6000 32400
rect 5920 32332 5932 32388
rect 5988 32332 6000 32388
rect 5920 32068 6000 32332
rect 5920 32012 5932 32068
rect 5988 32012 6000 32068
rect 5920 31748 6000 32012
rect 5920 31692 5932 31748
rect 5988 31692 6000 31748
rect 5920 31428 6000 31692
rect 5920 31372 5932 31428
rect 5988 31372 6000 31428
rect 5920 31108 6000 31372
rect 5920 31052 5932 31108
rect 5988 31052 6000 31108
rect 5920 30788 6000 31052
rect 5920 30732 5932 30788
rect 5988 30732 6000 30788
rect 5920 30468 6000 30732
rect 5920 30412 5932 30468
rect 5988 30412 6000 30468
rect 5920 30400 6000 30412
rect 6080 32388 6160 32400
rect 6080 32332 6092 32388
rect 6148 32332 6160 32388
rect 6080 32068 6160 32332
rect 6080 32012 6092 32068
rect 6148 32012 6160 32068
rect 6080 31748 6160 32012
rect 6080 31692 6092 31748
rect 6148 31692 6160 31748
rect 6080 31428 6160 31692
rect 6080 31372 6092 31428
rect 6148 31372 6160 31428
rect 6080 31108 6160 31372
rect 6080 31052 6092 31108
rect 6148 31052 6160 31108
rect 6080 30788 6160 31052
rect 6080 30732 6092 30788
rect 6148 30732 6160 30788
rect 6080 30468 6160 30732
rect 6080 30412 6092 30468
rect 6148 30412 6160 30468
rect 6080 30400 6160 30412
rect 6240 32388 6320 32400
rect 6240 32332 6252 32388
rect 6308 32332 6320 32388
rect 6240 32068 6320 32332
rect 6240 32012 6252 32068
rect 6308 32012 6320 32068
rect 6240 31748 6320 32012
rect 6240 31692 6252 31748
rect 6308 31692 6320 31748
rect 6240 31428 6320 31692
rect 6240 31372 6252 31428
rect 6308 31372 6320 31428
rect 6240 31108 6320 31372
rect 6240 31052 6252 31108
rect 6308 31052 6320 31108
rect 6240 30788 6320 31052
rect 6240 30732 6252 30788
rect 6308 30732 6320 30788
rect 6240 30468 6320 30732
rect 6240 30412 6252 30468
rect 6308 30412 6320 30468
rect 6240 30400 6320 30412
rect 6400 32388 6480 32400
rect 6400 32332 6412 32388
rect 6468 32332 6480 32388
rect 6400 32068 6480 32332
rect 6400 32012 6412 32068
rect 6468 32012 6480 32068
rect 6400 31748 6480 32012
rect 6400 31692 6412 31748
rect 6468 31692 6480 31748
rect 6400 31428 6480 31692
rect 6400 31372 6412 31428
rect 6468 31372 6480 31428
rect 6400 31108 6480 31372
rect 6400 31052 6412 31108
rect 6468 31052 6480 31108
rect 6400 30788 6480 31052
rect 6400 30732 6412 30788
rect 6468 30732 6480 30788
rect 6400 30468 6480 30732
rect 6400 30412 6412 30468
rect 6468 30412 6480 30468
rect 6400 30400 6480 30412
rect 6560 32388 6640 32400
rect 6560 32332 6572 32388
rect 6628 32332 6640 32388
rect 6560 32068 6640 32332
rect 6560 32012 6572 32068
rect 6628 32012 6640 32068
rect 6560 31748 6640 32012
rect 6560 31692 6572 31748
rect 6628 31692 6640 31748
rect 6560 31428 6640 31692
rect 6560 31372 6572 31428
rect 6628 31372 6640 31428
rect 6560 31108 6640 31372
rect 6560 31052 6572 31108
rect 6628 31052 6640 31108
rect 6560 30788 6640 31052
rect 6560 30732 6572 30788
rect 6628 30732 6640 30788
rect 6560 30468 6640 30732
rect 6560 30412 6572 30468
rect 6628 30412 6640 30468
rect 6560 30400 6640 30412
rect 6720 32388 6800 32400
rect 6720 32332 6732 32388
rect 6788 32332 6800 32388
rect 6720 32068 6800 32332
rect 6720 32012 6732 32068
rect 6788 32012 6800 32068
rect 6720 31748 6800 32012
rect 6720 31692 6732 31748
rect 6788 31692 6800 31748
rect 6720 31428 6800 31692
rect 6720 31372 6732 31428
rect 6788 31372 6800 31428
rect 6720 31108 6800 31372
rect 6720 31052 6732 31108
rect 6788 31052 6800 31108
rect 6720 30788 6800 31052
rect 6720 30732 6732 30788
rect 6788 30732 6800 30788
rect 6720 30468 6800 30732
rect 6720 30412 6732 30468
rect 6788 30412 6800 30468
rect 6720 30400 6800 30412
rect 6880 32388 6960 32400
rect 6880 32332 6892 32388
rect 6948 32332 6960 32388
rect 6880 32068 6960 32332
rect 6880 32012 6892 32068
rect 6948 32012 6960 32068
rect 6880 31748 6960 32012
rect 6880 31692 6892 31748
rect 6948 31692 6960 31748
rect 6880 31428 6960 31692
rect 6880 31372 6892 31428
rect 6948 31372 6960 31428
rect 6880 31108 6960 31372
rect 6880 31052 6892 31108
rect 6948 31052 6960 31108
rect 6880 30788 6960 31052
rect 6880 30732 6892 30788
rect 6948 30732 6960 30788
rect 6880 30468 6960 30732
rect 6880 30412 6892 30468
rect 6948 30412 6960 30468
rect 6880 30400 6960 30412
rect 7040 32388 7120 32400
rect 7040 32332 7052 32388
rect 7108 32332 7120 32388
rect 7040 32068 7120 32332
rect 7040 32012 7052 32068
rect 7108 32012 7120 32068
rect 7040 31748 7120 32012
rect 7040 31692 7052 31748
rect 7108 31692 7120 31748
rect 7040 31428 7120 31692
rect 7040 31372 7052 31428
rect 7108 31372 7120 31428
rect 7040 31108 7120 31372
rect 7040 31052 7052 31108
rect 7108 31052 7120 31108
rect 7040 30788 7120 31052
rect 7040 30732 7052 30788
rect 7108 30732 7120 30788
rect 7040 30468 7120 30732
rect 7040 30412 7052 30468
rect 7108 30412 7120 30468
rect 7040 30400 7120 30412
rect 7200 32388 7280 32400
rect 7200 32332 7212 32388
rect 7268 32332 7280 32388
rect 7200 32068 7280 32332
rect 7200 32012 7212 32068
rect 7268 32012 7280 32068
rect 7200 31748 7280 32012
rect 7200 31692 7212 31748
rect 7268 31692 7280 31748
rect 7200 31428 7280 31692
rect 7200 31372 7212 31428
rect 7268 31372 7280 31428
rect 7200 31108 7280 31372
rect 7200 31052 7212 31108
rect 7268 31052 7280 31108
rect 7200 30788 7280 31052
rect 7200 30732 7212 30788
rect 7268 30732 7280 30788
rect 7200 30468 7280 30732
rect 7200 30412 7212 30468
rect 7268 30412 7280 30468
rect 7200 30400 7280 30412
rect 7360 32388 7440 32400
rect 7360 32332 7372 32388
rect 7428 32332 7440 32388
rect 7360 32068 7440 32332
rect 7360 32012 7372 32068
rect 7428 32012 7440 32068
rect 7360 31748 7440 32012
rect 7360 31692 7372 31748
rect 7428 31692 7440 31748
rect 7360 31428 7440 31692
rect 7360 31372 7372 31428
rect 7428 31372 7440 31428
rect 7360 31108 7440 31372
rect 7360 31052 7372 31108
rect 7428 31052 7440 31108
rect 7360 30788 7440 31052
rect 7360 30732 7372 30788
rect 7428 30732 7440 30788
rect 7360 30468 7440 30732
rect 7360 30412 7372 30468
rect 7428 30412 7440 30468
rect 7360 30400 7440 30412
rect 7520 32388 7600 32400
rect 7520 32332 7532 32388
rect 7588 32332 7600 32388
rect 7520 32068 7600 32332
rect 7520 32012 7532 32068
rect 7588 32012 7600 32068
rect 7520 31748 7600 32012
rect 7520 31692 7532 31748
rect 7588 31692 7600 31748
rect 7520 31428 7600 31692
rect 7520 31372 7532 31428
rect 7588 31372 7600 31428
rect 7520 31108 7600 31372
rect 7520 31052 7532 31108
rect 7588 31052 7600 31108
rect 7520 30788 7600 31052
rect 7520 30732 7532 30788
rect 7588 30732 7600 30788
rect 7520 30468 7600 30732
rect 7520 30412 7532 30468
rect 7588 30412 7600 30468
rect 7520 30400 7600 30412
rect 7680 32388 7760 32400
rect 7680 32332 7692 32388
rect 7748 32332 7760 32388
rect 7680 32068 7760 32332
rect 7680 32012 7692 32068
rect 7748 32012 7760 32068
rect 7680 31748 7760 32012
rect 7680 31692 7692 31748
rect 7748 31692 7760 31748
rect 7680 31428 7760 31692
rect 7680 31372 7692 31428
rect 7748 31372 7760 31428
rect 7680 31108 7760 31372
rect 7680 31052 7692 31108
rect 7748 31052 7760 31108
rect 7680 30788 7760 31052
rect 7680 30732 7692 30788
rect 7748 30732 7760 30788
rect 7680 30468 7760 30732
rect 7680 30412 7692 30468
rect 7748 30412 7760 30468
rect 7680 30400 7760 30412
rect 7840 32388 7920 32400
rect 7840 32332 7852 32388
rect 7908 32332 7920 32388
rect 7840 32068 7920 32332
rect 7840 32012 7852 32068
rect 7908 32012 7920 32068
rect 7840 31748 7920 32012
rect 7840 31692 7852 31748
rect 7908 31692 7920 31748
rect 7840 31428 7920 31692
rect 7840 31372 7852 31428
rect 7908 31372 7920 31428
rect 7840 31108 7920 31372
rect 7840 31052 7852 31108
rect 7908 31052 7920 31108
rect 7840 30788 7920 31052
rect 7840 30732 7852 30788
rect 7908 30732 7920 30788
rect 7840 30468 7920 30732
rect 7840 30412 7852 30468
rect 7908 30412 7920 30468
rect 7840 30400 7920 30412
rect 8000 32388 8080 32400
rect 8000 32332 8012 32388
rect 8068 32332 8080 32388
rect 8000 32068 8080 32332
rect 8000 32012 8012 32068
rect 8068 32012 8080 32068
rect 8000 31748 8080 32012
rect 8000 31692 8012 31748
rect 8068 31692 8080 31748
rect 8000 31428 8080 31692
rect 8000 31372 8012 31428
rect 8068 31372 8080 31428
rect 8000 31108 8080 31372
rect 8000 31052 8012 31108
rect 8068 31052 8080 31108
rect 8000 30788 8080 31052
rect 8000 30732 8012 30788
rect 8068 30732 8080 30788
rect 8000 30468 8080 30732
rect 8000 30412 8012 30468
rect 8068 30412 8080 30468
rect 8000 30400 8080 30412
rect 8160 32388 8240 32400
rect 8160 32332 8172 32388
rect 8228 32332 8240 32388
rect 8160 32068 8240 32332
rect 8160 32012 8172 32068
rect 8228 32012 8240 32068
rect 8160 31748 8240 32012
rect 8160 31692 8172 31748
rect 8228 31692 8240 31748
rect 8160 31428 8240 31692
rect 8160 31372 8172 31428
rect 8228 31372 8240 31428
rect 8160 31108 8240 31372
rect 8160 31052 8172 31108
rect 8228 31052 8240 31108
rect 8160 30788 8240 31052
rect 8160 30732 8172 30788
rect 8228 30732 8240 30788
rect 8160 30468 8240 30732
rect 8160 30412 8172 30468
rect 8228 30412 8240 30468
rect 8160 30400 8240 30412
rect 8320 32388 8400 32400
rect 8320 32332 8332 32388
rect 8388 32332 8400 32388
rect 8320 32068 8400 32332
rect 8320 32012 8332 32068
rect 8388 32012 8400 32068
rect 8320 31748 8400 32012
rect 8320 31692 8332 31748
rect 8388 31692 8400 31748
rect 8320 31428 8400 31692
rect 8320 31372 8332 31428
rect 8388 31372 8400 31428
rect 8320 31108 8400 31372
rect 8320 31052 8332 31108
rect 8388 31052 8400 31108
rect 8320 30788 8400 31052
rect 8320 30732 8332 30788
rect 8388 30732 8400 30788
rect 8320 30468 8400 30732
rect 8320 30412 8332 30468
rect 8388 30412 8400 30468
rect 8320 30400 8400 30412
rect 0 30308 80 30320
rect 0 30252 12 30308
rect 68 30252 80 30308
rect 0 29988 80 30252
rect 0 29932 12 29988
rect 68 29932 80 29988
rect 0 29920 80 29932
rect 160 30308 240 30320
rect 160 30252 172 30308
rect 228 30252 240 30308
rect 160 29988 240 30252
rect 160 29932 172 29988
rect 228 29932 240 29988
rect 160 29920 240 29932
rect 320 30308 400 30320
rect 320 30252 332 30308
rect 388 30252 400 30308
rect 320 29988 400 30252
rect 320 29932 332 29988
rect 388 29932 400 29988
rect 320 29920 400 29932
rect 480 30308 560 30320
rect 480 30252 492 30308
rect 548 30252 560 30308
rect 480 29988 560 30252
rect 480 29932 492 29988
rect 548 29932 560 29988
rect 480 29920 560 29932
rect 640 30308 720 30320
rect 640 30252 652 30308
rect 708 30252 720 30308
rect 640 29988 720 30252
rect 640 29932 652 29988
rect 708 29932 720 29988
rect 640 29920 720 29932
rect 800 30308 880 30320
rect 800 30252 812 30308
rect 868 30252 880 30308
rect 800 29988 880 30252
rect 800 29932 812 29988
rect 868 29932 880 29988
rect 800 29920 880 29932
rect 960 30308 1040 30320
rect 960 30252 972 30308
rect 1028 30252 1040 30308
rect 960 29988 1040 30252
rect 960 29932 972 29988
rect 1028 29932 1040 29988
rect 960 29920 1040 29932
rect 1120 30308 1200 30320
rect 1120 30252 1132 30308
rect 1188 30252 1200 30308
rect 1120 29988 1200 30252
rect 1120 29932 1132 29988
rect 1188 29932 1200 29988
rect 1120 29920 1200 29932
rect 1280 30308 1360 30320
rect 1280 30252 1292 30308
rect 1348 30252 1360 30308
rect 1280 29988 1360 30252
rect 1280 29932 1292 29988
rect 1348 29932 1360 29988
rect 1280 29920 1360 29932
rect 1440 30308 1520 30320
rect 1440 30252 1452 30308
rect 1508 30252 1520 30308
rect 1440 29988 1520 30252
rect 1440 29932 1452 29988
rect 1508 29932 1520 29988
rect 1440 29920 1520 29932
rect 1600 30308 1680 30320
rect 1600 30252 1612 30308
rect 1668 30252 1680 30308
rect 1600 29988 1680 30252
rect 1600 29932 1612 29988
rect 1668 29932 1680 29988
rect 1600 29920 1680 29932
rect 1760 30308 1840 30320
rect 1760 30252 1772 30308
rect 1828 30252 1840 30308
rect 1760 29988 1840 30252
rect 1760 29932 1772 29988
rect 1828 29932 1840 29988
rect 1760 29920 1840 29932
rect 1920 30308 2000 30320
rect 1920 30252 1932 30308
rect 1988 30252 2000 30308
rect 1920 29988 2000 30252
rect 1920 29932 1932 29988
rect 1988 29932 2000 29988
rect 1920 29920 2000 29932
rect 2080 30308 2160 30320
rect 2080 30252 2092 30308
rect 2148 30252 2160 30308
rect 2080 29988 2160 30252
rect 2080 29932 2092 29988
rect 2148 29932 2160 29988
rect 2080 29920 2160 29932
rect 2240 30308 2320 30320
rect 2240 30252 2252 30308
rect 2308 30252 2320 30308
rect 2240 29988 2320 30252
rect 2240 29932 2252 29988
rect 2308 29932 2320 29988
rect 2240 29920 2320 29932
rect 2400 30308 2480 30320
rect 2400 30252 2412 30308
rect 2468 30252 2480 30308
rect 2400 29988 2480 30252
rect 2400 29932 2412 29988
rect 2468 29932 2480 29988
rect 2400 29920 2480 29932
rect 2560 30308 2640 30320
rect 2560 30252 2572 30308
rect 2628 30252 2640 30308
rect 2560 29988 2640 30252
rect 2560 29932 2572 29988
rect 2628 29932 2640 29988
rect 2560 29920 2640 29932
rect 2720 30308 2800 30320
rect 2720 30252 2732 30308
rect 2788 30252 2800 30308
rect 2720 29988 2800 30252
rect 2720 29932 2732 29988
rect 2788 29932 2800 29988
rect 2720 29920 2800 29932
rect 2880 30308 2960 30320
rect 2880 30252 2892 30308
rect 2948 30252 2960 30308
rect 2880 29988 2960 30252
rect 2880 29932 2892 29988
rect 2948 29932 2960 29988
rect 2880 29920 2960 29932
rect 3040 30308 3120 30320
rect 3040 30252 3052 30308
rect 3108 30252 3120 30308
rect 3040 29988 3120 30252
rect 3040 29932 3052 29988
rect 3108 29932 3120 29988
rect 3040 29920 3120 29932
rect 3200 30308 3280 30320
rect 3200 30252 3212 30308
rect 3268 30252 3280 30308
rect 3200 29988 3280 30252
rect 3200 29932 3212 29988
rect 3268 29932 3280 29988
rect 3200 29920 3280 29932
rect 3360 30308 3440 30320
rect 3360 30252 3372 30308
rect 3428 30252 3440 30308
rect 3360 29988 3440 30252
rect 3360 29932 3372 29988
rect 3428 29932 3440 29988
rect 3360 29920 3440 29932
rect 3520 30308 3600 30320
rect 3520 30252 3532 30308
rect 3588 30252 3600 30308
rect 3520 29988 3600 30252
rect 3520 29932 3532 29988
rect 3588 29932 3600 29988
rect 3520 29920 3600 29932
rect 3680 30308 3760 30320
rect 3680 30252 3692 30308
rect 3748 30252 3760 30308
rect 3680 29988 3760 30252
rect 3680 29932 3692 29988
rect 3748 29932 3760 29988
rect 3680 29920 3760 29932
rect 3840 30308 3920 30320
rect 3840 30252 3852 30308
rect 3908 30252 3920 30308
rect 3840 29988 3920 30252
rect 3840 29932 3852 29988
rect 3908 29932 3920 29988
rect 3840 29920 3920 29932
rect 4000 30308 4080 30320
rect 4000 30252 4012 30308
rect 4068 30252 4080 30308
rect 4000 29988 4080 30252
rect 4000 29932 4012 29988
rect 4068 29932 4080 29988
rect 4000 29920 4080 29932
rect 4160 30308 4240 30320
rect 4160 30252 4172 30308
rect 4228 30252 4240 30308
rect 4160 29988 4240 30252
rect 4160 29932 4172 29988
rect 4228 29932 4240 29988
rect 4160 29920 4240 29932
rect 4320 30308 4400 30320
rect 4320 30252 4332 30308
rect 4388 30252 4400 30308
rect 4320 29988 4400 30252
rect 4320 29932 4332 29988
rect 4388 29932 4400 29988
rect 4320 29920 4400 29932
rect 4480 30308 4560 30320
rect 4480 30252 4492 30308
rect 4548 30252 4560 30308
rect 4480 29988 4560 30252
rect 4480 29932 4492 29988
rect 4548 29932 4560 29988
rect 4480 29920 4560 29932
rect 4640 30308 4720 30320
rect 4640 30252 4652 30308
rect 4708 30252 4720 30308
rect 4640 29988 4720 30252
rect 4640 29932 4652 29988
rect 4708 29932 4720 29988
rect 4640 29920 4720 29932
rect 4800 30308 4880 30320
rect 4800 30252 4812 30308
rect 4868 30252 4880 30308
rect 4800 29988 4880 30252
rect 4800 29932 4812 29988
rect 4868 29932 4880 29988
rect 4800 29920 4880 29932
rect 4960 30308 5040 30320
rect 4960 30252 4972 30308
rect 5028 30252 5040 30308
rect 4960 29988 5040 30252
rect 4960 29932 4972 29988
rect 5028 29932 5040 29988
rect 4960 29920 5040 29932
rect 5120 30308 5200 30320
rect 5120 30252 5132 30308
rect 5188 30252 5200 30308
rect 5120 29988 5200 30252
rect 5120 29932 5132 29988
rect 5188 29932 5200 29988
rect 5120 29920 5200 29932
rect 5280 30308 5360 30320
rect 5280 30252 5292 30308
rect 5348 30252 5360 30308
rect 5280 29988 5360 30252
rect 5280 29932 5292 29988
rect 5348 29932 5360 29988
rect 5280 29920 5360 29932
rect 5440 30308 5520 30320
rect 5440 30252 5452 30308
rect 5508 30252 5520 30308
rect 5440 29988 5520 30252
rect 5440 29932 5452 29988
rect 5508 29932 5520 29988
rect 5440 29920 5520 29932
rect 5600 30308 5680 30320
rect 5600 30252 5612 30308
rect 5668 30252 5680 30308
rect 5600 29988 5680 30252
rect 5600 29932 5612 29988
rect 5668 29932 5680 29988
rect 5600 29920 5680 29932
rect 5760 30308 5840 30320
rect 5760 30252 5772 30308
rect 5828 30252 5840 30308
rect 5760 29988 5840 30252
rect 5760 29932 5772 29988
rect 5828 29932 5840 29988
rect 5760 29920 5840 29932
rect 5920 30308 6000 30320
rect 5920 30252 5932 30308
rect 5988 30252 6000 30308
rect 5920 29988 6000 30252
rect 5920 29932 5932 29988
rect 5988 29932 6000 29988
rect 5920 29920 6000 29932
rect 6080 30308 6160 30320
rect 6080 30252 6092 30308
rect 6148 30252 6160 30308
rect 6080 29988 6160 30252
rect 6080 29932 6092 29988
rect 6148 29932 6160 29988
rect 6080 29920 6160 29932
rect 6240 30308 6320 30320
rect 6240 30252 6252 30308
rect 6308 30252 6320 30308
rect 6240 29988 6320 30252
rect 6240 29932 6252 29988
rect 6308 29932 6320 29988
rect 6240 29920 6320 29932
rect 6400 30308 6480 30320
rect 6400 30252 6412 30308
rect 6468 30252 6480 30308
rect 6400 29988 6480 30252
rect 6400 29932 6412 29988
rect 6468 29932 6480 29988
rect 6400 29920 6480 29932
rect 6560 30308 6640 30320
rect 6560 30252 6572 30308
rect 6628 30252 6640 30308
rect 6560 29988 6640 30252
rect 6560 29932 6572 29988
rect 6628 29932 6640 29988
rect 6560 29920 6640 29932
rect 6720 30308 6800 30320
rect 6720 30252 6732 30308
rect 6788 30252 6800 30308
rect 6720 29988 6800 30252
rect 6720 29932 6732 29988
rect 6788 29932 6800 29988
rect 6720 29920 6800 29932
rect 6880 30308 6960 30320
rect 6880 30252 6892 30308
rect 6948 30252 6960 30308
rect 6880 29988 6960 30252
rect 6880 29932 6892 29988
rect 6948 29932 6960 29988
rect 6880 29920 6960 29932
rect 7040 30308 7120 30320
rect 7040 30252 7052 30308
rect 7108 30252 7120 30308
rect 7040 29988 7120 30252
rect 7040 29932 7052 29988
rect 7108 29932 7120 29988
rect 7040 29920 7120 29932
rect 7200 30308 7280 30320
rect 7200 30252 7212 30308
rect 7268 30252 7280 30308
rect 7200 29988 7280 30252
rect 7200 29932 7212 29988
rect 7268 29932 7280 29988
rect 7200 29920 7280 29932
rect 7360 30308 7440 30320
rect 7360 30252 7372 30308
rect 7428 30252 7440 30308
rect 7360 29988 7440 30252
rect 7360 29932 7372 29988
rect 7428 29932 7440 29988
rect 7360 29920 7440 29932
rect 7520 30308 7600 30320
rect 7520 30252 7532 30308
rect 7588 30252 7600 30308
rect 7520 29988 7600 30252
rect 7520 29932 7532 29988
rect 7588 29932 7600 29988
rect 7520 29920 7600 29932
rect 7680 30308 7760 30320
rect 7680 30252 7692 30308
rect 7748 30252 7760 30308
rect 7680 29988 7760 30252
rect 7680 29932 7692 29988
rect 7748 29932 7760 29988
rect 7680 29920 7760 29932
rect 7840 30308 7920 30320
rect 7840 30252 7852 30308
rect 7908 30252 7920 30308
rect 7840 29988 7920 30252
rect 7840 29932 7852 29988
rect 7908 29932 7920 29988
rect 7840 29920 7920 29932
rect 8000 30308 8080 30320
rect 8000 30252 8012 30308
rect 8068 30252 8080 30308
rect 8000 29988 8080 30252
rect 8000 29932 8012 29988
rect 8068 29932 8080 29988
rect 8000 29920 8080 29932
rect 8160 30308 8240 30320
rect 8160 30252 8172 30308
rect 8228 30252 8240 30308
rect 8160 29988 8240 30252
rect 8160 29932 8172 29988
rect 8228 29932 8240 29988
rect 8160 29920 8240 29932
rect 8320 30308 8400 30320
rect 8320 30252 8332 30308
rect 8388 30252 8400 30308
rect 8320 29988 8400 30252
rect 8320 29932 8332 29988
rect 8388 29932 8400 29988
rect 8320 29920 8400 29932
rect 0 29828 80 29840
rect 0 29772 12 29828
rect 68 29772 80 29828
rect 0 29508 80 29772
rect 0 29452 12 29508
rect 68 29452 80 29508
rect 0 29440 80 29452
rect 160 29828 240 29840
rect 160 29772 172 29828
rect 228 29772 240 29828
rect 160 29508 240 29772
rect 160 29452 172 29508
rect 228 29452 240 29508
rect 160 29440 240 29452
rect 320 29828 400 29840
rect 320 29772 332 29828
rect 388 29772 400 29828
rect 320 29508 400 29772
rect 320 29452 332 29508
rect 388 29452 400 29508
rect 320 29440 400 29452
rect 480 29828 560 29840
rect 480 29772 492 29828
rect 548 29772 560 29828
rect 480 29508 560 29772
rect 480 29452 492 29508
rect 548 29452 560 29508
rect 480 29440 560 29452
rect 640 29828 720 29840
rect 640 29772 652 29828
rect 708 29772 720 29828
rect 640 29508 720 29772
rect 640 29452 652 29508
rect 708 29452 720 29508
rect 640 29440 720 29452
rect 800 29828 880 29840
rect 800 29772 812 29828
rect 868 29772 880 29828
rect 800 29508 880 29772
rect 800 29452 812 29508
rect 868 29452 880 29508
rect 800 29440 880 29452
rect 960 29828 1040 29840
rect 960 29772 972 29828
rect 1028 29772 1040 29828
rect 960 29508 1040 29772
rect 960 29452 972 29508
rect 1028 29452 1040 29508
rect 960 29440 1040 29452
rect 1120 29828 1200 29840
rect 1120 29772 1132 29828
rect 1188 29772 1200 29828
rect 1120 29508 1200 29772
rect 1120 29452 1132 29508
rect 1188 29452 1200 29508
rect 1120 29440 1200 29452
rect 1280 29828 1360 29840
rect 1280 29772 1292 29828
rect 1348 29772 1360 29828
rect 1280 29508 1360 29772
rect 1280 29452 1292 29508
rect 1348 29452 1360 29508
rect 1280 29440 1360 29452
rect 1440 29828 1520 29840
rect 1440 29772 1452 29828
rect 1508 29772 1520 29828
rect 1440 29508 1520 29772
rect 1440 29452 1452 29508
rect 1508 29452 1520 29508
rect 1440 29440 1520 29452
rect 1600 29828 1680 29840
rect 1600 29772 1612 29828
rect 1668 29772 1680 29828
rect 1600 29508 1680 29772
rect 1600 29452 1612 29508
rect 1668 29452 1680 29508
rect 1600 29440 1680 29452
rect 1760 29828 1840 29840
rect 1760 29772 1772 29828
rect 1828 29772 1840 29828
rect 1760 29508 1840 29772
rect 1760 29452 1772 29508
rect 1828 29452 1840 29508
rect 1760 29440 1840 29452
rect 1920 29828 2000 29840
rect 1920 29772 1932 29828
rect 1988 29772 2000 29828
rect 1920 29508 2000 29772
rect 1920 29452 1932 29508
rect 1988 29452 2000 29508
rect 1920 29440 2000 29452
rect 2080 29828 2160 29840
rect 2080 29772 2092 29828
rect 2148 29772 2160 29828
rect 2080 29508 2160 29772
rect 2080 29452 2092 29508
rect 2148 29452 2160 29508
rect 2080 29440 2160 29452
rect 2240 29828 2320 29840
rect 2240 29772 2252 29828
rect 2308 29772 2320 29828
rect 2240 29508 2320 29772
rect 2240 29452 2252 29508
rect 2308 29452 2320 29508
rect 2240 29440 2320 29452
rect 2400 29828 2480 29840
rect 2400 29772 2412 29828
rect 2468 29772 2480 29828
rect 2400 29508 2480 29772
rect 2400 29452 2412 29508
rect 2468 29452 2480 29508
rect 2400 29440 2480 29452
rect 2560 29828 2640 29840
rect 2560 29772 2572 29828
rect 2628 29772 2640 29828
rect 2560 29508 2640 29772
rect 2560 29452 2572 29508
rect 2628 29452 2640 29508
rect 2560 29440 2640 29452
rect 2720 29828 2800 29840
rect 2720 29772 2732 29828
rect 2788 29772 2800 29828
rect 2720 29508 2800 29772
rect 2720 29452 2732 29508
rect 2788 29452 2800 29508
rect 2720 29440 2800 29452
rect 2880 29828 2960 29840
rect 2880 29772 2892 29828
rect 2948 29772 2960 29828
rect 2880 29508 2960 29772
rect 2880 29452 2892 29508
rect 2948 29452 2960 29508
rect 2880 29440 2960 29452
rect 3040 29828 3120 29840
rect 3040 29772 3052 29828
rect 3108 29772 3120 29828
rect 3040 29508 3120 29772
rect 3040 29452 3052 29508
rect 3108 29452 3120 29508
rect 3040 29440 3120 29452
rect 3200 29828 3280 29840
rect 3200 29772 3212 29828
rect 3268 29772 3280 29828
rect 3200 29508 3280 29772
rect 3200 29452 3212 29508
rect 3268 29452 3280 29508
rect 3200 29440 3280 29452
rect 3360 29828 3440 29840
rect 3360 29772 3372 29828
rect 3428 29772 3440 29828
rect 3360 29508 3440 29772
rect 3360 29452 3372 29508
rect 3428 29452 3440 29508
rect 3360 29440 3440 29452
rect 3520 29828 3600 29840
rect 3520 29772 3532 29828
rect 3588 29772 3600 29828
rect 3520 29508 3600 29772
rect 3520 29452 3532 29508
rect 3588 29452 3600 29508
rect 3520 29440 3600 29452
rect 3680 29828 3760 29840
rect 3680 29772 3692 29828
rect 3748 29772 3760 29828
rect 3680 29508 3760 29772
rect 3680 29452 3692 29508
rect 3748 29452 3760 29508
rect 3680 29440 3760 29452
rect 3840 29828 3920 29840
rect 3840 29772 3852 29828
rect 3908 29772 3920 29828
rect 3840 29508 3920 29772
rect 3840 29452 3852 29508
rect 3908 29452 3920 29508
rect 3840 29440 3920 29452
rect 4000 29828 4080 29840
rect 4000 29772 4012 29828
rect 4068 29772 4080 29828
rect 4000 29508 4080 29772
rect 4000 29452 4012 29508
rect 4068 29452 4080 29508
rect 4000 29440 4080 29452
rect 4160 29828 4240 29840
rect 4160 29772 4172 29828
rect 4228 29772 4240 29828
rect 4160 29508 4240 29772
rect 4160 29452 4172 29508
rect 4228 29452 4240 29508
rect 4160 29440 4240 29452
rect 4320 29828 4400 29840
rect 4320 29772 4332 29828
rect 4388 29772 4400 29828
rect 4320 29508 4400 29772
rect 4320 29452 4332 29508
rect 4388 29452 4400 29508
rect 4320 29440 4400 29452
rect 4480 29828 4560 29840
rect 4480 29772 4492 29828
rect 4548 29772 4560 29828
rect 4480 29508 4560 29772
rect 4480 29452 4492 29508
rect 4548 29452 4560 29508
rect 4480 29440 4560 29452
rect 4640 29828 4720 29840
rect 4640 29772 4652 29828
rect 4708 29772 4720 29828
rect 4640 29508 4720 29772
rect 4640 29452 4652 29508
rect 4708 29452 4720 29508
rect 4640 29440 4720 29452
rect 4800 29828 4880 29840
rect 4800 29772 4812 29828
rect 4868 29772 4880 29828
rect 4800 29508 4880 29772
rect 4800 29452 4812 29508
rect 4868 29452 4880 29508
rect 4800 29440 4880 29452
rect 4960 29828 5040 29840
rect 4960 29772 4972 29828
rect 5028 29772 5040 29828
rect 4960 29508 5040 29772
rect 4960 29452 4972 29508
rect 5028 29452 5040 29508
rect 4960 29440 5040 29452
rect 5120 29828 5200 29840
rect 5120 29772 5132 29828
rect 5188 29772 5200 29828
rect 5120 29508 5200 29772
rect 5120 29452 5132 29508
rect 5188 29452 5200 29508
rect 5120 29440 5200 29452
rect 5280 29828 5360 29840
rect 5280 29772 5292 29828
rect 5348 29772 5360 29828
rect 5280 29508 5360 29772
rect 5280 29452 5292 29508
rect 5348 29452 5360 29508
rect 5280 29440 5360 29452
rect 5440 29828 5520 29840
rect 5440 29772 5452 29828
rect 5508 29772 5520 29828
rect 5440 29508 5520 29772
rect 5440 29452 5452 29508
rect 5508 29452 5520 29508
rect 5440 29440 5520 29452
rect 5600 29828 5680 29840
rect 5600 29772 5612 29828
rect 5668 29772 5680 29828
rect 5600 29508 5680 29772
rect 5600 29452 5612 29508
rect 5668 29452 5680 29508
rect 5600 29440 5680 29452
rect 5760 29828 5840 29840
rect 5760 29772 5772 29828
rect 5828 29772 5840 29828
rect 5760 29508 5840 29772
rect 5760 29452 5772 29508
rect 5828 29452 5840 29508
rect 5760 29440 5840 29452
rect 5920 29828 6000 29840
rect 5920 29772 5932 29828
rect 5988 29772 6000 29828
rect 5920 29508 6000 29772
rect 5920 29452 5932 29508
rect 5988 29452 6000 29508
rect 5920 29440 6000 29452
rect 6080 29828 6160 29840
rect 6080 29772 6092 29828
rect 6148 29772 6160 29828
rect 6080 29508 6160 29772
rect 6080 29452 6092 29508
rect 6148 29452 6160 29508
rect 6080 29440 6160 29452
rect 6240 29828 6320 29840
rect 6240 29772 6252 29828
rect 6308 29772 6320 29828
rect 6240 29508 6320 29772
rect 6240 29452 6252 29508
rect 6308 29452 6320 29508
rect 6240 29440 6320 29452
rect 6400 29828 6480 29840
rect 6400 29772 6412 29828
rect 6468 29772 6480 29828
rect 6400 29508 6480 29772
rect 6400 29452 6412 29508
rect 6468 29452 6480 29508
rect 6400 29440 6480 29452
rect 6560 29828 6640 29840
rect 6560 29772 6572 29828
rect 6628 29772 6640 29828
rect 6560 29508 6640 29772
rect 6560 29452 6572 29508
rect 6628 29452 6640 29508
rect 6560 29440 6640 29452
rect 6720 29828 6800 29840
rect 6720 29772 6732 29828
rect 6788 29772 6800 29828
rect 6720 29508 6800 29772
rect 6720 29452 6732 29508
rect 6788 29452 6800 29508
rect 6720 29440 6800 29452
rect 6880 29828 6960 29840
rect 6880 29772 6892 29828
rect 6948 29772 6960 29828
rect 6880 29508 6960 29772
rect 6880 29452 6892 29508
rect 6948 29452 6960 29508
rect 6880 29440 6960 29452
rect 7040 29828 7120 29840
rect 7040 29772 7052 29828
rect 7108 29772 7120 29828
rect 7040 29508 7120 29772
rect 7040 29452 7052 29508
rect 7108 29452 7120 29508
rect 7040 29440 7120 29452
rect 7200 29828 7280 29840
rect 7200 29772 7212 29828
rect 7268 29772 7280 29828
rect 7200 29508 7280 29772
rect 7200 29452 7212 29508
rect 7268 29452 7280 29508
rect 7200 29440 7280 29452
rect 7360 29828 7440 29840
rect 7360 29772 7372 29828
rect 7428 29772 7440 29828
rect 7360 29508 7440 29772
rect 7360 29452 7372 29508
rect 7428 29452 7440 29508
rect 7360 29440 7440 29452
rect 7520 29828 7600 29840
rect 7520 29772 7532 29828
rect 7588 29772 7600 29828
rect 7520 29508 7600 29772
rect 7520 29452 7532 29508
rect 7588 29452 7600 29508
rect 7520 29440 7600 29452
rect 7680 29828 7760 29840
rect 7680 29772 7692 29828
rect 7748 29772 7760 29828
rect 7680 29508 7760 29772
rect 7680 29452 7692 29508
rect 7748 29452 7760 29508
rect 7680 29440 7760 29452
rect 7840 29828 7920 29840
rect 7840 29772 7852 29828
rect 7908 29772 7920 29828
rect 7840 29508 7920 29772
rect 7840 29452 7852 29508
rect 7908 29452 7920 29508
rect 7840 29440 7920 29452
rect 8000 29828 8080 29840
rect 8000 29772 8012 29828
rect 8068 29772 8080 29828
rect 8000 29508 8080 29772
rect 8000 29452 8012 29508
rect 8068 29452 8080 29508
rect 8000 29440 8080 29452
rect 8160 29828 8240 29840
rect 8160 29772 8172 29828
rect 8228 29772 8240 29828
rect 8160 29508 8240 29772
rect 8160 29452 8172 29508
rect 8228 29452 8240 29508
rect 8160 29440 8240 29452
rect 8320 29828 8400 29840
rect 8320 29772 8332 29828
rect 8388 29772 8400 29828
rect 8320 29508 8400 29772
rect 8320 29452 8332 29508
rect 8388 29452 8400 29508
rect 8320 29440 8400 29452
rect 8480 29360 8560 32972
rect 8640 33188 8720 33360
rect 8640 33132 8652 33188
rect 8708 33132 8720 33188
rect 8640 29360 8720 33132
rect 8800 33348 8880 33360
rect 8800 33292 8812 33348
rect 8868 33292 8880 33348
rect 8800 33028 8880 33292
rect 8800 32972 8812 33028
rect 8868 32972 8880 33028
rect 8800 29360 8880 32972
rect 8960 32868 9040 33360
rect 8960 32812 8972 32868
rect 9028 32812 9040 32868
rect 8960 32548 9040 32812
rect 8960 32492 8972 32548
rect 9028 32492 9040 32548
rect 8960 29360 9040 32492
rect 9120 32708 9200 33360
rect 9120 32652 9132 32708
rect 9188 32652 9200 32708
rect 9120 29360 9200 32652
rect 9280 32868 9360 33360
rect 9280 32812 9292 32868
rect 9348 32812 9360 32868
rect 9280 32548 9360 32812
rect 9280 32492 9292 32548
rect 9348 32492 9360 32548
rect 9280 29360 9360 32492
rect 9440 32388 9520 33360
rect 9440 32332 9452 32388
rect 9508 32332 9520 32388
rect 9440 32068 9520 32332
rect 9440 32012 9452 32068
rect 9508 32012 9520 32068
rect 9440 31748 9520 32012
rect 9440 31692 9452 31748
rect 9508 31692 9520 31748
rect 9440 31428 9520 31692
rect 9440 31372 9452 31428
rect 9508 31372 9520 31428
rect 9440 31108 9520 31372
rect 9440 31052 9452 31108
rect 9508 31052 9520 31108
rect 9440 30788 9520 31052
rect 9440 30732 9452 30788
rect 9508 30732 9520 30788
rect 9440 30468 9520 30732
rect 9440 30412 9452 30468
rect 9508 30412 9520 30468
rect 9440 29360 9520 30412
rect 9600 32228 9680 33360
rect 9600 32172 9612 32228
rect 9668 32172 9680 32228
rect 9600 29360 9680 32172
rect 9760 32388 9840 33360
rect 9760 32332 9772 32388
rect 9828 32332 9840 32388
rect 9760 32068 9840 32332
rect 9760 32012 9772 32068
rect 9828 32012 9840 32068
rect 9760 31748 9840 32012
rect 9760 31692 9772 31748
rect 9828 31692 9840 31748
rect 9760 31428 9840 31692
rect 9760 31372 9772 31428
rect 9828 31372 9840 31428
rect 9760 31108 9840 31372
rect 9760 31052 9772 31108
rect 9828 31052 9840 31108
rect 9760 30788 9840 31052
rect 9760 30732 9772 30788
rect 9828 30732 9840 30788
rect 9760 30468 9840 30732
rect 9760 30412 9772 30468
rect 9828 30412 9840 30468
rect 9760 29360 9840 30412
rect 9920 31908 10000 33360
rect 9920 31852 9932 31908
rect 9988 31852 10000 31908
rect 9920 29360 10000 31852
rect 10080 32388 10160 33360
rect 10080 32332 10092 32388
rect 10148 32332 10160 32388
rect 10080 32068 10160 32332
rect 10080 32012 10092 32068
rect 10148 32012 10160 32068
rect 10080 31748 10160 32012
rect 10080 31692 10092 31748
rect 10148 31692 10160 31748
rect 10080 31428 10160 31692
rect 10080 31372 10092 31428
rect 10148 31372 10160 31428
rect 10080 31108 10160 31372
rect 10080 31052 10092 31108
rect 10148 31052 10160 31108
rect 10080 30788 10160 31052
rect 10080 30732 10092 30788
rect 10148 30732 10160 30788
rect 10080 30468 10160 30732
rect 10080 30412 10092 30468
rect 10148 30412 10160 30468
rect 10080 29360 10160 30412
rect 10240 31588 10320 33360
rect 10240 31532 10252 31588
rect 10308 31532 10320 31588
rect 10240 29360 10320 31532
rect 10400 32388 10480 33360
rect 10400 32332 10412 32388
rect 10468 32332 10480 32388
rect 10400 32068 10480 32332
rect 10400 32012 10412 32068
rect 10468 32012 10480 32068
rect 10400 31748 10480 32012
rect 10400 31692 10412 31748
rect 10468 31692 10480 31748
rect 10400 31428 10480 31692
rect 10400 31372 10412 31428
rect 10468 31372 10480 31428
rect 10400 31108 10480 31372
rect 10400 31052 10412 31108
rect 10468 31052 10480 31108
rect 10400 30788 10480 31052
rect 10400 30732 10412 30788
rect 10468 30732 10480 30788
rect 10400 30468 10480 30732
rect 10400 30412 10412 30468
rect 10468 30412 10480 30468
rect 10400 29360 10480 30412
rect 10560 31268 10640 33360
rect 10560 31212 10572 31268
rect 10628 31212 10640 31268
rect 10560 29360 10640 31212
rect 10720 32388 10800 33360
rect 10720 32332 10732 32388
rect 10788 32332 10800 32388
rect 10720 32068 10800 32332
rect 10720 32012 10732 32068
rect 10788 32012 10800 32068
rect 10720 31748 10800 32012
rect 10720 31692 10732 31748
rect 10788 31692 10800 31748
rect 10720 31428 10800 31692
rect 10720 31372 10732 31428
rect 10788 31372 10800 31428
rect 10720 31108 10800 31372
rect 10720 31052 10732 31108
rect 10788 31052 10800 31108
rect 10720 30788 10800 31052
rect 10720 30732 10732 30788
rect 10788 30732 10800 30788
rect 10720 30468 10800 30732
rect 10720 30412 10732 30468
rect 10788 30412 10800 30468
rect 10720 29360 10800 30412
rect 10880 30948 10960 33360
rect 10880 30892 10892 30948
rect 10948 30892 10960 30948
rect 10880 29360 10960 30892
rect 11040 32388 11120 33360
rect 11040 32332 11052 32388
rect 11108 32332 11120 32388
rect 11040 32068 11120 32332
rect 11040 32012 11052 32068
rect 11108 32012 11120 32068
rect 11040 31748 11120 32012
rect 11040 31692 11052 31748
rect 11108 31692 11120 31748
rect 11040 31428 11120 31692
rect 11040 31372 11052 31428
rect 11108 31372 11120 31428
rect 11040 31108 11120 31372
rect 11040 31052 11052 31108
rect 11108 31052 11120 31108
rect 11040 30788 11120 31052
rect 11040 30732 11052 30788
rect 11108 30732 11120 30788
rect 11040 30468 11120 30732
rect 11040 30412 11052 30468
rect 11108 30412 11120 30468
rect 11040 29360 11120 30412
rect 11200 30628 11280 33360
rect 11200 30572 11212 30628
rect 11268 30572 11280 30628
rect 11200 29360 11280 30572
rect 11360 32388 11440 33360
rect 11360 32332 11372 32388
rect 11428 32332 11440 32388
rect 11360 32068 11440 32332
rect 11360 32012 11372 32068
rect 11428 32012 11440 32068
rect 11360 31748 11440 32012
rect 11360 31692 11372 31748
rect 11428 31692 11440 31748
rect 11360 31428 11440 31692
rect 11360 31372 11372 31428
rect 11428 31372 11440 31428
rect 11360 31108 11440 31372
rect 11360 31052 11372 31108
rect 11428 31052 11440 31108
rect 11360 30788 11440 31052
rect 11360 30732 11372 30788
rect 11428 30732 11440 30788
rect 11360 30468 11440 30732
rect 11360 30412 11372 30468
rect 11428 30412 11440 30468
rect 11360 29360 11440 30412
rect 11520 30308 11600 33360
rect 11520 30252 11532 30308
rect 11588 30252 11600 30308
rect 11520 29988 11600 30252
rect 11520 29932 11532 29988
rect 11588 29932 11600 29988
rect 11520 29360 11600 29932
rect 11680 30148 11760 33360
rect 11680 30092 11692 30148
rect 11748 30092 11760 30148
rect 11680 29360 11760 30092
rect 11840 30308 11920 33360
rect 11840 30252 11852 30308
rect 11908 30252 11920 30308
rect 11840 29988 11920 30252
rect 11840 29932 11852 29988
rect 11908 29932 11920 29988
rect 11840 29360 11920 29932
rect 12000 29828 12080 33360
rect 12000 29772 12012 29828
rect 12068 29772 12080 29828
rect 12000 29508 12080 29772
rect 12000 29452 12012 29508
rect 12068 29452 12080 29508
rect 12000 29360 12080 29452
rect 12160 29668 12240 33360
rect 12160 29612 12172 29668
rect 12228 29612 12240 29668
rect 12160 29360 12240 29612
rect 12320 29828 12400 33360
rect 12480 33348 12560 33360
rect 12480 33292 12492 33348
rect 12548 33292 12560 33348
rect 12480 33028 12560 33292
rect 12480 32972 12492 33028
rect 12548 32972 12560 33028
rect 12480 32960 12560 32972
rect 12640 33348 12720 33360
rect 12640 33292 12652 33348
rect 12708 33292 12720 33348
rect 12640 33028 12720 33292
rect 12640 32972 12652 33028
rect 12708 32972 12720 33028
rect 12640 32960 12720 32972
rect 12800 33348 12880 33360
rect 12800 33292 12812 33348
rect 12868 33292 12880 33348
rect 12800 33028 12880 33292
rect 12800 32972 12812 33028
rect 12868 32972 12880 33028
rect 12800 32960 12880 32972
rect 12960 33348 13040 33360
rect 12960 33292 12972 33348
rect 13028 33292 13040 33348
rect 12960 33028 13040 33292
rect 12960 32972 12972 33028
rect 13028 32972 13040 33028
rect 12960 32960 13040 32972
rect 13120 33348 13200 33360
rect 13120 33292 13132 33348
rect 13188 33292 13200 33348
rect 13120 33028 13200 33292
rect 13120 32972 13132 33028
rect 13188 32972 13200 33028
rect 13120 32960 13200 32972
rect 13280 33348 13360 33360
rect 13280 33292 13292 33348
rect 13348 33292 13360 33348
rect 13280 33028 13360 33292
rect 13280 32972 13292 33028
rect 13348 32972 13360 33028
rect 13280 32960 13360 32972
rect 13440 33348 13520 33360
rect 13440 33292 13452 33348
rect 13508 33292 13520 33348
rect 13440 33028 13520 33292
rect 13440 32972 13452 33028
rect 13508 32972 13520 33028
rect 13440 32960 13520 32972
rect 13600 33348 13680 33360
rect 13600 33292 13612 33348
rect 13668 33292 13680 33348
rect 13600 33028 13680 33292
rect 13600 32972 13612 33028
rect 13668 32972 13680 33028
rect 13600 32960 13680 32972
rect 13760 33348 13840 33360
rect 13760 33292 13772 33348
rect 13828 33292 13840 33348
rect 13760 33028 13840 33292
rect 13760 32972 13772 33028
rect 13828 32972 13840 33028
rect 13760 32960 13840 32972
rect 13920 33348 14000 33360
rect 13920 33292 13932 33348
rect 13988 33292 14000 33348
rect 13920 33028 14000 33292
rect 13920 32972 13932 33028
rect 13988 32972 14000 33028
rect 13920 32960 14000 32972
rect 14080 33348 14160 33360
rect 14080 33292 14092 33348
rect 14148 33292 14160 33348
rect 14080 33028 14160 33292
rect 14080 32972 14092 33028
rect 14148 32972 14160 33028
rect 14080 32960 14160 32972
rect 14240 33348 14320 33360
rect 14240 33292 14252 33348
rect 14308 33292 14320 33348
rect 14240 33028 14320 33292
rect 14240 32972 14252 33028
rect 14308 32972 14320 33028
rect 14240 32960 14320 32972
rect 14400 33348 14480 33360
rect 14400 33292 14412 33348
rect 14468 33292 14480 33348
rect 14400 33028 14480 33292
rect 14400 32972 14412 33028
rect 14468 32972 14480 33028
rect 14400 32960 14480 32972
rect 14560 33348 14640 33360
rect 14560 33292 14572 33348
rect 14628 33292 14640 33348
rect 14560 33028 14640 33292
rect 14560 32972 14572 33028
rect 14628 32972 14640 33028
rect 14560 32960 14640 32972
rect 14720 33348 14800 33360
rect 14720 33292 14732 33348
rect 14788 33292 14800 33348
rect 14720 33028 14800 33292
rect 14720 32972 14732 33028
rect 14788 32972 14800 33028
rect 14720 32960 14800 32972
rect 14880 33348 14960 33360
rect 14880 33292 14892 33348
rect 14948 33292 14960 33348
rect 14880 33028 14960 33292
rect 14880 32972 14892 33028
rect 14948 32972 14960 33028
rect 14880 32960 14960 32972
rect 15040 33348 15120 33360
rect 15040 33292 15052 33348
rect 15108 33292 15120 33348
rect 15040 33028 15120 33292
rect 15040 32972 15052 33028
rect 15108 32972 15120 33028
rect 15040 32960 15120 32972
rect 15200 33348 15280 33360
rect 15200 33292 15212 33348
rect 15268 33292 15280 33348
rect 15200 33028 15280 33292
rect 15200 32972 15212 33028
rect 15268 32972 15280 33028
rect 15200 32960 15280 32972
rect 15360 33348 15440 33360
rect 15360 33292 15372 33348
rect 15428 33292 15440 33348
rect 15360 33028 15440 33292
rect 15360 32972 15372 33028
rect 15428 32972 15440 33028
rect 15360 32960 15440 32972
rect 15520 33348 15600 33360
rect 15520 33292 15532 33348
rect 15588 33292 15600 33348
rect 15520 33028 15600 33292
rect 15520 32972 15532 33028
rect 15588 32972 15600 33028
rect 15520 32960 15600 32972
rect 15680 33348 15760 33360
rect 15680 33292 15692 33348
rect 15748 33292 15760 33348
rect 15680 33028 15760 33292
rect 15680 32972 15692 33028
rect 15748 32972 15760 33028
rect 15680 32960 15760 32972
rect 15840 33348 15920 33360
rect 15840 33292 15852 33348
rect 15908 33292 15920 33348
rect 15840 33028 15920 33292
rect 15840 32972 15852 33028
rect 15908 32972 15920 33028
rect 15840 32960 15920 32972
rect 16000 33348 16080 33360
rect 16000 33292 16012 33348
rect 16068 33292 16080 33348
rect 16000 33028 16080 33292
rect 16000 32972 16012 33028
rect 16068 32972 16080 33028
rect 16000 32960 16080 32972
rect 16160 33348 16240 33360
rect 16160 33292 16172 33348
rect 16228 33292 16240 33348
rect 16160 33028 16240 33292
rect 16160 32972 16172 33028
rect 16228 32972 16240 33028
rect 16160 32960 16240 32972
rect 16320 33348 16400 33360
rect 16320 33292 16332 33348
rect 16388 33292 16400 33348
rect 16320 33028 16400 33292
rect 16320 32972 16332 33028
rect 16388 32972 16400 33028
rect 16320 32960 16400 32972
rect 16480 33348 16560 33360
rect 16480 33292 16492 33348
rect 16548 33292 16560 33348
rect 16480 33028 16560 33292
rect 16480 32972 16492 33028
rect 16548 32972 16560 33028
rect 16480 32960 16560 32972
rect 16640 33348 16720 33360
rect 16640 33292 16652 33348
rect 16708 33292 16720 33348
rect 16640 33028 16720 33292
rect 16640 32972 16652 33028
rect 16708 32972 16720 33028
rect 16640 32960 16720 32972
rect 16800 33348 16880 33360
rect 16800 33292 16812 33348
rect 16868 33292 16880 33348
rect 16800 33028 16880 33292
rect 16800 32972 16812 33028
rect 16868 32972 16880 33028
rect 16800 32960 16880 32972
rect 16960 33348 17040 33360
rect 16960 33292 16972 33348
rect 17028 33292 17040 33348
rect 16960 33028 17040 33292
rect 16960 32972 16972 33028
rect 17028 32972 17040 33028
rect 16960 32960 17040 32972
rect 17120 33348 17200 33360
rect 17120 33292 17132 33348
rect 17188 33292 17200 33348
rect 17120 33028 17200 33292
rect 17120 32972 17132 33028
rect 17188 32972 17200 33028
rect 17120 32960 17200 32972
rect 17280 33348 17360 33360
rect 17280 33292 17292 33348
rect 17348 33292 17360 33348
rect 17280 33028 17360 33292
rect 17280 32972 17292 33028
rect 17348 32972 17360 33028
rect 17280 32960 17360 32972
rect 17440 33348 17520 33360
rect 17440 33292 17452 33348
rect 17508 33292 17520 33348
rect 17440 33028 17520 33292
rect 17440 32972 17452 33028
rect 17508 32972 17520 33028
rect 17440 32960 17520 32972
rect 17600 33348 17680 33360
rect 17600 33292 17612 33348
rect 17668 33292 17680 33348
rect 17600 33028 17680 33292
rect 17600 32972 17612 33028
rect 17668 32972 17680 33028
rect 17600 32960 17680 32972
rect 17760 33348 17840 33360
rect 17760 33292 17772 33348
rect 17828 33292 17840 33348
rect 17760 33028 17840 33292
rect 17760 32972 17772 33028
rect 17828 32972 17840 33028
rect 17760 32960 17840 32972
rect 17920 33348 18000 33360
rect 17920 33292 17932 33348
rect 17988 33292 18000 33348
rect 17920 33028 18000 33292
rect 17920 32972 17932 33028
rect 17988 32972 18000 33028
rect 17920 32960 18000 32972
rect 18080 33348 18160 33360
rect 18080 33292 18092 33348
rect 18148 33292 18160 33348
rect 18080 33028 18160 33292
rect 18080 32972 18092 33028
rect 18148 32972 18160 33028
rect 18080 32960 18160 32972
rect 18240 33348 18320 33360
rect 18240 33292 18252 33348
rect 18308 33292 18320 33348
rect 18240 33028 18320 33292
rect 18240 32972 18252 33028
rect 18308 32972 18320 33028
rect 18240 32960 18320 32972
rect 18400 33348 18480 33360
rect 18400 33292 18412 33348
rect 18468 33292 18480 33348
rect 18400 33028 18480 33292
rect 18400 32972 18412 33028
rect 18468 32972 18480 33028
rect 18400 32960 18480 32972
rect 18560 33348 18640 33360
rect 18560 33292 18572 33348
rect 18628 33292 18640 33348
rect 18560 33028 18640 33292
rect 18560 32972 18572 33028
rect 18628 32972 18640 33028
rect 18560 32960 18640 32972
rect 18720 33348 18800 33360
rect 18720 33292 18732 33348
rect 18788 33292 18800 33348
rect 18720 33028 18800 33292
rect 18720 32972 18732 33028
rect 18788 32972 18800 33028
rect 18720 32960 18800 32972
rect 18880 33348 18960 33360
rect 18880 33292 18892 33348
rect 18948 33292 18960 33348
rect 18880 33028 18960 33292
rect 18880 32972 18892 33028
rect 18948 32972 18960 33028
rect 18880 32960 18960 32972
rect 19040 33348 19120 33452
rect 19040 33292 19052 33348
rect 19108 33292 19120 33348
rect 19040 33028 19120 33292
rect 19040 32972 19052 33028
rect 19108 32972 19120 33028
rect 12480 32868 12560 32880
rect 12480 32812 12492 32868
rect 12548 32812 12560 32868
rect 12480 32548 12560 32812
rect 12480 32492 12492 32548
rect 12548 32492 12560 32548
rect 12480 32480 12560 32492
rect 12640 32868 12720 32880
rect 12640 32812 12652 32868
rect 12708 32812 12720 32868
rect 12640 32548 12720 32812
rect 12640 32492 12652 32548
rect 12708 32492 12720 32548
rect 12640 32480 12720 32492
rect 12800 32868 12880 32880
rect 12800 32812 12812 32868
rect 12868 32812 12880 32868
rect 12800 32548 12880 32812
rect 12800 32492 12812 32548
rect 12868 32492 12880 32548
rect 12800 32480 12880 32492
rect 12960 32868 13040 32880
rect 12960 32812 12972 32868
rect 13028 32812 13040 32868
rect 12960 32548 13040 32812
rect 12960 32492 12972 32548
rect 13028 32492 13040 32548
rect 12960 32480 13040 32492
rect 13120 32868 13200 32880
rect 13120 32812 13132 32868
rect 13188 32812 13200 32868
rect 13120 32548 13200 32812
rect 13120 32492 13132 32548
rect 13188 32492 13200 32548
rect 13120 32480 13200 32492
rect 13280 32868 13360 32880
rect 13280 32812 13292 32868
rect 13348 32812 13360 32868
rect 13280 32548 13360 32812
rect 13280 32492 13292 32548
rect 13348 32492 13360 32548
rect 13280 32480 13360 32492
rect 13440 32868 13520 32880
rect 13440 32812 13452 32868
rect 13508 32812 13520 32868
rect 13440 32548 13520 32812
rect 13440 32492 13452 32548
rect 13508 32492 13520 32548
rect 13440 32480 13520 32492
rect 13600 32868 13680 32880
rect 13600 32812 13612 32868
rect 13668 32812 13680 32868
rect 13600 32548 13680 32812
rect 13600 32492 13612 32548
rect 13668 32492 13680 32548
rect 13600 32480 13680 32492
rect 13760 32868 13840 32880
rect 13760 32812 13772 32868
rect 13828 32812 13840 32868
rect 13760 32548 13840 32812
rect 13760 32492 13772 32548
rect 13828 32492 13840 32548
rect 13760 32480 13840 32492
rect 13920 32868 14000 32880
rect 13920 32812 13932 32868
rect 13988 32812 14000 32868
rect 13920 32548 14000 32812
rect 13920 32492 13932 32548
rect 13988 32492 14000 32548
rect 13920 32480 14000 32492
rect 14080 32868 14160 32880
rect 14080 32812 14092 32868
rect 14148 32812 14160 32868
rect 14080 32548 14160 32812
rect 14080 32492 14092 32548
rect 14148 32492 14160 32548
rect 14080 32480 14160 32492
rect 14240 32868 14320 32880
rect 14240 32812 14252 32868
rect 14308 32812 14320 32868
rect 14240 32548 14320 32812
rect 14240 32492 14252 32548
rect 14308 32492 14320 32548
rect 14240 32480 14320 32492
rect 14400 32868 14480 32880
rect 14400 32812 14412 32868
rect 14468 32812 14480 32868
rect 14400 32548 14480 32812
rect 14400 32492 14412 32548
rect 14468 32492 14480 32548
rect 14400 32480 14480 32492
rect 14560 32868 14640 32880
rect 14560 32812 14572 32868
rect 14628 32812 14640 32868
rect 14560 32548 14640 32812
rect 14560 32492 14572 32548
rect 14628 32492 14640 32548
rect 14560 32480 14640 32492
rect 14720 32868 14800 32880
rect 14720 32812 14732 32868
rect 14788 32812 14800 32868
rect 14720 32548 14800 32812
rect 14720 32492 14732 32548
rect 14788 32492 14800 32548
rect 14720 32480 14800 32492
rect 14880 32868 14960 32880
rect 14880 32812 14892 32868
rect 14948 32812 14960 32868
rect 14880 32548 14960 32812
rect 14880 32492 14892 32548
rect 14948 32492 14960 32548
rect 14880 32480 14960 32492
rect 15040 32868 15120 32880
rect 15040 32812 15052 32868
rect 15108 32812 15120 32868
rect 15040 32548 15120 32812
rect 15040 32492 15052 32548
rect 15108 32492 15120 32548
rect 15040 32480 15120 32492
rect 15200 32868 15280 32880
rect 15200 32812 15212 32868
rect 15268 32812 15280 32868
rect 15200 32548 15280 32812
rect 15200 32492 15212 32548
rect 15268 32492 15280 32548
rect 15200 32480 15280 32492
rect 15360 32868 15440 32880
rect 15360 32812 15372 32868
rect 15428 32812 15440 32868
rect 15360 32548 15440 32812
rect 15360 32492 15372 32548
rect 15428 32492 15440 32548
rect 15360 32480 15440 32492
rect 15520 32868 15600 32880
rect 15520 32812 15532 32868
rect 15588 32812 15600 32868
rect 15520 32548 15600 32812
rect 15520 32492 15532 32548
rect 15588 32492 15600 32548
rect 15520 32480 15600 32492
rect 15680 32868 15760 32880
rect 15680 32812 15692 32868
rect 15748 32812 15760 32868
rect 15680 32548 15760 32812
rect 15680 32492 15692 32548
rect 15748 32492 15760 32548
rect 15680 32480 15760 32492
rect 15840 32868 15920 32880
rect 15840 32812 15852 32868
rect 15908 32812 15920 32868
rect 15840 32548 15920 32812
rect 15840 32492 15852 32548
rect 15908 32492 15920 32548
rect 15840 32480 15920 32492
rect 16000 32868 16080 32880
rect 16000 32812 16012 32868
rect 16068 32812 16080 32868
rect 16000 32548 16080 32812
rect 16000 32492 16012 32548
rect 16068 32492 16080 32548
rect 16000 32480 16080 32492
rect 16160 32868 16240 32880
rect 16160 32812 16172 32868
rect 16228 32812 16240 32868
rect 16160 32548 16240 32812
rect 16160 32492 16172 32548
rect 16228 32492 16240 32548
rect 16160 32480 16240 32492
rect 16320 32868 16400 32880
rect 16320 32812 16332 32868
rect 16388 32812 16400 32868
rect 16320 32548 16400 32812
rect 16320 32492 16332 32548
rect 16388 32492 16400 32548
rect 16320 32480 16400 32492
rect 16480 32868 16560 32880
rect 16480 32812 16492 32868
rect 16548 32812 16560 32868
rect 16480 32548 16560 32812
rect 16480 32492 16492 32548
rect 16548 32492 16560 32548
rect 16480 32480 16560 32492
rect 16640 32868 16720 32880
rect 16640 32812 16652 32868
rect 16708 32812 16720 32868
rect 16640 32548 16720 32812
rect 16640 32492 16652 32548
rect 16708 32492 16720 32548
rect 16640 32480 16720 32492
rect 16800 32868 16880 32880
rect 16800 32812 16812 32868
rect 16868 32812 16880 32868
rect 16800 32548 16880 32812
rect 16800 32492 16812 32548
rect 16868 32492 16880 32548
rect 16800 32480 16880 32492
rect 16960 32868 17040 32880
rect 16960 32812 16972 32868
rect 17028 32812 17040 32868
rect 16960 32548 17040 32812
rect 16960 32492 16972 32548
rect 17028 32492 17040 32548
rect 16960 32480 17040 32492
rect 17120 32868 17200 32880
rect 17120 32812 17132 32868
rect 17188 32812 17200 32868
rect 17120 32548 17200 32812
rect 17120 32492 17132 32548
rect 17188 32492 17200 32548
rect 17120 32480 17200 32492
rect 17280 32868 17360 32880
rect 17280 32812 17292 32868
rect 17348 32812 17360 32868
rect 17280 32548 17360 32812
rect 17280 32492 17292 32548
rect 17348 32492 17360 32548
rect 17280 32480 17360 32492
rect 17440 32868 17520 32880
rect 17440 32812 17452 32868
rect 17508 32812 17520 32868
rect 17440 32548 17520 32812
rect 17440 32492 17452 32548
rect 17508 32492 17520 32548
rect 17440 32480 17520 32492
rect 17600 32868 17680 32880
rect 17600 32812 17612 32868
rect 17668 32812 17680 32868
rect 17600 32548 17680 32812
rect 17600 32492 17612 32548
rect 17668 32492 17680 32548
rect 17600 32480 17680 32492
rect 17760 32868 17840 32880
rect 17760 32812 17772 32868
rect 17828 32812 17840 32868
rect 17760 32548 17840 32812
rect 17760 32492 17772 32548
rect 17828 32492 17840 32548
rect 17760 32480 17840 32492
rect 17920 32868 18000 32880
rect 17920 32812 17932 32868
rect 17988 32812 18000 32868
rect 17920 32548 18000 32812
rect 17920 32492 17932 32548
rect 17988 32492 18000 32548
rect 17920 32480 18000 32492
rect 18080 32868 18160 32880
rect 18080 32812 18092 32868
rect 18148 32812 18160 32868
rect 18080 32548 18160 32812
rect 18080 32492 18092 32548
rect 18148 32492 18160 32548
rect 18080 32480 18160 32492
rect 18240 32868 18320 32880
rect 18240 32812 18252 32868
rect 18308 32812 18320 32868
rect 18240 32548 18320 32812
rect 18240 32492 18252 32548
rect 18308 32492 18320 32548
rect 18240 32480 18320 32492
rect 18400 32868 18480 32880
rect 18400 32812 18412 32868
rect 18468 32812 18480 32868
rect 18400 32548 18480 32812
rect 18400 32492 18412 32548
rect 18468 32492 18480 32548
rect 18400 32480 18480 32492
rect 18560 32868 18640 32880
rect 18560 32812 18572 32868
rect 18628 32812 18640 32868
rect 18560 32548 18640 32812
rect 18560 32492 18572 32548
rect 18628 32492 18640 32548
rect 18560 32480 18640 32492
rect 18720 32868 18800 32880
rect 18720 32812 18732 32868
rect 18788 32812 18800 32868
rect 18720 32548 18800 32812
rect 18720 32492 18732 32548
rect 18788 32492 18800 32548
rect 18720 32480 18800 32492
rect 18880 32868 18960 32880
rect 18880 32812 18892 32868
rect 18948 32812 18960 32868
rect 18880 32548 18960 32812
rect 18880 32492 18892 32548
rect 18948 32492 18960 32548
rect 18880 32480 18960 32492
rect 12480 32388 12560 32400
rect 12480 32332 12492 32388
rect 12548 32332 12560 32388
rect 12480 32068 12560 32332
rect 12480 32012 12492 32068
rect 12548 32012 12560 32068
rect 12480 31748 12560 32012
rect 12480 31692 12492 31748
rect 12548 31692 12560 31748
rect 12480 31428 12560 31692
rect 12480 31372 12492 31428
rect 12548 31372 12560 31428
rect 12480 31108 12560 31372
rect 12480 31052 12492 31108
rect 12548 31052 12560 31108
rect 12480 30788 12560 31052
rect 12480 30732 12492 30788
rect 12548 30732 12560 30788
rect 12480 30468 12560 30732
rect 12480 30412 12492 30468
rect 12548 30412 12560 30468
rect 12480 30400 12560 30412
rect 12640 32388 12720 32400
rect 12640 32332 12652 32388
rect 12708 32332 12720 32388
rect 12640 32068 12720 32332
rect 12640 32012 12652 32068
rect 12708 32012 12720 32068
rect 12640 31748 12720 32012
rect 12640 31692 12652 31748
rect 12708 31692 12720 31748
rect 12640 31428 12720 31692
rect 12640 31372 12652 31428
rect 12708 31372 12720 31428
rect 12640 31108 12720 31372
rect 12640 31052 12652 31108
rect 12708 31052 12720 31108
rect 12640 30788 12720 31052
rect 12640 30732 12652 30788
rect 12708 30732 12720 30788
rect 12640 30468 12720 30732
rect 12640 30412 12652 30468
rect 12708 30412 12720 30468
rect 12640 30400 12720 30412
rect 12800 32388 12880 32400
rect 12800 32332 12812 32388
rect 12868 32332 12880 32388
rect 12800 32068 12880 32332
rect 12800 32012 12812 32068
rect 12868 32012 12880 32068
rect 12800 31748 12880 32012
rect 12800 31692 12812 31748
rect 12868 31692 12880 31748
rect 12800 31428 12880 31692
rect 12800 31372 12812 31428
rect 12868 31372 12880 31428
rect 12800 31108 12880 31372
rect 12800 31052 12812 31108
rect 12868 31052 12880 31108
rect 12800 30788 12880 31052
rect 12800 30732 12812 30788
rect 12868 30732 12880 30788
rect 12800 30468 12880 30732
rect 12800 30412 12812 30468
rect 12868 30412 12880 30468
rect 12800 30400 12880 30412
rect 12960 32388 13040 32400
rect 12960 32332 12972 32388
rect 13028 32332 13040 32388
rect 12960 32068 13040 32332
rect 12960 32012 12972 32068
rect 13028 32012 13040 32068
rect 12960 31748 13040 32012
rect 12960 31692 12972 31748
rect 13028 31692 13040 31748
rect 12960 31428 13040 31692
rect 12960 31372 12972 31428
rect 13028 31372 13040 31428
rect 12960 31108 13040 31372
rect 12960 31052 12972 31108
rect 13028 31052 13040 31108
rect 12960 30788 13040 31052
rect 12960 30732 12972 30788
rect 13028 30732 13040 30788
rect 12960 30468 13040 30732
rect 12960 30412 12972 30468
rect 13028 30412 13040 30468
rect 12960 30400 13040 30412
rect 13120 32388 13200 32400
rect 13120 32332 13132 32388
rect 13188 32332 13200 32388
rect 13120 32068 13200 32332
rect 13120 32012 13132 32068
rect 13188 32012 13200 32068
rect 13120 31748 13200 32012
rect 13120 31692 13132 31748
rect 13188 31692 13200 31748
rect 13120 31428 13200 31692
rect 13120 31372 13132 31428
rect 13188 31372 13200 31428
rect 13120 31108 13200 31372
rect 13120 31052 13132 31108
rect 13188 31052 13200 31108
rect 13120 30788 13200 31052
rect 13120 30732 13132 30788
rect 13188 30732 13200 30788
rect 13120 30468 13200 30732
rect 13120 30412 13132 30468
rect 13188 30412 13200 30468
rect 13120 30400 13200 30412
rect 13280 32388 13360 32400
rect 13280 32332 13292 32388
rect 13348 32332 13360 32388
rect 13280 32068 13360 32332
rect 13280 32012 13292 32068
rect 13348 32012 13360 32068
rect 13280 31748 13360 32012
rect 13280 31692 13292 31748
rect 13348 31692 13360 31748
rect 13280 31428 13360 31692
rect 13280 31372 13292 31428
rect 13348 31372 13360 31428
rect 13280 31108 13360 31372
rect 13280 31052 13292 31108
rect 13348 31052 13360 31108
rect 13280 30788 13360 31052
rect 13280 30732 13292 30788
rect 13348 30732 13360 30788
rect 13280 30468 13360 30732
rect 13280 30412 13292 30468
rect 13348 30412 13360 30468
rect 13280 30400 13360 30412
rect 13440 32388 13520 32400
rect 13440 32332 13452 32388
rect 13508 32332 13520 32388
rect 13440 32068 13520 32332
rect 13440 32012 13452 32068
rect 13508 32012 13520 32068
rect 13440 31748 13520 32012
rect 13440 31692 13452 31748
rect 13508 31692 13520 31748
rect 13440 31428 13520 31692
rect 13440 31372 13452 31428
rect 13508 31372 13520 31428
rect 13440 31108 13520 31372
rect 13440 31052 13452 31108
rect 13508 31052 13520 31108
rect 13440 30788 13520 31052
rect 13440 30732 13452 30788
rect 13508 30732 13520 30788
rect 13440 30468 13520 30732
rect 13440 30412 13452 30468
rect 13508 30412 13520 30468
rect 13440 30400 13520 30412
rect 13600 32388 13680 32400
rect 13600 32332 13612 32388
rect 13668 32332 13680 32388
rect 13600 32068 13680 32332
rect 13600 32012 13612 32068
rect 13668 32012 13680 32068
rect 13600 31748 13680 32012
rect 13600 31692 13612 31748
rect 13668 31692 13680 31748
rect 13600 31428 13680 31692
rect 13600 31372 13612 31428
rect 13668 31372 13680 31428
rect 13600 31108 13680 31372
rect 13600 31052 13612 31108
rect 13668 31052 13680 31108
rect 13600 30788 13680 31052
rect 13600 30732 13612 30788
rect 13668 30732 13680 30788
rect 13600 30468 13680 30732
rect 13600 30412 13612 30468
rect 13668 30412 13680 30468
rect 13600 30400 13680 30412
rect 13760 32388 13840 32400
rect 13760 32332 13772 32388
rect 13828 32332 13840 32388
rect 13760 32068 13840 32332
rect 13760 32012 13772 32068
rect 13828 32012 13840 32068
rect 13760 31748 13840 32012
rect 13760 31692 13772 31748
rect 13828 31692 13840 31748
rect 13760 31428 13840 31692
rect 13760 31372 13772 31428
rect 13828 31372 13840 31428
rect 13760 31108 13840 31372
rect 13760 31052 13772 31108
rect 13828 31052 13840 31108
rect 13760 30788 13840 31052
rect 13760 30732 13772 30788
rect 13828 30732 13840 30788
rect 13760 30468 13840 30732
rect 13760 30412 13772 30468
rect 13828 30412 13840 30468
rect 13760 30400 13840 30412
rect 13920 32388 14000 32400
rect 13920 32332 13932 32388
rect 13988 32332 14000 32388
rect 13920 32068 14000 32332
rect 13920 32012 13932 32068
rect 13988 32012 14000 32068
rect 13920 31748 14000 32012
rect 13920 31692 13932 31748
rect 13988 31692 14000 31748
rect 13920 31428 14000 31692
rect 13920 31372 13932 31428
rect 13988 31372 14000 31428
rect 13920 31108 14000 31372
rect 13920 31052 13932 31108
rect 13988 31052 14000 31108
rect 13920 30788 14000 31052
rect 13920 30732 13932 30788
rect 13988 30732 14000 30788
rect 13920 30468 14000 30732
rect 13920 30412 13932 30468
rect 13988 30412 14000 30468
rect 13920 30400 14000 30412
rect 14080 32388 14160 32400
rect 14080 32332 14092 32388
rect 14148 32332 14160 32388
rect 14080 32068 14160 32332
rect 14080 32012 14092 32068
rect 14148 32012 14160 32068
rect 14080 31748 14160 32012
rect 14080 31692 14092 31748
rect 14148 31692 14160 31748
rect 14080 31428 14160 31692
rect 14080 31372 14092 31428
rect 14148 31372 14160 31428
rect 14080 31108 14160 31372
rect 14080 31052 14092 31108
rect 14148 31052 14160 31108
rect 14080 30788 14160 31052
rect 14080 30732 14092 30788
rect 14148 30732 14160 30788
rect 14080 30468 14160 30732
rect 14080 30412 14092 30468
rect 14148 30412 14160 30468
rect 14080 30400 14160 30412
rect 14240 32388 14320 32400
rect 14240 32332 14252 32388
rect 14308 32332 14320 32388
rect 14240 32068 14320 32332
rect 14240 32012 14252 32068
rect 14308 32012 14320 32068
rect 14240 31748 14320 32012
rect 14240 31692 14252 31748
rect 14308 31692 14320 31748
rect 14240 31428 14320 31692
rect 14240 31372 14252 31428
rect 14308 31372 14320 31428
rect 14240 31108 14320 31372
rect 14240 31052 14252 31108
rect 14308 31052 14320 31108
rect 14240 30788 14320 31052
rect 14240 30732 14252 30788
rect 14308 30732 14320 30788
rect 14240 30468 14320 30732
rect 14240 30412 14252 30468
rect 14308 30412 14320 30468
rect 14240 30400 14320 30412
rect 14400 32388 14480 32400
rect 14400 32332 14412 32388
rect 14468 32332 14480 32388
rect 14400 32068 14480 32332
rect 14400 32012 14412 32068
rect 14468 32012 14480 32068
rect 14400 31748 14480 32012
rect 14400 31692 14412 31748
rect 14468 31692 14480 31748
rect 14400 31428 14480 31692
rect 14400 31372 14412 31428
rect 14468 31372 14480 31428
rect 14400 31108 14480 31372
rect 14400 31052 14412 31108
rect 14468 31052 14480 31108
rect 14400 30788 14480 31052
rect 14400 30732 14412 30788
rect 14468 30732 14480 30788
rect 14400 30468 14480 30732
rect 14400 30412 14412 30468
rect 14468 30412 14480 30468
rect 14400 30400 14480 30412
rect 14560 32388 14640 32400
rect 14560 32332 14572 32388
rect 14628 32332 14640 32388
rect 14560 32068 14640 32332
rect 14560 32012 14572 32068
rect 14628 32012 14640 32068
rect 14560 31748 14640 32012
rect 14560 31692 14572 31748
rect 14628 31692 14640 31748
rect 14560 31428 14640 31692
rect 14560 31372 14572 31428
rect 14628 31372 14640 31428
rect 14560 31108 14640 31372
rect 14560 31052 14572 31108
rect 14628 31052 14640 31108
rect 14560 30788 14640 31052
rect 14560 30732 14572 30788
rect 14628 30732 14640 30788
rect 14560 30468 14640 30732
rect 14560 30412 14572 30468
rect 14628 30412 14640 30468
rect 14560 30400 14640 30412
rect 14720 32388 14800 32400
rect 14720 32332 14732 32388
rect 14788 32332 14800 32388
rect 14720 32068 14800 32332
rect 14720 32012 14732 32068
rect 14788 32012 14800 32068
rect 14720 31748 14800 32012
rect 14720 31692 14732 31748
rect 14788 31692 14800 31748
rect 14720 31428 14800 31692
rect 14720 31372 14732 31428
rect 14788 31372 14800 31428
rect 14720 31108 14800 31372
rect 14720 31052 14732 31108
rect 14788 31052 14800 31108
rect 14720 30788 14800 31052
rect 14720 30732 14732 30788
rect 14788 30732 14800 30788
rect 14720 30468 14800 30732
rect 14720 30412 14732 30468
rect 14788 30412 14800 30468
rect 14720 30400 14800 30412
rect 14880 32388 14960 32400
rect 14880 32332 14892 32388
rect 14948 32332 14960 32388
rect 14880 32068 14960 32332
rect 14880 32012 14892 32068
rect 14948 32012 14960 32068
rect 14880 31748 14960 32012
rect 14880 31692 14892 31748
rect 14948 31692 14960 31748
rect 14880 31428 14960 31692
rect 14880 31372 14892 31428
rect 14948 31372 14960 31428
rect 14880 31108 14960 31372
rect 14880 31052 14892 31108
rect 14948 31052 14960 31108
rect 14880 30788 14960 31052
rect 14880 30732 14892 30788
rect 14948 30732 14960 30788
rect 14880 30468 14960 30732
rect 14880 30412 14892 30468
rect 14948 30412 14960 30468
rect 14880 30400 14960 30412
rect 15040 32388 15120 32400
rect 15040 32332 15052 32388
rect 15108 32332 15120 32388
rect 15040 32068 15120 32332
rect 15040 32012 15052 32068
rect 15108 32012 15120 32068
rect 15040 31748 15120 32012
rect 15040 31692 15052 31748
rect 15108 31692 15120 31748
rect 15040 31428 15120 31692
rect 15040 31372 15052 31428
rect 15108 31372 15120 31428
rect 15040 31108 15120 31372
rect 15040 31052 15052 31108
rect 15108 31052 15120 31108
rect 15040 30788 15120 31052
rect 15040 30732 15052 30788
rect 15108 30732 15120 30788
rect 15040 30468 15120 30732
rect 15040 30412 15052 30468
rect 15108 30412 15120 30468
rect 15040 30400 15120 30412
rect 15200 32388 15280 32400
rect 15200 32332 15212 32388
rect 15268 32332 15280 32388
rect 15200 32068 15280 32332
rect 15200 32012 15212 32068
rect 15268 32012 15280 32068
rect 15200 31748 15280 32012
rect 15200 31692 15212 31748
rect 15268 31692 15280 31748
rect 15200 31428 15280 31692
rect 15200 31372 15212 31428
rect 15268 31372 15280 31428
rect 15200 31108 15280 31372
rect 15200 31052 15212 31108
rect 15268 31052 15280 31108
rect 15200 30788 15280 31052
rect 15200 30732 15212 30788
rect 15268 30732 15280 30788
rect 15200 30468 15280 30732
rect 15200 30412 15212 30468
rect 15268 30412 15280 30468
rect 15200 30400 15280 30412
rect 15360 32388 15440 32400
rect 15360 32332 15372 32388
rect 15428 32332 15440 32388
rect 15360 32068 15440 32332
rect 15360 32012 15372 32068
rect 15428 32012 15440 32068
rect 15360 31748 15440 32012
rect 15360 31692 15372 31748
rect 15428 31692 15440 31748
rect 15360 31428 15440 31692
rect 15360 31372 15372 31428
rect 15428 31372 15440 31428
rect 15360 31108 15440 31372
rect 15360 31052 15372 31108
rect 15428 31052 15440 31108
rect 15360 30788 15440 31052
rect 15360 30732 15372 30788
rect 15428 30732 15440 30788
rect 15360 30468 15440 30732
rect 15360 30412 15372 30468
rect 15428 30412 15440 30468
rect 15360 30400 15440 30412
rect 15520 32388 15600 32400
rect 15520 32332 15532 32388
rect 15588 32332 15600 32388
rect 15520 32068 15600 32332
rect 15520 32012 15532 32068
rect 15588 32012 15600 32068
rect 15520 31748 15600 32012
rect 15520 31692 15532 31748
rect 15588 31692 15600 31748
rect 15520 31428 15600 31692
rect 15520 31372 15532 31428
rect 15588 31372 15600 31428
rect 15520 31108 15600 31372
rect 15520 31052 15532 31108
rect 15588 31052 15600 31108
rect 15520 30788 15600 31052
rect 15520 30732 15532 30788
rect 15588 30732 15600 30788
rect 15520 30468 15600 30732
rect 15520 30412 15532 30468
rect 15588 30412 15600 30468
rect 15520 30400 15600 30412
rect 15680 32388 15760 32400
rect 15680 32332 15692 32388
rect 15748 32332 15760 32388
rect 15680 32068 15760 32332
rect 15680 32012 15692 32068
rect 15748 32012 15760 32068
rect 15680 31748 15760 32012
rect 15680 31692 15692 31748
rect 15748 31692 15760 31748
rect 15680 31428 15760 31692
rect 15680 31372 15692 31428
rect 15748 31372 15760 31428
rect 15680 31108 15760 31372
rect 15680 31052 15692 31108
rect 15748 31052 15760 31108
rect 15680 30788 15760 31052
rect 15680 30732 15692 30788
rect 15748 30732 15760 30788
rect 15680 30468 15760 30732
rect 15680 30412 15692 30468
rect 15748 30412 15760 30468
rect 15680 30400 15760 30412
rect 15840 32388 15920 32400
rect 15840 32332 15852 32388
rect 15908 32332 15920 32388
rect 15840 32068 15920 32332
rect 15840 32012 15852 32068
rect 15908 32012 15920 32068
rect 15840 31748 15920 32012
rect 15840 31692 15852 31748
rect 15908 31692 15920 31748
rect 15840 31428 15920 31692
rect 15840 31372 15852 31428
rect 15908 31372 15920 31428
rect 15840 31108 15920 31372
rect 15840 31052 15852 31108
rect 15908 31052 15920 31108
rect 15840 30788 15920 31052
rect 15840 30732 15852 30788
rect 15908 30732 15920 30788
rect 15840 30468 15920 30732
rect 15840 30412 15852 30468
rect 15908 30412 15920 30468
rect 15840 30400 15920 30412
rect 16000 32388 16080 32400
rect 16000 32332 16012 32388
rect 16068 32332 16080 32388
rect 16000 32068 16080 32332
rect 16000 32012 16012 32068
rect 16068 32012 16080 32068
rect 16000 31748 16080 32012
rect 16000 31692 16012 31748
rect 16068 31692 16080 31748
rect 16000 31428 16080 31692
rect 16000 31372 16012 31428
rect 16068 31372 16080 31428
rect 16000 31108 16080 31372
rect 16000 31052 16012 31108
rect 16068 31052 16080 31108
rect 16000 30788 16080 31052
rect 16000 30732 16012 30788
rect 16068 30732 16080 30788
rect 16000 30468 16080 30732
rect 16000 30412 16012 30468
rect 16068 30412 16080 30468
rect 16000 30400 16080 30412
rect 16160 32388 16240 32400
rect 16160 32332 16172 32388
rect 16228 32332 16240 32388
rect 16160 32068 16240 32332
rect 16160 32012 16172 32068
rect 16228 32012 16240 32068
rect 16160 31748 16240 32012
rect 16160 31692 16172 31748
rect 16228 31692 16240 31748
rect 16160 31428 16240 31692
rect 16160 31372 16172 31428
rect 16228 31372 16240 31428
rect 16160 31108 16240 31372
rect 16160 31052 16172 31108
rect 16228 31052 16240 31108
rect 16160 30788 16240 31052
rect 16160 30732 16172 30788
rect 16228 30732 16240 30788
rect 16160 30468 16240 30732
rect 16160 30412 16172 30468
rect 16228 30412 16240 30468
rect 16160 30400 16240 30412
rect 16320 32388 16400 32400
rect 16320 32332 16332 32388
rect 16388 32332 16400 32388
rect 16320 32068 16400 32332
rect 16320 32012 16332 32068
rect 16388 32012 16400 32068
rect 16320 31748 16400 32012
rect 16320 31692 16332 31748
rect 16388 31692 16400 31748
rect 16320 31428 16400 31692
rect 16320 31372 16332 31428
rect 16388 31372 16400 31428
rect 16320 31108 16400 31372
rect 16320 31052 16332 31108
rect 16388 31052 16400 31108
rect 16320 30788 16400 31052
rect 16320 30732 16332 30788
rect 16388 30732 16400 30788
rect 16320 30468 16400 30732
rect 16320 30412 16332 30468
rect 16388 30412 16400 30468
rect 16320 30400 16400 30412
rect 16480 32388 16560 32400
rect 16480 32332 16492 32388
rect 16548 32332 16560 32388
rect 16480 32068 16560 32332
rect 16480 32012 16492 32068
rect 16548 32012 16560 32068
rect 16480 31748 16560 32012
rect 16480 31692 16492 31748
rect 16548 31692 16560 31748
rect 16480 31428 16560 31692
rect 16480 31372 16492 31428
rect 16548 31372 16560 31428
rect 16480 31108 16560 31372
rect 16480 31052 16492 31108
rect 16548 31052 16560 31108
rect 16480 30788 16560 31052
rect 16480 30732 16492 30788
rect 16548 30732 16560 30788
rect 16480 30468 16560 30732
rect 16480 30412 16492 30468
rect 16548 30412 16560 30468
rect 16480 30400 16560 30412
rect 16640 32388 16720 32400
rect 16640 32332 16652 32388
rect 16708 32332 16720 32388
rect 16640 32068 16720 32332
rect 16640 32012 16652 32068
rect 16708 32012 16720 32068
rect 16640 31748 16720 32012
rect 16640 31692 16652 31748
rect 16708 31692 16720 31748
rect 16640 31428 16720 31692
rect 16640 31372 16652 31428
rect 16708 31372 16720 31428
rect 16640 31108 16720 31372
rect 16640 31052 16652 31108
rect 16708 31052 16720 31108
rect 16640 30788 16720 31052
rect 16640 30732 16652 30788
rect 16708 30732 16720 30788
rect 16640 30468 16720 30732
rect 16640 30412 16652 30468
rect 16708 30412 16720 30468
rect 16640 30400 16720 30412
rect 16800 32388 16880 32400
rect 16800 32332 16812 32388
rect 16868 32332 16880 32388
rect 16800 32068 16880 32332
rect 16800 32012 16812 32068
rect 16868 32012 16880 32068
rect 16800 31748 16880 32012
rect 16800 31692 16812 31748
rect 16868 31692 16880 31748
rect 16800 31428 16880 31692
rect 16800 31372 16812 31428
rect 16868 31372 16880 31428
rect 16800 31108 16880 31372
rect 16800 31052 16812 31108
rect 16868 31052 16880 31108
rect 16800 30788 16880 31052
rect 16800 30732 16812 30788
rect 16868 30732 16880 30788
rect 16800 30468 16880 30732
rect 16800 30412 16812 30468
rect 16868 30412 16880 30468
rect 16800 30400 16880 30412
rect 16960 32388 17040 32400
rect 16960 32332 16972 32388
rect 17028 32332 17040 32388
rect 16960 32068 17040 32332
rect 16960 32012 16972 32068
rect 17028 32012 17040 32068
rect 16960 31748 17040 32012
rect 16960 31692 16972 31748
rect 17028 31692 17040 31748
rect 16960 31428 17040 31692
rect 16960 31372 16972 31428
rect 17028 31372 17040 31428
rect 16960 31108 17040 31372
rect 16960 31052 16972 31108
rect 17028 31052 17040 31108
rect 16960 30788 17040 31052
rect 16960 30732 16972 30788
rect 17028 30732 17040 30788
rect 16960 30468 17040 30732
rect 16960 30412 16972 30468
rect 17028 30412 17040 30468
rect 16960 30400 17040 30412
rect 17120 32388 17200 32400
rect 17120 32332 17132 32388
rect 17188 32332 17200 32388
rect 17120 32068 17200 32332
rect 17120 32012 17132 32068
rect 17188 32012 17200 32068
rect 17120 31748 17200 32012
rect 17120 31692 17132 31748
rect 17188 31692 17200 31748
rect 17120 31428 17200 31692
rect 17120 31372 17132 31428
rect 17188 31372 17200 31428
rect 17120 31108 17200 31372
rect 17120 31052 17132 31108
rect 17188 31052 17200 31108
rect 17120 30788 17200 31052
rect 17120 30732 17132 30788
rect 17188 30732 17200 30788
rect 17120 30468 17200 30732
rect 17120 30412 17132 30468
rect 17188 30412 17200 30468
rect 17120 30400 17200 30412
rect 17280 32388 17360 32400
rect 17280 32332 17292 32388
rect 17348 32332 17360 32388
rect 17280 32068 17360 32332
rect 17280 32012 17292 32068
rect 17348 32012 17360 32068
rect 17280 31748 17360 32012
rect 17280 31692 17292 31748
rect 17348 31692 17360 31748
rect 17280 31428 17360 31692
rect 17280 31372 17292 31428
rect 17348 31372 17360 31428
rect 17280 31108 17360 31372
rect 17280 31052 17292 31108
rect 17348 31052 17360 31108
rect 17280 30788 17360 31052
rect 17280 30732 17292 30788
rect 17348 30732 17360 30788
rect 17280 30468 17360 30732
rect 17280 30412 17292 30468
rect 17348 30412 17360 30468
rect 17280 30400 17360 30412
rect 17440 32388 17520 32400
rect 17440 32332 17452 32388
rect 17508 32332 17520 32388
rect 17440 32068 17520 32332
rect 17440 32012 17452 32068
rect 17508 32012 17520 32068
rect 17440 31748 17520 32012
rect 17440 31692 17452 31748
rect 17508 31692 17520 31748
rect 17440 31428 17520 31692
rect 17440 31372 17452 31428
rect 17508 31372 17520 31428
rect 17440 31108 17520 31372
rect 17440 31052 17452 31108
rect 17508 31052 17520 31108
rect 17440 30788 17520 31052
rect 17440 30732 17452 30788
rect 17508 30732 17520 30788
rect 17440 30468 17520 30732
rect 17440 30412 17452 30468
rect 17508 30412 17520 30468
rect 17440 30400 17520 30412
rect 17600 32388 17680 32400
rect 17600 32332 17612 32388
rect 17668 32332 17680 32388
rect 17600 32068 17680 32332
rect 17600 32012 17612 32068
rect 17668 32012 17680 32068
rect 17600 31748 17680 32012
rect 17600 31692 17612 31748
rect 17668 31692 17680 31748
rect 17600 31428 17680 31692
rect 17600 31372 17612 31428
rect 17668 31372 17680 31428
rect 17600 31108 17680 31372
rect 17600 31052 17612 31108
rect 17668 31052 17680 31108
rect 17600 30788 17680 31052
rect 17600 30732 17612 30788
rect 17668 30732 17680 30788
rect 17600 30468 17680 30732
rect 17600 30412 17612 30468
rect 17668 30412 17680 30468
rect 17600 30400 17680 30412
rect 17760 32388 17840 32400
rect 17760 32332 17772 32388
rect 17828 32332 17840 32388
rect 17760 32068 17840 32332
rect 17760 32012 17772 32068
rect 17828 32012 17840 32068
rect 17760 31748 17840 32012
rect 17760 31692 17772 31748
rect 17828 31692 17840 31748
rect 17760 31428 17840 31692
rect 17760 31372 17772 31428
rect 17828 31372 17840 31428
rect 17760 31108 17840 31372
rect 17760 31052 17772 31108
rect 17828 31052 17840 31108
rect 17760 30788 17840 31052
rect 17760 30732 17772 30788
rect 17828 30732 17840 30788
rect 17760 30468 17840 30732
rect 17760 30412 17772 30468
rect 17828 30412 17840 30468
rect 17760 30400 17840 30412
rect 17920 32388 18000 32400
rect 17920 32332 17932 32388
rect 17988 32332 18000 32388
rect 17920 32068 18000 32332
rect 17920 32012 17932 32068
rect 17988 32012 18000 32068
rect 17920 31748 18000 32012
rect 17920 31692 17932 31748
rect 17988 31692 18000 31748
rect 17920 31428 18000 31692
rect 17920 31372 17932 31428
rect 17988 31372 18000 31428
rect 17920 31108 18000 31372
rect 17920 31052 17932 31108
rect 17988 31052 18000 31108
rect 17920 30788 18000 31052
rect 17920 30732 17932 30788
rect 17988 30732 18000 30788
rect 17920 30468 18000 30732
rect 17920 30412 17932 30468
rect 17988 30412 18000 30468
rect 17920 30400 18000 30412
rect 18080 32388 18160 32400
rect 18080 32332 18092 32388
rect 18148 32332 18160 32388
rect 18080 32068 18160 32332
rect 18080 32012 18092 32068
rect 18148 32012 18160 32068
rect 18080 31748 18160 32012
rect 18080 31692 18092 31748
rect 18148 31692 18160 31748
rect 18080 31428 18160 31692
rect 18080 31372 18092 31428
rect 18148 31372 18160 31428
rect 18080 31108 18160 31372
rect 18080 31052 18092 31108
rect 18148 31052 18160 31108
rect 18080 30788 18160 31052
rect 18080 30732 18092 30788
rect 18148 30732 18160 30788
rect 18080 30468 18160 30732
rect 18080 30412 18092 30468
rect 18148 30412 18160 30468
rect 18080 30400 18160 30412
rect 18240 32388 18320 32400
rect 18240 32332 18252 32388
rect 18308 32332 18320 32388
rect 18240 32068 18320 32332
rect 18240 32012 18252 32068
rect 18308 32012 18320 32068
rect 18240 31748 18320 32012
rect 18240 31692 18252 31748
rect 18308 31692 18320 31748
rect 18240 31428 18320 31692
rect 18240 31372 18252 31428
rect 18308 31372 18320 31428
rect 18240 31108 18320 31372
rect 18240 31052 18252 31108
rect 18308 31052 18320 31108
rect 18240 30788 18320 31052
rect 18240 30732 18252 30788
rect 18308 30732 18320 30788
rect 18240 30468 18320 30732
rect 18240 30412 18252 30468
rect 18308 30412 18320 30468
rect 18240 30400 18320 30412
rect 18400 32388 18480 32400
rect 18400 32332 18412 32388
rect 18468 32332 18480 32388
rect 18400 32068 18480 32332
rect 18400 32012 18412 32068
rect 18468 32012 18480 32068
rect 18400 31748 18480 32012
rect 18400 31692 18412 31748
rect 18468 31692 18480 31748
rect 18400 31428 18480 31692
rect 18400 31372 18412 31428
rect 18468 31372 18480 31428
rect 18400 31108 18480 31372
rect 18400 31052 18412 31108
rect 18468 31052 18480 31108
rect 18400 30788 18480 31052
rect 18400 30732 18412 30788
rect 18468 30732 18480 30788
rect 18400 30468 18480 30732
rect 18400 30412 18412 30468
rect 18468 30412 18480 30468
rect 18400 30400 18480 30412
rect 18560 32388 18640 32400
rect 18560 32332 18572 32388
rect 18628 32332 18640 32388
rect 18560 32068 18640 32332
rect 18560 32012 18572 32068
rect 18628 32012 18640 32068
rect 18560 31748 18640 32012
rect 18560 31692 18572 31748
rect 18628 31692 18640 31748
rect 18560 31428 18640 31692
rect 18560 31372 18572 31428
rect 18628 31372 18640 31428
rect 18560 31108 18640 31372
rect 18560 31052 18572 31108
rect 18628 31052 18640 31108
rect 18560 30788 18640 31052
rect 18560 30732 18572 30788
rect 18628 30732 18640 30788
rect 18560 30468 18640 30732
rect 18560 30412 18572 30468
rect 18628 30412 18640 30468
rect 18560 30400 18640 30412
rect 18720 32388 18800 32400
rect 18720 32332 18732 32388
rect 18788 32332 18800 32388
rect 18720 32068 18800 32332
rect 18720 32012 18732 32068
rect 18788 32012 18800 32068
rect 18720 31748 18800 32012
rect 18720 31692 18732 31748
rect 18788 31692 18800 31748
rect 18720 31428 18800 31692
rect 18720 31372 18732 31428
rect 18788 31372 18800 31428
rect 18720 31108 18800 31372
rect 18720 31052 18732 31108
rect 18788 31052 18800 31108
rect 18720 30788 18800 31052
rect 18720 30732 18732 30788
rect 18788 30732 18800 30788
rect 18720 30468 18800 30732
rect 18720 30412 18732 30468
rect 18788 30412 18800 30468
rect 18720 30400 18800 30412
rect 18880 32388 18960 32400
rect 18880 32332 18892 32388
rect 18948 32332 18960 32388
rect 18880 32068 18960 32332
rect 18880 32012 18892 32068
rect 18948 32012 18960 32068
rect 18880 31748 18960 32012
rect 18880 31692 18892 31748
rect 18948 31692 18960 31748
rect 18880 31428 18960 31692
rect 18880 31372 18892 31428
rect 18948 31372 18960 31428
rect 18880 31108 18960 31372
rect 18880 31052 18892 31108
rect 18948 31052 18960 31108
rect 18880 30788 18960 31052
rect 18880 30732 18892 30788
rect 18948 30732 18960 30788
rect 18880 30468 18960 30732
rect 18880 30412 18892 30468
rect 18948 30412 18960 30468
rect 18880 30400 18960 30412
rect 12480 30308 12560 30320
rect 12480 30252 12492 30308
rect 12548 30252 12560 30308
rect 12480 29988 12560 30252
rect 12480 29932 12492 29988
rect 12548 29932 12560 29988
rect 12480 29920 12560 29932
rect 12640 30308 12720 30320
rect 12640 30252 12652 30308
rect 12708 30252 12720 30308
rect 12640 29988 12720 30252
rect 12640 29932 12652 29988
rect 12708 29932 12720 29988
rect 12640 29920 12720 29932
rect 12800 30308 12880 30320
rect 12800 30252 12812 30308
rect 12868 30252 12880 30308
rect 12800 29988 12880 30252
rect 12800 29932 12812 29988
rect 12868 29932 12880 29988
rect 12800 29920 12880 29932
rect 12960 30308 13040 30320
rect 12960 30252 12972 30308
rect 13028 30252 13040 30308
rect 12960 29988 13040 30252
rect 12960 29932 12972 29988
rect 13028 29932 13040 29988
rect 12960 29920 13040 29932
rect 13120 30308 13200 30320
rect 13120 30252 13132 30308
rect 13188 30252 13200 30308
rect 13120 29988 13200 30252
rect 13120 29932 13132 29988
rect 13188 29932 13200 29988
rect 13120 29920 13200 29932
rect 13280 30308 13360 30320
rect 13280 30252 13292 30308
rect 13348 30252 13360 30308
rect 13280 29988 13360 30252
rect 13280 29932 13292 29988
rect 13348 29932 13360 29988
rect 13280 29920 13360 29932
rect 13440 30308 13520 30320
rect 13440 30252 13452 30308
rect 13508 30252 13520 30308
rect 13440 29988 13520 30252
rect 13440 29932 13452 29988
rect 13508 29932 13520 29988
rect 13440 29920 13520 29932
rect 13600 30308 13680 30320
rect 13600 30252 13612 30308
rect 13668 30252 13680 30308
rect 13600 29988 13680 30252
rect 13600 29932 13612 29988
rect 13668 29932 13680 29988
rect 13600 29920 13680 29932
rect 13760 30308 13840 30320
rect 13760 30252 13772 30308
rect 13828 30252 13840 30308
rect 13760 29988 13840 30252
rect 13760 29932 13772 29988
rect 13828 29932 13840 29988
rect 13760 29920 13840 29932
rect 13920 30308 14000 30320
rect 13920 30252 13932 30308
rect 13988 30252 14000 30308
rect 13920 29988 14000 30252
rect 13920 29932 13932 29988
rect 13988 29932 14000 29988
rect 13920 29920 14000 29932
rect 14080 30308 14160 30320
rect 14080 30252 14092 30308
rect 14148 30252 14160 30308
rect 14080 29988 14160 30252
rect 14080 29932 14092 29988
rect 14148 29932 14160 29988
rect 14080 29920 14160 29932
rect 14240 30308 14320 30320
rect 14240 30252 14252 30308
rect 14308 30252 14320 30308
rect 14240 29988 14320 30252
rect 14240 29932 14252 29988
rect 14308 29932 14320 29988
rect 14240 29920 14320 29932
rect 14400 30308 14480 30320
rect 14400 30252 14412 30308
rect 14468 30252 14480 30308
rect 14400 29988 14480 30252
rect 14400 29932 14412 29988
rect 14468 29932 14480 29988
rect 14400 29920 14480 29932
rect 14560 30308 14640 30320
rect 14560 30252 14572 30308
rect 14628 30252 14640 30308
rect 14560 29988 14640 30252
rect 14560 29932 14572 29988
rect 14628 29932 14640 29988
rect 14560 29920 14640 29932
rect 14720 30308 14800 30320
rect 14720 30252 14732 30308
rect 14788 30252 14800 30308
rect 14720 29988 14800 30252
rect 14720 29932 14732 29988
rect 14788 29932 14800 29988
rect 14720 29920 14800 29932
rect 14880 30308 14960 30320
rect 14880 30252 14892 30308
rect 14948 30252 14960 30308
rect 14880 29988 14960 30252
rect 14880 29932 14892 29988
rect 14948 29932 14960 29988
rect 14880 29920 14960 29932
rect 15040 30308 15120 30320
rect 15040 30252 15052 30308
rect 15108 30252 15120 30308
rect 15040 29988 15120 30252
rect 15040 29932 15052 29988
rect 15108 29932 15120 29988
rect 15040 29920 15120 29932
rect 15200 30308 15280 30320
rect 15200 30252 15212 30308
rect 15268 30252 15280 30308
rect 15200 29988 15280 30252
rect 15200 29932 15212 29988
rect 15268 29932 15280 29988
rect 15200 29920 15280 29932
rect 15360 30308 15440 30320
rect 15360 30252 15372 30308
rect 15428 30252 15440 30308
rect 15360 29988 15440 30252
rect 15360 29932 15372 29988
rect 15428 29932 15440 29988
rect 15360 29920 15440 29932
rect 15520 30308 15600 30320
rect 15520 30252 15532 30308
rect 15588 30252 15600 30308
rect 15520 29988 15600 30252
rect 15520 29932 15532 29988
rect 15588 29932 15600 29988
rect 15520 29920 15600 29932
rect 15680 30308 15760 30320
rect 15680 30252 15692 30308
rect 15748 30252 15760 30308
rect 15680 29988 15760 30252
rect 15680 29932 15692 29988
rect 15748 29932 15760 29988
rect 15680 29920 15760 29932
rect 15840 30308 15920 30320
rect 15840 30252 15852 30308
rect 15908 30252 15920 30308
rect 15840 29988 15920 30252
rect 15840 29932 15852 29988
rect 15908 29932 15920 29988
rect 15840 29920 15920 29932
rect 16000 30308 16080 30320
rect 16000 30252 16012 30308
rect 16068 30252 16080 30308
rect 16000 29988 16080 30252
rect 16000 29932 16012 29988
rect 16068 29932 16080 29988
rect 16000 29920 16080 29932
rect 16160 30308 16240 30320
rect 16160 30252 16172 30308
rect 16228 30252 16240 30308
rect 16160 29988 16240 30252
rect 16160 29932 16172 29988
rect 16228 29932 16240 29988
rect 16160 29920 16240 29932
rect 16320 30308 16400 30320
rect 16320 30252 16332 30308
rect 16388 30252 16400 30308
rect 16320 29988 16400 30252
rect 16320 29932 16332 29988
rect 16388 29932 16400 29988
rect 16320 29920 16400 29932
rect 16480 30308 16560 30320
rect 16480 30252 16492 30308
rect 16548 30252 16560 30308
rect 16480 29988 16560 30252
rect 16480 29932 16492 29988
rect 16548 29932 16560 29988
rect 16480 29920 16560 29932
rect 16640 30308 16720 30320
rect 16640 30252 16652 30308
rect 16708 30252 16720 30308
rect 16640 29988 16720 30252
rect 16640 29932 16652 29988
rect 16708 29932 16720 29988
rect 16640 29920 16720 29932
rect 16800 30308 16880 30320
rect 16800 30252 16812 30308
rect 16868 30252 16880 30308
rect 16800 29988 16880 30252
rect 16800 29932 16812 29988
rect 16868 29932 16880 29988
rect 16800 29920 16880 29932
rect 16960 30308 17040 30320
rect 16960 30252 16972 30308
rect 17028 30252 17040 30308
rect 16960 29988 17040 30252
rect 16960 29932 16972 29988
rect 17028 29932 17040 29988
rect 16960 29920 17040 29932
rect 17120 30308 17200 30320
rect 17120 30252 17132 30308
rect 17188 30252 17200 30308
rect 17120 29988 17200 30252
rect 17120 29932 17132 29988
rect 17188 29932 17200 29988
rect 17120 29920 17200 29932
rect 17280 30308 17360 30320
rect 17280 30252 17292 30308
rect 17348 30252 17360 30308
rect 17280 29988 17360 30252
rect 17280 29932 17292 29988
rect 17348 29932 17360 29988
rect 17280 29920 17360 29932
rect 17440 30308 17520 30320
rect 17440 30252 17452 30308
rect 17508 30252 17520 30308
rect 17440 29988 17520 30252
rect 17440 29932 17452 29988
rect 17508 29932 17520 29988
rect 17440 29920 17520 29932
rect 17600 30308 17680 30320
rect 17600 30252 17612 30308
rect 17668 30252 17680 30308
rect 17600 29988 17680 30252
rect 17600 29932 17612 29988
rect 17668 29932 17680 29988
rect 17600 29920 17680 29932
rect 17760 30308 17840 30320
rect 17760 30252 17772 30308
rect 17828 30252 17840 30308
rect 17760 29988 17840 30252
rect 17760 29932 17772 29988
rect 17828 29932 17840 29988
rect 17760 29920 17840 29932
rect 17920 30308 18000 30320
rect 17920 30252 17932 30308
rect 17988 30252 18000 30308
rect 17920 29988 18000 30252
rect 17920 29932 17932 29988
rect 17988 29932 18000 29988
rect 17920 29920 18000 29932
rect 18080 30308 18160 30320
rect 18080 30252 18092 30308
rect 18148 30252 18160 30308
rect 18080 29988 18160 30252
rect 18080 29932 18092 29988
rect 18148 29932 18160 29988
rect 18080 29920 18160 29932
rect 18240 30308 18320 30320
rect 18240 30252 18252 30308
rect 18308 30252 18320 30308
rect 18240 29988 18320 30252
rect 18240 29932 18252 29988
rect 18308 29932 18320 29988
rect 18240 29920 18320 29932
rect 18400 30308 18480 30320
rect 18400 30252 18412 30308
rect 18468 30252 18480 30308
rect 18400 29988 18480 30252
rect 18400 29932 18412 29988
rect 18468 29932 18480 29988
rect 18400 29920 18480 29932
rect 18560 30308 18640 30320
rect 18560 30252 18572 30308
rect 18628 30252 18640 30308
rect 18560 29988 18640 30252
rect 18560 29932 18572 29988
rect 18628 29932 18640 29988
rect 18560 29920 18640 29932
rect 18720 30308 18800 30320
rect 18720 30252 18732 30308
rect 18788 30252 18800 30308
rect 18720 29988 18800 30252
rect 18720 29932 18732 29988
rect 18788 29932 18800 29988
rect 18720 29920 18800 29932
rect 18880 30308 18960 30320
rect 18880 30252 18892 30308
rect 18948 30252 18960 30308
rect 18880 29988 18960 30252
rect 18880 29932 18892 29988
rect 18948 29932 18960 29988
rect 18880 29920 18960 29932
rect 12320 29772 12332 29828
rect 12388 29772 12400 29828
rect 12320 29508 12400 29772
rect 12320 29452 12332 29508
rect 12388 29452 12400 29508
rect 12320 29360 12400 29452
rect 12480 29828 12560 29840
rect 12480 29772 12492 29828
rect 12548 29772 12560 29828
rect 12480 29508 12560 29772
rect 12480 29452 12492 29508
rect 12548 29452 12560 29508
rect 12480 29440 12560 29452
rect 12640 29828 12720 29840
rect 12640 29772 12652 29828
rect 12708 29772 12720 29828
rect 12640 29508 12720 29772
rect 12640 29452 12652 29508
rect 12708 29452 12720 29508
rect 12640 29440 12720 29452
rect 12800 29828 12880 29840
rect 12800 29772 12812 29828
rect 12868 29772 12880 29828
rect 12800 29508 12880 29772
rect 12800 29452 12812 29508
rect 12868 29452 12880 29508
rect 12800 29440 12880 29452
rect 12960 29828 13040 29840
rect 12960 29772 12972 29828
rect 13028 29772 13040 29828
rect 12960 29508 13040 29772
rect 12960 29452 12972 29508
rect 13028 29452 13040 29508
rect 12960 29440 13040 29452
rect 13120 29828 13200 29840
rect 13120 29772 13132 29828
rect 13188 29772 13200 29828
rect 13120 29508 13200 29772
rect 13120 29452 13132 29508
rect 13188 29452 13200 29508
rect 13120 29440 13200 29452
rect 13280 29828 13360 29840
rect 13280 29772 13292 29828
rect 13348 29772 13360 29828
rect 13280 29508 13360 29772
rect 13280 29452 13292 29508
rect 13348 29452 13360 29508
rect 13280 29440 13360 29452
rect 13440 29828 13520 29840
rect 13440 29772 13452 29828
rect 13508 29772 13520 29828
rect 13440 29508 13520 29772
rect 13440 29452 13452 29508
rect 13508 29452 13520 29508
rect 13440 29440 13520 29452
rect 13600 29828 13680 29840
rect 13600 29772 13612 29828
rect 13668 29772 13680 29828
rect 13600 29508 13680 29772
rect 13600 29452 13612 29508
rect 13668 29452 13680 29508
rect 13600 29440 13680 29452
rect 13760 29828 13840 29840
rect 13760 29772 13772 29828
rect 13828 29772 13840 29828
rect 13760 29508 13840 29772
rect 13760 29452 13772 29508
rect 13828 29452 13840 29508
rect 13760 29440 13840 29452
rect 13920 29828 14000 29840
rect 13920 29772 13932 29828
rect 13988 29772 14000 29828
rect 13920 29508 14000 29772
rect 13920 29452 13932 29508
rect 13988 29452 14000 29508
rect 13920 29440 14000 29452
rect 14080 29828 14160 29840
rect 14080 29772 14092 29828
rect 14148 29772 14160 29828
rect 14080 29508 14160 29772
rect 14080 29452 14092 29508
rect 14148 29452 14160 29508
rect 14080 29440 14160 29452
rect 14240 29828 14320 29840
rect 14240 29772 14252 29828
rect 14308 29772 14320 29828
rect 14240 29508 14320 29772
rect 14240 29452 14252 29508
rect 14308 29452 14320 29508
rect 14240 29440 14320 29452
rect 14400 29828 14480 29840
rect 14400 29772 14412 29828
rect 14468 29772 14480 29828
rect 14400 29508 14480 29772
rect 14400 29452 14412 29508
rect 14468 29452 14480 29508
rect 14400 29440 14480 29452
rect 14560 29828 14640 29840
rect 14560 29772 14572 29828
rect 14628 29772 14640 29828
rect 14560 29508 14640 29772
rect 14560 29452 14572 29508
rect 14628 29452 14640 29508
rect 14560 29440 14640 29452
rect 14720 29828 14800 29840
rect 14720 29772 14732 29828
rect 14788 29772 14800 29828
rect 14720 29508 14800 29772
rect 14720 29452 14732 29508
rect 14788 29452 14800 29508
rect 14720 29440 14800 29452
rect 14880 29828 14960 29840
rect 14880 29772 14892 29828
rect 14948 29772 14960 29828
rect 14880 29508 14960 29772
rect 14880 29452 14892 29508
rect 14948 29452 14960 29508
rect 14880 29440 14960 29452
rect 15040 29828 15120 29840
rect 15040 29772 15052 29828
rect 15108 29772 15120 29828
rect 15040 29508 15120 29772
rect 15040 29452 15052 29508
rect 15108 29452 15120 29508
rect 15040 29440 15120 29452
rect 15200 29828 15280 29840
rect 15200 29772 15212 29828
rect 15268 29772 15280 29828
rect 15200 29508 15280 29772
rect 15200 29452 15212 29508
rect 15268 29452 15280 29508
rect 15200 29440 15280 29452
rect 15360 29828 15440 29840
rect 15360 29772 15372 29828
rect 15428 29772 15440 29828
rect 15360 29508 15440 29772
rect 15360 29452 15372 29508
rect 15428 29452 15440 29508
rect 15360 29440 15440 29452
rect 15520 29828 15600 29840
rect 15520 29772 15532 29828
rect 15588 29772 15600 29828
rect 15520 29508 15600 29772
rect 15520 29452 15532 29508
rect 15588 29452 15600 29508
rect 15520 29440 15600 29452
rect 15680 29828 15760 29840
rect 15680 29772 15692 29828
rect 15748 29772 15760 29828
rect 15680 29508 15760 29772
rect 15680 29452 15692 29508
rect 15748 29452 15760 29508
rect 15680 29440 15760 29452
rect 15840 29828 15920 29840
rect 15840 29772 15852 29828
rect 15908 29772 15920 29828
rect 15840 29508 15920 29772
rect 15840 29452 15852 29508
rect 15908 29452 15920 29508
rect 15840 29440 15920 29452
rect 16000 29828 16080 29840
rect 16000 29772 16012 29828
rect 16068 29772 16080 29828
rect 16000 29508 16080 29772
rect 16000 29452 16012 29508
rect 16068 29452 16080 29508
rect 16000 29440 16080 29452
rect 16160 29828 16240 29840
rect 16160 29772 16172 29828
rect 16228 29772 16240 29828
rect 16160 29508 16240 29772
rect 16160 29452 16172 29508
rect 16228 29452 16240 29508
rect 16160 29440 16240 29452
rect 16320 29828 16400 29840
rect 16320 29772 16332 29828
rect 16388 29772 16400 29828
rect 16320 29508 16400 29772
rect 16320 29452 16332 29508
rect 16388 29452 16400 29508
rect 16320 29440 16400 29452
rect 16480 29828 16560 29840
rect 16480 29772 16492 29828
rect 16548 29772 16560 29828
rect 16480 29508 16560 29772
rect 16480 29452 16492 29508
rect 16548 29452 16560 29508
rect 16480 29440 16560 29452
rect 16640 29828 16720 29840
rect 16640 29772 16652 29828
rect 16708 29772 16720 29828
rect 16640 29508 16720 29772
rect 16640 29452 16652 29508
rect 16708 29452 16720 29508
rect 16640 29440 16720 29452
rect 16800 29828 16880 29840
rect 16800 29772 16812 29828
rect 16868 29772 16880 29828
rect 16800 29508 16880 29772
rect 16800 29452 16812 29508
rect 16868 29452 16880 29508
rect 16800 29440 16880 29452
rect 16960 29828 17040 29840
rect 16960 29772 16972 29828
rect 17028 29772 17040 29828
rect 16960 29508 17040 29772
rect 16960 29452 16972 29508
rect 17028 29452 17040 29508
rect 16960 29440 17040 29452
rect 17120 29828 17200 29840
rect 17120 29772 17132 29828
rect 17188 29772 17200 29828
rect 17120 29508 17200 29772
rect 17120 29452 17132 29508
rect 17188 29452 17200 29508
rect 17120 29440 17200 29452
rect 17280 29828 17360 29840
rect 17280 29772 17292 29828
rect 17348 29772 17360 29828
rect 17280 29508 17360 29772
rect 17280 29452 17292 29508
rect 17348 29452 17360 29508
rect 17280 29440 17360 29452
rect 17440 29828 17520 29840
rect 17440 29772 17452 29828
rect 17508 29772 17520 29828
rect 17440 29508 17520 29772
rect 17440 29452 17452 29508
rect 17508 29452 17520 29508
rect 17440 29440 17520 29452
rect 17600 29828 17680 29840
rect 17600 29772 17612 29828
rect 17668 29772 17680 29828
rect 17600 29508 17680 29772
rect 17600 29452 17612 29508
rect 17668 29452 17680 29508
rect 17600 29440 17680 29452
rect 17760 29828 17840 29840
rect 17760 29772 17772 29828
rect 17828 29772 17840 29828
rect 17760 29508 17840 29772
rect 17760 29452 17772 29508
rect 17828 29452 17840 29508
rect 17760 29440 17840 29452
rect 17920 29828 18000 29840
rect 17920 29772 17932 29828
rect 17988 29772 18000 29828
rect 17920 29508 18000 29772
rect 17920 29452 17932 29508
rect 17988 29452 18000 29508
rect 17920 29440 18000 29452
rect 18080 29828 18160 29840
rect 18080 29772 18092 29828
rect 18148 29772 18160 29828
rect 18080 29508 18160 29772
rect 18080 29452 18092 29508
rect 18148 29452 18160 29508
rect 18080 29440 18160 29452
rect 18240 29828 18320 29840
rect 18240 29772 18252 29828
rect 18308 29772 18320 29828
rect 18240 29508 18320 29772
rect 18240 29452 18252 29508
rect 18308 29452 18320 29508
rect 18240 29440 18320 29452
rect 18400 29828 18480 29840
rect 18400 29772 18412 29828
rect 18468 29772 18480 29828
rect 18400 29508 18480 29772
rect 18400 29452 18412 29508
rect 18468 29452 18480 29508
rect 18400 29440 18480 29452
rect 18560 29828 18640 29840
rect 18560 29772 18572 29828
rect 18628 29772 18640 29828
rect 18560 29508 18640 29772
rect 18560 29452 18572 29508
rect 18628 29452 18640 29508
rect 18560 29440 18640 29452
rect 18720 29828 18800 29840
rect 18720 29772 18732 29828
rect 18788 29772 18800 29828
rect 18720 29508 18800 29772
rect 18720 29452 18732 29508
rect 18788 29452 18800 29508
rect 18720 29440 18800 29452
rect 18880 29828 18960 29840
rect 18880 29772 18892 29828
rect 18948 29772 18960 29828
rect 18880 29508 18960 29772
rect 18880 29452 18892 29508
rect 18948 29452 18960 29508
rect 18880 29440 18960 29452
rect 19040 29440 19120 32972
rect 19200 33668 19280 37360
rect 19200 33612 19212 33668
rect 19268 33612 19280 33668
rect 19200 33188 19280 33612
rect 19200 33132 19212 33188
rect 19268 33132 19280 33188
rect 19200 29440 19280 33132
rect 19360 33828 19440 37360
rect 19360 33772 19372 33828
rect 19428 33772 19440 33828
rect 19360 33508 19440 33772
rect 19360 33452 19372 33508
rect 19428 33452 19440 33508
rect 19360 33348 19440 33452
rect 19360 33292 19372 33348
rect 19428 33292 19440 33348
rect 19360 33028 19440 33292
rect 19360 32972 19372 33028
rect 19428 32972 19440 33028
rect 19360 29440 19440 32972
rect 19520 34308 19600 37360
rect 19520 34252 19532 34308
rect 19588 34252 19600 34308
rect 19520 33988 19600 34252
rect 19520 33932 19532 33988
rect 19588 33932 19600 33988
rect 19520 32868 19600 33932
rect 19520 32812 19532 32868
rect 19588 32812 19600 32868
rect 19520 32548 19600 32812
rect 19520 32492 19532 32548
rect 19588 32492 19600 32548
rect 19520 29440 19600 32492
rect 19680 34148 19760 37360
rect 19680 34092 19692 34148
rect 19748 34092 19760 34148
rect 19680 32708 19760 34092
rect 19680 32652 19692 32708
rect 19748 32652 19760 32708
rect 19680 29440 19760 32652
rect 19840 34308 19920 37360
rect 19840 34252 19852 34308
rect 19908 34252 19920 34308
rect 19840 33988 19920 34252
rect 19840 33932 19852 33988
rect 19908 33932 19920 33988
rect 19840 32868 19920 33932
rect 19840 32812 19852 32868
rect 19908 32812 19920 32868
rect 19840 32548 19920 32812
rect 19840 32492 19852 32548
rect 19908 32492 19920 32548
rect 19840 29440 19920 32492
rect 20000 36388 20080 37360
rect 20000 36332 20012 36388
rect 20068 36332 20080 36388
rect 20000 36068 20080 36332
rect 20000 36012 20012 36068
rect 20068 36012 20080 36068
rect 20000 35748 20080 36012
rect 20000 35692 20012 35748
rect 20068 35692 20080 35748
rect 20000 35428 20080 35692
rect 20000 35372 20012 35428
rect 20068 35372 20080 35428
rect 20000 35108 20080 35372
rect 20000 35052 20012 35108
rect 20068 35052 20080 35108
rect 20000 34788 20080 35052
rect 20000 34732 20012 34788
rect 20068 34732 20080 34788
rect 20000 34468 20080 34732
rect 20000 34412 20012 34468
rect 20068 34412 20080 34468
rect 20000 32388 20080 34412
rect 20000 32332 20012 32388
rect 20068 32332 20080 32388
rect 20000 32068 20080 32332
rect 20000 32012 20012 32068
rect 20068 32012 20080 32068
rect 20000 31748 20080 32012
rect 20000 31692 20012 31748
rect 20068 31692 20080 31748
rect 20000 31428 20080 31692
rect 20000 31372 20012 31428
rect 20068 31372 20080 31428
rect 20000 31108 20080 31372
rect 20000 31052 20012 31108
rect 20068 31052 20080 31108
rect 20000 30788 20080 31052
rect 20000 30732 20012 30788
rect 20068 30732 20080 30788
rect 20000 30468 20080 30732
rect 20000 30412 20012 30468
rect 20068 30412 20080 30468
rect 20000 29440 20080 30412
rect 20160 34628 20240 37360
rect 20160 34572 20172 34628
rect 20228 34572 20240 34628
rect 20160 32228 20240 34572
rect 20160 32172 20172 32228
rect 20228 32172 20240 32228
rect 20160 29440 20240 32172
rect 20320 36388 20400 37360
rect 20320 36332 20332 36388
rect 20388 36332 20400 36388
rect 20320 36068 20400 36332
rect 20320 36012 20332 36068
rect 20388 36012 20400 36068
rect 20320 35748 20400 36012
rect 20320 35692 20332 35748
rect 20388 35692 20400 35748
rect 20320 35428 20400 35692
rect 20320 35372 20332 35428
rect 20388 35372 20400 35428
rect 20320 35108 20400 35372
rect 20320 35052 20332 35108
rect 20388 35052 20400 35108
rect 20320 34788 20400 35052
rect 20320 34732 20332 34788
rect 20388 34732 20400 34788
rect 20320 34468 20400 34732
rect 20320 34412 20332 34468
rect 20388 34412 20400 34468
rect 20320 32388 20400 34412
rect 20320 32332 20332 32388
rect 20388 32332 20400 32388
rect 20320 32068 20400 32332
rect 20320 32012 20332 32068
rect 20388 32012 20400 32068
rect 20320 31748 20400 32012
rect 20320 31692 20332 31748
rect 20388 31692 20400 31748
rect 20320 31428 20400 31692
rect 20320 31372 20332 31428
rect 20388 31372 20400 31428
rect 20320 31108 20400 31372
rect 20320 31052 20332 31108
rect 20388 31052 20400 31108
rect 20320 30788 20400 31052
rect 20320 30732 20332 30788
rect 20388 30732 20400 30788
rect 20320 30468 20400 30732
rect 20320 30412 20332 30468
rect 20388 30412 20400 30468
rect 20320 29440 20400 30412
rect 20480 34948 20560 37360
rect 20480 34892 20492 34948
rect 20548 34892 20560 34948
rect 20480 31908 20560 34892
rect 20480 31852 20492 31908
rect 20548 31852 20560 31908
rect 20480 29440 20560 31852
rect 20640 36388 20720 37360
rect 20640 36332 20652 36388
rect 20708 36332 20720 36388
rect 20640 36068 20720 36332
rect 20640 36012 20652 36068
rect 20708 36012 20720 36068
rect 20640 35748 20720 36012
rect 20640 35692 20652 35748
rect 20708 35692 20720 35748
rect 20640 35428 20720 35692
rect 20640 35372 20652 35428
rect 20708 35372 20720 35428
rect 20640 35108 20720 35372
rect 20640 35052 20652 35108
rect 20708 35052 20720 35108
rect 20640 34788 20720 35052
rect 20640 34732 20652 34788
rect 20708 34732 20720 34788
rect 20640 34468 20720 34732
rect 20640 34412 20652 34468
rect 20708 34412 20720 34468
rect 20640 32388 20720 34412
rect 20640 32332 20652 32388
rect 20708 32332 20720 32388
rect 20640 32068 20720 32332
rect 20640 32012 20652 32068
rect 20708 32012 20720 32068
rect 20640 31748 20720 32012
rect 20640 31692 20652 31748
rect 20708 31692 20720 31748
rect 20640 31428 20720 31692
rect 20640 31372 20652 31428
rect 20708 31372 20720 31428
rect 20640 31108 20720 31372
rect 20640 31052 20652 31108
rect 20708 31052 20720 31108
rect 20640 30788 20720 31052
rect 20640 30732 20652 30788
rect 20708 30732 20720 30788
rect 20640 30468 20720 30732
rect 20640 30412 20652 30468
rect 20708 30412 20720 30468
rect 20640 29440 20720 30412
rect 20800 35268 20880 37360
rect 20800 35212 20812 35268
rect 20868 35212 20880 35268
rect 20800 31588 20880 35212
rect 20800 31532 20812 31588
rect 20868 31532 20880 31588
rect 20800 29440 20880 31532
rect 20960 36388 21040 37360
rect 20960 36332 20972 36388
rect 21028 36332 21040 36388
rect 20960 36068 21040 36332
rect 20960 36012 20972 36068
rect 21028 36012 21040 36068
rect 20960 35748 21040 36012
rect 20960 35692 20972 35748
rect 21028 35692 21040 35748
rect 20960 35428 21040 35692
rect 20960 35372 20972 35428
rect 21028 35372 21040 35428
rect 20960 35108 21040 35372
rect 20960 35052 20972 35108
rect 21028 35052 21040 35108
rect 20960 34788 21040 35052
rect 20960 34732 20972 34788
rect 21028 34732 21040 34788
rect 20960 34468 21040 34732
rect 20960 34412 20972 34468
rect 21028 34412 21040 34468
rect 20960 32388 21040 34412
rect 20960 32332 20972 32388
rect 21028 32332 21040 32388
rect 20960 32068 21040 32332
rect 20960 32012 20972 32068
rect 21028 32012 21040 32068
rect 20960 31748 21040 32012
rect 20960 31692 20972 31748
rect 21028 31692 21040 31748
rect 20960 31428 21040 31692
rect 20960 31372 20972 31428
rect 21028 31372 21040 31428
rect 20960 31108 21040 31372
rect 20960 31052 20972 31108
rect 21028 31052 21040 31108
rect 20960 30788 21040 31052
rect 20960 30732 20972 30788
rect 21028 30732 21040 30788
rect 20960 30468 21040 30732
rect 20960 30412 20972 30468
rect 21028 30412 21040 30468
rect 20960 29440 21040 30412
rect 21120 35588 21200 37360
rect 21120 35532 21132 35588
rect 21188 35532 21200 35588
rect 21120 31268 21200 35532
rect 21120 31212 21132 31268
rect 21188 31212 21200 31268
rect 21120 29440 21200 31212
rect 21280 36388 21360 37360
rect 21280 36332 21292 36388
rect 21348 36332 21360 36388
rect 21280 36068 21360 36332
rect 21280 36012 21292 36068
rect 21348 36012 21360 36068
rect 21280 35748 21360 36012
rect 21280 35692 21292 35748
rect 21348 35692 21360 35748
rect 21280 35428 21360 35692
rect 21280 35372 21292 35428
rect 21348 35372 21360 35428
rect 21280 35108 21360 35372
rect 21280 35052 21292 35108
rect 21348 35052 21360 35108
rect 21280 34788 21360 35052
rect 21280 34732 21292 34788
rect 21348 34732 21360 34788
rect 21280 34468 21360 34732
rect 21280 34412 21292 34468
rect 21348 34412 21360 34468
rect 21280 32388 21360 34412
rect 21280 32332 21292 32388
rect 21348 32332 21360 32388
rect 21280 32068 21360 32332
rect 21280 32012 21292 32068
rect 21348 32012 21360 32068
rect 21280 31748 21360 32012
rect 21280 31692 21292 31748
rect 21348 31692 21360 31748
rect 21280 31428 21360 31692
rect 21280 31372 21292 31428
rect 21348 31372 21360 31428
rect 21280 31108 21360 31372
rect 21280 31052 21292 31108
rect 21348 31052 21360 31108
rect 21280 30788 21360 31052
rect 21280 30732 21292 30788
rect 21348 30732 21360 30788
rect 21280 30468 21360 30732
rect 21280 30412 21292 30468
rect 21348 30412 21360 30468
rect 21280 29440 21360 30412
rect 21440 35908 21520 37360
rect 21440 35852 21452 35908
rect 21508 35852 21520 35908
rect 21440 30948 21520 35852
rect 21440 30892 21452 30948
rect 21508 30892 21520 30948
rect 21440 29440 21520 30892
rect 21600 36388 21680 37360
rect 21600 36332 21612 36388
rect 21668 36332 21680 36388
rect 21600 36068 21680 36332
rect 21600 36012 21612 36068
rect 21668 36012 21680 36068
rect 21600 35748 21680 36012
rect 21600 35692 21612 35748
rect 21668 35692 21680 35748
rect 21600 35428 21680 35692
rect 21600 35372 21612 35428
rect 21668 35372 21680 35428
rect 21600 35108 21680 35372
rect 21600 35052 21612 35108
rect 21668 35052 21680 35108
rect 21600 34788 21680 35052
rect 21600 34732 21612 34788
rect 21668 34732 21680 34788
rect 21600 34468 21680 34732
rect 21600 34412 21612 34468
rect 21668 34412 21680 34468
rect 21600 32388 21680 34412
rect 21600 32332 21612 32388
rect 21668 32332 21680 32388
rect 21600 32068 21680 32332
rect 21600 32012 21612 32068
rect 21668 32012 21680 32068
rect 21600 31748 21680 32012
rect 21600 31692 21612 31748
rect 21668 31692 21680 31748
rect 21600 31428 21680 31692
rect 21600 31372 21612 31428
rect 21668 31372 21680 31428
rect 21600 31108 21680 31372
rect 21600 31052 21612 31108
rect 21668 31052 21680 31108
rect 21600 30788 21680 31052
rect 21600 30732 21612 30788
rect 21668 30732 21680 30788
rect 21600 30468 21680 30732
rect 21600 30412 21612 30468
rect 21668 30412 21680 30468
rect 21600 29440 21680 30412
rect 21760 36228 21840 37360
rect 21760 36172 21772 36228
rect 21828 36172 21840 36228
rect 21760 30628 21840 36172
rect 21760 30572 21772 30628
rect 21828 30572 21840 30628
rect 21760 29440 21840 30572
rect 21920 36388 22000 37360
rect 21920 36332 21932 36388
rect 21988 36332 22000 36388
rect 21920 36068 22000 36332
rect 21920 36012 21932 36068
rect 21988 36012 22000 36068
rect 21920 35748 22000 36012
rect 21920 35692 21932 35748
rect 21988 35692 22000 35748
rect 21920 35428 22000 35692
rect 21920 35372 21932 35428
rect 21988 35372 22000 35428
rect 21920 35108 22000 35372
rect 21920 35052 21932 35108
rect 21988 35052 22000 35108
rect 21920 34788 22000 35052
rect 21920 34732 21932 34788
rect 21988 34732 22000 34788
rect 21920 34468 22000 34732
rect 21920 34412 21932 34468
rect 21988 34412 22000 34468
rect 21920 32388 22000 34412
rect 21920 32332 21932 32388
rect 21988 32332 22000 32388
rect 21920 32068 22000 32332
rect 21920 32012 21932 32068
rect 21988 32012 22000 32068
rect 21920 31748 22000 32012
rect 21920 31692 21932 31748
rect 21988 31692 22000 31748
rect 21920 31428 22000 31692
rect 21920 31372 21932 31428
rect 21988 31372 22000 31428
rect 21920 31108 22000 31372
rect 21920 31052 21932 31108
rect 21988 31052 22000 31108
rect 21920 30788 22000 31052
rect 21920 30732 21932 30788
rect 21988 30732 22000 30788
rect 21920 30468 22000 30732
rect 21920 30412 21932 30468
rect 21988 30412 22000 30468
rect 21920 29440 22000 30412
rect 22080 36868 22160 37360
rect 22080 36812 22092 36868
rect 22148 36812 22160 36868
rect 22080 36548 22160 36812
rect 22080 36492 22092 36548
rect 22148 36492 22160 36548
rect 22080 30308 22160 36492
rect 22080 30252 22092 30308
rect 22148 30252 22160 30308
rect 22080 29988 22160 30252
rect 22080 29932 22092 29988
rect 22148 29932 22160 29988
rect 22080 29440 22160 29932
rect 22240 36708 22320 37360
rect 22240 36652 22252 36708
rect 22308 36652 22320 36708
rect 22240 30148 22320 36652
rect 22240 30092 22252 30148
rect 22308 30092 22320 30148
rect 22240 29440 22320 30092
rect 22400 36868 22480 37360
rect 22400 36812 22412 36868
rect 22468 36812 22480 36868
rect 22400 36548 22480 36812
rect 22400 36492 22412 36548
rect 22468 36492 22480 36548
rect 22400 30308 22480 36492
rect 22400 30252 22412 30308
rect 22468 30252 22480 30308
rect 22400 29988 22480 30252
rect 22400 29932 22412 29988
rect 22468 29932 22480 29988
rect 22400 29440 22480 29932
rect 22560 37348 22640 37360
rect 22560 37292 22572 37348
rect 22628 37292 22640 37348
rect 22560 37028 22640 37292
rect 22560 36972 22572 37028
rect 22628 36972 22640 37028
rect 22560 29828 22640 36972
rect 22560 29772 22572 29828
rect 22628 29772 22640 29828
rect 22560 29508 22640 29772
rect 22560 29452 22572 29508
rect 22628 29452 22640 29508
rect 22560 29440 22640 29452
rect 22720 37188 22800 37360
rect 22720 37132 22732 37188
rect 22788 37132 22800 37188
rect 22720 29668 22800 37132
rect 22720 29612 22732 29668
rect 22788 29612 22800 29668
rect 22720 29440 22800 29612
rect 22880 37348 22960 37360
rect 22880 37292 22892 37348
rect 22948 37292 22960 37348
rect 22880 37028 22960 37292
rect 22880 36972 22892 37028
rect 22948 36972 22960 37028
rect 22880 29828 22960 36972
rect 23120 37348 23200 37360
rect 23120 37292 23132 37348
rect 23188 37292 23200 37348
rect 23120 37028 23200 37292
rect 23120 36972 23132 37028
rect 23188 36972 23200 37028
rect 23120 36960 23200 36972
rect 23280 37348 23360 37360
rect 23280 37292 23292 37348
rect 23348 37292 23360 37348
rect 23280 37028 23360 37292
rect 23280 36972 23292 37028
rect 23348 36972 23360 37028
rect 23280 36960 23360 36972
rect 23440 37348 23520 37360
rect 23440 37292 23452 37348
rect 23508 37292 23520 37348
rect 23440 37028 23520 37292
rect 23440 36972 23452 37028
rect 23508 36972 23520 37028
rect 23440 36960 23520 36972
rect 23600 37348 23680 37360
rect 23600 37292 23612 37348
rect 23668 37292 23680 37348
rect 23600 37028 23680 37292
rect 23600 36972 23612 37028
rect 23668 36972 23680 37028
rect 23600 36960 23680 36972
rect 23760 37348 23840 37360
rect 23760 37292 23772 37348
rect 23828 37292 23840 37348
rect 23760 37028 23840 37292
rect 23760 36972 23772 37028
rect 23828 36972 23840 37028
rect 23760 36960 23840 36972
rect 23920 37348 24000 37360
rect 23920 37292 23932 37348
rect 23988 37292 24000 37348
rect 23920 37028 24000 37292
rect 23920 36972 23932 37028
rect 23988 36972 24000 37028
rect 23920 36960 24000 36972
rect 24080 37348 24160 37360
rect 24080 37292 24092 37348
rect 24148 37292 24160 37348
rect 24080 37028 24160 37292
rect 24080 36972 24092 37028
rect 24148 36972 24160 37028
rect 24080 36960 24160 36972
rect 24240 37348 24320 37360
rect 24240 37292 24252 37348
rect 24308 37292 24320 37348
rect 24240 37028 24320 37292
rect 24240 36972 24252 37028
rect 24308 36972 24320 37028
rect 24240 36960 24320 36972
rect 24400 37348 24480 37360
rect 24400 37292 24412 37348
rect 24468 37292 24480 37348
rect 24400 37028 24480 37292
rect 24400 36972 24412 37028
rect 24468 36972 24480 37028
rect 24400 36960 24480 36972
rect 24560 37348 24640 37360
rect 24560 37292 24572 37348
rect 24628 37292 24640 37348
rect 24560 37028 24640 37292
rect 24560 36972 24572 37028
rect 24628 36972 24640 37028
rect 24560 36960 24640 36972
rect 24720 37348 24800 37360
rect 24720 37292 24732 37348
rect 24788 37292 24800 37348
rect 24720 37028 24800 37292
rect 24720 36972 24732 37028
rect 24788 36972 24800 37028
rect 24720 36960 24800 36972
rect 24880 37348 24960 37360
rect 24880 37292 24892 37348
rect 24948 37292 24960 37348
rect 24880 37028 24960 37292
rect 24880 36972 24892 37028
rect 24948 36972 24960 37028
rect 24880 36960 24960 36972
rect 25040 37348 25120 37360
rect 25040 37292 25052 37348
rect 25108 37292 25120 37348
rect 25040 37028 25120 37292
rect 25040 36972 25052 37028
rect 25108 36972 25120 37028
rect 25040 36960 25120 36972
rect 25200 37348 25280 37360
rect 25200 37292 25212 37348
rect 25268 37292 25280 37348
rect 25200 37028 25280 37292
rect 25200 36972 25212 37028
rect 25268 36972 25280 37028
rect 25200 36960 25280 36972
rect 25360 37348 25440 37360
rect 25360 37292 25372 37348
rect 25428 37292 25440 37348
rect 25360 37028 25440 37292
rect 25360 36972 25372 37028
rect 25428 36972 25440 37028
rect 25360 36960 25440 36972
rect 25520 37348 25600 37360
rect 25520 37292 25532 37348
rect 25588 37292 25600 37348
rect 25520 37028 25600 37292
rect 25520 36972 25532 37028
rect 25588 36972 25600 37028
rect 25520 36960 25600 36972
rect 25680 37348 25760 37360
rect 25680 37292 25692 37348
rect 25748 37292 25760 37348
rect 25680 37028 25760 37292
rect 25680 36972 25692 37028
rect 25748 36972 25760 37028
rect 25680 36960 25760 36972
rect 25840 37348 25920 37360
rect 25840 37292 25852 37348
rect 25908 37292 25920 37348
rect 25840 37028 25920 37292
rect 25840 36972 25852 37028
rect 25908 36972 25920 37028
rect 25840 36960 25920 36972
rect 26000 37348 26080 37360
rect 26000 37292 26012 37348
rect 26068 37292 26080 37348
rect 26000 37028 26080 37292
rect 26000 36972 26012 37028
rect 26068 36972 26080 37028
rect 26000 36960 26080 36972
rect 26160 37348 26240 37360
rect 26160 37292 26172 37348
rect 26228 37292 26240 37348
rect 26160 37028 26240 37292
rect 26160 36972 26172 37028
rect 26228 36972 26240 37028
rect 26160 36960 26240 36972
rect 26320 37348 26400 37360
rect 26320 37292 26332 37348
rect 26388 37292 26400 37348
rect 26320 37028 26400 37292
rect 26320 36972 26332 37028
rect 26388 36972 26400 37028
rect 26320 36960 26400 36972
rect 26480 37348 26560 37360
rect 26480 37292 26492 37348
rect 26548 37292 26560 37348
rect 26480 37028 26560 37292
rect 26480 36972 26492 37028
rect 26548 36972 26560 37028
rect 26480 36960 26560 36972
rect 26640 37348 26720 37360
rect 26640 37292 26652 37348
rect 26708 37292 26720 37348
rect 26640 37028 26720 37292
rect 26640 36972 26652 37028
rect 26708 36972 26720 37028
rect 26640 36960 26720 36972
rect 26800 37348 26880 37360
rect 26800 37292 26812 37348
rect 26868 37292 26880 37348
rect 26800 37028 26880 37292
rect 26800 36972 26812 37028
rect 26868 36972 26880 37028
rect 26800 36960 26880 36972
rect 26960 37348 27040 37360
rect 26960 37292 26972 37348
rect 27028 37292 27040 37348
rect 26960 37028 27040 37292
rect 26960 36972 26972 37028
rect 27028 36972 27040 37028
rect 26960 36960 27040 36972
rect 27120 37348 27200 37360
rect 27120 37292 27132 37348
rect 27188 37292 27200 37348
rect 27120 37028 27200 37292
rect 27120 36972 27132 37028
rect 27188 36972 27200 37028
rect 27120 36960 27200 36972
rect 27280 37348 27360 37360
rect 27280 37292 27292 37348
rect 27348 37292 27360 37348
rect 27280 37028 27360 37292
rect 27280 36972 27292 37028
rect 27348 36972 27360 37028
rect 27280 36960 27360 36972
rect 27440 37348 27520 37360
rect 27440 37292 27452 37348
rect 27508 37292 27520 37348
rect 27440 37028 27520 37292
rect 27440 36972 27452 37028
rect 27508 36972 27520 37028
rect 27440 36960 27520 36972
rect 27600 37348 27680 37360
rect 27600 37292 27612 37348
rect 27668 37292 27680 37348
rect 27600 37028 27680 37292
rect 27600 36972 27612 37028
rect 27668 36972 27680 37028
rect 27600 36960 27680 36972
rect 27760 37348 27840 37360
rect 27760 37292 27772 37348
rect 27828 37292 27840 37348
rect 27760 37028 27840 37292
rect 27760 36972 27772 37028
rect 27828 36972 27840 37028
rect 27760 36960 27840 36972
rect 27920 37348 28000 37360
rect 27920 37292 27932 37348
rect 27988 37292 28000 37348
rect 27920 37028 28000 37292
rect 27920 36972 27932 37028
rect 27988 36972 28000 37028
rect 27920 36960 28000 36972
rect 28080 37348 28160 37360
rect 28080 37292 28092 37348
rect 28148 37292 28160 37348
rect 28080 37028 28160 37292
rect 28080 36972 28092 37028
rect 28148 36972 28160 37028
rect 28080 36960 28160 36972
rect 28240 37348 28320 37360
rect 28240 37292 28252 37348
rect 28308 37292 28320 37348
rect 28240 37028 28320 37292
rect 28240 36972 28252 37028
rect 28308 36972 28320 37028
rect 28240 36960 28320 36972
rect 28400 37348 28480 37360
rect 28400 37292 28412 37348
rect 28468 37292 28480 37348
rect 28400 37028 28480 37292
rect 28400 36972 28412 37028
rect 28468 36972 28480 37028
rect 28400 36960 28480 36972
rect 28560 37348 28640 37360
rect 28560 37292 28572 37348
rect 28628 37292 28640 37348
rect 28560 37028 28640 37292
rect 28560 36972 28572 37028
rect 28628 36972 28640 37028
rect 28560 36960 28640 36972
rect 28720 37348 28800 37360
rect 28720 37292 28732 37348
rect 28788 37292 28800 37348
rect 28720 37028 28800 37292
rect 28720 36972 28732 37028
rect 28788 36972 28800 37028
rect 28720 36960 28800 36972
rect 28880 37348 28960 37360
rect 28880 37292 28892 37348
rect 28948 37292 28960 37348
rect 28880 37028 28960 37292
rect 28880 36972 28892 37028
rect 28948 36972 28960 37028
rect 28880 36960 28960 36972
rect 29040 37348 29120 37360
rect 29040 37292 29052 37348
rect 29108 37292 29120 37348
rect 29040 37028 29120 37292
rect 29040 36972 29052 37028
rect 29108 36972 29120 37028
rect 29040 36960 29120 36972
rect 29200 37348 29280 37360
rect 29200 37292 29212 37348
rect 29268 37292 29280 37348
rect 29200 37028 29280 37292
rect 29200 36972 29212 37028
rect 29268 36972 29280 37028
rect 29200 36960 29280 36972
rect 29360 37348 29440 37360
rect 29360 37292 29372 37348
rect 29428 37292 29440 37348
rect 29360 37028 29440 37292
rect 29360 36972 29372 37028
rect 29428 36972 29440 37028
rect 29360 36960 29440 36972
rect 23120 36868 23200 36880
rect 23120 36812 23132 36868
rect 23188 36812 23200 36868
rect 23120 36548 23200 36812
rect 23120 36492 23132 36548
rect 23188 36492 23200 36548
rect 23120 36480 23200 36492
rect 23280 36868 23360 36880
rect 23280 36812 23292 36868
rect 23348 36812 23360 36868
rect 23280 36548 23360 36812
rect 23280 36492 23292 36548
rect 23348 36492 23360 36548
rect 23280 36480 23360 36492
rect 23440 36868 23520 36880
rect 23440 36812 23452 36868
rect 23508 36812 23520 36868
rect 23440 36548 23520 36812
rect 23440 36492 23452 36548
rect 23508 36492 23520 36548
rect 23440 36480 23520 36492
rect 23600 36868 23680 36880
rect 23600 36812 23612 36868
rect 23668 36812 23680 36868
rect 23600 36548 23680 36812
rect 23600 36492 23612 36548
rect 23668 36492 23680 36548
rect 23600 36480 23680 36492
rect 23760 36868 23840 36880
rect 23760 36812 23772 36868
rect 23828 36812 23840 36868
rect 23760 36548 23840 36812
rect 23760 36492 23772 36548
rect 23828 36492 23840 36548
rect 23760 36480 23840 36492
rect 23920 36868 24000 36880
rect 23920 36812 23932 36868
rect 23988 36812 24000 36868
rect 23920 36548 24000 36812
rect 23920 36492 23932 36548
rect 23988 36492 24000 36548
rect 23920 36480 24000 36492
rect 24080 36868 24160 36880
rect 24080 36812 24092 36868
rect 24148 36812 24160 36868
rect 24080 36548 24160 36812
rect 24080 36492 24092 36548
rect 24148 36492 24160 36548
rect 24080 36480 24160 36492
rect 24240 36868 24320 36880
rect 24240 36812 24252 36868
rect 24308 36812 24320 36868
rect 24240 36548 24320 36812
rect 24240 36492 24252 36548
rect 24308 36492 24320 36548
rect 24240 36480 24320 36492
rect 24400 36868 24480 36880
rect 24400 36812 24412 36868
rect 24468 36812 24480 36868
rect 24400 36548 24480 36812
rect 24400 36492 24412 36548
rect 24468 36492 24480 36548
rect 24400 36480 24480 36492
rect 24560 36868 24640 36880
rect 24560 36812 24572 36868
rect 24628 36812 24640 36868
rect 24560 36548 24640 36812
rect 24560 36492 24572 36548
rect 24628 36492 24640 36548
rect 24560 36480 24640 36492
rect 24720 36868 24800 36880
rect 24720 36812 24732 36868
rect 24788 36812 24800 36868
rect 24720 36548 24800 36812
rect 24720 36492 24732 36548
rect 24788 36492 24800 36548
rect 24720 36480 24800 36492
rect 24880 36868 24960 36880
rect 24880 36812 24892 36868
rect 24948 36812 24960 36868
rect 24880 36548 24960 36812
rect 24880 36492 24892 36548
rect 24948 36492 24960 36548
rect 24880 36480 24960 36492
rect 25040 36868 25120 36880
rect 25040 36812 25052 36868
rect 25108 36812 25120 36868
rect 25040 36548 25120 36812
rect 25040 36492 25052 36548
rect 25108 36492 25120 36548
rect 25040 36480 25120 36492
rect 25200 36868 25280 36880
rect 25200 36812 25212 36868
rect 25268 36812 25280 36868
rect 25200 36548 25280 36812
rect 25200 36492 25212 36548
rect 25268 36492 25280 36548
rect 25200 36480 25280 36492
rect 25360 36868 25440 36880
rect 25360 36812 25372 36868
rect 25428 36812 25440 36868
rect 25360 36548 25440 36812
rect 25360 36492 25372 36548
rect 25428 36492 25440 36548
rect 25360 36480 25440 36492
rect 25520 36868 25600 36880
rect 25520 36812 25532 36868
rect 25588 36812 25600 36868
rect 25520 36548 25600 36812
rect 25520 36492 25532 36548
rect 25588 36492 25600 36548
rect 25520 36480 25600 36492
rect 25680 36868 25760 36880
rect 25680 36812 25692 36868
rect 25748 36812 25760 36868
rect 25680 36548 25760 36812
rect 25680 36492 25692 36548
rect 25748 36492 25760 36548
rect 25680 36480 25760 36492
rect 25840 36868 25920 36880
rect 25840 36812 25852 36868
rect 25908 36812 25920 36868
rect 25840 36548 25920 36812
rect 25840 36492 25852 36548
rect 25908 36492 25920 36548
rect 25840 36480 25920 36492
rect 26000 36868 26080 36880
rect 26000 36812 26012 36868
rect 26068 36812 26080 36868
rect 26000 36548 26080 36812
rect 26000 36492 26012 36548
rect 26068 36492 26080 36548
rect 26000 36480 26080 36492
rect 26160 36868 26240 36880
rect 26160 36812 26172 36868
rect 26228 36812 26240 36868
rect 26160 36548 26240 36812
rect 26160 36492 26172 36548
rect 26228 36492 26240 36548
rect 26160 36480 26240 36492
rect 26320 36868 26400 36880
rect 26320 36812 26332 36868
rect 26388 36812 26400 36868
rect 26320 36548 26400 36812
rect 26320 36492 26332 36548
rect 26388 36492 26400 36548
rect 26320 36480 26400 36492
rect 26480 36868 26560 36880
rect 26480 36812 26492 36868
rect 26548 36812 26560 36868
rect 26480 36548 26560 36812
rect 26480 36492 26492 36548
rect 26548 36492 26560 36548
rect 26480 36480 26560 36492
rect 26640 36868 26720 36880
rect 26640 36812 26652 36868
rect 26708 36812 26720 36868
rect 26640 36548 26720 36812
rect 26640 36492 26652 36548
rect 26708 36492 26720 36548
rect 26640 36480 26720 36492
rect 26800 36868 26880 36880
rect 26800 36812 26812 36868
rect 26868 36812 26880 36868
rect 26800 36548 26880 36812
rect 26800 36492 26812 36548
rect 26868 36492 26880 36548
rect 26800 36480 26880 36492
rect 26960 36868 27040 36880
rect 26960 36812 26972 36868
rect 27028 36812 27040 36868
rect 26960 36548 27040 36812
rect 26960 36492 26972 36548
rect 27028 36492 27040 36548
rect 26960 36480 27040 36492
rect 27120 36868 27200 36880
rect 27120 36812 27132 36868
rect 27188 36812 27200 36868
rect 27120 36548 27200 36812
rect 27120 36492 27132 36548
rect 27188 36492 27200 36548
rect 27120 36480 27200 36492
rect 27280 36868 27360 36880
rect 27280 36812 27292 36868
rect 27348 36812 27360 36868
rect 27280 36548 27360 36812
rect 27280 36492 27292 36548
rect 27348 36492 27360 36548
rect 27280 36480 27360 36492
rect 27440 36868 27520 36880
rect 27440 36812 27452 36868
rect 27508 36812 27520 36868
rect 27440 36548 27520 36812
rect 27440 36492 27452 36548
rect 27508 36492 27520 36548
rect 27440 36480 27520 36492
rect 27600 36868 27680 36880
rect 27600 36812 27612 36868
rect 27668 36812 27680 36868
rect 27600 36548 27680 36812
rect 27600 36492 27612 36548
rect 27668 36492 27680 36548
rect 27600 36480 27680 36492
rect 27760 36868 27840 36880
rect 27760 36812 27772 36868
rect 27828 36812 27840 36868
rect 27760 36548 27840 36812
rect 27760 36492 27772 36548
rect 27828 36492 27840 36548
rect 27760 36480 27840 36492
rect 27920 36868 28000 36880
rect 27920 36812 27932 36868
rect 27988 36812 28000 36868
rect 27920 36548 28000 36812
rect 27920 36492 27932 36548
rect 27988 36492 28000 36548
rect 27920 36480 28000 36492
rect 28080 36868 28160 36880
rect 28080 36812 28092 36868
rect 28148 36812 28160 36868
rect 28080 36548 28160 36812
rect 28080 36492 28092 36548
rect 28148 36492 28160 36548
rect 28080 36480 28160 36492
rect 28240 36868 28320 36880
rect 28240 36812 28252 36868
rect 28308 36812 28320 36868
rect 28240 36548 28320 36812
rect 28240 36492 28252 36548
rect 28308 36492 28320 36548
rect 28240 36480 28320 36492
rect 28400 36868 28480 36880
rect 28400 36812 28412 36868
rect 28468 36812 28480 36868
rect 28400 36548 28480 36812
rect 28400 36492 28412 36548
rect 28468 36492 28480 36548
rect 28400 36480 28480 36492
rect 28560 36868 28640 36880
rect 28560 36812 28572 36868
rect 28628 36812 28640 36868
rect 28560 36548 28640 36812
rect 28560 36492 28572 36548
rect 28628 36492 28640 36548
rect 28560 36480 28640 36492
rect 28720 36868 28800 36880
rect 28720 36812 28732 36868
rect 28788 36812 28800 36868
rect 28720 36548 28800 36812
rect 28720 36492 28732 36548
rect 28788 36492 28800 36548
rect 28720 36480 28800 36492
rect 28880 36868 28960 36880
rect 28880 36812 28892 36868
rect 28948 36812 28960 36868
rect 28880 36548 28960 36812
rect 28880 36492 28892 36548
rect 28948 36492 28960 36548
rect 28880 36480 28960 36492
rect 29040 36868 29120 36880
rect 29040 36812 29052 36868
rect 29108 36812 29120 36868
rect 29040 36548 29120 36812
rect 29040 36492 29052 36548
rect 29108 36492 29120 36548
rect 29040 36480 29120 36492
rect 29200 36868 29280 36880
rect 29200 36812 29212 36868
rect 29268 36812 29280 36868
rect 29200 36548 29280 36812
rect 29200 36492 29212 36548
rect 29268 36492 29280 36548
rect 29200 36480 29280 36492
rect 29360 36868 29440 36880
rect 29360 36812 29372 36868
rect 29428 36812 29440 36868
rect 29360 36548 29440 36812
rect 29360 36492 29372 36548
rect 29428 36492 29440 36548
rect 29360 36480 29440 36492
rect 23120 36388 23200 36400
rect 23120 36332 23132 36388
rect 23188 36332 23200 36388
rect 23120 36068 23200 36332
rect 23120 36012 23132 36068
rect 23188 36012 23200 36068
rect 23120 35748 23200 36012
rect 23120 35692 23132 35748
rect 23188 35692 23200 35748
rect 23120 35428 23200 35692
rect 23120 35372 23132 35428
rect 23188 35372 23200 35428
rect 23120 35108 23200 35372
rect 23120 35052 23132 35108
rect 23188 35052 23200 35108
rect 23120 34788 23200 35052
rect 23120 34732 23132 34788
rect 23188 34732 23200 34788
rect 23120 34468 23200 34732
rect 23120 34412 23132 34468
rect 23188 34412 23200 34468
rect 23120 34400 23200 34412
rect 23280 36388 23360 36400
rect 23280 36332 23292 36388
rect 23348 36332 23360 36388
rect 23280 36068 23360 36332
rect 23280 36012 23292 36068
rect 23348 36012 23360 36068
rect 23280 35748 23360 36012
rect 23280 35692 23292 35748
rect 23348 35692 23360 35748
rect 23280 35428 23360 35692
rect 23280 35372 23292 35428
rect 23348 35372 23360 35428
rect 23280 35108 23360 35372
rect 23280 35052 23292 35108
rect 23348 35052 23360 35108
rect 23280 34788 23360 35052
rect 23280 34732 23292 34788
rect 23348 34732 23360 34788
rect 23280 34468 23360 34732
rect 23280 34412 23292 34468
rect 23348 34412 23360 34468
rect 23280 34400 23360 34412
rect 23440 36388 23520 36400
rect 23440 36332 23452 36388
rect 23508 36332 23520 36388
rect 23440 36068 23520 36332
rect 23440 36012 23452 36068
rect 23508 36012 23520 36068
rect 23440 35748 23520 36012
rect 23440 35692 23452 35748
rect 23508 35692 23520 35748
rect 23440 35428 23520 35692
rect 23440 35372 23452 35428
rect 23508 35372 23520 35428
rect 23440 35108 23520 35372
rect 23440 35052 23452 35108
rect 23508 35052 23520 35108
rect 23440 34788 23520 35052
rect 23440 34732 23452 34788
rect 23508 34732 23520 34788
rect 23440 34468 23520 34732
rect 23440 34412 23452 34468
rect 23508 34412 23520 34468
rect 23440 34400 23520 34412
rect 23600 36388 23680 36400
rect 23600 36332 23612 36388
rect 23668 36332 23680 36388
rect 23600 36068 23680 36332
rect 23600 36012 23612 36068
rect 23668 36012 23680 36068
rect 23600 35748 23680 36012
rect 23600 35692 23612 35748
rect 23668 35692 23680 35748
rect 23600 35428 23680 35692
rect 23600 35372 23612 35428
rect 23668 35372 23680 35428
rect 23600 35108 23680 35372
rect 23600 35052 23612 35108
rect 23668 35052 23680 35108
rect 23600 34788 23680 35052
rect 23600 34732 23612 34788
rect 23668 34732 23680 34788
rect 23600 34468 23680 34732
rect 23600 34412 23612 34468
rect 23668 34412 23680 34468
rect 23600 34400 23680 34412
rect 23760 36388 23840 36400
rect 23760 36332 23772 36388
rect 23828 36332 23840 36388
rect 23760 36068 23840 36332
rect 23760 36012 23772 36068
rect 23828 36012 23840 36068
rect 23760 35748 23840 36012
rect 23760 35692 23772 35748
rect 23828 35692 23840 35748
rect 23760 35428 23840 35692
rect 23760 35372 23772 35428
rect 23828 35372 23840 35428
rect 23760 35108 23840 35372
rect 23760 35052 23772 35108
rect 23828 35052 23840 35108
rect 23760 34788 23840 35052
rect 23760 34732 23772 34788
rect 23828 34732 23840 34788
rect 23760 34468 23840 34732
rect 23760 34412 23772 34468
rect 23828 34412 23840 34468
rect 23760 34400 23840 34412
rect 23920 36388 24000 36400
rect 23920 36332 23932 36388
rect 23988 36332 24000 36388
rect 23920 36068 24000 36332
rect 23920 36012 23932 36068
rect 23988 36012 24000 36068
rect 23920 35748 24000 36012
rect 23920 35692 23932 35748
rect 23988 35692 24000 35748
rect 23920 35428 24000 35692
rect 23920 35372 23932 35428
rect 23988 35372 24000 35428
rect 23920 35108 24000 35372
rect 23920 35052 23932 35108
rect 23988 35052 24000 35108
rect 23920 34788 24000 35052
rect 23920 34732 23932 34788
rect 23988 34732 24000 34788
rect 23920 34468 24000 34732
rect 23920 34412 23932 34468
rect 23988 34412 24000 34468
rect 23920 34400 24000 34412
rect 24080 36388 24160 36400
rect 24080 36332 24092 36388
rect 24148 36332 24160 36388
rect 24080 36068 24160 36332
rect 24080 36012 24092 36068
rect 24148 36012 24160 36068
rect 24080 35748 24160 36012
rect 24080 35692 24092 35748
rect 24148 35692 24160 35748
rect 24080 35428 24160 35692
rect 24080 35372 24092 35428
rect 24148 35372 24160 35428
rect 24080 35108 24160 35372
rect 24080 35052 24092 35108
rect 24148 35052 24160 35108
rect 24080 34788 24160 35052
rect 24080 34732 24092 34788
rect 24148 34732 24160 34788
rect 24080 34468 24160 34732
rect 24080 34412 24092 34468
rect 24148 34412 24160 34468
rect 24080 34400 24160 34412
rect 24240 36388 24320 36400
rect 24240 36332 24252 36388
rect 24308 36332 24320 36388
rect 24240 36068 24320 36332
rect 24240 36012 24252 36068
rect 24308 36012 24320 36068
rect 24240 35748 24320 36012
rect 24240 35692 24252 35748
rect 24308 35692 24320 35748
rect 24240 35428 24320 35692
rect 24240 35372 24252 35428
rect 24308 35372 24320 35428
rect 24240 35108 24320 35372
rect 24240 35052 24252 35108
rect 24308 35052 24320 35108
rect 24240 34788 24320 35052
rect 24240 34732 24252 34788
rect 24308 34732 24320 34788
rect 24240 34468 24320 34732
rect 24240 34412 24252 34468
rect 24308 34412 24320 34468
rect 24240 34400 24320 34412
rect 24400 36388 24480 36400
rect 24400 36332 24412 36388
rect 24468 36332 24480 36388
rect 24400 36068 24480 36332
rect 24400 36012 24412 36068
rect 24468 36012 24480 36068
rect 24400 35748 24480 36012
rect 24400 35692 24412 35748
rect 24468 35692 24480 35748
rect 24400 35428 24480 35692
rect 24400 35372 24412 35428
rect 24468 35372 24480 35428
rect 24400 35108 24480 35372
rect 24400 35052 24412 35108
rect 24468 35052 24480 35108
rect 24400 34788 24480 35052
rect 24400 34732 24412 34788
rect 24468 34732 24480 34788
rect 24400 34468 24480 34732
rect 24400 34412 24412 34468
rect 24468 34412 24480 34468
rect 24400 34400 24480 34412
rect 24560 36388 24640 36400
rect 24560 36332 24572 36388
rect 24628 36332 24640 36388
rect 24560 36068 24640 36332
rect 24560 36012 24572 36068
rect 24628 36012 24640 36068
rect 24560 35748 24640 36012
rect 24560 35692 24572 35748
rect 24628 35692 24640 35748
rect 24560 35428 24640 35692
rect 24560 35372 24572 35428
rect 24628 35372 24640 35428
rect 24560 35108 24640 35372
rect 24560 35052 24572 35108
rect 24628 35052 24640 35108
rect 24560 34788 24640 35052
rect 24560 34732 24572 34788
rect 24628 34732 24640 34788
rect 24560 34468 24640 34732
rect 24560 34412 24572 34468
rect 24628 34412 24640 34468
rect 24560 34400 24640 34412
rect 24720 36388 24800 36400
rect 24720 36332 24732 36388
rect 24788 36332 24800 36388
rect 24720 36068 24800 36332
rect 24720 36012 24732 36068
rect 24788 36012 24800 36068
rect 24720 35748 24800 36012
rect 24720 35692 24732 35748
rect 24788 35692 24800 35748
rect 24720 35428 24800 35692
rect 24720 35372 24732 35428
rect 24788 35372 24800 35428
rect 24720 35108 24800 35372
rect 24720 35052 24732 35108
rect 24788 35052 24800 35108
rect 24720 34788 24800 35052
rect 24720 34732 24732 34788
rect 24788 34732 24800 34788
rect 24720 34468 24800 34732
rect 24720 34412 24732 34468
rect 24788 34412 24800 34468
rect 24720 34400 24800 34412
rect 24880 36388 24960 36400
rect 24880 36332 24892 36388
rect 24948 36332 24960 36388
rect 24880 36068 24960 36332
rect 24880 36012 24892 36068
rect 24948 36012 24960 36068
rect 24880 35748 24960 36012
rect 24880 35692 24892 35748
rect 24948 35692 24960 35748
rect 24880 35428 24960 35692
rect 24880 35372 24892 35428
rect 24948 35372 24960 35428
rect 24880 35108 24960 35372
rect 24880 35052 24892 35108
rect 24948 35052 24960 35108
rect 24880 34788 24960 35052
rect 24880 34732 24892 34788
rect 24948 34732 24960 34788
rect 24880 34468 24960 34732
rect 24880 34412 24892 34468
rect 24948 34412 24960 34468
rect 24880 34400 24960 34412
rect 25040 36388 25120 36400
rect 25040 36332 25052 36388
rect 25108 36332 25120 36388
rect 25040 36068 25120 36332
rect 25040 36012 25052 36068
rect 25108 36012 25120 36068
rect 25040 35748 25120 36012
rect 25040 35692 25052 35748
rect 25108 35692 25120 35748
rect 25040 35428 25120 35692
rect 25040 35372 25052 35428
rect 25108 35372 25120 35428
rect 25040 35108 25120 35372
rect 25040 35052 25052 35108
rect 25108 35052 25120 35108
rect 25040 34788 25120 35052
rect 25040 34732 25052 34788
rect 25108 34732 25120 34788
rect 25040 34468 25120 34732
rect 25040 34412 25052 34468
rect 25108 34412 25120 34468
rect 25040 34400 25120 34412
rect 25200 36388 25280 36400
rect 25200 36332 25212 36388
rect 25268 36332 25280 36388
rect 25200 36068 25280 36332
rect 25200 36012 25212 36068
rect 25268 36012 25280 36068
rect 25200 35748 25280 36012
rect 25200 35692 25212 35748
rect 25268 35692 25280 35748
rect 25200 35428 25280 35692
rect 25200 35372 25212 35428
rect 25268 35372 25280 35428
rect 25200 35108 25280 35372
rect 25200 35052 25212 35108
rect 25268 35052 25280 35108
rect 25200 34788 25280 35052
rect 25200 34732 25212 34788
rect 25268 34732 25280 34788
rect 25200 34468 25280 34732
rect 25200 34412 25212 34468
rect 25268 34412 25280 34468
rect 25200 34400 25280 34412
rect 25360 36388 25440 36400
rect 25360 36332 25372 36388
rect 25428 36332 25440 36388
rect 25360 36068 25440 36332
rect 25360 36012 25372 36068
rect 25428 36012 25440 36068
rect 25360 35748 25440 36012
rect 25360 35692 25372 35748
rect 25428 35692 25440 35748
rect 25360 35428 25440 35692
rect 25360 35372 25372 35428
rect 25428 35372 25440 35428
rect 25360 35108 25440 35372
rect 25360 35052 25372 35108
rect 25428 35052 25440 35108
rect 25360 34788 25440 35052
rect 25360 34732 25372 34788
rect 25428 34732 25440 34788
rect 25360 34468 25440 34732
rect 25360 34412 25372 34468
rect 25428 34412 25440 34468
rect 25360 34400 25440 34412
rect 25520 36388 25600 36400
rect 25520 36332 25532 36388
rect 25588 36332 25600 36388
rect 25520 36068 25600 36332
rect 25520 36012 25532 36068
rect 25588 36012 25600 36068
rect 25520 35748 25600 36012
rect 25520 35692 25532 35748
rect 25588 35692 25600 35748
rect 25520 35428 25600 35692
rect 25520 35372 25532 35428
rect 25588 35372 25600 35428
rect 25520 35108 25600 35372
rect 25520 35052 25532 35108
rect 25588 35052 25600 35108
rect 25520 34788 25600 35052
rect 25520 34732 25532 34788
rect 25588 34732 25600 34788
rect 25520 34468 25600 34732
rect 25520 34412 25532 34468
rect 25588 34412 25600 34468
rect 25520 34400 25600 34412
rect 25680 36388 25760 36400
rect 25680 36332 25692 36388
rect 25748 36332 25760 36388
rect 25680 36068 25760 36332
rect 25680 36012 25692 36068
rect 25748 36012 25760 36068
rect 25680 35748 25760 36012
rect 25680 35692 25692 35748
rect 25748 35692 25760 35748
rect 25680 35428 25760 35692
rect 25680 35372 25692 35428
rect 25748 35372 25760 35428
rect 25680 35108 25760 35372
rect 25680 35052 25692 35108
rect 25748 35052 25760 35108
rect 25680 34788 25760 35052
rect 25680 34732 25692 34788
rect 25748 34732 25760 34788
rect 25680 34468 25760 34732
rect 25680 34412 25692 34468
rect 25748 34412 25760 34468
rect 25680 34400 25760 34412
rect 25840 36388 25920 36400
rect 25840 36332 25852 36388
rect 25908 36332 25920 36388
rect 25840 36068 25920 36332
rect 25840 36012 25852 36068
rect 25908 36012 25920 36068
rect 25840 35748 25920 36012
rect 25840 35692 25852 35748
rect 25908 35692 25920 35748
rect 25840 35428 25920 35692
rect 25840 35372 25852 35428
rect 25908 35372 25920 35428
rect 25840 35108 25920 35372
rect 25840 35052 25852 35108
rect 25908 35052 25920 35108
rect 25840 34788 25920 35052
rect 25840 34732 25852 34788
rect 25908 34732 25920 34788
rect 25840 34468 25920 34732
rect 25840 34412 25852 34468
rect 25908 34412 25920 34468
rect 25840 34400 25920 34412
rect 26000 36388 26080 36400
rect 26000 36332 26012 36388
rect 26068 36332 26080 36388
rect 26000 36068 26080 36332
rect 26000 36012 26012 36068
rect 26068 36012 26080 36068
rect 26000 35748 26080 36012
rect 26000 35692 26012 35748
rect 26068 35692 26080 35748
rect 26000 35428 26080 35692
rect 26000 35372 26012 35428
rect 26068 35372 26080 35428
rect 26000 35108 26080 35372
rect 26000 35052 26012 35108
rect 26068 35052 26080 35108
rect 26000 34788 26080 35052
rect 26000 34732 26012 34788
rect 26068 34732 26080 34788
rect 26000 34468 26080 34732
rect 26000 34412 26012 34468
rect 26068 34412 26080 34468
rect 26000 34400 26080 34412
rect 26160 36388 26240 36400
rect 26160 36332 26172 36388
rect 26228 36332 26240 36388
rect 26160 36068 26240 36332
rect 26160 36012 26172 36068
rect 26228 36012 26240 36068
rect 26160 35748 26240 36012
rect 26160 35692 26172 35748
rect 26228 35692 26240 35748
rect 26160 35428 26240 35692
rect 26160 35372 26172 35428
rect 26228 35372 26240 35428
rect 26160 35108 26240 35372
rect 26160 35052 26172 35108
rect 26228 35052 26240 35108
rect 26160 34788 26240 35052
rect 26160 34732 26172 34788
rect 26228 34732 26240 34788
rect 26160 34468 26240 34732
rect 26160 34412 26172 34468
rect 26228 34412 26240 34468
rect 26160 34400 26240 34412
rect 26320 36388 26400 36400
rect 26320 36332 26332 36388
rect 26388 36332 26400 36388
rect 26320 36068 26400 36332
rect 26320 36012 26332 36068
rect 26388 36012 26400 36068
rect 26320 35748 26400 36012
rect 26320 35692 26332 35748
rect 26388 35692 26400 35748
rect 26320 35428 26400 35692
rect 26320 35372 26332 35428
rect 26388 35372 26400 35428
rect 26320 35108 26400 35372
rect 26320 35052 26332 35108
rect 26388 35052 26400 35108
rect 26320 34788 26400 35052
rect 26320 34732 26332 34788
rect 26388 34732 26400 34788
rect 26320 34468 26400 34732
rect 26320 34412 26332 34468
rect 26388 34412 26400 34468
rect 26320 34400 26400 34412
rect 26480 36388 26560 36400
rect 26480 36332 26492 36388
rect 26548 36332 26560 36388
rect 26480 36068 26560 36332
rect 26480 36012 26492 36068
rect 26548 36012 26560 36068
rect 26480 35748 26560 36012
rect 26480 35692 26492 35748
rect 26548 35692 26560 35748
rect 26480 35428 26560 35692
rect 26480 35372 26492 35428
rect 26548 35372 26560 35428
rect 26480 35108 26560 35372
rect 26480 35052 26492 35108
rect 26548 35052 26560 35108
rect 26480 34788 26560 35052
rect 26480 34732 26492 34788
rect 26548 34732 26560 34788
rect 26480 34468 26560 34732
rect 26480 34412 26492 34468
rect 26548 34412 26560 34468
rect 26480 34400 26560 34412
rect 26640 36388 26720 36400
rect 26640 36332 26652 36388
rect 26708 36332 26720 36388
rect 26640 36068 26720 36332
rect 26640 36012 26652 36068
rect 26708 36012 26720 36068
rect 26640 35748 26720 36012
rect 26640 35692 26652 35748
rect 26708 35692 26720 35748
rect 26640 35428 26720 35692
rect 26640 35372 26652 35428
rect 26708 35372 26720 35428
rect 26640 35108 26720 35372
rect 26640 35052 26652 35108
rect 26708 35052 26720 35108
rect 26640 34788 26720 35052
rect 26640 34732 26652 34788
rect 26708 34732 26720 34788
rect 26640 34468 26720 34732
rect 26640 34412 26652 34468
rect 26708 34412 26720 34468
rect 26640 34400 26720 34412
rect 26800 36388 26880 36400
rect 26800 36332 26812 36388
rect 26868 36332 26880 36388
rect 26800 36068 26880 36332
rect 26800 36012 26812 36068
rect 26868 36012 26880 36068
rect 26800 35748 26880 36012
rect 26800 35692 26812 35748
rect 26868 35692 26880 35748
rect 26800 35428 26880 35692
rect 26800 35372 26812 35428
rect 26868 35372 26880 35428
rect 26800 35108 26880 35372
rect 26800 35052 26812 35108
rect 26868 35052 26880 35108
rect 26800 34788 26880 35052
rect 26800 34732 26812 34788
rect 26868 34732 26880 34788
rect 26800 34468 26880 34732
rect 26800 34412 26812 34468
rect 26868 34412 26880 34468
rect 26800 34400 26880 34412
rect 26960 36388 27040 36400
rect 26960 36332 26972 36388
rect 27028 36332 27040 36388
rect 26960 36068 27040 36332
rect 26960 36012 26972 36068
rect 27028 36012 27040 36068
rect 26960 35748 27040 36012
rect 26960 35692 26972 35748
rect 27028 35692 27040 35748
rect 26960 35428 27040 35692
rect 26960 35372 26972 35428
rect 27028 35372 27040 35428
rect 26960 35108 27040 35372
rect 26960 35052 26972 35108
rect 27028 35052 27040 35108
rect 26960 34788 27040 35052
rect 26960 34732 26972 34788
rect 27028 34732 27040 34788
rect 26960 34468 27040 34732
rect 26960 34412 26972 34468
rect 27028 34412 27040 34468
rect 26960 34400 27040 34412
rect 27120 36388 27200 36400
rect 27120 36332 27132 36388
rect 27188 36332 27200 36388
rect 27120 36068 27200 36332
rect 27120 36012 27132 36068
rect 27188 36012 27200 36068
rect 27120 35748 27200 36012
rect 27120 35692 27132 35748
rect 27188 35692 27200 35748
rect 27120 35428 27200 35692
rect 27120 35372 27132 35428
rect 27188 35372 27200 35428
rect 27120 35108 27200 35372
rect 27120 35052 27132 35108
rect 27188 35052 27200 35108
rect 27120 34788 27200 35052
rect 27120 34732 27132 34788
rect 27188 34732 27200 34788
rect 27120 34468 27200 34732
rect 27120 34412 27132 34468
rect 27188 34412 27200 34468
rect 27120 34400 27200 34412
rect 27280 36388 27360 36400
rect 27280 36332 27292 36388
rect 27348 36332 27360 36388
rect 27280 36068 27360 36332
rect 27280 36012 27292 36068
rect 27348 36012 27360 36068
rect 27280 35748 27360 36012
rect 27280 35692 27292 35748
rect 27348 35692 27360 35748
rect 27280 35428 27360 35692
rect 27280 35372 27292 35428
rect 27348 35372 27360 35428
rect 27280 35108 27360 35372
rect 27280 35052 27292 35108
rect 27348 35052 27360 35108
rect 27280 34788 27360 35052
rect 27280 34732 27292 34788
rect 27348 34732 27360 34788
rect 27280 34468 27360 34732
rect 27280 34412 27292 34468
rect 27348 34412 27360 34468
rect 27280 34400 27360 34412
rect 27440 36388 27520 36400
rect 27440 36332 27452 36388
rect 27508 36332 27520 36388
rect 27440 36068 27520 36332
rect 27440 36012 27452 36068
rect 27508 36012 27520 36068
rect 27440 35748 27520 36012
rect 27440 35692 27452 35748
rect 27508 35692 27520 35748
rect 27440 35428 27520 35692
rect 27440 35372 27452 35428
rect 27508 35372 27520 35428
rect 27440 35108 27520 35372
rect 27440 35052 27452 35108
rect 27508 35052 27520 35108
rect 27440 34788 27520 35052
rect 27440 34732 27452 34788
rect 27508 34732 27520 34788
rect 27440 34468 27520 34732
rect 27440 34412 27452 34468
rect 27508 34412 27520 34468
rect 27440 34400 27520 34412
rect 27600 36388 27680 36400
rect 27600 36332 27612 36388
rect 27668 36332 27680 36388
rect 27600 36068 27680 36332
rect 27600 36012 27612 36068
rect 27668 36012 27680 36068
rect 27600 35748 27680 36012
rect 27600 35692 27612 35748
rect 27668 35692 27680 35748
rect 27600 35428 27680 35692
rect 27600 35372 27612 35428
rect 27668 35372 27680 35428
rect 27600 35108 27680 35372
rect 27600 35052 27612 35108
rect 27668 35052 27680 35108
rect 27600 34788 27680 35052
rect 27600 34732 27612 34788
rect 27668 34732 27680 34788
rect 27600 34468 27680 34732
rect 27600 34412 27612 34468
rect 27668 34412 27680 34468
rect 27600 34400 27680 34412
rect 27760 36388 27840 36400
rect 27760 36332 27772 36388
rect 27828 36332 27840 36388
rect 27760 36068 27840 36332
rect 27760 36012 27772 36068
rect 27828 36012 27840 36068
rect 27760 35748 27840 36012
rect 27760 35692 27772 35748
rect 27828 35692 27840 35748
rect 27760 35428 27840 35692
rect 27760 35372 27772 35428
rect 27828 35372 27840 35428
rect 27760 35108 27840 35372
rect 27760 35052 27772 35108
rect 27828 35052 27840 35108
rect 27760 34788 27840 35052
rect 27760 34732 27772 34788
rect 27828 34732 27840 34788
rect 27760 34468 27840 34732
rect 27760 34412 27772 34468
rect 27828 34412 27840 34468
rect 27760 34400 27840 34412
rect 27920 36388 28000 36400
rect 27920 36332 27932 36388
rect 27988 36332 28000 36388
rect 27920 36068 28000 36332
rect 27920 36012 27932 36068
rect 27988 36012 28000 36068
rect 27920 35748 28000 36012
rect 27920 35692 27932 35748
rect 27988 35692 28000 35748
rect 27920 35428 28000 35692
rect 27920 35372 27932 35428
rect 27988 35372 28000 35428
rect 27920 35108 28000 35372
rect 27920 35052 27932 35108
rect 27988 35052 28000 35108
rect 27920 34788 28000 35052
rect 27920 34732 27932 34788
rect 27988 34732 28000 34788
rect 27920 34468 28000 34732
rect 27920 34412 27932 34468
rect 27988 34412 28000 34468
rect 27920 34400 28000 34412
rect 28080 36388 28160 36400
rect 28080 36332 28092 36388
rect 28148 36332 28160 36388
rect 28080 36068 28160 36332
rect 28080 36012 28092 36068
rect 28148 36012 28160 36068
rect 28080 35748 28160 36012
rect 28080 35692 28092 35748
rect 28148 35692 28160 35748
rect 28080 35428 28160 35692
rect 28080 35372 28092 35428
rect 28148 35372 28160 35428
rect 28080 35108 28160 35372
rect 28080 35052 28092 35108
rect 28148 35052 28160 35108
rect 28080 34788 28160 35052
rect 28080 34732 28092 34788
rect 28148 34732 28160 34788
rect 28080 34468 28160 34732
rect 28080 34412 28092 34468
rect 28148 34412 28160 34468
rect 28080 34400 28160 34412
rect 28240 36388 28320 36400
rect 28240 36332 28252 36388
rect 28308 36332 28320 36388
rect 28240 36068 28320 36332
rect 28240 36012 28252 36068
rect 28308 36012 28320 36068
rect 28240 35748 28320 36012
rect 28240 35692 28252 35748
rect 28308 35692 28320 35748
rect 28240 35428 28320 35692
rect 28240 35372 28252 35428
rect 28308 35372 28320 35428
rect 28240 35108 28320 35372
rect 28240 35052 28252 35108
rect 28308 35052 28320 35108
rect 28240 34788 28320 35052
rect 28240 34732 28252 34788
rect 28308 34732 28320 34788
rect 28240 34468 28320 34732
rect 28240 34412 28252 34468
rect 28308 34412 28320 34468
rect 28240 34400 28320 34412
rect 28400 36388 28480 36400
rect 28400 36332 28412 36388
rect 28468 36332 28480 36388
rect 28400 36068 28480 36332
rect 28400 36012 28412 36068
rect 28468 36012 28480 36068
rect 28400 35748 28480 36012
rect 28400 35692 28412 35748
rect 28468 35692 28480 35748
rect 28400 35428 28480 35692
rect 28400 35372 28412 35428
rect 28468 35372 28480 35428
rect 28400 35108 28480 35372
rect 28400 35052 28412 35108
rect 28468 35052 28480 35108
rect 28400 34788 28480 35052
rect 28400 34732 28412 34788
rect 28468 34732 28480 34788
rect 28400 34468 28480 34732
rect 28400 34412 28412 34468
rect 28468 34412 28480 34468
rect 28400 34400 28480 34412
rect 28560 36388 28640 36400
rect 28560 36332 28572 36388
rect 28628 36332 28640 36388
rect 28560 36068 28640 36332
rect 28560 36012 28572 36068
rect 28628 36012 28640 36068
rect 28560 35748 28640 36012
rect 28560 35692 28572 35748
rect 28628 35692 28640 35748
rect 28560 35428 28640 35692
rect 28560 35372 28572 35428
rect 28628 35372 28640 35428
rect 28560 35108 28640 35372
rect 28560 35052 28572 35108
rect 28628 35052 28640 35108
rect 28560 34788 28640 35052
rect 28560 34732 28572 34788
rect 28628 34732 28640 34788
rect 28560 34468 28640 34732
rect 28560 34412 28572 34468
rect 28628 34412 28640 34468
rect 28560 34400 28640 34412
rect 28720 36388 28800 36400
rect 28720 36332 28732 36388
rect 28788 36332 28800 36388
rect 28720 36068 28800 36332
rect 28720 36012 28732 36068
rect 28788 36012 28800 36068
rect 28720 35748 28800 36012
rect 28720 35692 28732 35748
rect 28788 35692 28800 35748
rect 28720 35428 28800 35692
rect 28720 35372 28732 35428
rect 28788 35372 28800 35428
rect 28720 35108 28800 35372
rect 28720 35052 28732 35108
rect 28788 35052 28800 35108
rect 28720 34788 28800 35052
rect 28720 34732 28732 34788
rect 28788 34732 28800 34788
rect 28720 34468 28800 34732
rect 28720 34412 28732 34468
rect 28788 34412 28800 34468
rect 28720 34400 28800 34412
rect 28880 36388 28960 36400
rect 28880 36332 28892 36388
rect 28948 36332 28960 36388
rect 28880 36068 28960 36332
rect 28880 36012 28892 36068
rect 28948 36012 28960 36068
rect 28880 35748 28960 36012
rect 28880 35692 28892 35748
rect 28948 35692 28960 35748
rect 28880 35428 28960 35692
rect 28880 35372 28892 35428
rect 28948 35372 28960 35428
rect 28880 35108 28960 35372
rect 28880 35052 28892 35108
rect 28948 35052 28960 35108
rect 28880 34788 28960 35052
rect 28880 34732 28892 34788
rect 28948 34732 28960 34788
rect 28880 34468 28960 34732
rect 28880 34412 28892 34468
rect 28948 34412 28960 34468
rect 28880 34400 28960 34412
rect 29040 36388 29120 36400
rect 29040 36332 29052 36388
rect 29108 36332 29120 36388
rect 29040 36068 29120 36332
rect 29040 36012 29052 36068
rect 29108 36012 29120 36068
rect 29040 35748 29120 36012
rect 29040 35692 29052 35748
rect 29108 35692 29120 35748
rect 29040 35428 29120 35692
rect 29040 35372 29052 35428
rect 29108 35372 29120 35428
rect 29040 35108 29120 35372
rect 29040 35052 29052 35108
rect 29108 35052 29120 35108
rect 29040 34788 29120 35052
rect 29040 34732 29052 34788
rect 29108 34732 29120 34788
rect 29040 34468 29120 34732
rect 29040 34412 29052 34468
rect 29108 34412 29120 34468
rect 29040 34400 29120 34412
rect 29200 36388 29280 36400
rect 29200 36332 29212 36388
rect 29268 36332 29280 36388
rect 29200 36068 29280 36332
rect 29200 36012 29212 36068
rect 29268 36012 29280 36068
rect 29200 35748 29280 36012
rect 29200 35692 29212 35748
rect 29268 35692 29280 35748
rect 29200 35428 29280 35692
rect 29200 35372 29212 35428
rect 29268 35372 29280 35428
rect 29200 35108 29280 35372
rect 29200 35052 29212 35108
rect 29268 35052 29280 35108
rect 29200 34788 29280 35052
rect 29200 34732 29212 34788
rect 29268 34732 29280 34788
rect 29200 34468 29280 34732
rect 29200 34412 29212 34468
rect 29268 34412 29280 34468
rect 29200 34400 29280 34412
rect 29360 36388 29440 36400
rect 29360 36332 29372 36388
rect 29428 36332 29440 36388
rect 29360 36068 29440 36332
rect 29360 36012 29372 36068
rect 29428 36012 29440 36068
rect 29360 35748 29440 36012
rect 29360 35692 29372 35748
rect 29428 35692 29440 35748
rect 29360 35428 29440 35692
rect 29360 35372 29372 35428
rect 29428 35372 29440 35428
rect 29360 35108 29440 35372
rect 29360 35052 29372 35108
rect 29428 35052 29440 35108
rect 29360 34788 29440 35052
rect 29360 34732 29372 34788
rect 29428 34732 29440 34788
rect 29360 34468 29440 34732
rect 29360 34412 29372 34468
rect 29428 34412 29440 34468
rect 29360 34400 29440 34412
rect 23120 34308 23200 34320
rect 23120 34252 23132 34308
rect 23188 34252 23200 34308
rect 23120 33988 23200 34252
rect 23120 33932 23132 33988
rect 23188 33932 23200 33988
rect 23120 33920 23200 33932
rect 23280 34308 23360 34320
rect 23280 34252 23292 34308
rect 23348 34252 23360 34308
rect 23280 33988 23360 34252
rect 23280 33932 23292 33988
rect 23348 33932 23360 33988
rect 23280 33920 23360 33932
rect 23440 34308 23520 34320
rect 23440 34252 23452 34308
rect 23508 34252 23520 34308
rect 23440 33988 23520 34252
rect 23440 33932 23452 33988
rect 23508 33932 23520 33988
rect 23440 33920 23520 33932
rect 23600 34308 23680 34320
rect 23600 34252 23612 34308
rect 23668 34252 23680 34308
rect 23600 33988 23680 34252
rect 23600 33932 23612 33988
rect 23668 33932 23680 33988
rect 23600 33920 23680 33932
rect 23760 34308 23840 34320
rect 23760 34252 23772 34308
rect 23828 34252 23840 34308
rect 23760 33988 23840 34252
rect 23760 33932 23772 33988
rect 23828 33932 23840 33988
rect 23760 33920 23840 33932
rect 23920 34308 24000 34320
rect 23920 34252 23932 34308
rect 23988 34252 24000 34308
rect 23920 33988 24000 34252
rect 23920 33932 23932 33988
rect 23988 33932 24000 33988
rect 23920 33920 24000 33932
rect 24080 34308 24160 34320
rect 24080 34252 24092 34308
rect 24148 34252 24160 34308
rect 24080 33988 24160 34252
rect 24080 33932 24092 33988
rect 24148 33932 24160 33988
rect 24080 33920 24160 33932
rect 24240 34308 24320 34320
rect 24240 34252 24252 34308
rect 24308 34252 24320 34308
rect 24240 33988 24320 34252
rect 24240 33932 24252 33988
rect 24308 33932 24320 33988
rect 24240 33920 24320 33932
rect 24400 34308 24480 34320
rect 24400 34252 24412 34308
rect 24468 34252 24480 34308
rect 24400 33988 24480 34252
rect 24400 33932 24412 33988
rect 24468 33932 24480 33988
rect 24400 33920 24480 33932
rect 24560 34308 24640 34320
rect 24560 34252 24572 34308
rect 24628 34252 24640 34308
rect 24560 33988 24640 34252
rect 24560 33932 24572 33988
rect 24628 33932 24640 33988
rect 24560 33920 24640 33932
rect 24720 34308 24800 34320
rect 24720 34252 24732 34308
rect 24788 34252 24800 34308
rect 24720 33988 24800 34252
rect 24720 33932 24732 33988
rect 24788 33932 24800 33988
rect 24720 33920 24800 33932
rect 24880 34308 24960 34320
rect 24880 34252 24892 34308
rect 24948 34252 24960 34308
rect 24880 33988 24960 34252
rect 24880 33932 24892 33988
rect 24948 33932 24960 33988
rect 24880 33920 24960 33932
rect 25040 34308 25120 34320
rect 25040 34252 25052 34308
rect 25108 34252 25120 34308
rect 25040 33988 25120 34252
rect 25040 33932 25052 33988
rect 25108 33932 25120 33988
rect 25040 33920 25120 33932
rect 25200 34308 25280 34320
rect 25200 34252 25212 34308
rect 25268 34252 25280 34308
rect 25200 33988 25280 34252
rect 25200 33932 25212 33988
rect 25268 33932 25280 33988
rect 25200 33920 25280 33932
rect 25360 34308 25440 34320
rect 25360 34252 25372 34308
rect 25428 34252 25440 34308
rect 25360 33988 25440 34252
rect 25360 33932 25372 33988
rect 25428 33932 25440 33988
rect 25360 33920 25440 33932
rect 25520 34308 25600 34320
rect 25520 34252 25532 34308
rect 25588 34252 25600 34308
rect 25520 33988 25600 34252
rect 25520 33932 25532 33988
rect 25588 33932 25600 33988
rect 25520 33920 25600 33932
rect 25680 34308 25760 34320
rect 25680 34252 25692 34308
rect 25748 34252 25760 34308
rect 25680 33988 25760 34252
rect 25680 33932 25692 33988
rect 25748 33932 25760 33988
rect 25680 33920 25760 33932
rect 25840 34308 25920 34320
rect 25840 34252 25852 34308
rect 25908 34252 25920 34308
rect 25840 33988 25920 34252
rect 25840 33932 25852 33988
rect 25908 33932 25920 33988
rect 25840 33920 25920 33932
rect 26000 34308 26080 34320
rect 26000 34252 26012 34308
rect 26068 34252 26080 34308
rect 26000 33988 26080 34252
rect 26000 33932 26012 33988
rect 26068 33932 26080 33988
rect 26000 33920 26080 33932
rect 26160 34308 26240 34320
rect 26160 34252 26172 34308
rect 26228 34252 26240 34308
rect 26160 33988 26240 34252
rect 26160 33932 26172 33988
rect 26228 33932 26240 33988
rect 26160 33920 26240 33932
rect 26320 34308 26400 34320
rect 26320 34252 26332 34308
rect 26388 34252 26400 34308
rect 26320 33988 26400 34252
rect 26320 33932 26332 33988
rect 26388 33932 26400 33988
rect 26320 33920 26400 33932
rect 26480 34308 26560 34320
rect 26480 34252 26492 34308
rect 26548 34252 26560 34308
rect 26480 33988 26560 34252
rect 26480 33932 26492 33988
rect 26548 33932 26560 33988
rect 26480 33920 26560 33932
rect 26640 34308 26720 34320
rect 26640 34252 26652 34308
rect 26708 34252 26720 34308
rect 26640 33988 26720 34252
rect 26640 33932 26652 33988
rect 26708 33932 26720 33988
rect 26640 33920 26720 33932
rect 26800 34308 26880 34320
rect 26800 34252 26812 34308
rect 26868 34252 26880 34308
rect 26800 33988 26880 34252
rect 26800 33932 26812 33988
rect 26868 33932 26880 33988
rect 26800 33920 26880 33932
rect 26960 34308 27040 34320
rect 26960 34252 26972 34308
rect 27028 34252 27040 34308
rect 26960 33988 27040 34252
rect 26960 33932 26972 33988
rect 27028 33932 27040 33988
rect 26960 33920 27040 33932
rect 27120 34308 27200 34320
rect 27120 34252 27132 34308
rect 27188 34252 27200 34308
rect 27120 33988 27200 34252
rect 27120 33932 27132 33988
rect 27188 33932 27200 33988
rect 27120 33920 27200 33932
rect 27280 34308 27360 34320
rect 27280 34252 27292 34308
rect 27348 34252 27360 34308
rect 27280 33988 27360 34252
rect 27280 33932 27292 33988
rect 27348 33932 27360 33988
rect 27280 33920 27360 33932
rect 27440 34308 27520 34320
rect 27440 34252 27452 34308
rect 27508 34252 27520 34308
rect 27440 33988 27520 34252
rect 27440 33932 27452 33988
rect 27508 33932 27520 33988
rect 27440 33920 27520 33932
rect 27600 34308 27680 34320
rect 27600 34252 27612 34308
rect 27668 34252 27680 34308
rect 27600 33988 27680 34252
rect 27600 33932 27612 33988
rect 27668 33932 27680 33988
rect 27600 33920 27680 33932
rect 27760 34308 27840 34320
rect 27760 34252 27772 34308
rect 27828 34252 27840 34308
rect 27760 33988 27840 34252
rect 27760 33932 27772 33988
rect 27828 33932 27840 33988
rect 27760 33920 27840 33932
rect 27920 34308 28000 34320
rect 27920 34252 27932 34308
rect 27988 34252 28000 34308
rect 27920 33988 28000 34252
rect 27920 33932 27932 33988
rect 27988 33932 28000 33988
rect 27920 33920 28000 33932
rect 28080 34308 28160 34320
rect 28080 34252 28092 34308
rect 28148 34252 28160 34308
rect 28080 33988 28160 34252
rect 28080 33932 28092 33988
rect 28148 33932 28160 33988
rect 28080 33920 28160 33932
rect 28240 34308 28320 34320
rect 28240 34252 28252 34308
rect 28308 34252 28320 34308
rect 28240 33988 28320 34252
rect 28240 33932 28252 33988
rect 28308 33932 28320 33988
rect 28240 33920 28320 33932
rect 28400 34308 28480 34320
rect 28400 34252 28412 34308
rect 28468 34252 28480 34308
rect 28400 33988 28480 34252
rect 28400 33932 28412 33988
rect 28468 33932 28480 33988
rect 28400 33920 28480 33932
rect 28560 34308 28640 34320
rect 28560 34252 28572 34308
rect 28628 34252 28640 34308
rect 28560 33988 28640 34252
rect 28560 33932 28572 33988
rect 28628 33932 28640 33988
rect 28560 33920 28640 33932
rect 28720 34308 28800 34320
rect 28720 34252 28732 34308
rect 28788 34252 28800 34308
rect 28720 33988 28800 34252
rect 28720 33932 28732 33988
rect 28788 33932 28800 33988
rect 28720 33920 28800 33932
rect 28880 34308 28960 34320
rect 28880 34252 28892 34308
rect 28948 34252 28960 34308
rect 28880 33988 28960 34252
rect 28880 33932 28892 33988
rect 28948 33932 28960 33988
rect 28880 33920 28960 33932
rect 29040 34308 29120 34320
rect 29040 34252 29052 34308
rect 29108 34252 29120 34308
rect 29040 33988 29120 34252
rect 29040 33932 29052 33988
rect 29108 33932 29120 33988
rect 29040 33920 29120 33932
rect 29200 34308 29280 34320
rect 29200 34252 29212 34308
rect 29268 34252 29280 34308
rect 29200 33988 29280 34252
rect 29200 33932 29212 33988
rect 29268 33932 29280 33988
rect 29200 33920 29280 33932
rect 29360 34308 29440 34320
rect 29360 34252 29372 34308
rect 29428 34252 29440 34308
rect 29360 33988 29440 34252
rect 29360 33932 29372 33988
rect 29428 33932 29440 33988
rect 29360 33920 29440 33932
rect 23120 33828 23200 33840
rect 23120 33772 23132 33828
rect 23188 33772 23200 33828
rect 23120 33508 23200 33772
rect 23120 33452 23132 33508
rect 23188 33452 23200 33508
rect 23120 33440 23200 33452
rect 23280 33828 23360 33840
rect 23280 33772 23292 33828
rect 23348 33772 23360 33828
rect 23280 33508 23360 33772
rect 23280 33452 23292 33508
rect 23348 33452 23360 33508
rect 23280 33440 23360 33452
rect 23440 33828 23520 33840
rect 23440 33772 23452 33828
rect 23508 33772 23520 33828
rect 23440 33508 23520 33772
rect 23440 33452 23452 33508
rect 23508 33452 23520 33508
rect 23440 33440 23520 33452
rect 23600 33828 23680 33840
rect 23600 33772 23612 33828
rect 23668 33772 23680 33828
rect 23600 33508 23680 33772
rect 23600 33452 23612 33508
rect 23668 33452 23680 33508
rect 23600 33440 23680 33452
rect 23760 33828 23840 33840
rect 23760 33772 23772 33828
rect 23828 33772 23840 33828
rect 23760 33508 23840 33772
rect 23760 33452 23772 33508
rect 23828 33452 23840 33508
rect 23760 33440 23840 33452
rect 23920 33828 24000 33840
rect 23920 33772 23932 33828
rect 23988 33772 24000 33828
rect 23920 33508 24000 33772
rect 23920 33452 23932 33508
rect 23988 33452 24000 33508
rect 23920 33440 24000 33452
rect 24080 33828 24160 33840
rect 24080 33772 24092 33828
rect 24148 33772 24160 33828
rect 24080 33508 24160 33772
rect 24080 33452 24092 33508
rect 24148 33452 24160 33508
rect 24080 33440 24160 33452
rect 24240 33828 24320 33840
rect 24240 33772 24252 33828
rect 24308 33772 24320 33828
rect 24240 33508 24320 33772
rect 24240 33452 24252 33508
rect 24308 33452 24320 33508
rect 24240 33440 24320 33452
rect 24400 33828 24480 33840
rect 24400 33772 24412 33828
rect 24468 33772 24480 33828
rect 24400 33508 24480 33772
rect 24400 33452 24412 33508
rect 24468 33452 24480 33508
rect 24400 33440 24480 33452
rect 24560 33828 24640 33840
rect 24560 33772 24572 33828
rect 24628 33772 24640 33828
rect 24560 33508 24640 33772
rect 24560 33452 24572 33508
rect 24628 33452 24640 33508
rect 24560 33440 24640 33452
rect 24720 33828 24800 33840
rect 24720 33772 24732 33828
rect 24788 33772 24800 33828
rect 24720 33508 24800 33772
rect 24720 33452 24732 33508
rect 24788 33452 24800 33508
rect 24720 33440 24800 33452
rect 24880 33828 24960 33840
rect 24880 33772 24892 33828
rect 24948 33772 24960 33828
rect 24880 33508 24960 33772
rect 24880 33452 24892 33508
rect 24948 33452 24960 33508
rect 24880 33440 24960 33452
rect 25040 33828 25120 33840
rect 25040 33772 25052 33828
rect 25108 33772 25120 33828
rect 25040 33508 25120 33772
rect 25040 33452 25052 33508
rect 25108 33452 25120 33508
rect 25040 33440 25120 33452
rect 25200 33828 25280 33840
rect 25200 33772 25212 33828
rect 25268 33772 25280 33828
rect 25200 33508 25280 33772
rect 25200 33452 25212 33508
rect 25268 33452 25280 33508
rect 25200 33440 25280 33452
rect 25360 33828 25440 33840
rect 25360 33772 25372 33828
rect 25428 33772 25440 33828
rect 25360 33508 25440 33772
rect 25360 33452 25372 33508
rect 25428 33452 25440 33508
rect 25360 33440 25440 33452
rect 25520 33828 25600 33840
rect 25520 33772 25532 33828
rect 25588 33772 25600 33828
rect 25520 33508 25600 33772
rect 25520 33452 25532 33508
rect 25588 33452 25600 33508
rect 25520 33440 25600 33452
rect 25680 33828 25760 33840
rect 25680 33772 25692 33828
rect 25748 33772 25760 33828
rect 25680 33508 25760 33772
rect 25680 33452 25692 33508
rect 25748 33452 25760 33508
rect 25680 33440 25760 33452
rect 25840 33828 25920 33840
rect 25840 33772 25852 33828
rect 25908 33772 25920 33828
rect 25840 33508 25920 33772
rect 25840 33452 25852 33508
rect 25908 33452 25920 33508
rect 25840 33440 25920 33452
rect 26000 33828 26080 33840
rect 26000 33772 26012 33828
rect 26068 33772 26080 33828
rect 26000 33508 26080 33772
rect 26000 33452 26012 33508
rect 26068 33452 26080 33508
rect 26000 33440 26080 33452
rect 26160 33828 26240 33840
rect 26160 33772 26172 33828
rect 26228 33772 26240 33828
rect 26160 33508 26240 33772
rect 26160 33452 26172 33508
rect 26228 33452 26240 33508
rect 26160 33440 26240 33452
rect 26320 33828 26400 33840
rect 26320 33772 26332 33828
rect 26388 33772 26400 33828
rect 26320 33508 26400 33772
rect 26320 33452 26332 33508
rect 26388 33452 26400 33508
rect 26320 33440 26400 33452
rect 26480 33828 26560 33840
rect 26480 33772 26492 33828
rect 26548 33772 26560 33828
rect 26480 33508 26560 33772
rect 26480 33452 26492 33508
rect 26548 33452 26560 33508
rect 26480 33440 26560 33452
rect 26640 33828 26720 33840
rect 26640 33772 26652 33828
rect 26708 33772 26720 33828
rect 26640 33508 26720 33772
rect 26640 33452 26652 33508
rect 26708 33452 26720 33508
rect 26640 33440 26720 33452
rect 26800 33828 26880 33840
rect 26800 33772 26812 33828
rect 26868 33772 26880 33828
rect 26800 33508 26880 33772
rect 26800 33452 26812 33508
rect 26868 33452 26880 33508
rect 26800 33440 26880 33452
rect 26960 33828 27040 33840
rect 26960 33772 26972 33828
rect 27028 33772 27040 33828
rect 26960 33508 27040 33772
rect 26960 33452 26972 33508
rect 27028 33452 27040 33508
rect 26960 33440 27040 33452
rect 27120 33828 27200 33840
rect 27120 33772 27132 33828
rect 27188 33772 27200 33828
rect 27120 33508 27200 33772
rect 27120 33452 27132 33508
rect 27188 33452 27200 33508
rect 27120 33440 27200 33452
rect 27280 33828 27360 33840
rect 27280 33772 27292 33828
rect 27348 33772 27360 33828
rect 27280 33508 27360 33772
rect 27280 33452 27292 33508
rect 27348 33452 27360 33508
rect 27280 33440 27360 33452
rect 27440 33828 27520 33840
rect 27440 33772 27452 33828
rect 27508 33772 27520 33828
rect 27440 33508 27520 33772
rect 27440 33452 27452 33508
rect 27508 33452 27520 33508
rect 27440 33440 27520 33452
rect 27600 33828 27680 33840
rect 27600 33772 27612 33828
rect 27668 33772 27680 33828
rect 27600 33508 27680 33772
rect 27600 33452 27612 33508
rect 27668 33452 27680 33508
rect 27600 33440 27680 33452
rect 27760 33828 27840 33840
rect 27760 33772 27772 33828
rect 27828 33772 27840 33828
rect 27760 33508 27840 33772
rect 27760 33452 27772 33508
rect 27828 33452 27840 33508
rect 27760 33440 27840 33452
rect 27920 33828 28000 33840
rect 27920 33772 27932 33828
rect 27988 33772 28000 33828
rect 27920 33508 28000 33772
rect 27920 33452 27932 33508
rect 27988 33452 28000 33508
rect 27920 33440 28000 33452
rect 28080 33828 28160 33840
rect 28080 33772 28092 33828
rect 28148 33772 28160 33828
rect 28080 33508 28160 33772
rect 28080 33452 28092 33508
rect 28148 33452 28160 33508
rect 28080 33440 28160 33452
rect 28240 33828 28320 33840
rect 28240 33772 28252 33828
rect 28308 33772 28320 33828
rect 28240 33508 28320 33772
rect 28240 33452 28252 33508
rect 28308 33452 28320 33508
rect 28240 33440 28320 33452
rect 28400 33828 28480 33840
rect 28400 33772 28412 33828
rect 28468 33772 28480 33828
rect 28400 33508 28480 33772
rect 28400 33452 28412 33508
rect 28468 33452 28480 33508
rect 28400 33440 28480 33452
rect 28560 33828 28640 33840
rect 28560 33772 28572 33828
rect 28628 33772 28640 33828
rect 28560 33508 28640 33772
rect 28560 33452 28572 33508
rect 28628 33452 28640 33508
rect 28560 33440 28640 33452
rect 28720 33828 28800 33840
rect 28720 33772 28732 33828
rect 28788 33772 28800 33828
rect 28720 33508 28800 33772
rect 28720 33452 28732 33508
rect 28788 33452 28800 33508
rect 28720 33440 28800 33452
rect 28880 33828 28960 33840
rect 28880 33772 28892 33828
rect 28948 33772 28960 33828
rect 28880 33508 28960 33772
rect 28880 33452 28892 33508
rect 28948 33452 28960 33508
rect 28880 33440 28960 33452
rect 29040 33828 29120 33840
rect 29040 33772 29052 33828
rect 29108 33772 29120 33828
rect 29040 33508 29120 33772
rect 29040 33452 29052 33508
rect 29108 33452 29120 33508
rect 29040 33440 29120 33452
rect 29200 33828 29280 33840
rect 29200 33772 29212 33828
rect 29268 33772 29280 33828
rect 29200 33508 29280 33772
rect 29200 33452 29212 33508
rect 29268 33452 29280 33508
rect 29200 33440 29280 33452
rect 29360 33828 29440 33840
rect 29360 33772 29372 33828
rect 29428 33772 29440 33828
rect 29360 33508 29440 33772
rect 29360 33452 29372 33508
rect 29428 33452 29440 33508
rect 29360 33440 29440 33452
rect 29520 33828 29600 37440
rect 29520 33772 29532 33828
rect 29588 33772 29600 33828
rect 29520 33508 29600 33772
rect 29520 33452 29532 33508
rect 29588 33452 29600 33508
rect 29520 33440 29600 33452
rect 29680 33668 29760 37440
rect 29680 33612 29692 33668
rect 29748 33612 29760 33668
rect 29680 33440 29760 33612
rect 29840 33828 29920 37440
rect 29840 33772 29852 33828
rect 29908 33772 29920 33828
rect 29840 33508 29920 33772
rect 29840 33452 29852 33508
rect 29908 33452 29920 33508
rect 29840 33440 29920 33452
rect 30000 34308 30080 37440
rect 30000 34252 30012 34308
rect 30068 34252 30080 34308
rect 30000 33988 30080 34252
rect 30000 33932 30012 33988
rect 30068 33932 30080 33988
rect 30000 33440 30080 33932
rect 30160 34148 30240 37440
rect 30160 34092 30172 34148
rect 30228 34092 30240 34148
rect 30160 33440 30240 34092
rect 30320 34308 30400 37440
rect 30320 34252 30332 34308
rect 30388 34252 30400 34308
rect 30320 33988 30400 34252
rect 30320 33932 30332 33988
rect 30388 33932 30400 33988
rect 30320 33440 30400 33932
rect 30480 36388 30560 37440
rect 30480 36332 30492 36388
rect 30548 36332 30560 36388
rect 30480 36068 30560 36332
rect 30480 36012 30492 36068
rect 30548 36012 30560 36068
rect 30480 35748 30560 36012
rect 30480 35692 30492 35748
rect 30548 35692 30560 35748
rect 30480 35428 30560 35692
rect 30480 35372 30492 35428
rect 30548 35372 30560 35428
rect 30480 35108 30560 35372
rect 30480 35052 30492 35108
rect 30548 35052 30560 35108
rect 30480 34788 30560 35052
rect 30480 34732 30492 34788
rect 30548 34732 30560 34788
rect 30480 34468 30560 34732
rect 30480 34412 30492 34468
rect 30548 34412 30560 34468
rect 30480 33440 30560 34412
rect 30640 34628 30720 37440
rect 30640 34572 30652 34628
rect 30708 34572 30720 34628
rect 30640 33440 30720 34572
rect 30800 36388 30880 37440
rect 30800 36332 30812 36388
rect 30868 36332 30880 36388
rect 30800 36068 30880 36332
rect 30800 36012 30812 36068
rect 30868 36012 30880 36068
rect 30800 35748 30880 36012
rect 30800 35692 30812 35748
rect 30868 35692 30880 35748
rect 30800 35428 30880 35692
rect 30800 35372 30812 35428
rect 30868 35372 30880 35428
rect 30800 35108 30880 35372
rect 30800 35052 30812 35108
rect 30868 35052 30880 35108
rect 30800 34788 30880 35052
rect 30800 34732 30812 34788
rect 30868 34732 30880 34788
rect 30800 34468 30880 34732
rect 30800 34412 30812 34468
rect 30868 34412 30880 34468
rect 30800 33440 30880 34412
rect 30960 34948 31040 37440
rect 30960 34892 30972 34948
rect 31028 34892 31040 34948
rect 30960 33440 31040 34892
rect 31120 36388 31200 37440
rect 31120 36332 31132 36388
rect 31188 36332 31200 36388
rect 31120 36068 31200 36332
rect 31120 36012 31132 36068
rect 31188 36012 31200 36068
rect 31120 35748 31200 36012
rect 31120 35692 31132 35748
rect 31188 35692 31200 35748
rect 31120 35428 31200 35692
rect 31120 35372 31132 35428
rect 31188 35372 31200 35428
rect 31120 35108 31200 35372
rect 31120 35052 31132 35108
rect 31188 35052 31200 35108
rect 31120 34788 31200 35052
rect 31120 34732 31132 34788
rect 31188 34732 31200 34788
rect 31120 34468 31200 34732
rect 31120 34412 31132 34468
rect 31188 34412 31200 34468
rect 31120 33440 31200 34412
rect 31280 35268 31360 37440
rect 31280 35212 31292 35268
rect 31348 35212 31360 35268
rect 31280 33440 31360 35212
rect 31440 36388 31520 37440
rect 31440 36332 31452 36388
rect 31508 36332 31520 36388
rect 31440 36068 31520 36332
rect 31440 36012 31452 36068
rect 31508 36012 31520 36068
rect 31440 35748 31520 36012
rect 31440 35692 31452 35748
rect 31508 35692 31520 35748
rect 31440 35428 31520 35692
rect 31440 35372 31452 35428
rect 31508 35372 31520 35428
rect 31440 35108 31520 35372
rect 31440 35052 31452 35108
rect 31508 35052 31520 35108
rect 31440 34788 31520 35052
rect 31440 34732 31452 34788
rect 31508 34732 31520 34788
rect 31440 34468 31520 34732
rect 31440 34412 31452 34468
rect 31508 34412 31520 34468
rect 31440 33440 31520 34412
rect 31600 35588 31680 37440
rect 31600 35532 31612 35588
rect 31668 35532 31680 35588
rect 31600 33440 31680 35532
rect 31760 36388 31840 37440
rect 31760 36332 31772 36388
rect 31828 36332 31840 36388
rect 31760 36068 31840 36332
rect 31760 36012 31772 36068
rect 31828 36012 31840 36068
rect 31760 35748 31840 36012
rect 31760 35692 31772 35748
rect 31828 35692 31840 35748
rect 31760 35428 31840 35692
rect 31760 35372 31772 35428
rect 31828 35372 31840 35428
rect 31760 35108 31840 35372
rect 31760 35052 31772 35108
rect 31828 35052 31840 35108
rect 31760 34788 31840 35052
rect 31760 34732 31772 34788
rect 31828 34732 31840 34788
rect 31760 34468 31840 34732
rect 31760 34412 31772 34468
rect 31828 34412 31840 34468
rect 31760 33440 31840 34412
rect 31920 35908 32000 37440
rect 31920 35852 31932 35908
rect 31988 35852 32000 35908
rect 31920 33440 32000 35852
rect 32080 36388 32160 37440
rect 32080 36332 32092 36388
rect 32148 36332 32160 36388
rect 32080 36068 32160 36332
rect 32080 36012 32092 36068
rect 32148 36012 32160 36068
rect 32080 35748 32160 36012
rect 32080 35692 32092 35748
rect 32148 35692 32160 35748
rect 32080 35428 32160 35692
rect 32080 35372 32092 35428
rect 32148 35372 32160 35428
rect 32080 35108 32160 35372
rect 32080 35052 32092 35108
rect 32148 35052 32160 35108
rect 32080 34788 32160 35052
rect 32080 34732 32092 34788
rect 32148 34732 32160 34788
rect 32080 34468 32160 34732
rect 32080 34412 32092 34468
rect 32148 34412 32160 34468
rect 32080 33440 32160 34412
rect 32240 36228 32320 37440
rect 32240 36172 32252 36228
rect 32308 36172 32320 36228
rect 32240 33440 32320 36172
rect 32400 36388 32480 37440
rect 32400 36332 32412 36388
rect 32468 36332 32480 36388
rect 32400 36068 32480 36332
rect 32400 36012 32412 36068
rect 32468 36012 32480 36068
rect 32400 35748 32480 36012
rect 32400 35692 32412 35748
rect 32468 35692 32480 35748
rect 32400 35428 32480 35692
rect 32400 35372 32412 35428
rect 32468 35372 32480 35428
rect 32400 35108 32480 35372
rect 32400 35052 32412 35108
rect 32468 35052 32480 35108
rect 32400 34788 32480 35052
rect 32400 34732 32412 34788
rect 32468 34732 32480 34788
rect 32400 34468 32480 34732
rect 32400 34412 32412 34468
rect 32468 34412 32480 34468
rect 32400 33440 32480 34412
rect 32560 36868 32640 37440
rect 32560 36812 32572 36868
rect 32628 36812 32640 36868
rect 32560 36548 32640 36812
rect 32560 36492 32572 36548
rect 32628 36492 32640 36548
rect 32560 33440 32640 36492
rect 32720 36708 32800 37440
rect 32720 36652 32732 36708
rect 32788 36652 32800 36708
rect 32720 33440 32800 36652
rect 32880 36868 32960 37440
rect 32880 36812 32892 36868
rect 32948 36812 32960 36868
rect 32880 36548 32960 36812
rect 32880 36492 32892 36548
rect 32948 36492 32960 36548
rect 32880 33440 32960 36492
rect 33040 37348 33120 37440
rect 33040 37292 33052 37348
rect 33108 37292 33120 37348
rect 33040 37028 33120 37292
rect 33040 36972 33052 37028
rect 33108 36972 33120 37028
rect 33040 33440 33120 36972
rect 33200 37188 33280 37440
rect 33200 37132 33212 37188
rect 33268 37132 33280 37188
rect 33200 33440 33280 37132
rect 33360 37348 33440 37440
rect 33360 37292 33372 37348
rect 33428 37292 33440 37348
rect 33360 37028 33440 37292
rect 33360 36972 33372 37028
rect 33428 36972 33440 37028
rect 33360 33440 33440 36972
rect 33520 37348 33600 37360
rect 33520 37292 33532 37348
rect 33588 37292 33600 37348
rect 33520 37028 33600 37292
rect 33520 36972 33532 37028
rect 33588 36972 33600 37028
rect 33520 36960 33600 36972
rect 33680 37348 33760 37360
rect 33680 37292 33692 37348
rect 33748 37292 33760 37348
rect 33680 37028 33760 37292
rect 33680 36972 33692 37028
rect 33748 36972 33760 37028
rect 33680 36960 33760 36972
rect 33840 37348 33920 37360
rect 33840 37292 33852 37348
rect 33908 37292 33920 37348
rect 33840 37028 33920 37292
rect 33840 36972 33852 37028
rect 33908 36972 33920 37028
rect 33840 36960 33920 36972
rect 34000 37348 34080 37360
rect 34000 37292 34012 37348
rect 34068 37292 34080 37348
rect 34000 37028 34080 37292
rect 34000 36972 34012 37028
rect 34068 36972 34080 37028
rect 34000 36960 34080 36972
rect 34160 37348 34240 37360
rect 34160 37292 34172 37348
rect 34228 37292 34240 37348
rect 34160 37028 34240 37292
rect 34160 36972 34172 37028
rect 34228 36972 34240 37028
rect 34160 36960 34240 36972
rect 34320 37348 34400 37360
rect 34320 37292 34332 37348
rect 34388 37292 34400 37348
rect 34320 37028 34400 37292
rect 34320 36972 34332 37028
rect 34388 36972 34400 37028
rect 34320 36960 34400 36972
rect 34480 37348 34560 37360
rect 34480 37292 34492 37348
rect 34548 37292 34560 37348
rect 34480 37028 34560 37292
rect 34480 36972 34492 37028
rect 34548 36972 34560 37028
rect 34480 36960 34560 36972
rect 34640 37348 34720 37360
rect 34640 37292 34652 37348
rect 34708 37292 34720 37348
rect 34640 37028 34720 37292
rect 34640 36972 34652 37028
rect 34708 36972 34720 37028
rect 34640 36960 34720 36972
rect 34800 37348 34880 37360
rect 34800 37292 34812 37348
rect 34868 37292 34880 37348
rect 34800 37028 34880 37292
rect 34800 36972 34812 37028
rect 34868 36972 34880 37028
rect 34800 36960 34880 36972
rect 34960 37348 35040 37360
rect 34960 37292 34972 37348
rect 35028 37292 35040 37348
rect 34960 37028 35040 37292
rect 34960 36972 34972 37028
rect 35028 36972 35040 37028
rect 34960 36960 35040 36972
rect 35120 37348 35200 37360
rect 35120 37292 35132 37348
rect 35188 37292 35200 37348
rect 35120 37028 35200 37292
rect 35120 36972 35132 37028
rect 35188 36972 35200 37028
rect 35120 36960 35200 36972
rect 35280 37348 35360 37360
rect 35280 37292 35292 37348
rect 35348 37292 35360 37348
rect 35280 37028 35360 37292
rect 35280 36972 35292 37028
rect 35348 36972 35360 37028
rect 35280 36960 35360 36972
rect 35440 37348 35520 37360
rect 35440 37292 35452 37348
rect 35508 37292 35520 37348
rect 35440 37028 35520 37292
rect 35440 36972 35452 37028
rect 35508 36972 35520 37028
rect 35440 36960 35520 36972
rect 35600 37348 35680 37360
rect 35600 37292 35612 37348
rect 35668 37292 35680 37348
rect 35600 37028 35680 37292
rect 35600 36972 35612 37028
rect 35668 36972 35680 37028
rect 35600 36960 35680 36972
rect 35760 37348 35840 37360
rect 35760 37292 35772 37348
rect 35828 37292 35840 37348
rect 35760 37028 35840 37292
rect 35760 36972 35772 37028
rect 35828 36972 35840 37028
rect 35760 36960 35840 36972
rect 35920 37348 36000 37360
rect 35920 37292 35932 37348
rect 35988 37292 36000 37348
rect 35920 37028 36000 37292
rect 35920 36972 35932 37028
rect 35988 36972 36000 37028
rect 35920 36960 36000 36972
rect 36080 37348 36160 37360
rect 36080 37292 36092 37348
rect 36148 37292 36160 37348
rect 36080 37028 36160 37292
rect 36080 36972 36092 37028
rect 36148 36972 36160 37028
rect 36080 36960 36160 36972
rect 36240 37348 36320 37360
rect 36240 37292 36252 37348
rect 36308 37292 36320 37348
rect 36240 37028 36320 37292
rect 36240 36972 36252 37028
rect 36308 36972 36320 37028
rect 36240 36960 36320 36972
rect 36400 37348 36480 37360
rect 36400 37292 36412 37348
rect 36468 37292 36480 37348
rect 36400 37028 36480 37292
rect 36400 36972 36412 37028
rect 36468 36972 36480 37028
rect 36400 36960 36480 36972
rect 36560 37348 36640 37360
rect 36560 37292 36572 37348
rect 36628 37292 36640 37348
rect 36560 37028 36640 37292
rect 36560 36972 36572 37028
rect 36628 36972 36640 37028
rect 36560 36960 36640 36972
rect 36720 37348 36800 37360
rect 36720 37292 36732 37348
rect 36788 37292 36800 37348
rect 36720 37028 36800 37292
rect 36720 36972 36732 37028
rect 36788 36972 36800 37028
rect 36720 36960 36800 36972
rect 36880 37348 36960 37360
rect 36880 37292 36892 37348
rect 36948 37292 36960 37348
rect 36880 37028 36960 37292
rect 36880 36972 36892 37028
rect 36948 36972 36960 37028
rect 36880 36960 36960 36972
rect 37040 37348 37120 37360
rect 37040 37292 37052 37348
rect 37108 37292 37120 37348
rect 37040 37028 37120 37292
rect 37040 36972 37052 37028
rect 37108 36972 37120 37028
rect 37040 36960 37120 36972
rect 37200 37348 37280 37360
rect 37200 37292 37212 37348
rect 37268 37292 37280 37348
rect 37200 37028 37280 37292
rect 37200 36972 37212 37028
rect 37268 36972 37280 37028
rect 37200 36960 37280 36972
rect 37360 37348 37440 37360
rect 37360 37292 37372 37348
rect 37428 37292 37440 37348
rect 37360 37028 37440 37292
rect 37360 36972 37372 37028
rect 37428 36972 37440 37028
rect 37360 36960 37440 36972
rect 37520 37348 37600 37360
rect 37520 37292 37532 37348
rect 37588 37292 37600 37348
rect 37520 37028 37600 37292
rect 37520 36972 37532 37028
rect 37588 36972 37600 37028
rect 37520 36960 37600 36972
rect 37680 37348 37760 37360
rect 37680 37292 37692 37348
rect 37748 37292 37760 37348
rect 37680 37028 37760 37292
rect 37680 36972 37692 37028
rect 37748 36972 37760 37028
rect 37680 36960 37760 36972
rect 37840 37348 37920 37360
rect 37840 37292 37852 37348
rect 37908 37292 37920 37348
rect 37840 37028 37920 37292
rect 37840 36972 37852 37028
rect 37908 36972 37920 37028
rect 37840 36960 37920 36972
rect 38000 37348 38080 37360
rect 38000 37292 38012 37348
rect 38068 37292 38080 37348
rect 38000 37028 38080 37292
rect 38000 36972 38012 37028
rect 38068 36972 38080 37028
rect 38000 36960 38080 36972
rect 38160 37348 38240 37360
rect 38160 37292 38172 37348
rect 38228 37292 38240 37348
rect 38160 37028 38240 37292
rect 38160 36972 38172 37028
rect 38228 36972 38240 37028
rect 38160 36960 38240 36972
rect 38320 37348 38400 37360
rect 38320 37292 38332 37348
rect 38388 37292 38400 37348
rect 38320 37028 38400 37292
rect 38320 36972 38332 37028
rect 38388 36972 38400 37028
rect 38320 36960 38400 36972
rect 38480 37348 38560 37360
rect 38480 37292 38492 37348
rect 38548 37292 38560 37348
rect 38480 37028 38560 37292
rect 38480 36972 38492 37028
rect 38548 36972 38560 37028
rect 38480 36960 38560 36972
rect 38640 37348 38720 37360
rect 38640 37292 38652 37348
rect 38708 37292 38720 37348
rect 38640 37028 38720 37292
rect 38640 36972 38652 37028
rect 38708 36972 38720 37028
rect 38640 36960 38720 36972
rect 38800 37348 38880 37360
rect 38800 37292 38812 37348
rect 38868 37292 38880 37348
rect 38800 37028 38880 37292
rect 38800 36972 38812 37028
rect 38868 36972 38880 37028
rect 38800 36960 38880 36972
rect 38960 37348 39040 37360
rect 38960 37292 38972 37348
rect 39028 37292 39040 37348
rect 38960 37028 39040 37292
rect 38960 36972 38972 37028
rect 39028 36972 39040 37028
rect 38960 36960 39040 36972
rect 39120 37348 39200 37360
rect 39120 37292 39132 37348
rect 39188 37292 39200 37348
rect 39120 37028 39200 37292
rect 39120 36972 39132 37028
rect 39188 36972 39200 37028
rect 39120 36960 39200 36972
rect 39280 37348 39360 37360
rect 39280 37292 39292 37348
rect 39348 37292 39360 37348
rect 39280 37028 39360 37292
rect 39280 36972 39292 37028
rect 39348 36972 39360 37028
rect 39280 36960 39360 36972
rect 39440 37348 39520 37360
rect 39440 37292 39452 37348
rect 39508 37292 39520 37348
rect 39440 37028 39520 37292
rect 39440 36972 39452 37028
rect 39508 36972 39520 37028
rect 39440 36960 39520 36972
rect 39600 37348 39680 37360
rect 39600 37292 39612 37348
rect 39668 37292 39680 37348
rect 39600 37028 39680 37292
rect 39600 36972 39612 37028
rect 39668 36972 39680 37028
rect 39600 36960 39680 36972
rect 39760 37348 39840 37360
rect 39760 37292 39772 37348
rect 39828 37292 39840 37348
rect 39760 37028 39840 37292
rect 39760 36972 39772 37028
rect 39828 36972 39840 37028
rect 39760 36960 39840 36972
rect 39920 37348 40000 37360
rect 39920 37292 39932 37348
rect 39988 37292 40000 37348
rect 39920 37028 40000 37292
rect 39920 36972 39932 37028
rect 39988 36972 40000 37028
rect 39920 36960 40000 36972
rect 40080 37348 40160 37360
rect 40080 37292 40092 37348
rect 40148 37292 40160 37348
rect 40080 37028 40160 37292
rect 40080 36972 40092 37028
rect 40148 36972 40160 37028
rect 40080 36960 40160 36972
rect 40240 37348 40320 37360
rect 40240 37292 40252 37348
rect 40308 37292 40320 37348
rect 40240 37028 40320 37292
rect 40240 36972 40252 37028
rect 40308 36972 40320 37028
rect 40240 36960 40320 36972
rect 40400 37348 40480 37360
rect 40400 37292 40412 37348
rect 40468 37292 40480 37348
rect 40400 37028 40480 37292
rect 40400 36972 40412 37028
rect 40468 36972 40480 37028
rect 40400 36960 40480 36972
rect 40560 37348 40640 37360
rect 40560 37292 40572 37348
rect 40628 37292 40640 37348
rect 40560 37028 40640 37292
rect 40560 36972 40572 37028
rect 40628 36972 40640 37028
rect 40560 36960 40640 36972
rect 40720 37348 40800 37360
rect 40720 37292 40732 37348
rect 40788 37292 40800 37348
rect 40720 37028 40800 37292
rect 40720 36972 40732 37028
rect 40788 36972 40800 37028
rect 40720 36960 40800 36972
rect 40880 37348 40960 37360
rect 40880 37292 40892 37348
rect 40948 37292 40960 37348
rect 40880 37028 40960 37292
rect 40880 36972 40892 37028
rect 40948 36972 40960 37028
rect 40880 36960 40960 36972
rect 41040 37348 41120 37360
rect 41040 37292 41052 37348
rect 41108 37292 41120 37348
rect 41040 37028 41120 37292
rect 41040 36972 41052 37028
rect 41108 36972 41120 37028
rect 41040 36960 41120 36972
rect 41200 37348 41280 37360
rect 41200 37292 41212 37348
rect 41268 37292 41280 37348
rect 41200 37028 41280 37292
rect 41200 36972 41212 37028
rect 41268 36972 41280 37028
rect 41200 36960 41280 36972
rect 41360 37348 41440 37360
rect 41360 37292 41372 37348
rect 41428 37292 41440 37348
rect 41360 37028 41440 37292
rect 41360 36972 41372 37028
rect 41428 36972 41440 37028
rect 41360 36960 41440 36972
rect 41520 37348 41600 37360
rect 41520 37292 41532 37348
rect 41588 37292 41600 37348
rect 41520 37028 41600 37292
rect 41520 36972 41532 37028
rect 41588 36972 41600 37028
rect 41520 36960 41600 36972
rect 41680 37348 41760 37360
rect 41680 37292 41692 37348
rect 41748 37292 41760 37348
rect 41680 37028 41760 37292
rect 41680 36972 41692 37028
rect 41748 36972 41760 37028
rect 41680 36960 41760 36972
rect 41840 37348 41920 37360
rect 41840 37292 41852 37348
rect 41908 37292 41920 37348
rect 41840 37028 41920 37292
rect 41840 36972 41852 37028
rect 41908 36972 41920 37028
rect 41840 36960 41920 36972
rect 33520 36868 33600 36880
rect 33520 36812 33532 36868
rect 33588 36812 33600 36868
rect 33520 36548 33600 36812
rect 33520 36492 33532 36548
rect 33588 36492 33600 36548
rect 33520 36480 33600 36492
rect 33680 36868 33760 36880
rect 33680 36812 33692 36868
rect 33748 36812 33760 36868
rect 33680 36548 33760 36812
rect 33680 36492 33692 36548
rect 33748 36492 33760 36548
rect 33680 36480 33760 36492
rect 33840 36868 33920 36880
rect 33840 36812 33852 36868
rect 33908 36812 33920 36868
rect 33840 36548 33920 36812
rect 33840 36492 33852 36548
rect 33908 36492 33920 36548
rect 33840 36480 33920 36492
rect 34000 36868 34080 36880
rect 34000 36812 34012 36868
rect 34068 36812 34080 36868
rect 34000 36548 34080 36812
rect 34000 36492 34012 36548
rect 34068 36492 34080 36548
rect 34000 36480 34080 36492
rect 34160 36868 34240 36880
rect 34160 36812 34172 36868
rect 34228 36812 34240 36868
rect 34160 36548 34240 36812
rect 34160 36492 34172 36548
rect 34228 36492 34240 36548
rect 34160 36480 34240 36492
rect 34320 36868 34400 36880
rect 34320 36812 34332 36868
rect 34388 36812 34400 36868
rect 34320 36548 34400 36812
rect 34320 36492 34332 36548
rect 34388 36492 34400 36548
rect 34320 36480 34400 36492
rect 34480 36868 34560 36880
rect 34480 36812 34492 36868
rect 34548 36812 34560 36868
rect 34480 36548 34560 36812
rect 34480 36492 34492 36548
rect 34548 36492 34560 36548
rect 34480 36480 34560 36492
rect 34640 36868 34720 36880
rect 34640 36812 34652 36868
rect 34708 36812 34720 36868
rect 34640 36548 34720 36812
rect 34640 36492 34652 36548
rect 34708 36492 34720 36548
rect 34640 36480 34720 36492
rect 34800 36868 34880 36880
rect 34800 36812 34812 36868
rect 34868 36812 34880 36868
rect 34800 36548 34880 36812
rect 34800 36492 34812 36548
rect 34868 36492 34880 36548
rect 34800 36480 34880 36492
rect 34960 36868 35040 36880
rect 34960 36812 34972 36868
rect 35028 36812 35040 36868
rect 34960 36548 35040 36812
rect 34960 36492 34972 36548
rect 35028 36492 35040 36548
rect 34960 36480 35040 36492
rect 35120 36868 35200 36880
rect 35120 36812 35132 36868
rect 35188 36812 35200 36868
rect 35120 36548 35200 36812
rect 35120 36492 35132 36548
rect 35188 36492 35200 36548
rect 35120 36480 35200 36492
rect 35280 36868 35360 36880
rect 35280 36812 35292 36868
rect 35348 36812 35360 36868
rect 35280 36548 35360 36812
rect 35280 36492 35292 36548
rect 35348 36492 35360 36548
rect 35280 36480 35360 36492
rect 35440 36868 35520 36880
rect 35440 36812 35452 36868
rect 35508 36812 35520 36868
rect 35440 36548 35520 36812
rect 35440 36492 35452 36548
rect 35508 36492 35520 36548
rect 35440 36480 35520 36492
rect 35600 36868 35680 36880
rect 35600 36812 35612 36868
rect 35668 36812 35680 36868
rect 35600 36548 35680 36812
rect 35600 36492 35612 36548
rect 35668 36492 35680 36548
rect 35600 36480 35680 36492
rect 35760 36868 35840 36880
rect 35760 36812 35772 36868
rect 35828 36812 35840 36868
rect 35760 36548 35840 36812
rect 35760 36492 35772 36548
rect 35828 36492 35840 36548
rect 35760 36480 35840 36492
rect 35920 36868 36000 36880
rect 35920 36812 35932 36868
rect 35988 36812 36000 36868
rect 35920 36548 36000 36812
rect 35920 36492 35932 36548
rect 35988 36492 36000 36548
rect 35920 36480 36000 36492
rect 36080 36868 36160 36880
rect 36080 36812 36092 36868
rect 36148 36812 36160 36868
rect 36080 36548 36160 36812
rect 36080 36492 36092 36548
rect 36148 36492 36160 36548
rect 36080 36480 36160 36492
rect 36240 36868 36320 36880
rect 36240 36812 36252 36868
rect 36308 36812 36320 36868
rect 36240 36548 36320 36812
rect 36240 36492 36252 36548
rect 36308 36492 36320 36548
rect 36240 36480 36320 36492
rect 36400 36868 36480 36880
rect 36400 36812 36412 36868
rect 36468 36812 36480 36868
rect 36400 36548 36480 36812
rect 36400 36492 36412 36548
rect 36468 36492 36480 36548
rect 36400 36480 36480 36492
rect 36560 36868 36640 36880
rect 36560 36812 36572 36868
rect 36628 36812 36640 36868
rect 36560 36548 36640 36812
rect 36560 36492 36572 36548
rect 36628 36492 36640 36548
rect 36560 36480 36640 36492
rect 36720 36868 36800 36880
rect 36720 36812 36732 36868
rect 36788 36812 36800 36868
rect 36720 36548 36800 36812
rect 36720 36492 36732 36548
rect 36788 36492 36800 36548
rect 36720 36480 36800 36492
rect 36880 36868 36960 36880
rect 36880 36812 36892 36868
rect 36948 36812 36960 36868
rect 36880 36548 36960 36812
rect 36880 36492 36892 36548
rect 36948 36492 36960 36548
rect 36880 36480 36960 36492
rect 37040 36868 37120 36880
rect 37040 36812 37052 36868
rect 37108 36812 37120 36868
rect 37040 36548 37120 36812
rect 37040 36492 37052 36548
rect 37108 36492 37120 36548
rect 37040 36480 37120 36492
rect 37200 36868 37280 36880
rect 37200 36812 37212 36868
rect 37268 36812 37280 36868
rect 37200 36548 37280 36812
rect 37200 36492 37212 36548
rect 37268 36492 37280 36548
rect 37200 36480 37280 36492
rect 37360 36868 37440 36880
rect 37360 36812 37372 36868
rect 37428 36812 37440 36868
rect 37360 36548 37440 36812
rect 37360 36492 37372 36548
rect 37428 36492 37440 36548
rect 37360 36480 37440 36492
rect 37520 36868 37600 36880
rect 37520 36812 37532 36868
rect 37588 36812 37600 36868
rect 37520 36548 37600 36812
rect 37520 36492 37532 36548
rect 37588 36492 37600 36548
rect 37520 36480 37600 36492
rect 37680 36868 37760 36880
rect 37680 36812 37692 36868
rect 37748 36812 37760 36868
rect 37680 36548 37760 36812
rect 37680 36492 37692 36548
rect 37748 36492 37760 36548
rect 37680 36480 37760 36492
rect 37840 36868 37920 36880
rect 37840 36812 37852 36868
rect 37908 36812 37920 36868
rect 37840 36548 37920 36812
rect 37840 36492 37852 36548
rect 37908 36492 37920 36548
rect 37840 36480 37920 36492
rect 38000 36868 38080 36880
rect 38000 36812 38012 36868
rect 38068 36812 38080 36868
rect 38000 36548 38080 36812
rect 38000 36492 38012 36548
rect 38068 36492 38080 36548
rect 38000 36480 38080 36492
rect 38160 36868 38240 36880
rect 38160 36812 38172 36868
rect 38228 36812 38240 36868
rect 38160 36548 38240 36812
rect 38160 36492 38172 36548
rect 38228 36492 38240 36548
rect 38160 36480 38240 36492
rect 38320 36868 38400 36880
rect 38320 36812 38332 36868
rect 38388 36812 38400 36868
rect 38320 36548 38400 36812
rect 38320 36492 38332 36548
rect 38388 36492 38400 36548
rect 38320 36480 38400 36492
rect 38480 36868 38560 36880
rect 38480 36812 38492 36868
rect 38548 36812 38560 36868
rect 38480 36548 38560 36812
rect 38480 36492 38492 36548
rect 38548 36492 38560 36548
rect 38480 36480 38560 36492
rect 38640 36868 38720 36880
rect 38640 36812 38652 36868
rect 38708 36812 38720 36868
rect 38640 36548 38720 36812
rect 38640 36492 38652 36548
rect 38708 36492 38720 36548
rect 38640 36480 38720 36492
rect 38800 36868 38880 36880
rect 38800 36812 38812 36868
rect 38868 36812 38880 36868
rect 38800 36548 38880 36812
rect 38800 36492 38812 36548
rect 38868 36492 38880 36548
rect 38800 36480 38880 36492
rect 38960 36868 39040 36880
rect 38960 36812 38972 36868
rect 39028 36812 39040 36868
rect 38960 36548 39040 36812
rect 38960 36492 38972 36548
rect 39028 36492 39040 36548
rect 38960 36480 39040 36492
rect 39120 36868 39200 36880
rect 39120 36812 39132 36868
rect 39188 36812 39200 36868
rect 39120 36548 39200 36812
rect 39120 36492 39132 36548
rect 39188 36492 39200 36548
rect 39120 36480 39200 36492
rect 39280 36868 39360 36880
rect 39280 36812 39292 36868
rect 39348 36812 39360 36868
rect 39280 36548 39360 36812
rect 39280 36492 39292 36548
rect 39348 36492 39360 36548
rect 39280 36480 39360 36492
rect 39440 36868 39520 36880
rect 39440 36812 39452 36868
rect 39508 36812 39520 36868
rect 39440 36548 39520 36812
rect 39440 36492 39452 36548
rect 39508 36492 39520 36548
rect 39440 36480 39520 36492
rect 39600 36868 39680 36880
rect 39600 36812 39612 36868
rect 39668 36812 39680 36868
rect 39600 36548 39680 36812
rect 39600 36492 39612 36548
rect 39668 36492 39680 36548
rect 39600 36480 39680 36492
rect 39760 36868 39840 36880
rect 39760 36812 39772 36868
rect 39828 36812 39840 36868
rect 39760 36548 39840 36812
rect 39760 36492 39772 36548
rect 39828 36492 39840 36548
rect 39760 36480 39840 36492
rect 39920 36868 40000 36880
rect 39920 36812 39932 36868
rect 39988 36812 40000 36868
rect 39920 36548 40000 36812
rect 39920 36492 39932 36548
rect 39988 36492 40000 36548
rect 39920 36480 40000 36492
rect 40080 36868 40160 36880
rect 40080 36812 40092 36868
rect 40148 36812 40160 36868
rect 40080 36548 40160 36812
rect 40080 36492 40092 36548
rect 40148 36492 40160 36548
rect 40080 36480 40160 36492
rect 40240 36868 40320 36880
rect 40240 36812 40252 36868
rect 40308 36812 40320 36868
rect 40240 36548 40320 36812
rect 40240 36492 40252 36548
rect 40308 36492 40320 36548
rect 40240 36480 40320 36492
rect 40400 36868 40480 36880
rect 40400 36812 40412 36868
rect 40468 36812 40480 36868
rect 40400 36548 40480 36812
rect 40400 36492 40412 36548
rect 40468 36492 40480 36548
rect 40400 36480 40480 36492
rect 40560 36868 40640 36880
rect 40560 36812 40572 36868
rect 40628 36812 40640 36868
rect 40560 36548 40640 36812
rect 40560 36492 40572 36548
rect 40628 36492 40640 36548
rect 40560 36480 40640 36492
rect 40720 36868 40800 36880
rect 40720 36812 40732 36868
rect 40788 36812 40800 36868
rect 40720 36548 40800 36812
rect 40720 36492 40732 36548
rect 40788 36492 40800 36548
rect 40720 36480 40800 36492
rect 40880 36868 40960 36880
rect 40880 36812 40892 36868
rect 40948 36812 40960 36868
rect 40880 36548 40960 36812
rect 40880 36492 40892 36548
rect 40948 36492 40960 36548
rect 40880 36480 40960 36492
rect 41040 36868 41120 36880
rect 41040 36812 41052 36868
rect 41108 36812 41120 36868
rect 41040 36548 41120 36812
rect 41040 36492 41052 36548
rect 41108 36492 41120 36548
rect 41040 36480 41120 36492
rect 41200 36868 41280 36880
rect 41200 36812 41212 36868
rect 41268 36812 41280 36868
rect 41200 36548 41280 36812
rect 41200 36492 41212 36548
rect 41268 36492 41280 36548
rect 41200 36480 41280 36492
rect 41360 36868 41440 36880
rect 41360 36812 41372 36868
rect 41428 36812 41440 36868
rect 41360 36548 41440 36812
rect 41360 36492 41372 36548
rect 41428 36492 41440 36548
rect 41360 36480 41440 36492
rect 41520 36868 41600 36880
rect 41520 36812 41532 36868
rect 41588 36812 41600 36868
rect 41520 36548 41600 36812
rect 41520 36492 41532 36548
rect 41588 36492 41600 36548
rect 41520 36480 41600 36492
rect 41680 36868 41760 36880
rect 41680 36812 41692 36868
rect 41748 36812 41760 36868
rect 41680 36548 41760 36812
rect 41680 36492 41692 36548
rect 41748 36492 41760 36548
rect 41680 36480 41760 36492
rect 41840 36868 41920 36880
rect 41840 36812 41852 36868
rect 41908 36812 41920 36868
rect 41840 36548 41920 36812
rect 41840 36492 41852 36548
rect 41908 36492 41920 36548
rect 41840 36480 41920 36492
rect 33520 36388 33600 36400
rect 33520 36332 33532 36388
rect 33588 36332 33600 36388
rect 33520 36068 33600 36332
rect 33520 36012 33532 36068
rect 33588 36012 33600 36068
rect 33520 35748 33600 36012
rect 33520 35692 33532 35748
rect 33588 35692 33600 35748
rect 33520 35428 33600 35692
rect 33520 35372 33532 35428
rect 33588 35372 33600 35428
rect 33520 35108 33600 35372
rect 33520 35052 33532 35108
rect 33588 35052 33600 35108
rect 33520 34788 33600 35052
rect 33520 34732 33532 34788
rect 33588 34732 33600 34788
rect 33520 34468 33600 34732
rect 33520 34412 33532 34468
rect 33588 34412 33600 34468
rect 33520 34400 33600 34412
rect 33680 36388 33760 36400
rect 33680 36332 33692 36388
rect 33748 36332 33760 36388
rect 33680 36068 33760 36332
rect 33680 36012 33692 36068
rect 33748 36012 33760 36068
rect 33680 35748 33760 36012
rect 33680 35692 33692 35748
rect 33748 35692 33760 35748
rect 33680 35428 33760 35692
rect 33680 35372 33692 35428
rect 33748 35372 33760 35428
rect 33680 35108 33760 35372
rect 33680 35052 33692 35108
rect 33748 35052 33760 35108
rect 33680 34788 33760 35052
rect 33680 34732 33692 34788
rect 33748 34732 33760 34788
rect 33680 34468 33760 34732
rect 33680 34412 33692 34468
rect 33748 34412 33760 34468
rect 33680 34400 33760 34412
rect 33840 36388 33920 36400
rect 33840 36332 33852 36388
rect 33908 36332 33920 36388
rect 33840 36068 33920 36332
rect 33840 36012 33852 36068
rect 33908 36012 33920 36068
rect 33840 35748 33920 36012
rect 33840 35692 33852 35748
rect 33908 35692 33920 35748
rect 33840 35428 33920 35692
rect 33840 35372 33852 35428
rect 33908 35372 33920 35428
rect 33840 35108 33920 35372
rect 33840 35052 33852 35108
rect 33908 35052 33920 35108
rect 33840 34788 33920 35052
rect 33840 34732 33852 34788
rect 33908 34732 33920 34788
rect 33840 34468 33920 34732
rect 33840 34412 33852 34468
rect 33908 34412 33920 34468
rect 33840 34400 33920 34412
rect 34000 36388 34080 36400
rect 34000 36332 34012 36388
rect 34068 36332 34080 36388
rect 34000 36068 34080 36332
rect 34000 36012 34012 36068
rect 34068 36012 34080 36068
rect 34000 35748 34080 36012
rect 34000 35692 34012 35748
rect 34068 35692 34080 35748
rect 34000 35428 34080 35692
rect 34000 35372 34012 35428
rect 34068 35372 34080 35428
rect 34000 35108 34080 35372
rect 34000 35052 34012 35108
rect 34068 35052 34080 35108
rect 34000 34788 34080 35052
rect 34000 34732 34012 34788
rect 34068 34732 34080 34788
rect 34000 34468 34080 34732
rect 34000 34412 34012 34468
rect 34068 34412 34080 34468
rect 34000 34400 34080 34412
rect 34160 36388 34240 36400
rect 34160 36332 34172 36388
rect 34228 36332 34240 36388
rect 34160 36068 34240 36332
rect 34160 36012 34172 36068
rect 34228 36012 34240 36068
rect 34160 35748 34240 36012
rect 34160 35692 34172 35748
rect 34228 35692 34240 35748
rect 34160 35428 34240 35692
rect 34160 35372 34172 35428
rect 34228 35372 34240 35428
rect 34160 35108 34240 35372
rect 34160 35052 34172 35108
rect 34228 35052 34240 35108
rect 34160 34788 34240 35052
rect 34160 34732 34172 34788
rect 34228 34732 34240 34788
rect 34160 34468 34240 34732
rect 34160 34412 34172 34468
rect 34228 34412 34240 34468
rect 34160 34400 34240 34412
rect 34320 36388 34400 36400
rect 34320 36332 34332 36388
rect 34388 36332 34400 36388
rect 34320 36068 34400 36332
rect 34320 36012 34332 36068
rect 34388 36012 34400 36068
rect 34320 35748 34400 36012
rect 34320 35692 34332 35748
rect 34388 35692 34400 35748
rect 34320 35428 34400 35692
rect 34320 35372 34332 35428
rect 34388 35372 34400 35428
rect 34320 35108 34400 35372
rect 34320 35052 34332 35108
rect 34388 35052 34400 35108
rect 34320 34788 34400 35052
rect 34320 34732 34332 34788
rect 34388 34732 34400 34788
rect 34320 34468 34400 34732
rect 34320 34412 34332 34468
rect 34388 34412 34400 34468
rect 34320 34400 34400 34412
rect 34480 36388 34560 36400
rect 34480 36332 34492 36388
rect 34548 36332 34560 36388
rect 34480 36068 34560 36332
rect 34480 36012 34492 36068
rect 34548 36012 34560 36068
rect 34480 35748 34560 36012
rect 34480 35692 34492 35748
rect 34548 35692 34560 35748
rect 34480 35428 34560 35692
rect 34480 35372 34492 35428
rect 34548 35372 34560 35428
rect 34480 35108 34560 35372
rect 34480 35052 34492 35108
rect 34548 35052 34560 35108
rect 34480 34788 34560 35052
rect 34480 34732 34492 34788
rect 34548 34732 34560 34788
rect 34480 34468 34560 34732
rect 34480 34412 34492 34468
rect 34548 34412 34560 34468
rect 34480 34400 34560 34412
rect 34640 36388 34720 36400
rect 34640 36332 34652 36388
rect 34708 36332 34720 36388
rect 34640 36068 34720 36332
rect 34640 36012 34652 36068
rect 34708 36012 34720 36068
rect 34640 35748 34720 36012
rect 34640 35692 34652 35748
rect 34708 35692 34720 35748
rect 34640 35428 34720 35692
rect 34640 35372 34652 35428
rect 34708 35372 34720 35428
rect 34640 35108 34720 35372
rect 34640 35052 34652 35108
rect 34708 35052 34720 35108
rect 34640 34788 34720 35052
rect 34640 34732 34652 34788
rect 34708 34732 34720 34788
rect 34640 34468 34720 34732
rect 34640 34412 34652 34468
rect 34708 34412 34720 34468
rect 34640 34400 34720 34412
rect 34800 36388 34880 36400
rect 34800 36332 34812 36388
rect 34868 36332 34880 36388
rect 34800 36068 34880 36332
rect 34800 36012 34812 36068
rect 34868 36012 34880 36068
rect 34800 35748 34880 36012
rect 34800 35692 34812 35748
rect 34868 35692 34880 35748
rect 34800 35428 34880 35692
rect 34800 35372 34812 35428
rect 34868 35372 34880 35428
rect 34800 35108 34880 35372
rect 34800 35052 34812 35108
rect 34868 35052 34880 35108
rect 34800 34788 34880 35052
rect 34800 34732 34812 34788
rect 34868 34732 34880 34788
rect 34800 34468 34880 34732
rect 34800 34412 34812 34468
rect 34868 34412 34880 34468
rect 34800 34400 34880 34412
rect 34960 36388 35040 36400
rect 34960 36332 34972 36388
rect 35028 36332 35040 36388
rect 34960 36068 35040 36332
rect 34960 36012 34972 36068
rect 35028 36012 35040 36068
rect 34960 35748 35040 36012
rect 34960 35692 34972 35748
rect 35028 35692 35040 35748
rect 34960 35428 35040 35692
rect 34960 35372 34972 35428
rect 35028 35372 35040 35428
rect 34960 35108 35040 35372
rect 34960 35052 34972 35108
rect 35028 35052 35040 35108
rect 34960 34788 35040 35052
rect 34960 34732 34972 34788
rect 35028 34732 35040 34788
rect 34960 34468 35040 34732
rect 34960 34412 34972 34468
rect 35028 34412 35040 34468
rect 34960 34400 35040 34412
rect 35120 36388 35200 36400
rect 35120 36332 35132 36388
rect 35188 36332 35200 36388
rect 35120 36068 35200 36332
rect 35120 36012 35132 36068
rect 35188 36012 35200 36068
rect 35120 35748 35200 36012
rect 35120 35692 35132 35748
rect 35188 35692 35200 35748
rect 35120 35428 35200 35692
rect 35120 35372 35132 35428
rect 35188 35372 35200 35428
rect 35120 35108 35200 35372
rect 35120 35052 35132 35108
rect 35188 35052 35200 35108
rect 35120 34788 35200 35052
rect 35120 34732 35132 34788
rect 35188 34732 35200 34788
rect 35120 34468 35200 34732
rect 35120 34412 35132 34468
rect 35188 34412 35200 34468
rect 35120 34400 35200 34412
rect 35280 36388 35360 36400
rect 35280 36332 35292 36388
rect 35348 36332 35360 36388
rect 35280 36068 35360 36332
rect 35280 36012 35292 36068
rect 35348 36012 35360 36068
rect 35280 35748 35360 36012
rect 35280 35692 35292 35748
rect 35348 35692 35360 35748
rect 35280 35428 35360 35692
rect 35280 35372 35292 35428
rect 35348 35372 35360 35428
rect 35280 35108 35360 35372
rect 35280 35052 35292 35108
rect 35348 35052 35360 35108
rect 35280 34788 35360 35052
rect 35280 34732 35292 34788
rect 35348 34732 35360 34788
rect 35280 34468 35360 34732
rect 35280 34412 35292 34468
rect 35348 34412 35360 34468
rect 35280 34400 35360 34412
rect 35440 36388 35520 36400
rect 35440 36332 35452 36388
rect 35508 36332 35520 36388
rect 35440 36068 35520 36332
rect 35440 36012 35452 36068
rect 35508 36012 35520 36068
rect 35440 35748 35520 36012
rect 35440 35692 35452 35748
rect 35508 35692 35520 35748
rect 35440 35428 35520 35692
rect 35440 35372 35452 35428
rect 35508 35372 35520 35428
rect 35440 35108 35520 35372
rect 35440 35052 35452 35108
rect 35508 35052 35520 35108
rect 35440 34788 35520 35052
rect 35440 34732 35452 34788
rect 35508 34732 35520 34788
rect 35440 34468 35520 34732
rect 35440 34412 35452 34468
rect 35508 34412 35520 34468
rect 35440 34400 35520 34412
rect 35600 36388 35680 36400
rect 35600 36332 35612 36388
rect 35668 36332 35680 36388
rect 35600 36068 35680 36332
rect 35600 36012 35612 36068
rect 35668 36012 35680 36068
rect 35600 35748 35680 36012
rect 35600 35692 35612 35748
rect 35668 35692 35680 35748
rect 35600 35428 35680 35692
rect 35600 35372 35612 35428
rect 35668 35372 35680 35428
rect 35600 35108 35680 35372
rect 35600 35052 35612 35108
rect 35668 35052 35680 35108
rect 35600 34788 35680 35052
rect 35600 34732 35612 34788
rect 35668 34732 35680 34788
rect 35600 34468 35680 34732
rect 35600 34412 35612 34468
rect 35668 34412 35680 34468
rect 35600 34400 35680 34412
rect 35760 36388 35840 36400
rect 35760 36332 35772 36388
rect 35828 36332 35840 36388
rect 35760 36068 35840 36332
rect 35760 36012 35772 36068
rect 35828 36012 35840 36068
rect 35760 35748 35840 36012
rect 35760 35692 35772 35748
rect 35828 35692 35840 35748
rect 35760 35428 35840 35692
rect 35760 35372 35772 35428
rect 35828 35372 35840 35428
rect 35760 35108 35840 35372
rect 35760 35052 35772 35108
rect 35828 35052 35840 35108
rect 35760 34788 35840 35052
rect 35760 34732 35772 34788
rect 35828 34732 35840 34788
rect 35760 34468 35840 34732
rect 35760 34412 35772 34468
rect 35828 34412 35840 34468
rect 35760 34400 35840 34412
rect 35920 36388 36000 36400
rect 35920 36332 35932 36388
rect 35988 36332 36000 36388
rect 35920 36068 36000 36332
rect 35920 36012 35932 36068
rect 35988 36012 36000 36068
rect 35920 35748 36000 36012
rect 35920 35692 35932 35748
rect 35988 35692 36000 35748
rect 35920 35428 36000 35692
rect 35920 35372 35932 35428
rect 35988 35372 36000 35428
rect 35920 35108 36000 35372
rect 35920 35052 35932 35108
rect 35988 35052 36000 35108
rect 35920 34788 36000 35052
rect 35920 34732 35932 34788
rect 35988 34732 36000 34788
rect 35920 34468 36000 34732
rect 35920 34412 35932 34468
rect 35988 34412 36000 34468
rect 35920 34400 36000 34412
rect 36080 36388 36160 36400
rect 36080 36332 36092 36388
rect 36148 36332 36160 36388
rect 36080 36068 36160 36332
rect 36080 36012 36092 36068
rect 36148 36012 36160 36068
rect 36080 35748 36160 36012
rect 36080 35692 36092 35748
rect 36148 35692 36160 35748
rect 36080 35428 36160 35692
rect 36080 35372 36092 35428
rect 36148 35372 36160 35428
rect 36080 35108 36160 35372
rect 36080 35052 36092 35108
rect 36148 35052 36160 35108
rect 36080 34788 36160 35052
rect 36080 34732 36092 34788
rect 36148 34732 36160 34788
rect 36080 34468 36160 34732
rect 36080 34412 36092 34468
rect 36148 34412 36160 34468
rect 36080 34400 36160 34412
rect 36240 36388 36320 36400
rect 36240 36332 36252 36388
rect 36308 36332 36320 36388
rect 36240 36068 36320 36332
rect 36240 36012 36252 36068
rect 36308 36012 36320 36068
rect 36240 35748 36320 36012
rect 36240 35692 36252 35748
rect 36308 35692 36320 35748
rect 36240 35428 36320 35692
rect 36240 35372 36252 35428
rect 36308 35372 36320 35428
rect 36240 35108 36320 35372
rect 36240 35052 36252 35108
rect 36308 35052 36320 35108
rect 36240 34788 36320 35052
rect 36240 34732 36252 34788
rect 36308 34732 36320 34788
rect 36240 34468 36320 34732
rect 36240 34412 36252 34468
rect 36308 34412 36320 34468
rect 36240 34400 36320 34412
rect 36400 36388 36480 36400
rect 36400 36332 36412 36388
rect 36468 36332 36480 36388
rect 36400 36068 36480 36332
rect 36400 36012 36412 36068
rect 36468 36012 36480 36068
rect 36400 35748 36480 36012
rect 36400 35692 36412 35748
rect 36468 35692 36480 35748
rect 36400 35428 36480 35692
rect 36400 35372 36412 35428
rect 36468 35372 36480 35428
rect 36400 35108 36480 35372
rect 36400 35052 36412 35108
rect 36468 35052 36480 35108
rect 36400 34788 36480 35052
rect 36400 34732 36412 34788
rect 36468 34732 36480 34788
rect 36400 34468 36480 34732
rect 36400 34412 36412 34468
rect 36468 34412 36480 34468
rect 36400 34400 36480 34412
rect 36560 36388 36640 36400
rect 36560 36332 36572 36388
rect 36628 36332 36640 36388
rect 36560 36068 36640 36332
rect 36560 36012 36572 36068
rect 36628 36012 36640 36068
rect 36560 35748 36640 36012
rect 36560 35692 36572 35748
rect 36628 35692 36640 35748
rect 36560 35428 36640 35692
rect 36560 35372 36572 35428
rect 36628 35372 36640 35428
rect 36560 35108 36640 35372
rect 36560 35052 36572 35108
rect 36628 35052 36640 35108
rect 36560 34788 36640 35052
rect 36560 34732 36572 34788
rect 36628 34732 36640 34788
rect 36560 34468 36640 34732
rect 36560 34412 36572 34468
rect 36628 34412 36640 34468
rect 36560 34400 36640 34412
rect 36720 36388 36800 36400
rect 36720 36332 36732 36388
rect 36788 36332 36800 36388
rect 36720 36068 36800 36332
rect 36720 36012 36732 36068
rect 36788 36012 36800 36068
rect 36720 35748 36800 36012
rect 36720 35692 36732 35748
rect 36788 35692 36800 35748
rect 36720 35428 36800 35692
rect 36720 35372 36732 35428
rect 36788 35372 36800 35428
rect 36720 35108 36800 35372
rect 36720 35052 36732 35108
rect 36788 35052 36800 35108
rect 36720 34788 36800 35052
rect 36720 34732 36732 34788
rect 36788 34732 36800 34788
rect 36720 34468 36800 34732
rect 36720 34412 36732 34468
rect 36788 34412 36800 34468
rect 36720 34400 36800 34412
rect 36880 36388 36960 36400
rect 36880 36332 36892 36388
rect 36948 36332 36960 36388
rect 36880 36068 36960 36332
rect 36880 36012 36892 36068
rect 36948 36012 36960 36068
rect 36880 35748 36960 36012
rect 36880 35692 36892 35748
rect 36948 35692 36960 35748
rect 36880 35428 36960 35692
rect 36880 35372 36892 35428
rect 36948 35372 36960 35428
rect 36880 35108 36960 35372
rect 36880 35052 36892 35108
rect 36948 35052 36960 35108
rect 36880 34788 36960 35052
rect 36880 34732 36892 34788
rect 36948 34732 36960 34788
rect 36880 34468 36960 34732
rect 36880 34412 36892 34468
rect 36948 34412 36960 34468
rect 36880 34400 36960 34412
rect 37040 36388 37120 36400
rect 37040 36332 37052 36388
rect 37108 36332 37120 36388
rect 37040 36068 37120 36332
rect 37040 36012 37052 36068
rect 37108 36012 37120 36068
rect 37040 35748 37120 36012
rect 37040 35692 37052 35748
rect 37108 35692 37120 35748
rect 37040 35428 37120 35692
rect 37040 35372 37052 35428
rect 37108 35372 37120 35428
rect 37040 35108 37120 35372
rect 37040 35052 37052 35108
rect 37108 35052 37120 35108
rect 37040 34788 37120 35052
rect 37040 34732 37052 34788
rect 37108 34732 37120 34788
rect 37040 34468 37120 34732
rect 37040 34412 37052 34468
rect 37108 34412 37120 34468
rect 37040 34400 37120 34412
rect 37200 36388 37280 36400
rect 37200 36332 37212 36388
rect 37268 36332 37280 36388
rect 37200 36068 37280 36332
rect 37200 36012 37212 36068
rect 37268 36012 37280 36068
rect 37200 35748 37280 36012
rect 37200 35692 37212 35748
rect 37268 35692 37280 35748
rect 37200 35428 37280 35692
rect 37200 35372 37212 35428
rect 37268 35372 37280 35428
rect 37200 35108 37280 35372
rect 37200 35052 37212 35108
rect 37268 35052 37280 35108
rect 37200 34788 37280 35052
rect 37200 34732 37212 34788
rect 37268 34732 37280 34788
rect 37200 34468 37280 34732
rect 37200 34412 37212 34468
rect 37268 34412 37280 34468
rect 37200 34400 37280 34412
rect 37360 36388 37440 36400
rect 37360 36332 37372 36388
rect 37428 36332 37440 36388
rect 37360 36068 37440 36332
rect 37360 36012 37372 36068
rect 37428 36012 37440 36068
rect 37360 35748 37440 36012
rect 37360 35692 37372 35748
rect 37428 35692 37440 35748
rect 37360 35428 37440 35692
rect 37360 35372 37372 35428
rect 37428 35372 37440 35428
rect 37360 35108 37440 35372
rect 37360 35052 37372 35108
rect 37428 35052 37440 35108
rect 37360 34788 37440 35052
rect 37360 34732 37372 34788
rect 37428 34732 37440 34788
rect 37360 34468 37440 34732
rect 37360 34412 37372 34468
rect 37428 34412 37440 34468
rect 37360 34400 37440 34412
rect 37520 36388 37600 36400
rect 37520 36332 37532 36388
rect 37588 36332 37600 36388
rect 37520 36068 37600 36332
rect 37520 36012 37532 36068
rect 37588 36012 37600 36068
rect 37520 35748 37600 36012
rect 37520 35692 37532 35748
rect 37588 35692 37600 35748
rect 37520 35428 37600 35692
rect 37520 35372 37532 35428
rect 37588 35372 37600 35428
rect 37520 35108 37600 35372
rect 37520 35052 37532 35108
rect 37588 35052 37600 35108
rect 37520 34788 37600 35052
rect 37520 34732 37532 34788
rect 37588 34732 37600 34788
rect 37520 34468 37600 34732
rect 37520 34412 37532 34468
rect 37588 34412 37600 34468
rect 37520 34400 37600 34412
rect 37680 36388 37760 36400
rect 37680 36332 37692 36388
rect 37748 36332 37760 36388
rect 37680 36068 37760 36332
rect 37680 36012 37692 36068
rect 37748 36012 37760 36068
rect 37680 35748 37760 36012
rect 37680 35692 37692 35748
rect 37748 35692 37760 35748
rect 37680 35428 37760 35692
rect 37680 35372 37692 35428
rect 37748 35372 37760 35428
rect 37680 35108 37760 35372
rect 37680 35052 37692 35108
rect 37748 35052 37760 35108
rect 37680 34788 37760 35052
rect 37680 34732 37692 34788
rect 37748 34732 37760 34788
rect 37680 34468 37760 34732
rect 37680 34412 37692 34468
rect 37748 34412 37760 34468
rect 37680 34400 37760 34412
rect 37840 36388 37920 36400
rect 37840 36332 37852 36388
rect 37908 36332 37920 36388
rect 37840 36068 37920 36332
rect 37840 36012 37852 36068
rect 37908 36012 37920 36068
rect 37840 35748 37920 36012
rect 37840 35692 37852 35748
rect 37908 35692 37920 35748
rect 37840 35428 37920 35692
rect 37840 35372 37852 35428
rect 37908 35372 37920 35428
rect 37840 35108 37920 35372
rect 37840 35052 37852 35108
rect 37908 35052 37920 35108
rect 37840 34788 37920 35052
rect 37840 34732 37852 34788
rect 37908 34732 37920 34788
rect 37840 34468 37920 34732
rect 37840 34412 37852 34468
rect 37908 34412 37920 34468
rect 37840 34400 37920 34412
rect 38000 36388 38080 36400
rect 38000 36332 38012 36388
rect 38068 36332 38080 36388
rect 38000 36068 38080 36332
rect 38000 36012 38012 36068
rect 38068 36012 38080 36068
rect 38000 35748 38080 36012
rect 38000 35692 38012 35748
rect 38068 35692 38080 35748
rect 38000 35428 38080 35692
rect 38000 35372 38012 35428
rect 38068 35372 38080 35428
rect 38000 35108 38080 35372
rect 38000 35052 38012 35108
rect 38068 35052 38080 35108
rect 38000 34788 38080 35052
rect 38000 34732 38012 34788
rect 38068 34732 38080 34788
rect 38000 34468 38080 34732
rect 38000 34412 38012 34468
rect 38068 34412 38080 34468
rect 38000 34400 38080 34412
rect 38160 36388 38240 36400
rect 38160 36332 38172 36388
rect 38228 36332 38240 36388
rect 38160 36068 38240 36332
rect 38160 36012 38172 36068
rect 38228 36012 38240 36068
rect 38160 35748 38240 36012
rect 38160 35692 38172 35748
rect 38228 35692 38240 35748
rect 38160 35428 38240 35692
rect 38160 35372 38172 35428
rect 38228 35372 38240 35428
rect 38160 35108 38240 35372
rect 38160 35052 38172 35108
rect 38228 35052 38240 35108
rect 38160 34788 38240 35052
rect 38160 34732 38172 34788
rect 38228 34732 38240 34788
rect 38160 34468 38240 34732
rect 38160 34412 38172 34468
rect 38228 34412 38240 34468
rect 38160 34400 38240 34412
rect 38320 36388 38400 36400
rect 38320 36332 38332 36388
rect 38388 36332 38400 36388
rect 38320 36068 38400 36332
rect 38320 36012 38332 36068
rect 38388 36012 38400 36068
rect 38320 35748 38400 36012
rect 38320 35692 38332 35748
rect 38388 35692 38400 35748
rect 38320 35428 38400 35692
rect 38320 35372 38332 35428
rect 38388 35372 38400 35428
rect 38320 35108 38400 35372
rect 38320 35052 38332 35108
rect 38388 35052 38400 35108
rect 38320 34788 38400 35052
rect 38320 34732 38332 34788
rect 38388 34732 38400 34788
rect 38320 34468 38400 34732
rect 38320 34412 38332 34468
rect 38388 34412 38400 34468
rect 38320 34400 38400 34412
rect 38480 36388 38560 36400
rect 38480 36332 38492 36388
rect 38548 36332 38560 36388
rect 38480 36068 38560 36332
rect 38480 36012 38492 36068
rect 38548 36012 38560 36068
rect 38480 35748 38560 36012
rect 38480 35692 38492 35748
rect 38548 35692 38560 35748
rect 38480 35428 38560 35692
rect 38480 35372 38492 35428
rect 38548 35372 38560 35428
rect 38480 35108 38560 35372
rect 38480 35052 38492 35108
rect 38548 35052 38560 35108
rect 38480 34788 38560 35052
rect 38480 34732 38492 34788
rect 38548 34732 38560 34788
rect 38480 34468 38560 34732
rect 38480 34412 38492 34468
rect 38548 34412 38560 34468
rect 38480 34400 38560 34412
rect 38640 36388 38720 36400
rect 38640 36332 38652 36388
rect 38708 36332 38720 36388
rect 38640 36068 38720 36332
rect 38640 36012 38652 36068
rect 38708 36012 38720 36068
rect 38640 35748 38720 36012
rect 38640 35692 38652 35748
rect 38708 35692 38720 35748
rect 38640 35428 38720 35692
rect 38640 35372 38652 35428
rect 38708 35372 38720 35428
rect 38640 35108 38720 35372
rect 38640 35052 38652 35108
rect 38708 35052 38720 35108
rect 38640 34788 38720 35052
rect 38640 34732 38652 34788
rect 38708 34732 38720 34788
rect 38640 34468 38720 34732
rect 38640 34412 38652 34468
rect 38708 34412 38720 34468
rect 38640 34400 38720 34412
rect 38800 36388 38880 36400
rect 38800 36332 38812 36388
rect 38868 36332 38880 36388
rect 38800 36068 38880 36332
rect 38800 36012 38812 36068
rect 38868 36012 38880 36068
rect 38800 35748 38880 36012
rect 38800 35692 38812 35748
rect 38868 35692 38880 35748
rect 38800 35428 38880 35692
rect 38800 35372 38812 35428
rect 38868 35372 38880 35428
rect 38800 35108 38880 35372
rect 38800 35052 38812 35108
rect 38868 35052 38880 35108
rect 38800 34788 38880 35052
rect 38800 34732 38812 34788
rect 38868 34732 38880 34788
rect 38800 34468 38880 34732
rect 38800 34412 38812 34468
rect 38868 34412 38880 34468
rect 38800 34400 38880 34412
rect 38960 36388 39040 36400
rect 38960 36332 38972 36388
rect 39028 36332 39040 36388
rect 38960 36068 39040 36332
rect 38960 36012 38972 36068
rect 39028 36012 39040 36068
rect 38960 35748 39040 36012
rect 38960 35692 38972 35748
rect 39028 35692 39040 35748
rect 38960 35428 39040 35692
rect 38960 35372 38972 35428
rect 39028 35372 39040 35428
rect 38960 35108 39040 35372
rect 38960 35052 38972 35108
rect 39028 35052 39040 35108
rect 38960 34788 39040 35052
rect 38960 34732 38972 34788
rect 39028 34732 39040 34788
rect 38960 34468 39040 34732
rect 38960 34412 38972 34468
rect 39028 34412 39040 34468
rect 38960 34400 39040 34412
rect 39120 36388 39200 36400
rect 39120 36332 39132 36388
rect 39188 36332 39200 36388
rect 39120 36068 39200 36332
rect 39120 36012 39132 36068
rect 39188 36012 39200 36068
rect 39120 35748 39200 36012
rect 39120 35692 39132 35748
rect 39188 35692 39200 35748
rect 39120 35428 39200 35692
rect 39120 35372 39132 35428
rect 39188 35372 39200 35428
rect 39120 35108 39200 35372
rect 39120 35052 39132 35108
rect 39188 35052 39200 35108
rect 39120 34788 39200 35052
rect 39120 34732 39132 34788
rect 39188 34732 39200 34788
rect 39120 34468 39200 34732
rect 39120 34412 39132 34468
rect 39188 34412 39200 34468
rect 39120 34400 39200 34412
rect 39280 36388 39360 36400
rect 39280 36332 39292 36388
rect 39348 36332 39360 36388
rect 39280 36068 39360 36332
rect 39280 36012 39292 36068
rect 39348 36012 39360 36068
rect 39280 35748 39360 36012
rect 39280 35692 39292 35748
rect 39348 35692 39360 35748
rect 39280 35428 39360 35692
rect 39280 35372 39292 35428
rect 39348 35372 39360 35428
rect 39280 35108 39360 35372
rect 39280 35052 39292 35108
rect 39348 35052 39360 35108
rect 39280 34788 39360 35052
rect 39280 34732 39292 34788
rect 39348 34732 39360 34788
rect 39280 34468 39360 34732
rect 39280 34412 39292 34468
rect 39348 34412 39360 34468
rect 39280 34400 39360 34412
rect 39440 36388 39520 36400
rect 39440 36332 39452 36388
rect 39508 36332 39520 36388
rect 39440 36068 39520 36332
rect 39440 36012 39452 36068
rect 39508 36012 39520 36068
rect 39440 35748 39520 36012
rect 39440 35692 39452 35748
rect 39508 35692 39520 35748
rect 39440 35428 39520 35692
rect 39440 35372 39452 35428
rect 39508 35372 39520 35428
rect 39440 35108 39520 35372
rect 39440 35052 39452 35108
rect 39508 35052 39520 35108
rect 39440 34788 39520 35052
rect 39440 34732 39452 34788
rect 39508 34732 39520 34788
rect 39440 34468 39520 34732
rect 39440 34412 39452 34468
rect 39508 34412 39520 34468
rect 39440 34400 39520 34412
rect 39600 36388 39680 36400
rect 39600 36332 39612 36388
rect 39668 36332 39680 36388
rect 39600 36068 39680 36332
rect 39600 36012 39612 36068
rect 39668 36012 39680 36068
rect 39600 35748 39680 36012
rect 39600 35692 39612 35748
rect 39668 35692 39680 35748
rect 39600 35428 39680 35692
rect 39600 35372 39612 35428
rect 39668 35372 39680 35428
rect 39600 35108 39680 35372
rect 39600 35052 39612 35108
rect 39668 35052 39680 35108
rect 39600 34788 39680 35052
rect 39600 34732 39612 34788
rect 39668 34732 39680 34788
rect 39600 34468 39680 34732
rect 39600 34412 39612 34468
rect 39668 34412 39680 34468
rect 39600 34400 39680 34412
rect 39760 36388 39840 36400
rect 39760 36332 39772 36388
rect 39828 36332 39840 36388
rect 39760 36068 39840 36332
rect 39760 36012 39772 36068
rect 39828 36012 39840 36068
rect 39760 35748 39840 36012
rect 39760 35692 39772 35748
rect 39828 35692 39840 35748
rect 39760 35428 39840 35692
rect 39760 35372 39772 35428
rect 39828 35372 39840 35428
rect 39760 35108 39840 35372
rect 39760 35052 39772 35108
rect 39828 35052 39840 35108
rect 39760 34788 39840 35052
rect 39760 34732 39772 34788
rect 39828 34732 39840 34788
rect 39760 34468 39840 34732
rect 39760 34412 39772 34468
rect 39828 34412 39840 34468
rect 39760 34400 39840 34412
rect 39920 36388 40000 36400
rect 39920 36332 39932 36388
rect 39988 36332 40000 36388
rect 39920 36068 40000 36332
rect 39920 36012 39932 36068
rect 39988 36012 40000 36068
rect 39920 35748 40000 36012
rect 39920 35692 39932 35748
rect 39988 35692 40000 35748
rect 39920 35428 40000 35692
rect 39920 35372 39932 35428
rect 39988 35372 40000 35428
rect 39920 35108 40000 35372
rect 39920 35052 39932 35108
rect 39988 35052 40000 35108
rect 39920 34788 40000 35052
rect 39920 34732 39932 34788
rect 39988 34732 40000 34788
rect 39920 34468 40000 34732
rect 39920 34412 39932 34468
rect 39988 34412 40000 34468
rect 39920 34400 40000 34412
rect 40080 36388 40160 36400
rect 40080 36332 40092 36388
rect 40148 36332 40160 36388
rect 40080 36068 40160 36332
rect 40080 36012 40092 36068
rect 40148 36012 40160 36068
rect 40080 35748 40160 36012
rect 40080 35692 40092 35748
rect 40148 35692 40160 35748
rect 40080 35428 40160 35692
rect 40080 35372 40092 35428
rect 40148 35372 40160 35428
rect 40080 35108 40160 35372
rect 40080 35052 40092 35108
rect 40148 35052 40160 35108
rect 40080 34788 40160 35052
rect 40080 34732 40092 34788
rect 40148 34732 40160 34788
rect 40080 34468 40160 34732
rect 40080 34412 40092 34468
rect 40148 34412 40160 34468
rect 40080 34400 40160 34412
rect 40240 36388 40320 36400
rect 40240 36332 40252 36388
rect 40308 36332 40320 36388
rect 40240 36068 40320 36332
rect 40240 36012 40252 36068
rect 40308 36012 40320 36068
rect 40240 35748 40320 36012
rect 40240 35692 40252 35748
rect 40308 35692 40320 35748
rect 40240 35428 40320 35692
rect 40240 35372 40252 35428
rect 40308 35372 40320 35428
rect 40240 35108 40320 35372
rect 40240 35052 40252 35108
rect 40308 35052 40320 35108
rect 40240 34788 40320 35052
rect 40240 34732 40252 34788
rect 40308 34732 40320 34788
rect 40240 34468 40320 34732
rect 40240 34412 40252 34468
rect 40308 34412 40320 34468
rect 40240 34400 40320 34412
rect 40400 36388 40480 36400
rect 40400 36332 40412 36388
rect 40468 36332 40480 36388
rect 40400 36068 40480 36332
rect 40400 36012 40412 36068
rect 40468 36012 40480 36068
rect 40400 35748 40480 36012
rect 40400 35692 40412 35748
rect 40468 35692 40480 35748
rect 40400 35428 40480 35692
rect 40400 35372 40412 35428
rect 40468 35372 40480 35428
rect 40400 35108 40480 35372
rect 40400 35052 40412 35108
rect 40468 35052 40480 35108
rect 40400 34788 40480 35052
rect 40400 34732 40412 34788
rect 40468 34732 40480 34788
rect 40400 34468 40480 34732
rect 40400 34412 40412 34468
rect 40468 34412 40480 34468
rect 40400 34400 40480 34412
rect 40560 36388 40640 36400
rect 40560 36332 40572 36388
rect 40628 36332 40640 36388
rect 40560 36068 40640 36332
rect 40560 36012 40572 36068
rect 40628 36012 40640 36068
rect 40560 35748 40640 36012
rect 40560 35692 40572 35748
rect 40628 35692 40640 35748
rect 40560 35428 40640 35692
rect 40560 35372 40572 35428
rect 40628 35372 40640 35428
rect 40560 35108 40640 35372
rect 40560 35052 40572 35108
rect 40628 35052 40640 35108
rect 40560 34788 40640 35052
rect 40560 34732 40572 34788
rect 40628 34732 40640 34788
rect 40560 34468 40640 34732
rect 40560 34412 40572 34468
rect 40628 34412 40640 34468
rect 40560 34400 40640 34412
rect 40720 36388 40800 36400
rect 40720 36332 40732 36388
rect 40788 36332 40800 36388
rect 40720 36068 40800 36332
rect 40720 36012 40732 36068
rect 40788 36012 40800 36068
rect 40720 35748 40800 36012
rect 40720 35692 40732 35748
rect 40788 35692 40800 35748
rect 40720 35428 40800 35692
rect 40720 35372 40732 35428
rect 40788 35372 40800 35428
rect 40720 35108 40800 35372
rect 40720 35052 40732 35108
rect 40788 35052 40800 35108
rect 40720 34788 40800 35052
rect 40720 34732 40732 34788
rect 40788 34732 40800 34788
rect 40720 34468 40800 34732
rect 40720 34412 40732 34468
rect 40788 34412 40800 34468
rect 40720 34400 40800 34412
rect 40880 36388 40960 36400
rect 40880 36332 40892 36388
rect 40948 36332 40960 36388
rect 40880 36068 40960 36332
rect 40880 36012 40892 36068
rect 40948 36012 40960 36068
rect 40880 35748 40960 36012
rect 40880 35692 40892 35748
rect 40948 35692 40960 35748
rect 40880 35428 40960 35692
rect 40880 35372 40892 35428
rect 40948 35372 40960 35428
rect 40880 35108 40960 35372
rect 40880 35052 40892 35108
rect 40948 35052 40960 35108
rect 40880 34788 40960 35052
rect 40880 34732 40892 34788
rect 40948 34732 40960 34788
rect 40880 34468 40960 34732
rect 40880 34412 40892 34468
rect 40948 34412 40960 34468
rect 40880 34400 40960 34412
rect 41040 36388 41120 36400
rect 41040 36332 41052 36388
rect 41108 36332 41120 36388
rect 41040 36068 41120 36332
rect 41040 36012 41052 36068
rect 41108 36012 41120 36068
rect 41040 35748 41120 36012
rect 41040 35692 41052 35748
rect 41108 35692 41120 35748
rect 41040 35428 41120 35692
rect 41040 35372 41052 35428
rect 41108 35372 41120 35428
rect 41040 35108 41120 35372
rect 41040 35052 41052 35108
rect 41108 35052 41120 35108
rect 41040 34788 41120 35052
rect 41040 34732 41052 34788
rect 41108 34732 41120 34788
rect 41040 34468 41120 34732
rect 41040 34412 41052 34468
rect 41108 34412 41120 34468
rect 41040 34400 41120 34412
rect 41200 36388 41280 36400
rect 41200 36332 41212 36388
rect 41268 36332 41280 36388
rect 41200 36068 41280 36332
rect 41200 36012 41212 36068
rect 41268 36012 41280 36068
rect 41200 35748 41280 36012
rect 41200 35692 41212 35748
rect 41268 35692 41280 35748
rect 41200 35428 41280 35692
rect 41200 35372 41212 35428
rect 41268 35372 41280 35428
rect 41200 35108 41280 35372
rect 41200 35052 41212 35108
rect 41268 35052 41280 35108
rect 41200 34788 41280 35052
rect 41200 34732 41212 34788
rect 41268 34732 41280 34788
rect 41200 34468 41280 34732
rect 41200 34412 41212 34468
rect 41268 34412 41280 34468
rect 41200 34400 41280 34412
rect 41360 36388 41440 36400
rect 41360 36332 41372 36388
rect 41428 36332 41440 36388
rect 41360 36068 41440 36332
rect 41360 36012 41372 36068
rect 41428 36012 41440 36068
rect 41360 35748 41440 36012
rect 41360 35692 41372 35748
rect 41428 35692 41440 35748
rect 41360 35428 41440 35692
rect 41360 35372 41372 35428
rect 41428 35372 41440 35428
rect 41360 35108 41440 35372
rect 41360 35052 41372 35108
rect 41428 35052 41440 35108
rect 41360 34788 41440 35052
rect 41360 34732 41372 34788
rect 41428 34732 41440 34788
rect 41360 34468 41440 34732
rect 41360 34412 41372 34468
rect 41428 34412 41440 34468
rect 41360 34400 41440 34412
rect 41520 36388 41600 36400
rect 41520 36332 41532 36388
rect 41588 36332 41600 36388
rect 41520 36068 41600 36332
rect 41520 36012 41532 36068
rect 41588 36012 41600 36068
rect 41520 35748 41600 36012
rect 41520 35692 41532 35748
rect 41588 35692 41600 35748
rect 41520 35428 41600 35692
rect 41520 35372 41532 35428
rect 41588 35372 41600 35428
rect 41520 35108 41600 35372
rect 41520 35052 41532 35108
rect 41588 35052 41600 35108
rect 41520 34788 41600 35052
rect 41520 34732 41532 34788
rect 41588 34732 41600 34788
rect 41520 34468 41600 34732
rect 41520 34412 41532 34468
rect 41588 34412 41600 34468
rect 41520 34400 41600 34412
rect 41680 36388 41760 36400
rect 41680 36332 41692 36388
rect 41748 36332 41760 36388
rect 41680 36068 41760 36332
rect 41680 36012 41692 36068
rect 41748 36012 41760 36068
rect 41680 35748 41760 36012
rect 41680 35692 41692 35748
rect 41748 35692 41760 35748
rect 41680 35428 41760 35692
rect 41680 35372 41692 35428
rect 41748 35372 41760 35428
rect 41680 35108 41760 35372
rect 41680 35052 41692 35108
rect 41748 35052 41760 35108
rect 41680 34788 41760 35052
rect 41680 34732 41692 34788
rect 41748 34732 41760 34788
rect 41680 34468 41760 34732
rect 41680 34412 41692 34468
rect 41748 34412 41760 34468
rect 41680 34400 41760 34412
rect 41840 36388 41920 36400
rect 41840 36332 41852 36388
rect 41908 36332 41920 36388
rect 41840 36068 41920 36332
rect 41840 36012 41852 36068
rect 41908 36012 41920 36068
rect 41840 35748 41920 36012
rect 41840 35692 41852 35748
rect 41908 35692 41920 35748
rect 41840 35428 41920 35692
rect 41840 35372 41852 35428
rect 41908 35372 41920 35428
rect 41840 35108 41920 35372
rect 41840 35052 41852 35108
rect 41908 35052 41920 35108
rect 41840 34788 41920 35052
rect 41840 34732 41852 34788
rect 41908 34732 41920 34788
rect 41840 34468 41920 34732
rect 41840 34412 41852 34468
rect 41908 34412 41920 34468
rect 41840 34400 41920 34412
rect 33520 34308 33600 34320
rect 33520 34252 33532 34308
rect 33588 34252 33600 34308
rect 33520 33988 33600 34252
rect 33520 33932 33532 33988
rect 33588 33932 33600 33988
rect 33520 33920 33600 33932
rect 33680 34308 33760 34320
rect 33680 34252 33692 34308
rect 33748 34252 33760 34308
rect 33680 33988 33760 34252
rect 33680 33932 33692 33988
rect 33748 33932 33760 33988
rect 33680 33920 33760 33932
rect 33840 34308 33920 34320
rect 33840 34252 33852 34308
rect 33908 34252 33920 34308
rect 33840 33988 33920 34252
rect 33840 33932 33852 33988
rect 33908 33932 33920 33988
rect 33840 33920 33920 33932
rect 34000 34308 34080 34320
rect 34000 34252 34012 34308
rect 34068 34252 34080 34308
rect 34000 33988 34080 34252
rect 34000 33932 34012 33988
rect 34068 33932 34080 33988
rect 34000 33920 34080 33932
rect 34160 34308 34240 34320
rect 34160 34252 34172 34308
rect 34228 34252 34240 34308
rect 34160 33988 34240 34252
rect 34160 33932 34172 33988
rect 34228 33932 34240 33988
rect 34160 33920 34240 33932
rect 34320 34308 34400 34320
rect 34320 34252 34332 34308
rect 34388 34252 34400 34308
rect 34320 33988 34400 34252
rect 34320 33932 34332 33988
rect 34388 33932 34400 33988
rect 34320 33920 34400 33932
rect 34480 34308 34560 34320
rect 34480 34252 34492 34308
rect 34548 34252 34560 34308
rect 34480 33988 34560 34252
rect 34480 33932 34492 33988
rect 34548 33932 34560 33988
rect 34480 33920 34560 33932
rect 34640 34308 34720 34320
rect 34640 34252 34652 34308
rect 34708 34252 34720 34308
rect 34640 33988 34720 34252
rect 34640 33932 34652 33988
rect 34708 33932 34720 33988
rect 34640 33920 34720 33932
rect 34800 34308 34880 34320
rect 34800 34252 34812 34308
rect 34868 34252 34880 34308
rect 34800 33988 34880 34252
rect 34800 33932 34812 33988
rect 34868 33932 34880 33988
rect 34800 33920 34880 33932
rect 34960 34308 35040 34320
rect 34960 34252 34972 34308
rect 35028 34252 35040 34308
rect 34960 33988 35040 34252
rect 34960 33932 34972 33988
rect 35028 33932 35040 33988
rect 34960 33920 35040 33932
rect 35120 34308 35200 34320
rect 35120 34252 35132 34308
rect 35188 34252 35200 34308
rect 35120 33988 35200 34252
rect 35120 33932 35132 33988
rect 35188 33932 35200 33988
rect 35120 33920 35200 33932
rect 35280 34308 35360 34320
rect 35280 34252 35292 34308
rect 35348 34252 35360 34308
rect 35280 33988 35360 34252
rect 35280 33932 35292 33988
rect 35348 33932 35360 33988
rect 35280 33920 35360 33932
rect 35440 34308 35520 34320
rect 35440 34252 35452 34308
rect 35508 34252 35520 34308
rect 35440 33988 35520 34252
rect 35440 33932 35452 33988
rect 35508 33932 35520 33988
rect 35440 33920 35520 33932
rect 35600 34308 35680 34320
rect 35600 34252 35612 34308
rect 35668 34252 35680 34308
rect 35600 33988 35680 34252
rect 35600 33932 35612 33988
rect 35668 33932 35680 33988
rect 35600 33920 35680 33932
rect 35760 34308 35840 34320
rect 35760 34252 35772 34308
rect 35828 34252 35840 34308
rect 35760 33988 35840 34252
rect 35760 33932 35772 33988
rect 35828 33932 35840 33988
rect 35760 33920 35840 33932
rect 35920 34308 36000 34320
rect 35920 34252 35932 34308
rect 35988 34252 36000 34308
rect 35920 33988 36000 34252
rect 35920 33932 35932 33988
rect 35988 33932 36000 33988
rect 35920 33920 36000 33932
rect 36080 34308 36160 34320
rect 36080 34252 36092 34308
rect 36148 34252 36160 34308
rect 36080 33988 36160 34252
rect 36080 33932 36092 33988
rect 36148 33932 36160 33988
rect 36080 33920 36160 33932
rect 36240 34308 36320 34320
rect 36240 34252 36252 34308
rect 36308 34252 36320 34308
rect 36240 33988 36320 34252
rect 36240 33932 36252 33988
rect 36308 33932 36320 33988
rect 36240 33920 36320 33932
rect 36400 34308 36480 34320
rect 36400 34252 36412 34308
rect 36468 34252 36480 34308
rect 36400 33988 36480 34252
rect 36400 33932 36412 33988
rect 36468 33932 36480 33988
rect 36400 33920 36480 33932
rect 36560 34308 36640 34320
rect 36560 34252 36572 34308
rect 36628 34252 36640 34308
rect 36560 33988 36640 34252
rect 36560 33932 36572 33988
rect 36628 33932 36640 33988
rect 36560 33920 36640 33932
rect 36720 34308 36800 34320
rect 36720 34252 36732 34308
rect 36788 34252 36800 34308
rect 36720 33988 36800 34252
rect 36720 33932 36732 33988
rect 36788 33932 36800 33988
rect 36720 33920 36800 33932
rect 36880 34308 36960 34320
rect 36880 34252 36892 34308
rect 36948 34252 36960 34308
rect 36880 33988 36960 34252
rect 36880 33932 36892 33988
rect 36948 33932 36960 33988
rect 36880 33920 36960 33932
rect 37040 34308 37120 34320
rect 37040 34252 37052 34308
rect 37108 34252 37120 34308
rect 37040 33988 37120 34252
rect 37040 33932 37052 33988
rect 37108 33932 37120 33988
rect 37040 33920 37120 33932
rect 37200 34308 37280 34320
rect 37200 34252 37212 34308
rect 37268 34252 37280 34308
rect 37200 33988 37280 34252
rect 37200 33932 37212 33988
rect 37268 33932 37280 33988
rect 37200 33920 37280 33932
rect 37360 34308 37440 34320
rect 37360 34252 37372 34308
rect 37428 34252 37440 34308
rect 37360 33988 37440 34252
rect 37360 33932 37372 33988
rect 37428 33932 37440 33988
rect 37360 33920 37440 33932
rect 37520 34308 37600 34320
rect 37520 34252 37532 34308
rect 37588 34252 37600 34308
rect 37520 33988 37600 34252
rect 37520 33932 37532 33988
rect 37588 33932 37600 33988
rect 37520 33920 37600 33932
rect 37680 34308 37760 34320
rect 37680 34252 37692 34308
rect 37748 34252 37760 34308
rect 37680 33988 37760 34252
rect 37680 33932 37692 33988
rect 37748 33932 37760 33988
rect 37680 33920 37760 33932
rect 37840 34308 37920 34320
rect 37840 34252 37852 34308
rect 37908 34252 37920 34308
rect 37840 33988 37920 34252
rect 37840 33932 37852 33988
rect 37908 33932 37920 33988
rect 37840 33920 37920 33932
rect 38000 34308 38080 34320
rect 38000 34252 38012 34308
rect 38068 34252 38080 34308
rect 38000 33988 38080 34252
rect 38000 33932 38012 33988
rect 38068 33932 38080 33988
rect 38000 33920 38080 33932
rect 38160 34308 38240 34320
rect 38160 34252 38172 34308
rect 38228 34252 38240 34308
rect 38160 33988 38240 34252
rect 38160 33932 38172 33988
rect 38228 33932 38240 33988
rect 38160 33920 38240 33932
rect 38320 34308 38400 34320
rect 38320 34252 38332 34308
rect 38388 34252 38400 34308
rect 38320 33988 38400 34252
rect 38320 33932 38332 33988
rect 38388 33932 38400 33988
rect 38320 33920 38400 33932
rect 38480 34308 38560 34320
rect 38480 34252 38492 34308
rect 38548 34252 38560 34308
rect 38480 33988 38560 34252
rect 38480 33932 38492 33988
rect 38548 33932 38560 33988
rect 38480 33920 38560 33932
rect 38640 34308 38720 34320
rect 38640 34252 38652 34308
rect 38708 34252 38720 34308
rect 38640 33988 38720 34252
rect 38640 33932 38652 33988
rect 38708 33932 38720 33988
rect 38640 33920 38720 33932
rect 38800 34308 38880 34320
rect 38800 34252 38812 34308
rect 38868 34252 38880 34308
rect 38800 33988 38880 34252
rect 38800 33932 38812 33988
rect 38868 33932 38880 33988
rect 38800 33920 38880 33932
rect 38960 34308 39040 34320
rect 38960 34252 38972 34308
rect 39028 34252 39040 34308
rect 38960 33988 39040 34252
rect 38960 33932 38972 33988
rect 39028 33932 39040 33988
rect 38960 33920 39040 33932
rect 39120 34308 39200 34320
rect 39120 34252 39132 34308
rect 39188 34252 39200 34308
rect 39120 33988 39200 34252
rect 39120 33932 39132 33988
rect 39188 33932 39200 33988
rect 39120 33920 39200 33932
rect 39280 34308 39360 34320
rect 39280 34252 39292 34308
rect 39348 34252 39360 34308
rect 39280 33988 39360 34252
rect 39280 33932 39292 33988
rect 39348 33932 39360 33988
rect 39280 33920 39360 33932
rect 39440 34308 39520 34320
rect 39440 34252 39452 34308
rect 39508 34252 39520 34308
rect 39440 33988 39520 34252
rect 39440 33932 39452 33988
rect 39508 33932 39520 33988
rect 39440 33920 39520 33932
rect 39600 34308 39680 34320
rect 39600 34252 39612 34308
rect 39668 34252 39680 34308
rect 39600 33988 39680 34252
rect 39600 33932 39612 33988
rect 39668 33932 39680 33988
rect 39600 33920 39680 33932
rect 39760 34308 39840 34320
rect 39760 34252 39772 34308
rect 39828 34252 39840 34308
rect 39760 33988 39840 34252
rect 39760 33932 39772 33988
rect 39828 33932 39840 33988
rect 39760 33920 39840 33932
rect 39920 34308 40000 34320
rect 39920 34252 39932 34308
rect 39988 34252 40000 34308
rect 39920 33988 40000 34252
rect 39920 33932 39932 33988
rect 39988 33932 40000 33988
rect 39920 33920 40000 33932
rect 40080 34308 40160 34320
rect 40080 34252 40092 34308
rect 40148 34252 40160 34308
rect 40080 33988 40160 34252
rect 40080 33932 40092 33988
rect 40148 33932 40160 33988
rect 40080 33920 40160 33932
rect 40240 34308 40320 34320
rect 40240 34252 40252 34308
rect 40308 34252 40320 34308
rect 40240 33988 40320 34252
rect 40240 33932 40252 33988
rect 40308 33932 40320 33988
rect 40240 33920 40320 33932
rect 40400 34308 40480 34320
rect 40400 34252 40412 34308
rect 40468 34252 40480 34308
rect 40400 33988 40480 34252
rect 40400 33932 40412 33988
rect 40468 33932 40480 33988
rect 40400 33920 40480 33932
rect 40560 34308 40640 34320
rect 40560 34252 40572 34308
rect 40628 34252 40640 34308
rect 40560 33988 40640 34252
rect 40560 33932 40572 33988
rect 40628 33932 40640 33988
rect 40560 33920 40640 33932
rect 40720 34308 40800 34320
rect 40720 34252 40732 34308
rect 40788 34252 40800 34308
rect 40720 33988 40800 34252
rect 40720 33932 40732 33988
rect 40788 33932 40800 33988
rect 40720 33920 40800 33932
rect 40880 34308 40960 34320
rect 40880 34252 40892 34308
rect 40948 34252 40960 34308
rect 40880 33988 40960 34252
rect 40880 33932 40892 33988
rect 40948 33932 40960 33988
rect 40880 33920 40960 33932
rect 41040 34308 41120 34320
rect 41040 34252 41052 34308
rect 41108 34252 41120 34308
rect 41040 33988 41120 34252
rect 41040 33932 41052 33988
rect 41108 33932 41120 33988
rect 41040 33920 41120 33932
rect 41200 34308 41280 34320
rect 41200 34252 41212 34308
rect 41268 34252 41280 34308
rect 41200 33988 41280 34252
rect 41200 33932 41212 33988
rect 41268 33932 41280 33988
rect 41200 33920 41280 33932
rect 41360 34308 41440 34320
rect 41360 34252 41372 34308
rect 41428 34252 41440 34308
rect 41360 33988 41440 34252
rect 41360 33932 41372 33988
rect 41428 33932 41440 33988
rect 41360 33920 41440 33932
rect 41520 34308 41600 34320
rect 41520 34252 41532 34308
rect 41588 34252 41600 34308
rect 41520 33988 41600 34252
rect 41520 33932 41532 33988
rect 41588 33932 41600 33988
rect 41520 33920 41600 33932
rect 41680 34308 41760 34320
rect 41680 34252 41692 34308
rect 41748 34252 41760 34308
rect 41680 33988 41760 34252
rect 41680 33932 41692 33988
rect 41748 33932 41760 33988
rect 41680 33920 41760 33932
rect 41840 34308 41920 34320
rect 41840 34252 41852 34308
rect 41908 34252 41920 34308
rect 41840 33988 41920 34252
rect 41840 33932 41852 33988
rect 41908 33932 41920 33988
rect 41840 33920 41920 33932
rect 33520 33828 33600 33840
rect 33520 33772 33532 33828
rect 33588 33772 33600 33828
rect 33520 33508 33600 33772
rect 33520 33452 33532 33508
rect 33588 33452 33600 33508
rect 33520 33440 33600 33452
rect 33680 33828 33760 33840
rect 33680 33772 33692 33828
rect 33748 33772 33760 33828
rect 33680 33508 33760 33772
rect 33680 33452 33692 33508
rect 33748 33452 33760 33508
rect 33680 33440 33760 33452
rect 33840 33828 33920 33840
rect 33840 33772 33852 33828
rect 33908 33772 33920 33828
rect 33840 33508 33920 33772
rect 33840 33452 33852 33508
rect 33908 33452 33920 33508
rect 33840 33440 33920 33452
rect 34000 33828 34080 33840
rect 34000 33772 34012 33828
rect 34068 33772 34080 33828
rect 34000 33508 34080 33772
rect 34000 33452 34012 33508
rect 34068 33452 34080 33508
rect 34000 33440 34080 33452
rect 34160 33828 34240 33840
rect 34160 33772 34172 33828
rect 34228 33772 34240 33828
rect 34160 33508 34240 33772
rect 34160 33452 34172 33508
rect 34228 33452 34240 33508
rect 34160 33440 34240 33452
rect 34320 33828 34400 33840
rect 34320 33772 34332 33828
rect 34388 33772 34400 33828
rect 34320 33508 34400 33772
rect 34320 33452 34332 33508
rect 34388 33452 34400 33508
rect 34320 33440 34400 33452
rect 34480 33828 34560 33840
rect 34480 33772 34492 33828
rect 34548 33772 34560 33828
rect 34480 33508 34560 33772
rect 34480 33452 34492 33508
rect 34548 33452 34560 33508
rect 34480 33440 34560 33452
rect 34640 33828 34720 33840
rect 34640 33772 34652 33828
rect 34708 33772 34720 33828
rect 34640 33508 34720 33772
rect 34640 33452 34652 33508
rect 34708 33452 34720 33508
rect 34640 33440 34720 33452
rect 34800 33828 34880 33840
rect 34800 33772 34812 33828
rect 34868 33772 34880 33828
rect 34800 33508 34880 33772
rect 34800 33452 34812 33508
rect 34868 33452 34880 33508
rect 34800 33440 34880 33452
rect 34960 33828 35040 33840
rect 34960 33772 34972 33828
rect 35028 33772 35040 33828
rect 34960 33508 35040 33772
rect 34960 33452 34972 33508
rect 35028 33452 35040 33508
rect 34960 33440 35040 33452
rect 35120 33828 35200 33840
rect 35120 33772 35132 33828
rect 35188 33772 35200 33828
rect 35120 33508 35200 33772
rect 35120 33452 35132 33508
rect 35188 33452 35200 33508
rect 35120 33440 35200 33452
rect 35280 33828 35360 33840
rect 35280 33772 35292 33828
rect 35348 33772 35360 33828
rect 35280 33508 35360 33772
rect 35280 33452 35292 33508
rect 35348 33452 35360 33508
rect 35280 33440 35360 33452
rect 35440 33828 35520 33840
rect 35440 33772 35452 33828
rect 35508 33772 35520 33828
rect 35440 33508 35520 33772
rect 35440 33452 35452 33508
rect 35508 33452 35520 33508
rect 35440 33440 35520 33452
rect 35600 33828 35680 33840
rect 35600 33772 35612 33828
rect 35668 33772 35680 33828
rect 35600 33508 35680 33772
rect 35600 33452 35612 33508
rect 35668 33452 35680 33508
rect 35600 33440 35680 33452
rect 35760 33828 35840 33840
rect 35760 33772 35772 33828
rect 35828 33772 35840 33828
rect 35760 33508 35840 33772
rect 35760 33452 35772 33508
rect 35828 33452 35840 33508
rect 35760 33440 35840 33452
rect 35920 33828 36000 33840
rect 35920 33772 35932 33828
rect 35988 33772 36000 33828
rect 35920 33508 36000 33772
rect 35920 33452 35932 33508
rect 35988 33452 36000 33508
rect 35920 33440 36000 33452
rect 36080 33828 36160 33840
rect 36080 33772 36092 33828
rect 36148 33772 36160 33828
rect 36080 33508 36160 33772
rect 36080 33452 36092 33508
rect 36148 33452 36160 33508
rect 36080 33440 36160 33452
rect 36240 33828 36320 33840
rect 36240 33772 36252 33828
rect 36308 33772 36320 33828
rect 36240 33508 36320 33772
rect 36240 33452 36252 33508
rect 36308 33452 36320 33508
rect 36240 33440 36320 33452
rect 36400 33828 36480 33840
rect 36400 33772 36412 33828
rect 36468 33772 36480 33828
rect 36400 33508 36480 33772
rect 36400 33452 36412 33508
rect 36468 33452 36480 33508
rect 36400 33440 36480 33452
rect 36560 33828 36640 33840
rect 36560 33772 36572 33828
rect 36628 33772 36640 33828
rect 36560 33508 36640 33772
rect 36560 33452 36572 33508
rect 36628 33452 36640 33508
rect 36560 33440 36640 33452
rect 36720 33828 36800 33840
rect 36720 33772 36732 33828
rect 36788 33772 36800 33828
rect 36720 33508 36800 33772
rect 36720 33452 36732 33508
rect 36788 33452 36800 33508
rect 36720 33440 36800 33452
rect 36880 33828 36960 33840
rect 36880 33772 36892 33828
rect 36948 33772 36960 33828
rect 36880 33508 36960 33772
rect 36880 33452 36892 33508
rect 36948 33452 36960 33508
rect 36880 33440 36960 33452
rect 37040 33828 37120 33840
rect 37040 33772 37052 33828
rect 37108 33772 37120 33828
rect 37040 33508 37120 33772
rect 37040 33452 37052 33508
rect 37108 33452 37120 33508
rect 37040 33440 37120 33452
rect 37200 33828 37280 33840
rect 37200 33772 37212 33828
rect 37268 33772 37280 33828
rect 37200 33508 37280 33772
rect 37200 33452 37212 33508
rect 37268 33452 37280 33508
rect 37200 33440 37280 33452
rect 37360 33828 37440 33840
rect 37360 33772 37372 33828
rect 37428 33772 37440 33828
rect 37360 33508 37440 33772
rect 37360 33452 37372 33508
rect 37428 33452 37440 33508
rect 37360 33440 37440 33452
rect 37520 33828 37600 33840
rect 37520 33772 37532 33828
rect 37588 33772 37600 33828
rect 37520 33508 37600 33772
rect 37520 33452 37532 33508
rect 37588 33452 37600 33508
rect 37520 33440 37600 33452
rect 37680 33828 37760 33840
rect 37680 33772 37692 33828
rect 37748 33772 37760 33828
rect 37680 33508 37760 33772
rect 37680 33452 37692 33508
rect 37748 33452 37760 33508
rect 37680 33440 37760 33452
rect 37840 33828 37920 33840
rect 37840 33772 37852 33828
rect 37908 33772 37920 33828
rect 37840 33508 37920 33772
rect 37840 33452 37852 33508
rect 37908 33452 37920 33508
rect 37840 33440 37920 33452
rect 38000 33828 38080 33840
rect 38000 33772 38012 33828
rect 38068 33772 38080 33828
rect 38000 33508 38080 33772
rect 38000 33452 38012 33508
rect 38068 33452 38080 33508
rect 38000 33440 38080 33452
rect 38160 33828 38240 33840
rect 38160 33772 38172 33828
rect 38228 33772 38240 33828
rect 38160 33508 38240 33772
rect 38160 33452 38172 33508
rect 38228 33452 38240 33508
rect 38160 33440 38240 33452
rect 38320 33828 38400 33840
rect 38320 33772 38332 33828
rect 38388 33772 38400 33828
rect 38320 33508 38400 33772
rect 38320 33452 38332 33508
rect 38388 33452 38400 33508
rect 38320 33440 38400 33452
rect 38480 33828 38560 33840
rect 38480 33772 38492 33828
rect 38548 33772 38560 33828
rect 38480 33508 38560 33772
rect 38480 33452 38492 33508
rect 38548 33452 38560 33508
rect 38480 33440 38560 33452
rect 38640 33828 38720 33840
rect 38640 33772 38652 33828
rect 38708 33772 38720 33828
rect 38640 33508 38720 33772
rect 38640 33452 38652 33508
rect 38708 33452 38720 33508
rect 38640 33440 38720 33452
rect 38800 33828 38880 33840
rect 38800 33772 38812 33828
rect 38868 33772 38880 33828
rect 38800 33508 38880 33772
rect 38800 33452 38812 33508
rect 38868 33452 38880 33508
rect 38800 33440 38880 33452
rect 38960 33828 39040 33840
rect 38960 33772 38972 33828
rect 39028 33772 39040 33828
rect 38960 33508 39040 33772
rect 38960 33452 38972 33508
rect 39028 33452 39040 33508
rect 38960 33440 39040 33452
rect 39120 33828 39200 33840
rect 39120 33772 39132 33828
rect 39188 33772 39200 33828
rect 39120 33508 39200 33772
rect 39120 33452 39132 33508
rect 39188 33452 39200 33508
rect 39120 33440 39200 33452
rect 39280 33828 39360 33840
rect 39280 33772 39292 33828
rect 39348 33772 39360 33828
rect 39280 33508 39360 33772
rect 39280 33452 39292 33508
rect 39348 33452 39360 33508
rect 39280 33440 39360 33452
rect 39440 33828 39520 33840
rect 39440 33772 39452 33828
rect 39508 33772 39520 33828
rect 39440 33508 39520 33772
rect 39440 33452 39452 33508
rect 39508 33452 39520 33508
rect 39440 33440 39520 33452
rect 39600 33828 39680 33840
rect 39600 33772 39612 33828
rect 39668 33772 39680 33828
rect 39600 33508 39680 33772
rect 39600 33452 39612 33508
rect 39668 33452 39680 33508
rect 39600 33440 39680 33452
rect 39760 33828 39840 33840
rect 39760 33772 39772 33828
rect 39828 33772 39840 33828
rect 39760 33508 39840 33772
rect 39760 33452 39772 33508
rect 39828 33452 39840 33508
rect 39760 33440 39840 33452
rect 39920 33828 40000 33840
rect 39920 33772 39932 33828
rect 39988 33772 40000 33828
rect 39920 33508 40000 33772
rect 39920 33452 39932 33508
rect 39988 33452 40000 33508
rect 39920 33440 40000 33452
rect 40080 33828 40160 33840
rect 40080 33772 40092 33828
rect 40148 33772 40160 33828
rect 40080 33508 40160 33772
rect 40080 33452 40092 33508
rect 40148 33452 40160 33508
rect 40080 33440 40160 33452
rect 40240 33828 40320 33840
rect 40240 33772 40252 33828
rect 40308 33772 40320 33828
rect 40240 33508 40320 33772
rect 40240 33452 40252 33508
rect 40308 33452 40320 33508
rect 40240 33440 40320 33452
rect 40400 33828 40480 33840
rect 40400 33772 40412 33828
rect 40468 33772 40480 33828
rect 40400 33508 40480 33772
rect 40400 33452 40412 33508
rect 40468 33452 40480 33508
rect 40400 33440 40480 33452
rect 40560 33828 40640 33840
rect 40560 33772 40572 33828
rect 40628 33772 40640 33828
rect 40560 33508 40640 33772
rect 40560 33452 40572 33508
rect 40628 33452 40640 33508
rect 40560 33440 40640 33452
rect 40720 33828 40800 33840
rect 40720 33772 40732 33828
rect 40788 33772 40800 33828
rect 40720 33508 40800 33772
rect 40720 33452 40732 33508
rect 40788 33452 40800 33508
rect 40720 33440 40800 33452
rect 40880 33828 40960 33840
rect 40880 33772 40892 33828
rect 40948 33772 40960 33828
rect 40880 33508 40960 33772
rect 40880 33452 40892 33508
rect 40948 33452 40960 33508
rect 40880 33440 40960 33452
rect 41040 33828 41120 33840
rect 41040 33772 41052 33828
rect 41108 33772 41120 33828
rect 41040 33508 41120 33772
rect 41040 33452 41052 33508
rect 41108 33452 41120 33508
rect 41040 33440 41120 33452
rect 41200 33828 41280 33840
rect 41200 33772 41212 33828
rect 41268 33772 41280 33828
rect 41200 33508 41280 33772
rect 41200 33452 41212 33508
rect 41268 33452 41280 33508
rect 41200 33440 41280 33452
rect 41360 33828 41440 33840
rect 41360 33772 41372 33828
rect 41428 33772 41440 33828
rect 41360 33508 41440 33772
rect 41360 33452 41372 33508
rect 41428 33452 41440 33508
rect 41360 33440 41440 33452
rect 41520 33828 41600 33840
rect 41520 33772 41532 33828
rect 41588 33772 41600 33828
rect 41520 33508 41600 33772
rect 41520 33452 41532 33508
rect 41588 33452 41600 33508
rect 41520 33440 41600 33452
rect 41680 33828 41760 33840
rect 41680 33772 41692 33828
rect 41748 33772 41760 33828
rect 41680 33508 41760 33772
rect 41680 33452 41692 33508
rect 41748 33452 41760 33508
rect 41680 33440 41760 33452
rect 41840 33828 41920 33840
rect 41840 33772 41852 33828
rect 41908 33772 41920 33828
rect 41840 33508 41920 33772
rect 41840 33452 41852 33508
rect 41908 33452 41920 33508
rect 41840 33440 41920 33452
rect 23120 33348 23200 33360
rect 23120 33292 23132 33348
rect 23188 33292 23200 33348
rect 23120 33028 23200 33292
rect 23120 32972 23132 33028
rect 23188 32972 23200 33028
rect 23120 32960 23200 32972
rect 23280 33348 23360 33360
rect 23280 33292 23292 33348
rect 23348 33292 23360 33348
rect 23280 33028 23360 33292
rect 23280 32972 23292 33028
rect 23348 32972 23360 33028
rect 23280 32960 23360 32972
rect 23440 33348 23520 33360
rect 23440 33292 23452 33348
rect 23508 33292 23520 33348
rect 23440 33028 23520 33292
rect 23440 32972 23452 33028
rect 23508 32972 23520 33028
rect 23440 32960 23520 32972
rect 23600 33348 23680 33360
rect 23600 33292 23612 33348
rect 23668 33292 23680 33348
rect 23600 33028 23680 33292
rect 23600 32972 23612 33028
rect 23668 32972 23680 33028
rect 23600 32960 23680 32972
rect 23760 33348 23840 33360
rect 23760 33292 23772 33348
rect 23828 33292 23840 33348
rect 23760 33028 23840 33292
rect 23760 32972 23772 33028
rect 23828 32972 23840 33028
rect 23760 32960 23840 32972
rect 23920 33348 24000 33360
rect 23920 33292 23932 33348
rect 23988 33292 24000 33348
rect 23920 33028 24000 33292
rect 23920 32972 23932 33028
rect 23988 32972 24000 33028
rect 23920 32960 24000 32972
rect 24080 33348 24160 33360
rect 24080 33292 24092 33348
rect 24148 33292 24160 33348
rect 24080 33028 24160 33292
rect 24080 32972 24092 33028
rect 24148 32972 24160 33028
rect 24080 32960 24160 32972
rect 24240 33348 24320 33360
rect 24240 33292 24252 33348
rect 24308 33292 24320 33348
rect 24240 33028 24320 33292
rect 24240 32972 24252 33028
rect 24308 32972 24320 33028
rect 24240 32960 24320 32972
rect 24400 33348 24480 33360
rect 24400 33292 24412 33348
rect 24468 33292 24480 33348
rect 24400 33028 24480 33292
rect 24400 32972 24412 33028
rect 24468 32972 24480 33028
rect 24400 32960 24480 32972
rect 24560 33348 24640 33360
rect 24560 33292 24572 33348
rect 24628 33292 24640 33348
rect 24560 33028 24640 33292
rect 24560 32972 24572 33028
rect 24628 32972 24640 33028
rect 24560 32960 24640 32972
rect 24720 33348 24800 33360
rect 24720 33292 24732 33348
rect 24788 33292 24800 33348
rect 24720 33028 24800 33292
rect 24720 32972 24732 33028
rect 24788 32972 24800 33028
rect 24720 32960 24800 32972
rect 24880 33348 24960 33360
rect 24880 33292 24892 33348
rect 24948 33292 24960 33348
rect 24880 33028 24960 33292
rect 24880 32972 24892 33028
rect 24948 32972 24960 33028
rect 24880 32960 24960 32972
rect 25040 33348 25120 33360
rect 25040 33292 25052 33348
rect 25108 33292 25120 33348
rect 25040 33028 25120 33292
rect 25040 32972 25052 33028
rect 25108 32972 25120 33028
rect 25040 32960 25120 32972
rect 25200 33348 25280 33360
rect 25200 33292 25212 33348
rect 25268 33292 25280 33348
rect 25200 33028 25280 33292
rect 25200 32972 25212 33028
rect 25268 32972 25280 33028
rect 25200 32960 25280 32972
rect 25360 33348 25440 33360
rect 25360 33292 25372 33348
rect 25428 33292 25440 33348
rect 25360 33028 25440 33292
rect 25360 32972 25372 33028
rect 25428 32972 25440 33028
rect 25360 32960 25440 32972
rect 25520 33348 25600 33360
rect 25520 33292 25532 33348
rect 25588 33292 25600 33348
rect 25520 33028 25600 33292
rect 25520 32972 25532 33028
rect 25588 32972 25600 33028
rect 25520 32960 25600 32972
rect 25680 33348 25760 33360
rect 25680 33292 25692 33348
rect 25748 33292 25760 33348
rect 25680 33028 25760 33292
rect 25680 32972 25692 33028
rect 25748 32972 25760 33028
rect 25680 32960 25760 32972
rect 25840 33348 25920 33360
rect 25840 33292 25852 33348
rect 25908 33292 25920 33348
rect 25840 33028 25920 33292
rect 25840 32972 25852 33028
rect 25908 32972 25920 33028
rect 25840 32960 25920 32972
rect 26000 33348 26080 33360
rect 26000 33292 26012 33348
rect 26068 33292 26080 33348
rect 26000 33028 26080 33292
rect 26000 32972 26012 33028
rect 26068 32972 26080 33028
rect 26000 32960 26080 32972
rect 26160 33348 26240 33360
rect 26160 33292 26172 33348
rect 26228 33292 26240 33348
rect 26160 33028 26240 33292
rect 26160 32972 26172 33028
rect 26228 32972 26240 33028
rect 26160 32960 26240 32972
rect 26320 33348 26400 33360
rect 26320 33292 26332 33348
rect 26388 33292 26400 33348
rect 26320 33028 26400 33292
rect 26320 32972 26332 33028
rect 26388 32972 26400 33028
rect 26320 32960 26400 32972
rect 26480 33348 26560 33360
rect 26480 33292 26492 33348
rect 26548 33292 26560 33348
rect 26480 33028 26560 33292
rect 26480 32972 26492 33028
rect 26548 32972 26560 33028
rect 26480 32960 26560 32972
rect 26640 33348 26720 33360
rect 26640 33292 26652 33348
rect 26708 33292 26720 33348
rect 26640 33028 26720 33292
rect 26640 32972 26652 33028
rect 26708 32972 26720 33028
rect 26640 32960 26720 32972
rect 26800 33348 26880 33360
rect 26800 33292 26812 33348
rect 26868 33292 26880 33348
rect 26800 33028 26880 33292
rect 26800 32972 26812 33028
rect 26868 32972 26880 33028
rect 26800 32960 26880 32972
rect 26960 33348 27040 33360
rect 26960 33292 26972 33348
rect 27028 33292 27040 33348
rect 26960 33028 27040 33292
rect 26960 32972 26972 33028
rect 27028 32972 27040 33028
rect 26960 32960 27040 32972
rect 27120 33348 27200 33360
rect 27120 33292 27132 33348
rect 27188 33292 27200 33348
rect 27120 33028 27200 33292
rect 27120 32972 27132 33028
rect 27188 32972 27200 33028
rect 27120 32960 27200 32972
rect 27280 33348 27360 33360
rect 27280 33292 27292 33348
rect 27348 33292 27360 33348
rect 27280 33028 27360 33292
rect 27280 32972 27292 33028
rect 27348 32972 27360 33028
rect 27280 32960 27360 32972
rect 27440 33348 27520 33360
rect 27440 33292 27452 33348
rect 27508 33292 27520 33348
rect 27440 33028 27520 33292
rect 27440 32972 27452 33028
rect 27508 32972 27520 33028
rect 27440 32960 27520 32972
rect 27600 33348 27680 33360
rect 27600 33292 27612 33348
rect 27668 33292 27680 33348
rect 27600 33028 27680 33292
rect 27600 32972 27612 33028
rect 27668 32972 27680 33028
rect 27600 32960 27680 32972
rect 27760 33348 27840 33360
rect 27760 33292 27772 33348
rect 27828 33292 27840 33348
rect 27760 33028 27840 33292
rect 27760 32972 27772 33028
rect 27828 32972 27840 33028
rect 27760 32960 27840 32972
rect 27920 33348 28000 33360
rect 27920 33292 27932 33348
rect 27988 33292 28000 33348
rect 27920 33028 28000 33292
rect 27920 32972 27932 33028
rect 27988 32972 28000 33028
rect 27920 32960 28000 32972
rect 28080 33348 28160 33360
rect 28080 33292 28092 33348
rect 28148 33292 28160 33348
rect 28080 33028 28160 33292
rect 28080 32972 28092 33028
rect 28148 32972 28160 33028
rect 28080 32960 28160 32972
rect 28240 33348 28320 33360
rect 28240 33292 28252 33348
rect 28308 33292 28320 33348
rect 28240 33028 28320 33292
rect 28240 32972 28252 33028
rect 28308 32972 28320 33028
rect 28240 32960 28320 32972
rect 28400 33348 28480 33360
rect 28400 33292 28412 33348
rect 28468 33292 28480 33348
rect 28400 33028 28480 33292
rect 28400 32972 28412 33028
rect 28468 32972 28480 33028
rect 28400 32960 28480 32972
rect 28560 33348 28640 33360
rect 28560 33292 28572 33348
rect 28628 33292 28640 33348
rect 28560 33028 28640 33292
rect 28560 32972 28572 33028
rect 28628 32972 28640 33028
rect 28560 32960 28640 32972
rect 28720 33348 28800 33360
rect 28720 33292 28732 33348
rect 28788 33292 28800 33348
rect 28720 33028 28800 33292
rect 28720 32972 28732 33028
rect 28788 32972 28800 33028
rect 28720 32960 28800 32972
rect 28880 33348 28960 33360
rect 28880 33292 28892 33348
rect 28948 33292 28960 33348
rect 28880 33028 28960 33292
rect 28880 32972 28892 33028
rect 28948 32972 28960 33028
rect 28880 32960 28960 32972
rect 29040 33348 29120 33360
rect 29040 33292 29052 33348
rect 29108 33292 29120 33348
rect 29040 33028 29120 33292
rect 29040 32972 29052 33028
rect 29108 32972 29120 33028
rect 29040 32960 29120 32972
rect 29200 33348 29280 33360
rect 29200 33292 29212 33348
rect 29268 33292 29280 33348
rect 29200 33028 29280 33292
rect 29200 32972 29212 33028
rect 29268 32972 29280 33028
rect 29200 32960 29280 32972
rect 29360 33348 29440 33360
rect 29360 33292 29372 33348
rect 29428 33292 29440 33348
rect 29360 33028 29440 33292
rect 29360 32972 29372 33028
rect 29428 32972 29440 33028
rect 29360 32960 29440 32972
rect 23120 32868 23200 32880
rect 23120 32812 23132 32868
rect 23188 32812 23200 32868
rect 23120 32548 23200 32812
rect 23120 32492 23132 32548
rect 23188 32492 23200 32548
rect 23120 32480 23200 32492
rect 23280 32868 23360 32880
rect 23280 32812 23292 32868
rect 23348 32812 23360 32868
rect 23280 32548 23360 32812
rect 23280 32492 23292 32548
rect 23348 32492 23360 32548
rect 23280 32480 23360 32492
rect 23440 32868 23520 32880
rect 23440 32812 23452 32868
rect 23508 32812 23520 32868
rect 23440 32548 23520 32812
rect 23440 32492 23452 32548
rect 23508 32492 23520 32548
rect 23440 32480 23520 32492
rect 23600 32868 23680 32880
rect 23600 32812 23612 32868
rect 23668 32812 23680 32868
rect 23600 32548 23680 32812
rect 23600 32492 23612 32548
rect 23668 32492 23680 32548
rect 23600 32480 23680 32492
rect 23760 32868 23840 32880
rect 23760 32812 23772 32868
rect 23828 32812 23840 32868
rect 23760 32548 23840 32812
rect 23760 32492 23772 32548
rect 23828 32492 23840 32548
rect 23760 32480 23840 32492
rect 23920 32868 24000 32880
rect 23920 32812 23932 32868
rect 23988 32812 24000 32868
rect 23920 32548 24000 32812
rect 23920 32492 23932 32548
rect 23988 32492 24000 32548
rect 23920 32480 24000 32492
rect 24080 32868 24160 32880
rect 24080 32812 24092 32868
rect 24148 32812 24160 32868
rect 24080 32548 24160 32812
rect 24080 32492 24092 32548
rect 24148 32492 24160 32548
rect 24080 32480 24160 32492
rect 24240 32868 24320 32880
rect 24240 32812 24252 32868
rect 24308 32812 24320 32868
rect 24240 32548 24320 32812
rect 24240 32492 24252 32548
rect 24308 32492 24320 32548
rect 24240 32480 24320 32492
rect 24400 32868 24480 32880
rect 24400 32812 24412 32868
rect 24468 32812 24480 32868
rect 24400 32548 24480 32812
rect 24400 32492 24412 32548
rect 24468 32492 24480 32548
rect 24400 32480 24480 32492
rect 24560 32868 24640 32880
rect 24560 32812 24572 32868
rect 24628 32812 24640 32868
rect 24560 32548 24640 32812
rect 24560 32492 24572 32548
rect 24628 32492 24640 32548
rect 24560 32480 24640 32492
rect 24720 32868 24800 32880
rect 24720 32812 24732 32868
rect 24788 32812 24800 32868
rect 24720 32548 24800 32812
rect 24720 32492 24732 32548
rect 24788 32492 24800 32548
rect 24720 32480 24800 32492
rect 24880 32868 24960 32880
rect 24880 32812 24892 32868
rect 24948 32812 24960 32868
rect 24880 32548 24960 32812
rect 24880 32492 24892 32548
rect 24948 32492 24960 32548
rect 24880 32480 24960 32492
rect 25040 32868 25120 32880
rect 25040 32812 25052 32868
rect 25108 32812 25120 32868
rect 25040 32548 25120 32812
rect 25040 32492 25052 32548
rect 25108 32492 25120 32548
rect 25040 32480 25120 32492
rect 25200 32868 25280 32880
rect 25200 32812 25212 32868
rect 25268 32812 25280 32868
rect 25200 32548 25280 32812
rect 25200 32492 25212 32548
rect 25268 32492 25280 32548
rect 25200 32480 25280 32492
rect 25360 32868 25440 32880
rect 25360 32812 25372 32868
rect 25428 32812 25440 32868
rect 25360 32548 25440 32812
rect 25360 32492 25372 32548
rect 25428 32492 25440 32548
rect 25360 32480 25440 32492
rect 25520 32868 25600 32880
rect 25520 32812 25532 32868
rect 25588 32812 25600 32868
rect 25520 32548 25600 32812
rect 25520 32492 25532 32548
rect 25588 32492 25600 32548
rect 25520 32480 25600 32492
rect 25680 32868 25760 32880
rect 25680 32812 25692 32868
rect 25748 32812 25760 32868
rect 25680 32548 25760 32812
rect 25680 32492 25692 32548
rect 25748 32492 25760 32548
rect 25680 32480 25760 32492
rect 25840 32868 25920 32880
rect 25840 32812 25852 32868
rect 25908 32812 25920 32868
rect 25840 32548 25920 32812
rect 25840 32492 25852 32548
rect 25908 32492 25920 32548
rect 25840 32480 25920 32492
rect 26000 32868 26080 32880
rect 26000 32812 26012 32868
rect 26068 32812 26080 32868
rect 26000 32548 26080 32812
rect 26000 32492 26012 32548
rect 26068 32492 26080 32548
rect 26000 32480 26080 32492
rect 26160 32868 26240 32880
rect 26160 32812 26172 32868
rect 26228 32812 26240 32868
rect 26160 32548 26240 32812
rect 26160 32492 26172 32548
rect 26228 32492 26240 32548
rect 26160 32480 26240 32492
rect 26320 32868 26400 32880
rect 26320 32812 26332 32868
rect 26388 32812 26400 32868
rect 26320 32548 26400 32812
rect 26320 32492 26332 32548
rect 26388 32492 26400 32548
rect 26320 32480 26400 32492
rect 26480 32868 26560 32880
rect 26480 32812 26492 32868
rect 26548 32812 26560 32868
rect 26480 32548 26560 32812
rect 26480 32492 26492 32548
rect 26548 32492 26560 32548
rect 26480 32480 26560 32492
rect 26640 32868 26720 32880
rect 26640 32812 26652 32868
rect 26708 32812 26720 32868
rect 26640 32548 26720 32812
rect 26640 32492 26652 32548
rect 26708 32492 26720 32548
rect 26640 32480 26720 32492
rect 26800 32868 26880 32880
rect 26800 32812 26812 32868
rect 26868 32812 26880 32868
rect 26800 32548 26880 32812
rect 26800 32492 26812 32548
rect 26868 32492 26880 32548
rect 26800 32480 26880 32492
rect 26960 32868 27040 32880
rect 26960 32812 26972 32868
rect 27028 32812 27040 32868
rect 26960 32548 27040 32812
rect 26960 32492 26972 32548
rect 27028 32492 27040 32548
rect 26960 32480 27040 32492
rect 27120 32868 27200 32880
rect 27120 32812 27132 32868
rect 27188 32812 27200 32868
rect 27120 32548 27200 32812
rect 27120 32492 27132 32548
rect 27188 32492 27200 32548
rect 27120 32480 27200 32492
rect 27280 32868 27360 32880
rect 27280 32812 27292 32868
rect 27348 32812 27360 32868
rect 27280 32548 27360 32812
rect 27280 32492 27292 32548
rect 27348 32492 27360 32548
rect 27280 32480 27360 32492
rect 27440 32868 27520 32880
rect 27440 32812 27452 32868
rect 27508 32812 27520 32868
rect 27440 32548 27520 32812
rect 27440 32492 27452 32548
rect 27508 32492 27520 32548
rect 27440 32480 27520 32492
rect 27600 32868 27680 32880
rect 27600 32812 27612 32868
rect 27668 32812 27680 32868
rect 27600 32548 27680 32812
rect 27600 32492 27612 32548
rect 27668 32492 27680 32548
rect 27600 32480 27680 32492
rect 27760 32868 27840 32880
rect 27760 32812 27772 32868
rect 27828 32812 27840 32868
rect 27760 32548 27840 32812
rect 27760 32492 27772 32548
rect 27828 32492 27840 32548
rect 27760 32480 27840 32492
rect 27920 32868 28000 32880
rect 27920 32812 27932 32868
rect 27988 32812 28000 32868
rect 27920 32548 28000 32812
rect 27920 32492 27932 32548
rect 27988 32492 28000 32548
rect 27920 32480 28000 32492
rect 28080 32868 28160 32880
rect 28080 32812 28092 32868
rect 28148 32812 28160 32868
rect 28080 32548 28160 32812
rect 28080 32492 28092 32548
rect 28148 32492 28160 32548
rect 28080 32480 28160 32492
rect 28240 32868 28320 32880
rect 28240 32812 28252 32868
rect 28308 32812 28320 32868
rect 28240 32548 28320 32812
rect 28240 32492 28252 32548
rect 28308 32492 28320 32548
rect 28240 32480 28320 32492
rect 28400 32868 28480 32880
rect 28400 32812 28412 32868
rect 28468 32812 28480 32868
rect 28400 32548 28480 32812
rect 28400 32492 28412 32548
rect 28468 32492 28480 32548
rect 28400 32480 28480 32492
rect 28560 32868 28640 32880
rect 28560 32812 28572 32868
rect 28628 32812 28640 32868
rect 28560 32548 28640 32812
rect 28560 32492 28572 32548
rect 28628 32492 28640 32548
rect 28560 32480 28640 32492
rect 28720 32868 28800 32880
rect 28720 32812 28732 32868
rect 28788 32812 28800 32868
rect 28720 32548 28800 32812
rect 28720 32492 28732 32548
rect 28788 32492 28800 32548
rect 28720 32480 28800 32492
rect 28880 32868 28960 32880
rect 28880 32812 28892 32868
rect 28948 32812 28960 32868
rect 28880 32548 28960 32812
rect 28880 32492 28892 32548
rect 28948 32492 28960 32548
rect 28880 32480 28960 32492
rect 29040 32868 29120 32880
rect 29040 32812 29052 32868
rect 29108 32812 29120 32868
rect 29040 32548 29120 32812
rect 29040 32492 29052 32548
rect 29108 32492 29120 32548
rect 29040 32480 29120 32492
rect 29200 32868 29280 32880
rect 29200 32812 29212 32868
rect 29268 32812 29280 32868
rect 29200 32548 29280 32812
rect 29200 32492 29212 32548
rect 29268 32492 29280 32548
rect 29200 32480 29280 32492
rect 29360 32868 29440 32880
rect 29360 32812 29372 32868
rect 29428 32812 29440 32868
rect 29360 32548 29440 32812
rect 29360 32492 29372 32548
rect 29428 32492 29440 32548
rect 29360 32480 29440 32492
rect 23120 32388 23200 32400
rect 23120 32332 23132 32388
rect 23188 32332 23200 32388
rect 23120 32068 23200 32332
rect 23120 32012 23132 32068
rect 23188 32012 23200 32068
rect 23120 31748 23200 32012
rect 23120 31692 23132 31748
rect 23188 31692 23200 31748
rect 23120 31428 23200 31692
rect 23120 31372 23132 31428
rect 23188 31372 23200 31428
rect 23120 31108 23200 31372
rect 23120 31052 23132 31108
rect 23188 31052 23200 31108
rect 23120 30788 23200 31052
rect 23120 30732 23132 30788
rect 23188 30732 23200 30788
rect 23120 30468 23200 30732
rect 23120 30412 23132 30468
rect 23188 30412 23200 30468
rect 23120 30400 23200 30412
rect 23280 32388 23360 32400
rect 23280 32332 23292 32388
rect 23348 32332 23360 32388
rect 23280 32068 23360 32332
rect 23280 32012 23292 32068
rect 23348 32012 23360 32068
rect 23280 31748 23360 32012
rect 23280 31692 23292 31748
rect 23348 31692 23360 31748
rect 23280 31428 23360 31692
rect 23280 31372 23292 31428
rect 23348 31372 23360 31428
rect 23280 31108 23360 31372
rect 23280 31052 23292 31108
rect 23348 31052 23360 31108
rect 23280 30788 23360 31052
rect 23280 30732 23292 30788
rect 23348 30732 23360 30788
rect 23280 30468 23360 30732
rect 23280 30412 23292 30468
rect 23348 30412 23360 30468
rect 23280 30400 23360 30412
rect 23440 32388 23520 32400
rect 23440 32332 23452 32388
rect 23508 32332 23520 32388
rect 23440 32068 23520 32332
rect 23440 32012 23452 32068
rect 23508 32012 23520 32068
rect 23440 31748 23520 32012
rect 23440 31692 23452 31748
rect 23508 31692 23520 31748
rect 23440 31428 23520 31692
rect 23440 31372 23452 31428
rect 23508 31372 23520 31428
rect 23440 31108 23520 31372
rect 23440 31052 23452 31108
rect 23508 31052 23520 31108
rect 23440 30788 23520 31052
rect 23440 30732 23452 30788
rect 23508 30732 23520 30788
rect 23440 30468 23520 30732
rect 23440 30412 23452 30468
rect 23508 30412 23520 30468
rect 23440 30400 23520 30412
rect 23600 32388 23680 32400
rect 23600 32332 23612 32388
rect 23668 32332 23680 32388
rect 23600 32068 23680 32332
rect 23600 32012 23612 32068
rect 23668 32012 23680 32068
rect 23600 31748 23680 32012
rect 23600 31692 23612 31748
rect 23668 31692 23680 31748
rect 23600 31428 23680 31692
rect 23600 31372 23612 31428
rect 23668 31372 23680 31428
rect 23600 31108 23680 31372
rect 23600 31052 23612 31108
rect 23668 31052 23680 31108
rect 23600 30788 23680 31052
rect 23600 30732 23612 30788
rect 23668 30732 23680 30788
rect 23600 30468 23680 30732
rect 23600 30412 23612 30468
rect 23668 30412 23680 30468
rect 23600 30400 23680 30412
rect 23760 32388 23840 32400
rect 23760 32332 23772 32388
rect 23828 32332 23840 32388
rect 23760 32068 23840 32332
rect 23760 32012 23772 32068
rect 23828 32012 23840 32068
rect 23760 31748 23840 32012
rect 23760 31692 23772 31748
rect 23828 31692 23840 31748
rect 23760 31428 23840 31692
rect 23760 31372 23772 31428
rect 23828 31372 23840 31428
rect 23760 31108 23840 31372
rect 23760 31052 23772 31108
rect 23828 31052 23840 31108
rect 23760 30788 23840 31052
rect 23760 30732 23772 30788
rect 23828 30732 23840 30788
rect 23760 30468 23840 30732
rect 23760 30412 23772 30468
rect 23828 30412 23840 30468
rect 23760 30400 23840 30412
rect 23920 32388 24000 32400
rect 23920 32332 23932 32388
rect 23988 32332 24000 32388
rect 23920 32068 24000 32332
rect 23920 32012 23932 32068
rect 23988 32012 24000 32068
rect 23920 31748 24000 32012
rect 23920 31692 23932 31748
rect 23988 31692 24000 31748
rect 23920 31428 24000 31692
rect 23920 31372 23932 31428
rect 23988 31372 24000 31428
rect 23920 31108 24000 31372
rect 23920 31052 23932 31108
rect 23988 31052 24000 31108
rect 23920 30788 24000 31052
rect 23920 30732 23932 30788
rect 23988 30732 24000 30788
rect 23920 30468 24000 30732
rect 23920 30412 23932 30468
rect 23988 30412 24000 30468
rect 23920 30400 24000 30412
rect 24080 32388 24160 32400
rect 24080 32332 24092 32388
rect 24148 32332 24160 32388
rect 24080 32068 24160 32332
rect 24080 32012 24092 32068
rect 24148 32012 24160 32068
rect 24080 31748 24160 32012
rect 24080 31692 24092 31748
rect 24148 31692 24160 31748
rect 24080 31428 24160 31692
rect 24080 31372 24092 31428
rect 24148 31372 24160 31428
rect 24080 31108 24160 31372
rect 24080 31052 24092 31108
rect 24148 31052 24160 31108
rect 24080 30788 24160 31052
rect 24080 30732 24092 30788
rect 24148 30732 24160 30788
rect 24080 30468 24160 30732
rect 24080 30412 24092 30468
rect 24148 30412 24160 30468
rect 24080 30400 24160 30412
rect 24240 32388 24320 32400
rect 24240 32332 24252 32388
rect 24308 32332 24320 32388
rect 24240 32068 24320 32332
rect 24240 32012 24252 32068
rect 24308 32012 24320 32068
rect 24240 31748 24320 32012
rect 24240 31692 24252 31748
rect 24308 31692 24320 31748
rect 24240 31428 24320 31692
rect 24240 31372 24252 31428
rect 24308 31372 24320 31428
rect 24240 31108 24320 31372
rect 24240 31052 24252 31108
rect 24308 31052 24320 31108
rect 24240 30788 24320 31052
rect 24240 30732 24252 30788
rect 24308 30732 24320 30788
rect 24240 30468 24320 30732
rect 24240 30412 24252 30468
rect 24308 30412 24320 30468
rect 24240 30400 24320 30412
rect 24400 32388 24480 32400
rect 24400 32332 24412 32388
rect 24468 32332 24480 32388
rect 24400 32068 24480 32332
rect 24400 32012 24412 32068
rect 24468 32012 24480 32068
rect 24400 31748 24480 32012
rect 24400 31692 24412 31748
rect 24468 31692 24480 31748
rect 24400 31428 24480 31692
rect 24400 31372 24412 31428
rect 24468 31372 24480 31428
rect 24400 31108 24480 31372
rect 24400 31052 24412 31108
rect 24468 31052 24480 31108
rect 24400 30788 24480 31052
rect 24400 30732 24412 30788
rect 24468 30732 24480 30788
rect 24400 30468 24480 30732
rect 24400 30412 24412 30468
rect 24468 30412 24480 30468
rect 24400 30400 24480 30412
rect 24560 32388 24640 32400
rect 24560 32332 24572 32388
rect 24628 32332 24640 32388
rect 24560 32068 24640 32332
rect 24560 32012 24572 32068
rect 24628 32012 24640 32068
rect 24560 31748 24640 32012
rect 24560 31692 24572 31748
rect 24628 31692 24640 31748
rect 24560 31428 24640 31692
rect 24560 31372 24572 31428
rect 24628 31372 24640 31428
rect 24560 31108 24640 31372
rect 24560 31052 24572 31108
rect 24628 31052 24640 31108
rect 24560 30788 24640 31052
rect 24560 30732 24572 30788
rect 24628 30732 24640 30788
rect 24560 30468 24640 30732
rect 24560 30412 24572 30468
rect 24628 30412 24640 30468
rect 24560 30400 24640 30412
rect 24720 32388 24800 32400
rect 24720 32332 24732 32388
rect 24788 32332 24800 32388
rect 24720 32068 24800 32332
rect 24720 32012 24732 32068
rect 24788 32012 24800 32068
rect 24720 31748 24800 32012
rect 24720 31692 24732 31748
rect 24788 31692 24800 31748
rect 24720 31428 24800 31692
rect 24720 31372 24732 31428
rect 24788 31372 24800 31428
rect 24720 31108 24800 31372
rect 24720 31052 24732 31108
rect 24788 31052 24800 31108
rect 24720 30788 24800 31052
rect 24720 30732 24732 30788
rect 24788 30732 24800 30788
rect 24720 30468 24800 30732
rect 24720 30412 24732 30468
rect 24788 30412 24800 30468
rect 24720 30400 24800 30412
rect 24880 32388 24960 32400
rect 24880 32332 24892 32388
rect 24948 32332 24960 32388
rect 24880 32068 24960 32332
rect 24880 32012 24892 32068
rect 24948 32012 24960 32068
rect 24880 31748 24960 32012
rect 24880 31692 24892 31748
rect 24948 31692 24960 31748
rect 24880 31428 24960 31692
rect 24880 31372 24892 31428
rect 24948 31372 24960 31428
rect 24880 31108 24960 31372
rect 24880 31052 24892 31108
rect 24948 31052 24960 31108
rect 24880 30788 24960 31052
rect 24880 30732 24892 30788
rect 24948 30732 24960 30788
rect 24880 30468 24960 30732
rect 24880 30412 24892 30468
rect 24948 30412 24960 30468
rect 24880 30400 24960 30412
rect 25040 32388 25120 32400
rect 25040 32332 25052 32388
rect 25108 32332 25120 32388
rect 25040 32068 25120 32332
rect 25040 32012 25052 32068
rect 25108 32012 25120 32068
rect 25040 31748 25120 32012
rect 25040 31692 25052 31748
rect 25108 31692 25120 31748
rect 25040 31428 25120 31692
rect 25040 31372 25052 31428
rect 25108 31372 25120 31428
rect 25040 31108 25120 31372
rect 25040 31052 25052 31108
rect 25108 31052 25120 31108
rect 25040 30788 25120 31052
rect 25040 30732 25052 30788
rect 25108 30732 25120 30788
rect 25040 30468 25120 30732
rect 25040 30412 25052 30468
rect 25108 30412 25120 30468
rect 25040 30400 25120 30412
rect 25200 32388 25280 32400
rect 25200 32332 25212 32388
rect 25268 32332 25280 32388
rect 25200 32068 25280 32332
rect 25200 32012 25212 32068
rect 25268 32012 25280 32068
rect 25200 31748 25280 32012
rect 25200 31692 25212 31748
rect 25268 31692 25280 31748
rect 25200 31428 25280 31692
rect 25200 31372 25212 31428
rect 25268 31372 25280 31428
rect 25200 31108 25280 31372
rect 25200 31052 25212 31108
rect 25268 31052 25280 31108
rect 25200 30788 25280 31052
rect 25200 30732 25212 30788
rect 25268 30732 25280 30788
rect 25200 30468 25280 30732
rect 25200 30412 25212 30468
rect 25268 30412 25280 30468
rect 25200 30400 25280 30412
rect 25360 32388 25440 32400
rect 25360 32332 25372 32388
rect 25428 32332 25440 32388
rect 25360 32068 25440 32332
rect 25360 32012 25372 32068
rect 25428 32012 25440 32068
rect 25360 31748 25440 32012
rect 25360 31692 25372 31748
rect 25428 31692 25440 31748
rect 25360 31428 25440 31692
rect 25360 31372 25372 31428
rect 25428 31372 25440 31428
rect 25360 31108 25440 31372
rect 25360 31052 25372 31108
rect 25428 31052 25440 31108
rect 25360 30788 25440 31052
rect 25360 30732 25372 30788
rect 25428 30732 25440 30788
rect 25360 30468 25440 30732
rect 25360 30412 25372 30468
rect 25428 30412 25440 30468
rect 25360 30400 25440 30412
rect 25520 32388 25600 32400
rect 25520 32332 25532 32388
rect 25588 32332 25600 32388
rect 25520 32068 25600 32332
rect 25520 32012 25532 32068
rect 25588 32012 25600 32068
rect 25520 31748 25600 32012
rect 25520 31692 25532 31748
rect 25588 31692 25600 31748
rect 25520 31428 25600 31692
rect 25520 31372 25532 31428
rect 25588 31372 25600 31428
rect 25520 31108 25600 31372
rect 25520 31052 25532 31108
rect 25588 31052 25600 31108
rect 25520 30788 25600 31052
rect 25520 30732 25532 30788
rect 25588 30732 25600 30788
rect 25520 30468 25600 30732
rect 25520 30412 25532 30468
rect 25588 30412 25600 30468
rect 25520 30400 25600 30412
rect 25680 32388 25760 32400
rect 25680 32332 25692 32388
rect 25748 32332 25760 32388
rect 25680 32068 25760 32332
rect 25680 32012 25692 32068
rect 25748 32012 25760 32068
rect 25680 31748 25760 32012
rect 25680 31692 25692 31748
rect 25748 31692 25760 31748
rect 25680 31428 25760 31692
rect 25680 31372 25692 31428
rect 25748 31372 25760 31428
rect 25680 31108 25760 31372
rect 25680 31052 25692 31108
rect 25748 31052 25760 31108
rect 25680 30788 25760 31052
rect 25680 30732 25692 30788
rect 25748 30732 25760 30788
rect 25680 30468 25760 30732
rect 25680 30412 25692 30468
rect 25748 30412 25760 30468
rect 25680 30400 25760 30412
rect 25840 32388 25920 32400
rect 25840 32332 25852 32388
rect 25908 32332 25920 32388
rect 25840 32068 25920 32332
rect 25840 32012 25852 32068
rect 25908 32012 25920 32068
rect 25840 31748 25920 32012
rect 25840 31692 25852 31748
rect 25908 31692 25920 31748
rect 25840 31428 25920 31692
rect 25840 31372 25852 31428
rect 25908 31372 25920 31428
rect 25840 31108 25920 31372
rect 25840 31052 25852 31108
rect 25908 31052 25920 31108
rect 25840 30788 25920 31052
rect 25840 30732 25852 30788
rect 25908 30732 25920 30788
rect 25840 30468 25920 30732
rect 25840 30412 25852 30468
rect 25908 30412 25920 30468
rect 25840 30400 25920 30412
rect 26000 32388 26080 32400
rect 26000 32332 26012 32388
rect 26068 32332 26080 32388
rect 26000 32068 26080 32332
rect 26000 32012 26012 32068
rect 26068 32012 26080 32068
rect 26000 31748 26080 32012
rect 26000 31692 26012 31748
rect 26068 31692 26080 31748
rect 26000 31428 26080 31692
rect 26000 31372 26012 31428
rect 26068 31372 26080 31428
rect 26000 31108 26080 31372
rect 26000 31052 26012 31108
rect 26068 31052 26080 31108
rect 26000 30788 26080 31052
rect 26000 30732 26012 30788
rect 26068 30732 26080 30788
rect 26000 30468 26080 30732
rect 26000 30412 26012 30468
rect 26068 30412 26080 30468
rect 26000 30400 26080 30412
rect 26160 32388 26240 32400
rect 26160 32332 26172 32388
rect 26228 32332 26240 32388
rect 26160 32068 26240 32332
rect 26160 32012 26172 32068
rect 26228 32012 26240 32068
rect 26160 31748 26240 32012
rect 26160 31692 26172 31748
rect 26228 31692 26240 31748
rect 26160 31428 26240 31692
rect 26160 31372 26172 31428
rect 26228 31372 26240 31428
rect 26160 31108 26240 31372
rect 26160 31052 26172 31108
rect 26228 31052 26240 31108
rect 26160 30788 26240 31052
rect 26160 30732 26172 30788
rect 26228 30732 26240 30788
rect 26160 30468 26240 30732
rect 26160 30412 26172 30468
rect 26228 30412 26240 30468
rect 26160 30400 26240 30412
rect 26320 32388 26400 32400
rect 26320 32332 26332 32388
rect 26388 32332 26400 32388
rect 26320 32068 26400 32332
rect 26320 32012 26332 32068
rect 26388 32012 26400 32068
rect 26320 31748 26400 32012
rect 26320 31692 26332 31748
rect 26388 31692 26400 31748
rect 26320 31428 26400 31692
rect 26320 31372 26332 31428
rect 26388 31372 26400 31428
rect 26320 31108 26400 31372
rect 26320 31052 26332 31108
rect 26388 31052 26400 31108
rect 26320 30788 26400 31052
rect 26320 30732 26332 30788
rect 26388 30732 26400 30788
rect 26320 30468 26400 30732
rect 26320 30412 26332 30468
rect 26388 30412 26400 30468
rect 26320 30400 26400 30412
rect 26480 32388 26560 32400
rect 26480 32332 26492 32388
rect 26548 32332 26560 32388
rect 26480 32068 26560 32332
rect 26480 32012 26492 32068
rect 26548 32012 26560 32068
rect 26480 31748 26560 32012
rect 26480 31692 26492 31748
rect 26548 31692 26560 31748
rect 26480 31428 26560 31692
rect 26480 31372 26492 31428
rect 26548 31372 26560 31428
rect 26480 31108 26560 31372
rect 26480 31052 26492 31108
rect 26548 31052 26560 31108
rect 26480 30788 26560 31052
rect 26480 30732 26492 30788
rect 26548 30732 26560 30788
rect 26480 30468 26560 30732
rect 26480 30412 26492 30468
rect 26548 30412 26560 30468
rect 26480 30400 26560 30412
rect 26640 32388 26720 32400
rect 26640 32332 26652 32388
rect 26708 32332 26720 32388
rect 26640 32068 26720 32332
rect 26640 32012 26652 32068
rect 26708 32012 26720 32068
rect 26640 31748 26720 32012
rect 26640 31692 26652 31748
rect 26708 31692 26720 31748
rect 26640 31428 26720 31692
rect 26640 31372 26652 31428
rect 26708 31372 26720 31428
rect 26640 31108 26720 31372
rect 26640 31052 26652 31108
rect 26708 31052 26720 31108
rect 26640 30788 26720 31052
rect 26640 30732 26652 30788
rect 26708 30732 26720 30788
rect 26640 30468 26720 30732
rect 26640 30412 26652 30468
rect 26708 30412 26720 30468
rect 26640 30400 26720 30412
rect 26800 32388 26880 32400
rect 26800 32332 26812 32388
rect 26868 32332 26880 32388
rect 26800 32068 26880 32332
rect 26800 32012 26812 32068
rect 26868 32012 26880 32068
rect 26800 31748 26880 32012
rect 26800 31692 26812 31748
rect 26868 31692 26880 31748
rect 26800 31428 26880 31692
rect 26800 31372 26812 31428
rect 26868 31372 26880 31428
rect 26800 31108 26880 31372
rect 26800 31052 26812 31108
rect 26868 31052 26880 31108
rect 26800 30788 26880 31052
rect 26800 30732 26812 30788
rect 26868 30732 26880 30788
rect 26800 30468 26880 30732
rect 26800 30412 26812 30468
rect 26868 30412 26880 30468
rect 26800 30400 26880 30412
rect 26960 32388 27040 32400
rect 26960 32332 26972 32388
rect 27028 32332 27040 32388
rect 26960 32068 27040 32332
rect 26960 32012 26972 32068
rect 27028 32012 27040 32068
rect 26960 31748 27040 32012
rect 26960 31692 26972 31748
rect 27028 31692 27040 31748
rect 26960 31428 27040 31692
rect 26960 31372 26972 31428
rect 27028 31372 27040 31428
rect 26960 31108 27040 31372
rect 26960 31052 26972 31108
rect 27028 31052 27040 31108
rect 26960 30788 27040 31052
rect 26960 30732 26972 30788
rect 27028 30732 27040 30788
rect 26960 30468 27040 30732
rect 26960 30412 26972 30468
rect 27028 30412 27040 30468
rect 26960 30400 27040 30412
rect 27120 32388 27200 32400
rect 27120 32332 27132 32388
rect 27188 32332 27200 32388
rect 27120 32068 27200 32332
rect 27120 32012 27132 32068
rect 27188 32012 27200 32068
rect 27120 31748 27200 32012
rect 27120 31692 27132 31748
rect 27188 31692 27200 31748
rect 27120 31428 27200 31692
rect 27120 31372 27132 31428
rect 27188 31372 27200 31428
rect 27120 31108 27200 31372
rect 27120 31052 27132 31108
rect 27188 31052 27200 31108
rect 27120 30788 27200 31052
rect 27120 30732 27132 30788
rect 27188 30732 27200 30788
rect 27120 30468 27200 30732
rect 27120 30412 27132 30468
rect 27188 30412 27200 30468
rect 27120 30400 27200 30412
rect 27280 32388 27360 32400
rect 27280 32332 27292 32388
rect 27348 32332 27360 32388
rect 27280 32068 27360 32332
rect 27280 32012 27292 32068
rect 27348 32012 27360 32068
rect 27280 31748 27360 32012
rect 27280 31692 27292 31748
rect 27348 31692 27360 31748
rect 27280 31428 27360 31692
rect 27280 31372 27292 31428
rect 27348 31372 27360 31428
rect 27280 31108 27360 31372
rect 27280 31052 27292 31108
rect 27348 31052 27360 31108
rect 27280 30788 27360 31052
rect 27280 30732 27292 30788
rect 27348 30732 27360 30788
rect 27280 30468 27360 30732
rect 27280 30412 27292 30468
rect 27348 30412 27360 30468
rect 27280 30400 27360 30412
rect 27440 32388 27520 32400
rect 27440 32332 27452 32388
rect 27508 32332 27520 32388
rect 27440 32068 27520 32332
rect 27440 32012 27452 32068
rect 27508 32012 27520 32068
rect 27440 31748 27520 32012
rect 27440 31692 27452 31748
rect 27508 31692 27520 31748
rect 27440 31428 27520 31692
rect 27440 31372 27452 31428
rect 27508 31372 27520 31428
rect 27440 31108 27520 31372
rect 27440 31052 27452 31108
rect 27508 31052 27520 31108
rect 27440 30788 27520 31052
rect 27440 30732 27452 30788
rect 27508 30732 27520 30788
rect 27440 30468 27520 30732
rect 27440 30412 27452 30468
rect 27508 30412 27520 30468
rect 27440 30400 27520 30412
rect 27600 32388 27680 32400
rect 27600 32332 27612 32388
rect 27668 32332 27680 32388
rect 27600 32068 27680 32332
rect 27600 32012 27612 32068
rect 27668 32012 27680 32068
rect 27600 31748 27680 32012
rect 27600 31692 27612 31748
rect 27668 31692 27680 31748
rect 27600 31428 27680 31692
rect 27600 31372 27612 31428
rect 27668 31372 27680 31428
rect 27600 31108 27680 31372
rect 27600 31052 27612 31108
rect 27668 31052 27680 31108
rect 27600 30788 27680 31052
rect 27600 30732 27612 30788
rect 27668 30732 27680 30788
rect 27600 30468 27680 30732
rect 27600 30412 27612 30468
rect 27668 30412 27680 30468
rect 27600 30400 27680 30412
rect 27760 32388 27840 32400
rect 27760 32332 27772 32388
rect 27828 32332 27840 32388
rect 27760 32068 27840 32332
rect 27760 32012 27772 32068
rect 27828 32012 27840 32068
rect 27760 31748 27840 32012
rect 27760 31692 27772 31748
rect 27828 31692 27840 31748
rect 27760 31428 27840 31692
rect 27760 31372 27772 31428
rect 27828 31372 27840 31428
rect 27760 31108 27840 31372
rect 27760 31052 27772 31108
rect 27828 31052 27840 31108
rect 27760 30788 27840 31052
rect 27760 30732 27772 30788
rect 27828 30732 27840 30788
rect 27760 30468 27840 30732
rect 27760 30412 27772 30468
rect 27828 30412 27840 30468
rect 27760 30400 27840 30412
rect 27920 32388 28000 32400
rect 27920 32332 27932 32388
rect 27988 32332 28000 32388
rect 27920 32068 28000 32332
rect 27920 32012 27932 32068
rect 27988 32012 28000 32068
rect 27920 31748 28000 32012
rect 27920 31692 27932 31748
rect 27988 31692 28000 31748
rect 27920 31428 28000 31692
rect 27920 31372 27932 31428
rect 27988 31372 28000 31428
rect 27920 31108 28000 31372
rect 27920 31052 27932 31108
rect 27988 31052 28000 31108
rect 27920 30788 28000 31052
rect 27920 30732 27932 30788
rect 27988 30732 28000 30788
rect 27920 30468 28000 30732
rect 27920 30412 27932 30468
rect 27988 30412 28000 30468
rect 27920 30400 28000 30412
rect 28080 32388 28160 32400
rect 28080 32332 28092 32388
rect 28148 32332 28160 32388
rect 28080 32068 28160 32332
rect 28080 32012 28092 32068
rect 28148 32012 28160 32068
rect 28080 31748 28160 32012
rect 28080 31692 28092 31748
rect 28148 31692 28160 31748
rect 28080 31428 28160 31692
rect 28080 31372 28092 31428
rect 28148 31372 28160 31428
rect 28080 31108 28160 31372
rect 28080 31052 28092 31108
rect 28148 31052 28160 31108
rect 28080 30788 28160 31052
rect 28080 30732 28092 30788
rect 28148 30732 28160 30788
rect 28080 30468 28160 30732
rect 28080 30412 28092 30468
rect 28148 30412 28160 30468
rect 28080 30400 28160 30412
rect 28240 32388 28320 32400
rect 28240 32332 28252 32388
rect 28308 32332 28320 32388
rect 28240 32068 28320 32332
rect 28240 32012 28252 32068
rect 28308 32012 28320 32068
rect 28240 31748 28320 32012
rect 28240 31692 28252 31748
rect 28308 31692 28320 31748
rect 28240 31428 28320 31692
rect 28240 31372 28252 31428
rect 28308 31372 28320 31428
rect 28240 31108 28320 31372
rect 28240 31052 28252 31108
rect 28308 31052 28320 31108
rect 28240 30788 28320 31052
rect 28240 30732 28252 30788
rect 28308 30732 28320 30788
rect 28240 30468 28320 30732
rect 28240 30412 28252 30468
rect 28308 30412 28320 30468
rect 28240 30400 28320 30412
rect 28400 32388 28480 32400
rect 28400 32332 28412 32388
rect 28468 32332 28480 32388
rect 28400 32068 28480 32332
rect 28400 32012 28412 32068
rect 28468 32012 28480 32068
rect 28400 31748 28480 32012
rect 28400 31692 28412 31748
rect 28468 31692 28480 31748
rect 28400 31428 28480 31692
rect 28400 31372 28412 31428
rect 28468 31372 28480 31428
rect 28400 31108 28480 31372
rect 28400 31052 28412 31108
rect 28468 31052 28480 31108
rect 28400 30788 28480 31052
rect 28400 30732 28412 30788
rect 28468 30732 28480 30788
rect 28400 30468 28480 30732
rect 28400 30412 28412 30468
rect 28468 30412 28480 30468
rect 28400 30400 28480 30412
rect 28560 32388 28640 32400
rect 28560 32332 28572 32388
rect 28628 32332 28640 32388
rect 28560 32068 28640 32332
rect 28560 32012 28572 32068
rect 28628 32012 28640 32068
rect 28560 31748 28640 32012
rect 28560 31692 28572 31748
rect 28628 31692 28640 31748
rect 28560 31428 28640 31692
rect 28560 31372 28572 31428
rect 28628 31372 28640 31428
rect 28560 31108 28640 31372
rect 28560 31052 28572 31108
rect 28628 31052 28640 31108
rect 28560 30788 28640 31052
rect 28560 30732 28572 30788
rect 28628 30732 28640 30788
rect 28560 30468 28640 30732
rect 28560 30412 28572 30468
rect 28628 30412 28640 30468
rect 28560 30400 28640 30412
rect 28720 32388 28800 32400
rect 28720 32332 28732 32388
rect 28788 32332 28800 32388
rect 28720 32068 28800 32332
rect 28720 32012 28732 32068
rect 28788 32012 28800 32068
rect 28720 31748 28800 32012
rect 28720 31692 28732 31748
rect 28788 31692 28800 31748
rect 28720 31428 28800 31692
rect 28720 31372 28732 31428
rect 28788 31372 28800 31428
rect 28720 31108 28800 31372
rect 28720 31052 28732 31108
rect 28788 31052 28800 31108
rect 28720 30788 28800 31052
rect 28720 30732 28732 30788
rect 28788 30732 28800 30788
rect 28720 30468 28800 30732
rect 28720 30412 28732 30468
rect 28788 30412 28800 30468
rect 28720 30400 28800 30412
rect 28880 32388 28960 32400
rect 28880 32332 28892 32388
rect 28948 32332 28960 32388
rect 28880 32068 28960 32332
rect 28880 32012 28892 32068
rect 28948 32012 28960 32068
rect 28880 31748 28960 32012
rect 28880 31692 28892 31748
rect 28948 31692 28960 31748
rect 28880 31428 28960 31692
rect 28880 31372 28892 31428
rect 28948 31372 28960 31428
rect 28880 31108 28960 31372
rect 28880 31052 28892 31108
rect 28948 31052 28960 31108
rect 28880 30788 28960 31052
rect 28880 30732 28892 30788
rect 28948 30732 28960 30788
rect 28880 30468 28960 30732
rect 28880 30412 28892 30468
rect 28948 30412 28960 30468
rect 28880 30400 28960 30412
rect 29040 32388 29120 32400
rect 29040 32332 29052 32388
rect 29108 32332 29120 32388
rect 29040 32068 29120 32332
rect 29040 32012 29052 32068
rect 29108 32012 29120 32068
rect 29040 31748 29120 32012
rect 29040 31692 29052 31748
rect 29108 31692 29120 31748
rect 29040 31428 29120 31692
rect 29040 31372 29052 31428
rect 29108 31372 29120 31428
rect 29040 31108 29120 31372
rect 29040 31052 29052 31108
rect 29108 31052 29120 31108
rect 29040 30788 29120 31052
rect 29040 30732 29052 30788
rect 29108 30732 29120 30788
rect 29040 30468 29120 30732
rect 29040 30412 29052 30468
rect 29108 30412 29120 30468
rect 29040 30400 29120 30412
rect 29200 32388 29280 32400
rect 29200 32332 29212 32388
rect 29268 32332 29280 32388
rect 29200 32068 29280 32332
rect 29200 32012 29212 32068
rect 29268 32012 29280 32068
rect 29200 31748 29280 32012
rect 29200 31692 29212 31748
rect 29268 31692 29280 31748
rect 29200 31428 29280 31692
rect 29200 31372 29212 31428
rect 29268 31372 29280 31428
rect 29200 31108 29280 31372
rect 29200 31052 29212 31108
rect 29268 31052 29280 31108
rect 29200 30788 29280 31052
rect 29200 30732 29212 30788
rect 29268 30732 29280 30788
rect 29200 30468 29280 30732
rect 29200 30412 29212 30468
rect 29268 30412 29280 30468
rect 29200 30400 29280 30412
rect 29360 32388 29440 32400
rect 29360 32332 29372 32388
rect 29428 32332 29440 32388
rect 29360 32068 29440 32332
rect 29360 32012 29372 32068
rect 29428 32012 29440 32068
rect 29360 31748 29440 32012
rect 29360 31692 29372 31748
rect 29428 31692 29440 31748
rect 29360 31428 29440 31692
rect 29360 31372 29372 31428
rect 29428 31372 29440 31428
rect 29360 31108 29440 31372
rect 29360 31052 29372 31108
rect 29428 31052 29440 31108
rect 29360 30788 29440 31052
rect 29360 30732 29372 30788
rect 29428 30732 29440 30788
rect 29360 30468 29440 30732
rect 29360 30412 29372 30468
rect 29428 30412 29440 30468
rect 29360 30400 29440 30412
rect 23120 30308 23200 30320
rect 23120 30252 23132 30308
rect 23188 30252 23200 30308
rect 23120 29988 23200 30252
rect 23120 29932 23132 29988
rect 23188 29932 23200 29988
rect 23120 29920 23200 29932
rect 23280 30308 23360 30320
rect 23280 30252 23292 30308
rect 23348 30252 23360 30308
rect 23280 29988 23360 30252
rect 23280 29932 23292 29988
rect 23348 29932 23360 29988
rect 23280 29920 23360 29932
rect 23440 30308 23520 30320
rect 23440 30252 23452 30308
rect 23508 30252 23520 30308
rect 23440 29988 23520 30252
rect 23440 29932 23452 29988
rect 23508 29932 23520 29988
rect 23440 29920 23520 29932
rect 23600 30308 23680 30320
rect 23600 30252 23612 30308
rect 23668 30252 23680 30308
rect 23600 29988 23680 30252
rect 23600 29932 23612 29988
rect 23668 29932 23680 29988
rect 23600 29920 23680 29932
rect 23760 30308 23840 30320
rect 23760 30252 23772 30308
rect 23828 30252 23840 30308
rect 23760 29988 23840 30252
rect 23760 29932 23772 29988
rect 23828 29932 23840 29988
rect 23760 29920 23840 29932
rect 23920 30308 24000 30320
rect 23920 30252 23932 30308
rect 23988 30252 24000 30308
rect 23920 29988 24000 30252
rect 23920 29932 23932 29988
rect 23988 29932 24000 29988
rect 23920 29920 24000 29932
rect 24080 30308 24160 30320
rect 24080 30252 24092 30308
rect 24148 30252 24160 30308
rect 24080 29988 24160 30252
rect 24080 29932 24092 29988
rect 24148 29932 24160 29988
rect 24080 29920 24160 29932
rect 24240 30308 24320 30320
rect 24240 30252 24252 30308
rect 24308 30252 24320 30308
rect 24240 29988 24320 30252
rect 24240 29932 24252 29988
rect 24308 29932 24320 29988
rect 24240 29920 24320 29932
rect 24400 30308 24480 30320
rect 24400 30252 24412 30308
rect 24468 30252 24480 30308
rect 24400 29988 24480 30252
rect 24400 29932 24412 29988
rect 24468 29932 24480 29988
rect 24400 29920 24480 29932
rect 24560 30308 24640 30320
rect 24560 30252 24572 30308
rect 24628 30252 24640 30308
rect 24560 29988 24640 30252
rect 24560 29932 24572 29988
rect 24628 29932 24640 29988
rect 24560 29920 24640 29932
rect 24720 30308 24800 30320
rect 24720 30252 24732 30308
rect 24788 30252 24800 30308
rect 24720 29988 24800 30252
rect 24720 29932 24732 29988
rect 24788 29932 24800 29988
rect 24720 29920 24800 29932
rect 24880 30308 24960 30320
rect 24880 30252 24892 30308
rect 24948 30252 24960 30308
rect 24880 29988 24960 30252
rect 24880 29932 24892 29988
rect 24948 29932 24960 29988
rect 24880 29920 24960 29932
rect 25040 30308 25120 30320
rect 25040 30252 25052 30308
rect 25108 30252 25120 30308
rect 25040 29988 25120 30252
rect 25040 29932 25052 29988
rect 25108 29932 25120 29988
rect 25040 29920 25120 29932
rect 25200 30308 25280 30320
rect 25200 30252 25212 30308
rect 25268 30252 25280 30308
rect 25200 29988 25280 30252
rect 25200 29932 25212 29988
rect 25268 29932 25280 29988
rect 25200 29920 25280 29932
rect 25360 30308 25440 30320
rect 25360 30252 25372 30308
rect 25428 30252 25440 30308
rect 25360 29988 25440 30252
rect 25360 29932 25372 29988
rect 25428 29932 25440 29988
rect 25360 29920 25440 29932
rect 25520 30308 25600 30320
rect 25520 30252 25532 30308
rect 25588 30252 25600 30308
rect 25520 29988 25600 30252
rect 25520 29932 25532 29988
rect 25588 29932 25600 29988
rect 25520 29920 25600 29932
rect 25680 30308 25760 30320
rect 25680 30252 25692 30308
rect 25748 30252 25760 30308
rect 25680 29988 25760 30252
rect 25680 29932 25692 29988
rect 25748 29932 25760 29988
rect 25680 29920 25760 29932
rect 25840 30308 25920 30320
rect 25840 30252 25852 30308
rect 25908 30252 25920 30308
rect 25840 29988 25920 30252
rect 25840 29932 25852 29988
rect 25908 29932 25920 29988
rect 25840 29920 25920 29932
rect 26000 30308 26080 30320
rect 26000 30252 26012 30308
rect 26068 30252 26080 30308
rect 26000 29988 26080 30252
rect 26000 29932 26012 29988
rect 26068 29932 26080 29988
rect 26000 29920 26080 29932
rect 26160 30308 26240 30320
rect 26160 30252 26172 30308
rect 26228 30252 26240 30308
rect 26160 29988 26240 30252
rect 26160 29932 26172 29988
rect 26228 29932 26240 29988
rect 26160 29920 26240 29932
rect 26320 30308 26400 30320
rect 26320 30252 26332 30308
rect 26388 30252 26400 30308
rect 26320 29988 26400 30252
rect 26320 29932 26332 29988
rect 26388 29932 26400 29988
rect 26320 29920 26400 29932
rect 26480 30308 26560 30320
rect 26480 30252 26492 30308
rect 26548 30252 26560 30308
rect 26480 29988 26560 30252
rect 26480 29932 26492 29988
rect 26548 29932 26560 29988
rect 26480 29920 26560 29932
rect 26640 30308 26720 30320
rect 26640 30252 26652 30308
rect 26708 30252 26720 30308
rect 26640 29988 26720 30252
rect 26640 29932 26652 29988
rect 26708 29932 26720 29988
rect 26640 29920 26720 29932
rect 26800 30308 26880 30320
rect 26800 30252 26812 30308
rect 26868 30252 26880 30308
rect 26800 29988 26880 30252
rect 26800 29932 26812 29988
rect 26868 29932 26880 29988
rect 26800 29920 26880 29932
rect 26960 30308 27040 30320
rect 26960 30252 26972 30308
rect 27028 30252 27040 30308
rect 26960 29988 27040 30252
rect 26960 29932 26972 29988
rect 27028 29932 27040 29988
rect 26960 29920 27040 29932
rect 27120 30308 27200 30320
rect 27120 30252 27132 30308
rect 27188 30252 27200 30308
rect 27120 29988 27200 30252
rect 27120 29932 27132 29988
rect 27188 29932 27200 29988
rect 27120 29920 27200 29932
rect 27280 30308 27360 30320
rect 27280 30252 27292 30308
rect 27348 30252 27360 30308
rect 27280 29988 27360 30252
rect 27280 29932 27292 29988
rect 27348 29932 27360 29988
rect 27280 29920 27360 29932
rect 27440 30308 27520 30320
rect 27440 30252 27452 30308
rect 27508 30252 27520 30308
rect 27440 29988 27520 30252
rect 27440 29932 27452 29988
rect 27508 29932 27520 29988
rect 27440 29920 27520 29932
rect 27600 30308 27680 30320
rect 27600 30252 27612 30308
rect 27668 30252 27680 30308
rect 27600 29988 27680 30252
rect 27600 29932 27612 29988
rect 27668 29932 27680 29988
rect 27600 29920 27680 29932
rect 27760 30308 27840 30320
rect 27760 30252 27772 30308
rect 27828 30252 27840 30308
rect 27760 29988 27840 30252
rect 27760 29932 27772 29988
rect 27828 29932 27840 29988
rect 27760 29920 27840 29932
rect 27920 30308 28000 30320
rect 27920 30252 27932 30308
rect 27988 30252 28000 30308
rect 27920 29988 28000 30252
rect 27920 29932 27932 29988
rect 27988 29932 28000 29988
rect 27920 29920 28000 29932
rect 28080 30308 28160 30320
rect 28080 30252 28092 30308
rect 28148 30252 28160 30308
rect 28080 29988 28160 30252
rect 28080 29932 28092 29988
rect 28148 29932 28160 29988
rect 28080 29920 28160 29932
rect 28240 30308 28320 30320
rect 28240 30252 28252 30308
rect 28308 30252 28320 30308
rect 28240 29988 28320 30252
rect 28240 29932 28252 29988
rect 28308 29932 28320 29988
rect 28240 29920 28320 29932
rect 28400 30308 28480 30320
rect 28400 30252 28412 30308
rect 28468 30252 28480 30308
rect 28400 29988 28480 30252
rect 28400 29932 28412 29988
rect 28468 29932 28480 29988
rect 28400 29920 28480 29932
rect 28560 30308 28640 30320
rect 28560 30252 28572 30308
rect 28628 30252 28640 30308
rect 28560 29988 28640 30252
rect 28560 29932 28572 29988
rect 28628 29932 28640 29988
rect 28560 29920 28640 29932
rect 28720 30308 28800 30320
rect 28720 30252 28732 30308
rect 28788 30252 28800 30308
rect 28720 29988 28800 30252
rect 28720 29932 28732 29988
rect 28788 29932 28800 29988
rect 28720 29920 28800 29932
rect 28880 30308 28960 30320
rect 28880 30252 28892 30308
rect 28948 30252 28960 30308
rect 28880 29988 28960 30252
rect 28880 29932 28892 29988
rect 28948 29932 28960 29988
rect 28880 29920 28960 29932
rect 29040 30308 29120 30320
rect 29040 30252 29052 30308
rect 29108 30252 29120 30308
rect 29040 29988 29120 30252
rect 29040 29932 29052 29988
rect 29108 29932 29120 29988
rect 29040 29920 29120 29932
rect 29200 30308 29280 30320
rect 29200 30252 29212 30308
rect 29268 30252 29280 30308
rect 29200 29988 29280 30252
rect 29200 29932 29212 29988
rect 29268 29932 29280 29988
rect 29200 29920 29280 29932
rect 29360 30308 29440 30320
rect 29360 30252 29372 30308
rect 29428 30252 29440 30308
rect 29360 29988 29440 30252
rect 29360 29932 29372 29988
rect 29428 29932 29440 29988
rect 29360 29920 29440 29932
rect 22880 29772 22892 29828
rect 22948 29772 22960 29828
rect 22880 29508 22960 29772
rect 22880 29452 22892 29508
rect 22948 29452 22960 29508
rect 22880 29440 22960 29452
rect 23120 29828 23200 29840
rect 23120 29772 23132 29828
rect 23188 29772 23200 29828
rect 23120 29508 23200 29772
rect 23120 29452 23132 29508
rect 23188 29452 23200 29508
rect 23120 29440 23200 29452
rect 23280 29828 23360 29840
rect 23280 29772 23292 29828
rect 23348 29772 23360 29828
rect 23280 29508 23360 29772
rect 23280 29452 23292 29508
rect 23348 29452 23360 29508
rect 23280 29440 23360 29452
rect 23440 29828 23520 29840
rect 23440 29772 23452 29828
rect 23508 29772 23520 29828
rect 23440 29508 23520 29772
rect 23440 29452 23452 29508
rect 23508 29452 23520 29508
rect 23440 29440 23520 29452
rect 23600 29828 23680 29840
rect 23600 29772 23612 29828
rect 23668 29772 23680 29828
rect 23600 29508 23680 29772
rect 23600 29452 23612 29508
rect 23668 29452 23680 29508
rect 23600 29440 23680 29452
rect 23760 29828 23840 29840
rect 23760 29772 23772 29828
rect 23828 29772 23840 29828
rect 23760 29508 23840 29772
rect 23760 29452 23772 29508
rect 23828 29452 23840 29508
rect 23760 29440 23840 29452
rect 23920 29828 24000 29840
rect 23920 29772 23932 29828
rect 23988 29772 24000 29828
rect 23920 29508 24000 29772
rect 23920 29452 23932 29508
rect 23988 29452 24000 29508
rect 23920 29440 24000 29452
rect 24080 29828 24160 29840
rect 24080 29772 24092 29828
rect 24148 29772 24160 29828
rect 24080 29508 24160 29772
rect 24080 29452 24092 29508
rect 24148 29452 24160 29508
rect 24080 29440 24160 29452
rect 24240 29828 24320 29840
rect 24240 29772 24252 29828
rect 24308 29772 24320 29828
rect 24240 29508 24320 29772
rect 24240 29452 24252 29508
rect 24308 29452 24320 29508
rect 24240 29440 24320 29452
rect 24400 29828 24480 29840
rect 24400 29772 24412 29828
rect 24468 29772 24480 29828
rect 24400 29508 24480 29772
rect 24400 29452 24412 29508
rect 24468 29452 24480 29508
rect 24400 29440 24480 29452
rect 24560 29828 24640 29840
rect 24560 29772 24572 29828
rect 24628 29772 24640 29828
rect 24560 29508 24640 29772
rect 24560 29452 24572 29508
rect 24628 29452 24640 29508
rect 24560 29440 24640 29452
rect 24720 29828 24800 29840
rect 24720 29772 24732 29828
rect 24788 29772 24800 29828
rect 24720 29508 24800 29772
rect 24720 29452 24732 29508
rect 24788 29452 24800 29508
rect 24720 29440 24800 29452
rect 24880 29828 24960 29840
rect 24880 29772 24892 29828
rect 24948 29772 24960 29828
rect 24880 29508 24960 29772
rect 24880 29452 24892 29508
rect 24948 29452 24960 29508
rect 24880 29440 24960 29452
rect 25040 29828 25120 29840
rect 25040 29772 25052 29828
rect 25108 29772 25120 29828
rect 25040 29508 25120 29772
rect 25040 29452 25052 29508
rect 25108 29452 25120 29508
rect 25040 29440 25120 29452
rect 25200 29828 25280 29840
rect 25200 29772 25212 29828
rect 25268 29772 25280 29828
rect 25200 29508 25280 29772
rect 25200 29452 25212 29508
rect 25268 29452 25280 29508
rect 25200 29440 25280 29452
rect 25360 29828 25440 29840
rect 25360 29772 25372 29828
rect 25428 29772 25440 29828
rect 25360 29508 25440 29772
rect 25360 29452 25372 29508
rect 25428 29452 25440 29508
rect 25360 29440 25440 29452
rect 25520 29828 25600 29840
rect 25520 29772 25532 29828
rect 25588 29772 25600 29828
rect 25520 29508 25600 29772
rect 25520 29452 25532 29508
rect 25588 29452 25600 29508
rect 25520 29440 25600 29452
rect 25680 29828 25760 29840
rect 25680 29772 25692 29828
rect 25748 29772 25760 29828
rect 25680 29508 25760 29772
rect 25680 29452 25692 29508
rect 25748 29452 25760 29508
rect 25680 29440 25760 29452
rect 25840 29828 25920 29840
rect 25840 29772 25852 29828
rect 25908 29772 25920 29828
rect 25840 29508 25920 29772
rect 25840 29452 25852 29508
rect 25908 29452 25920 29508
rect 25840 29440 25920 29452
rect 26000 29828 26080 29840
rect 26000 29772 26012 29828
rect 26068 29772 26080 29828
rect 26000 29508 26080 29772
rect 26000 29452 26012 29508
rect 26068 29452 26080 29508
rect 26000 29440 26080 29452
rect 26160 29828 26240 29840
rect 26160 29772 26172 29828
rect 26228 29772 26240 29828
rect 26160 29508 26240 29772
rect 26160 29452 26172 29508
rect 26228 29452 26240 29508
rect 26160 29440 26240 29452
rect 26320 29828 26400 29840
rect 26320 29772 26332 29828
rect 26388 29772 26400 29828
rect 26320 29508 26400 29772
rect 26320 29452 26332 29508
rect 26388 29452 26400 29508
rect 26320 29440 26400 29452
rect 26480 29828 26560 29840
rect 26480 29772 26492 29828
rect 26548 29772 26560 29828
rect 26480 29508 26560 29772
rect 26480 29452 26492 29508
rect 26548 29452 26560 29508
rect 26480 29440 26560 29452
rect 26640 29828 26720 29840
rect 26640 29772 26652 29828
rect 26708 29772 26720 29828
rect 26640 29508 26720 29772
rect 26640 29452 26652 29508
rect 26708 29452 26720 29508
rect 26640 29440 26720 29452
rect 26800 29828 26880 29840
rect 26800 29772 26812 29828
rect 26868 29772 26880 29828
rect 26800 29508 26880 29772
rect 26800 29452 26812 29508
rect 26868 29452 26880 29508
rect 26800 29440 26880 29452
rect 26960 29828 27040 29840
rect 26960 29772 26972 29828
rect 27028 29772 27040 29828
rect 26960 29508 27040 29772
rect 26960 29452 26972 29508
rect 27028 29452 27040 29508
rect 26960 29440 27040 29452
rect 27120 29828 27200 29840
rect 27120 29772 27132 29828
rect 27188 29772 27200 29828
rect 27120 29508 27200 29772
rect 27120 29452 27132 29508
rect 27188 29452 27200 29508
rect 27120 29440 27200 29452
rect 27280 29828 27360 29840
rect 27280 29772 27292 29828
rect 27348 29772 27360 29828
rect 27280 29508 27360 29772
rect 27280 29452 27292 29508
rect 27348 29452 27360 29508
rect 27280 29440 27360 29452
rect 27440 29828 27520 29840
rect 27440 29772 27452 29828
rect 27508 29772 27520 29828
rect 27440 29508 27520 29772
rect 27440 29452 27452 29508
rect 27508 29452 27520 29508
rect 27440 29440 27520 29452
rect 27600 29828 27680 29840
rect 27600 29772 27612 29828
rect 27668 29772 27680 29828
rect 27600 29508 27680 29772
rect 27600 29452 27612 29508
rect 27668 29452 27680 29508
rect 27600 29440 27680 29452
rect 27760 29828 27840 29840
rect 27760 29772 27772 29828
rect 27828 29772 27840 29828
rect 27760 29508 27840 29772
rect 27760 29452 27772 29508
rect 27828 29452 27840 29508
rect 27760 29440 27840 29452
rect 27920 29828 28000 29840
rect 27920 29772 27932 29828
rect 27988 29772 28000 29828
rect 27920 29508 28000 29772
rect 27920 29452 27932 29508
rect 27988 29452 28000 29508
rect 27920 29440 28000 29452
rect 28080 29828 28160 29840
rect 28080 29772 28092 29828
rect 28148 29772 28160 29828
rect 28080 29508 28160 29772
rect 28080 29452 28092 29508
rect 28148 29452 28160 29508
rect 28080 29440 28160 29452
rect 28240 29828 28320 29840
rect 28240 29772 28252 29828
rect 28308 29772 28320 29828
rect 28240 29508 28320 29772
rect 28240 29452 28252 29508
rect 28308 29452 28320 29508
rect 28240 29440 28320 29452
rect 28400 29828 28480 29840
rect 28400 29772 28412 29828
rect 28468 29772 28480 29828
rect 28400 29508 28480 29772
rect 28400 29452 28412 29508
rect 28468 29452 28480 29508
rect 28400 29440 28480 29452
rect 28560 29828 28640 29840
rect 28560 29772 28572 29828
rect 28628 29772 28640 29828
rect 28560 29508 28640 29772
rect 28560 29452 28572 29508
rect 28628 29452 28640 29508
rect 28560 29440 28640 29452
rect 28720 29828 28800 29840
rect 28720 29772 28732 29828
rect 28788 29772 28800 29828
rect 28720 29508 28800 29772
rect 28720 29452 28732 29508
rect 28788 29452 28800 29508
rect 28720 29440 28800 29452
rect 28880 29828 28960 29840
rect 28880 29772 28892 29828
rect 28948 29772 28960 29828
rect 28880 29508 28960 29772
rect 28880 29452 28892 29508
rect 28948 29452 28960 29508
rect 28880 29440 28960 29452
rect 29040 29828 29120 29840
rect 29040 29772 29052 29828
rect 29108 29772 29120 29828
rect 29040 29508 29120 29772
rect 29040 29452 29052 29508
rect 29108 29452 29120 29508
rect 29040 29440 29120 29452
rect 29200 29828 29280 29840
rect 29200 29772 29212 29828
rect 29268 29772 29280 29828
rect 29200 29508 29280 29772
rect 29200 29452 29212 29508
rect 29268 29452 29280 29508
rect 29200 29440 29280 29452
rect 29360 29828 29440 29840
rect 29360 29772 29372 29828
rect 29428 29772 29440 29828
rect 29360 29508 29440 29772
rect 29360 29452 29372 29508
rect 29428 29452 29440 29508
rect 29360 29440 29440 29452
rect 29520 29828 29600 33360
rect 29520 29772 29532 29828
rect 29588 29772 29600 29828
rect 29520 29508 29600 29772
rect 29520 29452 29532 29508
rect 29588 29452 29600 29508
rect 29520 29360 29600 29452
rect 29680 29668 29760 33360
rect 29680 29612 29692 29668
rect 29748 29612 29760 29668
rect 29680 29360 29760 29612
rect 29840 29828 29920 33360
rect 29840 29772 29852 29828
rect 29908 29772 29920 29828
rect 29840 29508 29920 29772
rect 29840 29452 29852 29508
rect 29908 29452 29920 29508
rect 29840 29360 29920 29452
rect 30000 30308 30080 33360
rect 30000 30252 30012 30308
rect 30068 30252 30080 30308
rect 30000 29988 30080 30252
rect 30000 29932 30012 29988
rect 30068 29932 30080 29988
rect 30000 29360 30080 29932
rect 30160 30148 30240 33360
rect 30160 30092 30172 30148
rect 30228 30092 30240 30148
rect 30160 29360 30240 30092
rect 30320 30308 30400 33360
rect 30320 30252 30332 30308
rect 30388 30252 30400 30308
rect 30320 29988 30400 30252
rect 30320 29932 30332 29988
rect 30388 29932 30400 29988
rect 30320 29360 30400 29932
rect 30480 32388 30560 33360
rect 30480 32332 30492 32388
rect 30548 32332 30560 32388
rect 30480 32068 30560 32332
rect 30480 32012 30492 32068
rect 30548 32012 30560 32068
rect 30480 31748 30560 32012
rect 30480 31692 30492 31748
rect 30548 31692 30560 31748
rect 30480 31428 30560 31692
rect 30480 31372 30492 31428
rect 30548 31372 30560 31428
rect 30480 31108 30560 31372
rect 30480 31052 30492 31108
rect 30548 31052 30560 31108
rect 30480 30788 30560 31052
rect 30480 30732 30492 30788
rect 30548 30732 30560 30788
rect 30480 30468 30560 30732
rect 30480 30412 30492 30468
rect 30548 30412 30560 30468
rect 30480 29360 30560 30412
rect 30640 30628 30720 33360
rect 30640 30572 30652 30628
rect 30708 30572 30720 30628
rect 30640 29360 30720 30572
rect 30800 32388 30880 33360
rect 30800 32332 30812 32388
rect 30868 32332 30880 32388
rect 30800 32068 30880 32332
rect 30800 32012 30812 32068
rect 30868 32012 30880 32068
rect 30800 31748 30880 32012
rect 30800 31692 30812 31748
rect 30868 31692 30880 31748
rect 30800 31428 30880 31692
rect 30800 31372 30812 31428
rect 30868 31372 30880 31428
rect 30800 31108 30880 31372
rect 30800 31052 30812 31108
rect 30868 31052 30880 31108
rect 30800 30788 30880 31052
rect 30800 30732 30812 30788
rect 30868 30732 30880 30788
rect 30800 30468 30880 30732
rect 30800 30412 30812 30468
rect 30868 30412 30880 30468
rect 30800 29360 30880 30412
rect 30960 30948 31040 33360
rect 30960 30892 30972 30948
rect 31028 30892 31040 30948
rect 30960 29360 31040 30892
rect 31120 32388 31200 33360
rect 31120 32332 31132 32388
rect 31188 32332 31200 32388
rect 31120 32068 31200 32332
rect 31120 32012 31132 32068
rect 31188 32012 31200 32068
rect 31120 31748 31200 32012
rect 31120 31692 31132 31748
rect 31188 31692 31200 31748
rect 31120 31428 31200 31692
rect 31120 31372 31132 31428
rect 31188 31372 31200 31428
rect 31120 31108 31200 31372
rect 31120 31052 31132 31108
rect 31188 31052 31200 31108
rect 31120 30788 31200 31052
rect 31120 30732 31132 30788
rect 31188 30732 31200 30788
rect 31120 30468 31200 30732
rect 31120 30412 31132 30468
rect 31188 30412 31200 30468
rect 31120 29360 31200 30412
rect 31280 31268 31360 33360
rect 31280 31212 31292 31268
rect 31348 31212 31360 31268
rect 31280 29360 31360 31212
rect 31440 32388 31520 33360
rect 31440 32332 31452 32388
rect 31508 32332 31520 32388
rect 31440 32068 31520 32332
rect 31440 32012 31452 32068
rect 31508 32012 31520 32068
rect 31440 31748 31520 32012
rect 31440 31692 31452 31748
rect 31508 31692 31520 31748
rect 31440 31428 31520 31692
rect 31440 31372 31452 31428
rect 31508 31372 31520 31428
rect 31440 31108 31520 31372
rect 31440 31052 31452 31108
rect 31508 31052 31520 31108
rect 31440 30788 31520 31052
rect 31440 30732 31452 30788
rect 31508 30732 31520 30788
rect 31440 30468 31520 30732
rect 31440 30412 31452 30468
rect 31508 30412 31520 30468
rect 31440 29360 31520 30412
rect 31600 31588 31680 33360
rect 31600 31532 31612 31588
rect 31668 31532 31680 31588
rect 31600 29360 31680 31532
rect 31760 32388 31840 33360
rect 31760 32332 31772 32388
rect 31828 32332 31840 32388
rect 31760 32068 31840 32332
rect 31760 32012 31772 32068
rect 31828 32012 31840 32068
rect 31760 31748 31840 32012
rect 31760 31692 31772 31748
rect 31828 31692 31840 31748
rect 31760 31428 31840 31692
rect 31760 31372 31772 31428
rect 31828 31372 31840 31428
rect 31760 31108 31840 31372
rect 31760 31052 31772 31108
rect 31828 31052 31840 31108
rect 31760 30788 31840 31052
rect 31760 30732 31772 30788
rect 31828 30732 31840 30788
rect 31760 30468 31840 30732
rect 31760 30412 31772 30468
rect 31828 30412 31840 30468
rect 31760 29360 31840 30412
rect 31920 31908 32000 33360
rect 31920 31852 31932 31908
rect 31988 31852 32000 31908
rect 31920 29360 32000 31852
rect 32080 32388 32160 33360
rect 32080 32332 32092 32388
rect 32148 32332 32160 32388
rect 32080 32068 32160 32332
rect 32080 32012 32092 32068
rect 32148 32012 32160 32068
rect 32080 31748 32160 32012
rect 32080 31692 32092 31748
rect 32148 31692 32160 31748
rect 32080 31428 32160 31692
rect 32080 31372 32092 31428
rect 32148 31372 32160 31428
rect 32080 31108 32160 31372
rect 32080 31052 32092 31108
rect 32148 31052 32160 31108
rect 32080 30788 32160 31052
rect 32080 30732 32092 30788
rect 32148 30732 32160 30788
rect 32080 30468 32160 30732
rect 32080 30412 32092 30468
rect 32148 30412 32160 30468
rect 32080 29360 32160 30412
rect 32240 32228 32320 33360
rect 32240 32172 32252 32228
rect 32308 32172 32320 32228
rect 32240 29360 32320 32172
rect 32400 32388 32480 33360
rect 32400 32332 32412 32388
rect 32468 32332 32480 32388
rect 32400 32068 32480 32332
rect 32400 32012 32412 32068
rect 32468 32012 32480 32068
rect 32400 31748 32480 32012
rect 32400 31692 32412 31748
rect 32468 31692 32480 31748
rect 32400 31428 32480 31692
rect 32400 31372 32412 31428
rect 32468 31372 32480 31428
rect 32400 31108 32480 31372
rect 32400 31052 32412 31108
rect 32468 31052 32480 31108
rect 32400 30788 32480 31052
rect 32400 30732 32412 30788
rect 32468 30732 32480 30788
rect 32400 30468 32480 30732
rect 32400 30412 32412 30468
rect 32468 30412 32480 30468
rect 32400 29360 32480 30412
rect 32560 32868 32640 33360
rect 32560 32812 32572 32868
rect 32628 32812 32640 32868
rect 32560 32548 32640 32812
rect 32560 32492 32572 32548
rect 32628 32492 32640 32548
rect 32560 29360 32640 32492
rect 32720 32708 32800 33360
rect 32720 32652 32732 32708
rect 32788 32652 32800 32708
rect 32720 29360 32800 32652
rect 32880 32868 32960 33360
rect 32880 32812 32892 32868
rect 32948 32812 32960 32868
rect 32880 32548 32960 32812
rect 32880 32492 32892 32548
rect 32948 32492 32960 32548
rect 32880 29360 32960 32492
rect 33040 33348 33120 33360
rect 33040 33292 33052 33348
rect 33108 33292 33120 33348
rect 33040 33028 33120 33292
rect 33040 32972 33052 33028
rect 33108 32972 33120 33028
rect 33040 29360 33120 32972
rect 33200 33188 33280 33360
rect 33200 33132 33212 33188
rect 33268 33132 33280 33188
rect 33200 29360 33280 33132
rect 33360 33348 33440 33360
rect 33360 33292 33372 33348
rect 33428 33292 33440 33348
rect 33360 33028 33440 33292
rect 33360 32972 33372 33028
rect 33428 32972 33440 33028
rect 33360 29360 33440 32972
rect 33520 33348 33600 33360
rect 33520 33292 33532 33348
rect 33588 33292 33600 33348
rect 33520 33028 33600 33292
rect 33520 32972 33532 33028
rect 33588 32972 33600 33028
rect 33520 32960 33600 32972
rect 33680 33348 33760 33360
rect 33680 33292 33692 33348
rect 33748 33292 33760 33348
rect 33680 33028 33760 33292
rect 33680 32972 33692 33028
rect 33748 32972 33760 33028
rect 33680 32960 33760 32972
rect 33840 33348 33920 33360
rect 33840 33292 33852 33348
rect 33908 33292 33920 33348
rect 33840 33028 33920 33292
rect 33840 32972 33852 33028
rect 33908 32972 33920 33028
rect 33840 32960 33920 32972
rect 34000 33348 34080 33360
rect 34000 33292 34012 33348
rect 34068 33292 34080 33348
rect 34000 33028 34080 33292
rect 34000 32972 34012 33028
rect 34068 32972 34080 33028
rect 34000 32960 34080 32972
rect 34160 33348 34240 33360
rect 34160 33292 34172 33348
rect 34228 33292 34240 33348
rect 34160 33028 34240 33292
rect 34160 32972 34172 33028
rect 34228 32972 34240 33028
rect 34160 32960 34240 32972
rect 34320 33348 34400 33360
rect 34320 33292 34332 33348
rect 34388 33292 34400 33348
rect 34320 33028 34400 33292
rect 34320 32972 34332 33028
rect 34388 32972 34400 33028
rect 34320 32960 34400 32972
rect 34480 33348 34560 33360
rect 34480 33292 34492 33348
rect 34548 33292 34560 33348
rect 34480 33028 34560 33292
rect 34480 32972 34492 33028
rect 34548 32972 34560 33028
rect 34480 32960 34560 32972
rect 34640 33348 34720 33360
rect 34640 33292 34652 33348
rect 34708 33292 34720 33348
rect 34640 33028 34720 33292
rect 34640 32972 34652 33028
rect 34708 32972 34720 33028
rect 34640 32960 34720 32972
rect 34800 33348 34880 33360
rect 34800 33292 34812 33348
rect 34868 33292 34880 33348
rect 34800 33028 34880 33292
rect 34800 32972 34812 33028
rect 34868 32972 34880 33028
rect 34800 32960 34880 32972
rect 34960 33348 35040 33360
rect 34960 33292 34972 33348
rect 35028 33292 35040 33348
rect 34960 33028 35040 33292
rect 34960 32972 34972 33028
rect 35028 32972 35040 33028
rect 34960 32960 35040 32972
rect 35120 33348 35200 33360
rect 35120 33292 35132 33348
rect 35188 33292 35200 33348
rect 35120 33028 35200 33292
rect 35120 32972 35132 33028
rect 35188 32972 35200 33028
rect 35120 32960 35200 32972
rect 35280 33348 35360 33360
rect 35280 33292 35292 33348
rect 35348 33292 35360 33348
rect 35280 33028 35360 33292
rect 35280 32972 35292 33028
rect 35348 32972 35360 33028
rect 35280 32960 35360 32972
rect 35440 33348 35520 33360
rect 35440 33292 35452 33348
rect 35508 33292 35520 33348
rect 35440 33028 35520 33292
rect 35440 32972 35452 33028
rect 35508 32972 35520 33028
rect 35440 32960 35520 32972
rect 35600 33348 35680 33360
rect 35600 33292 35612 33348
rect 35668 33292 35680 33348
rect 35600 33028 35680 33292
rect 35600 32972 35612 33028
rect 35668 32972 35680 33028
rect 35600 32960 35680 32972
rect 35760 33348 35840 33360
rect 35760 33292 35772 33348
rect 35828 33292 35840 33348
rect 35760 33028 35840 33292
rect 35760 32972 35772 33028
rect 35828 32972 35840 33028
rect 35760 32960 35840 32972
rect 35920 33348 36000 33360
rect 35920 33292 35932 33348
rect 35988 33292 36000 33348
rect 35920 33028 36000 33292
rect 35920 32972 35932 33028
rect 35988 32972 36000 33028
rect 35920 32960 36000 32972
rect 36080 33348 36160 33360
rect 36080 33292 36092 33348
rect 36148 33292 36160 33348
rect 36080 33028 36160 33292
rect 36080 32972 36092 33028
rect 36148 32972 36160 33028
rect 36080 32960 36160 32972
rect 36240 33348 36320 33360
rect 36240 33292 36252 33348
rect 36308 33292 36320 33348
rect 36240 33028 36320 33292
rect 36240 32972 36252 33028
rect 36308 32972 36320 33028
rect 36240 32960 36320 32972
rect 36400 33348 36480 33360
rect 36400 33292 36412 33348
rect 36468 33292 36480 33348
rect 36400 33028 36480 33292
rect 36400 32972 36412 33028
rect 36468 32972 36480 33028
rect 36400 32960 36480 32972
rect 36560 33348 36640 33360
rect 36560 33292 36572 33348
rect 36628 33292 36640 33348
rect 36560 33028 36640 33292
rect 36560 32972 36572 33028
rect 36628 32972 36640 33028
rect 36560 32960 36640 32972
rect 36720 33348 36800 33360
rect 36720 33292 36732 33348
rect 36788 33292 36800 33348
rect 36720 33028 36800 33292
rect 36720 32972 36732 33028
rect 36788 32972 36800 33028
rect 36720 32960 36800 32972
rect 36880 33348 36960 33360
rect 36880 33292 36892 33348
rect 36948 33292 36960 33348
rect 36880 33028 36960 33292
rect 36880 32972 36892 33028
rect 36948 32972 36960 33028
rect 36880 32960 36960 32972
rect 37040 33348 37120 33360
rect 37040 33292 37052 33348
rect 37108 33292 37120 33348
rect 37040 33028 37120 33292
rect 37040 32972 37052 33028
rect 37108 32972 37120 33028
rect 37040 32960 37120 32972
rect 37200 33348 37280 33360
rect 37200 33292 37212 33348
rect 37268 33292 37280 33348
rect 37200 33028 37280 33292
rect 37200 32972 37212 33028
rect 37268 32972 37280 33028
rect 37200 32960 37280 32972
rect 37360 33348 37440 33360
rect 37360 33292 37372 33348
rect 37428 33292 37440 33348
rect 37360 33028 37440 33292
rect 37360 32972 37372 33028
rect 37428 32972 37440 33028
rect 37360 32960 37440 32972
rect 37520 33348 37600 33360
rect 37520 33292 37532 33348
rect 37588 33292 37600 33348
rect 37520 33028 37600 33292
rect 37520 32972 37532 33028
rect 37588 32972 37600 33028
rect 37520 32960 37600 32972
rect 37680 33348 37760 33360
rect 37680 33292 37692 33348
rect 37748 33292 37760 33348
rect 37680 33028 37760 33292
rect 37680 32972 37692 33028
rect 37748 32972 37760 33028
rect 37680 32960 37760 32972
rect 37840 33348 37920 33360
rect 37840 33292 37852 33348
rect 37908 33292 37920 33348
rect 37840 33028 37920 33292
rect 37840 32972 37852 33028
rect 37908 32972 37920 33028
rect 37840 32960 37920 32972
rect 38000 33348 38080 33360
rect 38000 33292 38012 33348
rect 38068 33292 38080 33348
rect 38000 33028 38080 33292
rect 38000 32972 38012 33028
rect 38068 32972 38080 33028
rect 38000 32960 38080 32972
rect 38160 33348 38240 33360
rect 38160 33292 38172 33348
rect 38228 33292 38240 33348
rect 38160 33028 38240 33292
rect 38160 32972 38172 33028
rect 38228 32972 38240 33028
rect 38160 32960 38240 32972
rect 38320 33348 38400 33360
rect 38320 33292 38332 33348
rect 38388 33292 38400 33348
rect 38320 33028 38400 33292
rect 38320 32972 38332 33028
rect 38388 32972 38400 33028
rect 38320 32960 38400 32972
rect 38480 33348 38560 33360
rect 38480 33292 38492 33348
rect 38548 33292 38560 33348
rect 38480 33028 38560 33292
rect 38480 32972 38492 33028
rect 38548 32972 38560 33028
rect 38480 32960 38560 32972
rect 38640 33348 38720 33360
rect 38640 33292 38652 33348
rect 38708 33292 38720 33348
rect 38640 33028 38720 33292
rect 38640 32972 38652 33028
rect 38708 32972 38720 33028
rect 38640 32960 38720 32972
rect 38800 33348 38880 33360
rect 38800 33292 38812 33348
rect 38868 33292 38880 33348
rect 38800 33028 38880 33292
rect 38800 32972 38812 33028
rect 38868 32972 38880 33028
rect 38800 32960 38880 32972
rect 38960 33348 39040 33360
rect 38960 33292 38972 33348
rect 39028 33292 39040 33348
rect 38960 33028 39040 33292
rect 38960 32972 38972 33028
rect 39028 32972 39040 33028
rect 38960 32960 39040 32972
rect 39120 33348 39200 33360
rect 39120 33292 39132 33348
rect 39188 33292 39200 33348
rect 39120 33028 39200 33292
rect 39120 32972 39132 33028
rect 39188 32972 39200 33028
rect 39120 32960 39200 32972
rect 39280 33348 39360 33360
rect 39280 33292 39292 33348
rect 39348 33292 39360 33348
rect 39280 33028 39360 33292
rect 39280 32972 39292 33028
rect 39348 32972 39360 33028
rect 39280 32960 39360 32972
rect 39440 33348 39520 33360
rect 39440 33292 39452 33348
rect 39508 33292 39520 33348
rect 39440 33028 39520 33292
rect 39440 32972 39452 33028
rect 39508 32972 39520 33028
rect 39440 32960 39520 32972
rect 39600 33348 39680 33360
rect 39600 33292 39612 33348
rect 39668 33292 39680 33348
rect 39600 33028 39680 33292
rect 39600 32972 39612 33028
rect 39668 32972 39680 33028
rect 39600 32960 39680 32972
rect 39760 33348 39840 33360
rect 39760 33292 39772 33348
rect 39828 33292 39840 33348
rect 39760 33028 39840 33292
rect 39760 32972 39772 33028
rect 39828 32972 39840 33028
rect 39760 32960 39840 32972
rect 39920 33348 40000 33360
rect 39920 33292 39932 33348
rect 39988 33292 40000 33348
rect 39920 33028 40000 33292
rect 39920 32972 39932 33028
rect 39988 32972 40000 33028
rect 39920 32960 40000 32972
rect 40080 33348 40160 33360
rect 40080 33292 40092 33348
rect 40148 33292 40160 33348
rect 40080 33028 40160 33292
rect 40080 32972 40092 33028
rect 40148 32972 40160 33028
rect 40080 32960 40160 32972
rect 40240 33348 40320 33360
rect 40240 33292 40252 33348
rect 40308 33292 40320 33348
rect 40240 33028 40320 33292
rect 40240 32972 40252 33028
rect 40308 32972 40320 33028
rect 40240 32960 40320 32972
rect 40400 33348 40480 33360
rect 40400 33292 40412 33348
rect 40468 33292 40480 33348
rect 40400 33028 40480 33292
rect 40400 32972 40412 33028
rect 40468 32972 40480 33028
rect 40400 32960 40480 32972
rect 40560 33348 40640 33360
rect 40560 33292 40572 33348
rect 40628 33292 40640 33348
rect 40560 33028 40640 33292
rect 40560 32972 40572 33028
rect 40628 32972 40640 33028
rect 40560 32960 40640 32972
rect 40720 33348 40800 33360
rect 40720 33292 40732 33348
rect 40788 33292 40800 33348
rect 40720 33028 40800 33292
rect 40720 32972 40732 33028
rect 40788 32972 40800 33028
rect 40720 32960 40800 32972
rect 40880 33348 40960 33360
rect 40880 33292 40892 33348
rect 40948 33292 40960 33348
rect 40880 33028 40960 33292
rect 40880 32972 40892 33028
rect 40948 32972 40960 33028
rect 40880 32960 40960 32972
rect 41040 33348 41120 33360
rect 41040 33292 41052 33348
rect 41108 33292 41120 33348
rect 41040 33028 41120 33292
rect 41040 32972 41052 33028
rect 41108 32972 41120 33028
rect 41040 32960 41120 32972
rect 41200 33348 41280 33360
rect 41200 33292 41212 33348
rect 41268 33292 41280 33348
rect 41200 33028 41280 33292
rect 41200 32972 41212 33028
rect 41268 32972 41280 33028
rect 41200 32960 41280 32972
rect 41360 33348 41440 33360
rect 41360 33292 41372 33348
rect 41428 33292 41440 33348
rect 41360 33028 41440 33292
rect 41360 32972 41372 33028
rect 41428 32972 41440 33028
rect 41360 32960 41440 32972
rect 41520 33348 41600 33360
rect 41520 33292 41532 33348
rect 41588 33292 41600 33348
rect 41520 33028 41600 33292
rect 41520 32972 41532 33028
rect 41588 32972 41600 33028
rect 41520 32960 41600 32972
rect 41680 33348 41760 33360
rect 41680 33292 41692 33348
rect 41748 33292 41760 33348
rect 41680 33028 41760 33292
rect 41680 32972 41692 33028
rect 41748 32972 41760 33028
rect 41680 32960 41760 32972
rect 41840 33348 41920 33360
rect 41840 33292 41852 33348
rect 41908 33292 41920 33348
rect 41840 33028 41920 33292
rect 41840 32972 41852 33028
rect 41908 32972 41920 33028
rect 41840 32960 41920 32972
rect 33520 32868 33600 32880
rect 33520 32812 33532 32868
rect 33588 32812 33600 32868
rect 33520 32548 33600 32812
rect 33520 32492 33532 32548
rect 33588 32492 33600 32548
rect 33520 32480 33600 32492
rect 33680 32868 33760 32880
rect 33680 32812 33692 32868
rect 33748 32812 33760 32868
rect 33680 32548 33760 32812
rect 33680 32492 33692 32548
rect 33748 32492 33760 32548
rect 33680 32480 33760 32492
rect 33840 32868 33920 32880
rect 33840 32812 33852 32868
rect 33908 32812 33920 32868
rect 33840 32548 33920 32812
rect 33840 32492 33852 32548
rect 33908 32492 33920 32548
rect 33840 32480 33920 32492
rect 34000 32868 34080 32880
rect 34000 32812 34012 32868
rect 34068 32812 34080 32868
rect 34000 32548 34080 32812
rect 34000 32492 34012 32548
rect 34068 32492 34080 32548
rect 34000 32480 34080 32492
rect 34160 32868 34240 32880
rect 34160 32812 34172 32868
rect 34228 32812 34240 32868
rect 34160 32548 34240 32812
rect 34160 32492 34172 32548
rect 34228 32492 34240 32548
rect 34160 32480 34240 32492
rect 34320 32868 34400 32880
rect 34320 32812 34332 32868
rect 34388 32812 34400 32868
rect 34320 32548 34400 32812
rect 34320 32492 34332 32548
rect 34388 32492 34400 32548
rect 34320 32480 34400 32492
rect 34480 32868 34560 32880
rect 34480 32812 34492 32868
rect 34548 32812 34560 32868
rect 34480 32548 34560 32812
rect 34480 32492 34492 32548
rect 34548 32492 34560 32548
rect 34480 32480 34560 32492
rect 34640 32868 34720 32880
rect 34640 32812 34652 32868
rect 34708 32812 34720 32868
rect 34640 32548 34720 32812
rect 34640 32492 34652 32548
rect 34708 32492 34720 32548
rect 34640 32480 34720 32492
rect 34800 32868 34880 32880
rect 34800 32812 34812 32868
rect 34868 32812 34880 32868
rect 34800 32548 34880 32812
rect 34800 32492 34812 32548
rect 34868 32492 34880 32548
rect 34800 32480 34880 32492
rect 34960 32868 35040 32880
rect 34960 32812 34972 32868
rect 35028 32812 35040 32868
rect 34960 32548 35040 32812
rect 34960 32492 34972 32548
rect 35028 32492 35040 32548
rect 34960 32480 35040 32492
rect 35120 32868 35200 32880
rect 35120 32812 35132 32868
rect 35188 32812 35200 32868
rect 35120 32548 35200 32812
rect 35120 32492 35132 32548
rect 35188 32492 35200 32548
rect 35120 32480 35200 32492
rect 35280 32868 35360 32880
rect 35280 32812 35292 32868
rect 35348 32812 35360 32868
rect 35280 32548 35360 32812
rect 35280 32492 35292 32548
rect 35348 32492 35360 32548
rect 35280 32480 35360 32492
rect 35440 32868 35520 32880
rect 35440 32812 35452 32868
rect 35508 32812 35520 32868
rect 35440 32548 35520 32812
rect 35440 32492 35452 32548
rect 35508 32492 35520 32548
rect 35440 32480 35520 32492
rect 35600 32868 35680 32880
rect 35600 32812 35612 32868
rect 35668 32812 35680 32868
rect 35600 32548 35680 32812
rect 35600 32492 35612 32548
rect 35668 32492 35680 32548
rect 35600 32480 35680 32492
rect 35760 32868 35840 32880
rect 35760 32812 35772 32868
rect 35828 32812 35840 32868
rect 35760 32548 35840 32812
rect 35760 32492 35772 32548
rect 35828 32492 35840 32548
rect 35760 32480 35840 32492
rect 35920 32868 36000 32880
rect 35920 32812 35932 32868
rect 35988 32812 36000 32868
rect 35920 32548 36000 32812
rect 35920 32492 35932 32548
rect 35988 32492 36000 32548
rect 35920 32480 36000 32492
rect 36080 32868 36160 32880
rect 36080 32812 36092 32868
rect 36148 32812 36160 32868
rect 36080 32548 36160 32812
rect 36080 32492 36092 32548
rect 36148 32492 36160 32548
rect 36080 32480 36160 32492
rect 36240 32868 36320 32880
rect 36240 32812 36252 32868
rect 36308 32812 36320 32868
rect 36240 32548 36320 32812
rect 36240 32492 36252 32548
rect 36308 32492 36320 32548
rect 36240 32480 36320 32492
rect 36400 32868 36480 32880
rect 36400 32812 36412 32868
rect 36468 32812 36480 32868
rect 36400 32548 36480 32812
rect 36400 32492 36412 32548
rect 36468 32492 36480 32548
rect 36400 32480 36480 32492
rect 36560 32868 36640 32880
rect 36560 32812 36572 32868
rect 36628 32812 36640 32868
rect 36560 32548 36640 32812
rect 36560 32492 36572 32548
rect 36628 32492 36640 32548
rect 36560 32480 36640 32492
rect 36720 32868 36800 32880
rect 36720 32812 36732 32868
rect 36788 32812 36800 32868
rect 36720 32548 36800 32812
rect 36720 32492 36732 32548
rect 36788 32492 36800 32548
rect 36720 32480 36800 32492
rect 36880 32868 36960 32880
rect 36880 32812 36892 32868
rect 36948 32812 36960 32868
rect 36880 32548 36960 32812
rect 36880 32492 36892 32548
rect 36948 32492 36960 32548
rect 36880 32480 36960 32492
rect 37040 32868 37120 32880
rect 37040 32812 37052 32868
rect 37108 32812 37120 32868
rect 37040 32548 37120 32812
rect 37040 32492 37052 32548
rect 37108 32492 37120 32548
rect 37040 32480 37120 32492
rect 37200 32868 37280 32880
rect 37200 32812 37212 32868
rect 37268 32812 37280 32868
rect 37200 32548 37280 32812
rect 37200 32492 37212 32548
rect 37268 32492 37280 32548
rect 37200 32480 37280 32492
rect 37360 32868 37440 32880
rect 37360 32812 37372 32868
rect 37428 32812 37440 32868
rect 37360 32548 37440 32812
rect 37360 32492 37372 32548
rect 37428 32492 37440 32548
rect 37360 32480 37440 32492
rect 37520 32868 37600 32880
rect 37520 32812 37532 32868
rect 37588 32812 37600 32868
rect 37520 32548 37600 32812
rect 37520 32492 37532 32548
rect 37588 32492 37600 32548
rect 37520 32480 37600 32492
rect 37680 32868 37760 32880
rect 37680 32812 37692 32868
rect 37748 32812 37760 32868
rect 37680 32548 37760 32812
rect 37680 32492 37692 32548
rect 37748 32492 37760 32548
rect 37680 32480 37760 32492
rect 37840 32868 37920 32880
rect 37840 32812 37852 32868
rect 37908 32812 37920 32868
rect 37840 32548 37920 32812
rect 37840 32492 37852 32548
rect 37908 32492 37920 32548
rect 37840 32480 37920 32492
rect 38000 32868 38080 32880
rect 38000 32812 38012 32868
rect 38068 32812 38080 32868
rect 38000 32548 38080 32812
rect 38000 32492 38012 32548
rect 38068 32492 38080 32548
rect 38000 32480 38080 32492
rect 38160 32868 38240 32880
rect 38160 32812 38172 32868
rect 38228 32812 38240 32868
rect 38160 32548 38240 32812
rect 38160 32492 38172 32548
rect 38228 32492 38240 32548
rect 38160 32480 38240 32492
rect 38320 32868 38400 32880
rect 38320 32812 38332 32868
rect 38388 32812 38400 32868
rect 38320 32548 38400 32812
rect 38320 32492 38332 32548
rect 38388 32492 38400 32548
rect 38320 32480 38400 32492
rect 38480 32868 38560 32880
rect 38480 32812 38492 32868
rect 38548 32812 38560 32868
rect 38480 32548 38560 32812
rect 38480 32492 38492 32548
rect 38548 32492 38560 32548
rect 38480 32480 38560 32492
rect 38640 32868 38720 32880
rect 38640 32812 38652 32868
rect 38708 32812 38720 32868
rect 38640 32548 38720 32812
rect 38640 32492 38652 32548
rect 38708 32492 38720 32548
rect 38640 32480 38720 32492
rect 38800 32868 38880 32880
rect 38800 32812 38812 32868
rect 38868 32812 38880 32868
rect 38800 32548 38880 32812
rect 38800 32492 38812 32548
rect 38868 32492 38880 32548
rect 38800 32480 38880 32492
rect 38960 32868 39040 32880
rect 38960 32812 38972 32868
rect 39028 32812 39040 32868
rect 38960 32548 39040 32812
rect 38960 32492 38972 32548
rect 39028 32492 39040 32548
rect 38960 32480 39040 32492
rect 39120 32868 39200 32880
rect 39120 32812 39132 32868
rect 39188 32812 39200 32868
rect 39120 32548 39200 32812
rect 39120 32492 39132 32548
rect 39188 32492 39200 32548
rect 39120 32480 39200 32492
rect 39280 32868 39360 32880
rect 39280 32812 39292 32868
rect 39348 32812 39360 32868
rect 39280 32548 39360 32812
rect 39280 32492 39292 32548
rect 39348 32492 39360 32548
rect 39280 32480 39360 32492
rect 39440 32868 39520 32880
rect 39440 32812 39452 32868
rect 39508 32812 39520 32868
rect 39440 32548 39520 32812
rect 39440 32492 39452 32548
rect 39508 32492 39520 32548
rect 39440 32480 39520 32492
rect 39600 32868 39680 32880
rect 39600 32812 39612 32868
rect 39668 32812 39680 32868
rect 39600 32548 39680 32812
rect 39600 32492 39612 32548
rect 39668 32492 39680 32548
rect 39600 32480 39680 32492
rect 39760 32868 39840 32880
rect 39760 32812 39772 32868
rect 39828 32812 39840 32868
rect 39760 32548 39840 32812
rect 39760 32492 39772 32548
rect 39828 32492 39840 32548
rect 39760 32480 39840 32492
rect 39920 32868 40000 32880
rect 39920 32812 39932 32868
rect 39988 32812 40000 32868
rect 39920 32548 40000 32812
rect 39920 32492 39932 32548
rect 39988 32492 40000 32548
rect 39920 32480 40000 32492
rect 40080 32868 40160 32880
rect 40080 32812 40092 32868
rect 40148 32812 40160 32868
rect 40080 32548 40160 32812
rect 40080 32492 40092 32548
rect 40148 32492 40160 32548
rect 40080 32480 40160 32492
rect 40240 32868 40320 32880
rect 40240 32812 40252 32868
rect 40308 32812 40320 32868
rect 40240 32548 40320 32812
rect 40240 32492 40252 32548
rect 40308 32492 40320 32548
rect 40240 32480 40320 32492
rect 40400 32868 40480 32880
rect 40400 32812 40412 32868
rect 40468 32812 40480 32868
rect 40400 32548 40480 32812
rect 40400 32492 40412 32548
rect 40468 32492 40480 32548
rect 40400 32480 40480 32492
rect 40560 32868 40640 32880
rect 40560 32812 40572 32868
rect 40628 32812 40640 32868
rect 40560 32548 40640 32812
rect 40560 32492 40572 32548
rect 40628 32492 40640 32548
rect 40560 32480 40640 32492
rect 40720 32868 40800 32880
rect 40720 32812 40732 32868
rect 40788 32812 40800 32868
rect 40720 32548 40800 32812
rect 40720 32492 40732 32548
rect 40788 32492 40800 32548
rect 40720 32480 40800 32492
rect 40880 32868 40960 32880
rect 40880 32812 40892 32868
rect 40948 32812 40960 32868
rect 40880 32548 40960 32812
rect 40880 32492 40892 32548
rect 40948 32492 40960 32548
rect 40880 32480 40960 32492
rect 41040 32868 41120 32880
rect 41040 32812 41052 32868
rect 41108 32812 41120 32868
rect 41040 32548 41120 32812
rect 41040 32492 41052 32548
rect 41108 32492 41120 32548
rect 41040 32480 41120 32492
rect 41200 32868 41280 32880
rect 41200 32812 41212 32868
rect 41268 32812 41280 32868
rect 41200 32548 41280 32812
rect 41200 32492 41212 32548
rect 41268 32492 41280 32548
rect 41200 32480 41280 32492
rect 41360 32868 41440 32880
rect 41360 32812 41372 32868
rect 41428 32812 41440 32868
rect 41360 32548 41440 32812
rect 41360 32492 41372 32548
rect 41428 32492 41440 32548
rect 41360 32480 41440 32492
rect 41520 32868 41600 32880
rect 41520 32812 41532 32868
rect 41588 32812 41600 32868
rect 41520 32548 41600 32812
rect 41520 32492 41532 32548
rect 41588 32492 41600 32548
rect 41520 32480 41600 32492
rect 41680 32868 41760 32880
rect 41680 32812 41692 32868
rect 41748 32812 41760 32868
rect 41680 32548 41760 32812
rect 41680 32492 41692 32548
rect 41748 32492 41760 32548
rect 41680 32480 41760 32492
rect 41840 32868 41920 32880
rect 41840 32812 41852 32868
rect 41908 32812 41920 32868
rect 41840 32548 41920 32812
rect 41840 32492 41852 32548
rect 41908 32492 41920 32548
rect 41840 32480 41920 32492
rect 33520 32388 33600 32400
rect 33520 32332 33532 32388
rect 33588 32332 33600 32388
rect 33520 32068 33600 32332
rect 33520 32012 33532 32068
rect 33588 32012 33600 32068
rect 33520 31748 33600 32012
rect 33520 31692 33532 31748
rect 33588 31692 33600 31748
rect 33520 31428 33600 31692
rect 33520 31372 33532 31428
rect 33588 31372 33600 31428
rect 33520 31108 33600 31372
rect 33520 31052 33532 31108
rect 33588 31052 33600 31108
rect 33520 30788 33600 31052
rect 33520 30732 33532 30788
rect 33588 30732 33600 30788
rect 33520 30468 33600 30732
rect 33520 30412 33532 30468
rect 33588 30412 33600 30468
rect 33520 30400 33600 30412
rect 33680 32388 33760 32400
rect 33680 32332 33692 32388
rect 33748 32332 33760 32388
rect 33680 32068 33760 32332
rect 33680 32012 33692 32068
rect 33748 32012 33760 32068
rect 33680 31748 33760 32012
rect 33680 31692 33692 31748
rect 33748 31692 33760 31748
rect 33680 31428 33760 31692
rect 33680 31372 33692 31428
rect 33748 31372 33760 31428
rect 33680 31108 33760 31372
rect 33680 31052 33692 31108
rect 33748 31052 33760 31108
rect 33680 30788 33760 31052
rect 33680 30732 33692 30788
rect 33748 30732 33760 30788
rect 33680 30468 33760 30732
rect 33680 30412 33692 30468
rect 33748 30412 33760 30468
rect 33680 30400 33760 30412
rect 33840 32388 33920 32400
rect 33840 32332 33852 32388
rect 33908 32332 33920 32388
rect 33840 32068 33920 32332
rect 33840 32012 33852 32068
rect 33908 32012 33920 32068
rect 33840 31748 33920 32012
rect 33840 31692 33852 31748
rect 33908 31692 33920 31748
rect 33840 31428 33920 31692
rect 33840 31372 33852 31428
rect 33908 31372 33920 31428
rect 33840 31108 33920 31372
rect 33840 31052 33852 31108
rect 33908 31052 33920 31108
rect 33840 30788 33920 31052
rect 33840 30732 33852 30788
rect 33908 30732 33920 30788
rect 33840 30468 33920 30732
rect 33840 30412 33852 30468
rect 33908 30412 33920 30468
rect 33840 30400 33920 30412
rect 34000 32388 34080 32400
rect 34000 32332 34012 32388
rect 34068 32332 34080 32388
rect 34000 32068 34080 32332
rect 34000 32012 34012 32068
rect 34068 32012 34080 32068
rect 34000 31748 34080 32012
rect 34000 31692 34012 31748
rect 34068 31692 34080 31748
rect 34000 31428 34080 31692
rect 34000 31372 34012 31428
rect 34068 31372 34080 31428
rect 34000 31108 34080 31372
rect 34000 31052 34012 31108
rect 34068 31052 34080 31108
rect 34000 30788 34080 31052
rect 34000 30732 34012 30788
rect 34068 30732 34080 30788
rect 34000 30468 34080 30732
rect 34000 30412 34012 30468
rect 34068 30412 34080 30468
rect 34000 30400 34080 30412
rect 34160 32388 34240 32400
rect 34160 32332 34172 32388
rect 34228 32332 34240 32388
rect 34160 32068 34240 32332
rect 34160 32012 34172 32068
rect 34228 32012 34240 32068
rect 34160 31748 34240 32012
rect 34160 31692 34172 31748
rect 34228 31692 34240 31748
rect 34160 31428 34240 31692
rect 34160 31372 34172 31428
rect 34228 31372 34240 31428
rect 34160 31108 34240 31372
rect 34160 31052 34172 31108
rect 34228 31052 34240 31108
rect 34160 30788 34240 31052
rect 34160 30732 34172 30788
rect 34228 30732 34240 30788
rect 34160 30468 34240 30732
rect 34160 30412 34172 30468
rect 34228 30412 34240 30468
rect 34160 30400 34240 30412
rect 34320 32388 34400 32400
rect 34320 32332 34332 32388
rect 34388 32332 34400 32388
rect 34320 32068 34400 32332
rect 34320 32012 34332 32068
rect 34388 32012 34400 32068
rect 34320 31748 34400 32012
rect 34320 31692 34332 31748
rect 34388 31692 34400 31748
rect 34320 31428 34400 31692
rect 34320 31372 34332 31428
rect 34388 31372 34400 31428
rect 34320 31108 34400 31372
rect 34320 31052 34332 31108
rect 34388 31052 34400 31108
rect 34320 30788 34400 31052
rect 34320 30732 34332 30788
rect 34388 30732 34400 30788
rect 34320 30468 34400 30732
rect 34320 30412 34332 30468
rect 34388 30412 34400 30468
rect 34320 30400 34400 30412
rect 34480 32388 34560 32400
rect 34480 32332 34492 32388
rect 34548 32332 34560 32388
rect 34480 32068 34560 32332
rect 34480 32012 34492 32068
rect 34548 32012 34560 32068
rect 34480 31748 34560 32012
rect 34480 31692 34492 31748
rect 34548 31692 34560 31748
rect 34480 31428 34560 31692
rect 34480 31372 34492 31428
rect 34548 31372 34560 31428
rect 34480 31108 34560 31372
rect 34480 31052 34492 31108
rect 34548 31052 34560 31108
rect 34480 30788 34560 31052
rect 34480 30732 34492 30788
rect 34548 30732 34560 30788
rect 34480 30468 34560 30732
rect 34480 30412 34492 30468
rect 34548 30412 34560 30468
rect 34480 30400 34560 30412
rect 34640 32388 34720 32400
rect 34640 32332 34652 32388
rect 34708 32332 34720 32388
rect 34640 32068 34720 32332
rect 34640 32012 34652 32068
rect 34708 32012 34720 32068
rect 34640 31748 34720 32012
rect 34640 31692 34652 31748
rect 34708 31692 34720 31748
rect 34640 31428 34720 31692
rect 34640 31372 34652 31428
rect 34708 31372 34720 31428
rect 34640 31108 34720 31372
rect 34640 31052 34652 31108
rect 34708 31052 34720 31108
rect 34640 30788 34720 31052
rect 34640 30732 34652 30788
rect 34708 30732 34720 30788
rect 34640 30468 34720 30732
rect 34640 30412 34652 30468
rect 34708 30412 34720 30468
rect 34640 30400 34720 30412
rect 34800 32388 34880 32400
rect 34800 32332 34812 32388
rect 34868 32332 34880 32388
rect 34800 32068 34880 32332
rect 34800 32012 34812 32068
rect 34868 32012 34880 32068
rect 34800 31748 34880 32012
rect 34800 31692 34812 31748
rect 34868 31692 34880 31748
rect 34800 31428 34880 31692
rect 34800 31372 34812 31428
rect 34868 31372 34880 31428
rect 34800 31108 34880 31372
rect 34800 31052 34812 31108
rect 34868 31052 34880 31108
rect 34800 30788 34880 31052
rect 34800 30732 34812 30788
rect 34868 30732 34880 30788
rect 34800 30468 34880 30732
rect 34800 30412 34812 30468
rect 34868 30412 34880 30468
rect 34800 30400 34880 30412
rect 34960 32388 35040 32400
rect 34960 32332 34972 32388
rect 35028 32332 35040 32388
rect 34960 32068 35040 32332
rect 34960 32012 34972 32068
rect 35028 32012 35040 32068
rect 34960 31748 35040 32012
rect 34960 31692 34972 31748
rect 35028 31692 35040 31748
rect 34960 31428 35040 31692
rect 34960 31372 34972 31428
rect 35028 31372 35040 31428
rect 34960 31108 35040 31372
rect 34960 31052 34972 31108
rect 35028 31052 35040 31108
rect 34960 30788 35040 31052
rect 34960 30732 34972 30788
rect 35028 30732 35040 30788
rect 34960 30468 35040 30732
rect 34960 30412 34972 30468
rect 35028 30412 35040 30468
rect 34960 30400 35040 30412
rect 35120 32388 35200 32400
rect 35120 32332 35132 32388
rect 35188 32332 35200 32388
rect 35120 32068 35200 32332
rect 35120 32012 35132 32068
rect 35188 32012 35200 32068
rect 35120 31748 35200 32012
rect 35120 31692 35132 31748
rect 35188 31692 35200 31748
rect 35120 31428 35200 31692
rect 35120 31372 35132 31428
rect 35188 31372 35200 31428
rect 35120 31108 35200 31372
rect 35120 31052 35132 31108
rect 35188 31052 35200 31108
rect 35120 30788 35200 31052
rect 35120 30732 35132 30788
rect 35188 30732 35200 30788
rect 35120 30468 35200 30732
rect 35120 30412 35132 30468
rect 35188 30412 35200 30468
rect 35120 30400 35200 30412
rect 35280 32388 35360 32400
rect 35280 32332 35292 32388
rect 35348 32332 35360 32388
rect 35280 32068 35360 32332
rect 35280 32012 35292 32068
rect 35348 32012 35360 32068
rect 35280 31748 35360 32012
rect 35280 31692 35292 31748
rect 35348 31692 35360 31748
rect 35280 31428 35360 31692
rect 35280 31372 35292 31428
rect 35348 31372 35360 31428
rect 35280 31108 35360 31372
rect 35280 31052 35292 31108
rect 35348 31052 35360 31108
rect 35280 30788 35360 31052
rect 35280 30732 35292 30788
rect 35348 30732 35360 30788
rect 35280 30468 35360 30732
rect 35280 30412 35292 30468
rect 35348 30412 35360 30468
rect 35280 30400 35360 30412
rect 35440 32388 35520 32400
rect 35440 32332 35452 32388
rect 35508 32332 35520 32388
rect 35440 32068 35520 32332
rect 35440 32012 35452 32068
rect 35508 32012 35520 32068
rect 35440 31748 35520 32012
rect 35440 31692 35452 31748
rect 35508 31692 35520 31748
rect 35440 31428 35520 31692
rect 35440 31372 35452 31428
rect 35508 31372 35520 31428
rect 35440 31108 35520 31372
rect 35440 31052 35452 31108
rect 35508 31052 35520 31108
rect 35440 30788 35520 31052
rect 35440 30732 35452 30788
rect 35508 30732 35520 30788
rect 35440 30468 35520 30732
rect 35440 30412 35452 30468
rect 35508 30412 35520 30468
rect 35440 30400 35520 30412
rect 35600 32388 35680 32400
rect 35600 32332 35612 32388
rect 35668 32332 35680 32388
rect 35600 32068 35680 32332
rect 35600 32012 35612 32068
rect 35668 32012 35680 32068
rect 35600 31748 35680 32012
rect 35600 31692 35612 31748
rect 35668 31692 35680 31748
rect 35600 31428 35680 31692
rect 35600 31372 35612 31428
rect 35668 31372 35680 31428
rect 35600 31108 35680 31372
rect 35600 31052 35612 31108
rect 35668 31052 35680 31108
rect 35600 30788 35680 31052
rect 35600 30732 35612 30788
rect 35668 30732 35680 30788
rect 35600 30468 35680 30732
rect 35600 30412 35612 30468
rect 35668 30412 35680 30468
rect 35600 30400 35680 30412
rect 35760 32388 35840 32400
rect 35760 32332 35772 32388
rect 35828 32332 35840 32388
rect 35760 32068 35840 32332
rect 35760 32012 35772 32068
rect 35828 32012 35840 32068
rect 35760 31748 35840 32012
rect 35760 31692 35772 31748
rect 35828 31692 35840 31748
rect 35760 31428 35840 31692
rect 35760 31372 35772 31428
rect 35828 31372 35840 31428
rect 35760 31108 35840 31372
rect 35760 31052 35772 31108
rect 35828 31052 35840 31108
rect 35760 30788 35840 31052
rect 35760 30732 35772 30788
rect 35828 30732 35840 30788
rect 35760 30468 35840 30732
rect 35760 30412 35772 30468
rect 35828 30412 35840 30468
rect 35760 30400 35840 30412
rect 35920 32388 36000 32400
rect 35920 32332 35932 32388
rect 35988 32332 36000 32388
rect 35920 32068 36000 32332
rect 35920 32012 35932 32068
rect 35988 32012 36000 32068
rect 35920 31748 36000 32012
rect 35920 31692 35932 31748
rect 35988 31692 36000 31748
rect 35920 31428 36000 31692
rect 35920 31372 35932 31428
rect 35988 31372 36000 31428
rect 35920 31108 36000 31372
rect 35920 31052 35932 31108
rect 35988 31052 36000 31108
rect 35920 30788 36000 31052
rect 35920 30732 35932 30788
rect 35988 30732 36000 30788
rect 35920 30468 36000 30732
rect 35920 30412 35932 30468
rect 35988 30412 36000 30468
rect 35920 30400 36000 30412
rect 36080 32388 36160 32400
rect 36080 32332 36092 32388
rect 36148 32332 36160 32388
rect 36080 32068 36160 32332
rect 36080 32012 36092 32068
rect 36148 32012 36160 32068
rect 36080 31748 36160 32012
rect 36080 31692 36092 31748
rect 36148 31692 36160 31748
rect 36080 31428 36160 31692
rect 36080 31372 36092 31428
rect 36148 31372 36160 31428
rect 36080 31108 36160 31372
rect 36080 31052 36092 31108
rect 36148 31052 36160 31108
rect 36080 30788 36160 31052
rect 36080 30732 36092 30788
rect 36148 30732 36160 30788
rect 36080 30468 36160 30732
rect 36080 30412 36092 30468
rect 36148 30412 36160 30468
rect 36080 30400 36160 30412
rect 36240 32388 36320 32400
rect 36240 32332 36252 32388
rect 36308 32332 36320 32388
rect 36240 32068 36320 32332
rect 36240 32012 36252 32068
rect 36308 32012 36320 32068
rect 36240 31748 36320 32012
rect 36240 31692 36252 31748
rect 36308 31692 36320 31748
rect 36240 31428 36320 31692
rect 36240 31372 36252 31428
rect 36308 31372 36320 31428
rect 36240 31108 36320 31372
rect 36240 31052 36252 31108
rect 36308 31052 36320 31108
rect 36240 30788 36320 31052
rect 36240 30732 36252 30788
rect 36308 30732 36320 30788
rect 36240 30468 36320 30732
rect 36240 30412 36252 30468
rect 36308 30412 36320 30468
rect 36240 30400 36320 30412
rect 36400 32388 36480 32400
rect 36400 32332 36412 32388
rect 36468 32332 36480 32388
rect 36400 32068 36480 32332
rect 36400 32012 36412 32068
rect 36468 32012 36480 32068
rect 36400 31748 36480 32012
rect 36400 31692 36412 31748
rect 36468 31692 36480 31748
rect 36400 31428 36480 31692
rect 36400 31372 36412 31428
rect 36468 31372 36480 31428
rect 36400 31108 36480 31372
rect 36400 31052 36412 31108
rect 36468 31052 36480 31108
rect 36400 30788 36480 31052
rect 36400 30732 36412 30788
rect 36468 30732 36480 30788
rect 36400 30468 36480 30732
rect 36400 30412 36412 30468
rect 36468 30412 36480 30468
rect 36400 30400 36480 30412
rect 36560 32388 36640 32400
rect 36560 32332 36572 32388
rect 36628 32332 36640 32388
rect 36560 32068 36640 32332
rect 36560 32012 36572 32068
rect 36628 32012 36640 32068
rect 36560 31748 36640 32012
rect 36560 31692 36572 31748
rect 36628 31692 36640 31748
rect 36560 31428 36640 31692
rect 36560 31372 36572 31428
rect 36628 31372 36640 31428
rect 36560 31108 36640 31372
rect 36560 31052 36572 31108
rect 36628 31052 36640 31108
rect 36560 30788 36640 31052
rect 36560 30732 36572 30788
rect 36628 30732 36640 30788
rect 36560 30468 36640 30732
rect 36560 30412 36572 30468
rect 36628 30412 36640 30468
rect 36560 30400 36640 30412
rect 36720 32388 36800 32400
rect 36720 32332 36732 32388
rect 36788 32332 36800 32388
rect 36720 32068 36800 32332
rect 36720 32012 36732 32068
rect 36788 32012 36800 32068
rect 36720 31748 36800 32012
rect 36720 31692 36732 31748
rect 36788 31692 36800 31748
rect 36720 31428 36800 31692
rect 36720 31372 36732 31428
rect 36788 31372 36800 31428
rect 36720 31108 36800 31372
rect 36720 31052 36732 31108
rect 36788 31052 36800 31108
rect 36720 30788 36800 31052
rect 36720 30732 36732 30788
rect 36788 30732 36800 30788
rect 36720 30468 36800 30732
rect 36720 30412 36732 30468
rect 36788 30412 36800 30468
rect 36720 30400 36800 30412
rect 36880 32388 36960 32400
rect 36880 32332 36892 32388
rect 36948 32332 36960 32388
rect 36880 32068 36960 32332
rect 36880 32012 36892 32068
rect 36948 32012 36960 32068
rect 36880 31748 36960 32012
rect 36880 31692 36892 31748
rect 36948 31692 36960 31748
rect 36880 31428 36960 31692
rect 36880 31372 36892 31428
rect 36948 31372 36960 31428
rect 36880 31108 36960 31372
rect 36880 31052 36892 31108
rect 36948 31052 36960 31108
rect 36880 30788 36960 31052
rect 36880 30732 36892 30788
rect 36948 30732 36960 30788
rect 36880 30468 36960 30732
rect 36880 30412 36892 30468
rect 36948 30412 36960 30468
rect 36880 30400 36960 30412
rect 37040 32388 37120 32400
rect 37040 32332 37052 32388
rect 37108 32332 37120 32388
rect 37040 32068 37120 32332
rect 37040 32012 37052 32068
rect 37108 32012 37120 32068
rect 37040 31748 37120 32012
rect 37040 31692 37052 31748
rect 37108 31692 37120 31748
rect 37040 31428 37120 31692
rect 37040 31372 37052 31428
rect 37108 31372 37120 31428
rect 37040 31108 37120 31372
rect 37040 31052 37052 31108
rect 37108 31052 37120 31108
rect 37040 30788 37120 31052
rect 37040 30732 37052 30788
rect 37108 30732 37120 30788
rect 37040 30468 37120 30732
rect 37040 30412 37052 30468
rect 37108 30412 37120 30468
rect 37040 30400 37120 30412
rect 37200 32388 37280 32400
rect 37200 32332 37212 32388
rect 37268 32332 37280 32388
rect 37200 32068 37280 32332
rect 37200 32012 37212 32068
rect 37268 32012 37280 32068
rect 37200 31748 37280 32012
rect 37200 31692 37212 31748
rect 37268 31692 37280 31748
rect 37200 31428 37280 31692
rect 37200 31372 37212 31428
rect 37268 31372 37280 31428
rect 37200 31108 37280 31372
rect 37200 31052 37212 31108
rect 37268 31052 37280 31108
rect 37200 30788 37280 31052
rect 37200 30732 37212 30788
rect 37268 30732 37280 30788
rect 37200 30468 37280 30732
rect 37200 30412 37212 30468
rect 37268 30412 37280 30468
rect 37200 30400 37280 30412
rect 37360 32388 37440 32400
rect 37360 32332 37372 32388
rect 37428 32332 37440 32388
rect 37360 32068 37440 32332
rect 37360 32012 37372 32068
rect 37428 32012 37440 32068
rect 37360 31748 37440 32012
rect 37360 31692 37372 31748
rect 37428 31692 37440 31748
rect 37360 31428 37440 31692
rect 37360 31372 37372 31428
rect 37428 31372 37440 31428
rect 37360 31108 37440 31372
rect 37360 31052 37372 31108
rect 37428 31052 37440 31108
rect 37360 30788 37440 31052
rect 37360 30732 37372 30788
rect 37428 30732 37440 30788
rect 37360 30468 37440 30732
rect 37360 30412 37372 30468
rect 37428 30412 37440 30468
rect 37360 30400 37440 30412
rect 37520 32388 37600 32400
rect 37520 32332 37532 32388
rect 37588 32332 37600 32388
rect 37520 32068 37600 32332
rect 37520 32012 37532 32068
rect 37588 32012 37600 32068
rect 37520 31748 37600 32012
rect 37520 31692 37532 31748
rect 37588 31692 37600 31748
rect 37520 31428 37600 31692
rect 37520 31372 37532 31428
rect 37588 31372 37600 31428
rect 37520 31108 37600 31372
rect 37520 31052 37532 31108
rect 37588 31052 37600 31108
rect 37520 30788 37600 31052
rect 37520 30732 37532 30788
rect 37588 30732 37600 30788
rect 37520 30468 37600 30732
rect 37520 30412 37532 30468
rect 37588 30412 37600 30468
rect 37520 30400 37600 30412
rect 37680 32388 37760 32400
rect 37680 32332 37692 32388
rect 37748 32332 37760 32388
rect 37680 32068 37760 32332
rect 37680 32012 37692 32068
rect 37748 32012 37760 32068
rect 37680 31748 37760 32012
rect 37680 31692 37692 31748
rect 37748 31692 37760 31748
rect 37680 31428 37760 31692
rect 37680 31372 37692 31428
rect 37748 31372 37760 31428
rect 37680 31108 37760 31372
rect 37680 31052 37692 31108
rect 37748 31052 37760 31108
rect 37680 30788 37760 31052
rect 37680 30732 37692 30788
rect 37748 30732 37760 30788
rect 37680 30468 37760 30732
rect 37680 30412 37692 30468
rect 37748 30412 37760 30468
rect 37680 30400 37760 30412
rect 37840 32388 37920 32400
rect 37840 32332 37852 32388
rect 37908 32332 37920 32388
rect 37840 32068 37920 32332
rect 37840 32012 37852 32068
rect 37908 32012 37920 32068
rect 37840 31748 37920 32012
rect 37840 31692 37852 31748
rect 37908 31692 37920 31748
rect 37840 31428 37920 31692
rect 37840 31372 37852 31428
rect 37908 31372 37920 31428
rect 37840 31108 37920 31372
rect 37840 31052 37852 31108
rect 37908 31052 37920 31108
rect 37840 30788 37920 31052
rect 37840 30732 37852 30788
rect 37908 30732 37920 30788
rect 37840 30468 37920 30732
rect 37840 30412 37852 30468
rect 37908 30412 37920 30468
rect 37840 30400 37920 30412
rect 38000 32388 38080 32400
rect 38000 32332 38012 32388
rect 38068 32332 38080 32388
rect 38000 32068 38080 32332
rect 38000 32012 38012 32068
rect 38068 32012 38080 32068
rect 38000 31748 38080 32012
rect 38000 31692 38012 31748
rect 38068 31692 38080 31748
rect 38000 31428 38080 31692
rect 38000 31372 38012 31428
rect 38068 31372 38080 31428
rect 38000 31108 38080 31372
rect 38000 31052 38012 31108
rect 38068 31052 38080 31108
rect 38000 30788 38080 31052
rect 38000 30732 38012 30788
rect 38068 30732 38080 30788
rect 38000 30468 38080 30732
rect 38000 30412 38012 30468
rect 38068 30412 38080 30468
rect 38000 30400 38080 30412
rect 38160 32388 38240 32400
rect 38160 32332 38172 32388
rect 38228 32332 38240 32388
rect 38160 32068 38240 32332
rect 38160 32012 38172 32068
rect 38228 32012 38240 32068
rect 38160 31748 38240 32012
rect 38160 31692 38172 31748
rect 38228 31692 38240 31748
rect 38160 31428 38240 31692
rect 38160 31372 38172 31428
rect 38228 31372 38240 31428
rect 38160 31108 38240 31372
rect 38160 31052 38172 31108
rect 38228 31052 38240 31108
rect 38160 30788 38240 31052
rect 38160 30732 38172 30788
rect 38228 30732 38240 30788
rect 38160 30468 38240 30732
rect 38160 30412 38172 30468
rect 38228 30412 38240 30468
rect 38160 30400 38240 30412
rect 38320 32388 38400 32400
rect 38320 32332 38332 32388
rect 38388 32332 38400 32388
rect 38320 32068 38400 32332
rect 38320 32012 38332 32068
rect 38388 32012 38400 32068
rect 38320 31748 38400 32012
rect 38320 31692 38332 31748
rect 38388 31692 38400 31748
rect 38320 31428 38400 31692
rect 38320 31372 38332 31428
rect 38388 31372 38400 31428
rect 38320 31108 38400 31372
rect 38320 31052 38332 31108
rect 38388 31052 38400 31108
rect 38320 30788 38400 31052
rect 38320 30732 38332 30788
rect 38388 30732 38400 30788
rect 38320 30468 38400 30732
rect 38320 30412 38332 30468
rect 38388 30412 38400 30468
rect 38320 30400 38400 30412
rect 38480 32388 38560 32400
rect 38480 32332 38492 32388
rect 38548 32332 38560 32388
rect 38480 32068 38560 32332
rect 38480 32012 38492 32068
rect 38548 32012 38560 32068
rect 38480 31748 38560 32012
rect 38480 31692 38492 31748
rect 38548 31692 38560 31748
rect 38480 31428 38560 31692
rect 38480 31372 38492 31428
rect 38548 31372 38560 31428
rect 38480 31108 38560 31372
rect 38480 31052 38492 31108
rect 38548 31052 38560 31108
rect 38480 30788 38560 31052
rect 38480 30732 38492 30788
rect 38548 30732 38560 30788
rect 38480 30468 38560 30732
rect 38480 30412 38492 30468
rect 38548 30412 38560 30468
rect 38480 30400 38560 30412
rect 38640 32388 38720 32400
rect 38640 32332 38652 32388
rect 38708 32332 38720 32388
rect 38640 32068 38720 32332
rect 38640 32012 38652 32068
rect 38708 32012 38720 32068
rect 38640 31748 38720 32012
rect 38640 31692 38652 31748
rect 38708 31692 38720 31748
rect 38640 31428 38720 31692
rect 38640 31372 38652 31428
rect 38708 31372 38720 31428
rect 38640 31108 38720 31372
rect 38640 31052 38652 31108
rect 38708 31052 38720 31108
rect 38640 30788 38720 31052
rect 38640 30732 38652 30788
rect 38708 30732 38720 30788
rect 38640 30468 38720 30732
rect 38640 30412 38652 30468
rect 38708 30412 38720 30468
rect 38640 30400 38720 30412
rect 38800 32388 38880 32400
rect 38800 32332 38812 32388
rect 38868 32332 38880 32388
rect 38800 32068 38880 32332
rect 38800 32012 38812 32068
rect 38868 32012 38880 32068
rect 38800 31748 38880 32012
rect 38800 31692 38812 31748
rect 38868 31692 38880 31748
rect 38800 31428 38880 31692
rect 38800 31372 38812 31428
rect 38868 31372 38880 31428
rect 38800 31108 38880 31372
rect 38800 31052 38812 31108
rect 38868 31052 38880 31108
rect 38800 30788 38880 31052
rect 38800 30732 38812 30788
rect 38868 30732 38880 30788
rect 38800 30468 38880 30732
rect 38800 30412 38812 30468
rect 38868 30412 38880 30468
rect 38800 30400 38880 30412
rect 38960 32388 39040 32400
rect 38960 32332 38972 32388
rect 39028 32332 39040 32388
rect 38960 32068 39040 32332
rect 38960 32012 38972 32068
rect 39028 32012 39040 32068
rect 38960 31748 39040 32012
rect 38960 31692 38972 31748
rect 39028 31692 39040 31748
rect 38960 31428 39040 31692
rect 38960 31372 38972 31428
rect 39028 31372 39040 31428
rect 38960 31108 39040 31372
rect 38960 31052 38972 31108
rect 39028 31052 39040 31108
rect 38960 30788 39040 31052
rect 38960 30732 38972 30788
rect 39028 30732 39040 30788
rect 38960 30468 39040 30732
rect 38960 30412 38972 30468
rect 39028 30412 39040 30468
rect 38960 30400 39040 30412
rect 39120 32388 39200 32400
rect 39120 32332 39132 32388
rect 39188 32332 39200 32388
rect 39120 32068 39200 32332
rect 39120 32012 39132 32068
rect 39188 32012 39200 32068
rect 39120 31748 39200 32012
rect 39120 31692 39132 31748
rect 39188 31692 39200 31748
rect 39120 31428 39200 31692
rect 39120 31372 39132 31428
rect 39188 31372 39200 31428
rect 39120 31108 39200 31372
rect 39120 31052 39132 31108
rect 39188 31052 39200 31108
rect 39120 30788 39200 31052
rect 39120 30732 39132 30788
rect 39188 30732 39200 30788
rect 39120 30468 39200 30732
rect 39120 30412 39132 30468
rect 39188 30412 39200 30468
rect 39120 30400 39200 30412
rect 39280 32388 39360 32400
rect 39280 32332 39292 32388
rect 39348 32332 39360 32388
rect 39280 32068 39360 32332
rect 39280 32012 39292 32068
rect 39348 32012 39360 32068
rect 39280 31748 39360 32012
rect 39280 31692 39292 31748
rect 39348 31692 39360 31748
rect 39280 31428 39360 31692
rect 39280 31372 39292 31428
rect 39348 31372 39360 31428
rect 39280 31108 39360 31372
rect 39280 31052 39292 31108
rect 39348 31052 39360 31108
rect 39280 30788 39360 31052
rect 39280 30732 39292 30788
rect 39348 30732 39360 30788
rect 39280 30468 39360 30732
rect 39280 30412 39292 30468
rect 39348 30412 39360 30468
rect 39280 30400 39360 30412
rect 39440 32388 39520 32400
rect 39440 32332 39452 32388
rect 39508 32332 39520 32388
rect 39440 32068 39520 32332
rect 39440 32012 39452 32068
rect 39508 32012 39520 32068
rect 39440 31748 39520 32012
rect 39440 31692 39452 31748
rect 39508 31692 39520 31748
rect 39440 31428 39520 31692
rect 39440 31372 39452 31428
rect 39508 31372 39520 31428
rect 39440 31108 39520 31372
rect 39440 31052 39452 31108
rect 39508 31052 39520 31108
rect 39440 30788 39520 31052
rect 39440 30732 39452 30788
rect 39508 30732 39520 30788
rect 39440 30468 39520 30732
rect 39440 30412 39452 30468
rect 39508 30412 39520 30468
rect 39440 30400 39520 30412
rect 39600 32388 39680 32400
rect 39600 32332 39612 32388
rect 39668 32332 39680 32388
rect 39600 32068 39680 32332
rect 39600 32012 39612 32068
rect 39668 32012 39680 32068
rect 39600 31748 39680 32012
rect 39600 31692 39612 31748
rect 39668 31692 39680 31748
rect 39600 31428 39680 31692
rect 39600 31372 39612 31428
rect 39668 31372 39680 31428
rect 39600 31108 39680 31372
rect 39600 31052 39612 31108
rect 39668 31052 39680 31108
rect 39600 30788 39680 31052
rect 39600 30732 39612 30788
rect 39668 30732 39680 30788
rect 39600 30468 39680 30732
rect 39600 30412 39612 30468
rect 39668 30412 39680 30468
rect 39600 30400 39680 30412
rect 39760 32388 39840 32400
rect 39760 32332 39772 32388
rect 39828 32332 39840 32388
rect 39760 32068 39840 32332
rect 39760 32012 39772 32068
rect 39828 32012 39840 32068
rect 39760 31748 39840 32012
rect 39760 31692 39772 31748
rect 39828 31692 39840 31748
rect 39760 31428 39840 31692
rect 39760 31372 39772 31428
rect 39828 31372 39840 31428
rect 39760 31108 39840 31372
rect 39760 31052 39772 31108
rect 39828 31052 39840 31108
rect 39760 30788 39840 31052
rect 39760 30732 39772 30788
rect 39828 30732 39840 30788
rect 39760 30468 39840 30732
rect 39760 30412 39772 30468
rect 39828 30412 39840 30468
rect 39760 30400 39840 30412
rect 39920 32388 40000 32400
rect 39920 32332 39932 32388
rect 39988 32332 40000 32388
rect 39920 32068 40000 32332
rect 39920 32012 39932 32068
rect 39988 32012 40000 32068
rect 39920 31748 40000 32012
rect 39920 31692 39932 31748
rect 39988 31692 40000 31748
rect 39920 31428 40000 31692
rect 39920 31372 39932 31428
rect 39988 31372 40000 31428
rect 39920 31108 40000 31372
rect 39920 31052 39932 31108
rect 39988 31052 40000 31108
rect 39920 30788 40000 31052
rect 39920 30732 39932 30788
rect 39988 30732 40000 30788
rect 39920 30468 40000 30732
rect 39920 30412 39932 30468
rect 39988 30412 40000 30468
rect 39920 30400 40000 30412
rect 40080 32388 40160 32400
rect 40080 32332 40092 32388
rect 40148 32332 40160 32388
rect 40080 32068 40160 32332
rect 40080 32012 40092 32068
rect 40148 32012 40160 32068
rect 40080 31748 40160 32012
rect 40080 31692 40092 31748
rect 40148 31692 40160 31748
rect 40080 31428 40160 31692
rect 40080 31372 40092 31428
rect 40148 31372 40160 31428
rect 40080 31108 40160 31372
rect 40080 31052 40092 31108
rect 40148 31052 40160 31108
rect 40080 30788 40160 31052
rect 40080 30732 40092 30788
rect 40148 30732 40160 30788
rect 40080 30468 40160 30732
rect 40080 30412 40092 30468
rect 40148 30412 40160 30468
rect 40080 30400 40160 30412
rect 40240 32388 40320 32400
rect 40240 32332 40252 32388
rect 40308 32332 40320 32388
rect 40240 32068 40320 32332
rect 40240 32012 40252 32068
rect 40308 32012 40320 32068
rect 40240 31748 40320 32012
rect 40240 31692 40252 31748
rect 40308 31692 40320 31748
rect 40240 31428 40320 31692
rect 40240 31372 40252 31428
rect 40308 31372 40320 31428
rect 40240 31108 40320 31372
rect 40240 31052 40252 31108
rect 40308 31052 40320 31108
rect 40240 30788 40320 31052
rect 40240 30732 40252 30788
rect 40308 30732 40320 30788
rect 40240 30468 40320 30732
rect 40240 30412 40252 30468
rect 40308 30412 40320 30468
rect 40240 30400 40320 30412
rect 40400 32388 40480 32400
rect 40400 32332 40412 32388
rect 40468 32332 40480 32388
rect 40400 32068 40480 32332
rect 40400 32012 40412 32068
rect 40468 32012 40480 32068
rect 40400 31748 40480 32012
rect 40400 31692 40412 31748
rect 40468 31692 40480 31748
rect 40400 31428 40480 31692
rect 40400 31372 40412 31428
rect 40468 31372 40480 31428
rect 40400 31108 40480 31372
rect 40400 31052 40412 31108
rect 40468 31052 40480 31108
rect 40400 30788 40480 31052
rect 40400 30732 40412 30788
rect 40468 30732 40480 30788
rect 40400 30468 40480 30732
rect 40400 30412 40412 30468
rect 40468 30412 40480 30468
rect 40400 30400 40480 30412
rect 40560 32388 40640 32400
rect 40560 32332 40572 32388
rect 40628 32332 40640 32388
rect 40560 32068 40640 32332
rect 40560 32012 40572 32068
rect 40628 32012 40640 32068
rect 40560 31748 40640 32012
rect 40560 31692 40572 31748
rect 40628 31692 40640 31748
rect 40560 31428 40640 31692
rect 40560 31372 40572 31428
rect 40628 31372 40640 31428
rect 40560 31108 40640 31372
rect 40560 31052 40572 31108
rect 40628 31052 40640 31108
rect 40560 30788 40640 31052
rect 40560 30732 40572 30788
rect 40628 30732 40640 30788
rect 40560 30468 40640 30732
rect 40560 30412 40572 30468
rect 40628 30412 40640 30468
rect 40560 30400 40640 30412
rect 40720 32388 40800 32400
rect 40720 32332 40732 32388
rect 40788 32332 40800 32388
rect 40720 32068 40800 32332
rect 40720 32012 40732 32068
rect 40788 32012 40800 32068
rect 40720 31748 40800 32012
rect 40720 31692 40732 31748
rect 40788 31692 40800 31748
rect 40720 31428 40800 31692
rect 40720 31372 40732 31428
rect 40788 31372 40800 31428
rect 40720 31108 40800 31372
rect 40720 31052 40732 31108
rect 40788 31052 40800 31108
rect 40720 30788 40800 31052
rect 40720 30732 40732 30788
rect 40788 30732 40800 30788
rect 40720 30468 40800 30732
rect 40720 30412 40732 30468
rect 40788 30412 40800 30468
rect 40720 30400 40800 30412
rect 40880 32388 40960 32400
rect 40880 32332 40892 32388
rect 40948 32332 40960 32388
rect 40880 32068 40960 32332
rect 40880 32012 40892 32068
rect 40948 32012 40960 32068
rect 40880 31748 40960 32012
rect 40880 31692 40892 31748
rect 40948 31692 40960 31748
rect 40880 31428 40960 31692
rect 40880 31372 40892 31428
rect 40948 31372 40960 31428
rect 40880 31108 40960 31372
rect 40880 31052 40892 31108
rect 40948 31052 40960 31108
rect 40880 30788 40960 31052
rect 40880 30732 40892 30788
rect 40948 30732 40960 30788
rect 40880 30468 40960 30732
rect 40880 30412 40892 30468
rect 40948 30412 40960 30468
rect 40880 30400 40960 30412
rect 41040 32388 41120 32400
rect 41040 32332 41052 32388
rect 41108 32332 41120 32388
rect 41040 32068 41120 32332
rect 41040 32012 41052 32068
rect 41108 32012 41120 32068
rect 41040 31748 41120 32012
rect 41040 31692 41052 31748
rect 41108 31692 41120 31748
rect 41040 31428 41120 31692
rect 41040 31372 41052 31428
rect 41108 31372 41120 31428
rect 41040 31108 41120 31372
rect 41040 31052 41052 31108
rect 41108 31052 41120 31108
rect 41040 30788 41120 31052
rect 41040 30732 41052 30788
rect 41108 30732 41120 30788
rect 41040 30468 41120 30732
rect 41040 30412 41052 30468
rect 41108 30412 41120 30468
rect 41040 30400 41120 30412
rect 41200 32388 41280 32400
rect 41200 32332 41212 32388
rect 41268 32332 41280 32388
rect 41200 32068 41280 32332
rect 41200 32012 41212 32068
rect 41268 32012 41280 32068
rect 41200 31748 41280 32012
rect 41200 31692 41212 31748
rect 41268 31692 41280 31748
rect 41200 31428 41280 31692
rect 41200 31372 41212 31428
rect 41268 31372 41280 31428
rect 41200 31108 41280 31372
rect 41200 31052 41212 31108
rect 41268 31052 41280 31108
rect 41200 30788 41280 31052
rect 41200 30732 41212 30788
rect 41268 30732 41280 30788
rect 41200 30468 41280 30732
rect 41200 30412 41212 30468
rect 41268 30412 41280 30468
rect 41200 30400 41280 30412
rect 41360 32388 41440 32400
rect 41360 32332 41372 32388
rect 41428 32332 41440 32388
rect 41360 32068 41440 32332
rect 41360 32012 41372 32068
rect 41428 32012 41440 32068
rect 41360 31748 41440 32012
rect 41360 31692 41372 31748
rect 41428 31692 41440 31748
rect 41360 31428 41440 31692
rect 41360 31372 41372 31428
rect 41428 31372 41440 31428
rect 41360 31108 41440 31372
rect 41360 31052 41372 31108
rect 41428 31052 41440 31108
rect 41360 30788 41440 31052
rect 41360 30732 41372 30788
rect 41428 30732 41440 30788
rect 41360 30468 41440 30732
rect 41360 30412 41372 30468
rect 41428 30412 41440 30468
rect 41360 30400 41440 30412
rect 41520 32388 41600 32400
rect 41520 32332 41532 32388
rect 41588 32332 41600 32388
rect 41520 32068 41600 32332
rect 41520 32012 41532 32068
rect 41588 32012 41600 32068
rect 41520 31748 41600 32012
rect 41520 31692 41532 31748
rect 41588 31692 41600 31748
rect 41520 31428 41600 31692
rect 41520 31372 41532 31428
rect 41588 31372 41600 31428
rect 41520 31108 41600 31372
rect 41520 31052 41532 31108
rect 41588 31052 41600 31108
rect 41520 30788 41600 31052
rect 41520 30732 41532 30788
rect 41588 30732 41600 30788
rect 41520 30468 41600 30732
rect 41520 30412 41532 30468
rect 41588 30412 41600 30468
rect 41520 30400 41600 30412
rect 41680 32388 41760 32400
rect 41680 32332 41692 32388
rect 41748 32332 41760 32388
rect 41680 32068 41760 32332
rect 41680 32012 41692 32068
rect 41748 32012 41760 32068
rect 41680 31748 41760 32012
rect 41680 31692 41692 31748
rect 41748 31692 41760 31748
rect 41680 31428 41760 31692
rect 41680 31372 41692 31428
rect 41748 31372 41760 31428
rect 41680 31108 41760 31372
rect 41680 31052 41692 31108
rect 41748 31052 41760 31108
rect 41680 30788 41760 31052
rect 41680 30732 41692 30788
rect 41748 30732 41760 30788
rect 41680 30468 41760 30732
rect 41680 30412 41692 30468
rect 41748 30412 41760 30468
rect 41680 30400 41760 30412
rect 41840 32388 41920 32400
rect 41840 32332 41852 32388
rect 41908 32332 41920 32388
rect 41840 32068 41920 32332
rect 41840 32012 41852 32068
rect 41908 32012 41920 32068
rect 41840 31748 41920 32012
rect 41840 31692 41852 31748
rect 41908 31692 41920 31748
rect 41840 31428 41920 31692
rect 41840 31372 41852 31428
rect 41908 31372 41920 31428
rect 41840 31108 41920 31372
rect 41840 31052 41852 31108
rect 41908 31052 41920 31108
rect 41840 30788 41920 31052
rect 41840 30732 41852 30788
rect 41908 30732 41920 30788
rect 41840 30468 41920 30732
rect 41840 30412 41852 30468
rect 41908 30412 41920 30468
rect 41840 30400 41920 30412
rect 33520 30308 33600 30320
rect 33520 30252 33532 30308
rect 33588 30252 33600 30308
rect 33520 29988 33600 30252
rect 33520 29932 33532 29988
rect 33588 29932 33600 29988
rect 33520 29920 33600 29932
rect 33680 30308 33760 30320
rect 33680 30252 33692 30308
rect 33748 30252 33760 30308
rect 33680 29988 33760 30252
rect 33680 29932 33692 29988
rect 33748 29932 33760 29988
rect 33680 29920 33760 29932
rect 33840 30308 33920 30320
rect 33840 30252 33852 30308
rect 33908 30252 33920 30308
rect 33840 29988 33920 30252
rect 33840 29932 33852 29988
rect 33908 29932 33920 29988
rect 33840 29920 33920 29932
rect 34000 30308 34080 30320
rect 34000 30252 34012 30308
rect 34068 30252 34080 30308
rect 34000 29988 34080 30252
rect 34000 29932 34012 29988
rect 34068 29932 34080 29988
rect 34000 29920 34080 29932
rect 34160 30308 34240 30320
rect 34160 30252 34172 30308
rect 34228 30252 34240 30308
rect 34160 29988 34240 30252
rect 34160 29932 34172 29988
rect 34228 29932 34240 29988
rect 34160 29920 34240 29932
rect 34320 30308 34400 30320
rect 34320 30252 34332 30308
rect 34388 30252 34400 30308
rect 34320 29988 34400 30252
rect 34320 29932 34332 29988
rect 34388 29932 34400 29988
rect 34320 29920 34400 29932
rect 34480 30308 34560 30320
rect 34480 30252 34492 30308
rect 34548 30252 34560 30308
rect 34480 29988 34560 30252
rect 34480 29932 34492 29988
rect 34548 29932 34560 29988
rect 34480 29920 34560 29932
rect 34640 30308 34720 30320
rect 34640 30252 34652 30308
rect 34708 30252 34720 30308
rect 34640 29988 34720 30252
rect 34640 29932 34652 29988
rect 34708 29932 34720 29988
rect 34640 29920 34720 29932
rect 34800 30308 34880 30320
rect 34800 30252 34812 30308
rect 34868 30252 34880 30308
rect 34800 29988 34880 30252
rect 34800 29932 34812 29988
rect 34868 29932 34880 29988
rect 34800 29920 34880 29932
rect 34960 30308 35040 30320
rect 34960 30252 34972 30308
rect 35028 30252 35040 30308
rect 34960 29988 35040 30252
rect 34960 29932 34972 29988
rect 35028 29932 35040 29988
rect 34960 29920 35040 29932
rect 35120 30308 35200 30320
rect 35120 30252 35132 30308
rect 35188 30252 35200 30308
rect 35120 29988 35200 30252
rect 35120 29932 35132 29988
rect 35188 29932 35200 29988
rect 35120 29920 35200 29932
rect 35280 30308 35360 30320
rect 35280 30252 35292 30308
rect 35348 30252 35360 30308
rect 35280 29988 35360 30252
rect 35280 29932 35292 29988
rect 35348 29932 35360 29988
rect 35280 29920 35360 29932
rect 35440 30308 35520 30320
rect 35440 30252 35452 30308
rect 35508 30252 35520 30308
rect 35440 29988 35520 30252
rect 35440 29932 35452 29988
rect 35508 29932 35520 29988
rect 35440 29920 35520 29932
rect 35600 30308 35680 30320
rect 35600 30252 35612 30308
rect 35668 30252 35680 30308
rect 35600 29988 35680 30252
rect 35600 29932 35612 29988
rect 35668 29932 35680 29988
rect 35600 29920 35680 29932
rect 35760 30308 35840 30320
rect 35760 30252 35772 30308
rect 35828 30252 35840 30308
rect 35760 29988 35840 30252
rect 35760 29932 35772 29988
rect 35828 29932 35840 29988
rect 35760 29920 35840 29932
rect 35920 30308 36000 30320
rect 35920 30252 35932 30308
rect 35988 30252 36000 30308
rect 35920 29988 36000 30252
rect 35920 29932 35932 29988
rect 35988 29932 36000 29988
rect 35920 29920 36000 29932
rect 36080 30308 36160 30320
rect 36080 30252 36092 30308
rect 36148 30252 36160 30308
rect 36080 29988 36160 30252
rect 36080 29932 36092 29988
rect 36148 29932 36160 29988
rect 36080 29920 36160 29932
rect 36240 30308 36320 30320
rect 36240 30252 36252 30308
rect 36308 30252 36320 30308
rect 36240 29988 36320 30252
rect 36240 29932 36252 29988
rect 36308 29932 36320 29988
rect 36240 29920 36320 29932
rect 36400 30308 36480 30320
rect 36400 30252 36412 30308
rect 36468 30252 36480 30308
rect 36400 29988 36480 30252
rect 36400 29932 36412 29988
rect 36468 29932 36480 29988
rect 36400 29920 36480 29932
rect 36560 30308 36640 30320
rect 36560 30252 36572 30308
rect 36628 30252 36640 30308
rect 36560 29988 36640 30252
rect 36560 29932 36572 29988
rect 36628 29932 36640 29988
rect 36560 29920 36640 29932
rect 36720 30308 36800 30320
rect 36720 30252 36732 30308
rect 36788 30252 36800 30308
rect 36720 29988 36800 30252
rect 36720 29932 36732 29988
rect 36788 29932 36800 29988
rect 36720 29920 36800 29932
rect 36880 30308 36960 30320
rect 36880 30252 36892 30308
rect 36948 30252 36960 30308
rect 36880 29988 36960 30252
rect 36880 29932 36892 29988
rect 36948 29932 36960 29988
rect 36880 29920 36960 29932
rect 37040 30308 37120 30320
rect 37040 30252 37052 30308
rect 37108 30252 37120 30308
rect 37040 29988 37120 30252
rect 37040 29932 37052 29988
rect 37108 29932 37120 29988
rect 37040 29920 37120 29932
rect 37200 30308 37280 30320
rect 37200 30252 37212 30308
rect 37268 30252 37280 30308
rect 37200 29988 37280 30252
rect 37200 29932 37212 29988
rect 37268 29932 37280 29988
rect 37200 29920 37280 29932
rect 37360 30308 37440 30320
rect 37360 30252 37372 30308
rect 37428 30252 37440 30308
rect 37360 29988 37440 30252
rect 37360 29932 37372 29988
rect 37428 29932 37440 29988
rect 37360 29920 37440 29932
rect 37520 30308 37600 30320
rect 37520 30252 37532 30308
rect 37588 30252 37600 30308
rect 37520 29988 37600 30252
rect 37520 29932 37532 29988
rect 37588 29932 37600 29988
rect 37520 29920 37600 29932
rect 37680 30308 37760 30320
rect 37680 30252 37692 30308
rect 37748 30252 37760 30308
rect 37680 29988 37760 30252
rect 37680 29932 37692 29988
rect 37748 29932 37760 29988
rect 37680 29920 37760 29932
rect 37840 30308 37920 30320
rect 37840 30252 37852 30308
rect 37908 30252 37920 30308
rect 37840 29988 37920 30252
rect 37840 29932 37852 29988
rect 37908 29932 37920 29988
rect 37840 29920 37920 29932
rect 38000 30308 38080 30320
rect 38000 30252 38012 30308
rect 38068 30252 38080 30308
rect 38000 29988 38080 30252
rect 38000 29932 38012 29988
rect 38068 29932 38080 29988
rect 38000 29920 38080 29932
rect 38160 30308 38240 30320
rect 38160 30252 38172 30308
rect 38228 30252 38240 30308
rect 38160 29988 38240 30252
rect 38160 29932 38172 29988
rect 38228 29932 38240 29988
rect 38160 29920 38240 29932
rect 38320 30308 38400 30320
rect 38320 30252 38332 30308
rect 38388 30252 38400 30308
rect 38320 29988 38400 30252
rect 38320 29932 38332 29988
rect 38388 29932 38400 29988
rect 38320 29920 38400 29932
rect 38480 30308 38560 30320
rect 38480 30252 38492 30308
rect 38548 30252 38560 30308
rect 38480 29988 38560 30252
rect 38480 29932 38492 29988
rect 38548 29932 38560 29988
rect 38480 29920 38560 29932
rect 38640 30308 38720 30320
rect 38640 30252 38652 30308
rect 38708 30252 38720 30308
rect 38640 29988 38720 30252
rect 38640 29932 38652 29988
rect 38708 29932 38720 29988
rect 38640 29920 38720 29932
rect 38800 30308 38880 30320
rect 38800 30252 38812 30308
rect 38868 30252 38880 30308
rect 38800 29988 38880 30252
rect 38800 29932 38812 29988
rect 38868 29932 38880 29988
rect 38800 29920 38880 29932
rect 38960 30308 39040 30320
rect 38960 30252 38972 30308
rect 39028 30252 39040 30308
rect 38960 29988 39040 30252
rect 38960 29932 38972 29988
rect 39028 29932 39040 29988
rect 38960 29920 39040 29932
rect 39120 30308 39200 30320
rect 39120 30252 39132 30308
rect 39188 30252 39200 30308
rect 39120 29988 39200 30252
rect 39120 29932 39132 29988
rect 39188 29932 39200 29988
rect 39120 29920 39200 29932
rect 39280 30308 39360 30320
rect 39280 30252 39292 30308
rect 39348 30252 39360 30308
rect 39280 29988 39360 30252
rect 39280 29932 39292 29988
rect 39348 29932 39360 29988
rect 39280 29920 39360 29932
rect 39440 30308 39520 30320
rect 39440 30252 39452 30308
rect 39508 30252 39520 30308
rect 39440 29988 39520 30252
rect 39440 29932 39452 29988
rect 39508 29932 39520 29988
rect 39440 29920 39520 29932
rect 39600 30308 39680 30320
rect 39600 30252 39612 30308
rect 39668 30252 39680 30308
rect 39600 29988 39680 30252
rect 39600 29932 39612 29988
rect 39668 29932 39680 29988
rect 39600 29920 39680 29932
rect 39760 30308 39840 30320
rect 39760 30252 39772 30308
rect 39828 30252 39840 30308
rect 39760 29988 39840 30252
rect 39760 29932 39772 29988
rect 39828 29932 39840 29988
rect 39760 29920 39840 29932
rect 39920 30308 40000 30320
rect 39920 30252 39932 30308
rect 39988 30252 40000 30308
rect 39920 29988 40000 30252
rect 39920 29932 39932 29988
rect 39988 29932 40000 29988
rect 39920 29920 40000 29932
rect 40080 30308 40160 30320
rect 40080 30252 40092 30308
rect 40148 30252 40160 30308
rect 40080 29988 40160 30252
rect 40080 29932 40092 29988
rect 40148 29932 40160 29988
rect 40080 29920 40160 29932
rect 40240 30308 40320 30320
rect 40240 30252 40252 30308
rect 40308 30252 40320 30308
rect 40240 29988 40320 30252
rect 40240 29932 40252 29988
rect 40308 29932 40320 29988
rect 40240 29920 40320 29932
rect 40400 30308 40480 30320
rect 40400 30252 40412 30308
rect 40468 30252 40480 30308
rect 40400 29988 40480 30252
rect 40400 29932 40412 29988
rect 40468 29932 40480 29988
rect 40400 29920 40480 29932
rect 40560 30308 40640 30320
rect 40560 30252 40572 30308
rect 40628 30252 40640 30308
rect 40560 29988 40640 30252
rect 40560 29932 40572 29988
rect 40628 29932 40640 29988
rect 40560 29920 40640 29932
rect 40720 30308 40800 30320
rect 40720 30252 40732 30308
rect 40788 30252 40800 30308
rect 40720 29988 40800 30252
rect 40720 29932 40732 29988
rect 40788 29932 40800 29988
rect 40720 29920 40800 29932
rect 40880 30308 40960 30320
rect 40880 30252 40892 30308
rect 40948 30252 40960 30308
rect 40880 29988 40960 30252
rect 40880 29932 40892 29988
rect 40948 29932 40960 29988
rect 40880 29920 40960 29932
rect 41040 30308 41120 30320
rect 41040 30252 41052 30308
rect 41108 30252 41120 30308
rect 41040 29988 41120 30252
rect 41040 29932 41052 29988
rect 41108 29932 41120 29988
rect 41040 29920 41120 29932
rect 41200 30308 41280 30320
rect 41200 30252 41212 30308
rect 41268 30252 41280 30308
rect 41200 29988 41280 30252
rect 41200 29932 41212 29988
rect 41268 29932 41280 29988
rect 41200 29920 41280 29932
rect 41360 30308 41440 30320
rect 41360 30252 41372 30308
rect 41428 30252 41440 30308
rect 41360 29988 41440 30252
rect 41360 29932 41372 29988
rect 41428 29932 41440 29988
rect 41360 29920 41440 29932
rect 41520 30308 41600 30320
rect 41520 30252 41532 30308
rect 41588 30252 41600 30308
rect 41520 29988 41600 30252
rect 41520 29932 41532 29988
rect 41588 29932 41600 29988
rect 41520 29920 41600 29932
rect 41680 30308 41760 30320
rect 41680 30252 41692 30308
rect 41748 30252 41760 30308
rect 41680 29988 41760 30252
rect 41680 29932 41692 29988
rect 41748 29932 41760 29988
rect 41680 29920 41760 29932
rect 41840 30308 41920 30320
rect 41840 30252 41852 30308
rect 41908 30252 41920 30308
rect 41840 29988 41920 30252
rect 41840 29932 41852 29988
rect 41908 29932 41920 29988
rect 41840 29920 41920 29932
rect 33520 29828 33600 29840
rect 33520 29772 33532 29828
rect 33588 29772 33600 29828
rect 33520 29508 33600 29772
rect 33520 29452 33532 29508
rect 33588 29452 33600 29508
rect 33520 29440 33600 29452
rect 33680 29828 33760 29840
rect 33680 29772 33692 29828
rect 33748 29772 33760 29828
rect 33680 29508 33760 29772
rect 33680 29452 33692 29508
rect 33748 29452 33760 29508
rect 33680 29440 33760 29452
rect 33840 29828 33920 29840
rect 33840 29772 33852 29828
rect 33908 29772 33920 29828
rect 33840 29508 33920 29772
rect 33840 29452 33852 29508
rect 33908 29452 33920 29508
rect 33840 29440 33920 29452
rect 34000 29828 34080 29840
rect 34000 29772 34012 29828
rect 34068 29772 34080 29828
rect 34000 29508 34080 29772
rect 34000 29452 34012 29508
rect 34068 29452 34080 29508
rect 34000 29440 34080 29452
rect 34160 29828 34240 29840
rect 34160 29772 34172 29828
rect 34228 29772 34240 29828
rect 34160 29508 34240 29772
rect 34160 29452 34172 29508
rect 34228 29452 34240 29508
rect 34160 29440 34240 29452
rect 34320 29828 34400 29840
rect 34320 29772 34332 29828
rect 34388 29772 34400 29828
rect 34320 29508 34400 29772
rect 34320 29452 34332 29508
rect 34388 29452 34400 29508
rect 34320 29440 34400 29452
rect 34480 29828 34560 29840
rect 34480 29772 34492 29828
rect 34548 29772 34560 29828
rect 34480 29508 34560 29772
rect 34480 29452 34492 29508
rect 34548 29452 34560 29508
rect 34480 29440 34560 29452
rect 34640 29828 34720 29840
rect 34640 29772 34652 29828
rect 34708 29772 34720 29828
rect 34640 29508 34720 29772
rect 34640 29452 34652 29508
rect 34708 29452 34720 29508
rect 34640 29440 34720 29452
rect 34800 29828 34880 29840
rect 34800 29772 34812 29828
rect 34868 29772 34880 29828
rect 34800 29508 34880 29772
rect 34800 29452 34812 29508
rect 34868 29452 34880 29508
rect 34800 29440 34880 29452
rect 34960 29828 35040 29840
rect 34960 29772 34972 29828
rect 35028 29772 35040 29828
rect 34960 29508 35040 29772
rect 34960 29452 34972 29508
rect 35028 29452 35040 29508
rect 34960 29440 35040 29452
rect 35120 29828 35200 29840
rect 35120 29772 35132 29828
rect 35188 29772 35200 29828
rect 35120 29508 35200 29772
rect 35120 29452 35132 29508
rect 35188 29452 35200 29508
rect 35120 29440 35200 29452
rect 35280 29828 35360 29840
rect 35280 29772 35292 29828
rect 35348 29772 35360 29828
rect 35280 29508 35360 29772
rect 35280 29452 35292 29508
rect 35348 29452 35360 29508
rect 35280 29440 35360 29452
rect 35440 29828 35520 29840
rect 35440 29772 35452 29828
rect 35508 29772 35520 29828
rect 35440 29508 35520 29772
rect 35440 29452 35452 29508
rect 35508 29452 35520 29508
rect 35440 29440 35520 29452
rect 35600 29828 35680 29840
rect 35600 29772 35612 29828
rect 35668 29772 35680 29828
rect 35600 29508 35680 29772
rect 35600 29452 35612 29508
rect 35668 29452 35680 29508
rect 35600 29440 35680 29452
rect 35760 29828 35840 29840
rect 35760 29772 35772 29828
rect 35828 29772 35840 29828
rect 35760 29508 35840 29772
rect 35760 29452 35772 29508
rect 35828 29452 35840 29508
rect 35760 29440 35840 29452
rect 35920 29828 36000 29840
rect 35920 29772 35932 29828
rect 35988 29772 36000 29828
rect 35920 29508 36000 29772
rect 35920 29452 35932 29508
rect 35988 29452 36000 29508
rect 35920 29440 36000 29452
rect 36080 29828 36160 29840
rect 36080 29772 36092 29828
rect 36148 29772 36160 29828
rect 36080 29508 36160 29772
rect 36080 29452 36092 29508
rect 36148 29452 36160 29508
rect 36080 29440 36160 29452
rect 36240 29828 36320 29840
rect 36240 29772 36252 29828
rect 36308 29772 36320 29828
rect 36240 29508 36320 29772
rect 36240 29452 36252 29508
rect 36308 29452 36320 29508
rect 36240 29440 36320 29452
rect 36400 29828 36480 29840
rect 36400 29772 36412 29828
rect 36468 29772 36480 29828
rect 36400 29508 36480 29772
rect 36400 29452 36412 29508
rect 36468 29452 36480 29508
rect 36400 29440 36480 29452
rect 36560 29828 36640 29840
rect 36560 29772 36572 29828
rect 36628 29772 36640 29828
rect 36560 29508 36640 29772
rect 36560 29452 36572 29508
rect 36628 29452 36640 29508
rect 36560 29440 36640 29452
rect 36720 29828 36800 29840
rect 36720 29772 36732 29828
rect 36788 29772 36800 29828
rect 36720 29508 36800 29772
rect 36720 29452 36732 29508
rect 36788 29452 36800 29508
rect 36720 29440 36800 29452
rect 36880 29828 36960 29840
rect 36880 29772 36892 29828
rect 36948 29772 36960 29828
rect 36880 29508 36960 29772
rect 36880 29452 36892 29508
rect 36948 29452 36960 29508
rect 36880 29440 36960 29452
rect 37040 29828 37120 29840
rect 37040 29772 37052 29828
rect 37108 29772 37120 29828
rect 37040 29508 37120 29772
rect 37040 29452 37052 29508
rect 37108 29452 37120 29508
rect 37040 29440 37120 29452
rect 37200 29828 37280 29840
rect 37200 29772 37212 29828
rect 37268 29772 37280 29828
rect 37200 29508 37280 29772
rect 37200 29452 37212 29508
rect 37268 29452 37280 29508
rect 37200 29440 37280 29452
rect 37360 29828 37440 29840
rect 37360 29772 37372 29828
rect 37428 29772 37440 29828
rect 37360 29508 37440 29772
rect 37360 29452 37372 29508
rect 37428 29452 37440 29508
rect 37360 29440 37440 29452
rect 37520 29828 37600 29840
rect 37520 29772 37532 29828
rect 37588 29772 37600 29828
rect 37520 29508 37600 29772
rect 37520 29452 37532 29508
rect 37588 29452 37600 29508
rect 37520 29440 37600 29452
rect 37680 29828 37760 29840
rect 37680 29772 37692 29828
rect 37748 29772 37760 29828
rect 37680 29508 37760 29772
rect 37680 29452 37692 29508
rect 37748 29452 37760 29508
rect 37680 29440 37760 29452
rect 37840 29828 37920 29840
rect 37840 29772 37852 29828
rect 37908 29772 37920 29828
rect 37840 29508 37920 29772
rect 37840 29452 37852 29508
rect 37908 29452 37920 29508
rect 37840 29440 37920 29452
rect 38000 29828 38080 29840
rect 38000 29772 38012 29828
rect 38068 29772 38080 29828
rect 38000 29508 38080 29772
rect 38000 29452 38012 29508
rect 38068 29452 38080 29508
rect 38000 29440 38080 29452
rect 38160 29828 38240 29840
rect 38160 29772 38172 29828
rect 38228 29772 38240 29828
rect 38160 29508 38240 29772
rect 38160 29452 38172 29508
rect 38228 29452 38240 29508
rect 38160 29440 38240 29452
rect 38320 29828 38400 29840
rect 38320 29772 38332 29828
rect 38388 29772 38400 29828
rect 38320 29508 38400 29772
rect 38320 29452 38332 29508
rect 38388 29452 38400 29508
rect 38320 29440 38400 29452
rect 38480 29828 38560 29840
rect 38480 29772 38492 29828
rect 38548 29772 38560 29828
rect 38480 29508 38560 29772
rect 38480 29452 38492 29508
rect 38548 29452 38560 29508
rect 38480 29440 38560 29452
rect 38640 29828 38720 29840
rect 38640 29772 38652 29828
rect 38708 29772 38720 29828
rect 38640 29508 38720 29772
rect 38640 29452 38652 29508
rect 38708 29452 38720 29508
rect 38640 29440 38720 29452
rect 38800 29828 38880 29840
rect 38800 29772 38812 29828
rect 38868 29772 38880 29828
rect 38800 29508 38880 29772
rect 38800 29452 38812 29508
rect 38868 29452 38880 29508
rect 38800 29440 38880 29452
rect 38960 29828 39040 29840
rect 38960 29772 38972 29828
rect 39028 29772 39040 29828
rect 38960 29508 39040 29772
rect 38960 29452 38972 29508
rect 39028 29452 39040 29508
rect 38960 29440 39040 29452
rect 39120 29828 39200 29840
rect 39120 29772 39132 29828
rect 39188 29772 39200 29828
rect 39120 29508 39200 29772
rect 39120 29452 39132 29508
rect 39188 29452 39200 29508
rect 39120 29440 39200 29452
rect 39280 29828 39360 29840
rect 39280 29772 39292 29828
rect 39348 29772 39360 29828
rect 39280 29508 39360 29772
rect 39280 29452 39292 29508
rect 39348 29452 39360 29508
rect 39280 29440 39360 29452
rect 39440 29828 39520 29840
rect 39440 29772 39452 29828
rect 39508 29772 39520 29828
rect 39440 29508 39520 29772
rect 39440 29452 39452 29508
rect 39508 29452 39520 29508
rect 39440 29440 39520 29452
rect 39600 29828 39680 29840
rect 39600 29772 39612 29828
rect 39668 29772 39680 29828
rect 39600 29508 39680 29772
rect 39600 29452 39612 29508
rect 39668 29452 39680 29508
rect 39600 29440 39680 29452
rect 39760 29828 39840 29840
rect 39760 29772 39772 29828
rect 39828 29772 39840 29828
rect 39760 29508 39840 29772
rect 39760 29452 39772 29508
rect 39828 29452 39840 29508
rect 39760 29440 39840 29452
rect 39920 29828 40000 29840
rect 39920 29772 39932 29828
rect 39988 29772 40000 29828
rect 39920 29508 40000 29772
rect 39920 29452 39932 29508
rect 39988 29452 40000 29508
rect 39920 29440 40000 29452
rect 40080 29828 40160 29840
rect 40080 29772 40092 29828
rect 40148 29772 40160 29828
rect 40080 29508 40160 29772
rect 40080 29452 40092 29508
rect 40148 29452 40160 29508
rect 40080 29440 40160 29452
rect 40240 29828 40320 29840
rect 40240 29772 40252 29828
rect 40308 29772 40320 29828
rect 40240 29508 40320 29772
rect 40240 29452 40252 29508
rect 40308 29452 40320 29508
rect 40240 29440 40320 29452
rect 40400 29828 40480 29840
rect 40400 29772 40412 29828
rect 40468 29772 40480 29828
rect 40400 29508 40480 29772
rect 40400 29452 40412 29508
rect 40468 29452 40480 29508
rect 40400 29440 40480 29452
rect 40560 29828 40640 29840
rect 40560 29772 40572 29828
rect 40628 29772 40640 29828
rect 40560 29508 40640 29772
rect 40560 29452 40572 29508
rect 40628 29452 40640 29508
rect 40560 29440 40640 29452
rect 40720 29828 40800 29840
rect 40720 29772 40732 29828
rect 40788 29772 40800 29828
rect 40720 29508 40800 29772
rect 40720 29452 40732 29508
rect 40788 29452 40800 29508
rect 40720 29440 40800 29452
rect 40880 29828 40960 29840
rect 40880 29772 40892 29828
rect 40948 29772 40960 29828
rect 40880 29508 40960 29772
rect 40880 29452 40892 29508
rect 40948 29452 40960 29508
rect 40880 29440 40960 29452
rect 41040 29828 41120 29840
rect 41040 29772 41052 29828
rect 41108 29772 41120 29828
rect 41040 29508 41120 29772
rect 41040 29452 41052 29508
rect 41108 29452 41120 29508
rect 41040 29440 41120 29452
rect 41200 29828 41280 29840
rect 41200 29772 41212 29828
rect 41268 29772 41280 29828
rect 41200 29508 41280 29772
rect 41200 29452 41212 29508
rect 41268 29452 41280 29508
rect 41200 29440 41280 29452
rect 41360 29828 41440 29840
rect 41360 29772 41372 29828
rect 41428 29772 41440 29828
rect 41360 29508 41440 29772
rect 41360 29452 41372 29508
rect 41428 29452 41440 29508
rect 41360 29440 41440 29452
rect 41520 29828 41600 29840
rect 41520 29772 41532 29828
rect 41588 29772 41600 29828
rect 41520 29508 41600 29772
rect 41520 29452 41532 29508
rect 41588 29452 41600 29508
rect 41520 29440 41600 29452
rect 41680 29828 41760 29840
rect 41680 29772 41692 29828
rect 41748 29772 41760 29828
rect 41680 29508 41760 29772
rect 41680 29452 41692 29508
rect 41748 29452 41760 29508
rect 41680 29440 41760 29452
rect 41840 29828 41920 29840
rect 41840 29772 41852 29828
rect 41908 29772 41920 29828
rect 41840 29508 41920 29772
rect 41840 29452 41852 29508
rect 41908 29452 41920 29508
rect 41840 29440 41920 29452
<< metal4 >>
rect 0 70480 80 70880
rect 20880 70480 21040 70880
rect 0 70000 80 70400
rect 20880 70000 21040 70400
rect 0 69520 80 69920
rect 20880 69520 21040 69920
rect 0 69040 80 69440
rect 20880 69040 21040 69440
rect 20880 -2640 21040 -2240
rect 20880 -3120 21040 -2720
rect 20880 -3600 21040 -3200
rect 20880 -4080 21040 -3680
<< metal5 >>
rect 160 29440 560 37360
rect 1120 29440 1520 37360
rect 2080 29440 2480 37360
rect 3040 29440 3440 37360
rect 4000 29440 4400 37360
rect 4960 29440 5360 37360
rect 5920 29440 6320 37360
rect 6880 29440 7280 37360
rect 7840 29440 8240 37360
rect 12640 29440 13040 37360
rect 13600 29440 14000 37360
rect 14560 29440 14960 37360
rect 15520 29440 15920 37360
rect 16480 29440 16880 37360
rect 17440 29440 17840 37360
rect 18400 29440 18800 37360
rect 19360 29440 19760 37360
rect 20320 29440 20720 37360
rect 21200 29440 21600 37360
rect 22160 29440 22560 37360
rect 23120 29440 23520 37360
rect 24080 29440 24480 37360
rect 25040 29440 25440 37360
rect 26000 29440 26400 37360
rect 26960 29440 27360 37360
rect 27920 29440 28320 37360
rect 28880 29440 29280 37360
rect 33680 29440 34080 37360
rect 34640 29440 35040 37360
rect 35600 29440 36000 37360
rect 36560 29440 36960 37360
rect 37520 29440 37920 37360
rect 38480 29440 38880 37360
rect 39440 29440 39840 37360
rect 40400 29440 40800 37360
rect 41360 29440 41760 37360
use ota_core  4
timestamp 1638148091
transform 1 0 21040 0 1 -2160
box -26 -4640 20906 31600
use ota_core  3
timestamp 1638148091
transform -1 0 20880 0 1 -2160
box -26 -4640 20906 31600
use ota_core  2
timestamp 1638148091
transform -1 0 41920 0 -1 68960
box -26 -4640 20906 31600
use ota_core  1
timestamp 1638148091
transform 1 0 0 0 -1 68960
box -26 -4640 20906 31600
<< labels >>
rlabel metal2 s 0 36640 80 36720 4 bp
rlabel metal2 s 0 35520 80 35600 4 x
rlabel metal2 s 0 35200 80 35280 4 y
rlabel metal4 s 0 69520 80 69920 4 vddx
rlabel metal3 s 11680 37360 11760 37440 4 z
rlabel metal2 s 0 32160 80 32240 4 im
port 1 nsew
rlabel metal2 s 0 36160 80 36240 4 ip
port 2 nsew
rlabel metal2 s 0 31840 80 31920 4 op
port 3 nsew
rlabel metal2 s 0 35840 80 35920 4 om
port 4 nsew
rlabel metal2 s 0 37120 80 37200 4 ib
port 5 nsew
rlabel metal2 s 0 33600 80 33680 4 q
port 6 nsew
rlabel metal4 s 0 69040 80 69440 4 vdda
port 7 nsew
rlabel metal4 s 0 70000 80 70400 4 gnda
port 8 nsew
rlabel metal4 s 0 70480 80 70880 4 vssa
port 9 nsew
<< end >>
