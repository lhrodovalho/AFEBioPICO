* SPICE3 file created from n1_8.ext - technology: sky130A

.option scale=10000u

.subckt n1_8 D G S B
X0 a1 G S B sky130_fd_pr__nfet_01v8_lvt ad=10000 pd=600 as=5000 ps=300 w=100 l=800
X1 a5 G a4 B sky130_fd_pr__nfet_01v8_lvt ad=10000 pd=600 as=10000 ps=600 w=100 l=800
X2 a3 G a2 B sky130_fd_pr__nfet_01v8_lvt ad=10000 pd=600 as=10000 ps=600 w=100 l=800
X3 a1 G a2 B sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=100 l=800
X4 a7 G D B sky130_fd_pr__nfet_01v8_lvt ad=10000 pd=600 as=5000 ps=300 w=100 l=800
X5 a5 G a6 B sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=10000 ps=600 w=100 l=800
X6 a3 G a4 B sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=100 l=800
X7 a7 G a6 B sky130_fd_pr__nfet_01v8_lvt ad=0 pd=0 as=0 ps=0 w=100 l=800
.ends
