magic
tech sky130A
magscale 1 2
timestamp 1634662791
<< nwell >>
rect -5740 -6580 -5640 -920
rect 47000 -6580 47100 -920
<< pwell >>
rect -5820 -880 -5640 -820
rect 47000 -880 47180 -820
rect -5840 -10300 -5620 -10240
rect 47000 -10300 47200 -10240
rect -5840 -12560 -5780 -10300
rect 47140 -12560 47200 -10300
<< psubdiff >>
rect -5840 -880 -5640 -820
rect 47000 -880 47200 -820
rect -5840 -6620 -5780 -880
rect 47140 -6620 47200 -880
rect -5840 -6680 -3620 -6620
rect 20540 -6680 20820 -6620
rect 44980 -6680 47200 -6620
rect -5840 -10240 -5780 -6680
rect 47140 -10240 47200 -6680
rect -5840 -10300 -5620 -10240
rect 47000 -10300 47200 -10240
rect -5840 -12560 -5780 -10300
rect 47140 -12560 47200 -10300
rect -5840 -12620 47200 -12560
<< psubdiffcont >>
rect -3620 -6680 20540 -6620
rect 20820 -6680 44980 -6620
<< locali >>
rect -12400 -8240 -12060 -440
rect -12000 -8240 -11660 -440
rect -11620 -8240 -11280 -440
rect -11220 -8240 -10880 -440
rect -10820 -8240 -10480 -440
rect -10420 -8240 -10100 -440
rect -10040 -8240 -9320 -440
rect -9260 -8240 -8920 -440
rect -8860 -8240 -8520 -440
rect -8480 -8240 -8140 -440
rect -8080 -8240 -7740 -440
rect -7700 -8240 -7360 -440
rect -7300 -6800 -6960 -440
rect -5840 -880 -5640 -820
rect 47000 -880 47200 -820
rect -5840 -6620 -5780 -880
rect -2020 -960 -1920 -940
rect -5700 -6540 -5640 -960
rect -2020 -1020 -2000 -960
rect -1940 -1020 -1920 -960
rect -2020 -1040 -1920 -1020
rect 43280 -960 43380 -940
rect 43280 -1020 43300 -960
rect 43360 -1020 43380 -960
rect 43280 -1040 43380 -1020
rect 47000 -6540 47060 -960
rect 47140 -6620 47200 -880
rect -5840 -6680 -3700 -6620
rect -3640 -6680 -3620 -6620
rect 20540 -6680 20820 -6620
rect 44980 -6680 45000 -6620
rect 45060 -6680 47200 -6620
rect -7300 -6980 47120 -6800
rect -7300 -7040 -6960 -6980
rect -7300 -7220 47120 -7040
rect -7300 -7280 -6960 -7220
rect -7300 -7460 47120 -7280
rect -7300 -7520 -6960 -7460
rect -7300 -7700 47120 -7520
rect -7300 -7760 -6960 -7700
rect -7300 -7940 47120 -7760
rect -7300 -8000 -6960 -7940
rect -7300 -8180 47120 -8000
rect -7300 -8240 -6960 -8180
rect -12400 -8300 48840 -8240
rect -12400 -8620 -3580 -8300
rect -3520 -8620 44880 -8300
rect 44940 -8320 48840 -8300
rect 44940 -8600 48540 -8320
rect 48820 -8600 48840 -8320
rect 44940 -8620 48840 -8600
rect -12400 -8660 48840 -8620
rect -12400 -13000 -12060 -8660
rect -12000 -13000 -11660 -8660
rect -11620 -13000 -11280 -8660
rect -11220 -13000 -10880 -8660
rect -10820 -13000 -10480 -8660
rect -10420 -13000 -10100 -8660
rect -10040 -13000 -9320 -8660
rect -9260 -13000 -8920 -8660
rect -8860 -13000 -8520 -8660
rect -8480 -13000 -8140 -8660
rect -8080 -13000 -7740 -8660
rect -7700 -13000 -7360 -8660
rect -7300 -8680 48840 -8660
rect -7300 -8740 -6960 -8680
rect -7300 -8920 47120 -8740
rect -7300 -8980 -6960 -8920
rect -7300 -9160 47120 -8980
rect -7300 -9220 -6960 -9160
rect -7300 -9400 47120 -9220
rect -7300 -9460 -6960 -9400
rect -7300 -9640 47120 -9460
rect -7300 -9700 -6960 -9640
rect -7300 -9880 47120 -9700
rect -7300 -9940 -6960 -9880
rect -7300 -10120 47120 -9940
rect -7300 -13000 -6960 -10120
rect -5840 -10300 -5620 -10240
rect 47000 -10300 47200 -10240
rect -5840 -12560 -5780 -10300
rect -3720 -12560 -3620 -12540
rect 44980 -12560 45080 -12540
rect 47140 -12560 47200 -10300
rect -5840 -12620 -3700 -12560
rect -3640 -12620 45000 -12560
rect 45060 -12620 47200 -12560
rect -3720 -12640 -3620 -12620
rect 44980 -12640 45080 -12620
<< viali >>
rect -2000 -1020 -1940 -960
rect 43300 -1020 43360 -960
rect -3700 -6680 -3640 -6620
rect 45000 -6680 45060 -6620
rect -3580 -8620 -3520 -8300
rect 44880 -8620 44940 -8300
rect 48540 -8600 48820 -8320
rect -3700 -12620 -3640 -12560
rect 45000 -12620 45060 -12560
<< metal1 >>
rect -12460 -10120 -12400 -440
rect -12460 -13000 -12400 -10180
rect -12060 -10120 -12000 -440
rect -12060 -13000 -12000 -10180
rect -11680 -10120 -11620 -440
rect -11680 -13000 -11620 -10180
rect -11280 -10120 -11220 -440
rect -11280 -13000 -11220 -10180
rect -10880 -10120 -10820 -440
rect -10880 -13000 -10820 -10180
rect -10480 -10120 -10420 -440
rect -10480 -13000 -10420 -10180
rect -10100 -10120 -10040 -440
rect -10100 -13000 -10040 -10180
rect -9320 -10120 -9260 -440
rect -9320 -13000 -9260 -10180
rect -8920 -10120 -8860 -440
rect -8920 -13000 -8860 -10180
rect -8540 -10120 -8480 -440
rect -8540 -13000 -8480 -10180
rect -8140 -10120 -8080 -440
rect -8140 -13000 -8080 -10180
rect -7760 -10120 -7700 -440
rect -7760 -13000 -7700 -10180
rect -7360 -10120 -7300 -440
rect -7360 -13000 -7300 -10180
rect -6960 -10120 -6900 -440
rect -5580 -460 -5520 -440
rect -5580 -6720 -5520 -740
rect -3880 -460 -3820 -440
rect -3880 -780 -3820 -740
rect -2000 -460 -1940 -440
rect -2000 -780 -1940 -740
rect 1760 -460 1820 -440
rect 1760 -900 1820 -740
rect 3640 -460 3700 -440
rect 3640 -900 3700 -740
rect 7400 -460 7460 -440
rect 7400 -780 7460 -740
rect 11160 -460 11220 -440
rect 11160 -780 11220 -740
rect 14920 -460 14980 -440
rect 14920 -780 14980 -740
rect 20560 -460 20620 -440
rect 20560 -780 20620 -740
rect 20740 -460 20800 -440
rect 20740 -780 20800 -740
rect 26380 -460 26440 -440
rect 26380 -780 26440 -740
rect 30140 -460 30200 -440
rect 30140 -780 30200 -740
rect 33900 -460 33960 -440
rect 33900 -780 33960 -740
rect 37660 -460 37720 -440
rect 37660 -900 37720 -740
rect 39540 -460 39600 -440
rect 39540 -900 39600 -740
rect 43300 -460 43360 -440
rect 43300 -780 43360 -740
rect 45180 -460 45240 -440
rect 45180 -780 45240 -740
rect 46880 -460 46940 -440
rect -2020 -960 -1920 -940
rect -2020 -1020 -2000 -960
rect -1940 -1020 -1920 -960
rect -2020 -1040 -1920 -1020
rect 43280 -960 43380 -940
rect 43280 -1020 43300 -960
rect 43360 -1020 43380 -960
rect 43280 -1040 43380 -1020
rect 46880 -1080 46940 -740
rect -3720 -6620 -3620 -6600
rect -3720 -6680 -3700 -6620
rect -3640 -6680 -3620 -6620
rect -3720 -6700 -3620 -6680
rect -5340 -6860 -5280 -6720
rect -5340 -6940 -5280 -6920
rect -6960 -13000 -6900 -10180
rect -4120 -10000 -4060 -9980
rect -5580 -12700 -5520 -10200
rect -4120 -10220 -4060 -10060
rect -5580 -13000 -5520 -12980
rect -3880 -12700 -3820 -10200
rect -3700 -12540 -3640 -6700
rect -3580 -6740 -3520 -6720
rect -3580 -6980 -3520 -6800
rect -3460 -6860 -3400 -6720
rect -3460 -6940 -3400 -6920
rect -2000 -6860 -1940 -6720
rect -2000 -6940 -1940 -6920
rect -3580 -7220 -3520 -7040
rect -1820 -7100 -1760 -6720
rect -1820 -7180 -1760 -7160
rect -1580 -7100 -1520 -6720
rect -120 -6860 -60 -6300
rect 3640 -6320 3700 -6300
rect -120 -6940 -60 -6920
rect 300 -6860 360 -6720
rect 300 -6940 360 -6920
rect -1580 -7180 -1520 -7160
rect -3580 -7460 -3520 -7280
rect -3580 -7700 -3520 -7520
rect -3580 -7940 -3520 -7760
rect -3580 -8180 -3520 -8000
rect -3580 -8280 -3520 -8240
rect -3600 -8300 -3500 -8280
rect -3600 -8620 -3580 -8300
rect -3520 -8620 -3500 -8300
rect -3600 -8640 -3500 -8620
rect -3580 -8680 -3520 -8640
rect -3580 -8920 -3520 -8740
rect -3580 -9160 -3520 -8980
rect -3580 -9400 -3520 -9220
rect -3580 -9640 -3520 -9460
rect -3580 -9880 -3520 -9700
rect -3580 -10120 -3520 -9940
rect 1520 -9760 1580 -9740
rect -3580 -10200 -3520 -10180
rect -2240 -10000 -2180 -9980
rect -2240 -10200 -2180 -10060
rect -1820 -10000 -1760 -9980
rect -1820 -10200 -1760 -10060
rect -360 -10000 -300 -9980
rect -360 -10200 -300 -10060
rect 60 -10000 120 -9980
rect 60 -10480 120 -10060
rect 1520 -10200 1580 -9820
rect 1760 -9760 1820 -6720
rect 2180 -6860 2240 -6720
rect 2180 -6940 2240 -6920
rect 3640 -7340 3700 -6720
rect 3640 -7420 3700 -7400
rect 3820 -7340 3880 -6720
rect 3820 -7420 3880 -7400
rect 4060 -7580 4120 -6720
rect 4060 -7660 4120 -7640
rect 1760 -10200 1820 -9820
rect 1940 -8060 2000 -8040
rect 1940 -10200 2000 -8120
rect 3820 -8060 3880 -8040
rect 3400 -9040 3460 -9020
rect 3400 -10200 3460 -9100
rect 3820 -10480 3880 -8120
rect 5520 -8060 5580 -6300
rect 5940 -6860 6000 -6720
rect 5940 -6940 6000 -6920
rect 7400 -7340 7460 -6720
rect 7400 -7420 7460 -7400
rect 7580 -7340 7640 -6720
rect 7580 -7420 7640 -7400
rect 7820 -7820 7880 -6700
rect 7820 -7900 7880 -7880
rect 5520 -8140 5580 -8120
rect 5700 -8800 5760 -8780
rect 5280 -9040 5340 -9020
rect 5280 -10200 5340 -9100
rect 5520 -9040 5580 -9020
rect 5520 -10200 5580 -9100
rect 5700 -10200 5760 -8860
rect 7580 -8800 7640 -8780
rect 7160 -9040 7220 -9020
rect 7160 -10200 7220 -9100
rect 7580 -10480 7640 -8860
rect 9280 -8800 9340 -6300
rect 9700 -6860 9760 -6720
rect 9700 -6940 9760 -6920
rect 9280 -8880 9340 -8860
rect 9460 -8800 9520 -8780
rect 9040 -9040 9100 -9020
rect 9040 -10200 9100 -9100
rect 9280 -9520 9340 -9500
rect 9280 -10200 9340 -9580
rect 9460 -10200 9520 -8860
rect 10920 -9040 10980 -9020
rect 10920 -10200 10980 -9100
rect 11160 -9040 11220 -6720
rect 11340 -7340 11400 -6720
rect 11340 -7420 11400 -7400
rect 11580 -7820 11640 -6720
rect 11580 -7900 11640 -7880
rect 11160 -9120 11220 -9100
rect 11340 -8800 11400 -8780
rect 11340 -10480 11400 -8860
rect 13040 -8800 13100 -6300
rect 13460 -6860 13520 -6720
rect 13460 -6940 13520 -6920
rect 13040 -8880 13100 -8860
rect 13220 -8060 13280 -8040
rect 12800 -9040 12860 -9020
rect 12800 -10200 12860 -9100
rect 13040 -9520 13100 -9500
rect 13040 -10200 13100 -9580
rect 13220 -10200 13280 -8120
rect 14680 -9040 14740 -9020
rect 14680 -10200 14740 -9100
rect 14920 -9280 14980 -6720
rect 15100 -7340 15160 -6720
rect 15100 -7420 15160 -7400
rect 15340 -7580 15400 -6720
rect 15340 -7660 15400 -7640
rect 14920 -9360 14980 -9340
rect 15100 -8060 15160 -8040
rect 15100 -10480 15160 -8120
rect 16800 -8060 16860 -6300
rect 16800 -8140 16860 -8120
rect 16560 -9040 16620 -9020
rect 16560 -10200 16620 -9100
rect 16800 -9040 16860 -9020
rect 16800 -10200 16860 -9100
rect 16980 -9280 17040 -6720
rect 17220 -7100 17280 -6720
rect 17220 -7180 17280 -7160
rect 16980 -10480 17040 -9340
rect 18680 -9520 18740 -6300
rect 18860 -8320 18920 -6720
rect 18860 -8620 18920 -8600
rect 19100 -9280 19160 -6720
rect 19100 -9360 19160 -9340
rect 20560 -8320 20620 -8300
rect 18440 -9760 18500 -9740
rect 18440 -10200 18500 -9820
rect 18680 -10200 18740 -9580
rect 20320 -9520 20380 -9500
rect 20320 -10200 20380 -9580
rect 20560 -10200 20620 -8600
rect 20740 -8320 20800 -8300
rect 20740 -10200 20800 -8600
rect 22200 -9280 22260 -6720
rect 22440 -8320 22500 -6720
rect 22440 -8620 22500 -8600
rect 22200 -9360 22260 -9340
rect 20980 -9520 21040 -9500
rect 20980 -10200 21040 -9580
rect 22620 -9520 22680 -6300
rect 24080 -7100 24140 -6720
rect 24080 -7180 24140 -7160
rect 22620 -10200 22680 -9580
rect 24320 -9280 24380 -6720
rect 24500 -8060 24560 -6300
rect 25960 -7580 26020 -6720
rect 26200 -7340 26260 -6720
rect 26200 -7420 26260 -7400
rect 25960 -7660 26020 -7640
rect 24500 -8140 24560 -8120
rect 26200 -8060 26260 -8040
rect 22860 -9760 22920 -9740
rect 22860 -10200 22920 -9820
rect 24320 -10480 24380 -9340
rect 24500 -9040 24560 -9020
rect 24500 -10200 24560 -9100
rect 24740 -9040 24800 -9020
rect 24740 -10200 24800 -9100
rect 26200 -10480 26260 -8120
rect 26380 -9280 26440 -6720
rect 27840 -6860 27900 -6720
rect 27840 -6940 27900 -6920
rect 28080 -8060 28140 -8040
rect 26380 -9360 26440 -9340
rect 26620 -9040 26680 -9020
rect 26620 -10200 26680 -9100
rect 28080 -10200 28140 -8120
rect 28260 -8800 28320 -6300
rect 29720 -7820 29780 -6720
rect 29960 -7340 30020 -6720
rect 29960 -7420 30020 -7400
rect 29720 -7900 29780 -7880
rect 28260 -8880 28320 -8860
rect 29960 -8800 30020 -8780
rect 28500 -9040 28560 -9020
rect 28260 -9520 28320 -9500
rect 28260 -10200 28320 -9580
rect 28500 -10200 28560 -9100
rect 29960 -10480 30020 -8860
rect 30140 -9040 30200 -6720
rect 31600 -6860 31660 -6720
rect 31600 -6940 31660 -6920
rect 31840 -8800 31900 -8780
rect 30140 -9120 30200 -9100
rect 30380 -9040 30440 -9020
rect 30380 -10200 30440 -9100
rect 31840 -10200 31900 -8860
rect 32020 -8800 32080 -6300
rect 33480 -7820 33540 -6700
rect 33720 -7340 33780 -6720
rect 33720 -7420 33780 -7400
rect 33900 -7340 33960 -6720
rect 35360 -6860 35420 -6720
rect 35360 -6940 35420 -6920
rect 33900 -7420 33960 -7400
rect 33480 -7900 33540 -7880
rect 35780 -8060 35840 -6300
rect 37660 -6320 37720 -6300
rect 37240 -7580 37300 -6720
rect 37480 -7340 37540 -6720
rect 37480 -7420 37540 -7400
rect 37660 -7340 37720 -6720
rect 39120 -6860 39180 -6720
rect 39120 -6940 39180 -6920
rect 37660 -7420 37720 -7400
rect 37240 -7660 37300 -7640
rect 35780 -8140 35840 -8120
rect 37480 -8060 37540 -8040
rect 32020 -8880 32080 -8860
rect 33720 -8800 33780 -8780
rect 32260 -9040 32320 -9020
rect 32020 -9520 32080 -9500
rect 32020 -10200 32080 -9580
rect 32260 -10200 32320 -9100
rect 33720 -10480 33780 -8860
rect 35600 -8800 35660 -8780
rect 34140 -9040 34200 -9020
rect 34140 -10200 34200 -9100
rect 35600 -10200 35660 -8860
rect 35780 -9040 35840 -9020
rect 35780 -10200 35840 -9100
rect 36020 -9040 36080 -9020
rect 36020 -10200 36080 -9100
rect 37480 -10480 37540 -8120
rect 39360 -8060 39420 -8040
rect 37900 -9040 37960 -9020
rect 37900 -10200 37960 -9100
rect 39360 -10200 39420 -8120
rect 39540 -9760 39600 -6720
rect 41000 -6860 41060 -6720
rect 41000 -6940 41060 -6920
rect 41420 -6860 41480 -6300
rect 44980 -6620 45080 -6600
rect 44980 -6680 45000 -6620
rect 45060 -6680 45080 -6620
rect 44980 -6700 45080 -6680
rect 41420 -6940 41480 -6920
rect 42880 -7100 42940 -6720
rect 42880 -7180 42940 -7160
rect 43120 -7100 43180 -6720
rect 43300 -6860 43360 -6720
rect 43300 -6940 43360 -6920
rect 44760 -6860 44820 -6720
rect 44760 -6940 44820 -6920
rect 44880 -6740 44940 -6720
rect 43120 -7180 43180 -7160
rect 44880 -6980 44940 -6800
rect 44880 -7220 44940 -7040
rect 44880 -7460 44940 -7280
rect 44880 -7700 44940 -7520
rect 44880 -7940 44940 -7760
rect 44880 -8180 44940 -8000
rect 44880 -8280 44940 -8240
rect 44860 -8300 44960 -8280
rect 44860 -8620 44880 -8300
rect 44940 -8620 44960 -8300
rect 44860 -8640 44960 -8620
rect 44880 -8680 44940 -8640
rect 44880 -8920 44940 -8740
rect 44880 -9160 44940 -8980
rect 44880 -9400 44940 -9220
rect 44880 -9640 44940 -9460
rect 39540 -10200 39600 -9820
rect 39780 -9760 39840 -9740
rect 39780 -10200 39840 -9820
rect 44880 -9880 44940 -9700
rect 41240 -10000 41300 -9980
rect 41240 -10480 41300 -10060
rect 41660 -10000 41720 -9980
rect 41660 -10200 41720 -10060
rect 43120 -10000 43180 -9980
rect 43120 -10200 43180 -10060
rect 43540 -10000 43600 -9980
rect 43540 -10200 43600 -10060
rect 44880 -10120 44940 -9940
rect 44880 -10200 44940 -10180
rect 45000 -12540 45060 -6700
rect 46640 -6860 46700 -6660
rect 46640 -6940 46700 -6920
rect 48520 -8320 48840 -8300
rect 48520 -8600 48540 -8320
rect 48820 -8600 48840 -8320
rect 48520 -8620 48840 -8600
rect 45420 -10000 45480 -9980
rect 45420 -10200 45480 -10060
rect -3720 -12560 -3620 -12540
rect -3720 -12620 -3700 -12560
rect -3640 -12620 -3620 -12560
rect -3720 -12640 -3620 -12620
rect 44980 -12560 45080 -12540
rect 44980 -12620 45000 -12560
rect 45060 -12620 45080 -12560
rect 44980 -12640 45080 -12620
rect -3880 -13000 -3820 -12980
rect -3700 -12700 -3640 -12640
rect -3700 -13000 -3640 -12980
rect -1820 -12700 -1760 -12660
rect -1820 -13000 -1760 -12980
rect 1940 -12700 2000 -12660
rect 1940 -13000 2000 -12980
rect 5700 -12700 5760 -12660
rect 5700 -13000 5760 -12980
rect 9460 -12700 9520 -12660
rect 9460 -13000 9520 -12980
rect 13220 -12700 13280 -12660
rect 13220 -13000 13280 -12980
rect 18860 -12700 18920 -12660
rect 18860 -13000 18920 -12980
rect 22440 -12700 22500 -12660
rect 22440 -13000 22500 -12980
rect 28080 -12700 28140 -12660
rect 28080 -13000 28140 -12980
rect 31840 -12700 31900 -12660
rect 31840 -13000 31900 -12980
rect 35600 -12700 35660 -12660
rect 35600 -13000 35660 -12980
rect 39360 -12700 39420 -12660
rect 39360 -13000 39420 -12980
rect 43120 -12700 43180 -12660
rect 43120 -13000 43180 -12980
rect 45000 -12700 45060 -12640
rect 45000 -13000 45060 -12980
rect 45180 -12700 45240 -12500
rect 45180 -13000 45240 -12980
rect 46880 -12700 46940 -12660
rect 46880 -13000 46940 -12980
<< via1 >>
rect -12460 -10180 -12400 -10120
rect -12060 -10180 -12000 -10120
rect -11680 -10180 -11620 -10120
rect -11280 -10180 -11220 -10120
rect -10880 -10180 -10820 -10120
rect -10480 -10180 -10420 -10120
rect -10100 -10180 -10040 -10120
rect -9320 -10180 -9260 -10120
rect -8920 -10180 -8860 -10120
rect -8540 -10180 -8480 -10120
rect -8140 -10180 -8080 -10120
rect -7760 -10180 -7700 -10120
rect -7360 -10180 -7300 -10120
rect -5580 -740 -5520 -460
rect -3880 -740 -3820 -460
rect -2000 -740 -1940 -460
rect 1760 -740 1820 -460
rect 3640 -740 3700 -460
rect 7400 -740 7460 -460
rect 11160 -740 11220 -460
rect 14920 -740 14980 -460
rect 20560 -740 20620 -460
rect 20740 -740 20800 -460
rect 26380 -740 26440 -460
rect 30140 -740 30200 -460
rect 33900 -740 33960 -460
rect 37660 -740 37720 -460
rect 39540 -740 39600 -460
rect 43300 -740 43360 -460
rect 45180 -740 45240 -460
rect 46880 -740 46940 -460
rect -5340 -6920 -5280 -6860
rect -6960 -10180 -6900 -10120
rect -4120 -10060 -4060 -10000
rect -5580 -12980 -5520 -12700
rect -3580 -6800 -3520 -6740
rect -3460 -6920 -3400 -6860
rect -2000 -6920 -1940 -6860
rect -3580 -7040 -3520 -6980
rect -1820 -7160 -1760 -7100
rect -120 -6920 -60 -6860
rect 300 -6920 360 -6860
rect -1580 -7160 -1520 -7100
rect -3580 -7280 -3520 -7220
rect -3580 -7520 -3520 -7460
rect -3580 -7760 -3520 -7700
rect -3580 -8000 -3520 -7940
rect -3580 -8240 -3520 -8180
rect -3580 -8740 -3520 -8680
rect -3580 -8980 -3520 -8920
rect -3580 -9220 -3520 -9160
rect -3580 -9460 -3520 -9400
rect -3580 -9700 -3520 -9640
rect -3580 -9940 -3520 -9880
rect 1520 -9820 1580 -9760
rect -3580 -10180 -3520 -10120
rect -2240 -10060 -2180 -10000
rect -1820 -10060 -1760 -10000
rect -360 -10060 -300 -10000
rect 60 -10060 120 -10000
rect 2180 -6920 2240 -6860
rect 3640 -7400 3700 -7340
rect 3820 -7400 3880 -7340
rect 4060 -7640 4120 -7580
rect 1760 -9820 1820 -9760
rect 1940 -8120 2000 -8060
rect 3820 -8120 3880 -8060
rect 3400 -9100 3460 -9040
rect 5940 -6920 6000 -6860
rect 7400 -7400 7460 -7340
rect 7580 -7400 7640 -7340
rect 7820 -7880 7880 -7820
rect 5520 -8120 5580 -8060
rect 5700 -8860 5760 -8800
rect 5280 -9100 5340 -9040
rect 5520 -9100 5580 -9040
rect 7580 -8860 7640 -8800
rect 7160 -9100 7220 -9040
rect 9700 -6920 9760 -6860
rect 9280 -8860 9340 -8800
rect 9460 -8860 9520 -8800
rect 9040 -9100 9100 -9040
rect 9280 -9580 9340 -9520
rect 10920 -9100 10980 -9040
rect 11340 -7400 11400 -7340
rect 11580 -7880 11640 -7820
rect 11160 -9100 11220 -9040
rect 11340 -8860 11400 -8800
rect 13460 -6920 13520 -6860
rect 13040 -8860 13100 -8800
rect 13220 -8120 13280 -8060
rect 12800 -9100 12860 -9040
rect 13040 -9580 13100 -9520
rect 14680 -9100 14740 -9040
rect 15100 -7400 15160 -7340
rect 15340 -7640 15400 -7580
rect 14920 -9340 14980 -9280
rect 15100 -8120 15160 -8060
rect 16800 -8120 16860 -8060
rect 16560 -9100 16620 -9040
rect 16800 -9100 16860 -9040
rect 17220 -7160 17280 -7100
rect 16980 -9340 17040 -9280
rect 18860 -8600 18920 -8320
rect 19100 -9340 19160 -9280
rect 20560 -8600 20620 -8320
rect 18680 -9580 18740 -9520
rect 18440 -9820 18500 -9760
rect 20320 -9580 20380 -9520
rect 20740 -8600 20800 -8320
rect 22440 -8600 22500 -8320
rect 22200 -9340 22260 -9280
rect 20980 -9580 21040 -9520
rect 24080 -7160 24140 -7100
rect 22620 -9580 22680 -9520
rect 26200 -7400 26260 -7340
rect 25960 -7640 26020 -7580
rect 24500 -8120 24560 -8060
rect 26200 -8120 26260 -8060
rect 24320 -9340 24380 -9280
rect 22860 -9820 22920 -9760
rect 24500 -9100 24560 -9040
rect 24740 -9100 24800 -9040
rect 27840 -6920 27900 -6860
rect 28080 -8120 28140 -8060
rect 26380 -9340 26440 -9280
rect 26620 -9100 26680 -9040
rect 29960 -7400 30020 -7340
rect 29720 -7880 29780 -7820
rect 28260 -8860 28320 -8800
rect 29960 -8860 30020 -8800
rect 28500 -9100 28560 -9040
rect 28260 -9580 28320 -9520
rect 31600 -6920 31660 -6860
rect 31840 -8860 31900 -8800
rect 30140 -9100 30200 -9040
rect 30380 -9100 30440 -9040
rect 33720 -7400 33780 -7340
rect 35360 -6920 35420 -6860
rect 33900 -7400 33960 -7340
rect 33480 -7880 33540 -7820
rect 37480 -7400 37540 -7340
rect 39120 -6920 39180 -6860
rect 37660 -7400 37720 -7340
rect 37240 -7640 37300 -7580
rect 35780 -8120 35840 -8060
rect 37480 -8120 37540 -8060
rect 32020 -8860 32080 -8800
rect 33720 -8860 33780 -8800
rect 32260 -9100 32320 -9040
rect 32020 -9580 32080 -9520
rect 35600 -8860 35660 -8800
rect 34140 -9100 34200 -9040
rect 35780 -9100 35840 -9040
rect 36020 -9100 36080 -9040
rect 39360 -8120 39420 -8060
rect 37900 -9100 37960 -9040
rect 41000 -6920 41060 -6860
rect 41420 -6920 41480 -6860
rect 42880 -7160 42940 -7100
rect 43300 -6920 43360 -6860
rect 44760 -6920 44820 -6860
rect 44880 -6800 44940 -6740
rect 43120 -7160 43180 -7100
rect 44880 -7040 44940 -6980
rect 44880 -7280 44940 -7220
rect 44880 -7520 44940 -7460
rect 44880 -7760 44940 -7700
rect 44880 -8000 44940 -7940
rect 44880 -8240 44940 -8180
rect 44880 -8740 44940 -8680
rect 44880 -8980 44940 -8920
rect 44880 -9220 44940 -9160
rect 44880 -9460 44940 -9400
rect 44880 -9700 44940 -9640
rect 39540 -9820 39600 -9760
rect 39780 -9820 39840 -9760
rect 44880 -9940 44940 -9880
rect 41240 -10060 41300 -10000
rect 41660 -10060 41720 -10000
rect 43120 -10060 43180 -10000
rect 43540 -10060 43600 -10000
rect 44880 -10180 44940 -10120
rect 46640 -6920 46700 -6860
rect 48540 -8600 48820 -8320
rect 45420 -10060 45480 -10000
rect -3880 -12980 -3820 -12700
rect -3700 -12980 -3640 -12700
rect -1820 -12980 -1760 -12700
rect 1940 -12980 2000 -12700
rect 5700 -12980 5760 -12700
rect 9460 -12980 9520 -12700
rect 13220 -12980 13280 -12700
rect 18860 -12980 18920 -12700
rect 22440 -12980 22500 -12700
rect 28080 -12980 28140 -12700
rect 31840 -12980 31900 -12700
rect 35600 -12980 35660 -12700
rect 39360 -12980 39420 -12700
rect 43120 -12980 43180 -12700
rect 45000 -12980 45060 -12700
rect 45180 -12980 45240 -12700
rect 46880 -12980 46940 -12700
<< metal2 >>
rect 18240 480 18340 490
rect 18240 370 18340 380
rect -6840 -460 48840 -440
rect -6840 -740 -6820 -460
rect -6540 -740 -5580 -460
rect -5520 -740 -3880 -460
rect -3820 -740 -2000 -460
rect -1940 -740 1760 -460
rect 1820 -740 3640 -460
rect 3700 -740 7400 -460
rect 7460 -740 11160 -460
rect 11220 -740 14920 -460
rect 14980 -740 20560 -460
rect 20620 -740 20740 -460
rect 20800 -740 26380 -460
rect 26440 -740 30140 -460
rect 30200 -740 33900 -460
rect 33960 -740 37660 -460
rect 37720 -740 39540 -460
rect 39600 -740 43300 -460
rect 43360 -740 45180 -460
rect 45240 -740 46880 -460
rect 46940 -740 47900 -460
rect 48180 -740 48840 -460
rect -6840 -760 48840 -740
rect -12460 -6800 -3580 -6740
rect -3520 -6800 44880 -6740
rect 44940 -6800 47240 -6740
rect -12280 -6860 -12180 -6840
rect -12460 -6920 -12260 -6860
rect -12200 -6920 -5340 -6860
rect -5280 -6920 -3460 -6860
rect -3400 -6920 -2000 -6860
rect -1940 -6920 -120 -6860
rect -60 -6920 300 -6860
rect 360 -6920 2180 -6860
rect 2240 -6920 5940 -6860
rect 6000 -6920 9700 -6860
rect 9760 -6920 13460 -6860
rect 13520 -6920 27840 -6860
rect 27900 -6920 31600 -6860
rect 31660 -6920 35360 -6860
rect 35420 -6920 39120 -6860
rect 39180 -6920 41000 -6860
rect 41060 -6920 41420 -6860
rect 41480 -6920 43300 -6860
rect 43360 -6920 44760 -6860
rect 44820 -6920 46640 -6860
rect 46700 -6920 47240 -6860
rect -12280 -6940 -12180 -6920
rect -12460 -7040 -3580 -6980
rect -3520 -7040 44880 -6980
rect 44940 -7040 47240 -6980
rect -11880 -7100 -11780 -7080
rect -12460 -7160 -11860 -7100
rect -11800 -7160 -1820 -7100
rect -1760 -7160 -1580 -7100
rect -1520 -7160 17220 -7100
rect 17280 -7160 24080 -7100
rect 24140 -7160 42880 -7100
rect 42940 -7160 43120 -7100
rect 43180 -7160 47240 -7100
rect -11880 -7180 -11780 -7160
rect -12460 -7280 -3580 -7220
rect -3520 -7280 44880 -7220
rect 44940 -7280 47240 -7220
rect -11500 -7340 -11400 -7320
rect -12460 -7400 -11480 -7340
rect -11420 -7400 3640 -7340
rect 3700 -7400 3820 -7340
rect 3880 -7400 7400 -7340
rect 7460 -7400 7580 -7340
rect 7640 -7400 11340 -7340
rect 11400 -7400 15100 -7340
rect 15160 -7400 26200 -7340
rect 26260 -7400 29960 -7340
rect 30020 -7400 33720 -7340
rect 33780 -7400 33900 -7340
rect 33960 -7400 37480 -7340
rect 37540 -7400 37660 -7340
rect 37720 -7400 47240 -7340
rect -11500 -7420 -11400 -7400
rect -12460 -7520 -3580 -7460
rect -3520 -7520 44880 -7460
rect 44940 -7520 47240 -7460
rect -11100 -7580 -11000 -7560
rect -12480 -7640 -11080 -7580
rect -11020 -7640 4060 -7580
rect 4120 -7640 15340 -7580
rect 15400 -7640 25960 -7580
rect 26020 -7640 37240 -7580
rect 37300 -7640 47240 -7580
rect -11100 -7660 -11000 -7640
rect -12460 -7760 -3580 -7700
rect -3520 -7760 44880 -7700
rect 44940 -7760 47240 -7700
rect -10700 -7820 -10600 -7800
rect -12460 -7880 -10680 -7820
rect -10620 -7880 7820 -7820
rect 7880 -7880 11580 -7820
rect 11640 -7880 29720 -7820
rect 29780 -7880 33480 -7820
rect 33540 -7880 47240 -7820
rect -10700 -7900 -10600 -7880
rect -12460 -8000 -3580 -7940
rect -3520 -8000 44880 -7940
rect 44940 -8000 47240 -7940
rect -10300 -8060 -10200 -8040
rect -12460 -8120 -10280 -8060
rect -10220 -8120 1940 -8060
rect 2000 -8120 3820 -8060
rect 3880 -8120 5520 -8060
rect 5580 -8120 13220 -8060
rect 13280 -8120 15100 -8060
rect 15160 -8120 16800 -8060
rect 16860 -8120 24500 -8060
rect 24560 -8120 26200 -8060
rect 26260 -8120 28080 -8060
rect 28140 -8120 35780 -8060
rect 35840 -8120 37480 -8060
rect 37540 -8120 39360 -8060
rect 39420 -8120 47240 -8060
rect -10300 -8140 -10200 -8120
rect -12460 -8240 -3580 -8180
rect -3520 -8240 44880 -8180
rect 44940 -8240 47240 -8180
rect -12460 -8320 47240 -8300
rect -12460 -8600 -9880 -8320
rect -9460 -8600 18860 -8320
rect 18920 -8600 20560 -8320
rect 20620 -8600 20740 -8320
rect 20800 -8600 22440 -8320
rect 22500 -8600 47240 -8320
rect -12460 -8620 47240 -8600
rect 48520 -8320 48840 -8300
rect 48520 -8600 48540 -8320
rect 48820 -8600 48840 -8320
rect 48520 -8620 48840 -8600
rect -12460 -8740 -3580 -8680
rect -3520 -8740 44880 -8680
rect 44940 -8740 47240 -8680
rect -9140 -8800 -9040 -8780
rect -12460 -8860 -9120 -8800
rect -9060 -8860 5700 -8800
rect 5760 -8860 7580 -8800
rect 7640 -8860 9280 -8800
rect 9340 -8860 9460 -8800
rect 9520 -8860 11340 -8800
rect 11400 -8860 13040 -8800
rect 13100 -8860 28260 -8800
rect 28320 -8860 29960 -8800
rect 30020 -8860 31840 -8800
rect 31900 -8860 32020 -8800
rect 32080 -8860 33720 -8800
rect 33780 -8860 35600 -8800
rect 35660 -8860 47240 -8800
rect -9140 -8880 -9040 -8860
rect -12460 -8980 -3580 -8920
rect -3520 -8980 44880 -8920
rect 44940 -8980 47240 -8920
rect -8740 -9040 -8640 -9020
rect -12460 -9100 -8720 -9040
rect -8660 -9100 3400 -9040
rect 3460 -9100 5280 -9040
rect 5340 -9100 5520 -9040
rect 5580 -9100 7160 -9040
rect 7220 -9100 9040 -9040
rect 9100 -9100 10920 -9040
rect 10980 -9100 11160 -9040
rect 11220 -9100 12800 -9040
rect 12860 -9100 14680 -9040
rect 14740 -9100 16560 -9040
rect 16620 -9100 16800 -9040
rect 16860 -9100 24500 -9040
rect 24560 -9100 24740 -9040
rect 24800 -9100 26620 -9040
rect 26680 -9100 28500 -9040
rect 28560 -9100 30140 -9040
rect 30200 -9100 30380 -9040
rect 30440 -9100 32260 -9040
rect 32320 -9100 34140 -9040
rect 34200 -9100 35780 -9040
rect 35840 -9100 36020 -9040
rect 36080 -9100 37900 -9040
rect 37960 -9100 47240 -9040
rect -8740 -9120 -8640 -9100
rect -12460 -9220 -3580 -9160
rect -3520 -9220 44880 -9160
rect 44940 -9220 47240 -9160
rect -8360 -9280 -8260 -9260
rect -12460 -9340 -8340 -9280
rect -8280 -9340 14920 -9280
rect 14980 -9340 16980 -9280
rect 17040 -9340 19100 -9280
rect 19160 -9340 22200 -9280
rect 22260 -9340 24320 -9280
rect 24380 -9340 26380 -9280
rect 26440 -9340 47240 -9280
rect -8360 -9360 -8260 -9340
rect -12460 -9460 -3580 -9400
rect -3520 -9460 44880 -9400
rect 44940 -9460 47240 -9400
rect -7960 -9520 -7860 -9500
rect -12460 -9580 -7940 -9520
rect -7880 -9580 9280 -9520
rect 9340 -9580 13040 -9520
rect 13100 -9580 18680 -9520
rect 18740 -9580 20320 -9520
rect 20380 -9580 20980 -9520
rect 21040 -9580 22620 -9520
rect 22680 -9580 28260 -9520
rect 28320 -9580 32020 -9520
rect 32080 -9580 47240 -9520
rect -7960 -9600 -7860 -9580
rect -12460 -9700 -3580 -9640
rect -3520 -9700 44880 -9640
rect 44940 -9700 47240 -9640
rect -7580 -9760 -7480 -9740
rect -12460 -9820 -7560 -9760
rect -7500 -9820 1520 -9760
rect 1580 -9820 1760 -9760
rect 1820 -9820 18440 -9760
rect 18500 -9820 22860 -9760
rect 22920 -9820 39540 -9760
rect 39600 -9820 39780 -9760
rect 39840 -9820 47240 -9760
rect -7580 -9840 -7480 -9820
rect -12460 -9940 -3580 -9880
rect -3520 -9940 44880 -9880
rect 44940 -9940 47240 -9880
rect -7180 -10000 -7080 -9980
rect -12460 -10060 -7160 -10000
rect -7100 -10060 -4120 -10000
rect -4060 -10060 -2240 -10000
rect -2180 -10060 -1820 -10000
rect -1760 -10060 -360 -10000
rect -300 -10060 60 -10000
rect 120 -10060 41240 -10000
rect 41300 -10060 41660 -10000
rect 41720 -10060 43120 -10000
rect 43180 -10060 43540 -10000
rect 43600 -10060 45420 -10000
rect 45480 -10060 47240 -10000
rect -7180 -10080 -7080 -10060
rect -12480 -10180 -12460 -10120
rect -12400 -10180 -12060 -10120
rect -12000 -10180 -11680 -10120
rect -11620 -10180 -11280 -10120
rect -11220 -10180 -10880 -10120
rect -10820 -10180 -10480 -10120
rect -10420 -10180 -10100 -10120
rect -10040 -10180 -9320 -10120
rect -9260 -10180 -8920 -10120
rect -8860 -10180 -8540 -10120
rect -8480 -10180 -8140 -10120
rect -8080 -10180 -7760 -10120
rect -7700 -10180 -7360 -10120
rect -7300 -10180 -6960 -10120
rect -6900 -10180 -3580 -10120
rect -3520 -10180 44880 -10120
rect 44940 -10180 47240 -10120
rect -6200 -12700 48840 -12680
rect -6200 -12980 -6180 -12700
rect -5900 -12980 -5580 -12700
rect -5520 -12980 -3880 -12700
rect -3820 -12980 -3700 -12700
rect -3640 -12980 -1820 -12700
rect -1760 -12980 1940 -12700
rect 2000 -12980 5700 -12700
rect 5760 -12980 9460 -12700
rect 9520 -12980 13220 -12700
rect 13280 -12980 18860 -12700
rect 18920 -12980 22440 -12700
rect 22500 -12980 28080 -12700
rect 28140 -12980 31840 -12700
rect 31900 -12980 35600 -12700
rect 35660 -12980 39360 -12700
rect 39420 -12980 43120 -12700
rect 43180 -12980 45000 -12700
rect 45060 -12980 45180 -12700
rect 45240 -12980 46880 -12700
rect 46940 -12980 47260 -12700
rect 47540 -12980 48840 -12700
rect -6200 -13000 48840 -12980
<< via2 >>
rect 18240 380 18340 480
rect -6820 -740 -6540 -460
rect 47900 -740 48180 -460
rect -12260 -6920 -12200 -6860
rect -11860 -7160 -11800 -7100
rect -11480 -7400 -11420 -7340
rect -11080 -7640 -11020 -7580
rect -10680 -7880 -10620 -7820
rect -10280 -8120 -10220 -8060
rect -9880 -8600 -9460 -8320
rect 48540 -8600 48820 -8320
rect -9120 -8860 -9060 -8800
rect -8720 -9100 -8660 -9040
rect -8340 -9340 -8280 -9280
rect -7940 -9580 -7880 -9520
rect -7560 -9820 -7500 -9760
rect -7160 -10060 -7100 -10000
rect -6180 -12980 -5900 -12700
rect 47260 -12980 47540 -12700
<< metal3 >>
rect 18230 480 18350 485
rect 18230 380 18240 480
rect 18340 380 18350 480
rect 18230 375 18350 380
rect -12460 -13000 -12400 -440
rect -12260 -6840 -12200 -380
rect -12280 -6860 -12180 -6840
rect -12280 -6920 -12260 -6860
rect -12200 -6920 -12180 -6860
rect -12280 -6940 -12180 -6920
rect -12260 -13000 -12200 -6940
rect -12060 -13000 -12000 -440
rect -11860 -7080 -11800 -380
rect -11880 -7100 -11780 -7080
rect -11880 -7160 -11860 -7100
rect -11800 -7160 -11780 -7100
rect -11880 -7180 -11780 -7160
rect -11860 -13000 -11800 -7180
rect -11680 -13000 -11620 -440
rect -11480 -7320 -11420 -380
rect -11500 -7340 -11400 -7320
rect -11500 -7400 -11480 -7340
rect -11420 -7400 -11400 -7340
rect -11500 -7420 -11400 -7400
rect -11480 -13000 -11420 -7420
rect -11280 -13000 -11220 -440
rect -11080 -7560 -11020 -380
rect -11100 -7580 -11000 -7560
rect -11100 -7640 -11080 -7580
rect -11020 -7640 -11000 -7580
rect -11100 -7660 -11000 -7640
rect -11080 -13000 -11020 -7660
rect -10880 -13000 -10820 -440
rect -10680 -7800 -10620 -380
rect -10700 -7820 -10600 -7800
rect -10700 -7880 -10680 -7820
rect -10620 -7880 -10600 -7820
rect -10700 -7900 -10600 -7880
rect -10680 -13000 -10620 -7900
rect -10480 -13000 -10420 -440
rect -10280 -8040 -10220 -380
rect -10300 -8060 -10200 -8040
rect -10300 -8120 -10280 -8060
rect -10220 -8120 -10200 -8060
rect -10300 -8140 -10200 -8120
rect -10280 -13000 -10220 -8140
rect -10100 -13000 -10040 -440
rect -9900 -8320 -9440 -380
rect -9900 -8600 -9880 -8320
rect -9460 -8600 -9440 -8320
rect -9900 -13000 -9440 -8600
rect -9320 -13000 -9260 -440
rect -9120 -8780 -9060 -380
rect -9140 -8800 -9040 -8780
rect -9140 -8860 -9120 -8800
rect -9060 -8860 -9040 -8800
rect -9140 -8880 -9040 -8860
rect -9120 -13000 -9060 -8880
rect -8920 -13000 -8860 -440
rect -8720 -9020 -8660 -380
rect -8740 -9040 -8640 -9020
rect -8740 -9100 -8720 -9040
rect -8660 -9100 -8640 -9040
rect -8740 -9120 -8640 -9100
rect -8720 -13000 -8660 -9120
rect -8540 -13000 -8480 -440
rect -8340 -9260 -8280 -380
rect -8360 -9280 -8260 -9260
rect -8360 -9340 -8340 -9280
rect -8280 -9340 -8260 -9280
rect -8360 -9360 -8260 -9340
rect -8340 -13000 -8280 -9360
rect -8140 -13000 -8080 -440
rect -7940 -9500 -7880 -380
rect -7960 -9520 -7860 -9500
rect -7960 -9580 -7940 -9520
rect -7880 -9580 -7860 -9520
rect -7960 -9600 -7860 -9580
rect -7940 -13000 -7880 -9600
rect -7760 -13000 -7700 -440
rect -7560 -9740 -7500 -380
rect -7580 -9760 -7480 -9740
rect -7580 -9820 -7560 -9760
rect -7500 -9820 -7480 -9760
rect -7580 -9840 -7480 -9820
rect -7560 -13000 -7500 -9840
rect -7360 -13000 -7300 -440
rect -7160 -9980 -7100 -380
rect -7180 -10000 -7080 -9980
rect -7180 -10060 -7160 -10000
rect -7100 -10060 -7080 -10000
rect -7180 -10080 -7080 -10060
rect -7160 -13000 -7100 -10080
rect -6960 -13000 -6900 -440
rect -6840 -460 -6520 -440
rect -6840 -740 -6820 -460
rect -6540 -740 -6520 -460
rect -6840 -13000 -6520 -740
rect -6200 -12700 -5880 -440
rect -6200 -12980 -6180 -12700
rect -5900 -12980 -5880 -12700
rect -6200 -13000 -5880 -12980
rect 47240 -12700 47560 -380
rect 47240 -12980 47260 -12700
rect 47540 -12980 47560 -12700
rect 47240 -13000 47560 -12980
rect 47880 -460 48200 -380
rect 47880 -740 47900 -460
rect 48180 -740 48200 -460
rect 47880 -13000 48200 -740
rect 48520 -6880 48840 -380
rect 48520 -7140 48540 -6880
rect 48820 -7140 48840 -6880
rect 48520 -7360 48840 -7140
rect 48520 -7620 48540 -7360
rect 48820 -7620 48840 -7360
rect 48520 -7840 48840 -7620
rect 48520 -8100 48540 -7840
rect 48820 -8100 48840 -7840
rect 48520 -8320 48840 -8100
rect 48520 -8600 48540 -8320
rect 48820 -8600 48840 -8320
rect 48520 -8820 48840 -8600
rect 48520 -9080 48540 -8820
rect 48820 -9080 48840 -8820
rect 48520 -9300 48840 -9080
rect 48520 -9560 48540 -9300
rect 48820 -9560 48840 -9300
rect 48520 -9780 48840 -9560
rect 48520 -10040 48540 -9780
rect 48820 -10040 48840 -9780
rect 48520 -13000 48840 -10040
<< via3 >>
rect 48540 -7140 48820 -6880
rect 48540 -7620 48820 -7360
rect 48540 -8100 48820 -7840
rect 48540 -8600 48820 -8320
rect 48540 -9080 48820 -8820
rect 48540 -9560 48820 -9300
rect 48540 -10040 48820 -9780
<< metal4 >>
rect -6960 -6880 48840 -6860
rect -6960 -7140 48540 -6880
rect 48820 -7140 48840 -6880
rect -6960 -7160 48840 -7140
rect -6960 -7360 48840 -7340
rect -6960 -7620 48540 -7360
rect 48820 -7620 48840 -7360
rect -6960 -7640 48840 -7620
rect -6960 -7840 48840 -7820
rect -6960 -8100 48540 -7840
rect 48820 -8100 48840 -7840
rect -6960 -8120 48840 -8100
rect -6960 -8320 48840 -8300
rect -6960 -8600 48540 -8320
rect 48820 -8600 48840 -8320
rect -6960 -8620 48840 -8600
rect -6960 -8820 48840 -8800
rect -6960 -9080 48540 -8820
rect 48820 -9080 48840 -8820
rect -6960 -9100 48840 -9080
rect -6960 -9300 48840 -9280
rect -6960 -9560 48540 -9300
rect 48820 -9560 48840 -9300
rect -6960 -9580 48840 -9560
rect -6960 -9780 48840 -9760
rect -6960 -10040 48540 -9780
rect 48820 -10040 48840 -9780
rect -6960 -10060 48840 -10040
<< metal5 >>
rect -12260 -13000 -11800 -440
rect -11480 -13000 -11020 -440
rect -10680 -13000 -10220 -440
rect -9900 -13000 -9440 -440
rect -9120 -13000 -8660 -440
rect -8340 -13000 -7880 -440
rect -7560 -13000 -7100 -440
use n8_1  n8_1_8
timestamp 1634429522
transform 1 0 -5640 0 1 -12660
box 0 0 1880 2460
use n1_8  na4_1
timestamp 1634337365
transform 1 0 -3760 0 1 -12660
box 0 0 1880 2460
use p1_8  pa1_1
timestamp 1634440922
transform 1 0 -3760 0 1 -6720
box 0 0 1880 5940
use p8_1  p8_1_7
timestamp 1634440961
transform 1 0 -5640 0 1 -6720
box 0 0 1880 5940
use n1_8  nb4_1
timestamp 1634337365
transform 1 0 -1880 0 1 -12660
box 0 0 1880 2460
use p8_1  pa2_1
timestamp 1634440961
transform 1 0 -1880 0 1 -6720
box 0 0 1880 5940
use n8_1  nb3_1
timestamp 1634429522
transform 1 0 0 0 1 -12660
box 0 0 1880 2460
use p1_8  pb1_1
timestamp 1634440922
transform 1 0 0 0 1 -6720
box 0 0 1880 5940
use n1_8  ne4_1
timestamp 1634337365
transform 1 0 1880 0 1 -12660
box 0 0 1880 2460
use p1_8  pc1_1
timestamp 1634440922
transform 1 0 1880 0 1 -6720
box 0 0 1880 5940
use n8_1  ne3_1
timestamp 1634429522
transform 1 0 3760 0 1 -12660
box 0 0 1880 2460
use p8_1  pc2_1
timestamp 1634440961
transform 1 0 3760 0 1 -6720
box 0 0 1880 5940
use n1_8  nf4_1
timestamp 1634337365
transform 1 0 5640 0 1 -12660
box 0 0 1880 2460
use p1_8  pd1_1
timestamp 1634440922
transform 1 0 5640 0 1 -6720
box 0 0 1880 5940
use n8_1  nf3_1
timestamp 1634429522
transform 1 0 7520 0 1 -12660
box 0 0 1880 2460
use p8_1  pd2_1
timestamp 1634440961
transform 1 0 7520 0 1 -6720
box 0 0 1880 5940
use n1_8  nf4_2
timestamp 1634337365
transform 1 0 9400 0 1 -12660
box 0 0 1880 2460
use p1_8  pe1_1
timestamp 1634440922
transform 1 0 9400 0 1 -6720
box 0 0 1880 5940
use n8_1  nf3_2
timestamp 1634429522
transform 1 0 11280 0 1 -12660
box 0 0 1880 2460
use p8_1  pd2_2
timestamp 1634440961
transform 1 0 11280 0 1 -6720
box 0 0 1880 5940
use n1_8  ne4_2
timestamp 1634337365
transform 1 0 13160 0 1 -12660
box 0 0 1880 2460
use p1_8  pf1_1
timestamp 1634440922
transform 1 0 13160 0 1 -6720
box 0 0 1880 5940
use n8_1  ne3_2
timestamp 1634429522
transform 1 0 15040 0 1 -12660
box 0 0 1880 2460
use p8_1  pc2_2
timestamp 1634440961
transform 1 0 15040 0 1 -6720
box 0 0 1880 5940
use n8_1  nf2_1
timestamp 1634429522
transform 1 0 16920 0 1 -12660
box 0 0 1880 2460
use p8_1  pf2_1
timestamp 1634440961
transform 1 0 16920 0 1 -6720
box 0 0 1880 5940
use n8_1  ng4_1
timestamp 1634429522
transform 1 0 18800 0 1 -12660
box 0 0 1880 2460
use p8_1  pg1_1
timestamp 1634440961
transform 1 0 18800 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_6
timestamp 1634429522
transform -1 0 22560 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_6
timestamp 1634440961
transform -1 0 22560 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_5
timestamp 1634429522
transform -1 0 24440 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_5
timestamp 1634440961
transform -1 0 24440 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_4
timestamp 1634429522
transform -1 0 26320 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_4
timestamp 1634440961
transform -1 0 26320 0 1 -6720
box 0 0 1880 5940
use n1_8  n1_8_5
timestamp 1634337365
transform -1 0 28200 0 1 -12660
box 0 0 1880 2460
use p1_8  p1_8_5
timestamp 1634440922
transform -1 0 28200 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_3
timestamp 1634429522
transform -1 0 30080 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_3
timestamp 1634440961
transform -1 0 30080 0 1 -6720
box 0 0 1880 5940
use n1_8  n1_8_4
timestamp 1634337365
transform -1 0 31960 0 1 -12660
box 0 0 1880 2460
use p1_8  p1_8_4
timestamp 1634440922
transform -1 0 31960 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_2
timestamp 1634429522
transform -1 0 33840 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_2
timestamp 1634440961
transform -1 0 33840 0 1 -6720
box 0 0 1880 5940
use n1_8  n1_8_3
timestamp 1634337365
transform -1 0 35720 0 1 -12660
box 0 0 1880 2460
use p1_8  p1_8_3
timestamp 1634440922
transform -1 0 35720 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_1
timestamp 1634429522
transform -1 0 37600 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_1
timestamp 1634440961
transform -1 0 37600 0 1 -6720
box 0 0 1880 5940
use n1_8  n1_8_2
timestamp 1634337365
transform -1 0 39480 0 1 -12660
box 0 0 1880 2460
use p1_8  p1_8_2
timestamp 1634440922
transform -1 0 39480 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_0
timestamp 1634429522
transform -1 0 41360 0 1 -12660
box 0 0 1880 2460
use p1_8  p1_8_1
timestamp 1634440922
transform -1 0 41360 0 1 -6720
box 0 0 1880 5940
use n1_8  n1_8_0
timestamp 1634337365
transform -1 0 43240 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_0
timestamp 1634440961
transform -1 0 43240 0 1 -6720
box 0 0 1880 5940
use n1_8  n1_8_1
timestamp 1634337365
transform -1 0 45120 0 1 -12660
box 0 0 1880 2460
use p1_8  p1_8_0
timestamp 1634440922
transform -1 0 45120 0 1 -6720
box 0 0 1880 5940
use n8_1  n8_1_7
timestamp 1634429522
transform -1 0 47000 0 1 -12660
box 0 0 1880 2460
use p8_1  p8_1_8
timestamp 1634440961
transform -1 0 47000 0 1 -6720
box 0 0 1880 5940
<< labels >>
rlabel metal2 -12480 -7640 -12460 -7580 3 inm
rlabel metal3 -12260 -440 -12200 -380 1 p1
rlabel metal3 -11080 -440 -11020 -380 1 inm
port 1 n
rlabel metal3 -10680 -440 -10620 -380 1 inp
port 2 n
rlabel metal3 -10280 -440 -10220 -380 1 xm
rlabel metal3 -9900 -440 -9440 -380 1 out
port 3 n
rlabel metal3 -11860 -440 -11800 -380 1 ib
port 4 n
rlabel metal3 -11480 -440 -11420 -380 1 x
rlabel metal3 -9120 -440 -9060 -380 1 xp
rlabel metal3 -8720 -440 -8660 -380 1 a
rlabel metal3 -8340 -440 -8280 -380 1 b
rlabel metal3 -7940 -440 -7880 -380 1 c
rlabel metal3 -7560 -440 -7500 -380 1 n2
rlabel metal3 -7160 -440 -7100 -380 1 n1
rlabel metal3 47880 -440 48200 -380 1 vdda
port 5 n
rlabel metal3 48520 -440 48840 -380 1 gnda
port 6 n
rlabel metal3 47240 -440 47560 -380 1 vssa
port 7 n
<< end >>
