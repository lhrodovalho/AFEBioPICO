magic
tech sky130A
timestamp 1637789704
<< nwell >>
rect -180 -700 5180 -140
<< mvnmos >>
rect 0 -1440 200 -1340
rect 320 -1440 520 -1340
rect 640 -1440 840 -1340
rect 960 -1440 1160 -1340
rect 1280 -1440 1480 -1340
rect 1600 -1440 1800 -1340
rect 1920 -1440 2120 -1340
rect 2240 -1440 2440 -1340
rect 2560 -1440 2760 -1340
rect 2880 -1440 3080 -1340
rect 3200 -1440 3400 -1340
rect 3520 -1440 3720 -1340
rect 3840 -1440 4040 -1340
rect 4160 -1440 4360 -1340
rect 4480 -1440 4680 -1340
rect 4800 -1440 5000 -1340
<< mvpmos >>
rect 0 -540 200 -240
rect 320 -540 520 -240
rect 640 -540 840 -240
rect 960 -540 1160 -240
rect 1280 -540 1480 -240
rect 1600 -540 1800 -240
rect 1920 -540 2120 -240
rect 2240 -540 2440 -240
rect 2560 -540 2760 -240
rect 2880 -540 3080 -240
rect 3200 -540 3400 -240
rect 3520 -540 3720 -240
rect 3840 -540 4040 -240
rect 4160 -540 4360 -240
rect 4480 -540 4680 -240
rect 4800 -540 5000 -240
<< mvndiff >>
rect -80 -1350 0 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 0 -1350
rect -80 -1440 0 -1430
rect 200 -1350 320 -1340
rect 200 -1430 245 -1350
rect 275 -1430 320 -1350
rect 200 -1440 320 -1430
rect 520 -1350 640 -1340
rect 520 -1430 565 -1350
rect 595 -1430 640 -1350
rect 520 -1440 640 -1430
rect 840 -1350 960 -1340
rect 840 -1430 885 -1350
rect 915 -1430 960 -1350
rect 840 -1440 960 -1430
rect 1160 -1350 1280 -1340
rect 1160 -1430 1205 -1350
rect 1235 -1430 1280 -1350
rect 1160 -1440 1280 -1430
rect 1480 -1350 1600 -1340
rect 1480 -1430 1525 -1350
rect 1555 -1430 1600 -1350
rect 1480 -1440 1600 -1430
rect 1800 -1350 1920 -1340
rect 1800 -1430 1845 -1350
rect 1875 -1430 1920 -1350
rect 1800 -1440 1920 -1430
rect 2120 -1350 2240 -1340
rect 2120 -1430 2165 -1350
rect 2195 -1430 2240 -1350
rect 2120 -1440 2240 -1430
rect 2440 -1350 2560 -1340
rect 2440 -1430 2485 -1350
rect 2515 -1430 2560 -1350
rect 2440 -1440 2560 -1430
rect 2760 -1350 2880 -1340
rect 2760 -1430 2805 -1350
rect 2835 -1430 2880 -1350
rect 2760 -1440 2880 -1430
rect 3080 -1350 3200 -1340
rect 3080 -1430 3125 -1350
rect 3155 -1430 3200 -1350
rect 3080 -1440 3200 -1430
rect 3400 -1350 3520 -1340
rect 3400 -1430 3445 -1350
rect 3475 -1430 3520 -1350
rect 3400 -1440 3520 -1430
rect 3720 -1350 3840 -1340
rect 3720 -1430 3765 -1350
rect 3795 -1430 3840 -1350
rect 3720 -1440 3840 -1430
rect 4040 -1350 4160 -1340
rect 4040 -1430 4085 -1350
rect 4115 -1430 4160 -1350
rect 4040 -1440 4160 -1430
rect 4360 -1350 4480 -1340
rect 4360 -1430 4405 -1350
rect 4435 -1430 4480 -1350
rect 4360 -1440 4480 -1430
rect 4680 -1350 4800 -1340
rect 4680 -1430 4725 -1350
rect 4755 -1430 4800 -1350
rect 4680 -1440 4800 -1430
rect 5000 -1350 5080 -1340
rect 5000 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5000 -1440 5080 -1430
<< mvpdiff >>
rect -80 -250 0 -240
rect -80 -530 -75 -250
rect -45 -530 0 -250
rect -80 -540 0 -530
rect 200 -250 320 -240
rect 200 -530 245 -250
rect 275 -530 320 -250
rect 200 -540 320 -530
rect 520 -250 640 -240
rect 520 -530 565 -250
rect 595 -530 640 -250
rect 520 -540 640 -530
rect 840 -250 960 -240
rect 840 -530 885 -250
rect 915 -530 960 -250
rect 840 -540 960 -530
rect 1160 -250 1280 -240
rect 1160 -530 1205 -250
rect 1235 -530 1280 -250
rect 1160 -540 1280 -530
rect 1480 -250 1600 -240
rect 1480 -530 1525 -250
rect 1555 -530 1600 -250
rect 1480 -540 1600 -530
rect 1800 -250 1920 -240
rect 1800 -530 1845 -250
rect 1875 -530 1920 -250
rect 1800 -540 1920 -530
rect 2120 -250 2240 -240
rect 2120 -530 2165 -250
rect 2195 -530 2240 -250
rect 2120 -540 2240 -530
rect 2440 -250 2560 -240
rect 2440 -530 2485 -250
rect 2515 -530 2560 -250
rect 2440 -540 2560 -530
rect 2760 -250 2880 -240
rect 2760 -530 2805 -250
rect 2835 -530 2880 -250
rect 2760 -540 2880 -530
rect 3080 -250 3200 -240
rect 3080 -530 3125 -250
rect 3155 -530 3200 -250
rect 3080 -540 3200 -530
rect 3400 -250 3520 -240
rect 3400 -530 3445 -250
rect 3475 -530 3520 -250
rect 3400 -540 3520 -530
rect 3720 -250 3840 -240
rect 3720 -530 3765 -250
rect 3795 -530 3840 -250
rect 3720 -540 3840 -530
rect 4040 -250 4160 -240
rect 4040 -530 4085 -250
rect 4115 -530 4160 -250
rect 4040 -540 4160 -530
rect 4360 -250 4480 -240
rect 4360 -530 4405 -250
rect 4435 -530 4480 -250
rect 4360 -540 4480 -530
rect 4680 -250 4800 -240
rect 4680 -530 4725 -250
rect 4755 -530 4800 -250
rect 4680 -540 4800 -530
rect 5000 -250 5080 -240
rect 5000 -530 5045 -250
rect 5075 -530 5080 -250
rect 5000 -540 5080 -530
<< mvndiffc >>
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
<< mvpdiffc >>
rect -75 -530 -45 -250
rect 245 -530 275 -250
rect 565 -530 595 -250
rect 885 -530 915 -250
rect 1205 -530 1235 -250
rect 1525 -530 1555 -250
rect 1845 -530 1875 -250
rect 2165 -530 2195 -250
rect 2485 -530 2515 -250
rect 2805 -530 2835 -250
rect 3125 -530 3155 -250
rect 3445 -530 3475 -250
rect 3765 -530 3795 -250
rect 4085 -530 4115 -250
rect 4405 -530 4435 -250
rect 4725 -530 4755 -250
rect 5045 -530 5075 -250
<< psubdiff >>
rect -240 -120 -180 -80
rect 5180 -120 5240 -80
rect -240 -140 -200 -120
rect 5200 -140 5240 -120
rect -200 -760 -180 -720
rect 5180 -760 5200 -720
rect -200 -1240 -180 -1200
rect 5180 -1240 5200 -1200
rect -240 -1480 -200 -1460
rect 5200 -1480 5240 -1460
rect -240 -1520 -180 -1480
rect 5180 -1520 5240 -1480
<< nsubdiff >>
rect -160 -200 -100 -160
rect 5100 -200 5160 -160
rect -160 -220 -120 -200
rect 5120 -220 5160 -200
rect -160 -640 -120 -620
rect 5120 -640 5160 -620
rect -160 -680 -100 -640
rect 5100 -680 5160 -640
<< psubdiffcont >>
rect -180 -120 5180 -80
rect -240 -1460 -200 -140
rect -180 -760 5180 -720
rect -180 -1240 5180 -1200
rect 5200 -1460 5240 -140
rect -180 -1520 5180 -1480
<< nsubdiffcont >>
rect -100 -200 5100 -160
rect -160 -620 -120 -220
rect 5120 -620 5160 -220
rect -100 -680 5100 -640
<< poly >>
rect 0 -240 200 -220
rect 320 -240 520 -220
rect 640 -240 840 -220
rect 960 -240 1160 -220
rect 1280 -240 1480 -220
rect 1600 -240 1800 -220
rect 1920 -240 2120 -220
rect 2240 -240 2440 -220
rect 2560 -240 2760 -220
rect 2880 -240 3080 -220
rect 3200 -240 3400 -220
rect 3520 -240 3720 -220
rect 3840 -240 4040 -220
rect 4160 -240 4360 -220
rect 4480 -240 4680 -220
rect 4800 -240 5000 -220
rect 0 -565 200 -540
rect 0 -595 10 -565
rect 190 -595 200 -565
rect 0 -600 200 -595
rect 320 -565 520 -540
rect 320 -595 330 -565
rect 510 -595 520 -565
rect 320 -600 520 -595
rect 640 -565 840 -540
rect 640 -595 650 -565
rect 830 -595 840 -565
rect 640 -600 840 -595
rect 960 -565 1160 -540
rect 960 -595 970 -565
rect 1150 -595 1160 -565
rect 960 -600 1160 -595
rect 1280 -565 1480 -540
rect 1280 -595 1290 -565
rect 1470 -595 1480 -565
rect 1280 -600 1480 -595
rect 1600 -565 1800 -540
rect 1600 -595 1610 -565
rect 1790 -595 1800 -565
rect 1600 -600 1800 -595
rect 1920 -565 2120 -540
rect 1920 -595 1930 -565
rect 2110 -595 2120 -565
rect 1920 -600 2120 -595
rect 2240 -565 2440 -540
rect 2240 -595 2250 -565
rect 2430 -595 2440 -565
rect 2240 -600 2440 -595
rect 2560 -565 2760 -540
rect 2560 -595 2570 -565
rect 2750 -595 2760 -565
rect 2560 -600 2760 -595
rect 2880 -565 3080 -540
rect 2880 -595 2890 -565
rect 3070 -595 3080 -565
rect 2880 -600 3080 -595
rect 3200 -565 3400 -540
rect 3200 -595 3210 -565
rect 3390 -595 3400 -565
rect 3200 -600 3400 -595
rect 3520 -565 3720 -540
rect 3520 -595 3530 -565
rect 3710 -595 3720 -565
rect 3520 -600 3720 -595
rect 3840 -565 4040 -540
rect 3840 -595 3850 -565
rect 4030 -595 4040 -565
rect 3840 -600 4040 -595
rect 4160 -565 4360 -540
rect 4160 -595 4170 -565
rect 4350 -595 4360 -565
rect 4160 -600 4360 -595
rect 4480 -565 4680 -540
rect 4480 -595 4490 -565
rect 4670 -595 4680 -565
rect 4480 -600 4680 -595
rect 4800 -565 5000 -540
rect 4800 -595 4810 -565
rect 4990 -595 5000 -565
rect 4800 -600 5000 -595
rect 0 -1285 200 -1280
rect 0 -1315 10 -1285
rect 190 -1315 200 -1285
rect 0 -1340 200 -1315
rect 320 -1285 520 -1280
rect 320 -1315 330 -1285
rect 510 -1315 520 -1285
rect 320 -1340 520 -1315
rect 640 -1285 840 -1280
rect 640 -1315 650 -1285
rect 830 -1315 840 -1285
rect 640 -1340 840 -1315
rect 960 -1285 1160 -1280
rect 960 -1315 970 -1285
rect 1150 -1315 1160 -1285
rect 960 -1340 1160 -1315
rect 1280 -1285 1480 -1280
rect 1280 -1315 1290 -1285
rect 1470 -1315 1480 -1285
rect 1280 -1340 1480 -1315
rect 1600 -1285 1800 -1280
rect 1600 -1315 1610 -1285
rect 1790 -1315 1800 -1285
rect 1600 -1340 1800 -1315
rect 1920 -1285 2120 -1280
rect 1920 -1315 1930 -1285
rect 2110 -1315 2120 -1285
rect 1920 -1340 2120 -1315
rect 2240 -1285 2440 -1280
rect 2240 -1315 2250 -1285
rect 2430 -1315 2440 -1285
rect 2240 -1340 2440 -1315
rect 2560 -1285 2760 -1280
rect 2560 -1315 2570 -1285
rect 2750 -1315 2760 -1285
rect 2560 -1340 2760 -1315
rect 2880 -1285 3080 -1280
rect 2880 -1315 2890 -1285
rect 3070 -1315 3080 -1285
rect 2880 -1340 3080 -1315
rect 3200 -1285 3400 -1280
rect 3200 -1315 3210 -1285
rect 3390 -1315 3400 -1285
rect 3200 -1340 3400 -1315
rect 3520 -1285 3720 -1280
rect 3520 -1315 3530 -1285
rect 3710 -1315 3720 -1285
rect 3520 -1340 3720 -1315
rect 3840 -1285 4040 -1280
rect 3840 -1315 3850 -1285
rect 4030 -1315 4040 -1285
rect 3840 -1340 4040 -1315
rect 4160 -1285 4360 -1280
rect 4160 -1315 4170 -1285
rect 4350 -1315 4360 -1285
rect 4160 -1340 4360 -1315
rect 4480 -1285 4680 -1280
rect 4480 -1315 4490 -1285
rect 4670 -1315 4680 -1285
rect 4480 -1340 4680 -1315
rect 4800 -1285 5000 -1280
rect 4800 -1315 4810 -1285
rect 4990 -1315 5000 -1285
rect 4800 -1340 5000 -1315
rect 0 -1460 200 -1440
rect 320 -1460 520 -1440
rect 640 -1460 840 -1440
rect 960 -1460 1160 -1440
rect 1280 -1460 1480 -1440
rect 1600 -1460 1800 -1440
rect 1920 -1460 2120 -1440
rect 2240 -1460 2440 -1440
rect 2560 -1460 2760 -1440
rect 2880 -1460 3080 -1440
rect 3200 -1460 3400 -1440
rect 3520 -1460 3720 -1440
rect 3840 -1460 4040 -1440
rect 4160 -1460 4360 -1440
rect 4480 -1460 4680 -1440
rect 4800 -1460 5000 -1440
<< polycont >>
rect 10 -595 190 -565
rect 330 -595 510 -565
rect 650 -595 830 -565
rect 970 -595 1150 -565
rect 1290 -595 1470 -565
rect 1610 -595 1790 -565
rect 1930 -595 2110 -565
rect 2250 -595 2430 -565
rect 2570 -595 2750 -565
rect 2890 -595 3070 -565
rect 3210 -595 3390 -565
rect 3530 -595 3710 -565
rect 3850 -595 4030 -565
rect 4170 -595 4350 -565
rect 4490 -595 4670 -565
rect 4810 -595 4990 -565
rect 10 -1315 190 -1285
rect 330 -1315 510 -1285
rect 650 -1315 830 -1285
rect 970 -1315 1150 -1285
rect 1290 -1315 1470 -1285
rect 1610 -1315 1790 -1285
rect 1930 -1315 2110 -1285
rect 2250 -1315 2430 -1285
rect 2570 -1315 2750 -1285
rect 2890 -1315 3070 -1285
rect 3210 -1315 3390 -1285
rect 3530 -1315 3710 -1285
rect 3850 -1315 4030 -1285
rect 4170 -1315 4350 -1285
rect 4490 -1315 4670 -1285
rect 4810 -1315 4990 -1285
<< locali >>
rect -240 -120 -180 -80
rect 5180 -120 5240 -80
rect -240 -140 -200 -120
rect 5200 -140 5240 -120
rect -160 -200 -100 -160
rect 5100 -200 5160 -160
rect -160 -220 -120 -200
rect 5120 -220 5160 -200
rect -80 -250 -40 -240
rect -80 -530 -75 -250
rect -45 -530 -40 -250
rect -80 -540 -40 -530
rect 240 -250 280 -240
rect 240 -530 245 -250
rect 275 -530 280 -250
rect 240 -540 280 -530
rect 560 -250 600 -240
rect 560 -530 565 -250
rect 595 -530 600 -250
rect 560 -540 600 -530
rect 880 -250 920 -240
rect 880 -530 885 -250
rect 915 -530 920 -250
rect 880 -540 920 -530
rect 1200 -250 1240 -240
rect 1200 -530 1205 -250
rect 1235 -530 1240 -250
rect 1200 -540 1240 -530
rect 1520 -250 1560 -240
rect 1520 -530 1525 -250
rect 1555 -530 1560 -250
rect 1520 -540 1560 -530
rect 1840 -250 1880 -240
rect 1840 -530 1845 -250
rect 1875 -530 1880 -250
rect 1840 -540 1880 -530
rect 2160 -250 2200 -240
rect 2160 -530 2165 -250
rect 2195 -530 2200 -250
rect 2160 -540 2200 -530
rect 2480 -250 2520 -240
rect 2480 -530 2485 -250
rect 2515 -530 2520 -250
rect 2480 -540 2520 -530
rect 2800 -250 2840 -240
rect 2800 -530 2805 -250
rect 2835 -530 2840 -250
rect 2800 -540 2840 -530
rect 3120 -250 3160 -240
rect 3120 -530 3125 -250
rect 3155 -530 3160 -250
rect 3120 -540 3160 -530
rect 3440 -250 3480 -240
rect 3440 -530 3445 -250
rect 3475 -530 3480 -250
rect 3440 -540 3480 -530
rect 3760 -250 3800 -240
rect 3760 -530 3765 -250
rect 3795 -530 3800 -250
rect 3760 -540 3800 -530
rect 4080 -250 4120 -240
rect 4080 -530 4085 -250
rect 4115 -530 4120 -250
rect 4080 -540 4120 -530
rect 4400 -250 4440 -240
rect 4400 -530 4405 -250
rect 4435 -530 4440 -250
rect 4400 -540 4440 -530
rect 4720 -250 4760 -240
rect 4720 -530 4725 -250
rect 4755 -530 4760 -250
rect 4720 -540 4760 -530
rect 5040 -250 5080 -240
rect 5040 -530 5045 -250
rect 5075 -530 5080 -250
rect 5040 -540 5080 -530
rect 0 -565 200 -560
rect 0 -595 10 -565
rect 190 -595 200 -565
rect 0 -600 200 -595
rect 320 -565 520 -560
rect 320 -595 330 -565
rect 510 -595 520 -565
rect 320 -600 520 -595
rect 640 -565 840 -560
rect 640 -595 650 -565
rect 830 -595 840 -565
rect 640 -600 840 -595
rect 960 -565 1160 -560
rect 960 -595 970 -565
rect 1150 -595 1160 -565
rect 960 -600 1160 -595
rect 1280 -565 1480 -560
rect 1280 -595 1290 -565
rect 1470 -595 1480 -565
rect 1280 -600 1480 -595
rect 1600 -565 1800 -560
rect 1600 -595 1610 -565
rect 1790 -595 1800 -565
rect 1600 -600 1800 -595
rect 1920 -565 2120 -560
rect 1920 -595 1930 -565
rect 2110 -595 2120 -565
rect 1920 -600 2120 -595
rect 2240 -565 2440 -560
rect 2240 -595 2250 -565
rect 2430 -595 2440 -565
rect 2240 -600 2440 -595
rect 2560 -565 2760 -560
rect 2560 -595 2570 -565
rect 2750 -595 2760 -565
rect 2560 -600 2760 -595
rect 2880 -565 3080 -560
rect 2880 -595 2890 -565
rect 3070 -595 3080 -565
rect 2880 -600 3080 -595
rect 3200 -565 3400 -560
rect 3200 -595 3210 -565
rect 3390 -595 3400 -565
rect 3200 -600 3400 -595
rect 3520 -565 3720 -560
rect 3520 -595 3530 -565
rect 3710 -595 3720 -565
rect 3520 -600 3720 -595
rect 3840 -565 4040 -560
rect 3840 -595 3850 -565
rect 4030 -595 4040 -565
rect 3840 -600 4040 -595
rect 4160 -565 4360 -560
rect 4160 -595 4170 -565
rect 4350 -595 4360 -565
rect 4160 -600 4360 -595
rect 4480 -565 4680 -560
rect 4480 -595 4490 -565
rect 4670 -595 4680 -565
rect 4480 -600 4680 -595
rect 4800 -565 5000 -560
rect 4800 -595 4810 -565
rect 4990 -595 5000 -565
rect 4800 -600 5000 -595
rect -160 -640 -120 -620
rect 5120 -640 5160 -620
rect -160 -680 -100 -640
rect 5100 -680 5160 -640
rect -200 -760 -180 -720
rect 5180 -760 5200 -720
rect -160 -1200 -120 -760
rect 0 -1200 40 -760
rect 80 -1200 120 -760
rect 160 -1200 200 -760
rect 320 -1200 360 -760
rect 400 -1200 440 -760
rect 480 -1200 520 -760
rect 640 -1200 680 -760
rect 720 -1200 760 -760
rect 800 -1200 840 -760
rect 960 -1200 1000 -760
rect 1040 -1200 1080 -760
rect 1120 -1200 1160 -760
rect 1280 -1200 1320 -760
rect 1360 -1200 1400 -760
rect 1440 -1200 1480 -760
rect 1600 -1200 1640 -760
rect 1680 -1200 1720 -760
rect 1760 -1200 1800 -760
rect 1920 -1200 1960 -760
rect 2000 -1200 2040 -760
rect 2080 -1200 2120 -760
rect 2240 -1200 2280 -760
rect 2320 -1200 2360 -760
rect 2400 -1200 2440 -760
rect 2560 -1200 2600 -760
rect 2640 -1200 2680 -760
rect 2720 -1200 2760 -760
rect 2880 -1200 2920 -760
rect 2960 -1200 3000 -760
rect 3040 -1200 3080 -760
rect 3200 -1200 3240 -760
rect 3280 -1200 3320 -760
rect 3360 -1200 3400 -760
rect 3520 -1200 3560 -760
rect 3600 -1200 3640 -760
rect 3680 -1200 3720 -760
rect 3840 -1200 3880 -760
rect 3920 -1200 3960 -760
rect 4000 -1200 4040 -760
rect 4160 -1200 4200 -760
rect 4240 -1200 4280 -760
rect 4320 -1200 4360 -760
rect 4480 -1200 4520 -760
rect 4560 -1200 4600 -760
rect 4640 -1200 4680 -760
rect 4800 -1200 4840 -760
rect 4880 -1200 4920 -760
rect 4960 -1200 5000 -760
rect 5120 -1200 5160 -760
rect -200 -1240 -180 -1200
rect 5180 -1240 5200 -1200
rect 0 -1285 200 -1280
rect 0 -1315 10 -1285
rect 190 -1315 200 -1285
rect 0 -1320 200 -1315
rect 320 -1285 520 -1280
rect 320 -1315 330 -1285
rect 510 -1315 520 -1285
rect 320 -1320 520 -1315
rect 640 -1285 840 -1280
rect 640 -1315 650 -1285
rect 830 -1315 840 -1285
rect 640 -1320 840 -1315
rect 960 -1285 1160 -1280
rect 960 -1315 970 -1285
rect 1150 -1315 1160 -1285
rect 960 -1320 1160 -1315
rect 1280 -1285 1480 -1280
rect 1280 -1315 1290 -1285
rect 1470 -1315 1480 -1285
rect 1280 -1320 1480 -1315
rect 1600 -1285 1800 -1280
rect 1600 -1315 1610 -1285
rect 1790 -1315 1800 -1285
rect 1600 -1320 1800 -1315
rect 1920 -1285 2120 -1280
rect 1920 -1315 1930 -1285
rect 2110 -1315 2120 -1285
rect 1920 -1320 2120 -1315
rect 2240 -1285 2440 -1280
rect 2240 -1315 2250 -1285
rect 2430 -1315 2440 -1285
rect 2240 -1320 2440 -1315
rect 2560 -1285 2760 -1280
rect 2560 -1315 2570 -1285
rect 2750 -1315 2760 -1285
rect 2560 -1320 2760 -1315
rect 2880 -1285 3080 -1280
rect 2880 -1315 2890 -1285
rect 3070 -1315 3080 -1285
rect 2880 -1320 3080 -1315
rect 3200 -1285 3400 -1280
rect 3200 -1315 3210 -1285
rect 3390 -1315 3400 -1285
rect 3200 -1320 3400 -1315
rect 3520 -1285 3720 -1280
rect 3520 -1315 3530 -1285
rect 3710 -1315 3720 -1285
rect 3520 -1320 3720 -1315
rect 3840 -1285 4040 -1280
rect 3840 -1315 3850 -1285
rect 4030 -1315 4040 -1285
rect 3840 -1320 4040 -1315
rect 4160 -1285 4360 -1280
rect 4160 -1315 4170 -1285
rect 4350 -1315 4360 -1285
rect 4160 -1320 4360 -1315
rect 4480 -1285 4680 -1280
rect 4480 -1315 4490 -1285
rect 4670 -1315 4680 -1285
rect 4480 -1320 4680 -1315
rect 4800 -1285 5000 -1280
rect 4800 -1315 4810 -1285
rect 4990 -1315 5000 -1285
rect 4800 -1320 5000 -1315
rect -80 -1350 -40 -1340
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1440 -40 -1430
rect 240 -1350 280 -1340
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1340
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -1340
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1340
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1440 1240 -1430
rect 1520 -1350 1560 -1340
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1340
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -1340
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1340
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1440 2520 -1430
rect 2800 -1350 2840 -1340
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1340
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -1340
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1340
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1440 3800 -1430
rect 4080 -1350 4120 -1340
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1340
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -1340
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1340
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1440 5080 -1430
rect -240 -1510 -235 -1460
rect -205 -1480 -200 -1460
rect 5200 -1480 5205 -1460
rect -205 -1510 -180 -1480
rect -240 -1520 -180 -1510
rect 5180 -1510 5205 -1480
rect 5235 -1510 5240 -1460
rect 5180 -1520 5240 -1510
<< viali >>
rect -70 -190 -50 -170
rect 570 -190 590 -170
rect 1210 -190 1230 -170
rect 1850 -190 1870 -170
rect 2490 -190 2510 -170
rect 3130 -190 3150 -170
rect 3770 -190 3790 -170
rect 4410 -190 4430 -170
rect 5050 -190 5070 -170
rect -75 -530 -45 -250
rect 245 -530 275 -250
rect 565 -530 595 -250
rect 885 -530 915 -250
rect 1205 -530 1235 -250
rect 1525 -530 1555 -250
rect 1845 -530 1875 -250
rect 2165 -530 2195 -250
rect 2485 -530 2515 -250
rect 2805 -530 2835 -250
rect 3125 -530 3155 -250
rect 3445 -530 3475 -250
rect 3765 -530 3795 -250
rect 4085 -530 4115 -250
rect 4405 -530 4435 -250
rect 4725 -530 4755 -250
rect 5045 -530 5075 -250
rect 10 -595 190 -565
rect 330 -595 510 -565
rect 650 -595 830 -565
rect 970 -595 1150 -565
rect 1290 -595 1470 -565
rect 1610 -595 1790 -565
rect 1930 -595 2110 -565
rect 2250 -595 2430 -565
rect 2570 -595 2750 -565
rect 2890 -595 3070 -565
rect 3210 -595 3390 -565
rect 3530 -595 3710 -565
rect 3850 -595 4030 -565
rect 4170 -595 4350 -565
rect 4490 -595 4670 -565
rect 4810 -595 4990 -565
rect 10 -1315 190 -1285
rect 330 -1315 510 -1285
rect 650 -1315 830 -1285
rect 970 -1315 1150 -1285
rect 1290 -1315 1470 -1285
rect 1610 -1315 1790 -1285
rect 1930 -1315 2110 -1285
rect 2250 -1315 2430 -1285
rect 2570 -1315 2750 -1285
rect 2890 -1315 3070 -1285
rect 3210 -1315 3390 -1285
rect 3530 -1315 3710 -1285
rect 3850 -1315 4030 -1285
rect 4170 -1315 4350 -1285
rect 4490 -1315 4670 -1285
rect 4810 -1315 4990 -1285
rect -235 -1460 -205 -1330
rect -75 -1430 -45 -1350
rect 245 -1430 275 -1350
rect 565 -1430 595 -1350
rect 885 -1430 915 -1350
rect 1205 -1430 1235 -1350
rect 1525 -1430 1555 -1350
rect 1845 -1430 1875 -1350
rect 2165 -1430 2195 -1350
rect 2485 -1430 2515 -1350
rect 2805 -1430 2835 -1350
rect 3125 -1430 3155 -1350
rect 3445 -1430 3475 -1350
rect 3765 -1430 3795 -1350
rect 4085 -1430 4115 -1350
rect 4405 -1430 4435 -1350
rect 4725 -1430 4755 -1350
rect 5045 -1430 5075 -1350
rect -235 -1510 -205 -1460
rect 5205 -1460 5235 -1330
rect 5205 -1510 5235 -1460
<< metal1 >>
rect -80 -165 -40 -160
rect -80 -195 -75 -165
rect -45 -195 -40 -165
rect -80 -200 -40 -195
rect 560 -165 600 -160
rect 560 -195 565 -165
rect 595 -195 600 -165
rect 560 -200 600 -195
rect 1200 -165 1240 -160
rect 1200 -195 1205 -165
rect 1235 -195 1240 -165
rect 1200 -200 1240 -195
rect 1840 -165 1880 -160
rect 1840 -195 1845 -165
rect 1875 -195 1880 -165
rect 1840 -200 1880 -195
rect 2480 -165 2520 -160
rect 2480 -195 2485 -165
rect 2515 -195 2520 -165
rect 2480 -200 2520 -195
rect 3120 -165 3160 -160
rect 3120 -195 3125 -165
rect 3155 -195 3160 -165
rect 3120 -200 3160 -195
rect 3760 -165 3800 -160
rect 3760 -195 3765 -165
rect 3795 -195 3800 -165
rect 3760 -200 3800 -195
rect 4400 -165 4440 -160
rect 4400 -195 4405 -165
rect 4435 -195 4440 -165
rect 4400 -200 4440 -195
rect 5040 -165 5080 -160
rect 5040 -195 5045 -165
rect 5075 -195 5080 -165
rect 5040 -200 5080 -195
rect -80 -250 -40 -240
rect -80 -530 -75 -250
rect -45 -530 -40 -250
rect -160 -805 -120 -800
rect -160 -835 -155 -805
rect -125 -835 -120 -805
rect -160 -965 -120 -835
rect -160 -995 -155 -965
rect -125 -995 -120 -965
rect -160 -1125 -120 -995
rect -160 -1155 -155 -1125
rect -125 -1155 -120 -1125
rect -160 -1160 -120 -1155
rect -80 -1045 -40 -530
rect 240 -250 280 -240
rect 240 -530 245 -250
rect 275 -530 280 -250
rect 0 -565 200 -560
rect 0 -595 10 -565
rect 190 -595 200 -565
rect 0 -600 200 -595
rect -80 -1075 -75 -1045
rect -45 -1075 -40 -1045
rect -240 -1330 -200 -1320
rect -240 -1510 -235 -1330
rect -205 -1510 -200 -1330
rect -80 -1350 -40 -1075
rect 0 -805 40 -800
rect 0 -835 5 -805
rect 35 -835 40 -805
rect 0 -965 40 -835
rect 0 -995 5 -965
rect 35 -995 40 -965
rect 0 -1125 40 -995
rect 0 -1155 5 -1125
rect 35 -1155 40 -1125
rect 0 -1160 40 -1155
rect 80 -805 120 -800
rect 80 -835 85 -805
rect 115 -835 120 -805
rect 80 -965 120 -835
rect 80 -995 85 -965
rect 115 -995 120 -965
rect 80 -1125 120 -995
rect 80 -1155 85 -1125
rect 115 -1155 120 -1125
rect 80 -1160 120 -1155
rect 160 -805 200 -800
rect 160 -835 165 -805
rect 195 -835 200 -805
rect 160 -965 200 -835
rect 160 -995 165 -965
rect 195 -995 200 -965
rect 160 -1125 200 -995
rect 160 -1155 165 -1125
rect 195 -1155 200 -1125
rect 160 -1160 200 -1155
rect 240 -885 280 -530
rect 560 -250 600 -240
rect 560 -530 565 -250
rect 595 -530 600 -250
rect 320 -565 520 -560
rect 320 -595 330 -565
rect 510 -595 520 -565
rect 320 -600 520 -595
rect 240 -915 245 -885
rect 275 -915 280 -885
rect 0 -1285 200 -1280
rect 0 -1315 10 -1285
rect 190 -1315 200 -1285
rect 0 -1320 200 -1315
rect -80 -1430 -75 -1350
rect -45 -1430 -40 -1350
rect -80 -1440 -40 -1430
rect 240 -1350 280 -915
rect 320 -805 360 -800
rect 320 -835 325 -805
rect 355 -835 360 -805
rect 320 -965 360 -835
rect 320 -995 325 -965
rect 355 -995 360 -965
rect 320 -1125 360 -995
rect 320 -1155 325 -1125
rect 355 -1155 360 -1125
rect 320 -1160 360 -1155
rect 400 -805 440 -800
rect 400 -835 405 -805
rect 435 -835 440 -805
rect 400 -965 440 -835
rect 400 -995 405 -965
rect 435 -995 440 -965
rect 400 -1125 440 -995
rect 400 -1155 405 -1125
rect 435 -1155 440 -1125
rect 400 -1160 440 -1155
rect 480 -805 520 -800
rect 480 -835 485 -805
rect 515 -835 520 -805
rect 480 -965 520 -835
rect 480 -995 485 -965
rect 515 -995 520 -965
rect 480 -1125 520 -995
rect 480 -1155 485 -1125
rect 515 -1155 520 -1125
rect 480 -1160 520 -1155
rect 560 -1045 600 -530
rect 880 -250 920 -240
rect 880 -530 885 -250
rect 915 -530 920 -250
rect 640 -565 840 -560
rect 640 -595 650 -565
rect 830 -595 840 -565
rect 640 -600 840 -595
rect 560 -1075 565 -1045
rect 595 -1075 600 -1045
rect 320 -1285 520 -1280
rect 320 -1315 330 -1285
rect 510 -1315 520 -1285
rect 320 -1320 520 -1315
rect 240 -1430 245 -1350
rect 275 -1430 280 -1350
rect 240 -1440 280 -1430
rect 560 -1350 600 -1075
rect 640 -805 680 -800
rect 640 -835 645 -805
rect 675 -835 680 -805
rect 640 -965 680 -835
rect 640 -995 645 -965
rect 675 -995 680 -965
rect 640 -1125 680 -995
rect 640 -1155 645 -1125
rect 675 -1155 680 -1125
rect 640 -1160 680 -1155
rect 720 -805 760 -800
rect 720 -835 725 -805
rect 755 -835 760 -805
rect 720 -965 760 -835
rect 720 -995 725 -965
rect 755 -995 760 -965
rect 720 -1125 760 -995
rect 720 -1155 725 -1125
rect 755 -1155 760 -1125
rect 720 -1160 760 -1155
rect 800 -805 840 -800
rect 800 -835 805 -805
rect 835 -835 840 -805
rect 800 -965 840 -835
rect 800 -995 805 -965
rect 835 -995 840 -965
rect 800 -1125 840 -995
rect 800 -1155 805 -1125
rect 835 -1155 840 -1125
rect 800 -1160 840 -1155
rect 880 -885 920 -530
rect 1200 -250 1240 -240
rect 1200 -530 1205 -250
rect 1235 -530 1240 -250
rect 960 -565 1160 -560
rect 960 -595 970 -565
rect 1150 -595 1160 -565
rect 960 -600 1160 -595
rect 880 -915 885 -885
rect 915 -915 920 -885
rect 640 -1285 840 -1280
rect 640 -1315 650 -1285
rect 830 -1315 840 -1285
rect 640 -1320 840 -1315
rect 560 -1430 565 -1350
rect 595 -1430 600 -1350
rect 560 -1440 600 -1430
rect 880 -1350 920 -915
rect 960 -805 1000 -800
rect 960 -835 965 -805
rect 995 -835 1000 -805
rect 960 -965 1000 -835
rect 960 -995 965 -965
rect 995 -995 1000 -965
rect 960 -1125 1000 -995
rect 960 -1155 965 -1125
rect 995 -1155 1000 -1125
rect 960 -1160 1000 -1155
rect 1040 -805 1080 -800
rect 1040 -835 1045 -805
rect 1075 -835 1080 -805
rect 1040 -965 1080 -835
rect 1040 -995 1045 -965
rect 1075 -995 1080 -965
rect 1040 -1125 1080 -995
rect 1040 -1155 1045 -1125
rect 1075 -1155 1080 -1125
rect 1040 -1160 1080 -1155
rect 1120 -805 1160 -800
rect 1120 -835 1125 -805
rect 1155 -835 1160 -805
rect 1120 -965 1160 -835
rect 1120 -995 1125 -965
rect 1155 -995 1160 -965
rect 1120 -1125 1160 -995
rect 1120 -1155 1125 -1125
rect 1155 -1155 1160 -1125
rect 1120 -1160 1160 -1155
rect 1200 -1045 1240 -530
rect 1520 -250 1560 -240
rect 1520 -530 1525 -250
rect 1555 -530 1560 -250
rect 1280 -565 1480 -560
rect 1280 -595 1290 -565
rect 1470 -595 1480 -565
rect 1280 -600 1480 -595
rect 1200 -1075 1205 -1045
rect 1235 -1075 1240 -1045
rect 960 -1285 1160 -1280
rect 960 -1315 970 -1285
rect 1150 -1315 1160 -1285
rect 960 -1320 1160 -1315
rect 880 -1430 885 -1350
rect 915 -1430 920 -1350
rect 880 -1440 920 -1430
rect 1200 -1350 1240 -1075
rect 1280 -805 1320 -800
rect 1280 -835 1285 -805
rect 1315 -835 1320 -805
rect 1280 -965 1320 -835
rect 1280 -995 1285 -965
rect 1315 -995 1320 -965
rect 1280 -1125 1320 -995
rect 1280 -1155 1285 -1125
rect 1315 -1155 1320 -1125
rect 1280 -1160 1320 -1155
rect 1360 -805 1400 -800
rect 1360 -835 1365 -805
rect 1395 -835 1400 -805
rect 1360 -965 1400 -835
rect 1360 -995 1365 -965
rect 1395 -995 1400 -965
rect 1360 -1125 1400 -995
rect 1360 -1155 1365 -1125
rect 1395 -1155 1400 -1125
rect 1360 -1160 1400 -1155
rect 1440 -805 1480 -800
rect 1440 -835 1445 -805
rect 1475 -835 1480 -805
rect 1440 -965 1480 -835
rect 1440 -995 1445 -965
rect 1475 -995 1480 -965
rect 1440 -1125 1480 -995
rect 1440 -1155 1445 -1125
rect 1475 -1155 1480 -1125
rect 1440 -1160 1480 -1155
rect 1520 -885 1560 -530
rect 1840 -250 1880 -240
rect 1840 -530 1845 -250
rect 1875 -530 1880 -250
rect 1600 -565 1800 -560
rect 1600 -595 1610 -565
rect 1790 -595 1800 -565
rect 1600 -600 1800 -595
rect 1520 -915 1525 -885
rect 1555 -915 1560 -885
rect 1280 -1285 1480 -1280
rect 1280 -1315 1290 -1285
rect 1470 -1315 1480 -1285
rect 1280 -1320 1480 -1315
rect 1200 -1430 1205 -1350
rect 1235 -1430 1240 -1350
rect 1200 -1440 1240 -1430
rect 1520 -1350 1560 -915
rect 1600 -805 1640 -800
rect 1600 -835 1605 -805
rect 1635 -835 1640 -805
rect 1600 -965 1640 -835
rect 1600 -995 1605 -965
rect 1635 -995 1640 -965
rect 1600 -1125 1640 -995
rect 1600 -1155 1605 -1125
rect 1635 -1155 1640 -1125
rect 1600 -1160 1640 -1155
rect 1680 -805 1720 -800
rect 1680 -835 1685 -805
rect 1715 -835 1720 -805
rect 1680 -965 1720 -835
rect 1680 -995 1685 -965
rect 1715 -995 1720 -965
rect 1680 -1125 1720 -995
rect 1680 -1155 1685 -1125
rect 1715 -1155 1720 -1125
rect 1680 -1160 1720 -1155
rect 1760 -805 1800 -800
rect 1760 -835 1765 -805
rect 1795 -835 1800 -805
rect 1760 -965 1800 -835
rect 1760 -995 1765 -965
rect 1795 -995 1800 -965
rect 1760 -1125 1800 -995
rect 1760 -1155 1765 -1125
rect 1795 -1155 1800 -1125
rect 1760 -1160 1800 -1155
rect 1840 -1045 1880 -530
rect 2160 -250 2200 -240
rect 2160 -530 2165 -250
rect 2195 -530 2200 -250
rect 1920 -565 2120 -560
rect 1920 -595 1930 -565
rect 2110 -595 2120 -565
rect 1920 -600 2120 -595
rect 1840 -1075 1845 -1045
rect 1875 -1075 1880 -1045
rect 1600 -1285 1800 -1280
rect 1600 -1315 1610 -1285
rect 1790 -1315 1800 -1285
rect 1600 -1320 1800 -1315
rect 1520 -1430 1525 -1350
rect 1555 -1430 1560 -1350
rect 1520 -1440 1560 -1430
rect 1840 -1350 1880 -1075
rect 1920 -805 1960 -800
rect 1920 -835 1925 -805
rect 1955 -835 1960 -805
rect 1920 -965 1960 -835
rect 1920 -995 1925 -965
rect 1955 -995 1960 -965
rect 1920 -1125 1960 -995
rect 1920 -1155 1925 -1125
rect 1955 -1155 1960 -1125
rect 1920 -1160 1960 -1155
rect 2000 -805 2040 -800
rect 2000 -835 2005 -805
rect 2035 -835 2040 -805
rect 2000 -965 2040 -835
rect 2000 -995 2005 -965
rect 2035 -995 2040 -965
rect 2000 -1125 2040 -995
rect 2000 -1155 2005 -1125
rect 2035 -1155 2040 -1125
rect 2000 -1160 2040 -1155
rect 2080 -805 2120 -800
rect 2080 -835 2085 -805
rect 2115 -835 2120 -805
rect 2080 -965 2120 -835
rect 2080 -995 2085 -965
rect 2115 -995 2120 -965
rect 2080 -1125 2120 -995
rect 2080 -1155 2085 -1125
rect 2115 -1155 2120 -1125
rect 2080 -1160 2120 -1155
rect 2160 -885 2200 -530
rect 2480 -250 2520 -240
rect 2480 -530 2485 -250
rect 2515 -530 2520 -250
rect 2240 -565 2440 -560
rect 2240 -595 2250 -565
rect 2430 -595 2440 -565
rect 2240 -600 2440 -595
rect 2160 -915 2165 -885
rect 2195 -915 2200 -885
rect 1920 -1285 2120 -1280
rect 1920 -1315 1930 -1285
rect 2110 -1315 2120 -1285
rect 1920 -1320 2120 -1315
rect 1840 -1430 1845 -1350
rect 1875 -1430 1880 -1350
rect 1840 -1440 1880 -1430
rect 2160 -1350 2200 -915
rect 2240 -805 2280 -800
rect 2240 -835 2245 -805
rect 2275 -835 2280 -805
rect 2240 -965 2280 -835
rect 2240 -995 2245 -965
rect 2275 -995 2280 -965
rect 2240 -1125 2280 -995
rect 2240 -1155 2245 -1125
rect 2275 -1155 2280 -1125
rect 2240 -1160 2280 -1155
rect 2320 -805 2360 -800
rect 2320 -835 2325 -805
rect 2355 -835 2360 -805
rect 2320 -965 2360 -835
rect 2320 -995 2325 -965
rect 2355 -995 2360 -965
rect 2320 -1125 2360 -995
rect 2320 -1155 2325 -1125
rect 2355 -1155 2360 -1125
rect 2320 -1160 2360 -1155
rect 2400 -805 2440 -800
rect 2400 -835 2405 -805
rect 2435 -835 2440 -805
rect 2400 -965 2440 -835
rect 2400 -995 2405 -965
rect 2435 -995 2440 -965
rect 2400 -1125 2440 -995
rect 2400 -1155 2405 -1125
rect 2435 -1155 2440 -1125
rect 2400 -1160 2440 -1155
rect 2480 -1045 2520 -530
rect 2800 -250 2840 -240
rect 2800 -530 2805 -250
rect 2835 -530 2840 -250
rect 2560 -565 2760 -560
rect 2560 -595 2570 -565
rect 2750 -595 2760 -565
rect 2560 -600 2760 -595
rect 2480 -1075 2485 -1045
rect 2515 -1075 2520 -1045
rect 2240 -1285 2440 -1280
rect 2240 -1315 2250 -1285
rect 2430 -1315 2440 -1285
rect 2240 -1320 2440 -1315
rect 2160 -1430 2165 -1350
rect 2195 -1430 2200 -1350
rect 2160 -1440 2200 -1430
rect 2480 -1350 2520 -1075
rect 2560 -805 2600 -800
rect 2560 -835 2565 -805
rect 2595 -835 2600 -805
rect 2560 -965 2600 -835
rect 2560 -995 2565 -965
rect 2595 -995 2600 -965
rect 2560 -1125 2600 -995
rect 2560 -1155 2565 -1125
rect 2595 -1155 2600 -1125
rect 2560 -1160 2600 -1155
rect 2640 -805 2680 -800
rect 2640 -835 2645 -805
rect 2675 -835 2680 -805
rect 2640 -965 2680 -835
rect 2640 -995 2645 -965
rect 2675 -995 2680 -965
rect 2640 -1125 2680 -995
rect 2640 -1155 2645 -1125
rect 2675 -1155 2680 -1125
rect 2640 -1160 2680 -1155
rect 2720 -805 2760 -800
rect 2720 -835 2725 -805
rect 2755 -835 2760 -805
rect 2720 -965 2760 -835
rect 2720 -995 2725 -965
rect 2755 -995 2760 -965
rect 2720 -1125 2760 -995
rect 2720 -1155 2725 -1125
rect 2755 -1155 2760 -1125
rect 2720 -1160 2760 -1155
rect 2800 -885 2840 -530
rect 3120 -250 3160 -240
rect 3120 -530 3125 -250
rect 3155 -530 3160 -250
rect 2880 -565 3080 -560
rect 2880 -595 2890 -565
rect 3070 -595 3080 -565
rect 2880 -600 3080 -595
rect 2800 -915 2805 -885
rect 2835 -915 2840 -885
rect 2560 -1285 2760 -1280
rect 2560 -1315 2570 -1285
rect 2750 -1315 2760 -1285
rect 2560 -1320 2760 -1315
rect 2480 -1430 2485 -1350
rect 2515 -1430 2520 -1350
rect 2480 -1440 2520 -1430
rect 2800 -1350 2840 -915
rect 2880 -805 2920 -800
rect 2880 -835 2885 -805
rect 2915 -835 2920 -805
rect 2880 -965 2920 -835
rect 2880 -995 2885 -965
rect 2915 -995 2920 -965
rect 2880 -1125 2920 -995
rect 2880 -1155 2885 -1125
rect 2915 -1155 2920 -1125
rect 2880 -1160 2920 -1155
rect 2960 -805 3000 -800
rect 2960 -835 2965 -805
rect 2995 -835 3000 -805
rect 2960 -965 3000 -835
rect 2960 -995 2965 -965
rect 2995 -995 3000 -965
rect 2960 -1125 3000 -995
rect 2960 -1155 2965 -1125
rect 2995 -1155 3000 -1125
rect 2960 -1160 3000 -1155
rect 3040 -805 3080 -800
rect 3040 -835 3045 -805
rect 3075 -835 3080 -805
rect 3040 -965 3080 -835
rect 3040 -995 3045 -965
rect 3075 -995 3080 -965
rect 3040 -1125 3080 -995
rect 3040 -1155 3045 -1125
rect 3075 -1155 3080 -1125
rect 3040 -1160 3080 -1155
rect 3120 -1045 3160 -530
rect 3440 -250 3480 -240
rect 3440 -530 3445 -250
rect 3475 -530 3480 -250
rect 3200 -565 3400 -560
rect 3200 -595 3210 -565
rect 3390 -595 3400 -565
rect 3200 -600 3400 -595
rect 3120 -1075 3125 -1045
rect 3155 -1075 3160 -1045
rect 2880 -1285 3080 -1280
rect 2880 -1315 2890 -1285
rect 3070 -1315 3080 -1285
rect 2880 -1320 3080 -1315
rect 2800 -1430 2805 -1350
rect 2835 -1430 2840 -1350
rect 2800 -1440 2840 -1430
rect 3120 -1350 3160 -1075
rect 3200 -805 3240 -800
rect 3200 -835 3205 -805
rect 3235 -835 3240 -805
rect 3200 -965 3240 -835
rect 3200 -995 3205 -965
rect 3235 -995 3240 -965
rect 3200 -1125 3240 -995
rect 3200 -1155 3205 -1125
rect 3235 -1155 3240 -1125
rect 3200 -1160 3240 -1155
rect 3280 -805 3320 -800
rect 3280 -835 3285 -805
rect 3315 -835 3320 -805
rect 3280 -965 3320 -835
rect 3280 -995 3285 -965
rect 3315 -995 3320 -965
rect 3280 -1125 3320 -995
rect 3280 -1155 3285 -1125
rect 3315 -1155 3320 -1125
rect 3280 -1160 3320 -1155
rect 3360 -805 3400 -800
rect 3360 -835 3365 -805
rect 3395 -835 3400 -805
rect 3360 -965 3400 -835
rect 3360 -995 3365 -965
rect 3395 -995 3400 -965
rect 3360 -1125 3400 -995
rect 3360 -1155 3365 -1125
rect 3395 -1155 3400 -1125
rect 3360 -1160 3400 -1155
rect 3440 -885 3480 -530
rect 3760 -250 3800 -240
rect 3760 -530 3765 -250
rect 3795 -530 3800 -250
rect 3520 -565 3720 -560
rect 3520 -595 3530 -565
rect 3710 -595 3720 -565
rect 3520 -600 3720 -595
rect 3440 -915 3445 -885
rect 3475 -915 3480 -885
rect 3200 -1285 3400 -1280
rect 3200 -1315 3210 -1285
rect 3390 -1315 3400 -1285
rect 3200 -1320 3400 -1315
rect 3120 -1430 3125 -1350
rect 3155 -1430 3160 -1350
rect 3120 -1440 3160 -1430
rect 3440 -1350 3480 -915
rect 3520 -805 3560 -800
rect 3520 -835 3525 -805
rect 3555 -835 3560 -805
rect 3520 -965 3560 -835
rect 3520 -995 3525 -965
rect 3555 -995 3560 -965
rect 3520 -1125 3560 -995
rect 3520 -1155 3525 -1125
rect 3555 -1155 3560 -1125
rect 3520 -1160 3560 -1155
rect 3600 -805 3640 -800
rect 3600 -835 3605 -805
rect 3635 -835 3640 -805
rect 3600 -965 3640 -835
rect 3600 -995 3605 -965
rect 3635 -995 3640 -965
rect 3600 -1125 3640 -995
rect 3600 -1155 3605 -1125
rect 3635 -1155 3640 -1125
rect 3600 -1160 3640 -1155
rect 3680 -805 3720 -800
rect 3680 -835 3685 -805
rect 3715 -835 3720 -805
rect 3680 -965 3720 -835
rect 3680 -995 3685 -965
rect 3715 -995 3720 -965
rect 3680 -1125 3720 -995
rect 3680 -1155 3685 -1125
rect 3715 -1155 3720 -1125
rect 3680 -1160 3720 -1155
rect 3760 -1045 3800 -530
rect 4080 -250 4120 -240
rect 4080 -530 4085 -250
rect 4115 -530 4120 -250
rect 3840 -565 4040 -560
rect 3840 -595 3850 -565
rect 4030 -595 4040 -565
rect 3840 -600 4040 -595
rect 3760 -1075 3765 -1045
rect 3795 -1075 3800 -1045
rect 3520 -1285 3720 -1280
rect 3520 -1315 3530 -1285
rect 3710 -1315 3720 -1285
rect 3520 -1320 3720 -1315
rect 3440 -1430 3445 -1350
rect 3475 -1430 3480 -1350
rect 3440 -1440 3480 -1430
rect 3760 -1350 3800 -1075
rect 3840 -805 3880 -800
rect 3840 -835 3845 -805
rect 3875 -835 3880 -805
rect 3840 -965 3880 -835
rect 3840 -995 3845 -965
rect 3875 -995 3880 -965
rect 3840 -1125 3880 -995
rect 3840 -1155 3845 -1125
rect 3875 -1155 3880 -1125
rect 3840 -1160 3880 -1155
rect 3920 -805 3960 -800
rect 3920 -835 3925 -805
rect 3955 -835 3960 -805
rect 3920 -965 3960 -835
rect 3920 -995 3925 -965
rect 3955 -995 3960 -965
rect 3920 -1125 3960 -995
rect 3920 -1155 3925 -1125
rect 3955 -1155 3960 -1125
rect 3920 -1160 3960 -1155
rect 4000 -805 4040 -800
rect 4000 -835 4005 -805
rect 4035 -835 4040 -805
rect 4000 -965 4040 -835
rect 4000 -995 4005 -965
rect 4035 -995 4040 -965
rect 4000 -1125 4040 -995
rect 4000 -1155 4005 -1125
rect 4035 -1155 4040 -1125
rect 4000 -1160 4040 -1155
rect 4080 -885 4120 -530
rect 4400 -250 4440 -240
rect 4400 -530 4405 -250
rect 4435 -530 4440 -250
rect 4160 -565 4360 -560
rect 4160 -595 4170 -565
rect 4350 -595 4360 -565
rect 4160 -600 4360 -595
rect 4080 -915 4085 -885
rect 4115 -915 4120 -885
rect 3840 -1285 4040 -1280
rect 3840 -1315 3850 -1285
rect 4030 -1315 4040 -1285
rect 3840 -1320 4040 -1315
rect 3760 -1430 3765 -1350
rect 3795 -1430 3800 -1350
rect 3760 -1440 3800 -1430
rect 4080 -1350 4120 -915
rect 4160 -805 4200 -800
rect 4160 -835 4165 -805
rect 4195 -835 4200 -805
rect 4160 -965 4200 -835
rect 4160 -995 4165 -965
rect 4195 -995 4200 -965
rect 4160 -1125 4200 -995
rect 4160 -1155 4165 -1125
rect 4195 -1155 4200 -1125
rect 4160 -1160 4200 -1155
rect 4240 -805 4280 -800
rect 4240 -835 4245 -805
rect 4275 -835 4280 -805
rect 4240 -965 4280 -835
rect 4240 -995 4245 -965
rect 4275 -995 4280 -965
rect 4240 -1125 4280 -995
rect 4240 -1155 4245 -1125
rect 4275 -1155 4280 -1125
rect 4240 -1160 4280 -1155
rect 4320 -805 4360 -800
rect 4320 -835 4325 -805
rect 4355 -835 4360 -805
rect 4320 -965 4360 -835
rect 4320 -995 4325 -965
rect 4355 -995 4360 -965
rect 4320 -1125 4360 -995
rect 4320 -1155 4325 -1125
rect 4355 -1155 4360 -1125
rect 4320 -1160 4360 -1155
rect 4400 -1045 4440 -530
rect 4720 -250 4760 -240
rect 4720 -530 4725 -250
rect 4755 -530 4760 -250
rect 4480 -565 4680 -560
rect 4480 -595 4490 -565
rect 4670 -595 4680 -565
rect 4480 -600 4680 -595
rect 4400 -1075 4405 -1045
rect 4435 -1075 4440 -1045
rect 4160 -1285 4360 -1280
rect 4160 -1315 4170 -1285
rect 4350 -1315 4360 -1285
rect 4160 -1320 4360 -1315
rect 4080 -1430 4085 -1350
rect 4115 -1430 4120 -1350
rect 4080 -1440 4120 -1430
rect 4400 -1350 4440 -1075
rect 4480 -805 4520 -800
rect 4480 -835 4485 -805
rect 4515 -835 4520 -805
rect 4480 -965 4520 -835
rect 4480 -995 4485 -965
rect 4515 -995 4520 -965
rect 4480 -1125 4520 -995
rect 4480 -1155 4485 -1125
rect 4515 -1155 4520 -1125
rect 4480 -1160 4520 -1155
rect 4560 -805 4600 -800
rect 4560 -835 4565 -805
rect 4595 -835 4600 -805
rect 4560 -965 4600 -835
rect 4560 -995 4565 -965
rect 4595 -995 4600 -965
rect 4560 -1125 4600 -995
rect 4560 -1155 4565 -1125
rect 4595 -1155 4600 -1125
rect 4560 -1160 4600 -1155
rect 4640 -805 4680 -800
rect 4640 -835 4645 -805
rect 4675 -835 4680 -805
rect 4640 -965 4680 -835
rect 4640 -995 4645 -965
rect 4675 -995 4680 -965
rect 4640 -1125 4680 -995
rect 4640 -1155 4645 -1125
rect 4675 -1155 4680 -1125
rect 4640 -1160 4680 -1155
rect 4720 -885 4760 -530
rect 5040 -250 5080 -240
rect 5040 -530 5045 -250
rect 5075 -530 5080 -250
rect 4800 -565 5000 -560
rect 4800 -595 4810 -565
rect 4990 -595 5000 -565
rect 4800 -600 5000 -595
rect 4720 -915 4725 -885
rect 4755 -915 4760 -885
rect 4480 -1285 4680 -1280
rect 4480 -1315 4490 -1285
rect 4670 -1315 4680 -1285
rect 4480 -1320 4680 -1315
rect 4400 -1430 4405 -1350
rect 4435 -1430 4440 -1350
rect 4400 -1440 4440 -1430
rect 4720 -1350 4760 -915
rect 4800 -805 4840 -800
rect 4800 -835 4805 -805
rect 4835 -835 4840 -805
rect 4800 -965 4840 -835
rect 4800 -995 4805 -965
rect 4835 -995 4840 -965
rect 4800 -1125 4840 -995
rect 4800 -1155 4805 -1125
rect 4835 -1155 4840 -1125
rect 4800 -1160 4840 -1155
rect 4880 -805 4920 -800
rect 4880 -835 4885 -805
rect 4915 -835 4920 -805
rect 4880 -965 4920 -835
rect 4880 -995 4885 -965
rect 4915 -995 4920 -965
rect 4880 -1125 4920 -995
rect 4880 -1155 4885 -1125
rect 4915 -1155 4920 -1125
rect 4880 -1160 4920 -1155
rect 4960 -805 5000 -800
rect 4960 -835 4965 -805
rect 4995 -835 5000 -805
rect 4960 -965 5000 -835
rect 4960 -995 4965 -965
rect 4995 -995 5000 -965
rect 4960 -1125 5000 -995
rect 4960 -1155 4965 -1125
rect 4995 -1155 5000 -1125
rect 4960 -1160 5000 -1155
rect 5040 -1045 5080 -530
rect 5040 -1075 5045 -1045
rect 5075 -1075 5080 -1045
rect 4800 -1285 5000 -1280
rect 4800 -1315 4810 -1285
rect 4990 -1315 5000 -1285
rect 4800 -1320 5000 -1315
rect 4720 -1430 4725 -1350
rect 4755 -1430 4760 -1350
rect 4720 -1440 4760 -1430
rect 5040 -1350 5080 -1075
rect 5120 -805 5160 -800
rect 5120 -835 5125 -805
rect 5155 -835 5160 -805
rect 5120 -965 5160 -835
rect 5120 -995 5125 -965
rect 5155 -995 5160 -965
rect 5120 -1125 5160 -995
rect 5120 -1155 5125 -1125
rect 5155 -1155 5160 -1125
rect 5120 -1160 5160 -1155
rect 5040 -1430 5045 -1350
rect 5075 -1430 5080 -1350
rect 5040 -1440 5080 -1430
rect 5200 -1330 5240 -1320
rect -240 -1520 -200 -1510
rect 5200 -1510 5205 -1330
rect 5235 -1510 5240 -1330
rect 5200 -1520 5240 -1510
<< via1 >>
rect -75 -170 -45 -165
rect -75 -190 -70 -170
rect -70 -190 -50 -170
rect -50 -190 -45 -170
rect -75 -195 -45 -190
rect 565 -170 595 -165
rect 565 -190 570 -170
rect 570 -190 590 -170
rect 590 -190 595 -170
rect 565 -195 595 -190
rect 1205 -170 1235 -165
rect 1205 -190 1210 -170
rect 1210 -190 1230 -170
rect 1230 -190 1235 -170
rect 1205 -195 1235 -190
rect 1845 -170 1875 -165
rect 1845 -190 1850 -170
rect 1850 -190 1870 -170
rect 1870 -190 1875 -170
rect 1845 -195 1875 -190
rect 2485 -170 2515 -165
rect 2485 -190 2490 -170
rect 2490 -190 2510 -170
rect 2510 -190 2515 -170
rect 2485 -195 2515 -190
rect 3125 -170 3155 -165
rect 3125 -190 3130 -170
rect 3130 -190 3150 -170
rect 3150 -190 3155 -170
rect 3125 -195 3155 -190
rect 3765 -170 3795 -165
rect 3765 -190 3770 -170
rect 3770 -190 3790 -170
rect 3790 -190 3795 -170
rect 3765 -195 3795 -190
rect 4405 -170 4435 -165
rect 4405 -190 4410 -170
rect 4410 -190 4430 -170
rect 4430 -190 4435 -170
rect 4405 -195 4435 -190
rect 5045 -170 5075 -165
rect 5045 -190 5050 -170
rect 5050 -190 5070 -170
rect 5070 -190 5075 -170
rect 5045 -195 5075 -190
rect -155 -835 -125 -805
rect -155 -995 -125 -965
rect -155 -1155 -125 -1125
rect 10 -595 190 -565
rect -75 -1075 -45 -1045
rect -235 -1510 -205 -1360
rect 5 -835 35 -805
rect 5 -995 35 -965
rect 5 -1155 35 -1125
rect 85 -835 115 -805
rect 85 -995 115 -965
rect 85 -1155 115 -1125
rect 165 -835 195 -805
rect 165 -995 195 -965
rect 165 -1155 195 -1125
rect 330 -595 510 -565
rect 245 -915 275 -885
rect 10 -1315 190 -1285
rect 325 -835 355 -805
rect 325 -995 355 -965
rect 325 -1155 355 -1125
rect 405 -835 435 -805
rect 405 -995 435 -965
rect 405 -1155 435 -1125
rect 485 -835 515 -805
rect 485 -995 515 -965
rect 485 -1155 515 -1125
rect 650 -595 830 -565
rect 565 -1075 595 -1045
rect 330 -1315 510 -1285
rect 645 -835 675 -805
rect 645 -995 675 -965
rect 645 -1155 675 -1125
rect 725 -835 755 -805
rect 725 -995 755 -965
rect 725 -1155 755 -1125
rect 805 -835 835 -805
rect 805 -995 835 -965
rect 805 -1155 835 -1125
rect 970 -595 1150 -565
rect 885 -915 915 -885
rect 650 -1315 830 -1285
rect 965 -835 995 -805
rect 965 -995 995 -965
rect 965 -1155 995 -1125
rect 1045 -835 1075 -805
rect 1045 -995 1075 -965
rect 1045 -1155 1075 -1125
rect 1125 -835 1155 -805
rect 1125 -995 1155 -965
rect 1125 -1155 1155 -1125
rect 1290 -595 1470 -565
rect 1205 -1075 1235 -1045
rect 970 -1315 1150 -1285
rect 1285 -835 1315 -805
rect 1285 -995 1315 -965
rect 1285 -1155 1315 -1125
rect 1365 -835 1395 -805
rect 1365 -995 1395 -965
rect 1365 -1155 1395 -1125
rect 1445 -835 1475 -805
rect 1445 -995 1475 -965
rect 1445 -1155 1475 -1125
rect 1610 -595 1790 -565
rect 1525 -915 1555 -885
rect 1290 -1315 1470 -1285
rect 1605 -835 1635 -805
rect 1605 -995 1635 -965
rect 1605 -1155 1635 -1125
rect 1685 -835 1715 -805
rect 1685 -995 1715 -965
rect 1685 -1155 1715 -1125
rect 1765 -835 1795 -805
rect 1765 -995 1795 -965
rect 1765 -1155 1795 -1125
rect 1930 -595 2110 -565
rect 1845 -1075 1875 -1045
rect 1610 -1315 1790 -1285
rect 1925 -835 1955 -805
rect 1925 -995 1955 -965
rect 1925 -1155 1955 -1125
rect 2005 -835 2035 -805
rect 2005 -995 2035 -965
rect 2005 -1155 2035 -1125
rect 2085 -835 2115 -805
rect 2085 -995 2115 -965
rect 2085 -1155 2115 -1125
rect 2250 -595 2430 -565
rect 2165 -915 2195 -885
rect 1930 -1315 2110 -1285
rect 2245 -835 2275 -805
rect 2245 -995 2275 -965
rect 2245 -1155 2275 -1125
rect 2325 -835 2355 -805
rect 2325 -995 2355 -965
rect 2325 -1155 2355 -1125
rect 2405 -835 2435 -805
rect 2405 -995 2435 -965
rect 2405 -1155 2435 -1125
rect 2570 -595 2750 -565
rect 2485 -1075 2515 -1045
rect 2250 -1315 2430 -1285
rect 2565 -835 2595 -805
rect 2565 -995 2595 -965
rect 2565 -1155 2595 -1125
rect 2645 -835 2675 -805
rect 2645 -995 2675 -965
rect 2645 -1155 2675 -1125
rect 2725 -835 2755 -805
rect 2725 -995 2755 -965
rect 2725 -1155 2755 -1125
rect 2890 -595 3070 -565
rect 2805 -915 2835 -885
rect 2570 -1315 2750 -1285
rect 2885 -835 2915 -805
rect 2885 -995 2915 -965
rect 2885 -1155 2915 -1125
rect 2965 -835 2995 -805
rect 2965 -995 2995 -965
rect 2965 -1155 2995 -1125
rect 3045 -835 3075 -805
rect 3045 -995 3075 -965
rect 3045 -1155 3075 -1125
rect 3210 -595 3390 -565
rect 3125 -1075 3155 -1045
rect 2890 -1315 3070 -1285
rect 3205 -835 3235 -805
rect 3205 -995 3235 -965
rect 3205 -1155 3235 -1125
rect 3285 -835 3315 -805
rect 3285 -995 3315 -965
rect 3285 -1155 3315 -1125
rect 3365 -835 3395 -805
rect 3365 -995 3395 -965
rect 3365 -1155 3395 -1125
rect 3530 -595 3710 -565
rect 3445 -915 3475 -885
rect 3210 -1315 3390 -1285
rect 3525 -835 3555 -805
rect 3525 -995 3555 -965
rect 3525 -1155 3555 -1125
rect 3605 -835 3635 -805
rect 3605 -995 3635 -965
rect 3605 -1155 3635 -1125
rect 3685 -835 3715 -805
rect 3685 -995 3715 -965
rect 3685 -1155 3715 -1125
rect 3850 -595 4030 -565
rect 3765 -1075 3795 -1045
rect 3530 -1315 3710 -1285
rect 3845 -835 3875 -805
rect 3845 -995 3875 -965
rect 3845 -1155 3875 -1125
rect 3925 -835 3955 -805
rect 3925 -995 3955 -965
rect 3925 -1155 3955 -1125
rect 4005 -835 4035 -805
rect 4005 -995 4035 -965
rect 4005 -1155 4035 -1125
rect 4170 -595 4350 -565
rect 4085 -915 4115 -885
rect 3850 -1315 4030 -1285
rect 4165 -835 4195 -805
rect 4165 -995 4195 -965
rect 4165 -1155 4195 -1125
rect 4245 -835 4275 -805
rect 4245 -995 4275 -965
rect 4245 -1155 4275 -1125
rect 4325 -835 4355 -805
rect 4325 -995 4355 -965
rect 4325 -1155 4355 -1125
rect 4490 -595 4670 -565
rect 4405 -1075 4435 -1045
rect 4170 -1315 4350 -1285
rect 4485 -835 4515 -805
rect 4485 -995 4515 -965
rect 4485 -1155 4515 -1125
rect 4565 -835 4595 -805
rect 4565 -995 4595 -965
rect 4565 -1155 4595 -1125
rect 4645 -835 4675 -805
rect 4645 -995 4675 -965
rect 4645 -1155 4675 -1125
rect 4810 -595 4990 -565
rect 4725 -915 4755 -885
rect 4490 -1315 4670 -1285
rect 4805 -835 4835 -805
rect 4805 -995 4835 -965
rect 4805 -1155 4835 -1125
rect 4885 -835 4915 -805
rect 4885 -995 4915 -965
rect 4885 -1155 4915 -1125
rect 4965 -835 4995 -805
rect 4965 -995 4995 -965
rect 4965 -1155 4995 -1125
rect 5045 -1075 5075 -1045
rect 4810 -1315 4990 -1285
rect 5125 -835 5155 -805
rect 5125 -995 5155 -965
rect 5125 -1155 5155 -1125
rect 5205 -1510 5235 -1360
<< metal2 >>
rect -240 -165 5240 -160
rect -240 -195 -75 -165
rect -45 -195 565 -165
rect 595 -195 1205 -165
rect 1235 -195 1845 -165
rect 1875 -195 2485 -165
rect 2515 -195 3125 -165
rect 3155 -195 3765 -165
rect 3795 -195 4405 -165
rect 4435 -195 5045 -165
rect 5075 -195 5240 -165
rect -240 -200 5240 -195
rect -240 -485 5240 -480
rect -240 -515 -235 -485
rect -205 -515 5205 -485
rect 5235 -515 5240 -485
rect -240 -520 5240 -515
rect -240 -565 5240 -560
rect -240 -595 10 -565
rect 190 -595 330 -565
rect 510 -595 650 -565
rect 830 -595 970 -565
rect 1150 -595 1290 -565
rect 1470 -595 1610 -565
rect 1790 -595 1930 -565
rect 2110 -595 2250 -565
rect 2430 -595 2570 -565
rect 2750 -595 2890 -565
rect 3070 -595 3210 -565
rect 3390 -595 3530 -565
rect 3710 -595 3850 -565
rect 4030 -595 4170 -565
rect 4350 -595 4490 -565
rect 4670 -595 4810 -565
rect 4990 -595 5240 -565
rect -240 -600 5240 -595
rect -240 -645 5240 -640
rect -240 -675 -235 -645
rect -205 -675 5205 -645
rect 5235 -675 5240 -645
rect -240 -680 5240 -675
rect -240 -725 5240 -720
rect -240 -755 -235 -725
rect -205 -755 5205 -725
rect 5235 -755 5240 -725
rect -240 -760 5240 -755
rect -240 -805 5240 -800
rect -240 -835 -155 -805
rect -125 -835 5 -805
rect 35 -835 85 -805
rect 115 -835 165 -805
rect 195 -835 325 -805
rect 355 -835 405 -805
rect 435 -835 485 -805
rect 515 -835 645 -805
rect 675 -835 725 -805
rect 755 -835 805 -805
rect 835 -835 965 -805
rect 995 -835 1045 -805
rect 1075 -835 1125 -805
rect 1155 -835 1285 -805
rect 1315 -835 1365 -805
rect 1395 -835 1445 -805
rect 1475 -835 1605 -805
rect 1635 -835 1685 -805
rect 1715 -835 1765 -805
rect 1795 -835 1925 -805
rect 1955 -835 2005 -805
rect 2035 -835 2085 -805
rect 2115 -835 2245 -805
rect 2275 -835 2325 -805
rect 2355 -835 2405 -805
rect 2435 -835 2565 -805
rect 2595 -835 2645 -805
rect 2675 -835 2725 -805
rect 2755 -835 2885 -805
rect 2915 -835 2965 -805
rect 2995 -835 3045 -805
rect 3075 -835 3205 -805
rect 3235 -835 3285 -805
rect 3315 -835 3365 -805
rect 3395 -835 3525 -805
rect 3555 -835 3605 -805
rect 3635 -835 3685 -805
rect 3715 -835 3845 -805
rect 3875 -835 3925 -805
rect 3955 -835 4005 -805
rect 4035 -835 4165 -805
rect 4195 -835 4245 -805
rect 4275 -835 4325 -805
rect 4355 -835 4485 -805
rect 4515 -835 4565 -805
rect 4595 -835 4645 -805
rect 4675 -835 4805 -805
rect 4835 -835 4885 -805
rect 4915 -835 4965 -805
rect 4995 -835 5125 -805
rect 5155 -835 5240 -805
rect -240 -840 5240 -835
rect -240 -885 5240 -880
rect -240 -915 245 -885
rect 275 -915 885 -885
rect 915 -915 1525 -885
rect 1555 -915 2165 -885
rect 2195 -915 2805 -885
rect 2835 -915 3445 -885
rect 3475 -915 4085 -885
rect 4115 -915 4725 -885
rect 4755 -915 5240 -885
rect -240 -920 5240 -915
rect -240 -965 5240 -960
rect -240 -995 -155 -965
rect -125 -995 5 -965
rect 35 -995 85 -965
rect 115 -995 165 -965
rect 195 -995 325 -965
rect 355 -995 405 -965
rect 435 -995 485 -965
rect 515 -995 645 -965
rect 675 -995 725 -965
rect 755 -995 805 -965
rect 835 -995 965 -965
rect 995 -995 1045 -965
rect 1075 -995 1125 -965
rect 1155 -995 1285 -965
rect 1315 -995 1365 -965
rect 1395 -995 1445 -965
rect 1475 -995 1605 -965
rect 1635 -995 1685 -965
rect 1715 -995 1765 -965
rect 1795 -995 1925 -965
rect 1955 -995 2005 -965
rect 2035 -995 2085 -965
rect 2115 -995 2245 -965
rect 2275 -995 2325 -965
rect 2355 -995 2405 -965
rect 2435 -995 2565 -965
rect 2595 -995 2645 -965
rect 2675 -995 2725 -965
rect 2755 -995 2885 -965
rect 2915 -995 2965 -965
rect 2995 -995 3045 -965
rect 3075 -995 3205 -965
rect 3235 -995 3285 -965
rect 3315 -995 3365 -965
rect 3395 -995 3525 -965
rect 3555 -995 3605 -965
rect 3635 -995 3685 -965
rect 3715 -995 3845 -965
rect 3875 -995 3925 -965
rect 3955 -995 4005 -965
rect 4035 -995 4165 -965
rect 4195 -995 4245 -965
rect 4275 -995 4325 -965
rect 4355 -995 4485 -965
rect 4515 -995 4565 -965
rect 4595 -995 4645 -965
rect 4675 -995 4805 -965
rect 4835 -995 4885 -965
rect 4915 -995 4965 -965
rect 4995 -995 5125 -965
rect 5155 -995 5240 -965
rect -240 -1000 5240 -995
rect -240 -1045 5240 -1040
rect -240 -1075 -75 -1045
rect -45 -1075 565 -1045
rect 595 -1075 1205 -1045
rect 1235 -1075 1845 -1045
rect 1875 -1075 2485 -1045
rect 2515 -1075 3125 -1045
rect 3155 -1075 3765 -1045
rect 3795 -1075 4405 -1045
rect 4435 -1075 5045 -1045
rect 5075 -1075 5240 -1045
rect -240 -1080 5240 -1075
rect -240 -1125 5240 -1120
rect -240 -1155 -155 -1125
rect -125 -1155 5 -1125
rect 35 -1155 85 -1125
rect 115 -1155 165 -1125
rect 195 -1155 325 -1125
rect 355 -1155 405 -1125
rect 435 -1155 485 -1125
rect 515 -1155 645 -1125
rect 675 -1155 725 -1125
rect 755 -1155 805 -1125
rect 835 -1155 965 -1125
rect 995 -1155 1045 -1125
rect 1075 -1155 1125 -1125
rect 1155 -1155 1285 -1125
rect 1315 -1155 1365 -1125
rect 1395 -1155 1445 -1125
rect 1475 -1155 1605 -1125
rect 1635 -1155 1685 -1125
rect 1715 -1155 1765 -1125
rect 1795 -1155 1925 -1125
rect 1955 -1155 2005 -1125
rect 2035 -1155 2085 -1125
rect 2115 -1155 2245 -1125
rect 2275 -1155 2325 -1125
rect 2355 -1155 2405 -1125
rect 2435 -1155 2565 -1125
rect 2595 -1155 2645 -1125
rect 2675 -1155 2725 -1125
rect 2755 -1155 2885 -1125
rect 2915 -1155 2965 -1125
rect 2995 -1155 3045 -1125
rect 3075 -1155 3205 -1125
rect 3235 -1155 3285 -1125
rect 3315 -1155 3365 -1125
rect 3395 -1155 3525 -1125
rect 3555 -1155 3605 -1125
rect 3635 -1155 3685 -1125
rect 3715 -1155 3845 -1125
rect 3875 -1155 3925 -1125
rect 3955 -1155 4005 -1125
rect 4035 -1155 4165 -1125
rect 4195 -1155 4245 -1125
rect 4275 -1155 4325 -1125
rect 4355 -1155 4485 -1125
rect 4515 -1155 4565 -1125
rect 4595 -1155 4645 -1125
rect 4675 -1155 4805 -1125
rect 4835 -1155 4885 -1125
rect 4915 -1155 4965 -1125
rect 4995 -1155 5125 -1125
rect 5155 -1155 5240 -1125
rect -240 -1160 5240 -1155
rect -240 -1205 5240 -1200
rect -240 -1235 -235 -1205
rect -205 -1235 5205 -1205
rect 5235 -1235 5240 -1205
rect -240 -1240 5240 -1235
rect -240 -1285 5240 -1280
rect -240 -1315 10 -1285
rect 190 -1315 330 -1285
rect 510 -1315 650 -1285
rect 830 -1315 970 -1285
rect 1150 -1315 1290 -1285
rect 1470 -1315 1610 -1285
rect 1790 -1315 1930 -1285
rect 2110 -1315 2250 -1285
rect 2430 -1315 2570 -1285
rect 2750 -1315 2890 -1285
rect 3070 -1315 3210 -1285
rect 3390 -1315 3530 -1285
rect 3710 -1315 3850 -1285
rect 4030 -1315 4170 -1285
rect 4350 -1315 4490 -1285
rect 4670 -1315 4810 -1285
rect 4990 -1315 5240 -1285
rect -240 -1320 5240 -1315
rect -240 -1510 -235 -1360
rect -205 -1400 5205 -1360
rect -205 -1510 -200 -1400
rect -240 -1520 -200 -1510
rect 5200 -1510 5205 -1400
rect 5235 -1510 5240 -1360
rect 5200 -1520 5240 -1510
<< via2 >>
rect -235 -515 -205 -485
rect 5205 -515 5235 -485
rect -235 -675 -205 -645
rect 5205 -675 5235 -645
rect -235 -755 -205 -725
rect 5205 -755 5235 -725
rect -155 -835 -125 -805
rect 5 -835 35 -805
rect 85 -835 115 -805
rect 165 -835 195 -805
rect 325 -835 355 -805
rect 405 -835 435 -805
rect 485 -835 515 -805
rect 645 -835 675 -805
rect 725 -835 755 -805
rect 805 -835 835 -805
rect 965 -835 995 -805
rect 1045 -835 1075 -805
rect 1125 -835 1155 -805
rect 1285 -835 1315 -805
rect 1365 -835 1395 -805
rect 1445 -835 1475 -805
rect 1605 -835 1635 -805
rect 1685 -835 1715 -805
rect 1765 -835 1795 -805
rect 1925 -835 1955 -805
rect 2005 -835 2035 -805
rect 2085 -835 2115 -805
rect 2245 -835 2275 -805
rect 2325 -835 2355 -805
rect 2405 -835 2435 -805
rect 2565 -835 2595 -805
rect 2645 -835 2675 -805
rect 2725 -835 2755 -805
rect 2885 -835 2915 -805
rect 2965 -835 2995 -805
rect 3045 -835 3075 -805
rect 3205 -835 3235 -805
rect 3285 -835 3315 -805
rect 3365 -835 3395 -805
rect 3525 -835 3555 -805
rect 3605 -835 3635 -805
rect 3685 -835 3715 -805
rect 3845 -835 3875 -805
rect 3925 -835 3955 -805
rect 4005 -835 4035 -805
rect 4165 -835 4195 -805
rect 4245 -835 4275 -805
rect 4325 -835 4355 -805
rect 4485 -835 4515 -805
rect 4565 -835 4595 -805
rect 4645 -835 4675 -805
rect 4805 -835 4835 -805
rect 4885 -835 4915 -805
rect 4965 -835 4995 -805
rect 5125 -835 5155 -805
rect -155 -995 -125 -965
rect 5 -995 35 -965
rect 85 -995 115 -965
rect 165 -995 195 -965
rect 325 -995 355 -965
rect 405 -995 435 -965
rect 485 -995 515 -965
rect 645 -995 675 -965
rect 725 -995 755 -965
rect 805 -995 835 -965
rect 965 -995 995 -965
rect 1045 -995 1075 -965
rect 1125 -995 1155 -965
rect 1285 -995 1315 -965
rect 1365 -995 1395 -965
rect 1445 -995 1475 -965
rect 1605 -995 1635 -965
rect 1685 -995 1715 -965
rect 1765 -995 1795 -965
rect 1925 -995 1955 -965
rect 2005 -995 2035 -965
rect 2085 -995 2115 -965
rect 2245 -995 2275 -965
rect 2325 -995 2355 -965
rect 2405 -995 2435 -965
rect 2565 -995 2595 -965
rect 2645 -995 2675 -965
rect 2725 -995 2755 -965
rect 2885 -995 2915 -965
rect 2965 -995 2995 -965
rect 3045 -995 3075 -965
rect 3205 -995 3235 -965
rect 3285 -995 3315 -965
rect 3365 -995 3395 -965
rect 3525 -995 3555 -965
rect 3605 -995 3635 -965
rect 3685 -995 3715 -965
rect 3845 -995 3875 -965
rect 3925 -995 3955 -965
rect 4005 -995 4035 -965
rect 4165 -995 4195 -965
rect 4245 -995 4275 -965
rect 4325 -995 4355 -965
rect 4485 -995 4515 -965
rect 4565 -995 4595 -965
rect 4645 -995 4675 -965
rect 4805 -995 4835 -965
rect 4885 -995 4915 -965
rect 4965 -995 4995 -965
rect 5125 -995 5155 -965
rect -155 -1155 -125 -1125
rect 5 -1155 35 -1125
rect 85 -1155 115 -1125
rect 165 -1155 195 -1125
rect 325 -1155 355 -1125
rect 405 -1155 435 -1125
rect 485 -1155 515 -1125
rect 645 -1155 675 -1125
rect 725 -1155 755 -1125
rect 805 -1155 835 -1125
rect 965 -1155 995 -1125
rect 1045 -1155 1075 -1125
rect 1125 -1155 1155 -1125
rect 1285 -1155 1315 -1125
rect 1365 -1155 1395 -1125
rect 1445 -1155 1475 -1125
rect 1605 -1155 1635 -1125
rect 1685 -1155 1715 -1125
rect 1765 -1155 1795 -1125
rect 1925 -1155 1955 -1125
rect 2005 -1155 2035 -1125
rect 2085 -1155 2115 -1125
rect 2245 -1155 2275 -1125
rect 2325 -1155 2355 -1125
rect 2405 -1155 2435 -1125
rect 2565 -1155 2595 -1125
rect 2645 -1155 2675 -1125
rect 2725 -1155 2755 -1125
rect 2885 -1155 2915 -1125
rect 2965 -1155 2995 -1125
rect 3045 -1155 3075 -1125
rect 3205 -1155 3235 -1125
rect 3285 -1155 3315 -1125
rect 3365 -1155 3395 -1125
rect 3525 -1155 3555 -1125
rect 3605 -1155 3635 -1125
rect 3685 -1155 3715 -1125
rect 3845 -1155 3875 -1125
rect 3925 -1155 3955 -1125
rect 4005 -1155 4035 -1125
rect 4165 -1155 4195 -1125
rect 4245 -1155 4275 -1125
rect 4325 -1155 4355 -1125
rect 4485 -1155 4515 -1125
rect 4565 -1155 4595 -1125
rect 4645 -1155 4675 -1125
rect 4805 -1155 4835 -1125
rect 4885 -1155 4915 -1125
rect 4965 -1155 4995 -1125
rect 5125 -1155 5155 -1125
rect -235 -1235 -205 -1205
rect 5205 -1235 5235 -1205
rect -235 -1510 -205 -1360
rect 5205 -1510 5235 -1360
<< metal3 >>
rect -240 -485 -200 -480
rect -240 -515 -235 -485
rect -205 -515 -200 -485
rect -240 -645 -200 -515
rect -240 -675 -235 -645
rect -205 -675 -200 -645
rect -240 -725 -200 -675
rect -240 -755 -235 -725
rect -205 -755 -200 -725
rect -240 -1205 -200 -755
rect 5200 -485 5240 -480
rect 5200 -515 5205 -485
rect 5235 -515 5240 -485
rect 5200 -645 5240 -515
rect 5200 -675 5205 -645
rect 5235 -675 5240 -645
rect 5200 -725 5240 -675
rect 5200 -755 5205 -725
rect 5235 -755 5240 -725
rect -160 -805 -120 -800
rect -160 -835 -155 -805
rect -125 -835 -120 -805
rect -160 -965 -120 -835
rect -160 -995 -155 -965
rect -125 -995 -120 -965
rect -160 -1125 -120 -995
rect -160 -1155 -155 -1125
rect -125 -1155 -120 -1125
rect -160 -1160 -120 -1155
rect -80 -1160 -40 -800
rect 0 -805 40 -800
rect 0 -835 5 -805
rect 35 -835 40 -805
rect 0 -965 40 -835
rect 0 -995 5 -965
rect 35 -995 40 -965
rect 0 -1125 40 -995
rect 0 -1155 5 -1125
rect 35 -1155 40 -1125
rect 0 -1160 40 -1155
rect 80 -805 120 -800
rect 80 -835 85 -805
rect 115 -835 120 -805
rect 80 -965 120 -835
rect 80 -995 85 -965
rect 115 -995 120 -965
rect 80 -1125 120 -995
rect 80 -1155 85 -1125
rect 115 -1155 120 -1125
rect 80 -1160 120 -1155
rect 160 -805 200 -800
rect 160 -835 165 -805
rect 195 -835 200 -805
rect 160 -965 200 -835
rect 160 -995 165 -965
rect 195 -995 200 -965
rect 160 -1125 200 -995
rect 160 -1155 165 -1125
rect 195 -1155 200 -1125
rect 160 -1160 200 -1155
rect 320 -805 360 -800
rect 320 -835 325 -805
rect 355 -835 360 -805
rect 320 -965 360 -835
rect 320 -995 325 -965
rect 355 -995 360 -965
rect 320 -1125 360 -995
rect 320 -1155 325 -1125
rect 355 -1155 360 -1125
rect 320 -1160 360 -1155
rect 400 -805 440 -800
rect 400 -835 405 -805
rect 435 -835 440 -805
rect 400 -965 440 -835
rect 400 -995 405 -965
rect 435 -995 440 -965
rect 400 -1125 440 -995
rect 400 -1155 405 -1125
rect 435 -1155 440 -1125
rect 400 -1160 440 -1155
rect 480 -805 520 -800
rect 480 -835 485 -805
rect 515 -835 520 -805
rect 480 -965 520 -835
rect 480 -995 485 -965
rect 515 -995 520 -965
rect 480 -1125 520 -995
rect 480 -1155 485 -1125
rect 515 -1155 520 -1125
rect 480 -1160 520 -1155
rect 560 -1160 600 -800
rect 640 -805 680 -800
rect 640 -835 645 -805
rect 675 -835 680 -805
rect 640 -965 680 -835
rect 640 -995 645 -965
rect 675 -995 680 -965
rect 640 -1125 680 -995
rect 640 -1155 645 -1125
rect 675 -1155 680 -1125
rect 640 -1160 680 -1155
rect 720 -805 760 -800
rect 720 -835 725 -805
rect 755 -835 760 -805
rect 720 -965 760 -835
rect 720 -995 725 -965
rect 755 -995 760 -965
rect 720 -1125 760 -995
rect 720 -1155 725 -1125
rect 755 -1155 760 -1125
rect 720 -1160 760 -1155
rect 800 -805 840 -800
rect 800 -835 805 -805
rect 835 -835 840 -805
rect 800 -965 840 -835
rect 800 -995 805 -965
rect 835 -995 840 -965
rect 800 -1125 840 -995
rect 800 -1155 805 -1125
rect 835 -1155 840 -1125
rect 800 -1160 840 -1155
rect 960 -805 1000 -800
rect 960 -835 965 -805
rect 995 -835 1000 -805
rect 960 -965 1000 -835
rect 960 -995 965 -965
rect 995 -995 1000 -965
rect 960 -1125 1000 -995
rect 960 -1155 965 -1125
rect 995 -1155 1000 -1125
rect 960 -1160 1000 -1155
rect 1040 -805 1080 -800
rect 1040 -835 1045 -805
rect 1075 -835 1080 -805
rect 1040 -965 1080 -835
rect 1040 -995 1045 -965
rect 1075 -995 1080 -965
rect 1040 -1125 1080 -995
rect 1040 -1155 1045 -1125
rect 1075 -1155 1080 -1125
rect 1040 -1160 1080 -1155
rect 1120 -805 1160 -800
rect 1120 -835 1125 -805
rect 1155 -835 1160 -805
rect 1120 -965 1160 -835
rect 1120 -995 1125 -965
rect 1155 -995 1160 -965
rect 1120 -1125 1160 -995
rect 1120 -1155 1125 -1125
rect 1155 -1155 1160 -1125
rect 1120 -1160 1160 -1155
rect 1200 -1160 1240 -800
rect 1280 -805 1320 -800
rect 1280 -835 1285 -805
rect 1315 -835 1320 -805
rect 1280 -965 1320 -835
rect 1280 -995 1285 -965
rect 1315 -995 1320 -965
rect 1280 -1125 1320 -995
rect 1280 -1155 1285 -1125
rect 1315 -1155 1320 -1125
rect 1280 -1160 1320 -1155
rect 1360 -805 1400 -800
rect 1360 -835 1365 -805
rect 1395 -835 1400 -805
rect 1360 -965 1400 -835
rect 1360 -995 1365 -965
rect 1395 -995 1400 -965
rect 1360 -1125 1400 -995
rect 1360 -1155 1365 -1125
rect 1395 -1155 1400 -1125
rect 1360 -1160 1400 -1155
rect 1440 -805 1480 -800
rect 1440 -835 1445 -805
rect 1475 -835 1480 -805
rect 1440 -965 1480 -835
rect 1440 -995 1445 -965
rect 1475 -995 1480 -965
rect 1440 -1125 1480 -995
rect 1440 -1155 1445 -1125
rect 1475 -1155 1480 -1125
rect 1440 -1160 1480 -1155
rect 1600 -805 1640 -800
rect 1600 -835 1605 -805
rect 1635 -835 1640 -805
rect 1600 -965 1640 -835
rect 1600 -995 1605 -965
rect 1635 -995 1640 -965
rect 1600 -1125 1640 -995
rect 1600 -1155 1605 -1125
rect 1635 -1155 1640 -1125
rect 1600 -1160 1640 -1155
rect 1680 -805 1720 -800
rect 1680 -835 1685 -805
rect 1715 -835 1720 -805
rect 1680 -965 1720 -835
rect 1680 -995 1685 -965
rect 1715 -995 1720 -965
rect 1680 -1125 1720 -995
rect 1680 -1155 1685 -1125
rect 1715 -1155 1720 -1125
rect 1680 -1160 1720 -1155
rect 1760 -805 1800 -800
rect 1760 -835 1765 -805
rect 1795 -835 1800 -805
rect 1760 -965 1800 -835
rect 1760 -995 1765 -965
rect 1795 -995 1800 -965
rect 1760 -1125 1800 -995
rect 1760 -1155 1765 -1125
rect 1795 -1155 1800 -1125
rect 1760 -1160 1800 -1155
rect 1840 -1160 1880 -800
rect 1920 -805 1960 -800
rect 1920 -835 1925 -805
rect 1955 -835 1960 -805
rect 1920 -965 1960 -835
rect 1920 -995 1925 -965
rect 1955 -995 1960 -965
rect 1920 -1125 1960 -995
rect 1920 -1155 1925 -1125
rect 1955 -1155 1960 -1125
rect 1920 -1160 1960 -1155
rect 2000 -805 2040 -800
rect 2000 -835 2005 -805
rect 2035 -835 2040 -805
rect 2000 -965 2040 -835
rect 2000 -995 2005 -965
rect 2035 -995 2040 -965
rect 2000 -1125 2040 -995
rect 2000 -1155 2005 -1125
rect 2035 -1155 2040 -1125
rect 2000 -1160 2040 -1155
rect 2080 -805 2120 -800
rect 2080 -835 2085 -805
rect 2115 -835 2120 -805
rect 2080 -965 2120 -835
rect 2080 -995 2085 -965
rect 2115 -995 2120 -965
rect 2080 -1125 2120 -995
rect 2080 -1155 2085 -1125
rect 2115 -1155 2120 -1125
rect 2080 -1160 2120 -1155
rect 2240 -805 2280 -800
rect 2240 -835 2245 -805
rect 2275 -835 2280 -805
rect 2240 -965 2280 -835
rect 2240 -995 2245 -965
rect 2275 -995 2280 -965
rect 2240 -1125 2280 -995
rect 2240 -1155 2245 -1125
rect 2275 -1155 2280 -1125
rect 2240 -1160 2280 -1155
rect 2320 -805 2360 -800
rect 2320 -835 2325 -805
rect 2355 -835 2360 -805
rect 2320 -965 2360 -835
rect 2320 -995 2325 -965
rect 2355 -995 2360 -965
rect 2320 -1125 2360 -995
rect 2320 -1155 2325 -1125
rect 2355 -1155 2360 -1125
rect 2320 -1160 2360 -1155
rect 2400 -805 2440 -800
rect 2400 -835 2405 -805
rect 2435 -835 2440 -805
rect 2400 -965 2440 -835
rect 2400 -995 2405 -965
rect 2435 -995 2440 -965
rect 2400 -1125 2440 -995
rect 2400 -1155 2405 -1125
rect 2435 -1155 2440 -1125
rect 2400 -1160 2440 -1155
rect 2480 -1160 2520 -800
rect 2560 -805 2600 -800
rect 2560 -835 2565 -805
rect 2595 -835 2600 -805
rect 2560 -965 2600 -835
rect 2560 -995 2565 -965
rect 2595 -995 2600 -965
rect 2560 -1125 2600 -995
rect 2560 -1155 2565 -1125
rect 2595 -1155 2600 -1125
rect 2560 -1160 2600 -1155
rect 2640 -805 2680 -800
rect 2640 -835 2645 -805
rect 2675 -835 2680 -805
rect 2640 -965 2680 -835
rect 2640 -995 2645 -965
rect 2675 -995 2680 -965
rect 2640 -1125 2680 -995
rect 2640 -1155 2645 -1125
rect 2675 -1155 2680 -1125
rect 2640 -1160 2680 -1155
rect 2720 -805 2760 -800
rect 2720 -835 2725 -805
rect 2755 -835 2760 -805
rect 2720 -965 2760 -835
rect 2720 -995 2725 -965
rect 2755 -995 2760 -965
rect 2720 -1125 2760 -995
rect 2720 -1155 2725 -1125
rect 2755 -1155 2760 -1125
rect 2720 -1160 2760 -1155
rect 2880 -805 2920 -800
rect 2880 -835 2885 -805
rect 2915 -835 2920 -805
rect 2880 -965 2920 -835
rect 2880 -995 2885 -965
rect 2915 -995 2920 -965
rect 2880 -1125 2920 -995
rect 2880 -1155 2885 -1125
rect 2915 -1155 2920 -1125
rect 2880 -1160 2920 -1155
rect 2960 -805 3000 -800
rect 2960 -835 2965 -805
rect 2995 -835 3000 -805
rect 2960 -965 3000 -835
rect 2960 -995 2965 -965
rect 2995 -995 3000 -965
rect 2960 -1125 3000 -995
rect 2960 -1155 2965 -1125
rect 2995 -1155 3000 -1125
rect 2960 -1160 3000 -1155
rect 3040 -805 3080 -800
rect 3040 -835 3045 -805
rect 3075 -835 3080 -805
rect 3040 -965 3080 -835
rect 3040 -995 3045 -965
rect 3075 -995 3080 -965
rect 3040 -1125 3080 -995
rect 3040 -1155 3045 -1125
rect 3075 -1155 3080 -1125
rect 3040 -1160 3080 -1155
rect 3120 -1160 3160 -800
rect 3200 -805 3240 -800
rect 3200 -835 3205 -805
rect 3235 -835 3240 -805
rect 3200 -965 3240 -835
rect 3200 -995 3205 -965
rect 3235 -995 3240 -965
rect 3200 -1125 3240 -995
rect 3200 -1155 3205 -1125
rect 3235 -1155 3240 -1125
rect 3200 -1160 3240 -1155
rect 3280 -805 3320 -800
rect 3280 -835 3285 -805
rect 3315 -835 3320 -805
rect 3280 -965 3320 -835
rect 3280 -995 3285 -965
rect 3315 -995 3320 -965
rect 3280 -1125 3320 -995
rect 3280 -1155 3285 -1125
rect 3315 -1155 3320 -1125
rect 3280 -1160 3320 -1155
rect 3360 -805 3400 -800
rect 3360 -835 3365 -805
rect 3395 -835 3400 -805
rect 3360 -965 3400 -835
rect 3360 -995 3365 -965
rect 3395 -995 3400 -965
rect 3360 -1125 3400 -995
rect 3360 -1155 3365 -1125
rect 3395 -1155 3400 -1125
rect 3360 -1160 3400 -1155
rect 3520 -805 3560 -800
rect 3520 -835 3525 -805
rect 3555 -835 3560 -805
rect 3520 -965 3560 -835
rect 3520 -995 3525 -965
rect 3555 -995 3560 -965
rect 3520 -1125 3560 -995
rect 3520 -1155 3525 -1125
rect 3555 -1155 3560 -1125
rect 3520 -1160 3560 -1155
rect 3600 -805 3640 -800
rect 3600 -835 3605 -805
rect 3635 -835 3640 -805
rect 3600 -965 3640 -835
rect 3600 -995 3605 -965
rect 3635 -995 3640 -965
rect 3600 -1125 3640 -995
rect 3600 -1155 3605 -1125
rect 3635 -1155 3640 -1125
rect 3600 -1160 3640 -1155
rect 3680 -805 3720 -800
rect 3680 -835 3685 -805
rect 3715 -835 3720 -805
rect 3680 -965 3720 -835
rect 3680 -995 3685 -965
rect 3715 -995 3720 -965
rect 3680 -1125 3720 -995
rect 3680 -1155 3685 -1125
rect 3715 -1155 3720 -1125
rect 3680 -1160 3720 -1155
rect 3760 -1160 3800 -800
rect 3840 -805 3880 -800
rect 3840 -835 3845 -805
rect 3875 -835 3880 -805
rect 3840 -965 3880 -835
rect 3840 -995 3845 -965
rect 3875 -995 3880 -965
rect 3840 -1125 3880 -995
rect 3840 -1155 3845 -1125
rect 3875 -1155 3880 -1125
rect 3840 -1160 3880 -1155
rect 3920 -805 3960 -800
rect 3920 -835 3925 -805
rect 3955 -835 3960 -805
rect 3920 -965 3960 -835
rect 3920 -995 3925 -965
rect 3955 -995 3960 -965
rect 3920 -1125 3960 -995
rect 3920 -1155 3925 -1125
rect 3955 -1155 3960 -1125
rect 3920 -1160 3960 -1155
rect 4000 -805 4040 -800
rect 4000 -835 4005 -805
rect 4035 -835 4040 -805
rect 4000 -965 4040 -835
rect 4000 -995 4005 -965
rect 4035 -995 4040 -965
rect 4000 -1125 4040 -995
rect 4000 -1155 4005 -1125
rect 4035 -1155 4040 -1125
rect 4000 -1160 4040 -1155
rect 4160 -805 4200 -800
rect 4160 -835 4165 -805
rect 4195 -835 4200 -805
rect 4160 -965 4200 -835
rect 4160 -995 4165 -965
rect 4195 -995 4200 -965
rect 4160 -1125 4200 -995
rect 4160 -1155 4165 -1125
rect 4195 -1155 4200 -1125
rect 4160 -1160 4200 -1155
rect 4240 -805 4280 -800
rect 4240 -835 4245 -805
rect 4275 -835 4280 -805
rect 4240 -965 4280 -835
rect 4240 -995 4245 -965
rect 4275 -995 4280 -965
rect 4240 -1125 4280 -995
rect 4240 -1155 4245 -1125
rect 4275 -1155 4280 -1125
rect 4240 -1160 4280 -1155
rect 4320 -805 4360 -800
rect 4320 -835 4325 -805
rect 4355 -835 4360 -805
rect 4320 -965 4360 -835
rect 4320 -995 4325 -965
rect 4355 -995 4360 -965
rect 4320 -1125 4360 -995
rect 4320 -1155 4325 -1125
rect 4355 -1155 4360 -1125
rect 4320 -1160 4360 -1155
rect 4400 -1160 4440 -800
rect 4480 -805 4520 -800
rect 4480 -835 4485 -805
rect 4515 -835 4520 -805
rect 4480 -965 4520 -835
rect 4480 -995 4485 -965
rect 4515 -995 4520 -965
rect 4480 -1125 4520 -995
rect 4480 -1155 4485 -1125
rect 4515 -1155 4520 -1125
rect 4480 -1160 4520 -1155
rect 4560 -805 4600 -800
rect 4560 -835 4565 -805
rect 4595 -835 4600 -805
rect 4560 -965 4600 -835
rect 4560 -995 4565 -965
rect 4595 -995 4600 -965
rect 4560 -1125 4600 -995
rect 4560 -1155 4565 -1125
rect 4595 -1155 4600 -1125
rect 4560 -1160 4600 -1155
rect 4640 -805 4680 -800
rect 4640 -835 4645 -805
rect 4675 -835 4680 -805
rect 4640 -965 4680 -835
rect 4640 -995 4645 -965
rect 4675 -995 4680 -965
rect 4640 -1125 4680 -995
rect 4640 -1155 4645 -1125
rect 4675 -1155 4680 -1125
rect 4640 -1160 4680 -1155
rect 4800 -805 4840 -800
rect 4800 -835 4805 -805
rect 4835 -835 4840 -805
rect 4800 -965 4840 -835
rect 4800 -995 4805 -965
rect 4835 -995 4840 -965
rect 4800 -1125 4840 -995
rect 4800 -1155 4805 -1125
rect 4835 -1155 4840 -1125
rect 4800 -1160 4840 -1155
rect 4880 -805 4920 -800
rect 4880 -835 4885 -805
rect 4915 -835 4920 -805
rect 4880 -965 4920 -835
rect 4880 -995 4885 -965
rect 4915 -995 4920 -965
rect 4880 -1125 4920 -995
rect 4880 -1155 4885 -1125
rect 4915 -1155 4920 -1125
rect 4880 -1160 4920 -1155
rect 4960 -805 5000 -800
rect 4960 -835 4965 -805
rect 4995 -835 5000 -805
rect 4960 -965 5000 -835
rect 4960 -995 4965 -965
rect 4995 -995 5000 -965
rect 4960 -1125 5000 -995
rect 4960 -1155 4965 -1125
rect 4995 -1155 5000 -1125
rect 4960 -1160 5000 -1155
rect 5040 -1160 5080 -800
rect 5120 -805 5160 -800
rect 5120 -835 5125 -805
rect 5155 -835 5160 -805
rect 5120 -965 5160 -835
rect 5120 -995 5125 -965
rect 5155 -995 5160 -965
rect 5120 -1125 5160 -995
rect 5120 -1155 5125 -1125
rect 5155 -1155 5160 -1125
rect 5120 -1160 5160 -1155
rect -240 -1235 -235 -1205
rect -205 -1235 -200 -1205
rect -240 -1329 -200 -1235
rect -240 -1511 -236 -1329
rect -204 -1511 -200 -1329
rect -240 -1520 -200 -1511
rect 5200 -1205 5240 -755
rect 5200 -1235 5205 -1205
rect 5235 -1235 5240 -1205
rect 5200 -1329 5240 -1235
rect 5200 -1511 5204 -1329
rect 5236 -1511 5240 -1329
rect 5200 -1520 5240 -1511
<< via3 >>
rect -236 -1360 -204 -1329
rect -236 -1510 -235 -1360
rect -235 -1510 -205 -1360
rect -205 -1510 -204 -1360
rect -236 -1511 -204 -1510
rect 5204 -1360 5236 -1329
rect 5204 -1510 5205 -1360
rect 5205 -1510 5235 -1360
rect 5235 -1510 5236 -1360
rect 5204 -1511 5236 -1510
<< metal4 >>
rect -240 -280 5240 -240
rect -240 -400 -120 -280
rect 0 -400 1160 -280
rect 1280 -400 2440 -280
rect 2560 -400 3720 -280
rect 3840 -400 5000 -280
rect 5120 -400 5240 -280
rect -240 -440 5240 -400
rect -240 -1329 5240 -1320
rect -240 -1511 -236 -1329
rect -204 -1360 5204 -1329
rect -204 -1480 520 -1360
rect 640 -1480 1800 -1360
rect 1920 -1480 3080 -1360
rect 3200 -1480 4360 -1360
rect 4480 -1480 5204 -1360
rect -204 -1511 5204 -1480
rect 5236 -1511 5240 -1329
rect -240 -1520 5240 -1511
<< via4 >>
rect -120 -400 0 -280
rect 1160 -400 1280 -280
rect 2440 -400 2560 -280
rect 3720 -400 3840 -280
rect 5000 -400 5120 -280
rect 520 -1480 640 -1360
rect 1800 -1480 1920 -1360
rect 3080 -1480 3200 -1360
rect 4360 -1480 4480 -1360
<< metal5 >>
rect -160 -280 40 -80
rect -160 -400 -120 -280
rect 0 -400 40 -280
rect -160 -1520 40 -400
rect 480 -1360 680 -80
rect 480 -1480 520 -1360
rect 640 -1480 680 -1360
rect 480 -1520 680 -1480
rect 1120 -280 1320 -80
rect 1120 -400 1160 -280
rect 1280 -400 1320 -280
rect 1120 -1520 1320 -400
rect 1760 -1360 1960 -80
rect 1760 -1480 1800 -1360
rect 1920 -1480 1960 -1360
rect 1760 -1520 1960 -1480
rect 2400 -280 2600 -80
rect 2400 -400 2440 -280
rect 2560 -400 2600 -280
rect 2400 -1520 2600 -400
rect 3040 -1360 3240 -80
rect 3040 -1480 3080 -1360
rect 3200 -1480 3240 -1360
rect 3040 -1520 3240 -1480
rect 3680 -280 3880 -80
rect 3680 -400 3720 -280
rect 3840 -400 3880 -280
rect 3680 -1520 3880 -400
rect 4320 -1360 4520 -80
rect 4320 -1480 4360 -1360
rect 4480 -1480 4520 -1360
rect 4320 -1520 4520 -1480
rect 4960 -280 5160 -80
rect 4960 -400 5000 -280
rect 5120 -400 5160 -280
rect 4960 -1520 5160 -400
<< labels >>
rlabel metal2 5200 -200 5240 -160 0 gpa
port 0 nsew
rlabel metal2 5200 -600 5240 -560 0 gpb
port 1 nsew
rlabel metal2 5200 -920 5240 -880 0 dp
port 2 nsew
rlabel metal2 5200 -1000 5240 -960 0 out
port 3 nsew
rlabel metal2 5200 -1080 5240 -1040 0 dn
port 4 nsew
rlabel metal2 5200 -1320 5240 -1280 0 gnb
port 5 nsew
rlabel metal5 -160 -120 40 -80 0 vdda
port 6 nsew
rlabel metal5 480 -120 680 -80 0 vssa
port 7 nsew
<< end >>
