magic
tech sky130A
timestamp 1623884123
<< nwell >>
rect -420 640 11285 1200
<< nmos >>
rect -310 1690 -260 1790
rect -220 1690 -170 1790
rect -130 1690 -80 1790
rect -40 1690 10 1790
rect 50 1690 100 1790
rect 140 1690 190 1790
rect 230 1690 280 1790
rect 320 1690 370 1790
rect 410 1690 460 1790
rect 500 1690 550 1790
rect 590 1690 640 1790
rect 680 1690 730 1790
rect 770 1690 820 1790
rect 860 1690 910 1790
rect 950 1690 1000 1790
rect 1040 1690 1090 1790
rect 1130 1690 1180 1790
rect 1220 1690 1270 1790
rect 1310 1690 1360 1790
rect 1400 1690 1450 1790
rect 1490 1690 1540 1790
rect 1580 1690 1630 1790
rect 1670 1690 1720 1790
rect 1760 1690 1810 1790
rect 1850 1690 1900 1790
rect 1940 1690 1990 1790
rect 2030 1690 2080 1790
rect 2120 1690 2170 1790
rect 2210 1690 2260 1790
rect 2300 1690 2350 1790
rect 2390 1690 2440 1790
rect 2480 1690 2530 1790
rect 2570 1690 2620 1790
rect 2660 1690 2710 1790
rect 2750 1690 2800 1790
rect 2840 1690 2890 1790
rect 2930 1690 2980 1790
rect 3020 1690 3070 1790
rect 3115 1690 3165 1790
rect 3205 1690 3255 1790
rect 3295 1690 3345 1790
rect 3385 1690 3435 1790
rect 3475 1690 3525 1790
rect 3565 1690 3615 1790
rect 3655 1690 3705 1790
rect 3745 1690 3795 1790
rect 3835 1690 3885 1790
rect 3925 1690 3975 1790
rect 4015 1690 4065 1790
rect 4105 1690 4155 1790
rect 4195 1690 4245 1790
rect 4285 1690 4335 1790
rect 4375 1690 4425 1790
rect 4465 1690 4515 1790
rect 4555 1690 4605 1790
rect 4645 1690 4695 1790
rect 4735 1690 4785 1790
rect 4825 1690 4875 1790
rect 4915 1690 4965 1790
rect 5005 1690 5055 1790
rect 5095 1690 5145 1790
rect 5185 1690 5235 1790
rect 5275 1690 5325 1790
rect 5365 1690 5415 1790
rect 5455 1690 5505 1790
rect 5545 1690 5595 1790
rect 5635 1690 5685 1790
rect 5725 1690 5775 1790
rect 5815 1690 5865 1790
rect 5905 1690 5955 1790
rect 5995 1690 6045 1790
rect 6085 1690 6135 1790
rect 6175 1690 6225 1790
rect 6265 1690 6315 1790
rect 6355 1690 6405 1790
rect 6445 1690 6495 1790
rect 6535 1690 6585 1790
rect 6625 1690 6675 1790
rect 6715 1690 6765 1790
rect 6805 1690 6855 1790
rect 6895 1690 6945 1790
rect 6985 1690 7035 1790
rect 7075 1690 7125 1790
rect 7165 1690 7215 1790
rect 7255 1690 7305 1790
rect 7345 1690 7395 1790
rect 7435 1690 7485 1790
rect 7525 1690 7575 1790
rect 7615 1690 7665 1790
rect 7705 1690 7755 1790
rect 7795 1690 7845 1790
rect 7885 1690 7935 1790
rect 7975 1690 8025 1790
rect 8065 1690 8115 1790
rect 8155 1690 8205 1790
rect 8245 1690 8295 1790
rect 8335 1690 8385 1790
rect 8425 1690 8475 1790
rect 8515 1690 8565 1790
rect 8605 1690 8655 1790
rect 8695 1690 8745 1790
rect 8785 1690 8835 1790
rect 8875 1690 8925 1790
rect 8965 1690 9015 1790
rect 9055 1690 9105 1790
rect 9145 1690 9195 1790
rect 9235 1690 9285 1790
rect 9325 1690 9375 1790
rect 9415 1690 9465 1790
rect 9505 1690 9555 1790
rect 9595 1690 9645 1790
rect 9685 1690 9735 1790
rect 9775 1690 9825 1790
rect 9865 1690 9915 1790
rect 9955 1690 10005 1790
rect 10045 1690 10095 1790
rect 10135 1690 10185 1790
rect 10225 1690 10275 1790
rect 10315 1690 10365 1790
rect 10405 1690 10455 1790
rect 10495 1690 10545 1790
rect 10585 1690 10635 1790
rect 10675 1690 10725 1790
rect 10765 1690 10815 1790
rect 10855 1690 10905 1790
rect 10945 1690 10995 1790
rect 11035 1690 11085 1790
rect 11125 1690 11175 1790
rect -310 50 -260 150
rect -220 50 -170 150
rect -130 50 -80 150
rect -40 50 10 150
rect 50 50 100 150
rect 140 50 190 150
rect 230 50 280 150
rect 320 50 370 150
rect 410 50 460 150
rect 500 50 550 150
rect 590 50 640 150
rect 680 50 730 150
rect 770 50 820 150
rect 860 50 910 150
rect 950 50 1000 150
rect 1040 50 1090 150
rect 1130 50 1180 150
rect 1220 50 1270 150
rect 1310 50 1360 150
rect 1400 50 1450 150
rect 1490 50 1540 150
rect 1580 50 1630 150
rect 1670 50 1720 150
rect 1760 50 1810 150
rect 1850 50 1900 150
rect 1940 50 1990 150
rect 2030 50 2080 150
rect 2120 50 2170 150
rect 2210 50 2260 150
rect 2300 50 2350 150
rect 2390 50 2440 150
rect 2480 50 2530 150
rect 2570 50 2620 150
rect 2660 50 2710 150
rect 2750 50 2800 150
rect 2840 50 2890 150
rect 2930 50 2980 150
rect 3020 50 3070 150
rect 3110 50 3160 150
rect 3200 50 3250 150
rect 3290 50 3340 150
rect 3380 50 3430 150
rect 3470 50 3520 150
rect 3560 50 3610 150
rect 3650 50 3700 150
rect 3740 50 3790 150
rect 3830 50 3880 150
rect 3920 50 3970 150
rect 4010 50 4060 150
rect 4100 50 4150 150
rect 4190 50 4240 150
rect 4280 50 4330 150
rect 4370 50 4420 150
rect 4460 50 4510 150
rect 4550 50 4600 150
rect 4640 50 4690 150
rect 4730 50 4780 150
rect 4820 50 4870 150
rect 4910 50 4960 150
rect 5000 50 5050 150
rect 5090 50 5140 150
rect 5180 50 5230 150
rect 5270 50 5320 150
rect 5360 50 5410 150
rect 5450 50 5500 150
rect 5540 50 5590 150
rect 5630 50 5680 150
rect 5720 50 5770 150
rect 5810 50 5860 150
rect 5900 50 5950 150
rect 5990 50 6040 150
rect 6080 50 6130 150
rect 6170 50 6220 150
rect 6260 50 6310 150
rect 6350 50 6400 150
rect 6440 50 6490 150
rect 6530 50 6580 150
rect 6620 50 6670 150
rect 6710 50 6760 150
rect 6800 50 6850 150
rect 6890 50 6940 150
rect 6980 50 7030 150
rect 7070 50 7120 150
rect 7160 50 7210 150
rect 7250 50 7300 150
rect 7340 50 7390 150
rect 7430 50 7480 150
rect 7520 50 7570 150
rect 7610 50 7660 150
rect 7700 50 7750 150
rect 7795 50 7845 150
rect 7885 50 7935 150
rect 7975 50 8025 150
rect 8065 50 8115 150
rect 8155 50 8205 150
rect 8245 50 8295 150
rect 8335 50 8385 150
rect 8425 50 8475 150
rect 8515 50 8565 150
rect 8605 50 8655 150
rect 8695 50 8745 150
rect 8785 50 8835 150
rect 8875 50 8925 150
rect 8965 50 9015 150
rect 9055 50 9105 150
rect 9145 50 9195 150
rect 9235 50 9285 150
rect 9325 50 9375 150
rect 9415 50 9465 150
rect 9505 50 9555 150
rect 9595 50 9645 150
rect 9685 50 9735 150
rect 9775 50 9825 150
rect 9865 50 9915 150
rect 9955 50 10005 150
rect 10045 50 10095 150
rect 10135 50 10185 150
rect 10225 50 10275 150
rect 10315 50 10365 150
rect 10405 50 10455 150
rect 10495 50 10545 150
rect 10585 50 10635 150
rect 10675 50 10725 150
rect 10765 50 10815 150
rect 10855 50 10905 150
rect 10945 50 10995 150
rect 11035 50 11085 150
rect 11125 50 11175 150
<< pmos >>
rect -310 990 -260 1090
rect -220 990 -170 1090
rect -130 990 -80 1090
rect -40 990 10 1090
rect 50 990 100 1090
rect 140 990 190 1090
rect 230 990 280 1090
rect 320 990 370 1090
rect 410 990 460 1090
rect 500 990 550 1090
rect 590 990 640 1090
rect 680 990 730 1090
rect 770 990 820 1090
rect 860 990 910 1090
rect 950 990 1000 1090
rect 1040 990 1090 1090
rect 1130 990 1180 1090
rect 1220 990 1270 1090
rect 1310 990 1360 1090
rect 1400 990 1450 1090
rect 1490 990 1540 1090
rect 1580 990 1630 1090
rect 1670 990 1720 1090
rect 1760 990 1810 1090
rect 1850 990 1900 1090
rect 1940 990 1990 1090
rect 2030 990 2080 1090
rect 2120 990 2170 1090
rect 2210 990 2260 1090
rect 2300 990 2350 1090
rect 2390 990 2440 1090
rect 2480 990 2530 1090
rect 2570 990 2620 1090
rect 2660 990 2710 1090
rect 2750 990 2800 1090
rect 2840 990 2890 1090
rect 2930 990 2980 1090
rect 3020 990 3070 1090
rect 3115 990 3165 1090
rect 3205 990 3255 1090
rect 3295 990 3345 1090
rect 3385 990 3435 1090
rect 3475 990 3525 1090
rect 3565 990 3615 1090
rect 3655 990 3705 1090
rect 3745 990 3795 1090
rect 3835 990 3885 1090
rect 3925 990 3975 1090
rect 4015 990 4065 1090
rect 4105 990 4155 1090
rect 4195 990 4245 1090
rect 4285 990 4335 1090
rect 4375 990 4425 1090
rect 4465 990 4515 1090
rect 4555 990 4605 1090
rect 4645 990 4695 1090
rect 4735 990 4785 1090
rect 4825 990 4875 1090
rect 4915 990 4965 1090
rect 5005 990 5055 1090
rect 5095 990 5145 1090
rect 5185 990 5235 1090
rect 5275 990 5325 1090
rect 5365 990 5415 1090
rect 5455 990 5505 1090
rect 5545 990 5595 1090
rect 5635 990 5685 1090
rect 5725 990 5775 1090
rect 5815 990 5865 1090
rect 5905 990 5955 1090
rect 5995 990 6045 1090
rect 6085 990 6135 1090
rect 6175 990 6225 1090
rect 6265 990 6315 1090
rect 6355 990 6405 1090
rect 6445 990 6495 1090
rect 6535 990 6585 1090
rect 6625 990 6675 1090
rect 6715 990 6765 1090
rect 6805 990 6855 1090
rect 6895 990 6945 1090
rect 6985 990 7035 1090
rect 7075 990 7125 1090
rect 7165 990 7215 1090
rect 7255 990 7305 1090
rect 7345 990 7395 1090
rect 7435 990 7485 1090
rect 7525 990 7575 1090
rect 7615 990 7665 1090
rect 7705 990 7755 1090
rect 7795 990 7845 1090
rect 7885 990 7935 1090
rect 7975 990 8025 1090
rect 8065 990 8115 1090
rect 8155 990 8205 1090
rect 8245 990 8295 1090
rect 8335 990 8385 1090
rect 8425 990 8475 1090
rect 8515 990 8565 1090
rect 8605 990 8655 1090
rect 8695 990 8745 1090
rect 8785 990 8835 1090
rect 8875 990 8925 1090
rect 8965 990 9015 1090
rect 9055 990 9105 1090
rect 9145 990 9195 1090
rect 9235 990 9285 1090
rect 9325 990 9375 1090
rect 9415 990 9465 1090
rect 9505 990 9555 1090
rect 9595 990 9645 1090
rect 9685 990 9735 1090
rect 9775 990 9825 1090
rect 9865 990 9915 1090
rect 9955 990 10005 1090
rect 10045 990 10095 1090
rect 10135 990 10185 1090
rect 10225 990 10275 1090
rect 10315 990 10365 1090
rect 10405 990 10455 1090
rect 10495 990 10545 1090
rect 10585 990 10635 1090
rect 10675 990 10725 1090
rect 10765 990 10815 1090
rect 10855 990 10905 1090
rect 10945 990 10995 1090
rect 11035 990 11085 1090
rect 11125 990 11175 1090
rect -310 750 -260 850
rect -220 750 -170 850
rect -130 750 -80 850
rect -40 750 10 850
rect 50 750 100 850
rect 140 750 190 850
rect 230 750 280 850
rect 320 750 370 850
rect 410 750 460 850
rect 500 750 550 850
rect 590 750 640 850
rect 680 750 730 850
rect 770 750 820 850
rect 860 750 910 850
rect 950 750 1000 850
rect 1040 750 1090 850
rect 1130 750 1180 850
rect 1220 750 1270 850
rect 1310 750 1360 850
rect 1400 750 1450 850
rect 1490 750 1540 850
rect 1580 750 1630 850
rect 1670 750 1720 850
rect 1760 750 1810 850
rect 1850 750 1900 850
rect 1940 750 1990 850
rect 2030 750 2080 850
rect 2120 750 2170 850
rect 2210 750 2260 850
rect 2300 750 2350 850
rect 2390 750 2440 850
rect 2480 750 2530 850
rect 2570 750 2620 850
rect 2660 750 2710 850
rect 2750 750 2800 850
rect 2840 750 2890 850
rect 2930 750 2980 850
rect 3020 750 3070 850
rect 3110 750 3160 850
rect 3200 750 3250 850
rect 3290 750 3340 850
rect 3380 750 3430 850
rect 3470 750 3520 850
rect 3560 750 3610 850
rect 3650 750 3700 850
rect 3740 750 3790 850
rect 3830 750 3880 850
rect 3920 750 3970 850
rect 4010 750 4060 850
rect 4100 750 4150 850
rect 4190 750 4240 850
rect 4280 750 4330 850
rect 4370 750 4420 850
rect 4460 750 4510 850
rect 4550 750 4600 850
rect 4640 750 4690 850
rect 4730 750 4780 850
rect 4820 750 4870 850
rect 4910 750 4960 850
rect 5000 750 5050 850
rect 5090 750 5140 850
rect 5180 750 5230 850
rect 5270 750 5320 850
rect 5360 750 5410 850
rect 5450 750 5500 850
rect 5540 750 5590 850
rect 5630 750 5680 850
rect 5720 750 5770 850
rect 5810 750 5860 850
rect 5900 750 5950 850
rect 5990 750 6040 850
rect 6080 750 6130 850
rect 6170 750 6220 850
rect 6260 750 6310 850
rect 6350 750 6400 850
rect 6440 750 6490 850
rect 6530 750 6580 850
rect 6620 750 6670 850
rect 6710 750 6760 850
rect 6800 750 6850 850
rect 6890 750 6940 850
rect 6980 750 7030 850
rect 7070 750 7120 850
rect 7160 750 7210 850
rect 7250 750 7300 850
rect 7340 750 7390 850
rect 7430 750 7480 850
rect 7520 750 7570 850
rect 7610 750 7660 850
rect 7700 750 7750 850
rect 7795 750 7845 850
rect 7885 750 7935 850
rect 7975 750 8025 850
rect 8065 750 8115 850
rect 8155 750 8205 850
rect 8245 750 8295 850
rect 8335 750 8385 850
rect 8425 750 8475 850
rect 8515 750 8565 850
rect 8605 750 8655 850
rect 8695 750 8745 850
rect 8785 750 8835 850
rect 8875 750 8925 850
rect 8965 750 9015 850
rect 9055 750 9105 850
rect 9145 750 9195 850
rect 9235 750 9285 850
rect 9325 750 9375 850
rect 9415 750 9465 850
rect 9505 750 9555 850
rect 9595 750 9645 850
rect 9685 750 9735 850
rect 9775 750 9825 850
rect 9865 750 9915 850
rect 9955 750 10005 850
rect 10045 750 10095 850
rect 10135 750 10185 850
rect 10225 750 10275 850
rect 10315 750 10365 850
rect 10405 750 10455 850
rect 10495 750 10545 850
rect 10585 750 10635 850
rect 10675 750 10725 850
rect 10765 750 10815 850
rect 10855 750 10905 850
rect 10945 750 10995 850
rect 11035 750 11085 850
rect 11125 750 11175 850
<< ndiff >>
rect -350 1780 -310 1790
rect -350 1700 -340 1780
rect -320 1700 -310 1780
rect -350 1690 -310 1700
rect -260 1780 -220 1790
rect -260 1700 -250 1780
rect -230 1700 -220 1780
rect -260 1690 -220 1700
rect -170 1780 -130 1790
rect -170 1700 -160 1780
rect -140 1700 -130 1780
rect -170 1690 -130 1700
rect -80 1780 -40 1790
rect -80 1700 -70 1780
rect -50 1700 -40 1780
rect -80 1690 -40 1700
rect 10 1780 50 1790
rect 10 1700 20 1780
rect 40 1700 50 1780
rect 10 1690 50 1700
rect 100 1780 140 1790
rect 100 1700 110 1780
rect 130 1700 140 1780
rect 100 1690 140 1700
rect 190 1780 230 1790
rect 190 1700 200 1780
rect 220 1700 230 1780
rect 190 1690 230 1700
rect 280 1780 320 1790
rect 280 1700 290 1780
rect 310 1700 320 1780
rect 280 1690 320 1700
rect 370 1780 410 1790
rect 370 1700 380 1780
rect 400 1700 410 1780
rect 370 1690 410 1700
rect 460 1780 500 1790
rect 460 1700 470 1780
rect 490 1700 500 1780
rect 460 1690 500 1700
rect 550 1780 590 1790
rect 550 1700 560 1780
rect 580 1700 590 1780
rect 550 1690 590 1700
rect 640 1780 680 1790
rect 640 1700 650 1780
rect 670 1700 680 1780
rect 640 1690 680 1700
rect 730 1780 770 1790
rect 730 1700 740 1780
rect 760 1700 770 1780
rect 730 1690 770 1700
rect 820 1780 860 1790
rect 820 1700 830 1780
rect 850 1700 860 1780
rect 820 1690 860 1700
rect 910 1780 950 1790
rect 910 1700 920 1780
rect 940 1700 950 1780
rect 910 1690 950 1700
rect 1000 1780 1040 1790
rect 1000 1700 1010 1780
rect 1030 1700 1040 1780
rect 1000 1690 1040 1700
rect 1090 1780 1130 1790
rect 1090 1700 1100 1780
rect 1120 1700 1130 1780
rect 1090 1690 1130 1700
rect 1180 1780 1220 1790
rect 1180 1700 1190 1780
rect 1210 1700 1220 1780
rect 1180 1690 1220 1700
rect 1270 1780 1310 1790
rect 1270 1700 1280 1780
rect 1300 1700 1310 1780
rect 1270 1690 1310 1700
rect 1360 1780 1400 1790
rect 1360 1700 1370 1780
rect 1390 1700 1400 1780
rect 1360 1690 1400 1700
rect 1450 1780 1490 1790
rect 1450 1700 1460 1780
rect 1480 1700 1490 1780
rect 1450 1690 1490 1700
rect 1540 1780 1580 1790
rect 1540 1700 1550 1780
rect 1570 1700 1580 1780
rect 1540 1690 1580 1700
rect 1630 1780 1670 1790
rect 1630 1700 1640 1780
rect 1660 1700 1670 1780
rect 1630 1690 1670 1700
rect 1720 1780 1760 1790
rect 1720 1700 1730 1780
rect 1750 1700 1760 1780
rect 1720 1690 1760 1700
rect 1810 1780 1850 1790
rect 1810 1700 1820 1780
rect 1840 1700 1850 1780
rect 1810 1690 1850 1700
rect 1900 1780 1940 1790
rect 1900 1700 1910 1780
rect 1930 1700 1940 1780
rect 1900 1690 1940 1700
rect 1990 1780 2030 1790
rect 1990 1700 2000 1780
rect 2020 1700 2030 1780
rect 1990 1690 2030 1700
rect 2080 1780 2120 1790
rect 2080 1700 2090 1780
rect 2110 1700 2120 1780
rect 2080 1690 2120 1700
rect 2170 1780 2210 1790
rect 2170 1700 2180 1780
rect 2200 1700 2210 1780
rect 2170 1690 2210 1700
rect 2260 1780 2300 1790
rect 2260 1700 2270 1780
rect 2290 1700 2300 1780
rect 2260 1690 2300 1700
rect 2350 1780 2390 1790
rect 2350 1700 2360 1780
rect 2380 1700 2390 1780
rect 2350 1690 2390 1700
rect 2440 1780 2480 1790
rect 2440 1700 2450 1780
rect 2470 1700 2480 1780
rect 2440 1690 2480 1700
rect 2530 1780 2570 1790
rect 2530 1700 2540 1780
rect 2560 1700 2570 1780
rect 2530 1690 2570 1700
rect 2620 1780 2660 1790
rect 2620 1700 2630 1780
rect 2650 1700 2660 1780
rect 2620 1690 2660 1700
rect 2710 1780 2750 1790
rect 2710 1700 2720 1780
rect 2740 1700 2750 1780
rect 2710 1690 2750 1700
rect 2800 1780 2840 1790
rect 2800 1700 2810 1780
rect 2830 1700 2840 1780
rect 2800 1690 2840 1700
rect 2890 1780 2930 1790
rect 2890 1700 2900 1780
rect 2920 1700 2930 1780
rect 2890 1690 2930 1700
rect 2980 1780 3020 1790
rect 2980 1700 2990 1780
rect 3010 1700 3020 1780
rect 2980 1690 3020 1700
rect 3070 1780 3115 1790
rect 3070 1700 3085 1780
rect 3105 1700 3115 1780
rect 3070 1690 3115 1700
rect 3165 1780 3205 1790
rect 3165 1700 3175 1780
rect 3195 1700 3205 1780
rect 3165 1690 3205 1700
rect 3255 1780 3295 1790
rect 3255 1700 3265 1780
rect 3285 1700 3295 1780
rect 3255 1690 3295 1700
rect 3345 1780 3385 1790
rect 3345 1700 3355 1780
rect 3375 1700 3385 1780
rect 3345 1690 3385 1700
rect 3435 1780 3475 1790
rect 3435 1700 3445 1780
rect 3465 1700 3475 1780
rect 3435 1690 3475 1700
rect 3525 1780 3565 1790
rect 3525 1700 3535 1780
rect 3555 1700 3565 1780
rect 3525 1690 3565 1700
rect 3615 1780 3655 1790
rect 3615 1700 3625 1780
rect 3645 1700 3655 1780
rect 3615 1690 3655 1700
rect 3705 1780 3745 1790
rect 3705 1700 3715 1780
rect 3735 1700 3745 1780
rect 3705 1690 3745 1700
rect 3795 1780 3835 1790
rect 3795 1700 3805 1780
rect 3825 1700 3835 1780
rect 3795 1690 3835 1700
rect 3885 1780 3925 1790
rect 3885 1700 3895 1780
rect 3915 1700 3925 1780
rect 3885 1690 3925 1700
rect 3975 1780 4015 1790
rect 3975 1700 3985 1780
rect 4005 1700 4015 1780
rect 3975 1690 4015 1700
rect 4065 1780 4105 1790
rect 4065 1700 4075 1780
rect 4095 1700 4105 1780
rect 4065 1690 4105 1700
rect 4155 1780 4195 1790
rect 4155 1700 4165 1780
rect 4185 1700 4195 1780
rect 4155 1690 4195 1700
rect 4245 1780 4285 1790
rect 4245 1700 4255 1780
rect 4275 1700 4285 1780
rect 4245 1690 4285 1700
rect 4335 1780 4375 1790
rect 4335 1700 4345 1780
rect 4365 1700 4375 1780
rect 4335 1690 4375 1700
rect 4425 1780 4465 1790
rect 4425 1700 4435 1780
rect 4455 1700 4465 1780
rect 4425 1690 4465 1700
rect 4515 1780 4555 1790
rect 4515 1700 4525 1780
rect 4545 1700 4555 1780
rect 4515 1690 4555 1700
rect 4605 1780 4645 1790
rect 4605 1700 4615 1780
rect 4635 1700 4645 1780
rect 4605 1690 4645 1700
rect 4695 1780 4735 1790
rect 4695 1700 4705 1780
rect 4725 1700 4735 1780
rect 4695 1690 4735 1700
rect 4785 1780 4825 1790
rect 4785 1700 4795 1780
rect 4815 1700 4825 1780
rect 4785 1690 4825 1700
rect 4875 1780 4915 1790
rect 4875 1700 4885 1780
rect 4905 1700 4915 1780
rect 4875 1690 4915 1700
rect 4965 1780 5005 1790
rect 4965 1700 4975 1780
rect 4995 1700 5005 1780
rect 4965 1690 5005 1700
rect 5055 1780 5095 1790
rect 5055 1700 5065 1780
rect 5085 1700 5095 1780
rect 5055 1690 5095 1700
rect 5145 1780 5185 1790
rect 5145 1700 5155 1780
rect 5175 1700 5185 1780
rect 5145 1690 5185 1700
rect 5235 1780 5275 1790
rect 5235 1700 5245 1780
rect 5265 1700 5275 1780
rect 5235 1690 5275 1700
rect 5325 1780 5365 1790
rect 5325 1700 5335 1780
rect 5355 1700 5365 1780
rect 5325 1690 5365 1700
rect 5415 1780 5455 1790
rect 5415 1700 5425 1780
rect 5445 1700 5455 1780
rect 5415 1690 5455 1700
rect 5505 1780 5545 1790
rect 5505 1700 5515 1780
rect 5535 1700 5545 1780
rect 5505 1690 5545 1700
rect 5595 1780 5635 1790
rect 5595 1700 5605 1780
rect 5625 1700 5635 1780
rect 5595 1690 5635 1700
rect 5685 1780 5725 1790
rect 5685 1700 5695 1780
rect 5715 1700 5725 1780
rect 5685 1690 5725 1700
rect 5775 1780 5815 1790
rect 5775 1700 5785 1780
rect 5805 1700 5815 1780
rect 5775 1690 5815 1700
rect 5865 1780 5905 1790
rect 5865 1700 5875 1780
rect 5895 1700 5905 1780
rect 5865 1690 5905 1700
rect 5955 1780 5995 1790
rect 5955 1700 5965 1780
rect 5985 1700 5995 1780
rect 5955 1690 5995 1700
rect 6045 1780 6085 1790
rect 6045 1700 6055 1780
rect 6075 1700 6085 1780
rect 6045 1690 6085 1700
rect 6135 1780 6175 1790
rect 6135 1700 6145 1780
rect 6165 1700 6175 1780
rect 6135 1690 6175 1700
rect 6225 1780 6265 1790
rect 6225 1700 6235 1780
rect 6255 1700 6265 1780
rect 6225 1690 6265 1700
rect 6315 1780 6355 1790
rect 6315 1700 6325 1780
rect 6345 1700 6355 1780
rect 6315 1690 6355 1700
rect 6405 1780 6445 1790
rect 6405 1700 6415 1780
rect 6435 1700 6445 1780
rect 6405 1690 6445 1700
rect 6495 1780 6535 1790
rect 6495 1700 6505 1780
rect 6525 1700 6535 1780
rect 6495 1690 6535 1700
rect 6585 1780 6625 1790
rect 6585 1700 6595 1780
rect 6615 1700 6625 1780
rect 6585 1690 6625 1700
rect 6675 1780 6715 1790
rect 6675 1700 6685 1780
rect 6705 1700 6715 1780
rect 6675 1690 6715 1700
rect 6765 1780 6805 1790
rect 6765 1700 6775 1780
rect 6795 1700 6805 1780
rect 6765 1690 6805 1700
rect 6855 1780 6895 1790
rect 6855 1700 6865 1780
rect 6885 1700 6895 1780
rect 6855 1690 6895 1700
rect 6945 1780 6985 1790
rect 6945 1700 6955 1780
rect 6975 1700 6985 1780
rect 6945 1690 6985 1700
rect 7035 1780 7075 1790
rect 7035 1700 7045 1780
rect 7065 1700 7075 1780
rect 7035 1690 7075 1700
rect 7125 1780 7165 1790
rect 7125 1700 7135 1780
rect 7155 1700 7165 1780
rect 7125 1690 7165 1700
rect 7215 1780 7255 1790
rect 7215 1700 7225 1780
rect 7245 1700 7255 1780
rect 7215 1690 7255 1700
rect 7305 1780 7345 1790
rect 7305 1700 7315 1780
rect 7335 1700 7345 1780
rect 7305 1690 7345 1700
rect 7395 1780 7435 1790
rect 7395 1700 7405 1780
rect 7425 1700 7435 1780
rect 7395 1690 7435 1700
rect 7485 1780 7525 1790
rect 7485 1700 7495 1780
rect 7515 1700 7525 1780
rect 7485 1690 7525 1700
rect 7575 1780 7615 1790
rect 7575 1700 7585 1780
rect 7605 1700 7615 1780
rect 7575 1690 7615 1700
rect 7665 1780 7705 1790
rect 7665 1700 7675 1780
rect 7695 1700 7705 1780
rect 7665 1690 7705 1700
rect 7755 1780 7795 1790
rect 7755 1700 7765 1780
rect 7785 1700 7795 1780
rect 7755 1690 7795 1700
rect 7845 1780 7885 1790
rect 7845 1700 7855 1780
rect 7875 1700 7885 1780
rect 7845 1690 7885 1700
rect 7935 1780 7975 1790
rect 7935 1700 7945 1780
rect 7965 1700 7975 1780
rect 7935 1690 7975 1700
rect 8025 1780 8065 1790
rect 8025 1700 8035 1780
rect 8055 1700 8065 1780
rect 8025 1690 8065 1700
rect 8115 1780 8155 1790
rect 8115 1700 8125 1780
rect 8145 1700 8155 1780
rect 8115 1690 8155 1700
rect 8205 1780 8245 1790
rect 8205 1700 8215 1780
rect 8235 1700 8245 1780
rect 8205 1690 8245 1700
rect 8295 1780 8335 1790
rect 8295 1700 8305 1780
rect 8325 1700 8335 1780
rect 8295 1690 8335 1700
rect 8385 1780 8425 1790
rect 8385 1700 8395 1780
rect 8415 1700 8425 1780
rect 8385 1690 8425 1700
rect 8475 1780 8515 1790
rect 8475 1700 8485 1780
rect 8505 1700 8515 1780
rect 8475 1690 8515 1700
rect 8565 1780 8605 1790
rect 8565 1700 8575 1780
rect 8595 1700 8605 1780
rect 8565 1690 8605 1700
rect 8655 1780 8695 1790
rect 8655 1700 8665 1780
rect 8685 1700 8695 1780
rect 8655 1690 8695 1700
rect 8745 1780 8785 1790
rect 8745 1700 8755 1780
rect 8775 1700 8785 1780
rect 8745 1690 8785 1700
rect 8835 1780 8875 1790
rect 8835 1700 8845 1780
rect 8865 1700 8875 1780
rect 8835 1690 8875 1700
rect 8925 1780 8965 1790
rect 8925 1700 8935 1780
rect 8955 1700 8965 1780
rect 8925 1690 8965 1700
rect 9015 1780 9055 1790
rect 9015 1700 9025 1780
rect 9045 1700 9055 1780
rect 9015 1690 9055 1700
rect 9105 1780 9145 1790
rect 9105 1700 9115 1780
rect 9135 1700 9145 1780
rect 9105 1690 9145 1700
rect 9195 1780 9235 1790
rect 9195 1700 9205 1780
rect 9225 1700 9235 1780
rect 9195 1690 9235 1700
rect 9285 1780 9325 1790
rect 9285 1700 9295 1780
rect 9315 1700 9325 1780
rect 9285 1690 9325 1700
rect 9375 1780 9415 1790
rect 9375 1700 9385 1780
rect 9405 1700 9415 1780
rect 9375 1690 9415 1700
rect 9465 1780 9505 1790
rect 9465 1700 9475 1780
rect 9495 1700 9505 1780
rect 9465 1690 9505 1700
rect 9555 1780 9595 1790
rect 9555 1700 9565 1780
rect 9585 1700 9595 1780
rect 9555 1690 9595 1700
rect 9645 1780 9685 1790
rect 9645 1700 9655 1780
rect 9675 1700 9685 1780
rect 9645 1690 9685 1700
rect 9735 1780 9775 1790
rect 9735 1700 9745 1780
rect 9765 1700 9775 1780
rect 9735 1690 9775 1700
rect 9825 1780 9865 1790
rect 9825 1700 9835 1780
rect 9855 1700 9865 1780
rect 9825 1690 9865 1700
rect 9915 1780 9955 1790
rect 9915 1700 9925 1780
rect 9945 1700 9955 1780
rect 9915 1690 9955 1700
rect 10005 1780 10045 1790
rect 10005 1700 10015 1780
rect 10035 1700 10045 1780
rect 10005 1690 10045 1700
rect 10095 1780 10135 1790
rect 10095 1700 10105 1780
rect 10125 1700 10135 1780
rect 10095 1690 10135 1700
rect 10185 1780 10225 1790
rect 10185 1700 10195 1780
rect 10215 1700 10225 1780
rect 10185 1690 10225 1700
rect 10275 1780 10315 1790
rect 10275 1700 10285 1780
rect 10305 1700 10315 1780
rect 10275 1690 10315 1700
rect 10365 1780 10405 1790
rect 10365 1700 10375 1780
rect 10395 1700 10405 1780
rect 10365 1690 10405 1700
rect 10455 1780 10495 1790
rect 10455 1700 10465 1780
rect 10485 1700 10495 1780
rect 10455 1690 10495 1700
rect 10545 1780 10585 1790
rect 10545 1700 10555 1780
rect 10575 1700 10585 1780
rect 10545 1690 10585 1700
rect 10635 1780 10675 1790
rect 10635 1700 10645 1780
rect 10665 1700 10675 1780
rect 10635 1690 10675 1700
rect 10725 1780 10765 1790
rect 10725 1700 10735 1780
rect 10755 1700 10765 1780
rect 10725 1690 10765 1700
rect 10815 1780 10855 1790
rect 10815 1700 10825 1780
rect 10845 1700 10855 1780
rect 10815 1690 10855 1700
rect 10905 1780 10945 1790
rect 10905 1700 10915 1780
rect 10935 1700 10945 1780
rect 10905 1690 10945 1700
rect 10995 1780 11035 1790
rect 10995 1700 11005 1780
rect 11025 1700 11035 1780
rect 10995 1690 11035 1700
rect 11085 1780 11125 1790
rect 11085 1700 11095 1780
rect 11115 1700 11125 1780
rect 11085 1690 11125 1700
rect 11175 1780 11215 1790
rect 11175 1700 11185 1780
rect 11205 1700 11215 1780
rect 11175 1690 11215 1700
rect -350 140 -310 150
rect -350 60 -340 140
rect -320 60 -310 140
rect -350 50 -310 60
rect -260 140 -220 150
rect -260 60 -250 140
rect -230 60 -220 140
rect -260 50 -220 60
rect -170 140 -130 150
rect -170 60 -160 140
rect -140 60 -130 140
rect -170 50 -130 60
rect -80 140 -40 150
rect -80 60 -70 140
rect -50 60 -40 140
rect -80 50 -40 60
rect 10 140 50 150
rect 10 60 20 140
rect 40 60 50 140
rect 10 50 50 60
rect 100 140 140 150
rect 100 60 110 140
rect 130 60 140 140
rect 100 50 140 60
rect 190 140 230 150
rect 190 60 200 140
rect 220 60 230 140
rect 190 50 230 60
rect 280 140 320 150
rect 280 60 290 140
rect 310 60 320 140
rect 280 50 320 60
rect 370 140 410 150
rect 370 60 380 140
rect 400 60 410 140
rect 370 50 410 60
rect 460 140 500 150
rect 460 60 470 140
rect 490 60 500 140
rect 460 50 500 60
rect 550 140 590 150
rect 550 60 560 140
rect 580 60 590 140
rect 550 50 590 60
rect 640 140 680 150
rect 640 60 650 140
rect 670 60 680 140
rect 640 50 680 60
rect 730 140 770 150
rect 730 60 740 140
rect 760 60 770 140
rect 730 50 770 60
rect 820 140 860 150
rect 820 60 830 140
rect 850 60 860 140
rect 820 50 860 60
rect 910 140 950 150
rect 910 60 920 140
rect 940 60 950 140
rect 910 50 950 60
rect 1000 140 1040 150
rect 1000 60 1010 140
rect 1030 60 1040 140
rect 1000 50 1040 60
rect 1090 140 1130 150
rect 1090 60 1100 140
rect 1120 60 1130 140
rect 1090 50 1130 60
rect 1180 140 1220 150
rect 1180 60 1190 140
rect 1210 60 1220 140
rect 1180 50 1220 60
rect 1270 140 1310 150
rect 1270 60 1280 140
rect 1300 60 1310 140
rect 1270 50 1310 60
rect 1360 140 1400 150
rect 1360 60 1370 140
rect 1390 60 1400 140
rect 1360 50 1400 60
rect 1450 140 1490 150
rect 1450 60 1460 140
rect 1480 60 1490 140
rect 1450 50 1490 60
rect 1540 140 1580 150
rect 1540 60 1550 140
rect 1570 60 1580 140
rect 1540 50 1580 60
rect 1630 140 1670 150
rect 1630 60 1640 140
rect 1660 60 1670 140
rect 1630 50 1670 60
rect 1720 140 1760 150
rect 1720 60 1730 140
rect 1750 60 1760 140
rect 1720 50 1760 60
rect 1810 140 1850 150
rect 1810 60 1820 140
rect 1840 60 1850 140
rect 1810 50 1850 60
rect 1900 140 1940 150
rect 1900 60 1910 140
rect 1930 60 1940 140
rect 1900 50 1940 60
rect 1990 140 2030 150
rect 1990 60 2000 140
rect 2020 60 2030 140
rect 1990 50 2030 60
rect 2080 140 2120 150
rect 2080 60 2090 140
rect 2110 60 2120 140
rect 2080 50 2120 60
rect 2170 140 2210 150
rect 2170 60 2180 140
rect 2200 60 2210 140
rect 2170 50 2210 60
rect 2260 140 2300 150
rect 2260 60 2270 140
rect 2290 60 2300 140
rect 2260 50 2300 60
rect 2350 140 2390 150
rect 2350 60 2360 140
rect 2380 60 2390 140
rect 2350 50 2390 60
rect 2440 140 2480 150
rect 2440 60 2450 140
rect 2470 60 2480 140
rect 2440 50 2480 60
rect 2530 140 2570 150
rect 2530 60 2540 140
rect 2560 60 2570 140
rect 2530 50 2570 60
rect 2620 140 2660 150
rect 2620 60 2630 140
rect 2650 60 2660 140
rect 2620 50 2660 60
rect 2710 140 2750 150
rect 2710 60 2720 140
rect 2740 60 2750 140
rect 2710 50 2750 60
rect 2800 140 2840 150
rect 2800 60 2810 140
rect 2830 60 2840 140
rect 2800 50 2840 60
rect 2890 140 2930 150
rect 2890 60 2900 140
rect 2920 60 2930 140
rect 2890 50 2930 60
rect 2980 140 3020 150
rect 2980 60 2990 140
rect 3010 60 3020 140
rect 2980 50 3020 60
rect 3070 140 3110 150
rect 3070 60 3080 140
rect 3100 60 3110 140
rect 3070 50 3110 60
rect 3160 140 3200 150
rect 3160 60 3170 140
rect 3190 60 3200 140
rect 3160 50 3200 60
rect 3250 140 3290 150
rect 3250 60 3260 140
rect 3280 60 3290 140
rect 3250 50 3290 60
rect 3340 140 3380 150
rect 3340 60 3350 140
rect 3370 60 3380 140
rect 3340 50 3380 60
rect 3430 140 3470 150
rect 3430 60 3440 140
rect 3460 60 3470 140
rect 3430 50 3470 60
rect 3520 140 3560 150
rect 3520 60 3530 140
rect 3550 60 3560 140
rect 3520 50 3560 60
rect 3610 140 3650 150
rect 3610 60 3620 140
rect 3640 60 3650 140
rect 3610 50 3650 60
rect 3700 140 3740 150
rect 3700 60 3710 140
rect 3730 60 3740 140
rect 3700 50 3740 60
rect 3790 140 3830 150
rect 3790 60 3800 140
rect 3820 60 3830 140
rect 3790 50 3830 60
rect 3880 140 3920 150
rect 3880 60 3890 140
rect 3910 60 3920 140
rect 3880 50 3920 60
rect 3970 140 4010 150
rect 3970 60 3980 140
rect 4000 60 4010 140
rect 3970 50 4010 60
rect 4060 140 4100 150
rect 4060 60 4070 140
rect 4090 60 4100 140
rect 4060 50 4100 60
rect 4150 140 4190 150
rect 4150 60 4160 140
rect 4180 60 4190 140
rect 4150 50 4190 60
rect 4240 140 4280 150
rect 4240 60 4250 140
rect 4270 60 4280 140
rect 4240 50 4280 60
rect 4330 140 4370 150
rect 4330 60 4340 140
rect 4360 60 4370 140
rect 4330 50 4370 60
rect 4420 140 4460 150
rect 4420 60 4430 140
rect 4450 60 4460 140
rect 4420 50 4460 60
rect 4510 140 4550 150
rect 4510 60 4520 140
rect 4540 60 4550 140
rect 4510 50 4550 60
rect 4600 140 4640 150
rect 4600 60 4610 140
rect 4630 60 4640 140
rect 4600 50 4640 60
rect 4690 140 4730 150
rect 4690 60 4700 140
rect 4720 60 4730 140
rect 4690 50 4730 60
rect 4780 140 4820 150
rect 4780 60 4790 140
rect 4810 60 4820 140
rect 4780 50 4820 60
rect 4870 140 4910 150
rect 4870 60 4880 140
rect 4900 60 4910 140
rect 4870 50 4910 60
rect 4960 140 5000 150
rect 4960 60 4970 140
rect 4990 60 5000 140
rect 4960 50 5000 60
rect 5050 140 5090 150
rect 5050 60 5060 140
rect 5080 60 5090 140
rect 5050 50 5090 60
rect 5140 140 5180 150
rect 5140 60 5150 140
rect 5170 60 5180 140
rect 5140 50 5180 60
rect 5230 140 5270 150
rect 5230 60 5240 140
rect 5260 60 5270 140
rect 5230 50 5270 60
rect 5320 140 5360 150
rect 5320 60 5330 140
rect 5350 60 5360 140
rect 5320 50 5360 60
rect 5410 140 5450 150
rect 5410 60 5420 140
rect 5440 60 5450 140
rect 5410 50 5450 60
rect 5500 140 5540 150
rect 5500 60 5510 140
rect 5530 60 5540 140
rect 5500 50 5540 60
rect 5590 140 5630 150
rect 5590 60 5600 140
rect 5620 60 5630 140
rect 5590 50 5630 60
rect 5680 140 5720 150
rect 5680 60 5690 140
rect 5710 60 5720 140
rect 5680 50 5720 60
rect 5770 140 5810 150
rect 5770 60 5780 140
rect 5800 60 5810 140
rect 5770 50 5810 60
rect 5860 140 5900 150
rect 5860 60 5870 140
rect 5890 60 5900 140
rect 5860 50 5900 60
rect 5950 140 5990 150
rect 5950 60 5960 140
rect 5980 60 5990 140
rect 5950 50 5990 60
rect 6040 140 6080 150
rect 6040 60 6050 140
rect 6070 60 6080 140
rect 6040 50 6080 60
rect 6130 140 6170 150
rect 6130 60 6140 140
rect 6160 60 6170 140
rect 6130 50 6170 60
rect 6220 140 6260 150
rect 6220 60 6230 140
rect 6250 60 6260 140
rect 6220 50 6260 60
rect 6310 140 6350 150
rect 6310 60 6320 140
rect 6340 60 6350 140
rect 6310 50 6350 60
rect 6400 140 6440 150
rect 6400 60 6410 140
rect 6430 60 6440 140
rect 6400 50 6440 60
rect 6490 140 6530 150
rect 6490 60 6500 140
rect 6520 60 6530 140
rect 6490 50 6530 60
rect 6580 140 6620 150
rect 6580 60 6590 140
rect 6610 60 6620 140
rect 6580 50 6620 60
rect 6670 140 6710 150
rect 6670 60 6680 140
rect 6700 60 6710 140
rect 6670 50 6710 60
rect 6760 140 6800 150
rect 6760 60 6770 140
rect 6790 60 6800 140
rect 6760 50 6800 60
rect 6850 140 6890 150
rect 6850 60 6860 140
rect 6880 60 6890 140
rect 6850 50 6890 60
rect 6940 140 6980 150
rect 6940 60 6950 140
rect 6970 60 6980 140
rect 6940 50 6980 60
rect 7030 140 7070 150
rect 7030 60 7040 140
rect 7060 60 7070 140
rect 7030 50 7070 60
rect 7120 140 7160 150
rect 7120 60 7130 140
rect 7150 60 7160 140
rect 7120 50 7160 60
rect 7210 140 7250 150
rect 7210 60 7220 140
rect 7240 60 7250 140
rect 7210 50 7250 60
rect 7300 140 7340 150
rect 7300 60 7310 140
rect 7330 60 7340 140
rect 7300 50 7340 60
rect 7390 140 7430 150
rect 7390 60 7400 140
rect 7420 60 7430 140
rect 7390 50 7430 60
rect 7480 140 7520 150
rect 7480 60 7490 140
rect 7510 60 7520 140
rect 7480 50 7520 60
rect 7570 140 7610 150
rect 7570 60 7580 140
rect 7600 60 7610 140
rect 7570 50 7610 60
rect 7660 140 7700 150
rect 7660 60 7670 140
rect 7690 60 7700 140
rect 7660 50 7700 60
rect 7750 140 7795 150
rect 7750 60 7760 140
rect 7780 60 7795 140
rect 7750 50 7795 60
rect 7845 140 7885 150
rect 7845 60 7855 140
rect 7875 60 7885 140
rect 7845 50 7885 60
rect 7935 140 7975 150
rect 7935 60 7945 140
rect 7965 60 7975 140
rect 7935 50 7975 60
rect 8025 140 8065 150
rect 8025 60 8035 140
rect 8055 60 8065 140
rect 8025 50 8065 60
rect 8115 140 8155 150
rect 8115 60 8125 140
rect 8145 60 8155 140
rect 8115 50 8155 60
rect 8205 140 8245 150
rect 8205 60 8215 140
rect 8235 60 8245 140
rect 8205 50 8245 60
rect 8295 140 8335 150
rect 8295 60 8305 140
rect 8325 60 8335 140
rect 8295 50 8335 60
rect 8385 140 8425 150
rect 8385 60 8395 140
rect 8415 60 8425 140
rect 8385 50 8425 60
rect 8475 140 8515 150
rect 8475 60 8485 140
rect 8505 60 8515 140
rect 8475 50 8515 60
rect 8565 140 8605 150
rect 8565 60 8575 140
rect 8595 60 8605 140
rect 8565 50 8605 60
rect 8655 140 8695 150
rect 8655 60 8665 140
rect 8685 60 8695 140
rect 8655 50 8695 60
rect 8745 140 8785 150
rect 8745 60 8755 140
rect 8775 60 8785 140
rect 8745 50 8785 60
rect 8835 140 8875 150
rect 8835 60 8845 140
rect 8865 60 8875 140
rect 8835 50 8875 60
rect 8925 140 8965 150
rect 8925 60 8935 140
rect 8955 60 8965 140
rect 8925 50 8965 60
rect 9015 140 9055 150
rect 9015 60 9025 140
rect 9045 60 9055 140
rect 9015 50 9055 60
rect 9105 140 9145 150
rect 9105 60 9115 140
rect 9135 60 9145 140
rect 9105 50 9145 60
rect 9195 140 9235 150
rect 9195 60 9205 140
rect 9225 60 9235 140
rect 9195 50 9235 60
rect 9285 140 9325 150
rect 9285 60 9295 140
rect 9315 60 9325 140
rect 9285 50 9325 60
rect 9375 140 9415 150
rect 9375 60 9385 140
rect 9405 60 9415 140
rect 9375 50 9415 60
rect 9465 140 9505 150
rect 9465 60 9475 140
rect 9495 60 9505 140
rect 9465 50 9505 60
rect 9555 140 9595 150
rect 9555 60 9565 140
rect 9585 60 9595 140
rect 9555 50 9595 60
rect 9645 140 9685 150
rect 9645 60 9655 140
rect 9675 60 9685 140
rect 9645 50 9685 60
rect 9735 140 9775 150
rect 9735 60 9745 140
rect 9765 60 9775 140
rect 9735 50 9775 60
rect 9825 140 9865 150
rect 9825 60 9835 140
rect 9855 60 9865 140
rect 9825 50 9865 60
rect 9915 140 9955 150
rect 9915 60 9925 140
rect 9945 60 9955 140
rect 9915 50 9955 60
rect 10005 140 10045 150
rect 10005 60 10015 140
rect 10035 60 10045 140
rect 10005 50 10045 60
rect 10095 140 10135 150
rect 10095 60 10105 140
rect 10125 60 10135 140
rect 10095 50 10135 60
rect 10185 140 10225 150
rect 10185 60 10195 140
rect 10215 60 10225 140
rect 10185 50 10225 60
rect 10275 140 10315 150
rect 10275 60 10285 140
rect 10305 60 10315 140
rect 10275 50 10315 60
rect 10365 140 10405 150
rect 10365 60 10375 140
rect 10395 60 10405 140
rect 10365 50 10405 60
rect 10455 140 10495 150
rect 10455 60 10465 140
rect 10485 60 10495 140
rect 10455 50 10495 60
rect 10545 140 10585 150
rect 10545 60 10555 140
rect 10575 60 10585 140
rect 10545 50 10585 60
rect 10635 140 10675 150
rect 10635 60 10645 140
rect 10665 60 10675 140
rect 10635 50 10675 60
rect 10725 140 10765 150
rect 10725 60 10735 140
rect 10755 60 10765 140
rect 10725 50 10765 60
rect 10815 140 10855 150
rect 10815 60 10825 140
rect 10845 60 10855 140
rect 10815 50 10855 60
rect 10905 140 10945 150
rect 10905 60 10915 140
rect 10935 60 10945 140
rect 10905 50 10945 60
rect 10995 140 11035 150
rect 10995 60 11005 140
rect 11025 60 11035 140
rect 10995 50 11035 60
rect 11085 140 11125 150
rect 11085 60 11095 140
rect 11115 60 11125 140
rect 11085 50 11125 60
rect 11175 140 11215 150
rect 11175 60 11185 140
rect 11205 60 11215 140
rect 11175 50 11215 60
<< pdiff >>
rect -350 1080 -310 1090
rect -350 1000 -340 1080
rect -320 1000 -310 1080
rect -350 990 -310 1000
rect -260 1080 -220 1090
rect -260 1000 -250 1080
rect -230 1000 -220 1080
rect -260 990 -220 1000
rect -170 1080 -130 1090
rect -170 1000 -160 1080
rect -140 1000 -130 1080
rect -170 990 -130 1000
rect -80 1080 -40 1090
rect -80 1000 -70 1080
rect -50 1000 -40 1080
rect -80 990 -40 1000
rect 10 1080 50 1090
rect 10 1000 20 1080
rect 40 1000 50 1080
rect 10 990 50 1000
rect 100 1080 140 1090
rect 100 1000 110 1080
rect 130 1000 140 1080
rect 100 990 140 1000
rect 190 1080 230 1090
rect 190 1000 200 1080
rect 220 1000 230 1080
rect 190 990 230 1000
rect 280 1080 320 1090
rect 280 1000 290 1080
rect 310 1000 320 1080
rect 280 990 320 1000
rect 370 1080 410 1090
rect 370 1000 380 1080
rect 400 1000 410 1080
rect 370 990 410 1000
rect 460 1080 500 1090
rect 460 1000 470 1080
rect 490 1000 500 1080
rect 460 990 500 1000
rect 550 1080 590 1090
rect 550 1000 560 1080
rect 580 1000 590 1080
rect 550 990 590 1000
rect 640 1080 680 1090
rect 640 1000 650 1080
rect 670 1000 680 1080
rect 640 990 680 1000
rect 730 1080 770 1090
rect 730 1000 740 1080
rect 760 1000 770 1080
rect 730 990 770 1000
rect 820 1080 860 1090
rect 820 1000 830 1080
rect 850 1000 860 1080
rect 820 990 860 1000
rect 910 1080 950 1090
rect 910 1000 920 1080
rect 940 1000 950 1080
rect 910 990 950 1000
rect 1000 1080 1040 1090
rect 1000 1000 1010 1080
rect 1030 1000 1040 1080
rect 1000 990 1040 1000
rect 1090 1080 1130 1090
rect 1090 1000 1100 1080
rect 1120 1000 1130 1080
rect 1090 990 1130 1000
rect 1180 1080 1220 1090
rect 1180 1000 1190 1080
rect 1210 1000 1220 1080
rect 1180 990 1220 1000
rect 1270 1080 1310 1090
rect 1270 1000 1280 1080
rect 1300 1000 1310 1080
rect 1270 990 1310 1000
rect 1360 1080 1400 1090
rect 1360 1000 1370 1080
rect 1390 1000 1400 1080
rect 1360 990 1400 1000
rect 1450 1080 1490 1090
rect 1450 1000 1460 1080
rect 1480 1000 1490 1080
rect 1450 990 1490 1000
rect 1540 1080 1580 1090
rect 1540 1000 1550 1080
rect 1570 1000 1580 1080
rect 1540 990 1580 1000
rect 1630 1080 1670 1090
rect 1630 1000 1640 1080
rect 1660 1000 1670 1080
rect 1630 990 1670 1000
rect 1720 1080 1760 1090
rect 1720 1000 1730 1080
rect 1750 1000 1760 1080
rect 1720 990 1760 1000
rect 1810 1080 1850 1090
rect 1810 1000 1820 1080
rect 1840 1000 1850 1080
rect 1810 990 1850 1000
rect 1900 1080 1940 1090
rect 1900 1000 1910 1080
rect 1930 1000 1940 1080
rect 1900 990 1940 1000
rect 1990 1080 2030 1090
rect 1990 1000 2000 1080
rect 2020 1000 2030 1080
rect 1990 990 2030 1000
rect 2080 1080 2120 1090
rect 2080 1000 2090 1080
rect 2110 1000 2120 1080
rect 2080 990 2120 1000
rect 2170 1080 2210 1090
rect 2170 1000 2180 1080
rect 2200 1000 2210 1080
rect 2170 990 2210 1000
rect 2260 1080 2300 1090
rect 2260 1000 2270 1080
rect 2290 1000 2300 1080
rect 2260 990 2300 1000
rect 2350 1080 2390 1090
rect 2350 1000 2360 1080
rect 2380 1000 2390 1080
rect 2350 990 2390 1000
rect 2440 1080 2480 1090
rect 2440 1000 2450 1080
rect 2470 1000 2480 1080
rect 2440 990 2480 1000
rect 2530 1080 2570 1090
rect 2530 1000 2540 1080
rect 2560 1000 2570 1080
rect 2530 990 2570 1000
rect 2620 1080 2660 1090
rect 2620 1000 2630 1080
rect 2650 1000 2660 1080
rect 2620 990 2660 1000
rect 2710 1080 2750 1090
rect 2710 1000 2720 1080
rect 2740 1000 2750 1080
rect 2710 990 2750 1000
rect 2800 1080 2840 1090
rect 2800 1000 2810 1080
rect 2830 1000 2840 1080
rect 2800 990 2840 1000
rect 2890 1080 2930 1090
rect 2890 1000 2900 1080
rect 2920 1000 2930 1080
rect 2890 990 2930 1000
rect 2980 1080 3020 1090
rect 2980 1000 2990 1080
rect 3010 1000 3020 1080
rect 2980 990 3020 1000
rect 3070 1080 3115 1090
rect 3070 1000 3085 1080
rect 3105 1000 3115 1080
rect 3070 990 3115 1000
rect 3165 1080 3205 1090
rect 3165 1000 3175 1080
rect 3195 1000 3205 1080
rect 3165 990 3205 1000
rect 3255 1080 3295 1090
rect 3255 1000 3265 1080
rect 3285 1000 3295 1080
rect 3255 990 3295 1000
rect 3345 1080 3385 1090
rect 3345 1000 3355 1080
rect 3375 1000 3385 1080
rect 3345 990 3385 1000
rect 3435 1080 3475 1090
rect 3435 1000 3445 1080
rect 3465 1000 3475 1080
rect 3435 990 3475 1000
rect 3525 1080 3565 1090
rect 3525 1000 3535 1080
rect 3555 1000 3565 1080
rect 3525 990 3565 1000
rect 3615 1080 3655 1090
rect 3615 1000 3625 1080
rect 3645 1000 3655 1080
rect 3615 990 3655 1000
rect 3705 1080 3745 1090
rect 3705 1000 3715 1080
rect 3735 1000 3745 1080
rect 3705 990 3745 1000
rect 3795 1080 3835 1090
rect 3795 1000 3805 1080
rect 3825 1000 3835 1080
rect 3795 990 3835 1000
rect 3885 1080 3925 1090
rect 3885 1000 3895 1080
rect 3915 1000 3925 1080
rect 3885 990 3925 1000
rect 3975 1080 4015 1090
rect 3975 1000 3985 1080
rect 4005 1000 4015 1080
rect 3975 990 4015 1000
rect 4065 1080 4105 1090
rect 4065 1000 4075 1080
rect 4095 1000 4105 1080
rect 4065 990 4105 1000
rect 4155 1080 4195 1090
rect 4155 1000 4165 1080
rect 4185 1000 4195 1080
rect 4155 990 4195 1000
rect 4245 1080 4285 1090
rect 4245 1000 4255 1080
rect 4275 1000 4285 1080
rect 4245 990 4285 1000
rect 4335 1080 4375 1090
rect 4335 1000 4345 1080
rect 4365 1000 4375 1080
rect 4335 990 4375 1000
rect 4425 1080 4465 1090
rect 4425 1000 4435 1080
rect 4455 1000 4465 1080
rect 4425 990 4465 1000
rect 4515 1080 4555 1090
rect 4515 1000 4525 1080
rect 4545 1000 4555 1080
rect 4515 990 4555 1000
rect 4605 1080 4645 1090
rect 4605 1000 4615 1080
rect 4635 1000 4645 1080
rect 4605 990 4645 1000
rect 4695 1080 4735 1090
rect 4695 1000 4705 1080
rect 4725 1000 4735 1080
rect 4695 990 4735 1000
rect 4785 1080 4825 1090
rect 4785 1000 4795 1080
rect 4815 1000 4825 1080
rect 4785 990 4825 1000
rect 4875 1080 4915 1090
rect 4875 1000 4885 1080
rect 4905 1000 4915 1080
rect 4875 990 4915 1000
rect 4965 1080 5005 1090
rect 4965 1000 4975 1080
rect 4995 1000 5005 1080
rect 4965 990 5005 1000
rect 5055 1080 5095 1090
rect 5055 1000 5065 1080
rect 5085 1000 5095 1080
rect 5055 990 5095 1000
rect 5145 1080 5185 1090
rect 5145 1000 5155 1080
rect 5175 1000 5185 1080
rect 5145 990 5185 1000
rect 5235 1080 5275 1090
rect 5235 1000 5245 1080
rect 5265 1000 5275 1080
rect 5235 990 5275 1000
rect 5325 1080 5365 1090
rect 5325 1000 5335 1080
rect 5355 1000 5365 1080
rect 5325 990 5365 1000
rect 5415 1080 5455 1090
rect 5415 1000 5425 1080
rect 5445 1000 5455 1080
rect 5415 990 5455 1000
rect 5505 1080 5545 1090
rect 5505 1000 5515 1080
rect 5535 1000 5545 1080
rect 5505 990 5545 1000
rect 5595 1080 5635 1090
rect 5595 1000 5605 1080
rect 5625 1000 5635 1080
rect 5595 990 5635 1000
rect 5685 1080 5725 1090
rect 5685 1000 5695 1080
rect 5715 1000 5725 1080
rect 5685 990 5725 1000
rect 5775 1080 5815 1090
rect 5775 1000 5785 1080
rect 5805 1000 5815 1080
rect 5775 990 5815 1000
rect 5865 1080 5905 1090
rect 5865 1000 5875 1080
rect 5895 1000 5905 1080
rect 5865 990 5905 1000
rect 5955 1080 5995 1090
rect 5955 1000 5965 1080
rect 5985 1000 5995 1080
rect 5955 990 5995 1000
rect 6045 1080 6085 1090
rect 6045 1000 6055 1080
rect 6075 1000 6085 1080
rect 6045 990 6085 1000
rect 6135 1080 6175 1090
rect 6135 1000 6145 1080
rect 6165 1000 6175 1080
rect 6135 990 6175 1000
rect 6225 1080 6265 1090
rect 6225 1000 6235 1080
rect 6255 1000 6265 1080
rect 6225 990 6265 1000
rect 6315 1080 6355 1090
rect 6315 1000 6325 1080
rect 6345 1000 6355 1080
rect 6315 990 6355 1000
rect 6405 1080 6445 1090
rect 6405 1000 6415 1080
rect 6435 1000 6445 1080
rect 6405 990 6445 1000
rect 6495 1080 6535 1090
rect 6495 1000 6505 1080
rect 6525 1000 6535 1080
rect 6495 990 6535 1000
rect 6585 1080 6625 1090
rect 6585 1000 6595 1080
rect 6615 1000 6625 1080
rect 6585 990 6625 1000
rect 6675 1080 6715 1090
rect 6675 1000 6685 1080
rect 6705 1000 6715 1080
rect 6675 990 6715 1000
rect 6765 1080 6805 1090
rect 6765 1000 6775 1080
rect 6795 1000 6805 1080
rect 6765 990 6805 1000
rect 6855 1080 6895 1090
rect 6855 1000 6865 1080
rect 6885 1000 6895 1080
rect 6855 990 6895 1000
rect 6945 1080 6985 1090
rect 6945 1000 6955 1080
rect 6975 1000 6985 1080
rect 6945 990 6985 1000
rect 7035 1080 7075 1090
rect 7035 1000 7045 1080
rect 7065 1000 7075 1080
rect 7035 990 7075 1000
rect 7125 1080 7165 1090
rect 7125 1000 7135 1080
rect 7155 1000 7165 1080
rect 7125 990 7165 1000
rect 7215 1080 7255 1090
rect 7215 1000 7225 1080
rect 7245 1000 7255 1080
rect 7215 990 7255 1000
rect 7305 1080 7345 1090
rect 7305 1000 7315 1080
rect 7335 1000 7345 1080
rect 7305 990 7345 1000
rect 7395 1080 7435 1090
rect 7395 1000 7405 1080
rect 7425 1000 7435 1080
rect 7395 990 7435 1000
rect 7485 1080 7525 1090
rect 7485 1000 7495 1080
rect 7515 1000 7525 1080
rect 7485 990 7525 1000
rect 7575 1080 7615 1090
rect 7575 1000 7585 1080
rect 7605 1000 7615 1080
rect 7575 990 7615 1000
rect 7665 1080 7705 1090
rect 7665 1000 7675 1080
rect 7695 1000 7705 1080
rect 7665 990 7705 1000
rect 7755 1080 7795 1090
rect 7755 1000 7765 1080
rect 7785 1000 7795 1080
rect 7755 990 7795 1000
rect 7845 1080 7885 1090
rect 7845 1000 7855 1080
rect 7875 1000 7885 1080
rect 7845 990 7885 1000
rect 7935 1080 7975 1090
rect 7935 1000 7945 1080
rect 7965 1000 7975 1080
rect 7935 990 7975 1000
rect 8025 1080 8065 1090
rect 8025 1000 8035 1080
rect 8055 1000 8065 1080
rect 8025 990 8065 1000
rect 8115 1080 8155 1090
rect 8115 1000 8125 1080
rect 8145 1000 8155 1080
rect 8115 990 8155 1000
rect 8205 1080 8245 1090
rect 8205 1000 8215 1080
rect 8235 1000 8245 1080
rect 8205 990 8245 1000
rect 8295 1080 8335 1090
rect 8295 1000 8305 1080
rect 8325 1000 8335 1080
rect 8295 990 8335 1000
rect 8385 1080 8425 1090
rect 8385 1000 8395 1080
rect 8415 1000 8425 1080
rect 8385 990 8425 1000
rect 8475 1080 8515 1090
rect 8475 1000 8485 1080
rect 8505 1000 8515 1080
rect 8475 990 8515 1000
rect 8565 1080 8605 1090
rect 8565 1000 8575 1080
rect 8595 1000 8605 1080
rect 8565 990 8605 1000
rect 8655 1080 8695 1090
rect 8655 1000 8665 1080
rect 8685 1000 8695 1080
rect 8655 990 8695 1000
rect 8745 1080 8785 1090
rect 8745 1000 8755 1080
rect 8775 1000 8785 1080
rect 8745 990 8785 1000
rect 8835 1080 8875 1090
rect 8835 1000 8845 1080
rect 8865 1000 8875 1080
rect 8835 990 8875 1000
rect 8925 1080 8965 1090
rect 8925 1000 8935 1080
rect 8955 1000 8965 1080
rect 8925 990 8965 1000
rect 9015 1080 9055 1090
rect 9015 1000 9025 1080
rect 9045 1000 9055 1080
rect 9015 990 9055 1000
rect 9105 1080 9145 1090
rect 9105 1000 9115 1080
rect 9135 1000 9145 1080
rect 9105 990 9145 1000
rect 9195 1080 9235 1090
rect 9195 1000 9205 1080
rect 9225 1000 9235 1080
rect 9195 990 9235 1000
rect 9285 1080 9325 1090
rect 9285 1000 9295 1080
rect 9315 1000 9325 1080
rect 9285 990 9325 1000
rect 9375 1080 9415 1090
rect 9375 1000 9385 1080
rect 9405 1000 9415 1080
rect 9375 990 9415 1000
rect 9465 1080 9505 1090
rect 9465 1000 9475 1080
rect 9495 1000 9505 1080
rect 9465 990 9505 1000
rect 9555 1080 9595 1090
rect 9555 1000 9565 1080
rect 9585 1000 9595 1080
rect 9555 990 9595 1000
rect 9645 1080 9685 1090
rect 9645 1000 9655 1080
rect 9675 1000 9685 1080
rect 9645 990 9685 1000
rect 9735 1080 9775 1090
rect 9735 1000 9745 1080
rect 9765 1000 9775 1080
rect 9735 990 9775 1000
rect 9825 1080 9865 1090
rect 9825 1000 9835 1080
rect 9855 1000 9865 1080
rect 9825 990 9865 1000
rect 9915 1080 9955 1090
rect 9915 1000 9925 1080
rect 9945 1000 9955 1080
rect 9915 990 9955 1000
rect 10005 1080 10045 1090
rect 10005 1000 10015 1080
rect 10035 1000 10045 1080
rect 10005 990 10045 1000
rect 10095 1080 10135 1090
rect 10095 1000 10105 1080
rect 10125 1000 10135 1080
rect 10095 990 10135 1000
rect 10185 1080 10225 1090
rect 10185 1000 10195 1080
rect 10215 1000 10225 1080
rect 10185 990 10225 1000
rect 10275 1080 10315 1090
rect 10275 1000 10285 1080
rect 10305 1000 10315 1080
rect 10275 990 10315 1000
rect 10365 1080 10405 1090
rect 10365 1000 10375 1080
rect 10395 1000 10405 1080
rect 10365 990 10405 1000
rect 10455 1080 10495 1090
rect 10455 1000 10465 1080
rect 10485 1000 10495 1080
rect 10455 990 10495 1000
rect 10545 1080 10585 1090
rect 10545 1000 10555 1080
rect 10575 1000 10585 1080
rect 10545 990 10585 1000
rect 10635 1080 10675 1090
rect 10635 1000 10645 1080
rect 10665 1000 10675 1080
rect 10635 990 10675 1000
rect 10725 1080 10765 1090
rect 10725 1000 10735 1080
rect 10755 1000 10765 1080
rect 10725 990 10765 1000
rect 10815 1080 10855 1090
rect 10815 1000 10825 1080
rect 10845 1000 10855 1080
rect 10815 990 10855 1000
rect 10905 1080 10945 1090
rect 10905 1000 10915 1080
rect 10935 1000 10945 1080
rect 10905 990 10945 1000
rect 10995 1080 11035 1090
rect 10995 1000 11005 1080
rect 11025 1000 11035 1080
rect 10995 990 11035 1000
rect 11085 1080 11125 1090
rect 11085 1000 11095 1080
rect 11115 1000 11125 1080
rect 11085 990 11125 1000
rect 11175 1080 11215 1090
rect 11175 1000 11185 1080
rect 11205 1000 11215 1080
rect 11175 990 11215 1000
rect -350 840 -310 850
rect -350 760 -340 840
rect -320 760 -310 840
rect -350 750 -310 760
rect -260 840 -220 850
rect -260 760 -250 840
rect -230 760 -220 840
rect -260 750 -220 760
rect -170 840 -130 850
rect -170 760 -160 840
rect -140 760 -130 840
rect -170 750 -130 760
rect -80 840 -40 850
rect -80 760 -70 840
rect -50 760 -40 840
rect -80 750 -40 760
rect 10 840 50 850
rect 10 760 20 840
rect 40 760 50 840
rect 10 750 50 760
rect 100 840 140 850
rect 100 760 110 840
rect 130 760 140 840
rect 100 750 140 760
rect 190 840 230 850
rect 190 760 200 840
rect 220 760 230 840
rect 190 750 230 760
rect 280 840 320 850
rect 280 760 290 840
rect 310 760 320 840
rect 280 750 320 760
rect 370 840 410 850
rect 370 760 380 840
rect 400 760 410 840
rect 370 750 410 760
rect 460 840 500 850
rect 460 760 470 840
rect 490 760 500 840
rect 460 750 500 760
rect 550 840 590 850
rect 550 760 560 840
rect 580 760 590 840
rect 550 750 590 760
rect 640 840 680 850
rect 640 760 650 840
rect 670 760 680 840
rect 640 750 680 760
rect 730 840 770 850
rect 730 760 740 840
rect 760 760 770 840
rect 730 750 770 760
rect 820 840 860 850
rect 820 760 830 840
rect 850 760 860 840
rect 820 750 860 760
rect 910 840 950 850
rect 910 760 920 840
rect 940 760 950 840
rect 910 750 950 760
rect 1000 840 1040 850
rect 1000 760 1010 840
rect 1030 760 1040 840
rect 1000 750 1040 760
rect 1090 840 1130 850
rect 1090 760 1100 840
rect 1120 760 1130 840
rect 1090 750 1130 760
rect 1180 840 1220 850
rect 1180 760 1190 840
rect 1210 760 1220 840
rect 1180 750 1220 760
rect 1270 840 1310 850
rect 1270 760 1280 840
rect 1300 760 1310 840
rect 1270 750 1310 760
rect 1360 840 1400 850
rect 1360 760 1370 840
rect 1390 760 1400 840
rect 1360 750 1400 760
rect 1450 840 1490 850
rect 1450 760 1460 840
rect 1480 760 1490 840
rect 1450 750 1490 760
rect 1540 840 1580 850
rect 1540 760 1550 840
rect 1570 760 1580 840
rect 1540 750 1580 760
rect 1630 840 1670 850
rect 1630 760 1640 840
rect 1660 760 1670 840
rect 1630 750 1670 760
rect 1720 840 1760 850
rect 1720 760 1730 840
rect 1750 760 1760 840
rect 1720 750 1760 760
rect 1810 840 1850 850
rect 1810 760 1820 840
rect 1840 760 1850 840
rect 1810 750 1850 760
rect 1900 840 1940 850
rect 1900 760 1910 840
rect 1930 760 1940 840
rect 1900 750 1940 760
rect 1990 840 2030 850
rect 1990 760 2000 840
rect 2020 760 2030 840
rect 1990 750 2030 760
rect 2080 840 2120 850
rect 2080 760 2090 840
rect 2110 760 2120 840
rect 2080 750 2120 760
rect 2170 840 2210 850
rect 2170 760 2180 840
rect 2200 760 2210 840
rect 2170 750 2210 760
rect 2260 840 2300 850
rect 2260 760 2270 840
rect 2290 760 2300 840
rect 2260 750 2300 760
rect 2350 840 2390 850
rect 2350 760 2360 840
rect 2380 760 2390 840
rect 2350 750 2390 760
rect 2440 840 2480 850
rect 2440 760 2450 840
rect 2470 760 2480 840
rect 2440 750 2480 760
rect 2530 840 2570 850
rect 2530 760 2540 840
rect 2560 760 2570 840
rect 2530 750 2570 760
rect 2620 840 2660 850
rect 2620 760 2630 840
rect 2650 760 2660 840
rect 2620 750 2660 760
rect 2710 840 2750 850
rect 2710 760 2720 840
rect 2740 760 2750 840
rect 2710 750 2750 760
rect 2800 840 2840 850
rect 2800 760 2810 840
rect 2830 760 2840 840
rect 2800 750 2840 760
rect 2890 840 2930 850
rect 2890 760 2900 840
rect 2920 760 2930 840
rect 2890 750 2930 760
rect 2980 840 3020 850
rect 2980 760 2990 840
rect 3010 760 3020 840
rect 2980 750 3020 760
rect 3070 840 3110 850
rect 3070 760 3080 840
rect 3100 760 3110 840
rect 3070 750 3110 760
rect 3160 840 3200 850
rect 3160 760 3170 840
rect 3190 760 3200 840
rect 3160 750 3200 760
rect 3250 840 3290 850
rect 3250 760 3260 840
rect 3280 760 3290 840
rect 3250 750 3290 760
rect 3340 840 3380 850
rect 3340 760 3350 840
rect 3370 760 3380 840
rect 3340 750 3380 760
rect 3430 840 3470 850
rect 3430 760 3440 840
rect 3460 760 3470 840
rect 3430 750 3470 760
rect 3520 840 3560 850
rect 3520 760 3530 840
rect 3550 760 3560 840
rect 3520 750 3560 760
rect 3610 840 3650 850
rect 3610 760 3620 840
rect 3640 760 3650 840
rect 3610 750 3650 760
rect 3700 840 3740 850
rect 3700 760 3710 840
rect 3730 760 3740 840
rect 3700 750 3740 760
rect 3790 840 3830 850
rect 3790 760 3800 840
rect 3820 760 3830 840
rect 3790 750 3830 760
rect 3880 840 3920 850
rect 3880 760 3890 840
rect 3910 760 3920 840
rect 3880 750 3920 760
rect 3970 840 4010 850
rect 3970 760 3980 840
rect 4000 760 4010 840
rect 3970 750 4010 760
rect 4060 840 4100 850
rect 4060 760 4070 840
rect 4090 760 4100 840
rect 4060 750 4100 760
rect 4150 840 4190 850
rect 4150 760 4160 840
rect 4180 760 4190 840
rect 4150 750 4190 760
rect 4240 840 4280 850
rect 4240 760 4250 840
rect 4270 760 4280 840
rect 4240 750 4280 760
rect 4330 840 4370 850
rect 4330 760 4340 840
rect 4360 760 4370 840
rect 4330 750 4370 760
rect 4420 840 4460 850
rect 4420 760 4430 840
rect 4450 760 4460 840
rect 4420 750 4460 760
rect 4510 840 4550 850
rect 4510 760 4520 840
rect 4540 760 4550 840
rect 4510 750 4550 760
rect 4600 840 4640 850
rect 4600 760 4610 840
rect 4630 760 4640 840
rect 4600 750 4640 760
rect 4690 840 4730 850
rect 4690 760 4700 840
rect 4720 760 4730 840
rect 4690 750 4730 760
rect 4780 840 4820 850
rect 4780 760 4790 840
rect 4810 760 4820 840
rect 4780 750 4820 760
rect 4870 840 4910 850
rect 4870 760 4880 840
rect 4900 760 4910 840
rect 4870 750 4910 760
rect 4960 840 5000 850
rect 4960 760 4970 840
rect 4990 760 5000 840
rect 4960 750 5000 760
rect 5050 840 5090 850
rect 5050 760 5060 840
rect 5080 760 5090 840
rect 5050 750 5090 760
rect 5140 840 5180 850
rect 5140 760 5150 840
rect 5170 760 5180 840
rect 5140 750 5180 760
rect 5230 840 5270 850
rect 5230 760 5240 840
rect 5260 760 5270 840
rect 5230 750 5270 760
rect 5320 840 5360 850
rect 5320 760 5330 840
rect 5350 760 5360 840
rect 5320 750 5360 760
rect 5410 840 5450 850
rect 5410 760 5420 840
rect 5440 760 5450 840
rect 5410 750 5450 760
rect 5500 840 5540 850
rect 5500 760 5510 840
rect 5530 760 5540 840
rect 5500 750 5540 760
rect 5590 840 5630 850
rect 5590 760 5600 840
rect 5620 760 5630 840
rect 5590 750 5630 760
rect 5680 840 5720 850
rect 5680 760 5690 840
rect 5710 760 5720 840
rect 5680 750 5720 760
rect 5770 840 5810 850
rect 5770 760 5780 840
rect 5800 760 5810 840
rect 5770 750 5810 760
rect 5860 840 5900 850
rect 5860 760 5870 840
rect 5890 760 5900 840
rect 5860 750 5900 760
rect 5950 840 5990 850
rect 5950 760 5960 840
rect 5980 760 5990 840
rect 5950 750 5990 760
rect 6040 840 6080 850
rect 6040 760 6050 840
rect 6070 760 6080 840
rect 6040 750 6080 760
rect 6130 840 6170 850
rect 6130 760 6140 840
rect 6160 760 6170 840
rect 6130 750 6170 760
rect 6220 840 6260 850
rect 6220 760 6230 840
rect 6250 760 6260 840
rect 6220 750 6260 760
rect 6310 840 6350 850
rect 6310 760 6320 840
rect 6340 760 6350 840
rect 6310 750 6350 760
rect 6400 840 6440 850
rect 6400 760 6410 840
rect 6430 760 6440 840
rect 6400 750 6440 760
rect 6490 840 6530 850
rect 6490 760 6500 840
rect 6520 760 6530 840
rect 6490 750 6530 760
rect 6580 840 6620 850
rect 6580 760 6590 840
rect 6610 760 6620 840
rect 6580 750 6620 760
rect 6670 840 6710 850
rect 6670 760 6680 840
rect 6700 760 6710 840
rect 6670 750 6710 760
rect 6760 840 6800 850
rect 6760 760 6770 840
rect 6790 760 6800 840
rect 6760 750 6800 760
rect 6850 840 6890 850
rect 6850 760 6860 840
rect 6880 760 6890 840
rect 6850 750 6890 760
rect 6940 840 6980 850
rect 6940 760 6950 840
rect 6970 760 6980 840
rect 6940 750 6980 760
rect 7030 840 7070 850
rect 7030 760 7040 840
rect 7060 760 7070 840
rect 7030 750 7070 760
rect 7120 840 7160 850
rect 7120 760 7130 840
rect 7150 760 7160 840
rect 7120 750 7160 760
rect 7210 840 7250 850
rect 7210 760 7220 840
rect 7240 760 7250 840
rect 7210 750 7250 760
rect 7300 840 7340 850
rect 7300 760 7310 840
rect 7330 760 7340 840
rect 7300 750 7340 760
rect 7390 840 7430 850
rect 7390 760 7400 840
rect 7420 760 7430 840
rect 7390 750 7430 760
rect 7480 840 7520 850
rect 7480 760 7490 840
rect 7510 760 7520 840
rect 7480 750 7520 760
rect 7570 840 7610 850
rect 7570 760 7580 840
rect 7600 760 7610 840
rect 7570 750 7610 760
rect 7660 840 7700 850
rect 7660 760 7670 840
rect 7690 760 7700 840
rect 7660 750 7700 760
rect 7750 840 7795 850
rect 7750 760 7760 840
rect 7780 760 7795 840
rect 7750 750 7795 760
rect 7845 840 7885 850
rect 7845 760 7855 840
rect 7875 760 7885 840
rect 7845 750 7885 760
rect 7935 840 7975 850
rect 7935 760 7945 840
rect 7965 760 7975 840
rect 7935 750 7975 760
rect 8025 840 8065 850
rect 8025 760 8035 840
rect 8055 760 8065 840
rect 8025 750 8065 760
rect 8115 840 8155 850
rect 8115 760 8125 840
rect 8145 760 8155 840
rect 8115 750 8155 760
rect 8205 840 8245 850
rect 8205 760 8215 840
rect 8235 760 8245 840
rect 8205 750 8245 760
rect 8295 840 8335 850
rect 8295 760 8305 840
rect 8325 760 8335 840
rect 8295 750 8335 760
rect 8385 840 8425 850
rect 8385 760 8395 840
rect 8415 760 8425 840
rect 8385 750 8425 760
rect 8475 840 8515 850
rect 8475 760 8485 840
rect 8505 760 8515 840
rect 8475 750 8515 760
rect 8565 840 8605 850
rect 8565 760 8575 840
rect 8595 760 8605 840
rect 8565 750 8605 760
rect 8655 840 8695 850
rect 8655 760 8665 840
rect 8685 760 8695 840
rect 8655 750 8695 760
rect 8745 840 8785 850
rect 8745 760 8755 840
rect 8775 760 8785 840
rect 8745 750 8785 760
rect 8835 840 8875 850
rect 8835 760 8845 840
rect 8865 760 8875 840
rect 8835 750 8875 760
rect 8925 840 8965 850
rect 8925 760 8935 840
rect 8955 760 8965 840
rect 8925 750 8965 760
rect 9015 840 9055 850
rect 9015 760 9025 840
rect 9045 760 9055 840
rect 9015 750 9055 760
rect 9105 840 9145 850
rect 9105 760 9115 840
rect 9135 760 9145 840
rect 9105 750 9145 760
rect 9195 840 9235 850
rect 9195 760 9205 840
rect 9225 760 9235 840
rect 9195 750 9235 760
rect 9285 840 9325 850
rect 9285 760 9295 840
rect 9315 760 9325 840
rect 9285 750 9325 760
rect 9375 840 9415 850
rect 9375 760 9385 840
rect 9405 760 9415 840
rect 9375 750 9415 760
rect 9465 840 9505 850
rect 9465 760 9475 840
rect 9495 760 9505 840
rect 9465 750 9505 760
rect 9555 840 9595 850
rect 9555 760 9565 840
rect 9585 760 9595 840
rect 9555 750 9595 760
rect 9645 840 9685 850
rect 9645 760 9655 840
rect 9675 760 9685 840
rect 9645 750 9685 760
rect 9735 840 9775 850
rect 9735 760 9745 840
rect 9765 760 9775 840
rect 9735 750 9775 760
rect 9825 840 9865 850
rect 9825 760 9835 840
rect 9855 760 9865 840
rect 9825 750 9865 760
rect 9915 840 9955 850
rect 9915 760 9925 840
rect 9945 760 9955 840
rect 9915 750 9955 760
rect 10005 840 10045 850
rect 10005 760 10015 840
rect 10035 760 10045 840
rect 10005 750 10045 760
rect 10095 840 10135 850
rect 10095 760 10105 840
rect 10125 760 10135 840
rect 10095 750 10135 760
rect 10185 840 10225 850
rect 10185 760 10195 840
rect 10215 760 10225 840
rect 10185 750 10225 760
rect 10275 840 10315 850
rect 10275 760 10285 840
rect 10305 760 10315 840
rect 10275 750 10315 760
rect 10365 840 10405 850
rect 10365 760 10375 840
rect 10395 760 10405 840
rect 10365 750 10405 760
rect 10455 840 10495 850
rect 10455 760 10465 840
rect 10485 760 10495 840
rect 10455 750 10495 760
rect 10545 840 10585 850
rect 10545 760 10555 840
rect 10575 760 10585 840
rect 10545 750 10585 760
rect 10635 840 10675 850
rect 10635 760 10645 840
rect 10665 760 10675 840
rect 10635 750 10675 760
rect 10725 840 10765 850
rect 10725 760 10735 840
rect 10755 760 10765 840
rect 10725 750 10765 760
rect 10815 840 10855 850
rect 10815 760 10825 840
rect 10845 760 10855 840
rect 10815 750 10855 760
rect 10905 840 10945 850
rect 10905 760 10915 840
rect 10935 760 10945 840
rect 10905 750 10945 760
rect 10995 840 11035 850
rect 10995 760 11005 840
rect 11025 760 11035 840
rect 10995 750 11035 760
rect 11085 840 11125 850
rect 11085 760 11095 840
rect 11115 760 11125 840
rect 11085 750 11125 760
rect 11175 840 11215 850
rect 11175 760 11185 840
rect 11205 760 11215 840
rect 11175 750 11215 760
<< ndiffc >>
rect -340 1700 -320 1780
rect -250 1700 -230 1780
rect -160 1700 -140 1780
rect -70 1700 -50 1780
rect 20 1700 40 1780
rect 110 1700 130 1780
rect 200 1700 220 1780
rect 290 1700 310 1780
rect 380 1700 400 1780
rect 470 1700 490 1780
rect 560 1700 580 1780
rect 650 1700 670 1780
rect 740 1700 760 1780
rect 830 1700 850 1780
rect 920 1700 940 1780
rect 1010 1700 1030 1780
rect 1100 1700 1120 1780
rect 1190 1700 1210 1780
rect 1280 1700 1300 1780
rect 1370 1700 1390 1780
rect 1460 1700 1480 1780
rect 1550 1700 1570 1780
rect 1640 1700 1660 1780
rect 1730 1700 1750 1780
rect 1820 1700 1840 1780
rect 1910 1700 1930 1780
rect 2000 1700 2020 1780
rect 2090 1700 2110 1780
rect 2180 1700 2200 1780
rect 2270 1700 2290 1780
rect 2360 1700 2380 1780
rect 2450 1700 2470 1780
rect 2540 1700 2560 1780
rect 2630 1700 2650 1780
rect 2720 1700 2740 1780
rect 2810 1700 2830 1780
rect 2900 1700 2920 1780
rect 2990 1700 3010 1780
rect 3085 1700 3105 1780
rect 3175 1700 3195 1780
rect 3265 1700 3285 1780
rect 3355 1700 3375 1780
rect 3445 1700 3465 1780
rect 3535 1700 3555 1780
rect 3625 1700 3645 1780
rect 3715 1700 3735 1780
rect 3805 1700 3825 1780
rect 3895 1700 3915 1780
rect 3985 1700 4005 1780
rect 4075 1700 4095 1780
rect 4165 1700 4185 1780
rect 4255 1700 4275 1780
rect 4345 1700 4365 1780
rect 4435 1700 4455 1780
rect 4525 1700 4545 1780
rect 4615 1700 4635 1780
rect 4705 1700 4725 1780
rect 4795 1700 4815 1780
rect 4885 1700 4905 1780
rect 4975 1700 4995 1780
rect 5065 1700 5085 1780
rect 5155 1700 5175 1780
rect 5245 1700 5265 1780
rect 5335 1700 5355 1780
rect 5425 1700 5445 1780
rect 5515 1700 5535 1780
rect 5605 1700 5625 1780
rect 5695 1700 5715 1780
rect 5785 1700 5805 1780
rect 5875 1700 5895 1780
rect 5965 1700 5985 1780
rect 6055 1700 6075 1780
rect 6145 1700 6165 1780
rect 6235 1700 6255 1780
rect 6325 1700 6345 1780
rect 6415 1700 6435 1780
rect 6505 1700 6525 1780
rect 6595 1700 6615 1780
rect 6685 1700 6705 1780
rect 6775 1700 6795 1780
rect 6865 1700 6885 1780
rect 6955 1700 6975 1780
rect 7045 1700 7065 1780
rect 7135 1700 7155 1780
rect 7225 1700 7245 1780
rect 7315 1700 7335 1780
rect 7405 1700 7425 1780
rect 7495 1700 7515 1780
rect 7585 1700 7605 1780
rect 7675 1700 7695 1780
rect 7765 1700 7785 1780
rect 7855 1700 7875 1780
rect 7945 1700 7965 1780
rect 8035 1700 8055 1780
rect 8125 1700 8145 1780
rect 8215 1700 8235 1780
rect 8305 1700 8325 1780
rect 8395 1700 8415 1780
rect 8485 1700 8505 1780
rect 8575 1700 8595 1780
rect 8665 1700 8685 1780
rect 8755 1700 8775 1780
rect 8845 1700 8865 1780
rect 8935 1700 8955 1780
rect 9025 1700 9045 1780
rect 9115 1700 9135 1780
rect 9205 1700 9225 1780
rect 9295 1700 9315 1780
rect 9385 1700 9405 1780
rect 9475 1700 9495 1780
rect 9565 1700 9585 1780
rect 9655 1700 9675 1780
rect 9745 1700 9765 1780
rect 9835 1700 9855 1780
rect 9925 1700 9945 1780
rect 10015 1700 10035 1780
rect 10105 1700 10125 1780
rect 10195 1700 10215 1780
rect 10285 1700 10305 1780
rect 10375 1700 10395 1780
rect 10465 1700 10485 1780
rect 10555 1700 10575 1780
rect 10645 1700 10665 1780
rect 10735 1700 10755 1780
rect 10825 1700 10845 1780
rect 10915 1700 10935 1780
rect 11005 1700 11025 1780
rect 11095 1700 11115 1780
rect 11185 1700 11205 1780
rect -340 60 -320 140
rect -250 60 -230 140
rect -160 60 -140 140
rect -70 60 -50 140
rect 20 60 40 140
rect 110 60 130 140
rect 200 60 220 140
rect 290 60 310 140
rect 380 60 400 140
rect 470 60 490 140
rect 560 60 580 140
rect 650 60 670 140
rect 740 60 760 140
rect 830 60 850 140
rect 920 60 940 140
rect 1010 60 1030 140
rect 1100 60 1120 140
rect 1190 60 1210 140
rect 1280 60 1300 140
rect 1370 60 1390 140
rect 1460 60 1480 140
rect 1550 60 1570 140
rect 1640 60 1660 140
rect 1730 60 1750 140
rect 1820 60 1840 140
rect 1910 60 1930 140
rect 2000 60 2020 140
rect 2090 60 2110 140
rect 2180 60 2200 140
rect 2270 60 2290 140
rect 2360 60 2380 140
rect 2450 60 2470 140
rect 2540 60 2560 140
rect 2630 60 2650 140
rect 2720 60 2740 140
rect 2810 60 2830 140
rect 2900 60 2920 140
rect 2990 60 3010 140
rect 3080 60 3100 140
rect 3170 60 3190 140
rect 3260 60 3280 140
rect 3350 60 3370 140
rect 3440 60 3460 140
rect 3530 60 3550 140
rect 3620 60 3640 140
rect 3710 60 3730 140
rect 3800 60 3820 140
rect 3890 60 3910 140
rect 3980 60 4000 140
rect 4070 60 4090 140
rect 4160 60 4180 140
rect 4250 60 4270 140
rect 4340 60 4360 140
rect 4430 60 4450 140
rect 4520 60 4540 140
rect 4610 60 4630 140
rect 4700 60 4720 140
rect 4790 60 4810 140
rect 4880 60 4900 140
rect 4970 60 4990 140
rect 5060 60 5080 140
rect 5150 60 5170 140
rect 5240 60 5260 140
rect 5330 60 5350 140
rect 5420 60 5440 140
rect 5510 60 5530 140
rect 5600 60 5620 140
rect 5690 60 5710 140
rect 5780 60 5800 140
rect 5870 60 5890 140
rect 5960 60 5980 140
rect 6050 60 6070 140
rect 6140 60 6160 140
rect 6230 60 6250 140
rect 6320 60 6340 140
rect 6410 60 6430 140
rect 6500 60 6520 140
rect 6590 60 6610 140
rect 6680 60 6700 140
rect 6770 60 6790 140
rect 6860 60 6880 140
rect 6950 60 6970 140
rect 7040 60 7060 140
rect 7130 60 7150 140
rect 7220 60 7240 140
rect 7310 60 7330 140
rect 7400 60 7420 140
rect 7490 60 7510 140
rect 7580 60 7600 140
rect 7670 60 7690 140
rect 7760 60 7780 140
rect 7855 60 7875 140
rect 7945 60 7965 140
rect 8035 60 8055 140
rect 8125 60 8145 140
rect 8215 60 8235 140
rect 8305 60 8325 140
rect 8395 60 8415 140
rect 8485 60 8505 140
rect 8575 60 8595 140
rect 8665 60 8685 140
rect 8755 60 8775 140
rect 8845 60 8865 140
rect 8935 60 8955 140
rect 9025 60 9045 140
rect 9115 60 9135 140
rect 9205 60 9225 140
rect 9295 60 9315 140
rect 9385 60 9405 140
rect 9475 60 9495 140
rect 9565 60 9585 140
rect 9655 60 9675 140
rect 9745 60 9765 140
rect 9835 60 9855 140
rect 9925 60 9945 140
rect 10015 60 10035 140
rect 10105 60 10125 140
rect 10195 60 10215 140
rect 10285 60 10305 140
rect 10375 60 10395 140
rect 10465 60 10485 140
rect 10555 60 10575 140
rect 10645 60 10665 140
rect 10735 60 10755 140
rect 10825 60 10845 140
rect 10915 60 10935 140
rect 11005 60 11025 140
rect 11095 60 11115 140
rect 11185 60 11205 140
<< pdiffc >>
rect -340 1000 -320 1080
rect -250 1000 -230 1080
rect -160 1000 -140 1080
rect -70 1000 -50 1080
rect 20 1000 40 1080
rect 110 1000 130 1080
rect 200 1000 220 1080
rect 290 1000 310 1080
rect 380 1000 400 1080
rect 470 1000 490 1080
rect 560 1000 580 1080
rect 650 1000 670 1080
rect 740 1000 760 1080
rect 830 1000 850 1080
rect 920 1000 940 1080
rect 1010 1000 1030 1080
rect 1100 1000 1120 1080
rect 1190 1000 1210 1080
rect 1280 1000 1300 1080
rect 1370 1000 1390 1080
rect 1460 1000 1480 1080
rect 1550 1000 1570 1080
rect 1640 1000 1660 1080
rect 1730 1000 1750 1080
rect 1820 1000 1840 1080
rect 1910 1000 1930 1080
rect 2000 1000 2020 1080
rect 2090 1000 2110 1080
rect 2180 1000 2200 1080
rect 2270 1000 2290 1080
rect 2360 1000 2380 1080
rect 2450 1000 2470 1080
rect 2540 1000 2560 1080
rect 2630 1000 2650 1080
rect 2720 1000 2740 1080
rect 2810 1000 2830 1080
rect 2900 1000 2920 1080
rect 2990 1000 3010 1080
rect 3085 1000 3105 1080
rect 3175 1000 3195 1080
rect 3265 1000 3285 1080
rect 3355 1000 3375 1080
rect 3445 1000 3465 1080
rect 3535 1000 3555 1080
rect 3625 1000 3645 1080
rect 3715 1000 3735 1080
rect 3805 1000 3825 1080
rect 3895 1000 3915 1080
rect 3985 1000 4005 1080
rect 4075 1000 4095 1080
rect 4165 1000 4185 1080
rect 4255 1000 4275 1080
rect 4345 1000 4365 1080
rect 4435 1000 4455 1080
rect 4525 1000 4545 1080
rect 4615 1000 4635 1080
rect 4705 1000 4725 1080
rect 4795 1000 4815 1080
rect 4885 1000 4905 1080
rect 4975 1000 4995 1080
rect 5065 1000 5085 1080
rect 5155 1000 5175 1080
rect 5245 1000 5265 1080
rect 5335 1000 5355 1080
rect 5425 1000 5445 1080
rect 5515 1000 5535 1080
rect 5605 1000 5625 1080
rect 5695 1000 5715 1080
rect 5785 1000 5805 1080
rect 5875 1000 5895 1080
rect 5965 1000 5985 1080
rect 6055 1000 6075 1080
rect 6145 1000 6165 1080
rect 6235 1000 6255 1080
rect 6325 1000 6345 1080
rect 6415 1000 6435 1080
rect 6505 1000 6525 1080
rect 6595 1000 6615 1080
rect 6685 1000 6705 1080
rect 6775 1000 6795 1080
rect 6865 1000 6885 1080
rect 6955 1000 6975 1080
rect 7045 1000 7065 1080
rect 7135 1000 7155 1080
rect 7225 1000 7245 1080
rect 7315 1000 7335 1080
rect 7405 1000 7425 1080
rect 7495 1000 7515 1080
rect 7585 1000 7605 1080
rect 7675 1000 7695 1080
rect 7765 1000 7785 1080
rect 7855 1000 7875 1080
rect 7945 1000 7965 1080
rect 8035 1000 8055 1080
rect 8125 1000 8145 1080
rect 8215 1000 8235 1080
rect 8305 1000 8325 1080
rect 8395 1000 8415 1080
rect 8485 1000 8505 1080
rect 8575 1000 8595 1080
rect 8665 1000 8685 1080
rect 8755 1000 8775 1080
rect 8845 1000 8865 1080
rect 8935 1000 8955 1080
rect 9025 1000 9045 1080
rect 9115 1000 9135 1080
rect 9205 1000 9225 1080
rect 9295 1000 9315 1080
rect 9385 1000 9405 1080
rect 9475 1000 9495 1080
rect 9565 1000 9585 1080
rect 9655 1000 9675 1080
rect 9745 1000 9765 1080
rect 9835 1000 9855 1080
rect 9925 1000 9945 1080
rect 10015 1000 10035 1080
rect 10105 1000 10125 1080
rect 10195 1000 10215 1080
rect 10285 1000 10305 1080
rect 10375 1000 10395 1080
rect 10465 1000 10485 1080
rect 10555 1000 10575 1080
rect 10645 1000 10665 1080
rect 10735 1000 10755 1080
rect 10825 1000 10845 1080
rect 10915 1000 10935 1080
rect 11005 1000 11025 1080
rect 11095 1000 11115 1080
rect 11185 1000 11205 1080
rect -340 760 -320 840
rect -250 760 -230 840
rect -160 760 -140 840
rect -70 760 -50 840
rect 20 760 40 840
rect 110 760 130 840
rect 200 760 220 840
rect 290 760 310 840
rect 380 760 400 840
rect 470 760 490 840
rect 560 760 580 840
rect 650 760 670 840
rect 740 760 760 840
rect 830 760 850 840
rect 920 760 940 840
rect 1010 760 1030 840
rect 1100 760 1120 840
rect 1190 760 1210 840
rect 1280 760 1300 840
rect 1370 760 1390 840
rect 1460 760 1480 840
rect 1550 760 1570 840
rect 1640 760 1660 840
rect 1730 760 1750 840
rect 1820 760 1840 840
rect 1910 760 1930 840
rect 2000 760 2020 840
rect 2090 760 2110 840
rect 2180 760 2200 840
rect 2270 760 2290 840
rect 2360 760 2380 840
rect 2450 760 2470 840
rect 2540 760 2560 840
rect 2630 760 2650 840
rect 2720 760 2740 840
rect 2810 760 2830 840
rect 2900 760 2920 840
rect 2990 760 3010 840
rect 3080 760 3100 840
rect 3170 760 3190 840
rect 3260 760 3280 840
rect 3350 760 3370 840
rect 3440 760 3460 840
rect 3530 760 3550 840
rect 3620 760 3640 840
rect 3710 760 3730 840
rect 3800 760 3820 840
rect 3890 760 3910 840
rect 3980 760 4000 840
rect 4070 760 4090 840
rect 4160 760 4180 840
rect 4250 760 4270 840
rect 4340 760 4360 840
rect 4430 760 4450 840
rect 4520 760 4540 840
rect 4610 760 4630 840
rect 4700 760 4720 840
rect 4790 760 4810 840
rect 4880 760 4900 840
rect 4970 760 4990 840
rect 5060 760 5080 840
rect 5150 760 5170 840
rect 5240 760 5260 840
rect 5330 760 5350 840
rect 5420 760 5440 840
rect 5510 760 5530 840
rect 5600 760 5620 840
rect 5690 760 5710 840
rect 5780 760 5800 840
rect 5870 760 5890 840
rect 5960 760 5980 840
rect 6050 760 6070 840
rect 6140 760 6160 840
rect 6230 760 6250 840
rect 6320 760 6340 840
rect 6410 760 6430 840
rect 6500 760 6520 840
rect 6590 760 6610 840
rect 6680 760 6700 840
rect 6770 760 6790 840
rect 6860 760 6880 840
rect 6950 760 6970 840
rect 7040 760 7060 840
rect 7130 760 7150 840
rect 7220 760 7240 840
rect 7310 760 7330 840
rect 7400 760 7420 840
rect 7490 760 7510 840
rect 7580 760 7600 840
rect 7670 760 7690 840
rect 7760 760 7780 840
rect 7855 760 7875 840
rect 7945 760 7965 840
rect 8035 760 8055 840
rect 8125 760 8145 840
rect 8215 760 8235 840
rect 8305 760 8325 840
rect 8395 760 8415 840
rect 8485 760 8505 840
rect 8575 760 8595 840
rect 8665 760 8685 840
rect 8755 760 8775 840
rect 8845 760 8865 840
rect 8935 760 8955 840
rect 9025 760 9045 840
rect 9115 760 9135 840
rect 9205 760 9225 840
rect 9295 760 9315 840
rect 9385 760 9405 840
rect 9475 760 9495 840
rect 9565 760 9585 840
rect 9655 760 9675 840
rect 9745 760 9765 840
rect 9835 760 9855 840
rect 9925 760 9945 840
rect 10015 760 10035 840
rect 10105 760 10125 840
rect 10195 760 10215 840
rect 10285 760 10305 840
rect 10375 760 10395 840
rect 10465 760 10485 840
rect 10555 760 10575 840
rect 10645 760 10665 840
rect 10735 760 10755 840
rect 10825 760 10845 840
rect 10915 760 10935 840
rect 11005 760 11025 840
rect 11095 760 11115 840
rect 11185 760 11205 840
<< psubdiff >>
rect -485 1820 -295 1840
rect -275 1820 -205 1840
rect -185 1820 -115 1840
rect -95 1820 -25 1840
rect -5 1820 65 1840
rect 85 1820 155 1840
rect 175 1820 245 1840
rect 265 1820 335 1840
rect 355 1820 425 1840
rect 445 1820 515 1840
rect 535 1820 605 1840
rect 625 1820 695 1840
rect 715 1820 785 1840
rect 805 1820 875 1840
rect 895 1820 965 1840
rect 985 1820 1055 1840
rect 1075 1820 1145 1840
rect 1165 1820 1235 1840
rect 1255 1820 1325 1840
rect 1345 1820 1415 1840
rect 1435 1820 1505 1840
rect 1525 1820 1595 1840
rect 1615 1820 1685 1840
rect 1705 1820 1775 1840
rect 1795 1820 1865 1840
rect 1885 1820 1955 1840
rect 1975 1820 2045 1840
rect 2065 1820 2135 1840
rect 2155 1820 2225 1840
rect 2245 1820 2315 1840
rect 2335 1820 2405 1840
rect 2425 1820 2495 1840
rect 2515 1820 2585 1840
rect 2605 1820 2675 1840
rect 2695 1820 2765 1840
rect 2785 1820 2855 1840
rect 2875 1820 2945 1840
rect 2965 1820 3035 1840
rect 3055 1820 3130 1840
rect 3150 1820 3220 1840
rect 3240 1820 3310 1840
rect 3330 1820 3400 1840
rect 3420 1820 3490 1840
rect 3510 1820 3580 1840
rect 3600 1820 3670 1840
rect 3690 1820 3760 1840
rect 3780 1820 3850 1840
rect 3870 1820 3940 1840
rect 3960 1820 4030 1840
rect 4050 1820 4120 1840
rect 4140 1820 4210 1840
rect 4230 1820 4300 1840
rect 4320 1820 4390 1840
rect 4410 1820 4480 1840
rect 4500 1820 4570 1840
rect 4590 1820 4660 1840
rect 4680 1820 4750 1840
rect 4770 1820 4840 1840
rect 4860 1820 4930 1840
rect 4950 1820 5020 1840
rect 5040 1820 5110 1840
rect 5130 1820 5200 1840
rect 5220 1820 5290 1840
rect 5310 1820 5380 1840
rect 5400 1820 5470 1840
rect 5490 1820 5560 1840
rect 5580 1820 5650 1840
rect 5670 1820 5740 1840
rect 5760 1820 5830 1840
rect 5850 1820 5920 1840
rect 5940 1820 6010 1840
rect 6030 1820 6100 1840
rect 6120 1820 6190 1840
rect 6210 1820 6280 1840
rect 6300 1820 6370 1840
rect 6390 1820 6460 1840
rect 6480 1820 6550 1840
rect 6570 1820 6640 1840
rect 6660 1820 6730 1840
rect 6750 1820 6820 1840
rect 6840 1820 6910 1840
rect 6930 1820 7000 1840
rect 7020 1820 7090 1840
rect 7110 1820 7180 1840
rect 7200 1820 7270 1840
rect 7290 1820 7360 1840
rect 7380 1820 7450 1840
rect 7470 1820 7540 1840
rect 7560 1820 7630 1840
rect 7650 1820 7720 1840
rect 7740 1820 7810 1840
rect 7830 1820 7900 1840
rect 7920 1820 7990 1840
rect 8010 1820 8080 1840
rect 8100 1820 8170 1840
rect 8190 1820 8260 1840
rect 8280 1820 8350 1840
rect 8370 1820 8440 1840
rect 8460 1820 8530 1840
rect 8550 1820 8620 1840
rect 8640 1820 8710 1840
rect 8730 1820 8800 1840
rect 8820 1820 8890 1840
rect 8910 1820 8980 1840
rect 9000 1820 9070 1840
rect 9090 1820 9160 1840
rect 9180 1820 9250 1840
rect 9270 1820 9340 1840
rect 9360 1820 9430 1840
rect 9450 1820 9520 1840
rect 9540 1820 9610 1840
rect 9630 1820 9700 1840
rect 9720 1820 9790 1840
rect 9810 1820 9880 1840
rect 9900 1820 9970 1840
rect 9990 1820 10060 1840
rect 10080 1820 10150 1840
rect 10170 1820 10240 1840
rect 10260 1820 10330 1840
rect 10350 1820 10420 1840
rect 10440 1820 10510 1840
rect 10530 1820 10600 1840
rect 10620 1820 10690 1840
rect 10710 1820 10780 1840
rect 10800 1820 10870 1840
rect 10890 1820 10960 1840
rect 10980 1820 11050 1840
rect 11070 1820 11140 1840
rect 11160 1820 11350 1840
rect -475 1620 -455 1820
rect 11320 1620 11340 1820
rect -475 1600 -295 1620
rect -275 1600 -205 1620
rect -185 1600 -115 1620
rect -95 1600 -25 1620
rect -5 1600 65 1620
rect 85 1600 155 1620
rect 175 1600 245 1620
rect 265 1600 335 1620
rect 355 1600 425 1620
rect 445 1600 515 1620
rect 535 1600 605 1620
rect 625 1600 695 1620
rect 715 1600 785 1620
rect 805 1600 875 1620
rect 895 1600 965 1620
rect 985 1600 1055 1620
rect 1075 1600 1145 1620
rect 1165 1600 1235 1620
rect 1255 1600 1325 1620
rect 1345 1600 1415 1620
rect 1435 1600 1505 1620
rect 1525 1600 1595 1620
rect 1615 1600 1685 1620
rect 1705 1600 1775 1620
rect 1795 1600 1865 1620
rect 1885 1600 1955 1620
rect 1975 1600 2045 1620
rect 2065 1600 2135 1620
rect 2155 1600 2225 1620
rect 2245 1600 2315 1620
rect 2335 1600 2405 1620
rect 2425 1600 2495 1620
rect 2515 1600 2585 1620
rect 2605 1600 2675 1620
rect 2695 1600 2765 1620
rect 2785 1600 2855 1620
rect 2875 1600 2945 1620
rect 2965 1600 3035 1620
rect 3055 1600 3130 1620
rect 3150 1600 3220 1620
rect 3240 1600 3310 1620
rect 3330 1600 3400 1620
rect 3420 1600 3490 1620
rect 3510 1600 3580 1620
rect 3600 1600 3670 1620
rect 3690 1600 3760 1620
rect 3780 1600 3850 1620
rect 3870 1600 3940 1620
rect 3960 1600 4030 1620
rect 4050 1600 4120 1620
rect 4140 1600 4210 1620
rect 4230 1600 4300 1620
rect 4320 1600 4390 1620
rect 4410 1600 4480 1620
rect 4500 1600 4570 1620
rect 4590 1600 4660 1620
rect 4680 1600 4750 1620
rect 4770 1600 4840 1620
rect 4860 1600 4930 1620
rect 4950 1600 5020 1620
rect 5040 1600 5110 1620
rect 5130 1600 5200 1620
rect 5220 1600 5290 1620
rect 5310 1600 5380 1620
rect 5400 1600 5470 1620
rect 5490 1600 5560 1620
rect 5580 1600 5650 1620
rect 5670 1600 5740 1620
rect 5760 1600 5830 1620
rect 5850 1600 5920 1620
rect 5940 1600 6010 1620
rect 6030 1600 6100 1620
rect 6120 1600 6190 1620
rect 6210 1600 6280 1620
rect 6300 1600 6370 1620
rect 6390 1600 6460 1620
rect 6480 1600 6550 1620
rect 6570 1600 6640 1620
rect 6660 1600 6730 1620
rect 6750 1600 6820 1620
rect 6840 1600 6910 1620
rect 6930 1600 7000 1620
rect 7020 1600 7090 1620
rect 7110 1600 7180 1620
rect 7200 1600 7270 1620
rect 7290 1600 7360 1620
rect 7380 1600 7450 1620
rect 7470 1600 7540 1620
rect 7560 1600 7630 1620
rect 7650 1600 7720 1620
rect 7740 1600 7810 1620
rect 7830 1600 7900 1620
rect 7920 1600 7990 1620
rect 8010 1600 8080 1620
rect 8100 1600 8170 1620
rect 8190 1600 8260 1620
rect 8280 1600 8350 1620
rect 8370 1600 8440 1620
rect 8460 1600 8530 1620
rect 8550 1600 8620 1620
rect 8640 1600 8710 1620
rect 8730 1600 8800 1620
rect 8820 1600 8890 1620
rect 8910 1600 8980 1620
rect 9000 1600 9070 1620
rect 9090 1600 9160 1620
rect 9180 1600 9250 1620
rect 9270 1600 9340 1620
rect 9360 1600 9430 1620
rect 9450 1600 9520 1620
rect 9540 1600 9610 1620
rect 9630 1600 9700 1620
rect 9720 1600 9790 1620
rect 9810 1600 9880 1620
rect 9900 1600 9970 1620
rect 9990 1600 10060 1620
rect 10080 1600 10150 1620
rect 10170 1600 10240 1620
rect 10260 1600 10330 1620
rect 10350 1600 10420 1620
rect 10440 1600 10510 1620
rect 10530 1600 10600 1620
rect 10620 1600 10690 1620
rect 10710 1600 10780 1620
rect 10800 1600 10870 1620
rect 10890 1600 10960 1620
rect 10980 1600 11050 1620
rect 11070 1600 11140 1620
rect 11160 1600 11340 1620
rect -475 1240 -295 1260
rect -275 1240 -205 1260
rect -185 1240 -115 1260
rect -95 1240 -25 1260
rect -5 1240 65 1260
rect 85 1240 155 1260
rect 175 1240 245 1260
rect 265 1240 335 1260
rect 355 1240 425 1260
rect 445 1240 515 1260
rect 535 1240 605 1260
rect 625 1240 695 1260
rect 715 1240 785 1260
rect 805 1240 875 1260
rect 895 1240 965 1260
rect 985 1240 1055 1260
rect 1075 1240 1145 1260
rect 1165 1240 1235 1260
rect 1255 1240 1325 1260
rect 1345 1240 1415 1260
rect 1435 1240 1505 1260
rect 1525 1240 1595 1260
rect 1615 1240 1685 1260
rect 1705 1240 1775 1260
rect 1795 1240 1865 1260
rect 1885 1240 1955 1260
rect 1975 1240 2045 1260
rect 2065 1240 2135 1260
rect 2155 1240 2225 1260
rect 2245 1240 2315 1260
rect 2335 1240 2405 1260
rect 2425 1240 2495 1260
rect 2515 1240 2585 1260
rect 2605 1240 2675 1260
rect 2695 1240 2765 1260
rect 2785 1240 2855 1260
rect 2875 1240 2945 1260
rect 2965 1240 3035 1260
rect 3055 1240 3130 1260
rect 3150 1240 3220 1260
rect 3240 1240 3310 1260
rect 3330 1240 3400 1260
rect 3420 1240 3490 1260
rect 3510 1240 3580 1260
rect 3600 1240 3670 1260
rect 3690 1240 3760 1260
rect 3780 1240 3850 1260
rect 3870 1240 3940 1260
rect 3960 1240 4030 1260
rect 4050 1240 4120 1260
rect 4140 1240 4210 1260
rect 4230 1240 4300 1260
rect 4320 1240 4390 1260
rect 4410 1240 4480 1260
rect 4500 1240 4570 1260
rect 4590 1240 4660 1260
rect 4680 1240 4750 1260
rect 4770 1240 4840 1260
rect 4860 1240 4930 1260
rect 4950 1240 5020 1260
rect 5040 1240 5110 1260
rect 5130 1240 5200 1260
rect 5220 1240 5290 1260
rect 5310 1240 5380 1260
rect 5400 1240 5470 1260
rect 5490 1240 5560 1260
rect 5580 1240 5650 1260
rect 5670 1240 5740 1260
rect 5760 1240 5830 1260
rect 5850 1240 5920 1260
rect 5940 1240 6010 1260
rect 6030 1240 6100 1260
rect 6120 1240 6190 1260
rect 6210 1240 6280 1260
rect 6300 1240 6370 1260
rect 6390 1240 6460 1260
rect 6480 1240 6550 1260
rect 6570 1240 6640 1260
rect 6660 1240 6730 1260
rect 6750 1240 6820 1260
rect 6840 1240 6910 1260
rect 6930 1240 7000 1260
rect 7020 1240 7090 1260
rect 7110 1240 7180 1260
rect 7200 1240 7270 1260
rect 7290 1240 7360 1260
rect 7380 1240 7450 1260
rect 7470 1240 7540 1260
rect 7560 1240 7630 1260
rect 7650 1240 7720 1260
rect 7740 1240 7810 1260
rect 7830 1240 7900 1260
rect 7920 1240 7990 1260
rect 8010 1240 8080 1260
rect 8100 1240 8170 1260
rect 8190 1240 8260 1260
rect 8280 1240 8350 1260
rect 8370 1240 8440 1260
rect 8460 1240 8530 1260
rect 8550 1240 8620 1260
rect 8640 1240 8710 1260
rect 8730 1240 8800 1260
rect 8820 1240 8890 1260
rect 8910 1240 8980 1260
rect 9000 1240 9070 1260
rect 9090 1240 9160 1260
rect 9180 1240 9250 1260
rect 9270 1240 9340 1260
rect 9360 1240 9430 1260
rect 9450 1240 9520 1260
rect 9540 1240 9610 1260
rect 9630 1240 9700 1260
rect 9720 1240 9790 1260
rect 9810 1240 9880 1260
rect 9900 1240 9970 1260
rect 9990 1240 10060 1260
rect 10080 1240 10150 1260
rect 10170 1240 10240 1260
rect 10260 1240 10330 1260
rect 10350 1240 10420 1260
rect 10440 1240 10510 1260
rect 10530 1240 10600 1260
rect 10620 1240 10690 1260
rect 10710 1240 10780 1260
rect 10800 1240 10870 1260
rect 10890 1240 10960 1260
rect 10980 1240 11050 1260
rect 11070 1240 11140 1260
rect 11160 1240 11340 1260
rect -475 600 -455 1240
rect 11320 600 11340 1240
rect -475 580 -295 600
rect -275 580 -205 600
rect -185 580 -115 600
rect -95 580 -25 600
rect -5 580 65 600
rect 85 580 155 600
rect 175 580 245 600
rect 265 580 335 600
rect 355 580 425 600
rect 445 580 515 600
rect 535 580 605 600
rect 625 580 695 600
rect 715 580 785 600
rect 805 580 875 600
rect 895 580 965 600
rect 985 580 1055 600
rect 1075 580 1145 600
rect 1165 580 1235 600
rect 1255 580 1325 600
rect 1345 580 1415 600
rect 1435 580 1505 600
rect 1525 580 1595 600
rect 1615 580 1685 600
rect 1705 580 1775 600
rect 1795 580 1865 600
rect 1885 580 1955 600
rect 1975 580 2045 600
rect 2065 580 2135 600
rect 2155 580 2225 600
rect 2245 580 2315 600
rect 2335 580 2405 600
rect 2425 580 2495 600
rect 2515 580 2585 600
rect 2605 580 2675 600
rect 2695 580 2765 600
rect 2785 580 2855 600
rect 2875 580 2945 600
rect 2965 580 3035 600
rect 3055 580 3125 600
rect 3145 580 3215 600
rect 3235 580 3305 600
rect 3325 580 3395 600
rect 3415 580 3485 600
rect 3505 580 3575 600
rect 3595 580 3665 600
rect 3685 580 3755 600
rect 3775 580 3845 600
rect 3865 580 3935 600
rect 3955 580 4025 600
rect 4045 580 4115 600
rect 4135 580 4205 600
rect 4225 580 4295 600
rect 4315 580 4385 600
rect 4405 580 4475 600
rect 4495 580 4565 600
rect 4585 580 4655 600
rect 4675 580 4745 600
rect 4765 580 4835 600
rect 4855 580 4925 600
rect 4945 580 5015 600
rect 5035 580 5105 600
rect 5125 580 5195 600
rect 5215 580 5285 600
rect 5305 580 5375 600
rect 5395 580 5465 600
rect 5485 580 5555 600
rect 5575 580 5645 600
rect 5665 580 5735 600
rect 5755 580 5825 600
rect 5845 580 5915 600
rect 5935 580 6005 600
rect 6025 580 6095 600
rect 6115 580 6185 600
rect 6205 580 6275 600
rect 6295 580 6365 600
rect 6385 580 6455 600
rect 6475 580 6545 600
rect 6565 580 6635 600
rect 6655 580 6725 600
rect 6745 580 6815 600
rect 6835 580 6905 600
rect 6925 580 6995 600
rect 7015 580 7085 600
rect 7105 580 7175 600
rect 7195 580 7265 600
rect 7285 580 7355 600
rect 7375 580 7445 600
rect 7465 580 7535 600
rect 7555 580 7625 600
rect 7645 580 7715 600
rect 7735 580 7810 600
rect 7830 580 7900 600
rect 7920 580 7990 600
rect 8010 580 8080 600
rect 8100 580 8170 600
rect 8190 580 8260 600
rect 8280 580 8350 600
rect 8370 580 8440 600
rect 8460 580 8530 600
rect 8550 580 8620 600
rect 8640 580 8710 600
rect 8730 580 8800 600
rect 8820 580 8890 600
rect 8910 580 8980 600
rect 9000 580 9070 600
rect 9090 580 9160 600
rect 9180 580 9250 600
rect 9270 580 9340 600
rect 9360 580 9430 600
rect 9450 580 9520 600
rect 9540 580 9610 600
rect 9630 580 9700 600
rect 9720 580 9790 600
rect 9810 580 9880 600
rect 9900 580 9970 600
rect 9990 580 10060 600
rect 10080 580 10150 600
rect 10170 580 10240 600
rect 10260 580 10330 600
rect 10350 580 10420 600
rect 10440 580 10510 600
rect 10530 580 10600 600
rect 10620 580 10690 600
rect 10710 580 10780 600
rect 10800 580 10870 600
rect 10890 580 10960 600
rect 10980 580 11050 600
rect 11070 580 11140 600
rect 11160 580 11340 600
rect -475 220 -295 240
rect -275 220 -205 240
rect -185 220 -115 240
rect -95 220 -25 240
rect -5 220 65 240
rect 85 220 155 240
rect 175 220 245 240
rect 265 220 335 240
rect 355 220 425 240
rect 445 220 515 240
rect 535 220 605 240
rect 625 220 695 240
rect 715 220 785 240
rect 805 220 875 240
rect 895 220 965 240
rect 985 220 1055 240
rect 1075 220 1145 240
rect 1165 220 1235 240
rect 1255 220 1325 240
rect 1345 220 1415 240
rect 1435 220 1505 240
rect 1525 220 1595 240
rect 1615 220 1685 240
rect 1705 220 1775 240
rect 1795 220 1865 240
rect 1885 220 1955 240
rect 1975 220 2045 240
rect 2065 220 2135 240
rect 2155 220 2225 240
rect 2245 220 2315 240
rect 2335 220 2405 240
rect 2425 220 2495 240
rect 2515 220 2585 240
rect 2605 220 2675 240
rect 2695 220 2765 240
rect 2785 220 2855 240
rect 2875 220 2945 240
rect 2965 220 3035 240
rect 3055 220 3125 240
rect 3145 220 3215 240
rect 3235 220 3305 240
rect 3325 220 3395 240
rect 3415 220 3485 240
rect 3505 220 3575 240
rect 3595 220 3665 240
rect 3685 220 3755 240
rect 3775 220 3845 240
rect 3865 220 3935 240
rect 3955 220 4025 240
rect 4045 220 4115 240
rect 4135 220 4205 240
rect 4225 220 4295 240
rect 4315 220 4385 240
rect 4405 220 4475 240
rect 4495 220 4565 240
rect 4585 220 4655 240
rect 4675 220 4745 240
rect 4765 220 4835 240
rect 4855 220 4925 240
rect 4945 220 5015 240
rect 5035 220 5105 240
rect 5125 220 5195 240
rect 5215 220 5285 240
rect 5305 220 5375 240
rect 5395 220 5465 240
rect 5485 220 5555 240
rect 5575 220 5645 240
rect 5665 220 5735 240
rect 5755 220 5825 240
rect 5845 220 5915 240
rect 5935 220 6005 240
rect 6025 220 6095 240
rect 6115 220 6185 240
rect 6205 220 6275 240
rect 6295 220 6365 240
rect 6385 220 6455 240
rect 6475 220 6545 240
rect 6565 220 6635 240
rect 6655 220 6725 240
rect 6745 220 6815 240
rect 6835 220 6905 240
rect 6925 220 6995 240
rect 7015 220 7085 240
rect 7105 220 7175 240
rect 7195 220 7265 240
rect 7285 220 7355 240
rect 7375 220 7445 240
rect 7465 220 7535 240
rect 7555 220 7625 240
rect 7645 220 7715 240
rect 7735 220 7810 240
rect 7830 220 7900 240
rect 7920 220 7990 240
rect 8010 220 8080 240
rect 8100 220 8170 240
rect 8190 220 8260 240
rect 8280 220 8350 240
rect 8370 220 8440 240
rect 8460 220 8530 240
rect 8550 220 8620 240
rect 8640 220 8710 240
rect 8730 220 8800 240
rect 8820 220 8890 240
rect 8910 220 8980 240
rect 9000 220 9070 240
rect 9090 220 9160 240
rect 9180 220 9250 240
rect 9270 220 9340 240
rect 9360 220 9430 240
rect 9450 220 9520 240
rect 9540 220 9610 240
rect 9630 220 9700 240
rect 9720 220 9790 240
rect 9810 220 9880 240
rect 9900 220 9970 240
rect 9990 220 10060 240
rect 10080 220 10150 240
rect 10170 220 10240 240
rect 10260 220 10330 240
rect 10350 220 10420 240
rect 10440 220 10510 240
rect 10530 220 10600 240
rect 10620 220 10690 240
rect 10710 220 10780 240
rect 10800 220 10870 240
rect 10890 220 10960 240
rect 10980 220 11050 240
rect 11070 220 11140 240
rect 11160 220 11340 240
rect -475 20 -455 220
rect 11320 20 11340 220
rect -485 0 -295 20
rect -275 0 -205 20
rect -185 0 -115 20
rect -95 0 -25 20
rect -5 0 65 20
rect 85 0 155 20
rect 175 0 245 20
rect 265 0 335 20
rect 355 0 425 20
rect 445 0 515 20
rect 535 0 605 20
rect 625 0 695 20
rect 715 0 785 20
rect 805 0 875 20
rect 895 0 965 20
rect 985 0 1055 20
rect 1075 0 1145 20
rect 1165 0 1235 20
rect 1255 0 1325 20
rect 1345 0 1415 20
rect 1435 0 1505 20
rect 1525 0 1595 20
rect 1615 0 1685 20
rect 1705 0 1775 20
rect 1795 0 1865 20
rect 1885 0 1955 20
rect 1975 0 2045 20
rect 2065 0 2135 20
rect 2155 0 2225 20
rect 2245 0 2315 20
rect 2335 0 2405 20
rect 2425 0 2495 20
rect 2515 0 2585 20
rect 2605 0 2675 20
rect 2695 0 2765 20
rect 2785 0 2855 20
rect 2875 0 2945 20
rect 2965 0 3035 20
rect 3055 0 3125 20
rect 3145 0 3215 20
rect 3235 0 3305 20
rect 3325 0 3395 20
rect 3415 0 3485 20
rect 3505 0 3575 20
rect 3595 0 3665 20
rect 3685 0 3755 20
rect 3775 0 3845 20
rect 3865 0 3935 20
rect 3955 0 4025 20
rect 4045 0 4115 20
rect 4135 0 4205 20
rect 4225 0 4295 20
rect 4315 0 4385 20
rect 4405 0 4475 20
rect 4495 0 4565 20
rect 4585 0 4655 20
rect 4675 0 4745 20
rect 4765 0 4835 20
rect 4855 0 4925 20
rect 4945 0 5015 20
rect 5035 0 5105 20
rect 5125 0 5195 20
rect 5215 0 5285 20
rect 5305 0 5375 20
rect 5395 0 5465 20
rect 5485 0 5555 20
rect 5575 0 5645 20
rect 5665 0 5735 20
rect 5755 0 5825 20
rect 5845 0 5915 20
rect 5935 0 6005 20
rect 6025 0 6095 20
rect 6115 0 6185 20
rect 6205 0 6275 20
rect 6295 0 6365 20
rect 6385 0 6455 20
rect 6475 0 6545 20
rect 6565 0 6635 20
rect 6655 0 6725 20
rect 6745 0 6815 20
rect 6835 0 6905 20
rect 6925 0 6995 20
rect 7015 0 7085 20
rect 7105 0 7175 20
rect 7195 0 7265 20
rect 7285 0 7355 20
rect 7375 0 7445 20
rect 7465 0 7535 20
rect 7555 0 7625 20
rect 7645 0 7715 20
rect 7735 0 7810 20
rect 7830 0 7900 20
rect 7920 0 7990 20
rect 8010 0 8080 20
rect 8100 0 8170 20
rect 8190 0 8260 20
rect 8280 0 8350 20
rect 8370 0 8440 20
rect 8460 0 8530 20
rect 8550 0 8620 20
rect 8640 0 8710 20
rect 8730 0 8800 20
rect 8820 0 8890 20
rect 8910 0 8980 20
rect 9000 0 9070 20
rect 9090 0 9160 20
rect 9180 0 9250 20
rect 9270 0 9340 20
rect 9360 0 9430 20
rect 9450 0 9520 20
rect 9540 0 9610 20
rect 9630 0 9700 20
rect 9720 0 9790 20
rect 9810 0 9880 20
rect 9900 0 9970 20
rect 9990 0 10060 20
rect 10080 0 10150 20
rect 10170 0 10240 20
rect 10260 0 10330 20
rect 10350 0 10420 20
rect 10440 0 10510 20
rect 10530 0 10600 20
rect 10620 0 10690 20
rect 10710 0 10780 20
rect 10800 0 10870 20
rect 10890 0 10960 20
rect 10980 0 11050 20
rect 11070 0 11140 20
rect 11160 0 11350 20
<< nsubdiff >>
rect -400 1160 -295 1180
rect -275 1160 -205 1180
rect -185 1160 -115 1180
rect -95 1160 -25 1180
rect -5 1160 65 1180
rect 85 1160 155 1180
rect 175 1160 245 1180
rect 265 1160 335 1180
rect 355 1160 425 1180
rect 445 1160 515 1180
rect 535 1160 605 1180
rect 625 1160 695 1180
rect 715 1160 785 1180
rect 805 1160 875 1180
rect 895 1160 965 1180
rect 985 1160 1055 1180
rect 1075 1160 1145 1180
rect 1165 1160 1235 1180
rect 1255 1160 1325 1180
rect 1345 1160 1415 1180
rect 1435 1160 1505 1180
rect 1525 1160 1595 1180
rect 1615 1160 1685 1180
rect 1705 1160 1775 1180
rect 1795 1160 1865 1180
rect 1885 1160 1955 1180
rect 1975 1160 2045 1180
rect 2065 1160 2135 1180
rect 2155 1160 2225 1180
rect 2245 1160 2315 1180
rect 2335 1160 2405 1180
rect 2425 1160 2495 1180
rect 2515 1160 2585 1180
rect 2605 1160 2675 1180
rect 2695 1160 2765 1180
rect 2785 1160 2855 1180
rect 2875 1160 2945 1180
rect 2965 1160 3035 1180
rect 3055 1160 3130 1180
rect 3150 1160 3220 1180
rect 3240 1160 3310 1180
rect 3330 1160 3400 1180
rect 3420 1160 3490 1180
rect 3510 1160 3580 1180
rect 3600 1160 3670 1180
rect 3690 1160 3760 1180
rect 3780 1160 3850 1180
rect 3870 1160 3940 1180
rect 3960 1160 4030 1180
rect 4050 1160 4120 1180
rect 4140 1160 4210 1180
rect 4230 1160 4300 1180
rect 4320 1160 4390 1180
rect 4410 1160 4480 1180
rect 4500 1160 4570 1180
rect 4590 1160 4660 1180
rect 4680 1160 4750 1180
rect 4770 1160 4840 1180
rect 4860 1160 4930 1180
rect 4950 1160 5020 1180
rect 5040 1160 5110 1180
rect 5130 1160 5200 1180
rect 5220 1160 5290 1180
rect 5310 1160 5380 1180
rect 5400 1160 5470 1180
rect 5490 1160 5560 1180
rect 5580 1160 5650 1180
rect 5670 1160 5740 1180
rect 5760 1160 5830 1180
rect 5850 1160 5920 1180
rect 5940 1160 6010 1180
rect 6030 1160 6100 1180
rect 6120 1160 6190 1180
rect 6210 1160 6280 1180
rect 6300 1160 6370 1180
rect 6390 1160 6460 1180
rect 6480 1160 6550 1180
rect 6570 1160 6640 1180
rect 6660 1160 6730 1180
rect 6750 1160 6820 1180
rect 6840 1160 6910 1180
rect 6930 1160 7000 1180
rect 7020 1160 7090 1180
rect 7110 1160 7180 1180
rect 7200 1160 7270 1180
rect 7290 1160 7360 1180
rect 7380 1160 7450 1180
rect 7470 1160 7540 1180
rect 7560 1160 7630 1180
rect 7650 1160 7720 1180
rect 7740 1160 7810 1180
rect 7830 1160 7900 1180
rect 7920 1160 7990 1180
rect 8010 1160 8080 1180
rect 8100 1160 8170 1180
rect 8190 1160 8260 1180
rect 8280 1160 8350 1180
rect 8370 1160 8440 1180
rect 8460 1160 8530 1180
rect 8550 1160 8620 1180
rect 8640 1160 8710 1180
rect 8730 1160 8800 1180
rect 8820 1160 8890 1180
rect 8910 1160 8980 1180
rect 9000 1160 9070 1180
rect 9090 1160 9160 1180
rect 9180 1160 9250 1180
rect 9270 1160 9340 1180
rect 9360 1160 9430 1180
rect 9450 1160 9520 1180
rect 9540 1160 9610 1180
rect 9630 1160 9700 1180
rect 9720 1160 9790 1180
rect 9810 1160 9880 1180
rect 9900 1160 9970 1180
rect 9990 1160 10060 1180
rect 10080 1160 10150 1180
rect 10170 1160 10240 1180
rect 10260 1160 10330 1180
rect 10350 1160 10420 1180
rect 10440 1160 10510 1180
rect 10530 1160 10600 1180
rect 10620 1160 10690 1180
rect 10710 1160 10780 1180
rect 10800 1160 10870 1180
rect 10890 1160 10960 1180
rect 10980 1160 11050 1180
rect 11070 1160 11140 1180
rect 11160 1160 11265 1180
rect -400 960 -380 1160
rect 11245 960 11265 1160
rect -400 940 -295 960
rect -275 940 -205 960
rect -185 940 -115 960
rect -95 940 -25 960
rect -5 940 65 960
rect 85 940 155 960
rect 175 940 245 960
rect 265 940 335 960
rect 355 940 425 960
rect 445 940 515 960
rect 535 940 605 960
rect 625 940 695 960
rect 715 940 785 960
rect 805 940 875 960
rect 895 940 965 960
rect 985 940 1055 960
rect 1075 940 1145 960
rect 1165 940 1235 960
rect 1255 940 1325 960
rect 1345 940 1415 960
rect 1435 940 1505 960
rect 1525 940 1595 960
rect 1615 940 1685 960
rect 1705 940 1775 960
rect 1795 940 1865 960
rect 1885 940 1955 960
rect 1975 940 2045 960
rect 2065 940 2135 960
rect 2155 940 2225 960
rect 2245 940 2315 960
rect 2335 940 2405 960
rect 2425 940 2495 960
rect 2515 940 2585 960
rect 2605 940 2675 960
rect 2695 940 2765 960
rect 2785 940 2855 960
rect 2875 940 2945 960
rect 2965 940 3035 960
rect 3055 940 3130 960
rect 3150 940 3220 960
rect 3240 940 3310 960
rect 3330 940 3400 960
rect 3420 940 3490 960
rect 3510 940 3580 960
rect 3600 940 3670 960
rect 3690 940 3760 960
rect 3780 940 3850 960
rect 3870 940 3940 960
rect 3960 940 4030 960
rect 4050 940 4120 960
rect 4140 940 4210 960
rect 4230 940 4300 960
rect 4320 940 4390 960
rect 4410 940 4480 960
rect 4500 940 4570 960
rect 4590 940 4660 960
rect 4680 940 4750 960
rect 4770 940 4840 960
rect 4860 940 4930 960
rect 4950 940 5020 960
rect 5040 940 5110 960
rect 5130 940 5200 960
rect 5220 940 5290 960
rect 5310 940 5380 960
rect 5400 940 5470 960
rect 5490 940 5560 960
rect 5580 940 5650 960
rect 5670 940 5740 960
rect 5760 940 5830 960
rect 5850 940 5920 960
rect 5940 940 6010 960
rect 6030 940 6100 960
rect 6120 940 6190 960
rect 6210 940 6280 960
rect 6300 940 6370 960
rect 6390 940 6460 960
rect 6480 940 6550 960
rect 6570 940 6640 960
rect 6660 940 6730 960
rect 6750 940 6820 960
rect 6840 940 6910 960
rect 6930 940 7000 960
rect 7020 940 7090 960
rect 7110 940 7180 960
rect 7200 940 7270 960
rect 7290 940 7360 960
rect 7380 940 7450 960
rect 7470 940 7540 960
rect 7560 940 7630 960
rect 7650 940 7720 960
rect 7740 940 7810 960
rect 7830 940 7900 960
rect 7920 940 7990 960
rect 8010 940 8080 960
rect 8100 940 8170 960
rect 8190 940 8260 960
rect 8280 940 8350 960
rect 8370 940 8440 960
rect 8460 940 8530 960
rect 8550 940 8620 960
rect 8640 940 8710 960
rect 8730 940 8800 960
rect 8820 940 8890 960
rect 8910 940 8980 960
rect 9000 940 9070 960
rect 9090 940 9160 960
rect 9180 940 9250 960
rect 9270 940 9340 960
rect 9360 940 9430 960
rect 9450 940 9520 960
rect 9540 940 9610 960
rect 9630 940 9700 960
rect 9720 940 9790 960
rect 9810 940 9880 960
rect 9900 940 9970 960
rect 9990 940 10060 960
rect 10080 940 10150 960
rect 10170 940 10240 960
rect 10260 940 10330 960
rect 10350 940 10420 960
rect 10440 940 10510 960
rect 10530 940 10600 960
rect 10620 940 10690 960
rect 10710 940 10780 960
rect 10800 940 10870 960
rect 10890 940 10960 960
rect 10980 940 11050 960
rect 11070 940 11140 960
rect 11160 940 11265 960
rect -400 880 -295 900
rect -275 880 -205 900
rect -185 880 -115 900
rect -95 880 -25 900
rect -5 880 65 900
rect 85 880 155 900
rect 175 880 245 900
rect 265 880 335 900
rect 355 880 425 900
rect 445 880 515 900
rect 535 880 605 900
rect 625 880 695 900
rect 715 880 785 900
rect 805 880 875 900
rect 895 880 965 900
rect 985 880 1055 900
rect 1075 880 1145 900
rect 1165 880 1235 900
rect 1255 880 1325 900
rect 1345 880 1415 900
rect 1435 880 1505 900
rect 1525 880 1595 900
rect 1615 880 1685 900
rect 1705 880 1775 900
rect 1795 880 1865 900
rect 1885 880 1955 900
rect 1975 880 2045 900
rect 2065 880 2135 900
rect 2155 880 2225 900
rect 2245 880 2315 900
rect 2335 880 2405 900
rect 2425 880 2495 900
rect 2515 880 2585 900
rect 2605 880 2675 900
rect 2695 880 2765 900
rect 2785 880 2855 900
rect 2875 880 2945 900
rect 2965 880 3035 900
rect 3055 880 3125 900
rect 3145 880 3215 900
rect 3235 880 3305 900
rect 3325 880 3395 900
rect 3415 880 3485 900
rect 3505 880 3575 900
rect 3595 880 3665 900
rect 3685 880 3755 900
rect 3775 880 3845 900
rect 3865 880 3935 900
rect 3955 880 4025 900
rect 4045 880 4115 900
rect 4135 880 4205 900
rect 4225 880 4295 900
rect 4315 880 4385 900
rect 4405 880 4475 900
rect 4495 880 4565 900
rect 4585 880 4655 900
rect 4675 880 4745 900
rect 4765 880 4835 900
rect 4855 880 4925 900
rect 4945 880 5015 900
rect 5035 880 5105 900
rect 5125 880 5195 900
rect 5215 880 5285 900
rect 5305 880 5375 900
rect 5395 880 5465 900
rect 5485 880 5555 900
rect 5575 880 5645 900
rect 5665 880 5735 900
rect 5755 880 5825 900
rect 5845 880 5915 900
rect 5935 880 6005 900
rect 6025 880 6095 900
rect 6115 880 6185 900
rect 6205 880 6275 900
rect 6295 880 6365 900
rect 6385 880 6455 900
rect 6475 880 6545 900
rect 6565 880 6635 900
rect 6655 880 6725 900
rect 6745 880 6815 900
rect 6835 880 6905 900
rect 6925 880 6995 900
rect 7015 880 7085 900
rect 7105 880 7175 900
rect 7195 880 7265 900
rect 7285 880 7355 900
rect 7375 880 7445 900
rect 7465 880 7535 900
rect 7555 880 7625 900
rect 7645 880 7715 900
rect 7735 880 7810 900
rect 7830 880 7900 900
rect 7920 880 7990 900
rect 8010 880 8080 900
rect 8100 880 8170 900
rect 8190 880 8260 900
rect 8280 880 8350 900
rect 8370 880 8440 900
rect 8460 880 8530 900
rect 8550 880 8620 900
rect 8640 880 8710 900
rect 8730 880 8800 900
rect 8820 880 8890 900
rect 8910 880 8980 900
rect 9000 880 9070 900
rect 9090 880 9160 900
rect 9180 880 9250 900
rect 9270 880 9340 900
rect 9360 880 9430 900
rect 9450 880 9520 900
rect 9540 880 9610 900
rect 9630 880 9700 900
rect 9720 880 9790 900
rect 9810 880 9880 900
rect 9900 880 9970 900
rect 9990 880 10060 900
rect 10080 880 10150 900
rect 10170 880 10240 900
rect 10260 880 10330 900
rect 10350 880 10420 900
rect 10440 880 10510 900
rect 10530 880 10600 900
rect 10620 880 10690 900
rect 10710 880 10780 900
rect 10800 880 10870 900
rect 10890 880 10960 900
rect 10980 880 11050 900
rect 11070 880 11140 900
rect 11160 880 11265 900
rect -400 680 -380 880
rect 11245 680 11265 880
rect -400 660 -295 680
rect -275 660 -205 680
rect -185 660 -115 680
rect -95 660 -25 680
rect -5 660 65 680
rect 85 660 155 680
rect 175 660 245 680
rect 265 660 335 680
rect 355 660 425 680
rect 445 660 515 680
rect 535 660 605 680
rect 625 660 695 680
rect 715 660 785 680
rect 805 660 875 680
rect 895 660 965 680
rect 985 660 1055 680
rect 1075 660 1145 680
rect 1165 660 1235 680
rect 1255 660 1325 680
rect 1345 660 1415 680
rect 1435 660 1505 680
rect 1525 660 1595 680
rect 1615 660 1685 680
rect 1705 660 1775 680
rect 1795 660 1865 680
rect 1885 660 1955 680
rect 1975 660 2045 680
rect 2065 660 2135 680
rect 2155 660 2225 680
rect 2245 660 2315 680
rect 2335 660 2405 680
rect 2425 660 2495 680
rect 2515 660 2585 680
rect 2605 660 2675 680
rect 2695 660 2765 680
rect 2785 660 2855 680
rect 2875 660 2945 680
rect 2965 660 3035 680
rect 3055 660 3125 680
rect 3145 660 3215 680
rect 3235 660 3305 680
rect 3325 660 3395 680
rect 3415 660 3485 680
rect 3505 660 3575 680
rect 3595 660 3665 680
rect 3685 660 3755 680
rect 3775 660 3845 680
rect 3865 660 3935 680
rect 3955 660 4025 680
rect 4045 660 4115 680
rect 4135 660 4205 680
rect 4225 660 4295 680
rect 4315 660 4385 680
rect 4405 660 4475 680
rect 4495 660 4565 680
rect 4585 660 4655 680
rect 4675 660 4745 680
rect 4765 660 4835 680
rect 4855 660 4925 680
rect 4945 660 5015 680
rect 5035 660 5105 680
rect 5125 660 5195 680
rect 5215 660 5285 680
rect 5305 660 5375 680
rect 5395 660 5465 680
rect 5485 660 5555 680
rect 5575 660 5645 680
rect 5665 660 5735 680
rect 5755 660 5825 680
rect 5845 660 5915 680
rect 5935 660 6005 680
rect 6025 660 6095 680
rect 6115 660 6185 680
rect 6205 660 6275 680
rect 6295 660 6365 680
rect 6385 660 6455 680
rect 6475 660 6545 680
rect 6565 660 6635 680
rect 6655 660 6725 680
rect 6745 660 6815 680
rect 6835 660 6905 680
rect 6925 660 6995 680
rect 7015 660 7085 680
rect 7105 660 7175 680
rect 7195 660 7265 680
rect 7285 660 7355 680
rect 7375 660 7445 680
rect 7465 660 7535 680
rect 7555 660 7625 680
rect 7645 660 7715 680
rect 7735 660 7810 680
rect 7830 660 7900 680
rect 7920 660 7990 680
rect 8010 660 8080 680
rect 8100 660 8170 680
rect 8190 660 8260 680
rect 8280 660 8350 680
rect 8370 660 8440 680
rect 8460 660 8530 680
rect 8550 660 8620 680
rect 8640 660 8710 680
rect 8730 660 8800 680
rect 8820 660 8890 680
rect 8910 660 8980 680
rect 9000 660 9070 680
rect 9090 660 9160 680
rect 9180 660 9250 680
rect 9270 660 9340 680
rect 9360 660 9430 680
rect 9450 660 9520 680
rect 9540 660 9610 680
rect 9630 660 9700 680
rect 9720 660 9790 680
rect 9810 660 9880 680
rect 9900 660 9970 680
rect 9990 660 10060 680
rect 10080 660 10150 680
rect 10170 660 10240 680
rect 10260 660 10330 680
rect 10350 660 10420 680
rect 10440 660 10510 680
rect 10530 660 10600 680
rect 10620 660 10690 680
rect 10710 660 10780 680
rect 10800 660 10870 680
rect 10890 660 10960 680
rect 10980 660 11050 680
rect 11070 660 11140 680
rect 11160 660 11265 680
<< psubdiffcont >>
rect -295 1820 -275 1840
rect -205 1820 -185 1840
rect -115 1820 -95 1840
rect -25 1820 -5 1840
rect 65 1820 85 1840
rect 155 1820 175 1840
rect 245 1820 265 1840
rect 335 1820 355 1840
rect 425 1820 445 1840
rect 515 1820 535 1840
rect 605 1820 625 1840
rect 695 1820 715 1840
rect 785 1820 805 1840
rect 875 1820 895 1840
rect 965 1820 985 1840
rect 1055 1820 1075 1840
rect 1145 1820 1165 1840
rect 1235 1820 1255 1840
rect 1325 1820 1345 1840
rect 1415 1820 1435 1840
rect 1505 1820 1525 1840
rect 1595 1820 1615 1840
rect 1685 1820 1705 1840
rect 1775 1820 1795 1840
rect 1865 1820 1885 1840
rect 1955 1820 1975 1840
rect 2045 1820 2065 1840
rect 2135 1820 2155 1840
rect 2225 1820 2245 1840
rect 2315 1820 2335 1840
rect 2405 1820 2425 1840
rect 2495 1820 2515 1840
rect 2585 1820 2605 1840
rect 2675 1820 2695 1840
rect 2765 1820 2785 1840
rect 2855 1820 2875 1840
rect 2945 1820 2965 1840
rect 3035 1820 3055 1840
rect 3130 1820 3150 1840
rect 3220 1820 3240 1840
rect 3310 1820 3330 1840
rect 3400 1820 3420 1840
rect 3490 1820 3510 1840
rect 3580 1820 3600 1840
rect 3670 1820 3690 1840
rect 3760 1820 3780 1840
rect 3850 1820 3870 1840
rect 3940 1820 3960 1840
rect 4030 1820 4050 1840
rect 4120 1820 4140 1840
rect 4210 1820 4230 1840
rect 4300 1820 4320 1840
rect 4390 1820 4410 1840
rect 4480 1820 4500 1840
rect 4570 1820 4590 1840
rect 4660 1820 4680 1840
rect 4750 1820 4770 1840
rect 4840 1820 4860 1840
rect 4930 1820 4950 1840
rect 5020 1820 5040 1840
rect 5110 1820 5130 1840
rect 5200 1820 5220 1840
rect 5290 1820 5310 1840
rect 5380 1820 5400 1840
rect 5470 1820 5490 1840
rect 5560 1820 5580 1840
rect 5650 1820 5670 1840
rect 5740 1820 5760 1840
rect 5830 1820 5850 1840
rect 5920 1820 5940 1840
rect 6010 1820 6030 1840
rect 6100 1820 6120 1840
rect 6190 1820 6210 1840
rect 6280 1820 6300 1840
rect 6370 1820 6390 1840
rect 6460 1820 6480 1840
rect 6550 1820 6570 1840
rect 6640 1820 6660 1840
rect 6730 1820 6750 1840
rect 6820 1820 6840 1840
rect 6910 1820 6930 1840
rect 7000 1820 7020 1840
rect 7090 1820 7110 1840
rect 7180 1820 7200 1840
rect 7270 1820 7290 1840
rect 7360 1820 7380 1840
rect 7450 1820 7470 1840
rect 7540 1820 7560 1840
rect 7630 1820 7650 1840
rect 7720 1820 7740 1840
rect 7810 1820 7830 1840
rect 7900 1820 7920 1840
rect 7990 1820 8010 1840
rect 8080 1820 8100 1840
rect 8170 1820 8190 1840
rect 8260 1820 8280 1840
rect 8350 1820 8370 1840
rect 8440 1820 8460 1840
rect 8530 1820 8550 1840
rect 8620 1820 8640 1840
rect 8710 1820 8730 1840
rect 8800 1820 8820 1840
rect 8890 1820 8910 1840
rect 8980 1820 9000 1840
rect 9070 1820 9090 1840
rect 9160 1820 9180 1840
rect 9250 1820 9270 1840
rect 9340 1820 9360 1840
rect 9430 1820 9450 1840
rect 9520 1820 9540 1840
rect 9610 1820 9630 1840
rect 9700 1820 9720 1840
rect 9790 1820 9810 1840
rect 9880 1820 9900 1840
rect 9970 1820 9990 1840
rect 10060 1820 10080 1840
rect 10150 1820 10170 1840
rect 10240 1820 10260 1840
rect 10330 1820 10350 1840
rect 10420 1820 10440 1840
rect 10510 1820 10530 1840
rect 10600 1820 10620 1840
rect 10690 1820 10710 1840
rect 10780 1820 10800 1840
rect 10870 1820 10890 1840
rect 10960 1820 10980 1840
rect 11050 1820 11070 1840
rect 11140 1820 11160 1840
rect -295 1600 -275 1620
rect -205 1600 -185 1620
rect -115 1600 -95 1620
rect -25 1600 -5 1620
rect 65 1600 85 1620
rect 155 1600 175 1620
rect 245 1600 265 1620
rect 335 1600 355 1620
rect 425 1600 445 1620
rect 515 1600 535 1620
rect 605 1600 625 1620
rect 695 1600 715 1620
rect 785 1600 805 1620
rect 875 1600 895 1620
rect 965 1600 985 1620
rect 1055 1600 1075 1620
rect 1145 1600 1165 1620
rect 1235 1600 1255 1620
rect 1325 1600 1345 1620
rect 1415 1600 1435 1620
rect 1505 1600 1525 1620
rect 1595 1600 1615 1620
rect 1685 1600 1705 1620
rect 1775 1600 1795 1620
rect 1865 1600 1885 1620
rect 1955 1600 1975 1620
rect 2045 1600 2065 1620
rect 2135 1600 2155 1620
rect 2225 1600 2245 1620
rect 2315 1600 2335 1620
rect 2405 1600 2425 1620
rect 2495 1600 2515 1620
rect 2585 1600 2605 1620
rect 2675 1600 2695 1620
rect 2765 1600 2785 1620
rect 2855 1600 2875 1620
rect 2945 1600 2965 1620
rect 3035 1600 3055 1620
rect 3130 1600 3150 1620
rect 3220 1600 3240 1620
rect 3310 1600 3330 1620
rect 3400 1600 3420 1620
rect 3490 1600 3510 1620
rect 3580 1600 3600 1620
rect 3670 1600 3690 1620
rect 3760 1600 3780 1620
rect 3850 1600 3870 1620
rect 3940 1600 3960 1620
rect 4030 1600 4050 1620
rect 4120 1600 4140 1620
rect 4210 1600 4230 1620
rect 4300 1600 4320 1620
rect 4390 1600 4410 1620
rect 4480 1600 4500 1620
rect 4570 1600 4590 1620
rect 4660 1600 4680 1620
rect 4750 1600 4770 1620
rect 4840 1600 4860 1620
rect 4930 1600 4950 1620
rect 5020 1600 5040 1620
rect 5110 1600 5130 1620
rect 5200 1600 5220 1620
rect 5290 1600 5310 1620
rect 5380 1600 5400 1620
rect 5470 1600 5490 1620
rect 5560 1600 5580 1620
rect 5650 1600 5670 1620
rect 5740 1600 5760 1620
rect 5830 1600 5850 1620
rect 5920 1600 5940 1620
rect 6010 1600 6030 1620
rect 6100 1600 6120 1620
rect 6190 1600 6210 1620
rect 6280 1600 6300 1620
rect 6370 1600 6390 1620
rect 6460 1600 6480 1620
rect 6550 1600 6570 1620
rect 6640 1600 6660 1620
rect 6730 1600 6750 1620
rect 6820 1600 6840 1620
rect 6910 1600 6930 1620
rect 7000 1600 7020 1620
rect 7090 1600 7110 1620
rect 7180 1600 7200 1620
rect 7270 1600 7290 1620
rect 7360 1600 7380 1620
rect 7450 1600 7470 1620
rect 7540 1600 7560 1620
rect 7630 1600 7650 1620
rect 7720 1600 7740 1620
rect 7810 1600 7830 1620
rect 7900 1600 7920 1620
rect 7990 1600 8010 1620
rect 8080 1600 8100 1620
rect 8170 1600 8190 1620
rect 8260 1600 8280 1620
rect 8350 1600 8370 1620
rect 8440 1600 8460 1620
rect 8530 1600 8550 1620
rect 8620 1600 8640 1620
rect 8710 1600 8730 1620
rect 8800 1600 8820 1620
rect 8890 1600 8910 1620
rect 8980 1600 9000 1620
rect 9070 1600 9090 1620
rect 9160 1600 9180 1620
rect 9250 1600 9270 1620
rect 9340 1600 9360 1620
rect 9430 1600 9450 1620
rect 9520 1600 9540 1620
rect 9610 1600 9630 1620
rect 9700 1600 9720 1620
rect 9790 1600 9810 1620
rect 9880 1600 9900 1620
rect 9970 1600 9990 1620
rect 10060 1600 10080 1620
rect 10150 1600 10170 1620
rect 10240 1600 10260 1620
rect 10330 1600 10350 1620
rect 10420 1600 10440 1620
rect 10510 1600 10530 1620
rect 10600 1600 10620 1620
rect 10690 1600 10710 1620
rect 10780 1600 10800 1620
rect 10870 1600 10890 1620
rect 10960 1600 10980 1620
rect 11050 1600 11070 1620
rect 11140 1600 11160 1620
rect -295 1240 -275 1260
rect -205 1240 -185 1260
rect -115 1240 -95 1260
rect -25 1240 -5 1260
rect 65 1240 85 1260
rect 155 1240 175 1260
rect 245 1240 265 1260
rect 335 1240 355 1260
rect 425 1240 445 1260
rect 515 1240 535 1260
rect 605 1240 625 1260
rect 695 1240 715 1260
rect 785 1240 805 1260
rect 875 1240 895 1260
rect 965 1240 985 1260
rect 1055 1240 1075 1260
rect 1145 1240 1165 1260
rect 1235 1240 1255 1260
rect 1325 1240 1345 1260
rect 1415 1240 1435 1260
rect 1505 1240 1525 1260
rect 1595 1240 1615 1260
rect 1685 1240 1705 1260
rect 1775 1240 1795 1260
rect 1865 1240 1885 1260
rect 1955 1240 1975 1260
rect 2045 1240 2065 1260
rect 2135 1240 2155 1260
rect 2225 1240 2245 1260
rect 2315 1240 2335 1260
rect 2405 1240 2425 1260
rect 2495 1240 2515 1260
rect 2585 1240 2605 1260
rect 2675 1240 2695 1260
rect 2765 1240 2785 1260
rect 2855 1240 2875 1260
rect 2945 1240 2965 1260
rect 3035 1240 3055 1260
rect 3130 1240 3150 1260
rect 3220 1240 3240 1260
rect 3310 1240 3330 1260
rect 3400 1240 3420 1260
rect 3490 1240 3510 1260
rect 3580 1240 3600 1260
rect 3670 1240 3690 1260
rect 3760 1240 3780 1260
rect 3850 1240 3870 1260
rect 3940 1240 3960 1260
rect 4030 1240 4050 1260
rect 4120 1240 4140 1260
rect 4210 1240 4230 1260
rect 4300 1240 4320 1260
rect 4390 1240 4410 1260
rect 4480 1240 4500 1260
rect 4570 1240 4590 1260
rect 4660 1240 4680 1260
rect 4750 1240 4770 1260
rect 4840 1240 4860 1260
rect 4930 1240 4950 1260
rect 5020 1240 5040 1260
rect 5110 1240 5130 1260
rect 5200 1240 5220 1260
rect 5290 1240 5310 1260
rect 5380 1240 5400 1260
rect 5470 1240 5490 1260
rect 5560 1240 5580 1260
rect 5650 1240 5670 1260
rect 5740 1240 5760 1260
rect 5830 1240 5850 1260
rect 5920 1240 5940 1260
rect 6010 1240 6030 1260
rect 6100 1240 6120 1260
rect 6190 1240 6210 1260
rect 6280 1240 6300 1260
rect 6370 1240 6390 1260
rect 6460 1240 6480 1260
rect 6550 1240 6570 1260
rect 6640 1240 6660 1260
rect 6730 1240 6750 1260
rect 6820 1240 6840 1260
rect 6910 1240 6930 1260
rect 7000 1240 7020 1260
rect 7090 1240 7110 1260
rect 7180 1240 7200 1260
rect 7270 1240 7290 1260
rect 7360 1240 7380 1260
rect 7450 1240 7470 1260
rect 7540 1240 7560 1260
rect 7630 1240 7650 1260
rect 7720 1240 7740 1260
rect 7810 1240 7830 1260
rect 7900 1240 7920 1260
rect 7990 1240 8010 1260
rect 8080 1240 8100 1260
rect 8170 1240 8190 1260
rect 8260 1240 8280 1260
rect 8350 1240 8370 1260
rect 8440 1240 8460 1260
rect 8530 1240 8550 1260
rect 8620 1240 8640 1260
rect 8710 1240 8730 1260
rect 8800 1240 8820 1260
rect 8890 1240 8910 1260
rect 8980 1240 9000 1260
rect 9070 1240 9090 1260
rect 9160 1240 9180 1260
rect 9250 1240 9270 1260
rect 9340 1240 9360 1260
rect 9430 1240 9450 1260
rect 9520 1240 9540 1260
rect 9610 1240 9630 1260
rect 9700 1240 9720 1260
rect 9790 1240 9810 1260
rect 9880 1240 9900 1260
rect 9970 1240 9990 1260
rect 10060 1240 10080 1260
rect 10150 1240 10170 1260
rect 10240 1240 10260 1260
rect 10330 1240 10350 1260
rect 10420 1240 10440 1260
rect 10510 1240 10530 1260
rect 10600 1240 10620 1260
rect 10690 1240 10710 1260
rect 10780 1240 10800 1260
rect 10870 1240 10890 1260
rect 10960 1240 10980 1260
rect 11050 1240 11070 1260
rect 11140 1240 11160 1260
rect -295 580 -275 600
rect -205 580 -185 600
rect -115 580 -95 600
rect -25 580 -5 600
rect 65 580 85 600
rect 155 580 175 600
rect 245 580 265 600
rect 335 580 355 600
rect 425 580 445 600
rect 515 580 535 600
rect 605 580 625 600
rect 695 580 715 600
rect 785 580 805 600
rect 875 580 895 600
rect 965 580 985 600
rect 1055 580 1075 600
rect 1145 580 1165 600
rect 1235 580 1255 600
rect 1325 580 1345 600
rect 1415 580 1435 600
rect 1505 580 1525 600
rect 1595 580 1615 600
rect 1685 580 1705 600
rect 1775 580 1795 600
rect 1865 580 1885 600
rect 1955 580 1975 600
rect 2045 580 2065 600
rect 2135 580 2155 600
rect 2225 580 2245 600
rect 2315 580 2335 600
rect 2405 580 2425 600
rect 2495 580 2515 600
rect 2585 580 2605 600
rect 2675 580 2695 600
rect 2765 580 2785 600
rect 2855 580 2875 600
rect 2945 580 2965 600
rect 3035 580 3055 600
rect 3125 580 3145 600
rect 3215 580 3235 600
rect 3305 580 3325 600
rect 3395 580 3415 600
rect 3485 580 3505 600
rect 3575 580 3595 600
rect 3665 580 3685 600
rect 3755 580 3775 600
rect 3845 580 3865 600
rect 3935 580 3955 600
rect 4025 580 4045 600
rect 4115 580 4135 600
rect 4205 580 4225 600
rect 4295 580 4315 600
rect 4385 580 4405 600
rect 4475 580 4495 600
rect 4565 580 4585 600
rect 4655 580 4675 600
rect 4745 580 4765 600
rect 4835 580 4855 600
rect 4925 580 4945 600
rect 5015 580 5035 600
rect 5105 580 5125 600
rect 5195 580 5215 600
rect 5285 580 5305 600
rect 5375 580 5395 600
rect 5465 580 5485 600
rect 5555 580 5575 600
rect 5645 580 5665 600
rect 5735 580 5755 600
rect 5825 580 5845 600
rect 5915 580 5935 600
rect 6005 580 6025 600
rect 6095 580 6115 600
rect 6185 580 6205 600
rect 6275 580 6295 600
rect 6365 580 6385 600
rect 6455 580 6475 600
rect 6545 580 6565 600
rect 6635 580 6655 600
rect 6725 580 6745 600
rect 6815 580 6835 600
rect 6905 580 6925 600
rect 6995 580 7015 600
rect 7085 580 7105 600
rect 7175 580 7195 600
rect 7265 580 7285 600
rect 7355 580 7375 600
rect 7445 580 7465 600
rect 7535 580 7555 600
rect 7625 580 7645 600
rect 7715 580 7735 600
rect 7810 580 7830 600
rect 7900 580 7920 600
rect 7990 580 8010 600
rect 8080 580 8100 600
rect 8170 580 8190 600
rect 8260 580 8280 600
rect 8350 580 8370 600
rect 8440 580 8460 600
rect 8530 580 8550 600
rect 8620 580 8640 600
rect 8710 580 8730 600
rect 8800 580 8820 600
rect 8890 580 8910 600
rect 8980 580 9000 600
rect 9070 580 9090 600
rect 9160 580 9180 600
rect 9250 580 9270 600
rect 9340 580 9360 600
rect 9430 580 9450 600
rect 9520 580 9540 600
rect 9610 580 9630 600
rect 9700 580 9720 600
rect 9790 580 9810 600
rect 9880 580 9900 600
rect 9970 580 9990 600
rect 10060 580 10080 600
rect 10150 580 10170 600
rect 10240 580 10260 600
rect 10330 580 10350 600
rect 10420 580 10440 600
rect 10510 580 10530 600
rect 10600 580 10620 600
rect 10690 580 10710 600
rect 10780 580 10800 600
rect 10870 580 10890 600
rect 10960 580 10980 600
rect 11050 580 11070 600
rect 11140 580 11160 600
rect -295 220 -275 240
rect -205 220 -185 240
rect -115 220 -95 240
rect -25 220 -5 240
rect 65 220 85 240
rect 155 220 175 240
rect 245 220 265 240
rect 335 220 355 240
rect 425 220 445 240
rect 515 220 535 240
rect 605 220 625 240
rect 695 220 715 240
rect 785 220 805 240
rect 875 220 895 240
rect 965 220 985 240
rect 1055 220 1075 240
rect 1145 220 1165 240
rect 1235 220 1255 240
rect 1325 220 1345 240
rect 1415 220 1435 240
rect 1505 220 1525 240
rect 1595 220 1615 240
rect 1685 220 1705 240
rect 1775 220 1795 240
rect 1865 220 1885 240
rect 1955 220 1975 240
rect 2045 220 2065 240
rect 2135 220 2155 240
rect 2225 220 2245 240
rect 2315 220 2335 240
rect 2405 220 2425 240
rect 2495 220 2515 240
rect 2585 220 2605 240
rect 2675 220 2695 240
rect 2765 220 2785 240
rect 2855 220 2875 240
rect 2945 220 2965 240
rect 3035 220 3055 240
rect 3125 220 3145 240
rect 3215 220 3235 240
rect 3305 220 3325 240
rect 3395 220 3415 240
rect 3485 220 3505 240
rect 3575 220 3595 240
rect 3665 220 3685 240
rect 3755 220 3775 240
rect 3845 220 3865 240
rect 3935 220 3955 240
rect 4025 220 4045 240
rect 4115 220 4135 240
rect 4205 220 4225 240
rect 4295 220 4315 240
rect 4385 220 4405 240
rect 4475 220 4495 240
rect 4565 220 4585 240
rect 4655 220 4675 240
rect 4745 220 4765 240
rect 4835 220 4855 240
rect 4925 220 4945 240
rect 5015 220 5035 240
rect 5105 220 5125 240
rect 5195 220 5215 240
rect 5285 220 5305 240
rect 5375 220 5395 240
rect 5465 220 5485 240
rect 5555 220 5575 240
rect 5645 220 5665 240
rect 5735 220 5755 240
rect 5825 220 5845 240
rect 5915 220 5935 240
rect 6005 220 6025 240
rect 6095 220 6115 240
rect 6185 220 6205 240
rect 6275 220 6295 240
rect 6365 220 6385 240
rect 6455 220 6475 240
rect 6545 220 6565 240
rect 6635 220 6655 240
rect 6725 220 6745 240
rect 6815 220 6835 240
rect 6905 220 6925 240
rect 6995 220 7015 240
rect 7085 220 7105 240
rect 7175 220 7195 240
rect 7265 220 7285 240
rect 7355 220 7375 240
rect 7445 220 7465 240
rect 7535 220 7555 240
rect 7625 220 7645 240
rect 7715 220 7735 240
rect 7810 220 7830 240
rect 7900 220 7920 240
rect 7990 220 8010 240
rect 8080 220 8100 240
rect 8170 220 8190 240
rect 8260 220 8280 240
rect 8350 220 8370 240
rect 8440 220 8460 240
rect 8530 220 8550 240
rect 8620 220 8640 240
rect 8710 220 8730 240
rect 8800 220 8820 240
rect 8890 220 8910 240
rect 8980 220 9000 240
rect 9070 220 9090 240
rect 9160 220 9180 240
rect 9250 220 9270 240
rect 9340 220 9360 240
rect 9430 220 9450 240
rect 9520 220 9540 240
rect 9610 220 9630 240
rect 9700 220 9720 240
rect 9790 220 9810 240
rect 9880 220 9900 240
rect 9970 220 9990 240
rect 10060 220 10080 240
rect 10150 220 10170 240
rect 10240 220 10260 240
rect 10330 220 10350 240
rect 10420 220 10440 240
rect 10510 220 10530 240
rect 10600 220 10620 240
rect 10690 220 10710 240
rect 10780 220 10800 240
rect 10870 220 10890 240
rect 10960 220 10980 240
rect 11050 220 11070 240
rect 11140 220 11160 240
rect -295 0 -275 20
rect -205 0 -185 20
rect -115 0 -95 20
rect -25 0 -5 20
rect 65 0 85 20
rect 155 0 175 20
rect 245 0 265 20
rect 335 0 355 20
rect 425 0 445 20
rect 515 0 535 20
rect 605 0 625 20
rect 695 0 715 20
rect 785 0 805 20
rect 875 0 895 20
rect 965 0 985 20
rect 1055 0 1075 20
rect 1145 0 1165 20
rect 1235 0 1255 20
rect 1325 0 1345 20
rect 1415 0 1435 20
rect 1505 0 1525 20
rect 1595 0 1615 20
rect 1685 0 1705 20
rect 1775 0 1795 20
rect 1865 0 1885 20
rect 1955 0 1975 20
rect 2045 0 2065 20
rect 2135 0 2155 20
rect 2225 0 2245 20
rect 2315 0 2335 20
rect 2405 0 2425 20
rect 2495 0 2515 20
rect 2585 0 2605 20
rect 2675 0 2695 20
rect 2765 0 2785 20
rect 2855 0 2875 20
rect 2945 0 2965 20
rect 3035 0 3055 20
rect 3125 0 3145 20
rect 3215 0 3235 20
rect 3305 0 3325 20
rect 3395 0 3415 20
rect 3485 0 3505 20
rect 3575 0 3595 20
rect 3665 0 3685 20
rect 3755 0 3775 20
rect 3845 0 3865 20
rect 3935 0 3955 20
rect 4025 0 4045 20
rect 4115 0 4135 20
rect 4205 0 4225 20
rect 4295 0 4315 20
rect 4385 0 4405 20
rect 4475 0 4495 20
rect 4565 0 4585 20
rect 4655 0 4675 20
rect 4745 0 4765 20
rect 4835 0 4855 20
rect 4925 0 4945 20
rect 5015 0 5035 20
rect 5105 0 5125 20
rect 5195 0 5215 20
rect 5285 0 5305 20
rect 5375 0 5395 20
rect 5465 0 5485 20
rect 5555 0 5575 20
rect 5645 0 5665 20
rect 5735 0 5755 20
rect 5825 0 5845 20
rect 5915 0 5935 20
rect 6005 0 6025 20
rect 6095 0 6115 20
rect 6185 0 6205 20
rect 6275 0 6295 20
rect 6365 0 6385 20
rect 6455 0 6475 20
rect 6545 0 6565 20
rect 6635 0 6655 20
rect 6725 0 6745 20
rect 6815 0 6835 20
rect 6905 0 6925 20
rect 6995 0 7015 20
rect 7085 0 7105 20
rect 7175 0 7195 20
rect 7265 0 7285 20
rect 7355 0 7375 20
rect 7445 0 7465 20
rect 7535 0 7555 20
rect 7625 0 7645 20
rect 7715 0 7735 20
rect 7810 0 7830 20
rect 7900 0 7920 20
rect 7990 0 8010 20
rect 8080 0 8100 20
rect 8170 0 8190 20
rect 8260 0 8280 20
rect 8350 0 8370 20
rect 8440 0 8460 20
rect 8530 0 8550 20
rect 8620 0 8640 20
rect 8710 0 8730 20
rect 8800 0 8820 20
rect 8890 0 8910 20
rect 8980 0 9000 20
rect 9070 0 9090 20
rect 9160 0 9180 20
rect 9250 0 9270 20
rect 9340 0 9360 20
rect 9430 0 9450 20
rect 9520 0 9540 20
rect 9610 0 9630 20
rect 9700 0 9720 20
rect 9790 0 9810 20
rect 9880 0 9900 20
rect 9970 0 9990 20
rect 10060 0 10080 20
rect 10150 0 10170 20
rect 10240 0 10260 20
rect 10330 0 10350 20
rect 10420 0 10440 20
rect 10510 0 10530 20
rect 10600 0 10620 20
rect 10690 0 10710 20
rect 10780 0 10800 20
rect 10870 0 10890 20
rect 10960 0 10980 20
rect 11050 0 11070 20
rect 11140 0 11160 20
<< nsubdiffcont >>
rect -295 1160 -275 1180
rect -205 1160 -185 1180
rect -115 1160 -95 1180
rect -25 1160 -5 1180
rect 65 1160 85 1180
rect 155 1160 175 1180
rect 245 1160 265 1180
rect 335 1160 355 1180
rect 425 1160 445 1180
rect 515 1160 535 1180
rect 605 1160 625 1180
rect 695 1160 715 1180
rect 785 1160 805 1180
rect 875 1160 895 1180
rect 965 1160 985 1180
rect 1055 1160 1075 1180
rect 1145 1160 1165 1180
rect 1235 1160 1255 1180
rect 1325 1160 1345 1180
rect 1415 1160 1435 1180
rect 1505 1160 1525 1180
rect 1595 1160 1615 1180
rect 1685 1160 1705 1180
rect 1775 1160 1795 1180
rect 1865 1160 1885 1180
rect 1955 1160 1975 1180
rect 2045 1160 2065 1180
rect 2135 1160 2155 1180
rect 2225 1160 2245 1180
rect 2315 1160 2335 1180
rect 2405 1160 2425 1180
rect 2495 1160 2515 1180
rect 2585 1160 2605 1180
rect 2675 1160 2695 1180
rect 2765 1160 2785 1180
rect 2855 1160 2875 1180
rect 2945 1160 2965 1180
rect 3035 1160 3055 1180
rect 3130 1160 3150 1180
rect 3220 1160 3240 1180
rect 3310 1160 3330 1180
rect 3400 1160 3420 1180
rect 3490 1160 3510 1180
rect 3580 1160 3600 1180
rect 3670 1160 3690 1180
rect 3760 1160 3780 1180
rect 3850 1160 3870 1180
rect 3940 1160 3960 1180
rect 4030 1160 4050 1180
rect 4120 1160 4140 1180
rect 4210 1160 4230 1180
rect 4300 1160 4320 1180
rect 4390 1160 4410 1180
rect 4480 1160 4500 1180
rect 4570 1160 4590 1180
rect 4660 1160 4680 1180
rect 4750 1160 4770 1180
rect 4840 1160 4860 1180
rect 4930 1160 4950 1180
rect 5020 1160 5040 1180
rect 5110 1160 5130 1180
rect 5200 1160 5220 1180
rect 5290 1160 5310 1180
rect 5380 1160 5400 1180
rect 5470 1160 5490 1180
rect 5560 1160 5580 1180
rect 5650 1160 5670 1180
rect 5740 1160 5760 1180
rect 5830 1160 5850 1180
rect 5920 1160 5940 1180
rect 6010 1160 6030 1180
rect 6100 1160 6120 1180
rect 6190 1160 6210 1180
rect 6280 1160 6300 1180
rect 6370 1160 6390 1180
rect 6460 1160 6480 1180
rect 6550 1160 6570 1180
rect 6640 1160 6660 1180
rect 6730 1160 6750 1180
rect 6820 1160 6840 1180
rect 6910 1160 6930 1180
rect 7000 1160 7020 1180
rect 7090 1160 7110 1180
rect 7180 1160 7200 1180
rect 7270 1160 7290 1180
rect 7360 1160 7380 1180
rect 7450 1160 7470 1180
rect 7540 1160 7560 1180
rect 7630 1160 7650 1180
rect 7720 1160 7740 1180
rect 7810 1160 7830 1180
rect 7900 1160 7920 1180
rect 7990 1160 8010 1180
rect 8080 1160 8100 1180
rect 8170 1160 8190 1180
rect 8260 1160 8280 1180
rect 8350 1160 8370 1180
rect 8440 1160 8460 1180
rect 8530 1160 8550 1180
rect 8620 1160 8640 1180
rect 8710 1160 8730 1180
rect 8800 1160 8820 1180
rect 8890 1160 8910 1180
rect 8980 1160 9000 1180
rect 9070 1160 9090 1180
rect 9160 1160 9180 1180
rect 9250 1160 9270 1180
rect 9340 1160 9360 1180
rect 9430 1160 9450 1180
rect 9520 1160 9540 1180
rect 9610 1160 9630 1180
rect 9700 1160 9720 1180
rect 9790 1160 9810 1180
rect 9880 1160 9900 1180
rect 9970 1160 9990 1180
rect 10060 1160 10080 1180
rect 10150 1160 10170 1180
rect 10240 1160 10260 1180
rect 10330 1160 10350 1180
rect 10420 1160 10440 1180
rect 10510 1160 10530 1180
rect 10600 1160 10620 1180
rect 10690 1160 10710 1180
rect 10780 1160 10800 1180
rect 10870 1160 10890 1180
rect 10960 1160 10980 1180
rect 11050 1160 11070 1180
rect 11140 1160 11160 1180
rect -295 940 -275 960
rect -205 940 -185 960
rect -115 940 -95 960
rect -25 940 -5 960
rect 65 940 85 960
rect 155 940 175 960
rect 245 940 265 960
rect 335 940 355 960
rect 425 940 445 960
rect 515 940 535 960
rect 605 940 625 960
rect 695 940 715 960
rect 785 940 805 960
rect 875 940 895 960
rect 965 940 985 960
rect 1055 940 1075 960
rect 1145 940 1165 960
rect 1235 940 1255 960
rect 1325 940 1345 960
rect 1415 940 1435 960
rect 1505 940 1525 960
rect 1595 940 1615 960
rect 1685 940 1705 960
rect 1775 940 1795 960
rect 1865 940 1885 960
rect 1955 940 1975 960
rect 2045 940 2065 960
rect 2135 940 2155 960
rect 2225 940 2245 960
rect 2315 940 2335 960
rect 2405 940 2425 960
rect 2495 940 2515 960
rect 2585 940 2605 960
rect 2675 940 2695 960
rect 2765 940 2785 960
rect 2855 940 2875 960
rect 2945 940 2965 960
rect 3035 940 3055 960
rect 3130 940 3150 960
rect 3220 940 3240 960
rect 3310 940 3330 960
rect 3400 940 3420 960
rect 3490 940 3510 960
rect 3580 940 3600 960
rect 3670 940 3690 960
rect 3760 940 3780 960
rect 3850 940 3870 960
rect 3940 940 3960 960
rect 4030 940 4050 960
rect 4120 940 4140 960
rect 4210 940 4230 960
rect 4300 940 4320 960
rect 4390 940 4410 960
rect 4480 940 4500 960
rect 4570 940 4590 960
rect 4660 940 4680 960
rect 4750 940 4770 960
rect 4840 940 4860 960
rect 4930 940 4950 960
rect 5020 940 5040 960
rect 5110 940 5130 960
rect 5200 940 5220 960
rect 5290 940 5310 960
rect 5380 940 5400 960
rect 5470 940 5490 960
rect 5560 940 5580 960
rect 5650 940 5670 960
rect 5740 940 5760 960
rect 5830 940 5850 960
rect 5920 940 5940 960
rect 6010 940 6030 960
rect 6100 940 6120 960
rect 6190 940 6210 960
rect 6280 940 6300 960
rect 6370 940 6390 960
rect 6460 940 6480 960
rect 6550 940 6570 960
rect 6640 940 6660 960
rect 6730 940 6750 960
rect 6820 940 6840 960
rect 6910 940 6930 960
rect 7000 940 7020 960
rect 7090 940 7110 960
rect 7180 940 7200 960
rect 7270 940 7290 960
rect 7360 940 7380 960
rect 7450 940 7470 960
rect 7540 940 7560 960
rect 7630 940 7650 960
rect 7720 940 7740 960
rect 7810 940 7830 960
rect 7900 940 7920 960
rect 7990 940 8010 960
rect 8080 940 8100 960
rect 8170 940 8190 960
rect 8260 940 8280 960
rect 8350 940 8370 960
rect 8440 940 8460 960
rect 8530 940 8550 960
rect 8620 940 8640 960
rect 8710 940 8730 960
rect 8800 940 8820 960
rect 8890 940 8910 960
rect 8980 940 9000 960
rect 9070 940 9090 960
rect 9160 940 9180 960
rect 9250 940 9270 960
rect 9340 940 9360 960
rect 9430 940 9450 960
rect 9520 940 9540 960
rect 9610 940 9630 960
rect 9700 940 9720 960
rect 9790 940 9810 960
rect 9880 940 9900 960
rect 9970 940 9990 960
rect 10060 940 10080 960
rect 10150 940 10170 960
rect 10240 940 10260 960
rect 10330 940 10350 960
rect 10420 940 10440 960
rect 10510 940 10530 960
rect 10600 940 10620 960
rect 10690 940 10710 960
rect 10780 940 10800 960
rect 10870 940 10890 960
rect 10960 940 10980 960
rect 11050 940 11070 960
rect 11140 940 11160 960
rect -295 880 -275 900
rect -205 880 -185 900
rect -115 880 -95 900
rect -25 880 -5 900
rect 65 880 85 900
rect 155 880 175 900
rect 245 880 265 900
rect 335 880 355 900
rect 425 880 445 900
rect 515 880 535 900
rect 605 880 625 900
rect 695 880 715 900
rect 785 880 805 900
rect 875 880 895 900
rect 965 880 985 900
rect 1055 880 1075 900
rect 1145 880 1165 900
rect 1235 880 1255 900
rect 1325 880 1345 900
rect 1415 880 1435 900
rect 1505 880 1525 900
rect 1595 880 1615 900
rect 1685 880 1705 900
rect 1775 880 1795 900
rect 1865 880 1885 900
rect 1955 880 1975 900
rect 2045 880 2065 900
rect 2135 880 2155 900
rect 2225 880 2245 900
rect 2315 880 2335 900
rect 2405 880 2425 900
rect 2495 880 2515 900
rect 2585 880 2605 900
rect 2675 880 2695 900
rect 2765 880 2785 900
rect 2855 880 2875 900
rect 2945 880 2965 900
rect 3035 880 3055 900
rect 3125 880 3145 900
rect 3215 880 3235 900
rect 3305 880 3325 900
rect 3395 880 3415 900
rect 3485 880 3505 900
rect 3575 880 3595 900
rect 3665 880 3685 900
rect 3755 880 3775 900
rect 3845 880 3865 900
rect 3935 880 3955 900
rect 4025 880 4045 900
rect 4115 880 4135 900
rect 4205 880 4225 900
rect 4295 880 4315 900
rect 4385 880 4405 900
rect 4475 880 4495 900
rect 4565 880 4585 900
rect 4655 880 4675 900
rect 4745 880 4765 900
rect 4835 880 4855 900
rect 4925 880 4945 900
rect 5015 880 5035 900
rect 5105 880 5125 900
rect 5195 880 5215 900
rect 5285 880 5305 900
rect 5375 880 5395 900
rect 5465 880 5485 900
rect 5555 880 5575 900
rect 5645 880 5665 900
rect 5735 880 5755 900
rect 5825 880 5845 900
rect 5915 880 5935 900
rect 6005 880 6025 900
rect 6095 880 6115 900
rect 6185 880 6205 900
rect 6275 880 6295 900
rect 6365 880 6385 900
rect 6455 880 6475 900
rect 6545 880 6565 900
rect 6635 880 6655 900
rect 6725 880 6745 900
rect 6815 880 6835 900
rect 6905 880 6925 900
rect 6995 880 7015 900
rect 7085 880 7105 900
rect 7175 880 7195 900
rect 7265 880 7285 900
rect 7355 880 7375 900
rect 7445 880 7465 900
rect 7535 880 7555 900
rect 7625 880 7645 900
rect 7715 880 7735 900
rect 7810 880 7830 900
rect 7900 880 7920 900
rect 7990 880 8010 900
rect 8080 880 8100 900
rect 8170 880 8190 900
rect 8260 880 8280 900
rect 8350 880 8370 900
rect 8440 880 8460 900
rect 8530 880 8550 900
rect 8620 880 8640 900
rect 8710 880 8730 900
rect 8800 880 8820 900
rect 8890 880 8910 900
rect 8980 880 9000 900
rect 9070 880 9090 900
rect 9160 880 9180 900
rect 9250 880 9270 900
rect 9340 880 9360 900
rect 9430 880 9450 900
rect 9520 880 9540 900
rect 9610 880 9630 900
rect 9700 880 9720 900
rect 9790 880 9810 900
rect 9880 880 9900 900
rect 9970 880 9990 900
rect 10060 880 10080 900
rect 10150 880 10170 900
rect 10240 880 10260 900
rect 10330 880 10350 900
rect 10420 880 10440 900
rect 10510 880 10530 900
rect 10600 880 10620 900
rect 10690 880 10710 900
rect 10780 880 10800 900
rect 10870 880 10890 900
rect 10960 880 10980 900
rect 11050 880 11070 900
rect 11140 880 11160 900
rect -295 660 -275 680
rect -205 660 -185 680
rect -115 660 -95 680
rect -25 660 -5 680
rect 65 660 85 680
rect 155 660 175 680
rect 245 660 265 680
rect 335 660 355 680
rect 425 660 445 680
rect 515 660 535 680
rect 605 660 625 680
rect 695 660 715 680
rect 785 660 805 680
rect 875 660 895 680
rect 965 660 985 680
rect 1055 660 1075 680
rect 1145 660 1165 680
rect 1235 660 1255 680
rect 1325 660 1345 680
rect 1415 660 1435 680
rect 1505 660 1525 680
rect 1595 660 1615 680
rect 1685 660 1705 680
rect 1775 660 1795 680
rect 1865 660 1885 680
rect 1955 660 1975 680
rect 2045 660 2065 680
rect 2135 660 2155 680
rect 2225 660 2245 680
rect 2315 660 2335 680
rect 2405 660 2425 680
rect 2495 660 2515 680
rect 2585 660 2605 680
rect 2675 660 2695 680
rect 2765 660 2785 680
rect 2855 660 2875 680
rect 2945 660 2965 680
rect 3035 660 3055 680
rect 3125 660 3145 680
rect 3215 660 3235 680
rect 3305 660 3325 680
rect 3395 660 3415 680
rect 3485 660 3505 680
rect 3575 660 3595 680
rect 3665 660 3685 680
rect 3755 660 3775 680
rect 3845 660 3865 680
rect 3935 660 3955 680
rect 4025 660 4045 680
rect 4115 660 4135 680
rect 4205 660 4225 680
rect 4295 660 4315 680
rect 4385 660 4405 680
rect 4475 660 4495 680
rect 4565 660 4585 680
rect 4655 660 4675 680
rect 4745 660 4765 680
rect 4835 660 4855 680
rect 4925 660 4945 680
rect 5015 660 5035 680
rect 5105 660 5125 680
rect 5195 660 5215 680
rect 5285 660 5305 680
rect 5375 660 5395 680
rect 5465 660 5485 680
rect 5555 660 5575 680
rect 5645 660 5665 680
rect 5735 660 5755 680
rect 5825 660 5845 680
rect 5915 660 5935 680
rect 6005 660 6025 680
rect 6095 660 6115 680
rect 6185 660 6205 680
rect 6275 660 6295 680
rect 6365 660 6385 680
rect 6455 660 6475 680
rect 6545 660 6565 680
rect 6635 660 6655 680
rect 6725 660 6745 680
rect 6815 660 6835 680
rect 6905 660 6925 680
rect 6995 660 7015 680
rect 7085 660 7105 680
rect 7175 660 7195 680
rect 7265 660 7285 680
rect 7355 660 7375 680
rect 7445 660 7465 680
rect 7535 660 7555 680
rect 7625 660 7645 680
rect 7715 660 7735 680
rect 7810 660 7830 680
rect 7900 660 7920 680
rect 7990 660 8010 680
rect 8080 660 8100 680
rect 8170 660 8190 680
rect 8260 660 8280 680
rect 8350 660 8370 680
rect 8440 660 8460 680
rect 8530 660 8550 680
rect 8620 660 8640 680
rect 8710 660 8730 680
rect 8800 660 8820 680
rect 8890 660 8910 680
rect 8980 660 9000 680
rect 9070 660 9090 680
rect 9160 660 9180 680
rect 9250 660 9270 680
rect 9340 660 9360 680
rect 9430 660 9450 680
rect 9520 660 9540 680
rect 9610 660 9630 680
rect 9700 660 9720 680
rect 9790 660 9810 680
rect 9880 660 9900 680
rect 9970 660 9990 680
rect 10060 660 10080 680
rect 10150 660 10170 680
rect 10240 660 10260 680
rect 10330 660 10350 680
rect 10420 660 10440 680
rect 10510 660 10530 680
rect 10600 660 10620 680
rect 10690 660 10710 680
rect 10780 660 10800 680
rect 10870 660 10890 680
rect 10960 660 10980 680
rect 11050 660 11070 680
rect 11140 660 11160 680
<< poly >>
rect -310 1790 -260 1805
rect -220 1790 -170 1805
rect -130 1790 -80 1805
rect -40 1790 10 1805
rect 50 1790 100 1805
rect 140 1790 190 1805
rect 230 1790 280 1805
rect 320 1790 370 1805
rect 410 1790 460 1805
rect 500 1790 550 1805
rect 590 1790 640 1805
rect 680 1790 730 1805
rect 770 1790 820 1805
rect 860 1790 910 1805
rect 950 1790 1000 1805
rect 1040 1790 1090 1805
rect 1130 1790 1180 1805
rect 1220 1790 1270 1805
rect 1310 1790 1360 1805
rect 1400 1790 1450 1805
rect 1490 1790 1540 1805
rect 1580 1790 1630 1805
rect 1670 1790 1720 1805
rect 1760 1790 1810 1805
rect 1850 1790 1900 1805
rect 1940 1790 1990 1805
rect 2030 1790 2080 1805
rect 2120 1790 2170 1805
rect 2210 1790 2260 1805
rect 2300 1790 2350 1805
rect 2390 1790 2440 1805
rect 2480 1790 2530 1805
rect 2570 1790 2620 1805
rect 2660 1790 2710 1805
rect 2750 1790 2800 1805
rect 2840 1790 2890 1805
rect 2930 1790 2980 1805
rect 3020 1790 3070 1805
rect 3115 1790 3165 1805
rect 3205 1790 3255 1805
rect 3295 1790 3345 1805
rect 3385 1790 3435 1805
rect 3475 1790 3525 1805
rect 3565 1790 3615 1805
rect 3655 1790 3705 1805
rect 3745 1790 3795 1805
rect 3835 1790 3885 1805
rect 3925 1790 3975 1805
rect 4015 1790 4065 1805
rect 4105 1790 4155 1805
rect 4195 1790 4245 1805
rect 4285 1790 4335 1805
rect 4375 1790 4425 1805
rect 4465 1790 4515 1805
rect 4555 1790 4605 1805
rect 4645 1790 4695 1805
rect 4735 1790 4785 1805
rect 4825 1790 4875 1805
rect 4915 1790 4965 1805
rect 5005 1790 5055 1805
rect 5095 1790 5145 1805
rect 5185 1790 5235 1805
rect 5275 1790 5325 1805
rect 5365 1790 5415 1805
rect 5455 1790 5505 1805
rect 5545 1790 5595 1805
rect 5635 1790 5685 1805
rect 5725 1790 5775 1805
rect 5815 1790 5865 1805
rect 5905 1790 5955 1805
rect 5995 1790 6045 1805
rect 6085 1790 6135 1805
rect 6175 1790 6225 1805
rect 6265 1790 6315 1805
rect 6355 1790 6405 1805
rect 6445 1790 6495 1805
rect 6535 1790 6585 1805
rect 6625 1790 6675 1805
rect 6715 1790 6765 1805
rect 6805 1790 6855 1805
rect 6895 1790 6945 1805
rect 6985 1790 7035 1805
rect 7075 1790 7125 1805
rect 7165 1790 7215 1805
rect 7255 1790 7305 1805
rect 7345 1790 7395 1805
rect 7435 1790 7485 1805
rect 7525 1790 7575 1805
rect 7615 1790 7665 1805
rect 7705 1790 7755 1805
rect 7795 1790 7845 1805
rect 7885 1790 7935 1805
rect 7975 1790 8025 1805
rect 8065 1790 8115 1805
rect 8155 1790 8205 1805
rect 8245 1790 8295 1805
rect 8335 1790 8385 1805
rect 8425 1790 8475 1805
rect 8515 1790 8565 1805
rect 8605 1790 8655 1805
rect 8695 1790 8745 1805
rect 8785 1790 8835 1805
rect 8875 1790 8925 1805
rect 8965 1790 9015 1805
rect 9055 1790 9105 1805
rect 9145 1790 9195 1805
rect 9235 1790 9285 1805
rect 9325 1790 9375 1805
rect 9415 1790 9465 1805
rect 9505 1790 9555 1805
rect 9595 1790 9645 1805
rect 9685 1790 9735 1805
rect 9775 1790 9825 1805
rect 9865 1790 9915 1805
rect 9955 1790 10005 1805
rect 10045 1790 10095 1805
rect 10135 1790 10185 1805
rect 10225 1790 10275 1805
rect 10315 1790 10365 1805
rect 10405 1790 10455 1805
rect 10495 1790 10545 1805
rect 10585 1790 10635 1805
rect 10675 1790 10725 1805
rect 10765 1790 10815 1805
rect 10855 1790 10905 1805
rect 10945 1790 10995 1805
rect 11035 1790 11085 1805
rect 11125 1790 11175 1805
rect -310 1670 -260 1690
rect -220 1670 -170 1690
rect -310 1665 -170 1670
rect -310 1645 -295 1665
rect -275 1645 -205 1665
rect -185 1645 -170 1665
rect -310 1640 -170 1645
rect -130 1670 -80 1690
rect -40 1670 10 1690
rect -130 1665 10 1670
rect -130 1645 -115 1665
rect -95 1645 -25 1665
rect -5 1645 10 1665
rect -130 1640 10 1645
rect 50 1670 100 1690
rect 140 1670 190 1690
rect 50 1665 190 1670
rect 50 1645 65 1665
rect 85 1645 155 1665
rect 175 1645 190 1665
rect 50 1640 190 1645
rect 230 1670 280 1690
rect 320 1670 370 1690
rect 230 1665 370 1670
rect 230 1645 245 1665
rect 265 1645 335 1665
rect 355 1645 370 1665
rect 230 1640 370 1645
rect 410 1670 460 1690
rect 500 1670 550 1690
rect 410 1665 550 1670
rect 410 1645 425 1665
rect 445 1645 515 1665
rect 535 1645 550 1665
rect 410 1640 550 1645
rect 590 1670 640 1690
rect 680 1670 730 1690
rect 590 1665 730 1670
rect 590 1645 605 1665
rect 625 1645 695 1665
rect 715 1645 730 1665
rect 590 1640 730 1645
rect 770 1670 820 1690
rect 860 1670 910 1690
rect 770 1665 910 1670
rect 770 1645 785 1665
rect 805 1645 875 1665
rect 895 1645 910 1665
rect 770 1640 910 1645
rect 950 1670 1000 1690
rect 1040 1670 1090 1690
rect 950 1665 1090 1670
rect 950 1645 965 1665
rect 985 1645 1055 1665
rect 1075 1645 1090 1665
rect 950 1640 1090 1645
rect 1130 1670 1180 1690
rect 1220 1670 1270 1690
rect 1130 1665 1270 1670
rect 1130 1645 1145 1665
rect 1165 1645 1235 1665
rect 1255 1645 1270 1665
rect 1130 1640 1270 1645
rect 1310 1670 1360 1690
rect 1400 1670 1450 1690
rect 1310 1665 1450 1670
rect 1310 1645 1325 1665
rect 1345 1645 1415 1665
rect 1435 1645 1450 1665
rect 1310 1640 1450 1645
rect 1490 1670 1540 1690
rect 1580 1670 1630 1690
rect 1490 1665 1630 1670
rect 1490 1645 1505 1665
rect 1525 1645 1595 1665
rect 1615 1645 1630 1665
rect 1490 1640 1630 1645
rect 1670 1670 1720 1690
rect 1760 1670 1810 1690
rect 1670 1665 1810 1670
rect 1670 1645 1685 1665
rect 1705 1645 1775 1665
rect 1795 1645 1810 1665
rect 1670 1640 1810 1645
rect 1850 1670 1900 1690
rect 1940 1670 1990 1690
rect 1850 1665 1990 1670
rect 1850 1645 1865 1665
rect 1885 1645 1955 1665
rect 1975 1645 1990 1665
rect 1850 1640 1990 1645
rect 2030 1670 2080 1690
rect 2120 1670 2170 1690
rect 2030 1665 2170 1670
rect 2030 1645 2045 1665
rect 2065 1645 2135 1665
rect 2155 1645 2170 1665
rect 2030 1640 2170 1645
rect 2210 1670 2260 1690
rect 2300 1670 2350 1690
rect 2210 1665 2350 1670
rect 2210 1645 2225 1665
rect 2245 1645 2315 1665
rect 2335 1645 2350 1665
rect 2210 1640 2350 1645
rect 2390 1670 2440 1690
rect 2480 1670 2530 1690
rect 2390 1665 2530 1670
rect 2390 1645 2405 1665
rect 2425 1645 2495 1665
rect 2515 1645 2530 1665
rect 2390 1640 2530 1645
rect 2570 1670 2620 1690
rect 2660 1670 2710 1690
rect 2570 1665 2710 1670
rect 2570 1645 2585 1665
rect 2605 1645 2675 1665
rect 2695 1645 2710 1665
rect 2570 1640 2710 1645
rect 2750 1670 2800 1690
rect 2840 1670 2890 1690
rect 2750 1665 2890 1670
rect 2750 1645 2765 1665
rect 2785 1645 2855 1665
rect 2875 1645 2890 1665
rect 2750 1640 2890 1645
rect 2930 1670 2980 1690
rect 3020 1670 3070 1690
rect 2930 1665 3070 1670
rect 2930 1645 2945 1665
rect 2965 1645 3035 1665
rect 3055 1645 3070 1665
rect 2930 1640 3070 1645
rect 3115 1670 3165 1690
rect 3205 1670 3255 1690
rect 3115 1665 3255 1670
rect 3115 1645 3130 1665
rect 3150 1645 3220 1665
rect 3240 1645 3255 1665
rect 3115 1640 3255 1645
rect 3295 1670 3345 1690
rect 3385 1670 3435 1690
rect 3295 1665 3435 1670
rect 3295 1645 3310 1665
rect 3330 1645 3400 1665
rect 3420 1645 3435 1665
rect 3295 1640 3435 1645
rect 3475 1670 3525 1690
rect 3565 1670 3615 1690
rect 3475 1665 3615 1670
rect 3475 1645 3490 1665
rect 3510 1645 3580 1665
rect 3600 1645 3615 1665
rect 3475 1640 3615 1645
rect 3655 1670 3705 1690
rect 3745 1670 3795 1690
rect 3655 1665 3795 1670
rect 3655 1645 3670 1665
rect 3690 1645 3760 1665
rect 3780 1645 3795 1665
rect 3655 1640 3795 1645
rect 3835 1670 3885 1690
rect 3925 1670 3975 1690
rect 3835 1665 3975 1670
rect 3835 1645 3850 1665
rect 3870 1645 3940 1665
rect 3960 1645 3975 1665
rect 3835 1640 3975 1645
rect 4015 1670 4065 1690
rect 4105 1670 4155 1690
rect 4015 1665 4155 1670
rect 4015 1645 4030 1665
rect 4050 1645 4120 1665
rect 4140 1645 4155 1665
rect 4015 1640 4155 1645
rect 4195 1670 4245 1690
rect 4285 1670 4335 1690
rect 4195 1665 4335 1670
rect 4195 1645 4210 1665
rect 4230 1645 4300 1665
rect 4320 1645 4335 1665
rect 4195 1640 4335 1645
rect 4375 1670 4425 1690
rect 4465 1670 4515 1690
rect 4375 1665 4515 1670
rect 4375 1645 4390 1665
rect 4410 1645 4480 1665
rect 4500 1645 4515 1665
rect 4375 1640 4515 1645
rect 4555 1670 4605 1690
rect 4645 1670 4695 1690
rect 4555 1665 4695 1670
rect 4555 1645 4570 1665
rect 4590 1645 4660 1665
rect 4680 1645 4695 1665
rect 4555 1640 4695 1645
rect 4735 1670 4785 1690
rect 4825 1670 4875 1690
rect 4735 1665 4875 1670
rect 4735 1645 4750 1665
rect 4770 1645 4840 1665
rect 4860 1645 4875 1665
rect 4735 1640 4875 1645
rect 4915 1670 4965 1690
rect 5005 1670 5055 1690
rect 4915 1665 5055 1670
rect 4915 1645 4930 1665
rect 4950 1645 5020 1665
rect 5040 1645 5055 1665
rect 4915 1640 5055 1645
rect 5095 1670 5145 1690
rect 5185 1670 5235 1690
rect 5095 1665 5235 1670
rect 5095 1645 5110 1665
rect 5130 1645 5200 1665
rect 5220 1645 5235 1665
rect 5095 1640 5235 1645
rect 5275 1670 5325 1690
rect 5365 1670 5415 1690
rect 5275 1665 5415 1670
rect 5275 1645 5290 1665
rect 5310 1645 5380 1665
rect 5400 1645 5415 1665
rect 5275 1640 5415 1645
rect 5455 1670 5505 1690
rect 5545 1670 5595 1690
rect 5455 1665 5595 1670
rect 5455 1645 5470 1665
rect 5490 1645 5560 1665
rect 5580 1645 5595 1665
rect 5455 1640 5595 1645
rect 5635 1670 5685 1690
rect 5725 1670 5775 1690
rect 5635 1665 5775 1670
rect 5635 1645 5650 1665
rect 5670 1645 5740 1665
rect 5760 1645 5775 1665
rect 5635 1640 5775 1645
rect 5815 1670 5865 1690
rect 5905 1670 5955 1690
rect 5815 1665 5955 1670
rect 5815 1645 5830 1665
rect 5850 1645 5920 1665
rect 5940 1645 5955 1665
rect 5815 1640 5955 1645
rect 5995 1670 6045 1690
rect 6085 1670 6135 1690
rect 5995 1665 6135 1670
rect 5995 1645 6010 1665
rect 6030 1645 6100 1665
rect 6120 1645 6135 1665
rect 5995 1640 6135 1645
rect 6175 1670 6225 1690
rect 6265 1670 6315 1690
rect 6175 1665 6315 1670
rect 6175 1645 6190 1665
rect 6210 1645 6280 1665
rect 6300 1645 6315 1665
rect 6175 1640 6315 1645
rect 6355 1670 6405 1690
rect 6445 1670 6495 1690
rect 6355 1665 6495 1670
rect 6355 1645 6370 1665
rect 6390 1645 6460 1665
rect 6480 1645 6495 1665
rect 6355 1640 6495 1645
rect 6535 1670 6585 1690
rect 6625 1670 6675 1690
rect 6535 1665 6675 1670
rect 6535 1645 6550 1665
rect 6570 1645 6640 1665
rect 6660 1645 6675 1665
rect 6535 1640 6675 1645
rect 6715 1670 6765 1690
rect 6805 1670 6855 1690
rect 6715 1665 6855 1670
rect 6715 1645 6730 1665
rect 6750 1645 6820 1665
rect 6840 1645 6855 1665
rect 6715 1640 6855 1645
rect 6895 1670 6945 1690
rect 6985 1670 7035 1690
rect 6895 1665 7035 1670
rect 6895 1645 6910 1665
rect 6930 1645 7000 1665
rect 7020 1645 7035 1665
rect 6895 1640 7035 1645
rect 7075 1670 7125 1690
rect 7165 1670 7215 1690
rect 7075 1665 7215 1670
rect 7075 1645 7090 1665
rect 7110 1645 7180 1665
rect 7200 1645 7215 1665
rect 7075 1640 7215 1645
rect 7255 1670 7305 1690
rect 7345 1670 7395 1690
rect 7255 1665 7395 1670
rect 7255 1645 7270 1665
rect 7290 1645 7360 1665
rect 7380 1645 7395 1665
rect 7255 1640 7395 1645
rect 7435 1670 7485 1690
rect 7525 1670 7575 1690
rect 7435 1665 7575 1670
rect 7435 1645 7450 1665
rect 7470 1645 7540 1665
rect 7560 1645 7575 1665
rect 7435 1640 7575 1645
rect 7615 1670 7665 1690
rect 7705 1670 7755 1690
rect 7615 1665 7755 1670
rect 7615 1645 7630 1665
rect 7650 1645 7720 1665
rect 7740 1645 7755 1665
rect 7615 1640 7755 1645
rect 7795 1670 7845 1690
rect 7885 1670 7935 1690
rect 7795 1665 7935 1670
rect 7795 1645 7810 1665
rect 7830 1645 7900 1665
rect 7920 1645 7935 1665
rect 7795 1640 7935 1645
rect 7975 1670 8025 1690
rect 8065 1670 8115 1690
rect 7975 1665 8115 1670
rect 7975 1645 7990 1665
rect 8010 1645 8080 1665
rect 8100 1645 8115 1665
rect 7975 1640 8115 1645
rect 8155 1670 8205 1690
rect 8245 1670 8295 1690
rect 8155 1665 8295 1670
rect 8155 1645 8170 1665
rect 8190 1645 8260 1665
rect 8280 1645 8295 1665
rect 8155 1640 8295 1645
rect 8335 1670 8385 1690
rect 8425 1670 8475 1690
rect 8335 1665 8475 1670
rect 8335 1645 8350 1665
rect 8370 1645 8440 1665
rect 8460 1645 8475 1665
rect 8335 1640 8475 1645
rect 8515 1670 8565 1690
rect 8605 1670 8655 1690
rect 8515 1665 8655 1670
rect 8515 1645 8530 1665
rect 8550 1645 8620 1665
rect 8640 1645 8655 1665
rect 8515 1640 8655 1645
rect 8695 1670 8745 1690
rect 8785 1670 8835 1690
rect 8695 1665 8835 1670
rect 8695 1645 8710 1665
rect 8730 1645 8800 1665
rect 8820 1645 8835 1665
rect 8695 1640 8835 1645
rect 8875 1670 8925 1690
rect 8965 1670 9015 1690
rect 8875 1665 9015 1670
rect 8875 1645 8890 1665
rect 8910 1645 8980 1665
rect 9000 1645 9015 1665
rect 8875 1640 9015 1645
rect 9055 1670 9105 1690
rect 9145 1670 9195 1690
rect 9055 1665 9195 1670
rect 9055 1645 9070 1665
rect 9090 1645 9160 1665
rect 9180 1645 9195 1665
rect 9055 1640 9195 1645
rect 9235 1670 9285 1690
rect 9325 1670 9375 1690
rect 9235 1665 9375 1670
rect 9235 1645 9250 1665
rect 9270 1645 9340 1665
rect 9360 1645 9375 1665
rect 9235 1640 9375 1645
rect 9415 1670 9465 1690
rect 9505 1670 9555 1690
rect 9415 1665 9555 1670
rect 9415 1645 9430 1665
rect 9450 1645 9520 1665
rect 9540 1645 9555 1665
rect 9415 1640 9555 1645
rect 9595 1670 9645 1690
rect 9685 1670 9735 1690
rect 9595 1665 9735 1670
rect 9595 1645 9610 1665
rect 9630 1645 9700 1665
rect 9720 1645 9735 1665
rect 9595 1640 9735 1645
rect 9775 1670 9825 1690
rect 9865 1670 9915 1690
rect 9775 1665 9915 1670
rect 9775 1645 9790 1665
rect 9810 1645 9880 1665
rect 9900 1645 9915 1665
rect 9775 1640 9915 1645
rect 9955 1670 10005 1690
rect 10045 1670 10095 1690
rect 9955 1665 10095 1670
rect 9955 1645 9970 1665
rect 9990 1645 10060 1665
rect 10080 1645 10095 1665
rect 9955 1640 10095 1645
rect 10135 1670 10185 1690
rect 10225 1670 10275 1690
rect 10135 1665 10275 1670
rect 10135 1645 10150 1665
rect 10170 1645 10240 1665
rect 10260 1645 10275 1665
rect 10135 1640 10275 1645
rect 10315 1670 10365 1690
rect 10405 1670 10455 1690
rect 10315 1665 10455 1670
rect 10315 1645 10330 1665
rect 10350 1645 10420 1665
rect 10440 1645 10455 1665
rect 10315 1640 10455 1645
rect 10495 1670 10545 1690
rect 10585 1670 10635 1690
rect 10495 1665 10635 1670
rect 10495 1645 10510 1665
rect 10530 1645 10600 1665
rect 10620 1645 10635 1665
rect 10495 1640 10635 1645
rect 10675 1670 10725 1690
rect 10765 1670 10815 1690
rect 10675 1665 10815 1670
rect 10675 1645 10690 1665
rect 10710 1645 10780 1665
rect 10800 1645 10815 1665
rect 10675 1640 10815 1645
rect 10855 1670 10905 1690
rect 10945 1670 10995 1690
rect 10855 1665 10995 1670
rect 10855 1645 10870 1665
rect 10890 1645 10960 1665
rect 10980 1645 10995 1665
rect 10855 1640 10995 1645
rect 11035 1670 11085 1690
rect 11125 1670 11175 1690
rect 11035 1665 11175 1670
rect 11035 1645 11050 1665
rect 11070 1645 11140 1665
rect 11160 1645 11175 1665
rect 11035 1640 11175 1645
rect -310 1135 -170 1140
rect -310 1115 -295 1135
rect -275 1115 -205 1135
rect -185 1115 -170 1135
rect -310 1110 -170 1115
rect -310 1090 -260 1110
rect -220 1090 -170 1110
rect -130 1135 10 1140
rect -130 1115 -115 1135
rect -95 1115 -25 1135
rect -5 1115 10 1135
rect -130 1110 10 1115
rect -130 1090 -80 1110
rect -40 1090 10 1110
rect 50 1135 190 1140
rect 50 1115 65 1135
rect 85 1115 155 1135
rect 175 1115 190 1135
rect 50 1110 190 1115
rect 50 1090 100 1110
rect 140 1090 190 1110
rect 230 1135 370 1140
rect 230 1115 245 1135
rect 265 1115 335 1135
rect 355 1115 370 1135
rect 230 1110 370 1115
rect 230 1090 280 1110
rect 320 1090 370 1110
rect 410 1135 550 1140
rect 410 1115 425 1135
rect 445 1115 515 1135
rect 535 1115 550 1135
rect 410 1110 550 1115
rect 410 1090 460 1110
rect 500 1090 550 1110
rect 590 1135 730 1140
rect 590 1115 605 1135
rect 625 1115 695 1135
rect 715 1115 730 1135
rect 590 1110 730 1115
rect 590 1090 640 1110
rect 680 1090 730 1110
rect 770 1135 910 1140
rect 770 1115 785 1135
rect 805 1115 875 1135
rect 895 1115 910 1135
rect 770 1110 910 1115
rect 770 1090 820 1110
rect 860 1090 910 1110
rect 950 1135 1090 1140
rect 950 1115 965 1135
rect 985 1115 1055 1135
rect 1075 1115 1090 1135
rect 950 1110 1090 1115
rect 950 1090 1000 1110
rect 1040 1090 1090 1110
rect 1130 1135 1270 1140
rect 1130 1115 1145 1135
rect 1165 1115 1235 1135
rect 1255 1115 1270 1135
rect 1130 1110 1270 1115
rect 1130 1090 1180 1110
rect 1220 1090 1270 1110
rect 1310 1135 1450 1140
rect 1310 1115 1325 1135
rect 1345 1115 1415 1135
rect 1435 1115 1450 1135
rect 1310 1110 1450 1115
rect 1310 1090 1360 1110
rect 1400 1090 1450 1110
rect 1490 1135 1630 1140
rect 1490 1115 1505 1135
rect 1525 1115 1595 1135
rect 1615 1115 1630 1135
rect 1490 1110 1630 1115
rect 1490 1090 1540 1110
rect 1580 1090 1630 1110
rect 1670 1135 1810 1140
rect 1670 1115 1685 1135
rect 1705 1115 1775 1135
rect 1795 1115 1810 1135
rect 1670 1110 1810 1115
rect 1670 1090 1720 1110
rect 1760 1090 1810 1110
rect 1850 1135 1990 1140
rect 1850 1115 1865 1135
rect 1885 1115 1955 1135
rect 1975 1115 1990 1135
rect 1850 1110 1990 1115
rect 1850 1090 1900 1110
rect 1940 1090 1990 1110
rect 2030 1135 2170 1140
rect 2030 1115 2045 1135
rect 2065 1115 2135 1135
rect 2155 1115 2170 1135
rect 2030 1110 2170 1115
rect 2030 1090 2080 1110
rect 2120 1090 2170 1110
rect 2210 1135 2350 1140
rect 2210 1115 2225 1135
rect 2245 1115 2315 1135
rect 2335 1115 2350 1135
rect 2210 1110 2350 1115
rect 2210 1090 2260 1110
rect 2300 1090 2350 1110
rect 2390 1135 2530 1140
rect 2390 1115 2405 1135
rect 2425 1115 2495 1135
rect 2515 1115 2530 1135
rect 2390 1110 2530 1115
rect 2390 1090 2440 1110
rect 2480 1090 2530 1110
rect 2570 1135 2710 1140
rect 2570 1115 2585 1135
rect 2605 1115 2675 1135
rect 2695 1115 2710 1135
rect 2570 1110 2710 1115
rect 2570 1090 2620 1110
rect 2660 1090 2710 1110
rect 2750 1135 2890 1140
rect 2750 1115 2765 1135
rect 2785 1115 2855 1135
rect 2875 1115 2890 1135
rect 2750 1110 2890 1115
rect 2750 1090 2800 1110
rect 2840 1090 2890 1110
rect 2930 1135 3070 1140
rect 2930 1115 2945 1135
rect 2965 1115 3035 1135
rect 3055 1115 3070 1135
rect 2930 1110 3070 1115
rect 2930 1090 2980 1110
rect 3020 1090 3070 1110
rect 3115 1135 3255 1140
rect 3115 1115 3130 1135
rect 3150 1115 3220 1135
rect 3240 1115 3255 1135
rect 3115 1110 3255 1115
rect 3115 1090 3165 1110
rect 3205 1090 3255 1110
rect 3295 1135 3435 1140
rect 3295 1115 3310 1135
rect 3330 1115 3400 1135
rect 3420 1115 3435 1135
rect 3295 1110 3435 1115
rect 3295 1090 3345 1110
rect 3385 1090 3435 1110
rect 3475 1135 3615 1140
rect 3475 1115 3490 1135
rect 3510 1115 3580 1135
rect 3600 1115 3615 1135
rect 3475 1110 3615 1115
rect 3475 1090 3525 1110
rect 3565 1090 3615 1110
rect 3655 1135 3795 1140
rect 3655 1115 3670 1135
rect 3690 1115 3760 1135
rect 3780 1115 3795 1135
rect 3655 1110 3795 1115
rect 3655 1090 3705 1110
rect 3745 1090 3795 1110
rect 3835 1135 3975 1140
rect 3835 1115 3850 1135
rect 3870 1115 3940 1135
rect 3960 1115 3975 1135
rect 3835 1110 3975 1115
rect 3835 1090 3885 1110
rect 3925 1090 3975 1110
rect 4015 1135 4155 1140
rect 4015 1115 4030 1135
rect 4050 1115 4120 1135
rect 4140 1115 4155 1135
rect 4015 1110 4155 1115
rect 4015 1090 4065 1110
rect 4105 1090 4155 1110
rect 4195 1135 4335 1140
rect 4195 1115 4210 1135
rect 4230 1115 4300 1135
rect 4320 1115 4335 1135
rect 4195 1110 4335 1115
rect 4195 1090 4245 1110
rect 4285 1090 4335 1110
rect 4375 1135 4515 1140
rect 4375 1115 4390 1135
rect 4410 1115 4480 1135
rect 4500 1115 4515 1135
rect 4375 1110 4515 1115
rect 4375 1090 4425 1110
rect 4465 1090 4515 1110
rect 4555 1135 4695 1140
rect 4555 1115 4570 1135
rect 4590 1115 4660 1135
rect 4680 1115 4695 1135
rect 4555 1110 4695 1115
rect 4555 1090 4605 1110
rect 4645 1090 4695 1110
rect 4735 1135 4875 1140
rect 4735 1115 4750 1135
rect 4770 1115 4840 1135
rect 4860 1115 4875 1135
rect 4735 1110 4875 1115
rect 4735 1090 4785 1110
rect 4825 1090 4875 1110
rect 4915 1135 5055 1140
rect 4915 1115 4930 1135
rect 4950 1115 5020 1135
rect 5040 1115 5055 1135
rect 4915 1110 5055 1115
rect 4915 1090 4965 1110
rect 5005 1090 5055 1110
rect 5095 1135 5235 1140
rect 5095 1115 5110 1135
rect 5130 1115 5200 1135
rect 5220 1115 5235 1135
rect 5095 1110 5235 1115
rect 5095 1090 5145 1110
rect 5185 1090 5235 1110
rect 5275 1135 5415 1140
rect 5275 1115 5290 1135
rect 5310 1115 5380 1135
rect 5400 1115 5415 1135
rect 5275 1110 5415 1115
rect 5275 1090 5325 1110
rect 5365 1090 5415 1110
rect 5455 1135 5595 1140
rect 5455 1115 5470 1135
rect 5490 1115 5560 1135
rect 5580 1115 5595 1135
rect 5455 1110 5595 1115
rect 5455 1090 5505 1110
rect 5545 1090 5595 1110
rect 5635 1135 5775 1140
rect 5635 1115 5650 1135
rect 5670 1115 5740 1135
rect 5760 1115 5775 1135
rect 5635 1110 5775 1115
rect 5635 1090 5685 1110
rect 5725 1090 5775 1110
rect 5815 1135 5955 1140
rect 5815 1115 5830 1135
rect 5850 1115 5920 1135
rect 5940 1115 5955 1135
rect 5815 1110 5955 1115
rect 5815 1090 5865 1110
rect 5905 1090 5955 1110
rect 5995 1135 6135 1140
rect 5995 1115 6010 1135
rect 6030 1115 6100 1135
rect 6120 1115 6135 1135
rect 5995 1110 6135 1115
rect 5995 1090 6045 1110
rect 6085 1090 6135 1110
rect 6175 1135 6315 1140
rect 6175 1115 6190 1135
rect 6210 1115 6280 1135
rect 6300 1115 6315 1135
rect 6175 1110 6315 1115
rect 6175 1090 6225 1110
rect 6265 1090 6315 1110
rect 6355 1135 6495 1140
rect 6355 1115 6370 1135
rect 6390 1115 6460 1135
rect 6480 1115 6495 1135
rect 6355 1110 6495 1115
rect 6355 1090 6405 1110
rect 6445 1090 6495 1110
rect 6535 1135 6675 1140
rect 6535 1115 6550 1135
rect 6570 1115 6640 1135
rect 6660 1115 6675 1135
rect 6535 1110 6675 1115
rect 6535 1090 6585 1110
rect 6625 1090 6675 1110
rect 6715 1135 6855 1140
rect 6715 1115 6730 1135
rect 6750 1115 6820 1135
rect 6840 1115 6855 1135
rect 6715 1110 6855 1115
rect 6715 1090 6765 1110
rect 6805 1090 6855 1110
rect 6895 1135 7035 1140
rect 6895 1115 6910 1135
rect 6930 1115 7000 1135
rect 7020 1115 7035 1135
rect 6895 1110 7035 1115
rect 6895 1090 6945 1110
rect 6985 1090 7035 1110
rect 7075 1135 7215 1140
rect 7075 1115 7090 1135
rect 7110 1115 7180 1135
rect 7200 1115 7215 1135
rect 7075 1110 7215 1115
rect 7075 1090 7125 1110
rect 7165 1090 7215 1110
rect 7255 1135 7395 1140
rect 7255 1115 7270 1135
rect 7290 1115 7360 1135
rect 7380 1115 7395 1135
rect 7255 1110 7395 1115
rect 7255 1090 7305 1110
rect 7345 1090 7395 1110
rect 7435 1135 7575 1140
rect 7435 1115 7450 1135
rect 7470 1115 7540 1135
rect 7560 1115 7575 1135
rect 7435 1110 7575 1115
rect 7435 1090 7485 1110
rect 7525 1090 7575 1110
rect 7615 1135 7755 1140
rect 7615 1115 7630 1135
rect 7650 1115 7720 1135
rect 7740 1115 7755 1135
rect 7615 1110 7755 1115
rect 7615 1090 7665 1110
rect 7705 1090 7755 1110
rect 7795 1135 7935 1140
rect 7795 1115 7810 1135
rect 7830 1115 7900 1135
rect 7920 1115 7935 1135
rect 7795 1110 7935 1115
rect 7795 1090 7845 1110
rect 7885 1090 7935 1110
rect 7975 1135 8115 1140
rect 7975 1115 7990 1135
rect 8010 1115 8080 1135
rect 8100 1115 8115 1135
rect 7975 1110 8115 1115
rect 7975 1090 8025 1110
rect 8065 1090 8115 1110
rect 8155 1135 8295 1140
rect 8155 1115 8170 1135
rect 8190 1115 8260 1135
rect 8280 1115 8295 1135
rect 8155 1110 8295 1115
rect 8155 1090 8205 1110
rect 8245 1090 8295 1110
rect 8335 1135 8475 1140
rect 8335 1115 8350 1135
rect 8370 1115 8440 1135
rect 8460 1115 8475 1135
rect 8335 1110 8475 1115
rect 8335 1090 8385 1110
rect 8425 1090 8475 1110
rect 8515 1135 8655 1140
rect 8515 1115 8530 1135
rect 8550 1115 8620 1135
rect 8640 1115 8655 1135
rect 8515 1110 8655 1115
rect 8515 1090 8565 1110
rect 8605 1090 8655 1110
rect 8695 1135 8835 1140
rect 8695 1115 8710 1135
rect 8730 1115 8800 1135
rect 8820 1115 8835 1135
rect 8695 1110 8835 1115
rect 8695 1090 8745 1110
rect 8785 1090 8835 1110
rect 8875 1135 9015 1140
rect 8875 1115 8890 1135
rect 8910 1115 8980 1135
rect 9000 1115 9015 1135
rect 8875 1110 9015 1115
rect 8875 1090 8925 1110
rect 8965 1090 9015 1110
rect 9055 1135 9195 1140
rect 9055 1115 9070 1135
rect 9090 1115 9160 1135
rect 9180 1115 9195 1135
rect 9055 1110 9195 1115
rect 9055 1090 9105 1110
rect 9145 1090 9195 1110
rect 9235 1135 9375 1140
rect 9235 1115 9250 1135
rect 9270 1115 9340 1135
rect 9360 1115 9375 1135
rect 9235 1110 9375 1115
rect 9235 1090 9285 1110
rect 9325 1090 9375 1110
rect 9415 1135 9555 1140
rect 9415 1115 9430 1135
rect 9450 1115 9520 1135
rect 9540 1115 9555 1135
rect 9415 1110 9555 1115
rect 9415 1090 9465 1110
rect 9505 1090 9555 1110
rect 9595 1135 9735 1140
rect 9595 1115 9610 1135
rect 9630 1115 9700 1135
rect 9720 1115 9735 1135
rect 9595 1110 9735 1115
rect 9595 1090 9645 1110
rect 9685 1090 9735 1110
rect 9775 1135 9915 1140
rect 9775 1115 9790 1135
rect 9810 1115 9880 1135
rect 9900 1115 9915 1135
rect 9775 1110 9915 1115
rect 9775 1090 9825 1110
rect 9865 1090 9915 1110
rect 9955 1135 10095 1140
rect 9955 1115 9970 1135
rect 9990 1115 10060 1135
rect 10080 1115 10095 1135
rect 9955 1110 10095 1115
rect 9955 1090 10005 1110
rect 10045 1090 10095 1110
rect 10135 1135 10275 1140
rect 10135 1115 10150 1135
rect 10170 1115 10240 1135
rect 10260 1115 10275 1135
rect 10135 1110 10275 1115
rect 10135 1090 10185 1110
rect 10225 1090 10275 1110
rect 10315 1135 10455 1140
rect 10315 1115 10330 1135
rect 10350 1115 10420 1135
rect 10440 1115 10455 1135
rect 10315 1110 10455 1115
rect 10315 1090 10365 1110
rect 10405 1090 10455 1110
rect 10495 1135 10635 1140
rect 10495 1115 10510 1135
rect 10530 1115 10600 1135
rect 10620 1115 10635 1135
rect 10495 1110 10635 1115
rect 10495 1090 10545 1110
rect 10585 1090 10635 1110
rect 10675 1135 10815 1140
rect 10675 1115 10690 1135
rect 10710 1115 10780 1135
rect 10800 1115 10815 1135
rect 10675 1110 10815 1115
rect 10675 1090 10725 1110
rect 10765 1090 10815 1110
rect 10855 1135 10995 1140
rect 10855 1115 10870 1135
rect 10890 1115 10960 1135
rect 10980 1115 10995 1135
rect 10855 1110 10995 1115
rect 10855 1090 10905 1110
rect 10945 1090 10995 1110
rect 11035 1135 11175 1140
rect 11035 1115 11050 1135
rect 11070 1115 11140 1135
rect 11160 1115 11175 1135
rect 11035 1110 11175 1115
rect 11035 1090 11085 1110
rect 11125 1090 11175 1110
rect -310 975 -260 990
rect -220 975 -170 990
rect -130 975 -80 990
rect -40 975 10 990
rect 50 975 100 990
rect 140 975 190 990
rect 230 975 280 990
rect 320 975 370 990
rect 410 975 460 990
rect 500 975 550 990
rect 590 975 640 990
rect 680 975 730 990
rect 770 975 820 990
rect 860 975 910 990
rect 950 975 1000 990
rect 1040 975 1090 990
rect 1130 975 1180 990
rect 1220 975 1270 990
rect 1310 975 1360 990
rect 1400 975 1450 990
rect 1490 975 1540 990
rect 1580 975 1630 990
rect 1670 975 1720 990
rect 1760 975 1810 990
rect 1850 975 1900 990
rect 1940 975 1990 990
rect 2030 975 2080 990
rect 2120 975 2170 990
rect 2210 975 2260 990
rect 2300 975 2350 990
rect 2390 975 2440 990
rect 2480 975 2530 990
rect 2570 975 2620 990
rect 2660 975 2710 990
rect 2750 975 2800 990
rect 2840 975 2890 990
rect 2930 975 2980 990
rect 3020 975 3070 990
rect 3115 975 3165 990
rect 3205 975 3255 990
rect 3295 975 3345 990
rect 3385 975 3435 990
rect 3475 975 3525 990
rect 3565 975 3615 990
rect 3655 975 3705 990
rect 3745 975 3795 990
rect 3835 975 3885 990
rect 3925 975 3975 990
rect 4015 975 4065 990
rect 4105 975 4155 990
rect 4195 975 4245 990
rect 4285 975 4335 990
rect 4375 975 4425 990
rect 4465 975 4515 990
rect 4555 975 4605 990
rect 4645 975 4695 990
rect 4735 975 4785 990
rect 4825 975 4875 990
rect 4915 975 4965 990
rect 5005 975 5055 990
rect 5095 975 5145 990
rect 5185 975 5235 990
rect 5275 975 5325 990
rect 5365 975 5415 990
rect 5455 975 5505 990
rect 5545 975 5595 990
rect 5635 975 5685 990
rect 5725 975 5775 990
rect 5815 975 5865 990
rect 5905 975 5955 990
rect 5995 975 6045 990
rect 6085 975 6135 990
rect 6175 975 6225 990
rect 6265 975 6315 990
rect 6355 975 6405 990
rect 6445 975 6495 990
rect 6535 975 6585 990
rect 6625 975 6675 990
rect 6715 975 6765 990
rect 6805 975 6855 990
rect 6895 975 6945 990
rect 6985 975 7035 990
rect 7075 975 7125 990
rect 7165 975 7215 990
rect 7255 975 7305 990
rect 7345 975 7395 990
rect 7435 975 7485 990
rect 7525 975 7575 990
rect 7615 975 7665 990
rect 7705 975 7755 990
rect 7795 975 7845 990
rect 7885 975 7935 990
rect 7975 975 8025 990
rect 8065 975 8115 990
rect 8155 975 8205 990
rect 8245 975 8295 990
rect 8335 975 8385 990
rect 8425 975 8475 990
rect 8515 975 8565 990
rect 8605 975 8655 990
rect 8695 975 8745 990
rect 8785 975 8835 990
rect 8875 975 8925 990
rect 8965 975 9015 990
rect 9055 975 9105 990
rect 9145 975 9195 990
rect 9235 975 9285 990
rect 9325 975 9375 990
rect 9415 975 9465 990
rect 9505 975 9555 990
rect 9595 975 9645 990
rect 9685 975 9735 990
rect 9775 975 9825 990
rect 9865 975 9915 990
rect 9955 975 10005 990
rect 10045 975 10095 990
rect 10135 975 10185 990
rect 10225 975 10275 990
rect 10315 975 10365 990
rect 10405 975 10455 990
rect 10495 975 10545 990
rect 10585 975 10635 990
rect 10675 975 10725 990
rect 10765 975 10815 990
rect 10855 975 10905 990
rect 10945 975 10995 990
rect 11035 975 11085 990
rect 11125 975 11175 990
rect -310 850 -260 865
rect -220 850 -170 865
rect -130 850 -80 865
rect -40 850 10 865
rect 50 850 100 865
rect 140 850 190 865
rect 230 850 280 865
rect 320 850 370 865
rect 410 850 460 865
rect 500 850 550 865
rect 590 850 640 865
rect 680 850 730 865
rect 770 850 820 865
rect 860 850 910 865
rect 950 850 1000 865
rect 1040 850 1090 865
rect 1130 850 1180 865
rect 1220 850 1270 865
rect 1310 850 1360 865
rect 1400 850 1450 865
rect 1490 850 1540 865
rect 1580 850 1630 865
rect 1670 850 1720 865
rect 1760 850 1810 865
rect 1850 850 1900 865
rect 1940 850 1990 865
rect 2030 850 2080 865
rect 2120 850 2170 865
rect 2210 850 2260 865
rect 2300 850 2350 865
rect 2390 850 2440 865
rect 2480 850 2530 865
rect 2570 850 2620 865
rect 2660 850 2710 865
rect 2750 850 2800 865
rect 2840 850 2890 865
rect 2930 850 2980 865
rect 3020 850 3070 865
rect 3110 850 3160 865
rect 3200 850 3250 865
rect 3290 850 3340 865
rect 3380 850 3430 865
rect 3470 850 3520 865
rect 3560 850 3610 865
rect 3650 850 3700 865
rect 3740 850 3790 865
rect 3830 850 3880 865
rect 3920 850 3970 865
rect 4010 850 4060 865
rect 4100 850 4150 865
rect 4190 850 4240 865
rect 4280 850 4330 865
rect 4370 850 4420 865
rect 4460 850 4510 865
rect 4550 850 4600 865
rect 4640 850 4690 865
rect 4730 850 4780 865
rect 4820 850 4870 865
rect 4910 850 4960 865
rect 5000 850 5050 865
rect 5090 850 5140 865
rect 5180 850 5230 865
rect 5270 850 5320 865
rect 5360 850 5410 865
rect 5450 850 5500 865
rect 5540 850 5590 865
rect 5630 850 5680 865
rect 5720 850 5770 865
rect 5810 850 5860 865
rect 5900 850 5950 865
rect 5990 850 6040 865
rect 6080 850 6130 865
rect 6170 850 6220 865
rect 6260 850 6310 865
rect 6350 850 6400 865
rect 6440 850 6490 865
rect 6530 850 6580 865
rect 6620 850 6670 865
rect 6710 850 6760 865
rect 6800 850 6850 865
rect 6890 850 6940 865
rect 6980 850 7030 865
rect 7070 850 7120 865
rect 7160 850 7210 865
rect 7250 850 7300 865
rect 7340 850 7390 865
rect 7430 850 7480 865
rect 7520 850 7570 865
rect 7610 850 7660 865
rect 7700 850 7750 865
rect 7795 850 7845 865
rect 7885 850 7935 865
rect 7975 850 8025 865
rect 8065 850 8115 865
rect 8155 850 8205 865
rect 8245 850 8295 865
rect 8335 850 8385 865
rect 8425 850 8475 865
rect 8515 850 8565 865
rect 8605 850 8655 865
rect 8695 850 8745 865
rect 8785 850 8835 865
rect 8875 850 8925 865
rect 8965 850 9015 865
rect 9055 850 9105 865
rect 9145 850 9195 865
rect 9235 850 9285 865
rect 9325 850 9375 865
rect 9415 850 9465 865
rect 9505 850 9555 865
rect 9595 850 9645 865
rect 9685 850 9735 865
rect 9775 850 9825 865
rect 9865 850 9915 865
rect 9955 850 10005 865
rect 10045 850 10095 865
rect 10135 850 10185 865
rect 10225 850 10275 865
rect 10315 850 10365 865
rect 10405 850 10455 865
rect 10495 850 10545 865
rect 10585 850 10635 865
rect 10675 850 10725 865
rect 10765 850 10815 865
rect 10855 850 10905 865
rect 10945 850 10995 865
rect 11035 850 11085 865
rect 11125 850 11175 865
rect -310 730 -260 750
rect -220 730 -170 750
rect -310 725 -170 730
rect -310 705 -295 725
rect -275 705 -205 725
rect -185 705 -170 725
rect -310 700 -170 705
rect -130 730 -80 750
rect -40 730 10 750
rect -130 725 10 730
rect -130 705 -115 725
rect -95 705 -25 725
rect -5 705 10 725
rect -130 700 10 705
rect 50 730 100 750
rect 140 730 190 750
rect 50 725 190 730
rect 50 705 65 725
rect 85 705 155 725
rect 175 705 190 725
rect 50 700 190 705
rect 230 730 280 750
rect 320 730 370 750
rect 230 725 370 730
rect 230 705 245 725
rect 265 705 335 725
rect 355 705 370 725
rect 230 700 370 705
rect 410 730 460 750
rect 500 730 550 750
rect 410 725 550 730
rect 410 705 425 725
rect 445 705 515 725
rect 535 705 550 725
rect 410 700 550 705
rect 590 730 640 750
rect 680 730 730 750
rect 590 725 730 730
rect 590 705 605 725
rect 625 705 695 725
rect 715 705 730 725
rect 590 700 730 705
rect 770 730 820 750
rect 860 730 910 750
rect 770 725 910 730
rect 770 705 785 725
rect 805 705 875 725
rect 895 705 910 725
rect 770 700 910 705
rect 950 730 1000 750
rect 1040 730 1090 750
rect 950 725 1090 730
rect 950 705 965 725
rect 985 705 1055 725
rect 1075 705 1090 725
rect 950 700 1090 705
rect 1130 730 1180 750
rect 1220 730 1270 750
rect 1130 725 1270 730
rect 1130 705 1145 725
rect 1165 705 1235 725
rect 1255 705 1270 725
rect 1130 700 1270 705
rect 1310 730 1360 750
rect 1400 730 1450 750
rect 1310 725 1450 730
rect 1310 705 1325 725
rect 1345 705 1415 725
rect 1435 705 1450 725
rect 1310 700 1450 705
rect 1490 730 1540 750
rect 1580 730 1630 750
rect 1490 725 1630 730
rect 1490 705 1505 725
rect 1525 705 1595 725
rect 1615 705 1630 725
rect 1490 700 1630 705
rect 1670 730 1720 750
rect 1760 730 1810 750
rect 1670 725 1810 730
rect 1670 705 1685 725
rect 1705 705 1775 725
rect 1795 705 1810 725
rect 1670 700 1810 705
rect 1850 730 1900 750
rect 1940 730 1990 750
rect 1850 725 1990 730
rect 1850 705 1865 725
rect 1885 705 1955 725
rect 1975 705 1990 725
rect 1850 700 1990 705
rect 2030 730 2080 750
rect 2120 730 2170 750
rect 2030 725 2170 730
rect 2030 705 2045 725
rect 2065 705 2135 725
rect 2155 705 2170 725
rect 2030 700 2170 705
rect 2210 730 2260 750
rect 2300 730 2350 750
rect 2210 725 2350 730
rect 2210 705 2225 725
rect 2245 705 2315 725
rect 2335 705 2350 725
rect 2210 700 2350 705
rect 2390 730 2440 750
rect 2480 730 2530 750
rect 2390 725 2530 730
rect 2390 705 2405 725
rect 2425 705 2495 725
rect 2515 705 2530 725
rect 2390 700 2530 705
rect 2570 730 2620 750
rect 2660 730 2710 750
rect 2570 725 2710 730
rect 2570 705 2585 725
rect 2605 705 2675 725
rect 2695 705 2710 725
rect 2570 700 2710 705
rect 2750 730 2800 750
rect 2840 730 2890 750
rect 2750 725 2890 730
rect 2750 705 2765 725
rect 2785 705 2855 725
rect 2875 705 2890 725
rect 2750 700 2890 705
rect 2930 730 2980 750
rect 3020 730 3070 750
rect 2930 725 3070 730
rect 2930 705 2945 725
rect 2965 705 3035 725
rect 3055 705 3070 725
rect 2930 700 3070 705
rect 3110 730 3160 750
rect 3200 730 3250 750
rect 3110 725 3250 730
rect 3110 705 3125 725
rect 3145 705 3215 725
rect 3235 705 3250 725
rect 3110 700 3250 705
rect 3290 730 3340 750
rect 3380 730 3430 750
rect 3290 725 3430 730
rect 3290 705 3305 725
rect 3325 705 3395 725
rect 3415 705 3430 725
rect 3290 700 3430 705
rect 3470 730 3520 750
rect 3560 730 3610 750
rect 3470 725 3610 730
rect 3470 705 3485 725
rect 3505 705 3575 725
rect 3595 705 3610 725
rect 3470 700 3610 705
rect 3650 730 3700 750
rect 3740 730 3790 750
rect 3650 725 3790 730
rect 3650 705 3665 725
rect 3685 705 3755 725
rect 3775 705 3790 725
rect 3650 700 3790 705
rect 3830 730 3880 750
rect 3920 730 3970 750
rect 3830 725 3970 730
rect 3830 705 3845 725
rect 3865 705 3935 725
rect 3955 705 3970 725
rect 3830 700 3970 705
rect 4010 730 4060 750
rect 4100 730 4150 750
rect 4010 725 4150 730
rect 4010 705 4025 725
rect 4045 705 4115 725
rect 4135 705 4150 725
rect 4010 700 4150 705
rect 4190 730 4240 750
rect 4280 730 4330 750
rect 4190 725 4330 730
rect 4190 705 4205 725
rect 4225 705 4295 725
rect 4315 705 4330 725
rect 4190 700 4330 705
rect 4370 730 4420 750
rect 4460 730 4510 750
rect 4370 725 4510 730
rect 4370 705 4385 725
rect 4405 705 4475 725
rect 4495 705 4510 725
rect 4370 700 4510 705
rect 4550 730 4600 750
rect 4640 730 4690 750
rect 4550 725 4690 730
rect 4550 705 4565 725
rect 4585 705 4655 725
rect 4675 705 4690 725
rect 4550 700 4690 705
rect 4730 730 4780 750
rect 4820 730 4870 750
rect 4730 725 4870 730
rect 4730 705 4745 725
rect 4765 705 4835 725
rect 4855 705 4870 725
rect 4730 700 4870 705
rect 4910 730 4960 750
rect 5000 730 5050 750
rect 4910 725 5050 730
rect 4910 705 4925 725
rect 4945 705 5015 725
rect 5035 705 5050 725
rect 4910 700 5050 705
rect 5090 730 5140 750
rect 5180 730 5230 750
rect 5090 725 5230 730
rect 5090 705 5105 725
rect 5125 705 5195 725
rect 5215 705 5230 725
rect 5090 700 5230 705
rect 5270 730 5320 750
rect 5360 730 5410 750
rect 5270 725 5410 730
rect 5270 705 5285 725
rect 5305 705 5375 725
rect 5395 705 5410 725
rect 5270 700 5410 705
rect 5450 730 5500 750
rect 5540 730 5590 750
rect 5450 725 5590 730
rect 5450 705 5465 725
rect 5485 705 5555 725
rect 5575 705 5590 725
rect 5450 700 5590 705
rect 5630 730 5680 750
rect 5720 730 5770 750
rect 5630 725 5770 730
rect 5630 705 5645 725
rect 5665 705 5735 725
rect 5755 705 5770 725
rect 5630 700 5770 705
rect 5810 730 5860 750
rect 5900 730 5950 750
rect 5810 725 5950 730
rect 5810 705 5825 725
rect 5845 705 5915 725
rect 5935 705 5950 725
rect 5810 700 5950 705
rect 5990 730 6040 750
rect 6080 730 6130 750
rect 5990 725 6130 730
rect 5990 705 6005 725
rect 6025 705 6095 725
rect 6115 705 6130 725
rect 5990 700 6130 705
rect 6170 730 6220 750
rect 6260 730 6310 750
rect 6170 725 6310 730
rect 6170 705 6185 725
rect 6205 705 6275 725
rect 6295 705 6310 725
rect 6170 700 6310 705
rect 6350 730 6400 750
rect 6440 730 6490 750
rect 6350 725 6490 730
rect 6350 705 6365 725
rect 6385 705 6455 725
rect 6475 705 6490 725
rect 6350 700 6490 705
rect 6530 730 6580 750
rect 6620 730 6670 750
rect 6530 725 6670 730
rect 6530 705 6545 725
rect 6565 705 6635 725
rect 6655 705 6670 725
rect 6530 700 6670 705
rect 6710 730 6760 750
rect 6800 730 6850 750
rect 6710 725 6850 730
rect 6710 705 6725 725
rect 6745 705 6815 725
rect 6835 705 6850 725
rect 6710 700 6850 705
rect 6890 730 6940 750
rect 6980 730 7030 750
rect 6890 725 7030 730
rect 6890 705 6905 725
rect 6925 705 6995 725
rect 7015 705 7030 725
rect 6890 700 7030 705
rect 7070 730 7120 750
rect 7160 730 7210 750
rect 7070 725 7210 730
rect 7070 705 7085 725
rect 7105 705 7175 725
rect 7195 705 7210 725
rect 7070 700 7210 705
rect 7250 730 7300 750
rect 7340 730 7390 750
rect 7250 725 7390 730
rect 7250 705 7265 725
rect 7285 705 7355 725
rect 7375 705 7390 725
rect 7250 700 7390 705
rect 7430 730 7480 750
rect 7520 730 7570 750
rect 7430 725 7570 730
rect 7430 705 7445 725
rect 7465 705 7535 725
rect 7555 705 7570 725
rect 7430 700 7570 705
rect 7610 730 7660 750
rect 7700 730 7750 750
rect 7610 725 7750 730
rect 7610 705 7625 725
rect 7645 705 7715 725
rect 7735 705 7750 725
rect 7610 700 7750 705
rect 7795 730 7845 750
rect 7885 730 7935 750
rect 7795 725 7935 730
rect 7795 705 7810 725
rect 7830 705 7900 725
rect 7920 705 7935 725
rect 7795 700 7935 705
rect 7975 730 8025 750
rect 8065 730 8115 750
rect 7975 725 8115 730
rect 7975 705 7990 725
rect 8010 705 8080 725
rect 8100 705 8115 725
rect 7975 700 8115 705
rect 8155 730 8205 750
rect 8245 730 8295 750
rect 8155 725 8295 730
rect 8155 705 8170 725
rect 8190 705 8260 725
rect 8280 705 8295 725
rect 8155 700 8295 705
rect 8335 730 8385 750
rect 8425 730 8475 750
rect 8335 725 8475 730
rect 8335 705 8350 725
rect 8370 705 8440 725
rect 8460 705 8475 725
rect 8335 700 8475 705
rect 8515 730 8565 750
rect 8605 730 8655 750
rect 8515 725 8655 730
rect 8515 705 8530 725
rect 8550 705 8620 725
rect 8640 705 8655 725
rect 8515 700 8655 705
rect 8695 730 8745 750
rect 8785 730 8835 750
rect 8695 725 8835 730
rect 8695 705 8710 725
rect 8730 705 8800 725
rect 8820 705 8835 725
rect 8695 700 8835 705
rect 8875 730 8925 750
rect 8965 730 9015 750
rect 8875 725 9015 730
rect 8875 705 8890 725
rect 8910 705 8980 725
rect 9000 705 9015 725
rect 8875 700 9015 705
rect 9055 730 9105 750
rect 9145 730 9195 750
rect 9055 725 9195 730
rect 9055 705 9070 725
rect 9090 705 9160 725
rect 9180 705 9195 725
rect 9055 700 9195 705
rect 9235 730 9285 750
rect 9325 730 9375 750
rect 9235 725 9375 730
rect 9235 705 9250 725
rect 9270 705 9340 725
rect 9360 705 9375 725
rect 9235 700 9375 705
rect 9415 730 9465 750
rect 9505 730 9555 750
rect 9415 725 9555 730
rect 9415 705 9430 725
rect 9450 705 9520 725
rect 9540 705 9555 725
rect 9415 700 9555 705
rect 9595 730 9645 750
rect 9685 730 9735 750
rect 9595 725 9735 730
rect 9595 705 9610 725
rect 9630 705 9700 725
rect 9720 705 9735 725
rect 9595 700 9735 705
rect 9775 730 9825 750
rect 9865 730 9915 750
rect 9775 725 9915 730
rect 9775 705 9790 725
rect 9810 705 9880 725
rect 9900 705 9915 725
rect 9775 700 9915 705
rect 9955 730 10005 750
rect 10045 730 10095 750
rect 9955 725 10095 730
rect 9955 705 9970 725
rect 9990 705 10060 725
rect 10080 705 10095 725
rect 9955 700 10095 705
rect 10135 730 10185 750
rect 10225 730 10275 750
rect 10135 725 10275 730
rect 10135 705 10150 725
rect 10170 705 10240 725
rect 10260 705 10275 725
rect 10135 700 10275 705
rect 10315 730 10365 750
rect 10405 730 10455 750
rect 10315 725 10455 730
rect 10315 705 10330 725
rect 10350 705 10420 725
rect 10440 705 10455 725
rect 10315 700 10455 705
rect 10495 730 10545 750
rect 10585 730 10635 750
rect 10495 725 10635 730
rect 10495 705 10510 725
rect 10530 705 10600 725
rect 10620 705 10635 725
rect 10495 700 10635 705
rect 10675 730 10725 750
rect 10765 730 10815 750
rect 10675 725 10815 730
rect 10675 705 10690 725
rect 10710 705 10780 725
rect 10800 705 10815 725
rect 10675 700 10815 705
rect 10855 730 10905 750
rect 10945 730 10995 750
rect 10855 725 10995 730
rect 10855 705 10870 725
rect 10890 705 10960 725
rect 10980 705 10995 725
rect 10855 700 10995 705
rect 11035 730 11085 750
rect 11125 730 11175 750
rect 11035 725 11175 730
rect 11035 705 11050 725
rect 11070 705 11140 725
rect 11160 705 11175 725
rect 11035 700 11175 705
rect -310 195 -170 200
rect -310 175 -295 195
rect -275 175 -205 195
rect -185 175 -170 195
rect -310 170 -170 175
rect -310 150 -260 170
rect -220 150 -170 170
rect -130 195 10 200
rect -130 175 -115 195
rect -95 175 -25 195
rect -5 175 10 195
rect -130 170 10 175
rect -130 150 -80 170
rect -40 150 10 170
rect 50 195 190 200
rect 50 175 65 195
rect 85 175 155 195
rect 175 175 190 195
rect 50 170 190 175
rect 50 150 100 170
rect 140 150 190 170
rect 230 195 370 200
rect 230 175 245 195
rect 265 175 335 195
rect 355 175 370 195
rect 230 170 370 175
rect 230 150 280 170
rect 320 150 370 170
rect 410 195 550 200
rect 410 175 425 195
rect 445 175 515 195
rect 535 175 550 195
rect 410 170 550 175
rect 410 150 460 170
rect 500 150 550 170
rect 590 195 730 200
rect 590 175 605 195
rect 625 175 695 195
rect 715 175 730 195
rect 590 170 730 175
rect 590 150 640 170
rect 680 150 730 170
rect 770 195 910 200
rect 770 175 785 195
rect 805 175 875 195
rect 895 175 910 195
rect 770 170 910 175
rect 770 150 820 170
rect 860 150 910 170
rect 950 195 1090 200
rect 950 175 965 195
rect 985 175 1055 195
rect 1075 175 1090 195
rect 950 170 1090 175
rect 950 150 1000 170
rect 1040 150 1090 170
rect 1130 195 1270 200
rect 1130 175 1145 195
rect 1165 175 1235 195
rect 1255 175 1270 195
rect 1130 170 1270 175
rect 1130 150 1180 170
rect 1220 150 1270 170
rect 1310 195 1450 200
rect 1310 175 1325 195
rect 1345 175 1415 195
rect 1435 175 1450 195
rect 1310 170 1450 175
rect 1310 150 1360 170
rect 1400 150 1450 170
rect 1490 195 1630 200
rect 1490 175 1505 195
rect 1525 175 1595 195
rect 1615 175 1630 195
rect 1490 170 1630 175
rect 1490 150 1540 170
rect 1580 150 1630 170
rect 1670 195 1810 200
rect 1670 175 1685 195
rect 1705 175 1775 195
rect 1795 175 1810 195
rect 1670 170 1810 175
rect 1670 150 1720 170
rect 1760 150 1810 170
rect 1850 195 1990 200
rect 1850 175 1865 195
rect 1885 175 1955 195
rect 1975 175 1990 195
rect 1850 170 1990 175
rect 1850 150 1900 170
rect 1940 150 1990 170
rect 2030 195 2170 200
rect 2030 175 2045 195
rect 2065 175 2135 195
rect 2155 175 2170 195
rect 2030 170 2170 175
rect 2030 150 2080 170
rect 2120 150 2170 170
rect 2210 195 2350 200
rect 2210 175 2225 195
rect 2245 175 2315 195
rect 2335 175 2350 195
rect 2210 170 2350 175
rect 2210 150 2260 170
rect 2300 150 2350 170
rect 2390 195 2530 200
rect 2390 175 2405 195
rect 2425 175 2495 195
rect 2515 175 2530 195
rect 2390 170 2530 175
rect 2390 150 2440 170
rect 2480 150 2530 170
rect 2570 195 2710 200
rect 2570 175 2585 195
rect 2605 175 2675 195
rect 2695 175 2710 195
rect 2570 170 2710 175
rect 2570 150 2620 170
rect 2660 150 2710 170
rect 2750 195 2890 200
rect 2750 175 2765 195
rect 2785 175 2855 195
rect 2875 175 2890 195
rect 2750 170 2890 175
rect 2750 150 2800 170
rect 2840 150 2890 170
rect 2930 195 3070 200
rect 2930 175 2945 195
rect 2965 175 3035 195
rect 3055 175 3070 195
rect 2930 170 3070 175
rect 2930 150 2980 170
rect 3020 150 3070 170
rect 3110 195 3250 200
rect 3110 175 3125 195
rect 3145 175 3215 195
rect 3235 175 3250 195
rect 3110 170 3250 175
rect 3110 150 3160 170
rect 3200 150 3250 170
rect 3290 195 3430 200
rect 3290 175 3305 195
rect 3325 175 3395 195
rect 3415 175 3430 195
rect 3290 170 3430 175
rect 3290 150 3340 170
rect 3380 150 3430 170
rect 3470 195 3610 200
rect 3470 175 3485 195
rect 3505 175 3575 195
rect 3595 175 3610 195
rect 3470 170 3610 175
rect 3470 150 3520 170
rect 3560 150 3610 170
rect 3650 195 3790 200
rect 3650 175 3665 195
rect 3685 175 3755 195
rect 3775 175 3790 195
rect 3650 170 3790 175
rect 3650 150 3700 170
rect 3740 150 3790 170
rect 3830 195 3970 200
rect 3830 175 3845 195
rect 3865 175 3935 195
rect 3955 175 3970 195
rect 3830 170 3970 175
rect 3830 150 3880 170
rect 3920 150 3970 170
rect 4010 195 4150 200
rect 4010 175 4025 195
rect 4045 175 4115 195
rect 4135 175 4150 195
rect 4010 170 4150 175
rect 4010 150 4060 170
rect 4100 150 4150 170
rect 4190 195 4330 200
rect 4190 175 4205 195
rect 4225 175 4295 195
rect 4315 175 4330 195
rect 4190 170 4330 175
rect 4190 150 4240 170
rect 4280 150 4330 170
rect 4370 195 4510 200
rect 4370 175 4385 195
rect 4405 175 4475 195
rect 4495 175 4510 195
rect 4370 170 4510 175
rect 4370 150 4420 170
rect 4460 150 4510 170
rect 4550 195 4690 200
rect 4550 175 4565 195
rect 4585 175 4655 195
rect 4675 175 4690 195
rect 4550 170 4690 175
rect 4550 150 4600 170
rect 4640 150 4690 170
rect 4730 195 4870 200
rect 4730 175 4745 195
rect 4765 175 4835 195
rect 4855 175 4870 195
rect 4730 170 4870 175
rect 4730 150 4780 170
rect 4820 150 4870 170
rect 4910 195 5050 200
rect 4910 175 4925 195
rect 4945 175 5015 195
rect 5035 175 5050 195
rect 4910 170 5050 175
rect 4910 150 4960 170
rect 5000 150 5050 170
rect 5090 195 5230 200
rect 5090 175 5105 195
rect 5125 175 5195 195
rect 5215 175 5230 195
rect 5090 170 5230 175
rect 5090 150 5140 170
rect 5180 150 5230 170
rect 5270 195 5410 200
rect 5270 175 5285 195
rect 5305 175 5375 195
rect 5395 175 5410 195
rect 5270 170 5410 175
rect 5270 150 5320 170
rect 5360 150 5410 170
rect 5450 195 5590 200
rect 5450 175 5465 195
rect 5485 175 5555 195
rect 5575 175 5590 195
rect 5450 170 5590 175
rect 5450 150 5500 170
rect 5540 150 5590 170
rect 5630 195 5770 200
rect 5630 175 5645 195
rect 5665 175 5735 195
rect 5755 175 5770 195
rect 5630 170 5770 175
rect 5630 150 5680 170
rect 5720 150 5770 170
rect 5810 195 5950 200
rect 5810 175 5825 195
rect 5845 175 5915 195
rect 5935 175 5950 195
rect 5810 170 5950 175
rect 5810 150 5860 170
rect 5900 150 5950 170
rect 5990 195 6130 200
rect 5990 175 6005 195
rect 6025 175 6095 195
rect 6115 175 6130 195
rect 5990 170 6130 175
rect 5990 150 6040 170
rect 6080 150 6130 170
rect 6170 195 6310 200
rect 6170 175 6185 195
rect 6205 175 6275 195
rect 6295 175 6310 195
rect 6170 170 6310 175
rect 6170 150 6220 170
rect 6260 150 6310 170
rect 6350 195 6490 200
rect 6350 175 6365 195
rect 6385 175 6455 195
rect 6475 175 6490 195
rect 6350 170 6490 175
rect 6350 150 6400 170
rect 6440 150 6490 170
rect 6530 195 6670 200
rect 6530 175 6545 195
rect 6565 175 6635 195
rect 6655 175 6670 195
rect 6530 170 6670 175
rect 6530 150 6580 170
rect 6620 150 6670 170
rect 6710 195 6850 200
rect 6710 175 6725 195
rect 6745 175 6815 195
rect 6835 175 6850 195
rect 6710 170 6850 175
rect 6710 150 6760 170
rect 6800 150 6850 170
rect 6890 195 7030 200
rect 6890 175 6905 195
rect 6925 175 6995 195
rect 7015 175 7030 195
rect 6890 170 7030 175
rect 6890 150 6940 170
rect 6980 150 7030 170
rect 7070 195 7210 200
rect 7070 175 7085 195
rect 7105 175 7175 195
rect 7195 175 7210 195
rect 7070 170 7210 175
rect 7070 150 7120 170
rect 7160 150 7210 170
rect 7250 195 7390 200
rect 7250 175 7265 195
rect 7285 175 7355 195
rect 7375 175 7390 195
rect 7250 170 7390 175
rect 7250 150 7300 170
rect 7340 150 7390 170
rect 7430 195 7570 200
rect 7430 175 7445 195
rect 7465 175 7535 195
rect 7555 175 7570 195
rect 7430 170 7570 175
rect 7430 150 7480 170
rect 7520 150 7570 170
rect 7610 195 7750 200
rect 7610 175 7625 195
rect 7645 175 7715 195
rect 7735 175 7750 195
rect 7610 170 7750 175
rect 7610 150 7660 170
rect 7700 150 7750 170
rect 7795 195 7935 200
rect 7795 175 7810 195
rect 7830 175 7900 195
rect 7920 175 7935 195
rect 7795 170 7935 175
rect 7795 150 7845 170
rect 7885 150 7935 170
rect 7975 195 8115 200
rect 7975 175 7990 195
rect 8010 175 8080 195
rect 8100 175 8115 195
rect 7975 170 8115 175
rect 7975 150 8025 170
rect 8065 150 8115 170
rect 8155 195 8295 200
rect 8155 175 8170 195
rect 8190 175 8260 195
rect 8280 175 8295 195
rect 8155 170 8295 175
rect 8155 150 8205 170
rect 8245 150 8295 170
rect 8335 195 8475 200
rect 8335 175 8350 195
rect 8370 175 8440 195
rect 8460 175 8475 195
rect 8335 170 8475 175
rect 8335 150 8385 170
rect 8425 150 8475 170
rect 8515 195 8655 200
rect 8515 175 8530 195
rect 8550 175 8620 195
rect 8640 175 8655 195
rect 8515 170 8655 175
rect 8515 150 8565 170
rect 8605 150 8655 170
rect 8695 195 8835 200
rect 8695 175 8710 195
rect 8730 175 8800 195
rect 8820 175 8835 195
rect 8695 170 8835 175
rect 8695 150 8745 170
rect 8785 150 8835 170
rect 8875 195 9015 200
rect 8875 175 8890 195
rect 8910 175 8980 195
rect 9000 175 9015 195
rect 8875 170 9015 175
rect 8875 150 8925 170
rect 8965 150 9015 170
rect 9055 195 9195 200
rect 9055 175 9070 195
rect 9090 175 9160 195
rect 9180 175 9195 195
rect 9055 170 9195 175
rect 9055 150 9105 170
rect 9145 150 9195 170
rect 9235 195 9375 200
rect 9235 175 9250 195
rect 9270 175 9340 195
rect 9360 175 9375 195
rect 9235 170 9375 175
rect 9235 150 9285 170
rect 9325 150 9375 170
rect 9415 195 9555 200
rect 9415 175 9430 195
rect 9450 175 9520 195
rect 9540 175 9555 195
rect 9415 170 9555 175
rect 9415 150 9465 170
rect 9505 150 9555 170
rect 9595 195 9735 200
rect 9595 175 9610 195
rect 9630 175 9700 195
rect 9720 175 9735 195
rect 9595 170 9735 175
rect 9595 150 9645 170
rect 9685 150 9735 170
rect 9775 195 9915 200
rect 9775 175 9790 195
rect 9810 175 9880 195
rect 9900 175 9915 195
rect 9775 170 9915 175
rect 9775 150 9825 170
rect 9865 150 9915 170
rect 9955 195 10095 200
rect 9955 175 9970 195
rect 9990 175 10060 195
rect 10080 175 10095 195
rect 9955 170 10095 175
rect 9955 150 10005 170
rect 10045 150 10095 170
rect 10135 195 10275 200
rect 10135 175 10150 195
rect 10170 175 10240 195
rect 10260 175 10275 195
rect 10135 170 10275 175
rect 10135 150 10185 170
rect 10225 150 10275 170
rect 10315 195 10455 200
rect 10315 175 10330 195
rect 10350 175 10420 195
rect 10440 175 10455 195
rect 10315 170 10455 175
rect 10315 150 10365 170
rect 10405 150 10455 170
rect 10495 195 10635 200
rect 10495 175 10510 195
rect 10530 175 10600 195
rect 10620 175 10635 195
rect 10495 170 10635 175
rect 10495 150 10545 170
rect 10585 150 10635 170
rect 10675 195 10815 200
rect 10675 175 10690 195
rect 10710 175 10780 195
rect 10800 175 10815 195
rect 10675 170 10815 175
rect 10675 150 10725 170
rect 10765 150 10815 170
rect 10855 195 10995 200
rect 10855 175 10870 195
rect 10890 175 10960 195
rect 10980 175 10995 195
rect 10855 170 10995 175
rect 10855 150 10905 170
rect 10945 150 10995 170
rect 11035 195 11175 200
rect 11035 175 11050 195
rect 11070 175 11140 195
rect 11160 175 11175 195
rect 11035 170 11175 175
rect 11035 150 11085 170
rect 11125 150 11175 170
rect -310 35 -260 50
rect -220 35 -170 50
rect -130 35 -80 50
rect -40 35 10 50
rect 50 35 100 50
rect 140 35 190 50
rect 230 35 280 50
rect 320 35 370 50
rect 410 35 460 50
rect 500 35 550 50
rect 590 35 640 50
rect 680 35 730 50
rect 770 35 820 50
rect 860 35 910 50
rect 950 35 1000 50
rect 1040 35 1090 50
rect 1130 35 1180 50
rect 1220 35 1270 50
rect 1310 35 1360 50
rect 1400 35 1450 50
rect 1490 35 1540 50
rect 1580 35 1630 50
rect 1670 35 1720 50
rect 1760 35 1810 50
rect 1850 35 1900 50
rect 1940 35 1990 50
rect 2030 35 2080 50
rect 2120 35 2170 50
rect 2210 35 2260 50
rect 2300 35 2350 50
rect 2390 35 2440 50
rect 2480 35 2530 50
rect 2570 35 2620 50
rect 2660 35 2710 50
rect 2750 35 2800 50
rect 2840 35 2890 50
rect 2930 35 2980 50
rect 3020 35 3070 50
rect 3110 35 3160 50
rect 3200 35 3250 50
rect 3290 35 3340 50
rect 3380 35 3430 50
rect 3470 35 3520 50
rect 3560 35 3610 50
rect 3650 35 3700 50
rect 3740 35 3790 50
rect 3830 35 3880 50
rect 3920 35 3970 50
rect 4010 35 4060 50
rect 4100 35 4150 50
rect 4190 35 4240 50
rect 4280 35 4330 50
rect 4370 35 4420 50
rect 4460 35 4510 50
rect 4550 35 4600 50
rect 4640 35 4690 50
rect 4730 35 4780 50
rect 4820 35 4870 50
rect 4910 35 4960 50
rect 5000 35 5050 50
rect 5090 35 5140 50
rect 5180 35 5230 50
rect 5270 35 5320 50
rect 5360 35 5410 50
rect 5450 35 5500 50
rect 5540 35 5590 50
rect 5630 35 5680 50
rect 5720 35 5770 50
rect 5810 35 5860 50
rect 5900 35 5950 50
rect 5990 35 6040 50
rect 6080 35 6130 50
rect 6170 35 6220 50
rect 6260 35 6310 50
rect 6350 35 6400 50
rect 6440 35 6490 50
rect 6530 35 6580 50
rect 6620 35 6670 50
rect 6710 35 6760 50
rect 6800 35 6850 50
rect 6890 35 6940 50
rect 6980 35 7030 50
rect 7070 35 7120 50
rect 7160 35 7210 50
rect 7250 35 7300 50
rect 7340 35 7390 50
rect 7430 35 7480 50
rect 7520 35 7570 50
rect 7610 35 7660 50
rect 7700 35 7750 50
rect 7795 35 7845 50
rect 7885 35 7935 50
rect 7975 35 8025 50
rect 8065 35 8115 50
rect 8155 35 8205 50
rect 8245 35 8295 50
rect 8335 35 8385 50
rect 8425 35 8475 50
rect 8515 35 8565 50
rect 8605 35 8655 50
rect 8695 35 8745 50
rect 8785 35 8835 50
rect 8875 35 8925 50
rect 8965 35 9015 50
rect 9055 35 9105 50
rect 9145 35 9195 50
rect 9235 35 9285 50
rect 9325 35 9375 50
rect 9415 35 9465 50
rect 9505 35 9555 50
rect 9595 35 9645 50
rect 9685 35 9735 50
rect 9775 35 9825 50
rect 9865 35 9915 50
rect 9955 35 10005 50
rect 10045 35 10095 50
rect 10135 35 10185 50
rect 10225 35 10275 50
rect 10315 35 10365 50
rect 10405 35 10455 50
rect 10495 35 10545 50
rect 10585 35 10635 50
rect 10675 35 10725 50
rect 10765 35 10815 50
rect 10855 35 10905 50
rect 10945 35 10995 50
rect 11035 35 11085 50
rect 11125 35 11175 50
<< polycont >>
rect -295 1645 -275 1665
rect -205 1645 -185 1665
rect -115 1645 -95 1665
rect -25 1645 -5 1665
rect 65 1645 85 1665
rect 155 1645 175 1665
rect 245 1645 265 1665
rect 335 1645 355 1665
rect 425 1645 445 1665
rect 515 1645 535 1665
rect 605 1645 625 1665
rect 695 1645 715 1665
rect 785 1645 805 1665
rect 875 1645 895 1665
rect 965 1645 985 1665
rect 1055 1645 1075 1665
rect 1145 1645 1165 1665
rect 1235 1645 1255 1665
rect 1325 1645 1345 1665
rect 1415 1645 1435 1665
rect 1505 1645 1525 1665
rect 1595 1645 1615 1665
rect 1685 1645 1705 1665
rect 1775 1645 1795 1665
rect 1865 1645 1885 1665
rect 1955 1645 1975 1665
rect 2045 1645 2065 1665
rect 2135 1645 2155 1665
rect 2225 1645 2245 1665
rect 2315 1645 2335 1665
rect 2405 1645 2425 1665
rect 2495 1645 2515 1665
rect 2585 1645 2605 1665
rect 2675 1645 2695 1665
rect 2765 1645 2785 1665
rect 2855 1645 2875 1665
rect 2945 1645 2965 1665
rect 3035 1645 3055 1665
rect 3130 1645 3150 1665
rect 3220 1645 3240 1665
rect 3310 1645 3330 1665
rect 3400 1645 3420 1665
rect 3490 1645 3510 1665
rect 3580 1645 3600 1665
rect 3670 1645 3690 1665
rect 3760 1645 3780 1665
rect 3850 1645 3870 1665
rect 3940 1645 3960 1665
rect 4030 1645 4050 1665
rect 4120 1645 4140 1665
rect 4210 1645 4230 1665
rect 4300 1645 4320 1665
rect 4390 1645 4410 1665
rect 4480 1645 4500 1665
rect 4570 1645 4590 1665
rect 4660 1645 4680 1665
rect 4750 1645 4770 1665
rect 4840 1645 4860 1665
rect 4930 1645 4950 1665
rect 5020 1645 5040 1665
rect 5110 1645 5130 1665
rect 5200 1645 5220 1665
rect 5290 1645 5310 1665
rect 5380 1645 5400 1665
rect 5470 1645 5490 1665
rect 5560 1645 5580 1665
rect 5650 1645 5670 1665
rect 5740 1645 5760 1665
rect 5830 1645 5850 1665
rect 5920 1645 5940 1665
rect 6010 1645 6030 1665
rect 6100 1645 6120 1665
rect 6190 1645 6210 1665
rect 6280 1645 6300 1665
rect 6370 1645 6390 1665
rect 6460 1645 6480 1665
rect 6550 1645 6570 1665
rect 6640 1645 6660 1665
rect 6730 1645 6750 1665
rect 6820 1645 6840 1665
rect 6910 1645 6930 1665
rect 7000 1645 7020 1665
rect 7090 1645 7110 1665
rect 7180 1645 7200 1665
rect 7270 1645 7290 1665
rect 7360 1645 7380 1665
rect 7450 1645 7470 1665
rect 7540 1645 7560 1665
rect 7630 1645 7650 1665
rect 7720 1645 7740 1665
rect 7810 1645 7830 1665
rect 7900 1645 7920 1665
rect 7990 1645 8010 1665
rect 8080 1645 8100 1665
rect 8170 1645 8190 1665
rect 8260 1645 8280 1665
rect 8350 1645 8370 1665
rect 8440 1645 8460 1665
rect 8530 1645 8550 1665
rect 8620 1645 8640 1665
rect 8710 1645 8730 1665
rect 8800 1645 8820 1665
rect 8890 1645 8910 1665
rect 8980 1645 9000 1665
rect 9070 1645 9090 1665
rect 9160 1645 9180 1665
rect 9250 1645 9270 1665
rect 9340 1645 9360 1665
rect 9430 1645 9450 1665
rect 9520 1645 9540 1665
rect 9610 1645 9630 1665
rect 9700 1645 9720 1665
rect 9790 1645 9810 1665
rect 9880 1645 9900 1665
rect 9970 1645 9990 1665
rect 10060 1645 10080 1665
rect 10150 1645 10170 1665
rect 10240 1645 10260 1665
rect 10330 1645 10350 1665
rect 10420 1645 10440 1665
rect 10510 1645 10530 1665
rect 10600 1645 10620 1665
rect 10690 1645 10710 1665
rect 10780 1645 10800 1665
rect 10870 1645 10890 1665
rect 10960 1645 10980 1665
rect 11050 1645 11070 1665
rect 11140 1645 11160 1665
rect -295 1115 -275 1135
rect -205 1115 -185 1135
rect -115 1115 -95 1135
rect -25 1115 -5 1135
rect 65 1115 85 1135
rect 155 1115 175 1135
rect 245 1115 265 1135
rect 335 1115 355 1135
rect 425 1115 445 1135
rect 515 1115 535 1135
rect 605 1115 625 1135
rect 695 1115 715 1135
rect 785 1115 805 1135
rect 875 1115 895 1135
rect 965 1115 985 1135
rect 1055 1115 1075 1135
rect 1145 1115 1165 1135
rect 1235 1115 1255 1135
rect 1325 1115 1345 1135
rect 1415 1115 1435 1135
rect 1505 1115 1525 1135
rect 1595 1115 1615 1135
rect 1685 1115 1705 1135
rect 1775 1115 1795 1135
rect 1865 1115 1885 1135
rect 1955 1115 1975 1135
rect 2045 1115 2065 1135
rect 2135 1115 2155 1135
rect 2225 1115 2245 1135
rect 2315 1115 2335 1135
rect 2405 1115 2425 1135
rect 2495 1115 2515 1135
rect 2585 1115 2605 1135
rect 2675 1115 2695 1135
rect 2765 1115 2785 1135
rect 2855 1115 2875 1135
rect 2945 1115 2965 1135
rect 3035 1115 3055 1135
rect 3130 1115 3150 1135
rect 3220 1115 3240 1135
rect 3310 1115 3330 1135
rect 3400 1115 3420 1135
rect 3490 1115 3510 1135
rect 3580 1115 3600 1135
rect 3670 1115 3690 1135
rect 3760 1115 3780 1135
rect 3850 1115 3870 1135
rect 3940 1115 3960 1135
rect 4030 1115 4050 1135
rect 4120 1115 4140 1135
rect 4210 1115 4230 1135
rect 4300 1115 4320 1135
rect 4390 1115 4410 1135
rect 4480 1115 4500 1135
rect 4570 1115 4590 1135
rect 4660 1115 4680 1135
rect 4750 1115 4770 1135
rect 4840 1115 4860 1135
rect 4930 1115 4950 1135
rect 5020 1115 5040 1135
rect 5110 1115 5130 1135
rect 5200 1115 5220 1135
rect 5290 1115 5310 1135
rect 5380 1115 5400 1135
rect 5470 1115 5490 1135
rect 5560 1115 5580 1135
rect 5650 1115 5670 1135
rect 5740 1115 5760 1135
rect 5830 1115 5850 1135
rect 5920 1115 5940 1135
rect 6010 1115 6030 1135
rect 6100 1115 6120 1135
rect 6190 1115 6210 1135
rect 6280 1115 6300 1135
rect 6370 1115 6390 1135
rect 6460 1115 6480 1135
rect 6550 1115 6570 1135
rect 6640 1115 6660 1135
rect 6730 1115 6750 1135
rect 6820 1115 6840 1135
rect 6910 1115 6930 1135
rect 7000 1115 7020 1135
rect 7090 1115 7110 1135
rect 7180 1115 7200 1135
rect 7270 1115 7290 1135
rect 7360 1115 7380 1135
rect 7450 1115 7470 1135
rect 7540 1115 7560 1135
rect 7630 1115 7650 1135
rect 7720 1115 7740 1135
rect 7810 1115 7830 1135
rect 7900 1115 7920 1135
rect 7990 1115 8010 1135
rect 8080 1115 8100 1135
rect 8170 1115 8190 1135
rect 8260 1115 8280 1135
rect 8350 1115 8370 1135
rect 8440 1115 8460 1135
rect 8530 1115 8550 1135
rect 8620 1115 8640 1135
rect 8710 1115 8730 1135
rect 8800 1115 8820 1135
rect 8890 1115 8910 1135
rect 8980 1115 9000 1135
rect 9070 1115 9090 1135
rect 9160 1115 9180 1135
rect 9250 1115 9270 1135
rect 9340 1115 9360 1135
rect 9430 1115 9450 1135
rect 9520 1115 9540 1135
rect 9610 1115 9630 1135
rect 9700 1115 9720 1135
rect 9790 1115 9810 1135
rect 9880 1115 9900 1135
rect 9970 1115 9990 1135
rect 10060 1115 10080 1135
rect 10150 1115 10170 1135
rect 10240 1115 10260 1135
rect 10330 1115 10350 1135
rect 10420 1115 10440 1135
rect 10510 1115 10530 1135
rect 10600 1115 10620 1135
rect 10690 1115 10710 1135
rect 10780 1115 10800 1135
rect 10870 1115 10890 1135
rect 10960 1115 10980 1135
rect 11050 1115 11070 1135
rect 11140 1115 11160 1135
rect -295 705 -275 725
rect -205 705 -185 725
rect -115 705 -95 725
rect -25 705 -5 725
rect 65 705 85 725
rect 155 705 175 725
rect 245 705 265 725
rect 335 705 355 725
rect 425 705 445 725
rect 515 705 535 725
rect 605 705 625 725
rect 695 705 715 725
rect 785 705 805 725
rect 875 705 895 725
rect 965 705 985 725
rect 1055 705 1075 725
rect 1145 705 1165 725
rect 1235 705 1255 725
rect 1325 705 1345 725
rect 1415 705 1435 725
rect 1505 705 1525 725
rect 1595 705 1615 725
rect 1685 705 1705 725
rect 1775 705 1795 725
rect 1865 705 1885 725
rect 1955 705 1975 725
rect 2045 705 2065 725
rect 2135 705 2155 725
rect 2225 705 2245 725
rect 2315 705 2335 725
rect 2405 705 2425 725
rect 2495 705 2515 725
rect 2585 705 2605 725
rect 2675 705 2695 725
rect 2765 705 2785 725
rect 2855 705 2875 725
rect 2945 705 2965 725
rect 3035 705 3055 725
rect 3125 705 3145 725
rect 3215 705 3235 725
rect 3305 705 3325 725
rect 3395 705 3415 725
rect 3485 705 3505 725
rect 3575 705 3595 725
rect 3665 705 3685 725
rect 3755 705 3775 725
rect 3845 705 3865 725
rect 3935 705 3955 725
rect 4025 705 4045 725
rect 4115 705 4135 725
rect 4205 705 4225 725
rect 4295 705 4315 725
rect 4385 705 4405 725
rect 4475 705 4495 725
rect 4565 705 4585 725
rect 4655 705 4675 725
rect 4745 705 4765 725
rect 4835 705 4855 725
rect 4925 705 4945 725
rect 5015 705 5035 725
rect 5105 705 5125 725
rect 5195 705 5215 725
rect 5285 705 5305 725
rect 5375 705 5395 725
rect 5465 705 5485 725
rect 5555 705 5575 725
rect 5645 705 5665 725
rect 5735 705 5755 725
rect 5825 705 5845 725
rect 5915 705 5935 725
rect 6005 705 6025 725
rect 6095 705 6115 725
rect 6185 705 6205 725
rect 6275 705 6295 725
rect 6365 705 6385 725
rect 6455 705 6475 725
rect 6545 705 6565 725
rect 6635 705 6655 725
rect 6725 705 6745 725
rect 6815 705 6835 725
rect 6905 705 6925 725
rect 6995 705 7015 725
rect 7085 705 7105 725
rect 7175 705 7195 725
rect 7265 705 7285 725
rect 7355 705 7375 725
rect 7445 705 7465 725
rect 7535 705 7555 725
rect 7625 705 7645 725
rect 7715 705 7735 725
rect 7810 705 7830 725
rect 7900 705 7920 725
rect 7990 705 8010 725
rect 8080 705 8100 725
rect 8170 705 8190 725
rect 8260 705 8280 725
rect 8350 705 8370 725
rect 8440 705 8460 725
rect 8530 705 8550 725
rect 8620 705 8640 725
rect 8710 705 8730 725
rect 8800 705 8820 725
rect 8890 705 8910 725
rect 8980 705 9000 725
rect 9070 705 9090 725
rect 9160 705 9180 725
rect 9250 705 9270 725
rect 9340 705 9360 725
rect 9430 705 9450 725
rect 9520 705 9540 725
rect 9610 705 9630 725
rect 9700 705 9720 725
rect 9790 705 9810 725
rect 9880 705 9900 725
rect 9970 705 9990 725
rect 10060 705 10080 725
rect 10150 705 10170 725
rect 10240 705 10260 725
rect 10330 705 10350 725
rect 10420 705 10440 725
rect 10510 705 10530 725
rect 10600 705 10620 725
rect 10690 705 10710 725
rect 10780 705 10800 725
rect 10870 705 10890 725
rect 10960 705 10980 725
rect 11050 705 11070 725
rect 11140 705 11160 725
rect -295 175 -275 195
rect -205 175 -185 195
rect -115 175 -95 195
rect -25 175 -5 195
rect 65 175 85 195
rect 155 175 175 195
rect 245 175 265 195
rect 335 175 355 195
rect 425 175 445 195
rect 515 175 535 195
rect 605 175 625 195
rect 695 175 715 195
rect 785 175 805 195
rect 875 175 895 195
rect 965 175 985 195
rect 1055 175 1075 195
rect 1145 175 1165 195
rect 1235 175 1255 195
rect 1325 175 1345 195
rect 1415 175 1435 195
rect 1505 175 1525 195
rect 1595 175 1615 195
rect 1685 175 1705 195
rect 1775 175 1795 195
rect 1865 175 1885 195
rect 1955 175 1975 195
rect 2045 175 2065 195
rect 2135 175 2155 195
rect 2225 175 2245 195
rect 2315 175 2335 195
rect 2405 175 2425 195
rect 2495 175 2515 195
rect 2585 175 2605 195
rect 2675 175 2695 195
rect 2765 175 2785 195
rect 2855 175 2875 195
rect 2945 175 2965 195
rect 3035 175 3055 195
rect 3125 175 3145 195
rect 3215 175 3235 195
rect 3305 175 3325 195
rect 3395 175 3415 195
rect 3485 175 3505 195
rect 3575 175 3595 195
rect 3665 175 3685 195
rect 3755 175 3775 195
rect 3845 175 3865 195
rect 3935 175 3955 195
rect 4025 175 4045 195
rect 4115 175 4135 195
rect 4205 175 4225 195
rect 4295 175 4315 195
rect 4385 175 4405 195
rect 4475 175 4495 195
rect 4565 175 4585 195
rect 4655 175 4675 195
rect 4745 175 4765 195
rect 4835 175 4855 195
rect 4925 175 4945 195
rect 5015 175 5035 195
rect 5105 175 5125 195
rect 5195 175 5215 195
rect 5285 175 5305 195
rect 5375 175 5395 195
rect 5465 175 5485 195
rect 5555 175 5575 195
rect 5645 175 5665 195
rect 5735 175 5755 195
rect 5825 175 5845 195
rect 5915 175 5935 195
rect 6005 175 6025 195
rect 6095 175 6115 195
rect 6185 175 6205 195
rect 6275 175 6295 195
rect 6365 175 6385 195
rect 6455 175 6475 195
rect 6545 175 6565 195
rect 6635 175 6655 195
rect 6725 175 6745 195
rect 6815 175 6835 195
rect 6905 175 6925 195
rect 6995 175 7015 195
rect 7085 175 7105 195
rect 7175 175 7195 195
rect 7265 175 7285 195
rect 7355 175 7375 195
rect 7445 175 7465 195
rect 7535 175 7555 195
rect 7625 175 7645 195
rect 7715 175 7735 195
rect 7810 175 7830 195
rect 7900 175 7920 195
rect 7990 175 8010 195
rect 8080 175 8100 195
rect 8170 175 8190 195
rect 8260 175 8280 195
rect 8350 175 8370 195
rect 8440 175 8460 195
rect 8530 175 8550 195
rect 8620 175 8640 195
rect 8710 175 8730 195
rect 8800 175 8820 195
rect 8890 175 8910 195
rect 8980 175 9000 195
rect 9070 175 9090 195
rect 9160 175 9180 195
rect 9250 175 9270 195
rect 9340 175 9360 195
rect 9430 175 9450 195
rect 9520 175 9540 195
rect 9610 175 9630 195
rect 9700 175 9720 195
rect 9790 175 9810 195
rect 9880 175 9900 195
rect 9970 175 9990 195
rect 10060 175 10080 195
rect 10150 175 10170 195
rect 10240 175 10260 195
rect 10330 175 10350 195
rect 10420 175 10440 195
rect 10510 175 10530 195
rect 10600 175 10620 195
rect 10690 175 10710 195
rect 10780 175 10800 195
rect 10870 175 10890 195
rect 10960 175 10980 195
rect 11050 175 11070 195
rect 11140 175 11160 195
<< locali >>
rect -485 1820 -475 1840
rect -455 1820 -340 1840
rect -320 1820 -295 1840
rect -275 1820 -205 1840
rect -185 1820 -115 1840
rect -95 1820 -25 1840
rect -5 1820 65 1840
rect 85 1820 155 1840
rect 175 1820 200 1840
rect 220 1820 245 1840
rect 265 1820 335 1840
rect 355 1820 380 1840
rect 400 1820 425 1840
rect 445 1820 515 1840
rect 535 1820 560 1840
rect 580 1820 605 1840
rect 625 1820 695 1840
rect 715 1820 740 1840
rect 760 1820 785 1840
rect 805 1820 875 1840
rect 895 1820 920 1840
rect 940 1820 965 1840
rect 985 1820 1055 1840
rect 1075 1820 1100 1840
rect 1120 1820 1145 1840
rect 1165 1820 1235 1840
rect 1255 1820 1280 1840
rect 1300 1820 1325 1840
rect 1345 1820 1415 1840
rect 1435 1820 1460 1840
rect 1480 1820 1505 1840
rect 1525 1820 1595 1840
rect 1615 1820 1640 1840
rect 1660 1820 1685 1840
rect 1705 1820 1775 1840
rect 1795 1820 1820 1840
rect 1840 1820 1865 1840
rect 1885 1820 1955 1840
rect 1975 1820 2000 1840
rect 2020 1820 2045 1840
rect 2065 1820 2135 1840
rect 2155 1820 2180 1840
rect 2200 1820 2225 1840
rect 2245 1820 2315 1840
rect 2335 1820 2360 1840
rect 2380 1820 2405 1840
rect 2425 1820 2495 1840
rect 2515 1820 2540 1840
rect 2560 1820 2585 1840
rect 2605 1820 2675 1840
rect 2695 1820 2720 1840
rect 2740 1820 2765 1840
rect 2785 1820 2855 1840
rect 2875 1820 2900 1840
rect 2920 1820 2945 1840
rect 2965 1820 3035 1840
rect 3055 1820 3085 1840
rect 3105 1820 3130 1840
rect 3150 1820 3220 1840
rect 3240 1820 3265 1840
rect 3285 1820 3310 1840
rect 3330 1820 3400 1840
rect 3420 1820 3445 1840
rect 3465 1820 3490 1840
rect 3510 1820 3580 1840
rect 3600 1820 3625 1840
rect 3645 1820 3670 1840
rect 3690 1820 3760 1840
rect 3780 1820 3805 1840
rect 3825 1820 3850 1840
rect 3870 1820 3940 1840
rect 3960 1820 3985 1840
rect 4005 1820 4030 1840
rect 4050 1820 4120 1840
rect 4140 1820 4165 1840
rect 4185 1820 4210 1840
rect 4230 1820 4300 1840
rect 4320 1820 4345 1840
rect 4365 1820 4390 1840
rect 4410 1820 4480 1840
rect 4500 1820 4525 1840
rect 4545 1820 4570 1840
rect 4590 1820 4660 1840
rect 4680 1820 4705 1840
rect 4725 1820 4750 1840
rect 4770 1820 4840 1840
rect 4860 1820 4885 1840
rect 4905 1820 4930 1840
rect 4950 1820 5020 1840
rect 5040 1820 5065 1840
rect 5085 1820 5110 1840
rect 5130 1820 5200 1840
rect 5220 1820 5245 1840
rect 5265 1820 5290 1840
rect 5310 1820 5380 1840
rect 5400 1820 5425 1840
rect 5445 1820 5470 1840
rect 5490 1820 5560 1840
rect 5580 1820 5605 1840
rect 5625 1820 5650 1840
rect 5670 1820 5740 1840
rect 5760 1820 5785 1840
rect 5805 1820 5830 1840
rect 5850 1820 5920 1840
rect 5940 1820 5965 1840
rect 5985 1820 6010 1840
rect 6030 1820 6100 1840
rect 6120 1820 6145 1840
rect 6165 1820 6190 1840
rect 6210 1820 6280 1840
rect 6300 1820 6325 1840
rect 6345 1820 6370 1840
rect 6390 1820 6460 1840
rect 6480 1820 6505 1840
rect 6525 1820 6550 1840
rect 6570 1820 6640 1840
rect 6660 1820 6685 1840
rect 6705 1820 6730 1840
rect 6750 1820 6820 1840
rect 6840 1820 6865 1840
rect 6885 1820 6910 1840
rect 6930 1820 7000 1840
rect 7020 1820 7045 1840
rect 7065 1820 7090 1840
rect 7110 1820 7180 1840
rect 7200 1820 7225 1840
rect 7245 1820 7270 1840
rect 7290 1820 7360 1840
rect 7380 1820 7405 1840
rect 7425 1820 7450 1840
rect 7470 1820 7540 1840
rect 7560 1820 7585 1840
rect 7605 1820 7630 1840
rect 7650 1820 7720 1840
rect 7740 1820 7765 1840
rect 7785 1820 7810 1840
rect 7830 1820 7900 1840
rect 7920 1820 7945 1840
rect 7965 1820 7990 1840
rect 8010 1820 8080 1840
rect 8100 1820 8125 1840
rect 8145 1820 8170 1840
rect 8190 1820 8260 1840
rect 8280 1820 8305 1840
rect 8325 1820 8350 1840
rect 8370 1820 8440 1840
rect 8460 1820 8485 1840
rect 8505 1820 8530 1840
rect 8550 1820 8620 1840
rect 8640 1820 8665 1840
rect 8685 1820 8710 1840
rect 8730 1820 8800 1840
rect 8820 1820 8845 1840
rect 8865 1820 8890 1840
rect 8910 1820 8980 1840
rect 9000 1820 9025 1840
rect 9045 1820 9070 1840
rect 9090 1820 9160 1840
rect 9180 1820 9205 1840
rect 9225 1820 9250 1840
rect 9270 1820 9340 1840
rect 9360 1820 9385 1840
rect 9405 1820 9430 1840
rect 9450 1820 9520 1840
rect 9540 1820 9565 1840
rect 9585 1820 9610 1840
rect 9630 1820 9700 1840
rect 9720 1820 9745 1840
rect 9765 1820 9790 1840
rect 9810 1820 9880 1840
rect 9900 1820 9925 1840
rect 9945 1820 9970 1840
rect 9990 1820 10060 1840
rect 10080 1820 10105 1840
rect 10125 1820 10150 1840
rect 10170 1820 10240 1840
rect 10260 1820 10285 1840
rect 10305 1820 10330 1840
rect 10350 1820 10420 1840
rect 10440 1820 10465 1840
rect 10485 1820 10510 1840
rect 10530 1820 10600 1840
rect 10620 1820 10645 1840
rect 10665 1820 10690 1840
rect 10710 1820 10780 1840
rect 10800 1820 10870 1840
rect 10890 1820 10960 1840
rect 10980 1820 11050 1840
rect 11070 1820 11140 1840
rect 11160 1820 11185 1840
rect 11205 1820 11320 1840
rect 11340 1820 11350 1840
rect -475 1620 -455 1820
rect -340 1780 -320 1790
rect -340 1690 -320 1700
rect -250 1780 -230 1790
rect -250 1690 -230 1700
rect -160 1780 -140 1790
rect -160 1690 -140 1700
rect -70 1780 -50 1790
rect -70 1665 -50 1700
rect 20 1780 40 1790
rect 20 1690 40 1700
rect 110 1780 130 1790
rect 110 1690 130 1700
rect 200 1780 220 1790
rect 200 1690 220 1700
rect 290 1780 310 1790
rect 290 1690 310 1700
rect 380 1780 400 1790
rect 380 1690 400 1700
rect 470 1780 490 1790
rect 470 1690 490 1700
rect 560 1780 580 1790
rect 560 1690 580 1700
rect 650 1780 670 1790
rect 650 1690 670 1700
rect 740 1780 760 1790
rect 740 1690 760 1700
rect 830 1780 850 1790
rect 830 1690 850 1700
rect 920 1780 940 1790
rect 920 1690 940 1700
rect 1010 1780 1030 1790
rect 1010 1690 1030 1700
rect 1100 1780 1120 1790
rect 1100 1690 1120 1700
rect 1190 1780 1210 1790
rect 1190 1690 1210 1700
rect 1280 1780 1300 1790
rect 1280 1690 1300 1700
rect 1370 1780 1390 1790
rect 1370 1690 1390 1700
rect 1460 1780 1480 1790
rect 1460 1690 1480 1700
rect 1550 1780 1570 1790
rect 1550 1690 1570 1700
rect 1640 1780 1660 1790
rect 1640 1690 1660 1700
rect 1730 1780 1750 1790
rect 1730 1690 1750 1700
rect 1820 1780 1840 1790
rect 1820 1690 1840 1700
rect 1910 1780 1930 1790
rect 1910 1690 1930 1700
rect 2000 1780 2020 1790
rect 2000 1690 2020 1700
rect 2090 1780 2110 1790
rect 2090 1690 2110 1700
rect 2180 1780 2200 1790
rect 2180 1690 2200 1700
rect 2270 1780 2290 1790
rect 2270 1690 2290 1700
rect 2360 1780 2380 1790
rect 2360 1690 2380 1700
rect 2450 1780 2470 1790
rect 2450 1690 2470 1700
rect 2540 1780 2560 1790
rect 2540 1690 2560 1700
rect 2630 1780 2650 1790
rect 2630 1690 2650 1700
rect 2720 1780 2740 1790
rect 2720 1690 2740 1700
rect 2810 1780 2830 1790
rect 2810 1690 2830 1700
rect 2900 1780 2920 1790
rect 2900 1690 2920 1700
rect 2990 1780 3010 1790
rect 2990 1690 3010 1700
rect 3085 1780 3105 1790
rect 3085 1690 3105 1700
rect 3175 1780 3195 1790
rect 3175 1690 3195 1700
rect 3265 1780 3285 1790
rect 3265 1690 3285 1700
rect 3355 1780 3375 1790
rect 3355 1690 3375 1700
rect 3445 1780 3465 1790
rect 3445 1690 3465 1700
rect 3535 1780 3555 1790
rect 3535 1690 3555 1700
rect 3625 1780 3645 1790
rect 3625 1690 3645 1700
rect 3715 1780 3735 1790
rect 3715 1690 3735 1700
rect 3805 1780 3825 1790
rect 3805 1690 3825 1700
rect 3895 1780 3915 1790
rect 3895 1690 3915 1700
rect 3985 1780 4005 1790
rect 3985 1690 4005 1700
rect 4075 1780 4095 1790
rect 4075 1690 4095 1700
rect 4165 1780 4185 1790
rect 4165 1690 4185 1700
rect 4255 1780 4275 1790
rect 4255 1690 4275 1700
rect 4345 1780 4365 1790
rect 4345 1690 4365 1700
rect 4435 1780 4455 1790
rect 4435 1690 4455 1700
rect 4525 1780 4545 1790
rect 4525 1690 4545 1700
rect 4615 1780 4635 1790
rect 4615 1690 4635 1700
rect 4705 1780 4725 1790
rect 4705 1690 4725 1700
rect 4795 1780 4815 1790
rect 4795 1690 4815 1700
rect 4885 1780 4905 1790
rect 4885 1690 4905 1700
rect 4975 1780 4995 1790
rect 4975 1690 4995 1700
rect 5065 1780 5085 1790
rect 5065 1690 5085 1700
rect 5155 1780 5175 1790
rect 5155 1690 5175 1700
rect 5245 1780 5265 1790
rect 5245 1690 5265 1700
rect 5335 1780 5355 1790
rect 5335 1690 5355 1700
rect 5425 1780 5445 1790
rect 5425 1690 5445 1700
rect 5515 1780 5535 1790
rect 5515 1690 5535 1700
rect 5605 1780 5625 1790
rect 5605 1690 5625 1700
rect 5695 1780 5715 1790
rect 5695 1690 5715 1700
rect 5785 1780 5805 1790
rect 5785 1690 5805 1700
rect 5875 1780 5895 1790
rect 5875 1690 5895 1700
rect 5965 1780 5985 1790
rect 5965 1690 5985 1700
rect 6055 1780 6075 1790
rect 6055 1690 6075 1700
rect 6145 1780 6165 1790
rect 6145 1690 6165 1700
rect 6235 1780 6255 1790
rect 6235 1690 6255 1700
rect 6325 1780 6345 1790
rect 6325 1690 6345 1700
rect 6415 1780 6435 1790
rect 6415 1690 6435 1700
rect 6505 1780 6525 1790
rect 6505 1690 6525 1700
rect 6595 1780 6615 1790
rect 6595 1690 6615 1700
rect 6685 1780 6705 1790
rect 6685 1690 6705 1700
rect 6775 1780 6795 1790
rect 6775 1690 6795 1700
rect 6865 1780 6885 1790
rect 6865 1690 6885 1700
rect 6955 1780 6975 1790
rect 6955 1690 6975 1700
rect 7045 1780 7065 1790
rect 7045 1690 7065 1700
rect 7135 1780 7155 1790
rect 7135 1690 7155 1700
rect 7225 1780 7245 1790
rect 7225 1690 7245 1700
rect 7315 1780 7335 1790
rect 7315 1690 7335 1700
rect 7405 1780 7425 1790
rect 7405 1690 7425 1700
rect 7495 1780 7515 1790
rect 7495 1690 7515 1700
rect 7585 1780 7605 1790
rect 7585 1690 7605 1700
rect 7675 1780 7695 1790
rect 7675 1690 7695 1700
rect 7765 1780 7785 1790
rect 7765 1690 7785 1700
rect 7855 1780 7875 1790
rect 7855 1690 7875 1700
rect 7945 1780 7965 1790
rect 7945 1690 7965 1700
rect 8035 1780 8055 1790
rect 8035 1690 8055 1700
rect 8125 1780 8145 1790
rect 8125 1690 8145 1700
rect 8215 1780 8235 1790
rect 8215 1690 8235 1700
rect 8305 1780 8325 1790
rect 8305 1690 8325 1700
rect 8395 1780 8415 1790
rect 8395 1690 8415 1700
rect 8485 1780 8505 1790
rect 8485 1690 8505 1700
rect 8575 1780 8595 1790
rect 8575 1690 8595 1700
rect 8665 1780 8685 1790
rect 8665 1690 8685 1700
rect 8755 1780 8775 1790
rect 8755 1690 8775 1700
rect 8845 1780 8865 1790
rect 8845 1690 8865 1700
rect 8935 1780 8955 1790
rect 8935 1690 8955 1700
rect 9025 1780 9045 1790
rect 9025 1690 9045 1700
rect 9115 1780 9135 1790
rect 9115 1690 9135 1700
rect 9205 1780 9225 1790
rect 9205 1690 9225 1700
rect 9295 1780 9315 1790
rect 9295 1690 9315 1700
rect 9385 1780 9405 1790
rect 9385 1690 9405 1700
rect 9475 1780 9495 1790
rect 9475 1690 9495 1700
rect 9565 1780 9585 1790
rect 9565 1690 9585 1700
rect 9655 1780 9675 1790
rect 9655 1690 9675 1700
rect 9745 1780 9765 1790
rect 9745 1690 9765 1700
rect 9835 1780 9855 1790
rect 9835 1690 9855 1700
rect 9925 1780 9945 1790
rect 9925 1690 9945 1700
rect 10015 1780 10035 1790
rect 10015 1690 10035 1700
rect 10105 1780 10125 1790
rect 10105 1690 10125 1700
rect 10195 1780 10215 1790
rect 10195 1690 10215 1700
rect 10285 1780 10305 1790
rect 10285 1690 10305 1700
rect 10375 1780 10395 1790
rect 10375 1690 10395 1700
rect 10465 1780 10485 1790
rect 10465 1690 10485 1700
rect 10555 1780 10575 1790
rect 10555 1690 10575 1700
rect 10645 1780 10665 1790
rect 10645 1690 10665 1700
rect 10735 1780 10755 1790
rect 10735 1690 10755 1700
rect 10825 1780 10845 1790
rect 10825 1690 10845 1700
rect 10915 1780 10935 1790
rect 10915 1665 10935 1700
rect 11005 1780 11025 1790
rect 11005 1690 11025 1700
rect 11095 1780 11115 1790
rect 11095 1690 11115 1700
rect 11185 1780 11205 1790
rect 11185 1690 11205 1700
rect -305 1645 -295 1665
rect -275 1645 -205 1665
rect -185 1645 -115 1665
rect -95 1645 -25 1665
rect -5 1645 65 1665
rect 85 1645 155 1665
rect 175 1645 185 1665
rect 235 1645 245 1665
rect 265 1645 335 1665
rect 355 1645 365 1665
rect 415 1645 425 1665
rect 445 1645 515 1665
rect 535 1645 545 1665
rect 595 1645 605 1665
rect 625 1645 695 1665
rect 715 1645 725 1665
rect 775 1645 785 1665
rect 805 1645 875 1665
rect 895 1645 905 1665
rect 955 1645 965 1665
rect 985 1645 1055 1665
rect 1075 1645 1085 1665
rect 1135 1645 1145 1665
rect 1165 1645 1235 1665
rect 1255 1645 1265 1665
rect 1315 1645 1325 1665
rect 1345 1645 1415 1665
rect 1435 1645 1445 1665
rect 1495 1645 1505 1665
rect 1525 1645 1595 1665
rect 1615 1645 1625 1665
rect 1675 1645 1685 1665
rect 1705 1645 1775 1665
rect 1795 1645 1805 1665
rect 1855 1645 1865 1665
rect 1885 1645 1955 1665
rect 1975 1645 1985 1665
rect 2035 1645 2045 1665
rect 2065 1645 2135 1665
rect 2155 1645 2165 1665
rect 2215 1645 2225 1665
rect 2245 1645 2315 1665
rect 2335 1645 2345 1665
rect 2395 1645 2405 1665
rect 2425 1645 2495 1665
rect 2515 1645 2525 1665
rect 2575 1645 2585 1665
rect 2605 1645 2675 1665
rect 2695 1645 2705 1665
rect 2755 1645 2765 1665
rect 2785 1645 2855 1665
rect 2875 1645 2885 1665
rect 2935 1645 2945 1665
rect 2965 1645 3035 1665
rect 3055 1645 3065 1665
rect 3120 1645 3130 1665
rect 3150 1645 3220 1665
rect 3240 1645 3250 1665
rect 3300 1645 3310 1665
rect 3330 1645 3400 1665
rect 3420 1645 3430 1665
rect 3480 1645 3490 1665
rect 3510 1645 3580 1665
rect 3600 1645 3610 1665
rect 3660 1645 3670 1665
rect 3690 1645 3760 1665
rect 3780 1645 3790 1665
rect 3840 1645 3850 1665
rect 3870 1645 3940 1665
rect 3960 1645 3970 1665
rect 4020 1645 4030 1665
rect 4050 1645 4120 1665
rect 4140 1645 4150 1665
rect 4200 1645 4210 1665
rect 4230 1645 4300 1665
rect 4320 1645 4330 1665
rect 4380 1645 4390 1665
rect 4410 1645 4480 1665
rect 4500 1645 4510 1665
rect 4560 1645 4570 1665
rect 4590 1645 4660 1665
rect 4680 1645 4690 1665
rect 4740 1645 4750 1665
rect 4770 1645 4840 1665
rect 4860 1645 4870 1665
rect 4920 1645 4930 1665
rect 4950 1645 5020 1665
rect 5040 1645 5050 1665
rect 5100 1645 5110 1665
rect 5130 1645 5200 1665
rect 5220 1645 5230 1665
rect 5280 1645 5290 1665
rect 5310 1645 5380 1665
rect 5400 1645 5410 1665
rect 5460 1645 5470 1665
rect 5490 1645 5560 1665
rect 5580 1645 5590 1665
rect 5640 1645 5650 1665
rect 5670 1645 5740 1665
rect 5760 1645 5770 1665
rect 5820 1645 5830 1665
rect 5850 1645 5920 1665
rect 5940 1645 5950 1665
rect 6000 1645 6010 1665
rect 6030 1645 6100 1665
rect 6120 1645 6130 1665
rect 6180 1645 6190 1665
rect 6210 1645 6280 1665
rect 6300 1645 6310 1665
rect 6360 1645 6370 1665
rect 6390 1645 6460 1665
rect 6480 1645 6490 1665
rect 6540 1645 6550 1665
rect 6570 1645 6640 1665
rect 6660 1645 6670 1665
rect 6720 1645 6730 1665
rect 6750 1645 6820 1665
rect 6840 1645 6850 1665
rect 6900 1645 6910 1665
rect 6930 1645 7000 1665
rect 7020 1645 7030 1665
rect 7080 1645 7090 1665
rect 7110 1645 7180 1665
rect 7200 1645 7210 1665
rect 7260 1645 7270 1665
rect 7290 1645 7360 1665
rect 7380 1645 7390 1665
rect 7440 1645 7450 1665
rect 7470 1645 7540 1665
rect 7560 1645 7570 1665
rect 7620 1645 7630 1665
rect 7650 1645 7720 1665
rect 7740 1645 7750 1665
rect 7800 1645 7810 1665
rect 7830 1645 7900 1665
rect 7920 1645 7930 1665
rect 7980 1645 7990 1665
rect 8010 1645 8080 1665
rect 8100 1645 8110 1665
rect 8160 1645 8170 1665
rect 8190 1645 8260 1665
rect 8280 1645 8290 1665
rect 8340 1645 8350 1665
rect 8370 1645 8440 1665
rect 8460 1645 8470 1665
rect 8520 1645 8530 1665
rect 8550 1645 8620 1665
rect 8640 1645 8650 1665
rect 8700 1645 8710 1665
rect 8730 1645 8800 1665
rect 8820 1645 8830 1665
rect 8880 1645 8890 1665
rect 8910 1645 8980 1665
rect 9000 1645 9010 1665
rect 9060 1645 9070 1665
rect 9090 1645 9160 1665
rect 9180 1645 9190 1665
rect 9240 1645 9250 1665
rect 9270 1645 9340 1665
rect 9360 1645 9370 1665
rect 9420 1645 9430 1665
rect 9450 1645 9520 1665
rect 9540 1645 9550 1665
rect 9600 1645 9610 1665
rect 9630 1645 9700 1665
rect 9720 1645 9730 1665
rect 9780 1645 9790 1665
rect 9810 1645 9880 1665
rect 9900 1645 9910 1665
rect 9960 1645 9970 1665
rect 9990 1645 10060 1665
rect 10080 1645 10090 1665
rect 10140 1645 10150 1665
rect 10170 1645 10240 1665
rect 10260 1645 10270 1665
rect 10320 1645 10330 1665
rect 10350 1645 10420 1665
rect 10440 1645 10450 1665
rect 10500 1645 10510 1665
rect 10530 1645 10600 1665
rect 10620 1645 10630 1665
rect 10680 1645 10690 1665
rect 10710 1645 10780 1665
rect 10800 1645 10870 1665
rect 10890 1645 10960 1665
rect 10980 1645 11050 1665
rect 11070 1645 11140 1665
rect 11160 1645 11170 1665
rect 11320 1620 11340 1820
rect -475 1600 -295 1620
rect -275 1600 -205 1620
rect -185 1600 -115 1620
rect -95 1600 -25 1620
rect -5 1600 65 1620
rect 85 1600 155 1620
rect 175 1600 245 1620
rect 265 1600 335 1620
rect 355 1600 425 1620
rect 445 1600 515 1620
rect 535 1600 605 1620
rect 625 1600 695 1620
rect 715 1600 785 1620
rect 805 1600 875 1620
rect 895 1600 965 1620
rect 985 1600 1055 1620
rect 1075 1600 1145 1620
rect 1165 1600 1235 1620
rect 1255 1600 1325 1620
rect 1345 1600 1415 1620
rect 1435 1600 1505 1620
rect 1525 1600 1595 1620
rect 1615 1600 1685 1620
rect 1705 1600 1775 1620
rect 1795 1600 1865 1620
rect 1885 1600 1955 1620
rect 1975 1600 2045 1620
rect 2065 1600 2135 1620
rect 2155 1600 2225 1620
rect 2245 1600 2315 1620
rect 2335 1600 2405 1620
rect 2425 1600 2495 1620
rect 2515 1600 2585 1620
rect 2605 1600 2675 1620
rect 2695 1600 2765 1620
rect 2785 1600 2855 1620
rect 2875 1600 2945 1620
rect 2965 1600 3035 1620
rect 3055 1600 3130 1620
rect 3150 1600 3220 1620
rect 3240 1600 3310 1620
rect 3330 1600 3400 1620
rect 3420 1600 3490 1620
rect 3510 1600 3580 1620
rect 3600 1600 3670 1620
rect 3690 1600 3760 1620
rect 3780 1600 3850 1620
rect 3870 1600 3940 1620
rect 3960 1600 4030 1620
rect 4050 1600 4120 1620
rect 4140 1600 4210 1620
rect 4230 1600 4300 1620
rect 4320 1600 4390 1620
rect 4410 1600 4480 1620
rect 4500 1600 4570 1620
rect 4590 1600 4660 1620
rect 4680 1600 4750 1620
rect 4770 1600 4840 1620
rect 4860 1600 4930 1620
rect 4950 1600 5020 1620
rect 5040 1600 5110 1620
rect 5130 1600 5200 1620
rect 5220 1600 5290 1620
rect 5310 1600 5380 1620
rect 5400 1600 5470 1620
rect 5490 1600 5560 1620
rect 5580 1600 5650 1620
rect 5670 1600 5740 1620
rect 5760 1600 5830 1620
rect 5850 1600 5920 1620
rect 5940 1600 6010 1620
rect 6030 1600 6100 1620
rect 6120 1600 6190 1620
rect 6210 1600 6280 1620
rect 6300 1600 6370 1620
rect 6390 1600 6460 1620
rect 6480 1600 6550 1620
rect 6570 1600 6640 1620
rect 6660 1600 6730 1620
rect 6750 1600 6820 1620
rect 6840 1600 6910 1620
rect 6930 1600 7000 1620
rect 7020 1600 7090 1620
rect 7110 1600 7180 1620
rect 7200 1600 7270 1620
rect 7290 1600 7360 1620
rect 7380 1600 7450 1620
rect 7470 1600 7540 1620
rect 7560 1600 7630 1620
rect 7650 1600 7720 1620
rect 7740 1600 7810 1620
rect 7830 1600 7900 1620
rect 7920 1600 7990 1620
rect 8010 1600 8080 1620
rect 8100 1600 8170 1620
rect 8190 1600 8260 1620
rect 8280 1600 8350 1620
rect 8370 1600 8440 1620
rect 8460 1600 8530 1620
rect 8550 1600 8620 1620
rect 8640 1600 8710 1620
rect 8730 1600 8800 1620
rect 8820 1600 8890 1620
rect 8910 1600 8980 1620
rect 9000 1600 9070 1620
rect 9090 1600 9160 1620
rect 9180 1600 9250 1620
rect 9270 1600 9340 1620
rect 9360 1600 9430 1620
rect 9450 1600 9520 1620
rect 9540 1600 9610 1620
rect 9630 1600 9700 1620
rect 9720 1600 9790 1620
rect 9810 1600 9880 1620
rect 9900 1600 9970 1620
rect 9990 1600 10060 1620
rect 10080 1600 10150 1620
rect 10170 1600 10240 1620
rect 10260 1600 10330 1620
rect 10350 1600 10420 1620
rect 10440 1600 10510 1620
rect 10530 1600 10600 1620
rect 10620 1600 10690 1620
rect 10710 1600 10780 1620
rect 10800 1600 10870 1620
rect 10890 1600 10960 1620
rect 10980 1600 11050 1620
rect 11070 1600 11140 1620
rect 11160 1600 11340 1620
rect -350 1560 110 1580
rect 130 1560 6820 1580
rect 6840 1560 10510 1580
rect 10530 1560 10555 1580
rect 10575 1560 11215 1580
rect -350 1520 20 1540
rect 40 1520 335 1540
rect 355 1520 515 1540
rect 535 1520 695 1540
rect 715 1520 875 1540
rect 895 1520 1055 1540
rect 1075 1520 1235 1540
rect 1255 1520 1415 1540
rect 1435 1520 1595 1540
rect 1615 1520 7945 1540
rect 7965 1520 8665 1540
rect 8685 1520 9385 1540
rect 9405 1520 10105 1540
rect 10125 1520 11215 1540
rect -350 1480 -70 1500
rect -50 1480 4660 1500
rect 4680 1480 4840 1500
rect 4860 1480 5020 1500
rect 5040 1480 5200 1500
rect 5220 1480 5380 1500
rect 5400 1480 5560 1500
rect 5580 1480 5740 1500
rect 5760 1480 5920 1500
rect 5940 1480 8080 1500
rect 8100 1480 8260 1500
rect 8280 1480 8305 1500
rect 8325 1480 8440 1500
rect 8460 1480 8620 1500
rect 8640 1480 11215 1500
rect -350 1440 -160 1460
rect -140 1440 7720 1460
rect 7740 1440 7900 1460
rect 7920 1440 8800 1460
rect 8820 1440 8980 1460
rect 9000 1440 9160 1460
rect 9180 1440 9340 1460
rect 9360 1440 9385 1460
rect 9405 1440 9520 1460
rect 9540 1440 9700 1460
rect 9720 1440 9745 1460
rect 9765 1440 9880 1460
rect 9900 1440 10060 1460
rect 10080 1440 10105 1460
rect 10125 1440 10240 1460
rect 10260 1440 10420 1460
rect 10440 1440 11215 1460
rect -350 1400 -250 1420
rect -230 1400 1775 1420
rect 1795 1400 1955 1420
rect 1975 1400 2135 1420
rect 2155 1400 2315 1420
rect 2335 1400 2495 1420
rect 2515 1400 2675 1420
rect 2695 1400 2855 1420
rect 2875 1400 3035 1420
rect 3055 1400 3220 1420
rect 3240 1400 3400 1420
rect 3420 1400 3580 1420
rect 3600 1400 3760 1420
rect 3780 1400 3940 1420
rect 3960 1400 4120 1420
rect 4140 1400 4300 1420
rect 4320 1400 4480 1420
rect 4500 1400 6100 1420
rect 6120 1400 6280 1420
rect 6300 1400 6460 1420
rect 6480 1400 6640 1420
rect 6660 1400 6685 1420
rect 6705 1400 6730 1420
rect 6750 1400 6865 1420
rect 6885 1400 7000 1420
rect 7020 1400 7180 1420
rect 7200 1400 7360 1420
rect 7380 1400 7540 1420
rect 7560 1400 10600 1420
rect 10620 1400 11215 1420
rect -350 1360 920 1380
rect 940 1360 11005 1380
rect 11025 1360 11215 1380
rect -350 1320 605 1340
rect 625 1320 785 1340
rect 805 1320 965 1340
rect 985 1320 1145 1340
rect 1165 1320 1685 1340
rect 1705 1320 1865 1340
rect 1885 1320 2000 1340
rect 2020 1320 2045 1340
rect 2065 1320 2225 1340
rect 2245 1320 2360 1340
rect 2380 1320 2405 1340
rect 2425 1320 2585 1340
rect 2605 1320 2720 1340
rect 2740 1320 2765 1340
rect 2785 1320 2945 1340
rect 2965 1320 3490 1340
rect 3510 1320 3670 1340
rect 3690 1320 3850 1340
rect 3870 1320 4030 1340
rect 4050 1320 4930 1340
rect 4950 1320 5110 1340
rect 5130 1320 5290 1340
rect 5310 1320 5470 1340
rect 5490 1320 6370 1340
rect 6390 1320 6550 1340
rect 6570 1320 6910 1340
rect 6930 1320 7090 1340
rect 7110 1320 7990 1340
rect 8010 1320 8170 1340
rect 8190 1320 8350 1340
rect 8370 1320 8530 1340
rect 8550 1320 9250 1340
rect 9270 1320 9430 1340
rect 9450 1320 9970 1340
rect 9990 1320 10150 1340
rect 10170 1320 10915 1340
rect 10935 1320 11215 1340
rect -350 1280 245 1300
rect 265 1280 425 1300
rect 445 1280 1325 1300
rect 1345 1280 1505 1300
rect 1525 1280 3805 1300
rect 3825 1280 6010 1300
rect 6030 1280 6190 1300
rect 6210 1280 6775 1300
rect 6795 1280 7270 1300
rect 7290 1280 7450 1300
rect 7470 1280 7630 1300
rect 7650 1280 7810 1300
rect 7830 1280 8710 1300
rect 8730 1280 8890 1300
rect 8910 1280 9070 1300
rect 9090 1280 9610 1300
rect 9630 1280 9790 1300
rect 9810 1280 10330 1300
rect 10350 1280 10825 1300
rect 10845 1280 11215 1300
rect -475 1240 -295 1260
rect -275 1240 -205 1260
rect -185 1240 -115 1260
rect -95 1240 -25 1260
rect -5 1240 65 1260
rect 85 1240 155 1260
rect 175 1240 245 1260
rect 265 1240 335 1260
rect 355 1240 425 1260
rect 445 1240 515 1260
rect 535 1240 605 1260
rect 625 1240 695 1260
rect 715 1240 785 1260
rect 805 1240 875 1260
rect 895 1240 965 1260
rect 985 1240 1055 1260
rect 1075 1240 1145 1260
rect 1165 1240 1235 1260
rect 1255 1240 1325 1260
rect 1345 1240 1415 1260
rect 1435 1240 1505 1260
rect 1525 1240 1595 1260
rect 1615 1240 1685 1260
rect 1705 1240 1775 1260
rect 1795 1240 1865 1260
rect 1885 1240 1955 1260
rect 1975 1240 2045 1260
rect 2065 1240 2135 1260
rect 2155 1240 2225 1260
rect 2245 1240 2315 1260
rect 2335 1240 2405 1260
rect 2425 1240 2495 1260
rect 2515 1240 2585 1260
rect 2605 1240 2675 1260
rect 2695 1240 2765 1260
rect 2785 1240 2855 1260
rect 2875 1240 2945 1260
rect 2965 1240 3035 1260
rect 3055 1240 3130 1260
rect 3150 1240 3220 1260
rect 3240 1240 3310 1260
rect 3330 1240 3400 1260
rect 3420 1240 3490 1260
rect 3510 1240 3580 1260
rect 3600 1240 3670 1260
rect 3690 1240 3760 1260
rect 3780 1240 3850 1260
rect 3870 1240 3940 1260
rect 3960 1240 4030 1260
rect 4050 1240 4120 1260
rect 4140 1240 4210 1260
rect 4230 1240 4300 1260
rect 4320 1240 4390 1260
rect 4410 1240 4480 1260
rect 4500 1240 4570 1260
rect 4590 1240 4660 1260
rect 4680 1240 4750 1260
rect 4770 1240 4840 1260
rect 4860 1240 4930 1260
rect 4950 1240 5020 1260
rect 5040 1240 5110 1260
rect 5130 1240 5200 1260
rect 5220 1240 5290 1260
rect 5310 1240 5380 1260
rect 5400 1240 5470 1260
rect 5490 1240 5560 1260
rect 5580 1240 5650 1260
rect 5670 1240 5740 1260
rect 5760 1240 5830 1260
rect 5850 1240 5920 1260
rect 5940 1240 6010 1260
rect 6030 1240 6100 1260
rect 6120 1240 6190 1260
rect 6210 1240 6280 1260
rect 6300 1240 6370 1260
rect 6390 1240 6460 1260
rect 6480 1240 6550 1260
rect 6570 1240 6640 1260
rect 6660 1240 6730 1260
rect 6750 1240 6820 1260
rect 6840 1240 6910 1260
rect 6930 1240 7000 1260
rect 7020 1240 7090 1260
rect 7110 1240 7180 1260
rect 7200 1240 7270 1260
rect 7290 1240 7360 1260
rect 7380 1240 7450 1260
rect 7470 1240 7540 1260
rect 7560 1240 7630 1260
rect 7650 1240 7720 1260
rect 7740 1240 7810 1260
rect 7830 1240 7900 1260
rect 7920 1240 7990 1260
rect 8010 1240 8080 1260
rect 8100 1240 8170 1260
rect 8190 1240 8260 1260
rect 8280 1240 8350 1260
rect 8370 1240 8440 1260
rect 8460 1240 8530 1260
rect 8550 1240 8620 1260
rect 8640 1240 8710 1260
rect 8730 1240 8800 1260
rect 8820 1240 8890 1260
rect 8910 1240 8980 1260
rect 9000 1240 9070 1260
rect 9090 1240 9160 1260
rect 9180 1240 9250 1260
rect 9270 1240 9340 1260
rect 9360 1240 9430 1260
rect 9450 1240 9520 1260
rect 9540 1240 9610 1260
rect 9630 1240 9700 1260
rect 9720 1240 9790 1260
rect 9810 1240 9880 1260
rect 9900 1240 9970 1260
rect 9990 1240 10060 1260
rect 10080 1240 10150 1260
rect 10170 1240 10240 1260
rect 10260 1240 10330 1260
rect 10350 1240 10420 1260
rect 10440 1240 10510 1260
rect 10530 1240 10600 1260
rect 10620 1240 10690 1260
rect 10710 1240 10780 1260
rect 10800 1240 10870 1260
rect 10890 1240 10960 1260
rect 10980 1240 11050 1260
rect 11070 1240 11140 1260
rect 11160 1240 11340 1260
rect -475 600 -455 1240
rect -350 1200 3130 1220
rect 3150 1200 3310 1220
rect 3330 1200 4210 1220
rect 4230 1200 4390 1220
rect 4410 1200 4570 1220
rect 4590 1200 4750 1220
rect 4770 1200 5245 1220
rect 5265 1200 5650 1220
rect 5670 1200 5830 1220
rect 5850 1200 10735 1220
rect 10755 1200 11215 1220
rect -400 1160 -295 1180
rect -275 1160 -205 1180
rect -185 1160 -115 1180
rect -95 1160 -25 1180
rect -5 1160 65 1180
rect 85 1160 155 1180
rect 175 1160 245 1180
rect 265 1160 335 1180
rect 355 1160 425 1180
rect 445 1160 515 1180
rect 535 1160 605 1180
rect 625 1160 695 1180
rect 715 1160 785 1180
rect 805 1160 875 1180
rect 895 1160 965 1180
rect 985 1160 1055 1180
rect 1075 1160 1145 1180
rect 1165 1160 1235 1180
rect 1255 1160 1325 1180
rect 1345 1160 1415 1180
rect 1435 1160 1505 1180
rect 1525 1160 1595 1180
rect 1615 1160 1685 1180
rect 1705 1160 1775 1180
rect 1795 1160 1865 1180
rect 1885 1160 1955 1180
rect 1975 1160 2045 1180
rect 2065 1160 2135 1180
rect 2155 1160 2225 1180
rect 2245 1160 2315 1180
rect 2335 1160 2405 1180
rect 2425 1160 2495 1180
rect 2515 1160 2585 1180
rect 2605 1160 2675 1180
rect 2695 1160 2765 1180
rect 2785 1160 2855 1180
rect 2875 1160 2945 1180
rect 2965 1160 3035 1180
rect 3055 1160 3130 1180
rect 3150 1160 3220 1180
rect 3240 1160 3310 1180
rect 3330 1160 3400 1180
rect 3420 1160 3490 1180
rect 3510 1160 3580 1180
rect 3600 1160 3670 1180
rect 3690 1160 3760 1180
rect 3780 1160 3850 1180
rect 3870 1160 3940 1180
rect 3960 1160 4030 1180
rect 4050 1160 4120 1180
rect 4140 1160 4210 1180
rect 4230 1160 4300 1180
rect 4320 1160 4390 1180
rect 4410 1160 4480 1180
rect 4500 1160 4570 1180
rect 4590 1160 4660 1180
rect 4680 1160 4750 1180
rect 4770 1160 4840 1180
rect 4860 1160 4930 1180
rect 4950 1160 5020 1180
rect 5040 1160 5110 1180
rect 5130 1160 5200 1180
rect 5220 1160 5290 1180
rect 5310 1160 5380 1180
rect 5400 1160 5470 1180
rect 5490 1160 5560 1180
rect 5580 1160 5650 1180
rect 5670 1160 5740 1180
rect 5760 1160 5830 1180
rect 5850 1160 5920 1180
rect 5940 1160 6010 1180
rect 6030 1160 6100 1180
rect 6120 1160 6190 1180
rect 6210 1160 6280 1180
rect 6300 1160 6370 1180
rect 6390 1160 6460 1180
rect 6480 1160 6550 1180
rect 6570 1160 6640 1180
rect 6660 1160 6730 1180
rect 6750 1160 6820 1180
rect 6840 1160 6910 1180
rect 6930 1160 7000 1180
rect 7020 1160 7090 1180
rect 7110 1160 7180 1180
rect 7200 1160 7270 1180
rect 7290 1160 7360 1180
rect 7380 1160 7450 1180
rect 7470 1160 7540 1180
rect 7560 1160 7630 1180
rect 7650 1160 7720 1180
rect 7740 1160 7810 1180
rect 7830 1160 7900 1180
rect 7920 1160 7990 1180
rect 8010 1160 8080 1180
rect 8100 1160 8170 1180
rect 8190 1160 8260 1180
rect 8280 1160 8350 1180
rect 8370 1160 8440 1180
rect 8460 1160 8530 1180
rect 8550 1160 8620 1180
rect 8640 1160 8710 1180
rect 8730 1160 8800 1180
rect 8820 1160 8890 1180
rect 8910 1160 8980 1180
rect 9000 1160 9070 1180
rect 9090 1160 9160 1180
rect 9180 1160 9250 1180
rect 9270 1160 9340 1180
rect 9360 1160 9430 1180
rect 9450 1160 9520 1180
rect 9540 1160 9610 1180
rect 9630 1160 9700 1180
rect 9720 1160 9790 1180
rect 9810 1160 9880 1180
rect 9900 1160 9970 1180
rect 9990 1160 10060 1180
rect 10080 1160 10150 1180
rect 10170 1160 10240 1180
rect 10260 1160 10330 1180
rect 10350 1160 10420 1180
rect 10440 1160 10510 1180
rect 10530 1160 10600 1180
rect 10620 1160 10690 1180
rect 10710 1160 10780 1180
rect 10800 1160 10870 1180
rect 10890 1160 10960 1180
rect 10980 1160 11050 1180
rect 11070 1160 11140 1180
rect 11160 1160 11265 1180
rect -400 960 -380 1160
rect -305 1115 -295 1135
rect -275 1115 -205 1135
rect -185 1115 -115 1135
rect -95 1115 -25 1135
rect -5 1115 65 1135
rect 85 1115 155 1135
rect 175 1115 190 1135
rect 235 1115 245 1135
rect 265 1115 335 1135
rect 355 1115 365 1135
rect 415 1115 425 1135
rect 445 1115 515 1135
rect 535 1115 545 1135
rect 595 1115 605 1135
rect 625 1115 695 1135
rect 715 1115 725 1135
rect 775 1115 785 1135
rect 805 1115 875 1135
rect 895 1115 905 1135
rect 955 1115 965 1135
rect 985 1115 1055 1135
rect 1075 1115 1085 1135
rect 1135 1115 1145 1135
rect 1165 1115 1235 1135
rect 1255 1115 1265 1135
rect 1315 1115 1325 1135
rect 1345 1115 1415 1135
rect 1435 1115 1445 1135
rect 1495 1115 1505 1135
rect 1525 1115 1595 1135
rect 1615 1115 1625 1135
rect 1675 1115 1685 1135
rect 1705 1115 1775 1135
rect 1795 1115 1805 1135
rect 1855 1115 1865 1135
rect 1885 1115 1955 1135
rect 1975 1115 1985 1135
rect 2035 1115 2045 1135
rect 2065 1115 2135 1135
rect 2155 1115 2165 1135
rect 2215 1115 2225 1135
rect 2245 1115 2315 1135
rect 2335 1115 2345 1135
rect 2395 1115 2405 1135
rect 2425 1115 2495 1135
rect 2515 1115 2525 1135
rect 2575 1115 2585 1135
rect 2605 1115 2675 1135
rect 2695 1115 2705 1135
rect 2755 1115 2765 1135
rect 2785 1115 2855 1135
rect 2875 1115 2885 1135
rect 2935 1115 2945 1135
rect 2965 1115 3035 1135
rect 3055 1115 3065 1135
rect 3120 1115 3130 1135
rect 3150 1115 3220 1135
rect 3240 1115 3250 1135
rect 3300 1115 3310 1135
rect 3330 1115 3400 1135
rect 3420 1115 3430 1135
rect 3480 1115 3490 1135
rect 3510 1115 3580 1135
rect 3600 1115 3610 1135
rect 3660 1115 3670 1135
rect 3690 1115 3760 1135
rect 3780 1115 3790 1135
rect 3840 1115 3850 1135
rect 3870 1115 3940 1135
rect 3960 1115 3970 1135
rect 4020 1115 4030 1135
rect 4050 1115 4120 1135
rect 4140 1115 4150 1135
rect 4200 1115 4210 1135
rect 4230 1115 4300 1135
rect 4320 1115 4330 1135
rect 4380 1115 4390 1135
rect 4410 1115 4480 1135
rect 4500 1115 4510 1135
rect 4560 1115 4570 1135
rect 4590 1115 4660 1135
rect 4680 1115 4690 1135
rect 4740 1115 4750 1135
rect 4770 1115 4840 1135
rect 4860 1115 4870 1135
rect 4920 1115 4930 1135
rect 4950 1115 5020 1135
rect 5040 1115 5050 1135
rect 5100 1115 5110 1135
rect 5130 1115 5200 1135
rect 5220 1115 5230 1135
rect 5280 1115 5290 1135
rect 5310 1115 5380 1135
rect 5400 1115 5410 1135
rect 5460 1115 5470 1135
rect 5490 1115 5560 1135
rect 5580 1115 5590 1135
rect 5640 1115 5650 1135
rect 5670 1115 5740 1135
rect 5760 1115 5770 1135
rect 5820 1115 5830 1135
rect 5850 1115 5920 1135
rect 5940 1115 5950 1135
rect 6000 1115 6010 1135
rect 6030 1115 6100 1135
rect 6120 1115 6130 1135
rect 6180 1115 6190 1135
rect 6210 1115 6280 1135
rect 6300 1115 6310 1135
rect 6360 1115 6370 1135
rect 6390 1115 6460 1135
rect 6480 1115 6490 1135
rect 6540 1115 6550 1135
rect 6570 1115 6640 1135
rect 6660 1115 6670 1135
rect 6720 1115 6730 1135
rect 6750 1115 6820 1135
rect 6840 1115 6850 1135
rect 6900 1115 6910 1135
rect 6930 1115 7000 1135
rect 7020 1115 7030 1135
rect 7080 1115 7090 1135
rect 7110 1115 7180 1135
rect 7200 1115 7210 1135
rect 7260 1115 7270 1135
rect 7290 1115 7360 1135
rect 7380 1115 7390 1135
rect 7440 1115 7450 1135
rect 7470 1115 7540 1135
rect 7560 1115 7570 1135
rect 7620 1115 7630 1135
rect 7650 1115 7720 1135
rect 7740 1115 7750 1135
rect 7800 1115 7810 1135
rect 7830 1115 7900 1135
rect 7920 1115 7930 1135
rect 7980 1115 7990 1135
rect 8010 1115 8080 1135
rect 8100 1115 8110 1135
rect 8160 1115 8170 1135
rect 8190 1115 8260 1135
rect 8280 1115 8290 1135
rect 8340 1115 8350 1135
rect 8370 1115 8440 1135
rect 8460 1115 8470 1135
rect 8520 1115 8530 1135
rect 8550 1115 8620 1135
rect 8640 1115 8650 1135
rect 8700 1115 8710 1135
rect 8730 1115 8800 1135
rect 8820 1115 8830 1135
rect 8880 1115 8890 1135
rect 8910 1115 8980 1135
rect 9000 1115 9010 1135
rect 9060 1115 9070 1135
rect 9090 1115 9160 1135
rect 9180 1115 9190 1135
rect 9240 1115 9250 1135
rect 9270 1115 9340 1135
rect 9360 1115 9370 1135
rect 9420 1115 9430 1135
rect 9450 1115 9520 1135
rect 9540 1115 9550 1135
rect 9600 1115 9610 1135
rect 9630 1115 9700 1135
rect 9720 1115 9730 1135
rect 9780 1115 9790 1135
rect 9810 1115 9880 1135
rect 9900 1115 9910 1135
rect 9960 1115 9970 1135
rect 9990 1115 10060 1135
rect 10080 1115 10090 1135
rect 10140 1115 10150 1135
rect 10170 1115 10240 1135
rect 10260 1115 10270 1135
rect 10320 1115 10330 1135
rect 10350 1115 10420 1135
rect 10440 1115 10450 1135
rect 10500 1115 10510 1135
rect 10530 1115 10600 1135
rect 10620 1115 10635 1135
rect 10675 1115 10690 1135
rect 10710 1115 10780 1135
rect 10800 1115 10870 1135
rect 10890 1115 10960 1135
rect 10980 1115 11050 1135
rect 11070 1115 11140 1135
rect 11160 1115 11170 1135
rect -340 1080 -320 1090
rect -340 990 -320 1000
rect -250 1080 -230 1090
rect -250 990 -230 1000
rect -160 1080 -140 1090
rect -160 990 -140 1000
rect -70 1080 -50 1115
rect -70 990 -50 1000
rect 20 1080 40 1090
rect 20 990 40 1000
rect 110 1080 130 1090
rect 110 990 130 1000
rect 200 1080 220 1090
rect 200 990 220 1000
rect 290 1080 310 1090
rect 290 990 310 1000
rect 380 1080 400 1090
rect 380 990 400 1000
rect 470 1080 490 1090
rect 470 990 490 1000
rect 560 1080 580 1090
rect 560 990 580 1000
rect 650 1080 670 1090
rect 650 990 670 1000
rect 740 1080 760 1090
rect 740 990 760 1000
rect 830 1080 850 1090
rect 830 990 850 1000
rect 920 1080 940 1090
rect 920 990 940 1000
rect 1010 1080 1030 1090
rect 1010 990 1030 1000
rect 1100 1080 1120 1090
rect 1100 990 1120 1000
rect 1190 1080 1210 1090
rect 1190 990 1210 1000
rect 1280 1080 1300 1090
rect 1280 990 1300 1000
rect 1370 1080 1390 1090
rect 1370 990 1390 1000
rect 1460 1080 1480 1090
rect 1460 990 1480 1000
rect 1550 1080 1570 1090
rect 1550 990 1570 1000
rect 1640 1080 1660 1090
rect 1640 990 1660 1000
rect 1730 1080 1750 1090
rect 1730 990 1750 1000
rect 1820 1080 1840 1090
rect 1820 990 1840 1000
rect 1910 1080 1930 1090
rect 1910 990 1930 1000
rect 2000 1080 2020 1090
rect 2000 990 2020 1000
rect 2090 1080 2110 1090
rect 2090 990 2110 1000
rect 2180 1080 2200 1090
rect 2180 990 2200 1000
rect 2270 1080 2290 1090
rect 2270 990 2290 1000
rect 2360 1080 2380 1090
rect 2360 990 2380 1000
rect 2450 1080 2470 1090
rect 2450 990 2470 1000
rect 2540 1080 2560 1090
rect 2540 990 2560 1000
rect 2630 1080 2650 1090
rect 2630 990 2650 1000
rect 2720 1080 2740 1090
rect 2720 990 2740 1000
rect 2810 1080 2830 1090
rect 2810 990 2830 1000
rect 2900 1080 2920 1090
rect 2900 990 2920 1000
rect 2990 1080 3010 1090
rect 2990 990 3010 1000
rect 3085 1080 3105 1090
rect 3085 990 3105 1000
rect 3175 1080 3195 1090
rect 3175 990 3195 1000
rect 3265 1080 3285 1090
rect 3265 990 3285 1000
rect 3355 1080 3375 1090
rect 3355 990 3375 1000
rect 3445 1080 3465 1090
rect 3445 990 3465 1000
rect 3535 1080 3555 1090
rect 3535 990 3555 1000
rect 3625 1080 3645 1090
rect 3625 990 3645 1000
rect 3715 1080 3735 1090
rect 3715 990 3735 1000
rect 3805 1080 3825 1090
rect 3805 990 3825 1000
rect 3895 1080 3915 1090
rect 3895 990 3915 1000
rect 3985 1080 4005 1090
rect 3985 990 4005 1000
rect 4075 1080 4095 1090
rect 4075 990 4095 1000
rect 4165 1080 4185 1090
rect 4165 990 4185 1000
rect 4255 1080 4275 1090
rect 4255 990 4275 1000
rect 4345 1080 4365 1090
rect 4345 990 4365 1000
rect 4435 1080 4455 1090
rect 4435 990 4455 1000
rect 4525 1080 4545 1090
rect 4525 990 4545 1000
rect 4615 1080 4635 1090
rect 4615 990 4635 1000
rect 4705 1080 4725 1090
rect 4705 990 4725 1000
rect 4795 1080 4815 1090
rect 4795 990 4815 1000
rect 4885 1080 4905 1090
rect 4885 990 4905 1000
rect 4975 1080 4995 1090
rect 4975 990 4995 1000
rect 5065 1080 5085 1090
rect 5065 990 5085 1000
rect 5155 1080 5175 1090
rect 5155 990 5175 1000
rect 5245 1080 5265 1090
rect 5245 990 5265 1000
rect 5335 1080 5355 1090
rect 5335 990 5355 1000
rect 5425 1080 5445 1090
rect 5425 990 5445 1000
rect 5515 1080 5535 1090
rect 5515 990 5535 1000
rect 5605 1080 5625 1090
rect 5605 990 5625 1000
rect 5695 1080 5715 1090
rect 5695 990 5715 1000
rect 5785 1080 5805 1090
rect 5785 990 5805 1000
rect 5875 1080 5895 1090
rect 5875 990 5895 1000
rect 5965 1080 5985 1090
rect 5965 990 5985 1000
rect 6055 1080 6075 1090
rect 6055 990 6075 1000
rect 6145 1080 6165 1090
rect 6145 990 6165 1000
rect 6235 1080 6255 1090
rect 6235 990 6255 1000
rect 6325 1080 6345 1090
rect 6325 990 6345 1000
rect 6415 1080 6435 1090
rect 6415 990 6435 1000
rect 6505 1080 6525 1090
rect 6505 990 6525 1000
rect 6595 1080 6615 1090
rect 6595 990 6615 1000
rect 6685 1080 6705 1090
rect 6685 990 6705 1000
rect 6775 1080 6795 1090
rect 6775 990 6795 1000
rect 6865 1080 6885 1090
rect 6865 990 6885 1000
rect 6955 1080 6975 1090
rect 6955 990 6975 1000
rect 7045 1080 7065 1090
rect 7045 990 7065 1000
rect 7135 1080 7155 1090
rect 7135 990 7155 1000
rect 7225 1080 7245 1090
rect 7225 990 7245 1000
rect 7315 1080 7335 1090
rect 7315 990 7335 1000
rect 7405 1080 7425 1090
rect 7405 990 7425 1000
rect 7495 1080 7515 1090
rect 7495 990 7515 1000
rect 7585 1080 7605 1090
rect 7585 990 7605 1000
rect 7675 1080 7695 1090
rect 7675 990 7695 1000
rect 7765 1080 7785 1090
rect 7765 990 7785 1000
rect 7855 1080 7875 1090
rect 7855 990 7875 1000
rect 7945 1080 7965 1090
rect 7945 990 7965 1000
rect 8035 1080 8055 1090
rect 8035 990 8055 1000
rect 8125 1080 8145 1090
rect 8125 990 8145 1000
rect 8215 1080 8235 1090
rect 8215 990 8235 1000
rect 8305 1080 8325 1090
rect 8305 990 8325 1000
rect 8395 1080 8415 1090
rect 8395 990 8415 1000
rect 8485 1080 8505 1090
rect 8485 990 8505 1000
rect 8575 1080 8595 1090
rect 8575 990 8595 1000
rect 8665 1080 8685 1090
rect 8665 990 8685 1000
rect 8755 1080 8775 1090
rect 8755 990 8775 1000
rect 8845 1080 8865 1090
rect 8845 990 8865 1000
rect 8935 1080 8955 1090
rect 8935 990 8955 1000
rect 9025 1080 9045 1090
rect 9025 990 9045 1000
rect 9115 1080 9135 1090
rect 9115 990 9135 1000
rect 9205 1080 9225 1090
rect 9205 990 9225 1000
rect 9295 1080 9315 1090
rect 9295 990 9315 1000
rect 9385 1080 9405 1090
rect 9385 990 9405 1000
rect 9475 1080 9495 1090
rect 9475 990 9495 1000
rect 9565 1080 9585 1090
rect 9565 990 9585 1000
rect 9655 1080 9675 1090
rect 9655 990 9675 1000
rect 9745 1080 9765 1090
rect 9745 990 9765 1000
rect 9835 1080 9855 1090
rect 9835 990 9855 1000
rect 9925 1080 9945 1090
rect 9925 990 9945 1000
rect 10015 1080 10035 1090
rect 10015 990 10035 1000
rect 10105 1080 10125 1090
rect 10105 990 10125 1000
rect 10195 1080 10215 1090
rect 10195 990 10215 1000
rect 10285 1080 10305 1090
rect 10285 990 10305 1000
rect 10375 1080 10395 1090
rect 10375 990 10395 1000
rect 10465 1080 10485 1090
rect 10465 990 10485 1000
rect 10555 1080 10575 1090
rect 10555 990 10575 1000
rect 10645 1080 10665 1090
rect 10645 990 10665 1000
rect 10735 1080 10755 1090
rect 10735 990 10755 1000
rect 10825 1080 10845 1090
rect 10825 990 10845 1000
rect 10915 1080 10935 1115
rect 10915 990 10935 1000
rect 11005 1080 11025 1090
rect 11005 990 11025 1000
rect 11095 1080 11115 1090
rect 11095 990 11115 1000
rect 11185 1080 11205 1090
rect 11185 990 11205 1000
rect 11245 960 11265 1160
rect -400 940 -340 960
rect -320 940 -295 960
rect -275 940 -205 960
rect -185 940 -115 960
rect -95 940 -25 960
rect -5 940 65 960
rect 85 940 155 960
rect 175 940 200 960
rect 220 940 245 960
rect 265 940 335 960
rect 355 940 380 960
rect 400 940 425 960
rect 445 940 515 960
rect 535 940 560 960
rect 580 940 605 960
rect 625 940 695 960
rect 715 940 740 960
rect 760 940 785 960
rect 805 940 875 960
rect 895 940 920 960
rect 940 940 965 960
rect 985 940 1055 960
rect 1075 940 1100 960
rect 1120 940 1145 960
rect 1165 940 1235 960
rect 1255 940 1280 960
rect 1300 940 1325 960
rect 1345 940 1415 960
rect 1435 940 1460 960
rect 1480 940 1505 960
rect 1525 940 1595 960
rect 1615 940 1640 960
rect 1660 940 1685 960
rect 1705 940 1775 960
rect 1795 940 1820 960
rect 1840 940 1865 960
rect 1885 940 1955 960
rect 1975 940 2000 960
rect 2020 940 2045 960
rect 2065 940 2135 960
rect 2155 940 2180 960
rect 2200 940 2225 960
rect 2245 940 2315 960
rect 2335 940 2360 960
rect 2380 940 2405 960
rect 2425 940 2495 960
rect 2515 940 2540 960
rect 2560 940 2585 960
rect 2605 940 2675 960
rect 2695 940 2720 960
rect 2740 940 2765 960
rect 2785 940 2855 960
rect 2875 940 2900 960
rect 2920 940 2945 960
rect 2965 940 3035 960
rect 3055 940 3085 960
rect 3105 940 3130 960
rect 3150 940 3220 960
rect 3240 940 3265 960
rect 3285 940 3310 960
rect 3330 940 3400 960
rect 3420 940 3445 960
rect 3465 940 3490 960
rect 3510 940 3580 960
rect 3600 940 3625 960
rect 3645 940 3670 960
rect 3690 940 3760 960
rect 3780 940 3805 960
rect 3825 940 3850 960
rect 3870 940 3940 960
rect 3960 940 3985 960
rect 4005 940 4030 960
rect 4050 940 4120 960
rect 4140 940 4165 960
rect 4185 940 4210 960
rect 4230 940 4300 960
rect 4320 940 4345 960
rect 4365 940 4390 960
rect 4410 940 4480 960
rect 4500 940 4525 960
rect 4545 940 4570 960
rect 4590 940 4660 960
rect 4680 940 4705 960
rect 4725 940 4750 960
rect 4770 940 4840 960
rect 4860 940 4885 960
rect 4905 940 4930 960
rect 4950 940 5020 960
rect 5040 940 5065 960
rect 5085 940 5110 960
rect 5130 940 5200 960
rect 5220 940 5245 960
rect 5265 940 5290 960
rect 5310 940 5380 960
rect 5400 940 5425 960
rect 5445 940 5470 960
rect 5490 940 5560 960
rect 5580 940 5605 960
rect 5625 940 5650 960
rect 5670 940 5740 960
rect 5760 940 5785 960
rect 5805 940 5830 960
rect 5850 940 5920 960
rect 5940 940 5965 960
rect 5985 940 6010 960
rect 6030 940 6100 960
rect 6120 940 6145 960
rect 6165 940 6190 960
rect 6210 940 6280 960
rect 6300 940 6325 960
rect 6345 940 6370 960
rect 6390 940 6460 960
rect 6480 940 6505 960
rect 6525 940 6550 960
rect 6570 940 6640 960
rect 6660 940 6685 960
rect 6705 940 6730 960
rect 6750 940 6820 960
rect 6840 940 6865 960
rect 6885 940 6910 960
rect 6930 940 7000 960
rect 7020 940 7045 960
rect 7065 940 7090 960
rect 7110 940 7180 960
rect 7200 940 7225 960
rect 7245 940 7270 960
rect 7290 940 7360 960
rect 7380 940 7405 960
rect 7425 940 7450 960
rect 7470 940 7540 960
rect 7560 940 7585 960
rect 7605 940 7630 960
rect 7650 940 7720 960
rect 7740 940 7765 960
rect 7785 940 7810 960
rect 7830 940 7900 960
rect 7920 940 7945 960
rect 7965 940 7990 960
rect 8010 940 8080 960
rect 8100 940 8125 960
rect 8145 940 8170 960
rect 8190 940 8260 960
rect 8280 940 8305 960
rect 8325 940 8350 960
rect 8370 940 8440 960
rect 8460 940 8485 960
rect 8505 940 8530 960
rect 8550 940 8620 960
rect 8640 940 8665 960
rect 8685 940 8710 960
rect 8730 940 8800 960
rect 8820 940 8845 960
rect 8865 940 8890 960
rect 8910 940 8980 960
rect 9000 940 9025 960
rect 9045 940 9070 960
rect 9090 940 9160 960
rect 9180 940 9205 960
rect 9225 940 9250 960
rect 9270 940 9340 960
rect 9360 940 9385 960
rect 9405 940 9430 960
rect 9450 940 9520 960
rect 9540 940 9565 960
rect 9585 940 9610 960
rect 9630 940 9700 960
rect 9720 940 9745 960
rect 9765 940 9790 960
rect 9810 940 9880 960
rect 9900 940 9925 960
rect 9945 940 9970 960
rect 9990 940 10060 960
rect 10080 940 10105 960
rect 10125 940 10150 960
rect 10170 940 10240 960
rect 10260 940 10285 960
rect 10305 940 10330 960
rect 10350 940 10420 960
rect 10440 940 10465 960
rect 10485 940 10510 960
rect 10530 940 10600 960
rect 10620 940 10645 960
rect 10665 940 10690 960
rect 10710 940 10780 960
rect 10800 940 10870 960
rect 10890 940 10960 960
rect 10980 940 11050 960
rect 11070 940 11140 960
rect 11160 940 11185 960
rect 11205 940 11265 960
rect -400 880 -340 900
rect -320 880 -295 900
rect -275 880 -205 900
rect -185 880 -115 900
rect -95 880 -25 900
rect -5 880 65 900
rect 85 880 155 900
rect 175 880 200 900
rect 220 880 245 900
rect 265 880 335 900
rect 355 880 380 900
rect 400 880 425 900
rect 445 880 515 900
rect 535 880 560 900
rect 580 880 605 900
rect 625 880 695 900
rect 715 880 740 900
rect 760 880 785 900
rect 805 880 875 900
rect 895 880 920 900
rect 940 880 965 900
rect 985 880 1055 900
rect 1075 880 1100 900
rect 1120 880 1145 900
rect 1165 880 1235 900
rect 1255 880 1280 900
rect 1300 880 1325 900
rect 1345 880 1415 900
rect 1435 880 1460 900
rect 1480 880 1505 900
rect 1525 880 1595 900
rect 1615 880 1640 900
rect 1660 880 1685 900
rect 1705 880 1775 900
rect 1795 880 1820 900
rect 1840 880 1865 900
rect 1885 880 1955 900
rect 1975 880 2000 900
rect 2020 880 2045 900
rect 2065 880 2135 900
rect 2155 880 2180 900
rect 2200 880 2225 900
rect 2245 880 2315 900
rect 2335 880 2360 900
rect 2380 880 2405 900
rect 2425 880 2495 900
rect 2515 880 2540 900
rect 2560 880 2585 900
rect 2605 880 2675 900
rect 2695 880 2720 900
rect 2740 880 2765 900
rect 2785 880 2855 900
rect 2875 880 2900 900
rect 2920 880 2945 900
rect 2965 880 3035 900
rect 3055 880 3080 900
rect 3100 880 3125 900
rect 3145 880 3215 900
rect 3235 880 3260 900
rect 3280 880 3305 900
rect 3325 880 3395 900
rect 3415 880 3440 900
rect 3460 880 3485 900
rect 3505 880 3575 900
rect 3595 880 3620 900
rect 3640 880 3665 900
rect 3685 880 3755 900
rect 3775 880 3800 900
rect 3820 880 3845 900
rect 3865 880 3935 900
rect 3955 880 3980 900
rect 4000 880 4025 900
rect 4045 880 4115 900
rect 4135 880 4160 900
rect 4180 880 4205 900
rect 4225 880 4295 900
rect 4315 880 4340 900
rect 4360 880 4385 900
rect 4405 880 4475 900
rect 4495 880 4520 900
rect 4540 880 4565 900
rect 4585 880 4655 900
rect 4675 880 4700 900
rect 4720 880 4745 900
rect 4765 880 4835 900
rect 4855 880 4880 900
rect 4900 880 4925 900
rect 4945 880 5015 900
rect 5035 880 5060 900
rect 5080 880 5105 900
rect 5125 880 5195 900
rect 5215 880 5240 900
rect 5260 880 5285 900
rect 5305 880 5375 900
rect 5395 880 5420 900
rect 5440 880 5465 900
rect 5485 880 5555 900
rect 5575 880 5600 900
rect 5620 880 5645 900
rect 5665 880 5735 900
rect 5755 880 5780 900
rect 5800 880 5825 900
rect 5845 880 5915 900
rect 5935 880 5960 900
rect 5980 880 6005 900
rect 6025 880 6095 900
rect 6115 880 6140 900
rect 6160 880 6185 900
rect 6205 880 6275 900
rect 6295 880 6320 900
rect 6340 880 6365 900
rect 6385 880 6455 900
rect 6475 880 6500 900
rect 6520 880 6545 900
rect 6565 880 6635 900
rect 6655 880 6680 900
rect 6700 880 6725 900
rect 6745 880 6815 900
rect 6835 880 6860 900
rect 6880 880 6905 900
rect 6925 880 6995 900
rect 7015 880 7040 900
rect 7060 880 7085 900
rect 7105 880 7175 900
rect 7195 880 7220 900
rect 7240 880 7265 900
rect 7285 880 7355 900
rect 7375 880 7400 900
rect 7420 880 7445 900
rect 7465 880 7535 900
rect 7555 880 7580 900
rect 7600 880 7625 900
rect 7645 880 7715 900
rect 7735 880 7760 900
rect 7780 880 7810 900
rect 7830 880 7900 900
rect 7920 880 7945 900
rect 7965 880 7990 900
rect 8010 880 8080 900
rect 8100 880 8125 900
rect 8145 880 8170 900
rect 8190 880 8260 900
rect 8280 880 8305 900
rect 8325 880 8350 900
rect 8370 880 8440 900
rect 8460 880 8485 900
rect 8505 880 8530 900
rect 8550 880 8620 900
rect 8640 880 8665 900
rect 8685 880 8710 900
rect 8730 880 8800 900
rect 8820 880 8845 900
rect 8865 880 8890 900
rect 8910 880 8980 900
rect 9000 880 9025 900
rect 9045 880 9070 900
rect 9090 880 9160 900
rect 9180 880 9205 900
rect 9225 880 9250 900
rect 9270 880 9340 900
rect 9360 880 9385 900
rect 9405 880 9430 900
rect 9450 880 9520 900
rect 9540 880 9565 900
rect 9585 880 9610 900
rect 9630 880 9700 900
rect 9720 880 9745 900
rect 9765 880 9790 900
rect 9810 880 9880 900
rect 9900 880 9925 900
rect 9945 880 9970 900
rect 9990 880 10060 900
rect 10080 880 10105 900
rect 10125 880 10150 900
rect 10170 880 10240 900
rect 10260 880 10285 900
rect 10305 880 10330 900
rect 10350 880 10420 900
rect 10440 880 10465 900
rect 10485 880 10510 900
rect 10530 880 10600 900
rect 10620 880 10645 900
rect 10665 880 10690 900
rect 10710 880 10780 900
rect 10800 880 10870 900
rect 10890 880 10960 900
rect 10980 880 11050 900
rect 11070 880 11140 900
rect 11160 880 11185 900
rect 11205 880 11265 900
rect -400 680 -380 880
rect -340 840 -320 850
rect -340 750 -320 760
rect -250 840 -230 850
rect -250 750 -230 760
rect -160 840 -140 850
rect -160 750 -140 760
rect -70 840 -50 850
rect -70 725 -50 760
rect 20 840 40 850
rect 20 750 40 760
rect 110 840 130 850
rect 110 750 130 760
rect 200 840 220 850
rect 200 750 220 760
rect 290 840 310 850
rect 290 750 310 760
rect 380 840 400 850
rect 380 750 400 760
rect 470 840 490 850
rect 470 750 490 760
rect 560 840 580 850
rect 560 750 580 760
rect 650 840 670 850
rect 650 750 670 760
rect 740 840 760 850
rect 740 750 760 760
rect 830 840 850 850
rect 830 750 850 760
rect 920 840 940 850
rect 920 750 940 760
rect 1010 840 1030 850
rect 1010 750 1030 760
rect 1100 840 1120 850
rect 1100 750 1120 760
rect 1190 840 1210 850
rect 1190 750 1210 760
rect 1280 840 1300 850
rect 1280 750 1300 760
rect 1370 840 1390 850
rect 1370 750 1390 760
rect 1460 840 1480 850
rect 1460 750 1480 760
rect 1550 840 1570 850
rect 1550 750 1570 760
rect 1640 840 1660 850
rect 1640 750 1660 760
rect 1730 840 1750 850
rect 1730 750 1750 760
rect 1820 840 1840 850
rect 1820 750 1840 760
rect 1910 840 1930 850
rect 1910 750 1930 760
rect 2000 840 2020 850
rect 2000 750 2020 760
rect 2090 840 2110 850
rect 2090 750 2110 760
rect 2180 840 2200 850
rect 2180 750 2200 760
rect 2270 840 2290 850
rect 2270 750 2290 760
rect 2360 840 2380 850
rect 2360 750 2380 760
rect 2450 840 2470 850
rect 2450 750 2470 760
rect 2540 840 2560 850
rect 2540 750 2560 760
rect 2630 840 2650 850
rect 2630 750 2650 760
rect 2720 840 2740 850
rect 2720 750 2740 760
rect 2810 840 2830 850
rect 2810 750 2830 760
rect 2900 840 2920 850
rect 2900 750 2920 760
rect 2990 840 3010 850
rect 2990 750 3010 760
rect 3080 840 3100 850
rect 3080 750 3100 760
rect 3170 840 3190 850
rect 3170 750 3190 760
rect 3260 840 3280 850
rect 3260 750 3280 760
rect 3350 840 3370 850
rect 3350 750 3370 760
rect 3440 840 3460 850
rect 3440 750 3460 760
rect 3530 840 3550 850
rect 3530 750 3550 760
rect 3620 840 3640 850
rect 3620 750 3640 760
rect 3710 840 3730 850
rect 3710 750 3730 760
rect 3800 840 3820 850
rect 3800 750 3820 760
rect 3890 840 3910 850
rect 3890 750 3910 760
rect 3980 840 4000 850
rect 3980 750 4000 760
rect 4070 840 4090 850
rect 4070 750 4090 760
rect 4160 840 4180 850
rect 4160 750 4180 760
rect 4250 840 4270 850
rect 4250 750 4270 760
rect 4340 840 4360 850
rect 4340 750 4360 760
rect 4430 840 4450 850
rect 4430 750 4450 760
rect 4520 840 4540 850
rect 4520 750 4540 760
rect 4610 840 4630 850
rect 4610 750 4630 760
rect 4700 840 4720 850
rect 4700 750 4720 760
rect 4790 840 4810 850
rect 4790 750 4810 760
rect 4880 840 4900 850
rect 4880 750 4900 760
rect 4970 840 4990 850
rect 4970 750 4990 760
rect 5060 840 5080 850
rect 5060 750 5080 760
rect 5150 840 5170 850
rect 5150 750 5170 760
rect 5240 840 5260 850
rect 5240 750 5260 760
rect 5330 840 5350 850
rect 5330 750 5350 760
rect 5420 840 5440 850
rect 5420 750 5440 760
rect 5510 840 5530 850
rect 5510 750 5530 760
rect 5600 840 5620 850
rect 5600 750 5620 760
rect 5690 840 5710 850
rect 5690 750 5710 760
rect 5780 840 5800 850
rect 5780 750 5800 760
rect 5870 840 5890 850
rect 5870 750 5890 760
rect 5960 840 5980 850
rect 5960 750 5980 760
rect 6050 840 6070 850
rect 6050 750 6070 760
rect 6140 840 6160 850
rect 6140 750 6160 760
rect 6230 840 6250 850
rect 6230 750 6250 760
rect 6320 840 6340 850
rect 6320 750 6340 760
rect 6410 840 6430 850
rect 6410 750 6430 760
rect 6500 840 6520 850
rect 6500 750 6520 760
rect 6590 840 6610 850
rect 6590 750 6610 760
rect 6680 840 6700 850
rect 6680 750 6700 760
rect 6770 840 6790 850
rect 6770 750 6790 760
rect 6860 840 6880 850
rect 6860 750 6880 760
rect 6950 840 6970 850
rect 6950 750 6970 760
rect 7040 840 7060 850
rect 7040 750 7060 760
rect 7130 840 7150 850
rect 7130 750 7150 760
rect 7220 840 7240 850
rect 7220 750 7240 760
rect 7310 840 7330 850
rect 7310 750 7330 760
rect 7400 840 7420 850
rect 7400 750 7420 760
rect 7490 840 7510 850
rect 7490 750 7510 760
rect 7580 840 7600 850
rect 7580 750 7600 760
rect 7670 840 7690 850
rect 7670 750 7690 760
rect 7760 840 7780 850
rect 7760 750 7780 760
rect 7855 840 7875 850
rect 7855 750 7875 760
rect 7945 840 7965 850
rect 7945 750 7965 760
rect 8035 840 8055 850
rect 8035 750 8055 760
rect 8125 840 8145 850
rect 8125 750 8145 760
rect 8215 840 8235 850
rect 8215 750 8235 760
rect 8305 840 8325 850
rect 8305 750 8325 760
rect 8395 840 8415 850
rect 8395 750 8415 760
rect 8485 840 8505 850
rect 8485 750 8505 760
rect 8575 840 8595 850
rect 8575 750 8595 760
rect 8665 840 8685 850
rect 8665 750 8685 760
rect 8755 840 8775 850
rect 8755 750 8775 760
rect 8845 840 8865 850
rect 8845 750 8865 760
rect 8935 840 8955 850
rect 8935 750 8955 760
rect 9025 840 9045 850
rect 9025 750 9045 760
rect 9115 840 9135 850
rect 9115 750 9135 760
rect 9205 840 9225 850
rect 9205 750 9225 760
rect 9295 840 9315 850
rect 9295 750 9315 760
rect 9385 840 9405 850
rect 9385 750 9405 760
rect 9475 840 9495 850
rect 9475 750 9495 760
rect 9565 840 9585 850
rect 9565 750 9585 760
rect 9655 840 9675 850
rect 9655 750 9675 760
rect 9745 840 9765 850
rect 9745 750 9765 760
rect 9835 840 9855 850
rect 9835 750 9855 760
rect 9925 840 9945 850
rect 9925 750 9945 760
rect 10015 840 10035 850
rect 10015 750 10035 760
rect 10105 840 10125 850
rect 10105 750 10125 760
rect 10195 840 10215 850
rect 10195 750 10215 760
rect 10285 840 10305 850
rect 10285 750 10305 760
rect 10375 840 10395 850
rect 10375 750 10395 760
rect 10465 840 10485 850
rect 10465 750 10485 760
rect 10555 840 10575 850
rect 10555 750 10575 760
rect 10645 840 10665 850
rect 10645 750 10665 760
rect 10735 840 10755 850
rect 10735 750 10755 760
rect 10825 840 10845 850
rect 10825 750 10845 760
rect 10915 840 10935 850
rect 10915 725 10935 760
rect 11005 840 11025 850
rect 11005 750 11025 760
rect 11095 840 11115 850
rect 11095 750 11115 760
rect 11185 840 11205 850
rect 11185 750 11205 760
rect -305 705 -295 725
rect -275 705 -205 725
rect -185 705 -115 725
rect -95 705 -25 725
rect -5 705 65 725
rect 85 705 155 725
rect 175 705 190 725
rect 230 705 245 725
rect 265 705 335 725
rect 355 705 365 725
rect 415 705 425 725
rect 445 705 515 725
rect 535 705 545 725
rect 595 705 605 725
rect 625 705 695 725
rect 715 705 725 725
rect 775 705 785 725
rect 805 705 875 725
rect 895 705 905 725
rect 955 705 965 725
rect 985 705 1055 725
rect 1075 705 1085 725
rect 1135 705 1145 725
rect 1165 705 1235 725
rect 1255 705 1265 725
rect 1315 705 1325 725
rect 1345 705 1415 725
rect 1435 705 1445 725
rect 1495 705 1505 725
rect 1525 705 1595 725
rect 1615 705 1625 725
rect 1675 705 1685 725
rect 1705 705 1775 725
rect 1795 705 1805 725
rect 1855 705 1865 725
rect 1885 705 1955 725
rect 1975 705 1985 725
rect 2035 705 2045 725
rect 2065 705 2135 725
rect 2155 705 2165 725
rect 2215 705 2225 725
rect 2245 705 2315 725
rect 2335 705 2345 725
rect 2395 705 2405 725
rect 2425 705 2495 725
rect 2515 705 2525 725
rect 2575 705 2585 725
rect 2605 705 2675 725
rect 2695 705 2705 725
rect 2755 705 2765 725
rect 2785 705 2855 725
rect 2875 705 2885 725
rect 2935 705 2945 725
rect 2965 705 3035 725
rect 3055 705 3065 725
rect 3115 705 3125 725
rect 3145 705 3215 725
rect 3235 705 3245 725
rect 3295 705 3305 725
rect 3325 705 3395 725
rect 3415 705 3425 725
rect 3475 705 3485 725
rect 3505 705 3575 725
rect 3595 705 3605 725
rect 3655 705 3665 725
rect 3685 705 3755 725
rect 3775 705 3785 725
rect 3835 705 3845 725
rect 3865 705 3935 725
rect 3955 705 3965 725
rect 4015 705 4025 725
rect 4045 705 4115 725
rect 4135 705 4145 725
rect 4195 705 4205 725
rect 4225 705 4295 725
rect 4315 705 4325 725
rect 4375 705 4385 725
rect 4405 705 4475 725
rect 4495 705 4505 725
rect 4555 705 4565 725
rect 4585 705 4655 725
rect 4675 705 4685 725
rect 4735 705 4745 725
rect 4765 705 4835 725
rect 4855 705 4865 725
rect 4915 705 4925 725
rect 4945 705 5015 725
rect 5035 705 5045 725
rect 5095 705 5105 725
rect 5125 705 5195 725
rect 5215 705 5225 725
rect 5275 705 5285 725
rect 5305 705 5375 725
rect 5395 705 5405 725
rect 5455 705 5465 725
rect 5485 705 5555 725
rect 5575 705 5585 725
rect 5635 705 5645 725
rect 5665 705 5735 725
rect 5755 705 5765 725
rect 5815 705 5825 725
rect 5845 705 5915 725
rect 5935 705 5945 725
rect 5995 705 6005 725
rect 6025 705 6095 725
rect 6115 705 6125 725
rect 6175 705 6185 725
rect 6205 705 6275 725
rect 6295 705 6305 725
rect 6355 705 6365 725
rect 6385 705 6455 725
rect 6475 705 6485 725
rect 6535 705 6545 725
rect 6565 705 6635 725
rect 6655 705 6665 725
rect 6715 705 6725 725
rect 6745 705 6815 725
rect 6835 705 6845 725
rect 6895 705 6905 725
rect 6925 705 6995 725
rect 7015 705 7025 725
rect 7075 705 7085 725
rect 7105 705 7175 725
rect 7195 705 7205 725
rect 7255 705 7265 725
rect 7285 705 7355 725
rect 7375 705 7385 725
rect 7435 705 7445 725
rect 7465 705 7535 725
rect 7555 705 7565 725
rect 7615 705 7625 725
rect 7645 705 7715 725
rect 7735 705 7745 725
rect 7800 705 7810 725
rect 7830 705 7900 725
rect 7920 705 7930 725
rect 7980 705 7990 725
rect 8010 705 8080 725
rect 8100 705 8110 725
rect 8160 705 8170 725
rect 8190 705 8260 725
rect 8280 705 8290 725
rect 8340 705 8350 725
rect 8370 705 8440 725
rect 8460 705 8470 725
rect 8520 705 8530 725
rect 8550 705 8620 725
rect 8640 705 8650 725
rect 8700 705 8710 725
rect 8730 705 8800 725
rect 8820 705 8830 725
rect 8880 705 8890 725
rect 8910 705 8980 725
rect 9000 705 9010 725
rect 9060 705 9070 725
rect 9090 705 9160 725
rect 9180 705 9190 725
rect 9240 705 9250 725
rect 9270 705 9340 725
rect 9360 705 9370 725
rect 9420 705 9430 725
rect 9450 705 9520 725
rect 9540 705 9550 725
rect 9600 705 9610 725
rect 9630 705 9700 725
rect 9720 705 9730 725
rect 9780 705 9790 725
rect 9810 705 9880 725
rect 9900 705 9910 725
rect 9960 705 9970 725
rect 9990 705 10060 725
rect 10080 705 10090 725
rect 10140 705 10150 725
rect 10170 705 10240 725
rect 10260 705 10270 725
rect 10320 705 10330 725
rect 10350 705 10420 725
rect 10440 705 10450 725
rect 10500 705 10510 725
rect 10530 705 10600 725
rect 10620 705 10630 725
rect 10675 705 10690 725
rect 10710 705 10780 725
rect 10800 705 10870 725
rect 10890 705 10960 725
rect 10980 705 11050 725
rect 11070 705 11140 725
rect 11160 705 11170 725
rect 11245 680 11265 880
rect -400 660 -295 680
rect -275 660 -205 680
rect -185 660 -115 680
rect -95 660 -25 680
rect -5 660 65 680
rect 85 660 155 680
rect 175 660 245 680
rect 265 660 335 680
rect 355 660 425 680
rect 445 660 515 680
rect 535 660 605 680
rect 625 660 695 680
rect 715 660 785 680
rect 805 660 875 680
rect 895 660 965 680
rect 985 660 1055 680
rect 1075 660 1145 680
rect 1165 660 1235 680
rect 1255 660 1325 680
rect 1345 660 1415 680
rect 1435 660 1505 680
rect 1525 660 1595 680
rect 1615 660 1685 680
rect 1705 660 1775 680
rect 1795 660 1865 680
rect 1885 660 1955 680
rect 1975 660 2045 680
rect 2065 660 2135 680
rect 2155 660 2225 680
rect 2245 660 2315 680
rect 2335 660 2405 680
rect 2425 660 2495 680
rect 2515 660 2585 680
rect 2605 660 2675 680
rect 2695 660 2765 680
rect 2785 660 2855 680
rect 2875 660 2945 680
rect 2965 660 3035 680
rect 3055 660 3125 680
rect 3145 660 3215 680
rect 3235 660 3305 680
rect 3325 660 3395 680
rect 3415 660 3485 680
rect 3505 660 3575 680
rect 3595 660 3665 680
rect 3685 660 3755 680
rect 3775 660 3845 680
rect 3865 660 3935 680
rect 3955 660 4025 680
rect 4045 660 4115 680
rect 4135 660 4205 680
rect 4225 660 4295 680
rect 4315 660 4385 680
rect 4405 660 4475 680
rect 4495 660 4565 680
rect 4585 660 4655 680
rect 4675 660 4745 680
rect 4765 660 4835 680
rect 4855 660 4925 680
rect 4945 660 5015 680
rect 5035 660 5105 680
rect 5125 660 5195 680
rect 5215 660 5285 680
rect 5305 660 5375 680
rect 5395 660 5465 680
rect 5485 660 5555 680
rect 5575 660 5645 680
rect 5665 660 5735 680
rect 5755 660 5825 680
rect 5845 660 5915 680
rect 5935 660 6005 680
rect 6025 660 6095 680
rect 6115 660 6185 680
rect 6205 660 6275 680
rect 6295 660 6365 680
rect 6385 660 6455 680
rect 6475 660 6545 680
rect 6565 660 6635 680
rect 6655 660 6725 680
rect 6745 660 6815 680
rect 6835 660 6905 680
rect 6925 660 6995 680
rect 7015 660 7085 680
rect 7105 660 7175 680
rect 7195 660 7265 680
rect 7285 660 7355 680
rect 7375 660 7445 680
rect 7465 660 7535 680
rect 7555 660 7625 680
rect 7645 660 7715 680
rect 7735 660 7810 680
rect 7830 660 7900 680
rect 7920 660 7990 680
rect 8010 660 8080 680
rect 8100 660 8170 680
rect 8190 660 8260 680
rect 8280 660 8350 680
rect 8370 660 8440 680
rect 8460 660 8530 680
rect 8550 660 8620 680
rect 8640 660 8710 680
rect 8730 660 8800 680
rect 8820 660 8890 680
rect 8910 660 8980 680
rect 9000 660 9070 680
rect 9090 660 9160 680
rect 9180 660 9250 680
rect 9270 660 9340 680
rect 9360 660 9430 680
rect 9450 660 9520 680
rect 9540 660 9610 680
rect 9630 660 9700 680
rect 9720 660 9790 680
rect 9810 660 9880 680
rect 9900 660 9970 680
rect 9990 660 10060 680
rect 10080 660 10150 680
rect 10170 660 10240 680
rect 10260 660 10330 680
rect 10350 660 10420 680
rect 10440 660 10510 680
rect 10530 660 10600 680
rect 10620 660 10690 680
rect 10710 660 10780 680
rect 10800 660 10870 680
rect 10890 660 10960 680
rect 10980 660 11050 680
rect 11070 660 11140 680
rect 11160 660 11265 680
rect -350 620 5015 640
rect 5035 620 5195 640
rect 5215 620 5600 640
rect 5620 620 6095 640
rect 6115 620 6275 640
rect 6295 620 6455 640
rect 6475 620 6635 640
rect 6655 620 7535 640
rect 7555 620 7715 640
rect 7735 620 10735 640
rect 10755 620 11215 640
rect 11320 600 11340 1240
rect -475 580 -295 600
rect -275 580 -205 600
rect -185 580 -115 600
rect -95 580 -25 600
rect -5 580 65 600
rect 85 580 155 600
rect 175 580 245 600
rect 265 580 335 600
rect 355 580 425 600
rect 445 580 515 600
rect 535 580 605 600
rect 625 580 695 600
rect 715 580 785 600
rect 805 580 875 600
rect 895 580 965 600
rect 985 580 1055 600
rect 1075 580 1145 600
rect 1165 580 1235 600
rect 1255 580 1325 600
rect 1345 580 1415 600
rect 1435 580 1505 600
rect 1525 580 1595 600
rect 1615 580 1685 600
rect 1705 580 1775 600
rect 1795 580 1865 600
rect 1885 580 1955 600
rect 1975 580 2045 600
rect 2065 580 2135 600
rect 2155 580 2225 600
rect 2245 580 2315 600
rect 2335 580 2405 600
rect 2425 580 2495 600
rect 2515 580 2585 600
rect 2605 580 2675 600
rect 2695 580 2765 600
rect 2785 580 2855 600
rect 2875 580 2945 600
rect 2965 580 3035 600
rect 3055 580 3125 600
rect 3145 580 3215 600
rect 3235 580 3305 600
rect 3325 580 3395 600
rect 3415 580 3485 600
rect 3505 580 3575 600
rect 3595 580 3665 600
rect 3685 580 3755 600
rect 3775 580 3845 600
rect 3865 580 3935 600
rect 3955 580 4025 600
rect 4045 580 4115 600
rect 4135 580 4205 600
rect 4225 580 4295 600
rect 4315 580 4385 600
rect 4405 580 4475 600
rect 4495 580 4565 600
rect 4585 580 4655 600
rect 4675 580 4745 600
rect 4765 580 4835 600
rect 4855 580 4925 600
rect 4945 580 5015 600
rect 5035 580 5105 600
rect 5125 580 5195 600
rect 5215 580 5285 600
rect 5305 580 5375 600
rect 5395 580 5465 600
rect 5485 580 5555 600
rect 5575 580 5645 600
rect 5665 580 5735 600
rect 5755 580 5825 600
rect 5845 580 5915 600
rect 5935 580 6005 600
rect 6025 580 6095 600
rect 6115 580 6185 600
rect 6205 580 6275 600
rect 6295 580 6365 600
rect 6385 580 6455 600
rect 6475 580 6545 600
rect 6565 580 6635 600
rect 6655 580 6725 600
rect 6745 580 6815 600
rect 6835 580 6905 600
rect 6925 580 6995 600
rect 7015 580 7085 600
rect 7105 580 7175 600
rect 7195 580 7265 600
rect 7285 580 7355 600
rect 7375 580 7445 600
rect 7465 580 7535 600
rect 7555 580 7625 600
rect 7645 580 7715 600
rect 7735 580 7810 600
rect 7830 580 7900 600
rect 7920 580 7990 600
rect 8010 580 8080 600
rect 8100 580 8170 600
rect 8190 580 8260 600
rect 8280 580 8350 600
rect 8370 580 8440 600
rect 8460 580 8530 600
rect 8550 580 8620 600
rect 8640 580 8710 600
rect 8730 580 8800 600
rect 8820 580 8890 600
rect 8910 580 8980 600
rect 9000 580 9070 600
rect 9090 580 9160 600
rect 9180 580 9250 600
rect 9270 580 9340 600
rect 9360 580 9430 600
rect 9450 580 9520 600
rect 9540 580 9610 600
rect 9630 580 9700 600
rect 9720 580 9790 600
rect 9810 580 9880 600
rect 9900 580 9970 600
rect 9990 580 10060 600
rect 10080 580 10150 600
rect 10170 580 10240 600
rect 10260 580 10330 600
rect 10350 580 10420 600
rect 10440 580 10510 600
rect 10530 580 10600 600
rect 10620 580 10690 600
rect 10710 580 10780 600
rect 10800 580 10870 600
rect 10890 580 10960 600
rect 10980 580 11050 600
rect 11070 580 11140 600
rect 11160 580 11340 600
rect -350 540 515 560
rect 535 540 1055 560
rect 1075 540 1235 560
rect 1255 540 1775 560
rect 1795 540 1955 560
rect 1975 540 2135 560
rect 2155 540 3035 560
rect 3055 540 3215 560
rect 3235 540 3395 560
rect 3415 540 3575 560
rect 3595 540 4070 560
rect 4090 540 4655 560
rect 4675 540 4835 560
rect 4855 540 7040 560
rect 7060 540 9340 560
rect 9360 540 9520 560
rect 9540 540 10420 560
rect 10440 540 10600 560
rect 10620 540 10825 560
rect 10845 540 11215 560
rect -350 500 695 520
rect 715 500 875 520
rect 895 500 1415 520
rect 1435 500 1595 520
rect 1615 500 2315 520
rect 2335 500 2495 520
rect 2515 500 2675 520
rect 2695 500 2855 520
rect 2875 500 3755 520
rect 3775 500 3935 520
rect 3955 500 4295 520
rect 4315 500 4475 520
rect 4495 500 5375 520
rect 5395 500 5555 520
rect 5575 500 5735 520
rect 5755 500 5915 520
rect 5935 500 6815 520
rect 6835 500 6995 520
rect 7015 500 7175 520
rect 7195 500 7355 520
rect 7375 500 7900 520
rect 7920 500 8080 520
rect 8100 500 8125 520
rect 8145 500 8260 520
rect 8280 500 8440 520
rect 8460 500 8485 520
rect 8505 500 8620 520
rect 8640 500 8800 520
rect 8820 500 8845 520
rect 8865 500 8980 520
rect 9000 500 9160 520
rect 9180 500 9700 520
rect 9720 500 9880 520
rect 9900 500 10060 520
rect 10080 500 10240 520
rect 10260 500 10915 520
rect 10935 500 11215 520
rect -350 460 9925 480
rect 9945 460 11005 480
rect 11025 460 11215 480
rect -350 420 -250 440
rect -230 420 245 440
rect 265 420 3305 440
rect 3325 420 3485 440
rect 3505 420 3665 440
rect 3685 420 3845 440
rect 3865 420 3980 440
rect 4000 420 4115 440
rect 4135 420 4160 440
rect 4180 420 4205 440
rect 4225 420 4385 440
rect 4405 420 4565 440
rect 4585 420 4745 440
rect 4765 420 6365 440
rect 6385 420 6545 440
rect 6565 420 6725 440
rect 6745 420 6905 440
rect 6925 420 7085 440
rect 7105 420 7265 440
rect 7285 420 7445 440
rect 7465 420 7625 440
rect 7645 420 7810 440
rect 7830 420 7990 440
rect 8010 420 8170 440
rect 8190 420 8350 440
rect 8370 420 8530 440
rect 8550 420 8710 440
rect 8730 420 8890 440
rect 8910 420 9070 440
rect 9090 420 11215 440
rect -350 380 -160 400
rect -140 380 425 400
rect 445 380 605 400
rect 625 380 740 400
rect 760 380 785 400
rect 805 380 965 400
rect 985 380 1100 400
rect 1120 380 1145 400
rect 1165 380 1325 400
rect 1345 380 1460 400
rect 1480 380 1505 400
rect 1525 380 1685 400
rect 1705 380 1865 400
rect 1885 380 2045 400
rect 2065 380 2945 400
rect 2965 380 3125 400
rect 3145 380 11215 400
rect -350 340 -70 360
rect -50 340 2225 360
rect 2245 340 2405 360
rect 2425 340 2540 360
rect 2560 340 2585 360
rect 2605 340 2765 360
rect 2785 340 4925 360
rect 4945 340 5105 360
rect 5125 340 5285 360
rect 5305 340 5465 360
rect 5485 340 5645 360
rect 5665 340 5825 360
rect 5845 340 6005 360
rect 6025 340 6185 360
rect 6205 340 11215 360
rect -350 300 20 320
rect 40 300 740 320
rect 760 300 1460 320
rect 1480 300 2180 320
rect 2200 300 2900 320
rect 2920 300 9250 320
rect 9270 300 9430 320
rect 9450 300 9610 320
rect 9630 300 9790 320
rect 9810 300 9970 320
rect 9990 300 10150 320
rect 10170 300 10330 320
rect 10350 300 10510 320
rect 10530 300 11215 320
rect -350 260 110 280
rect 130 260 290 280
rect 310 260 335 280
rect 355 260 4025 280
rect 4045 260 11215 280
rect -475 220 -295 240
rect -275 220 -205 240
rect -185 220 -115 240
rect -95 220 -25 240
rect -5 220 65 240
rect 85 220 155 240
rect 175 220 245 240
rect 265 220 335 240
rect 355 220 425 240
rect 445 220 515 240
rect 535 220 605 240
rect 625 220 695 240
rect 715 220 785 240
rect 805 220 875 240
rect 895 220 965 240
rect 985 220 1055 240
rect 1075 220 1145 240
rect 1165 220 1235 240
rect 1255 220 1325 240
rect 1345 220 1415 240
rect 1435 220 1505 240
rect 1525 220 1595 240
rect 1615 220 1685 240
rect 1705 220 1775 240
rect 1795 220 1865 240
rect 1885 220 1955 240
rect 1975 220 2045 240
rect 2065 220 2135 240
rect 2155 220 2225 240
rect 2245 220 2315 240
rect 2335 220 2405 240
rect 2425 220 2495 240
rect 2515 220 2585 240
rect 2605 220 2675 240
rect 2695 220 2765 240
rect 2785 220 2855 240
rect 2875 220 2945 240
rect 2965 220 3035 240
rect 3055 220 3125 240
rect 3145 220 3215 240
rect 3235 220 3305 240
rect 3325 220 3395 240
rect 3415 220 3485 240
rect 3505 220 3575 240
rect 3595 220 3665 240
rect 3685 220 3755 240
rect 3775 220 3845 240
rect 3865 220 3935 240
rect 3955 220 4025 240
rect 4045 220 4115 240
rect 4135 220 4205 240
rect 4225 220 4295 240
rect 4315 220 4385 240
rect 4405 220 4475 240
rect 4495 220 4565 240
rect 4585 220 4655 240
rect 4675 220 4745 240
rect 4765 220 4835 240
rect 4855 220 4925 240
rect 4945 220 5015 240
rect 5035 220 5105 240
rect 5125 220 5195 240
rect 5215 220 5285 240
rect 5305 220 5375 240
rect 5395 220 5465 240
rect 5485 220 5555 240
rect 5575 220 5645 240
rect 5665 220 5735 240
rect 5755 220 5825 240
rect 5845 220 5915 240
rect 5935 220 6005 240
rect 6025 220 6095 240
rect 6115 220 6185 240
rect 6205 220 6275 240
rect 6295 220 6365 240
rect 6385 220 6455 240
rect 6475 220 6545 240
rect 6565 220 6635 240
rect 6655 220 6725 240
rect 6745 220 6815 240
rect 6835 220 6905 240
rect 6925 220 6995 240
rect 7015 220 7085 240
rect 7105 220 7175 240
rect 7195 220 7265 240
rect 7285 220 7355 240
rect 7375 220 7445 240
rect 7465 220 7535 240
rect 7555 220 7625 240
rect 7645 220 7715 240
rect 7735 220 7810 240
rect 7830 220 7900 240
rect 7920 220 7990 240
rect 8010 220 8080 240
rect 8100 220 8170 240
rect 8190 220 8260 240
rect 8280 220 8350 240
rect 8370 220 8440 240
rect 8460 220 8530 240
rect 8550 220 8620 240
rect 8640 220 8710 240
rect 8730 220 8800 240
rect 8820 220 8890 240
rect 8910 220 8980 240
rect 9000 220 9070 240
rect 9090 220 9160 240
rect 9180 220 9250 240
rect 9270 220 9340 240
rect 9360 220 9430 240
rect 9450 220 9520 240
rect 9540 220 9610 240
rect 9630 220 9700 240
rect 9720 220 9790 240
rect 9810 220 9880 240
rect 9900 220 9970 240
rect 9990 220 10060 240
rect 10080 220 10150 240
rect 10170 220 10240 240
rect 10260 220 10330 240
rect 10350 220 10420 240
rect 10440 220 10510 240
rect 10530 220 10600 240
rect 10620 220 10690 240
rect 10710 220 10780 240
rect 10800 220 10870 240
rect 10890 220 10960 240
rect 10980 220 11050 240
rect 11070 220 11140 240
rect 11160 220 11340 240
rect -475 20 -455 220
rect -305 175 -295 195
rect -275 175 -205 195
rect -185 175 -115 195
rect -95 175 -25 195
rect -5 175 65 195
rect 85 175 155 195
rect 175 175 185 195
rect 235 175 245 195
rect 265 175 335 195
rect 355 175 365 195
rect 415 175 425 195
rect 445 175 515 195
rect 535 175 545 195
rect 595 175 605 195
rect 625 175 695 195
rect 715 175 725 195
rect 775 175 785 195
rect 805 175 875 195
rect 895 175 905 195
rect 955 175 965 195
rect 985 175 1055 195
rect 1075 175 1085 195
rect 1135 175 1145 195
rect 1165 175 1235 195
rect 1255 175 1265 195
rect 1315 175 1325 195
rect 1345 175 1415 195
rect 1435 175 1445 195
rect 1495 175 1505 195
rect 1525 175 1595 195
rect 1615 175 1625 195
rect 1675 175 1685 195
rect 1705 175 1775 195
rect 1795 175 1805 195
rect 1855 175 1865 195
rect 1885 175 1955 195
rect 1975 175 1985 195
rect 2035 175 2045 195
rect 2065 175 2135 195
rect 2155 175 2165 195
rect 2215 175 2225 195
rect 2245 175 2315 195
rect 2335 175 2345 195
rect 2395 175 2405 195
rect 2425 175 2495 195
rect 2515 175 2525 195
rect 2575 175 2585 195
rect 2605 175 2675 195
rect 2695 175 2705 195
rect 2755 175 2765 195
rect 2785 175 2855 195
rect 2875 175 2885 195
rect 2935 175 2945 195
rect 2965 175 3035 195
rect 3055 175 3065 195
rect 3115 175 3125 195
rect 3145 175 3215 195
rect 3235 175 3245 195
rect 3295 175 3305 195
rect 3325 175 3395 195
rect 3415 175 3425 195
rect 3475 175 3485 195
rect 3505 175 3575 195
rect 3595 175 3605 195
rect 3655 175 3665 195
rect 3685 175 3755 195
rect 3775 175 3785 195
rect 3835 175 3845 195
rect 3865 175 3935 195
rect 3955 175 3965 195
rect 4015 175 4025 195
rect 4045 175 4115 195
rect 4135 175 4145 195
rect 4195 175 4205 195
rect 4225 175 4295 195
rect 4315 175 4325 195
rect 4375 175 4385 195
rect 4405 175 4475 195
rect 4495 175 4505 195
rect 4555 175 4565 195
rect 4585 175 4655 195
rect 4675 175 4685 195
rect 4735 175 4745 195
rect 4765 175 4835 195
rect 4855 175 4865 195
rect 4915 175 4925 195
rect 4945 175 5015 195
rect 5035 175 5045 195
rect 5095 175 5105 195
rect 5125 175 5195 195
rect 5215 175 5225 195
rect 5275 175 5285 195
rect 5305 175 5375 195
rect 5395 175 5405 195
rect 5455 175 5465 195
rect 5485 175 5555 195
rect 5575 175 5585 195
rect 5635 175 5645 195
rect 5665 175 5735 195
rect 5755 175 5765 195
rect 5815 175 5825 195
rect 5845 175 5915 195
rect 5935 175 5945 195
rect 5995 175 6005 195
rect 6025 175 6095 195
rect 6115 175 6125 195
rect 6175 175 6185 195
rect 6205 175 6275 195
rect 6295 175 6305 195
rect 6355 175 6365 195
rect 6385 175 6455 195
rect 6475 175 6485 195
rect 6535 175 6545 195
rect 6565 175 6635 195
rect 6655 175 6665 195
rect 6715 175 6725 195
rect 6745 175 6815 195
rect 6835 175 6845 195
rect 6895 175 6905 195
rect 6925 175 6995 195
rect 7015 175 7025 195
rect 7075 175 7085 195
rect 7105 175 7175 195
rect 7195 175 7205 195
rect 7255 175 7265 195
rect 7285 175 7355 195
rect 7375 175 7385 195
rect 7435 175 7445 195
rect 7465 175 7535 195
rect 7555 175 7565 195
rect 7615 175 7625 195
rect 7645 175 7715 195
rect 7735 175 7745 195
rect 7800 175 7810 195
rect 7830 175 7900 195
rect 7920 175 7930 195
rect 7980 175 7990 195
rect 8010 175 8080 195
rect 8100 175 8110 195
rect 8160 175 8170 195
rect 8190 175 8260 195
rect 8280 175 8290 195
rect 8340 175 8350 195
rect 8370 175 8440 195
rect 8460 175 8470 195
rect 8520 175 8530 195
rect 8550 175 8620 195
rect 8640 175 8650 195
rect 8700 175 8710 195
rect 8730 175 8800 195
rect 8820 175 8830 195
rect 8880 175 8890 195
rect 8910 175 8980 195
rect 9000 175 9010 195
rect 9060 175 9070 195
rect 9090 175 9160 195
rect 9180 175 9190 195
rect 9240 175 9250 195
rect 9270 175 9340 195
rect 9360 175 9370 195
rect 9420 175 9430 195
rect 9450 175 9520 195
rect 9540 175 9550 195
rect 9600 175 9610 195
rect 9630 175 9700 195
rect 9720 175 9730 195
rect 9780 175 9790 195
rect 9810 175 9880 195
rect 9900 175 9910 195
rect 9960 175 9970 195
rect 9990 175 10060 195
rect 10080 175 10090 195
rect 10140 175 10150 195
rect 10170 175 10240 195
rect 10260 175 10270 195
rect 10320 175 10330 195
rect 10350 175 10420 195
rect 10440 175 10450 195
rect 10500 175 10510 195
rect 10530 175 10600 195
rect 10620 175 10630 195
rect 10680 175 10690 195
rect 10710 175 10780 195
rect 10800 175 10870 195
rect 10890 175 10960 195
rect 10980 175 11050 195
rect 11070 175 11140 195
rect 11160 175 11170 195
rect -340 140 -320 150
rect -340 50 -320 60
rect -250 140 -230 150
rect -250 50 -230 60
rect -160 140 -140 150
rect -160 50 -140 60
rect -70 140 -50 175
rect -70 50 -50 60
rect 20 140 40 150
rect 20 50 40 60
rect 110 140 130 150
rect 110 50 130 60
rect 200 140 220 150
rect 200 50 220 60
rect 290 140 310 150
rect 290 50 310 60
rect 380 140 400 150
rect 380 50 400 60
rect 470 140 490 150
rect 470 50 490 60
rect 560 140 580 150
rect 560 50 580 60
rect 650 140 670 150
rect 650 50 670 60
rect 740 140 760 150
rect 740 50 760 60
rect 830 140 850 150
rect 830 50 850 60
rect 920 140 940 150
rect 920 50 940 60
rect 1010 140 1030 150
rect 1010 50 1030 60
rect 1100 140 1120 150
rect 1100 50 1120 60
rect 1190 140 1210 150
rect 1190 50 1210 60
rect 1280 140 1300 150
rect 1280 50 1300 60
rect 1370 140 1390 150
rect 1370 50 1390 60
rect 1460 140 1480 150
rect 1460 50 1480 60
rect 1550 140 1570 150
rect 1550 50 1570 60
rect 1640 140 1660 150
rect 1640 50 1660 60
rect 1730 140 1750 150
rect 1730 50 1750 60
rect 1820 140 1840 150
rect 1820 50 1840 60
rect 1910 140 1930 150
rect 1910 50 1930 60
rect 2000 140 2020 150
rect 2000 50 2020 60
rect 2090 140 2110 150
rect 2090 50 2110 60
rect 2180 140 2200 150
rect 2180 50 2200 60
rect 2270 140 2290 150
rect 2270 50 2290 60
rect 2360 140 2380 150
rect 2360 50 2380 60
rect 2450 140 2470 150
rect 2450 50 2470 60
rect 2540 140 2560 150
rect 2540 50 2560 60
rect 2630 140 2650 150
rect 2630 50 2650 60
rect 2720 140 2740 150
rect 2720 50 2740 60
rect 2810 140 2830 150
rect 2810 50 2830 60
rect 2900 140 2920 150
rect 2900 50 2920 60
rect 2990 140 3010 150
rect 2990 50 3010 60
rect 3080 140 3100 150
rect 3080 50 3100 60
rect 3170 140 3190 150
rect 3170 50 3190 60
rect 3260 140 3280 150
rect 3260 50 3280 60
rect 3350 140 3370 150
rect 3350 50 3370 60
rect 3440 140 3460 150
rect 3440 50 3460 60
rect 3530 140 3550 150
rect 3530 50 3550 60
rect 3620 140 3640 150
rect 3620 50 3640 60
rect 3710 140 3730 150
rect 3710 50 3730 60
rect 3800 140 3820 150
rect 3800 50 3820 60
rect 3890 140 3910 150
rect 3890 50 3910 60
rect 3980 140 4000 150
rect 3980 50 4000 60
rect 4070 140 4090 150
rect 4070 50 4090 60
rect 4160 140 4180 150
rect 4160 50 4180 60
rect 4250 140 4270 150
rect 4250 50 4270 60
rect 4340 140 4360 150
rect 4340 50 4360 60
rect 4430 140 4450 150
rect 4430 50 4450 60
rect 4520 140 4540 150
rect 4520 50 4540 60
rect 4610 140 4630 150
rect 4610 50 4630 60
rect 4700 140 4720 150
rect 4700 50 4720 60
rect 4790 140 4810 150
rect 4790 50 4810 60
rect 4880 140 4900 150
rect 4880 50 4900 60
rect 4970 140 4990 150
rect 4970 50 4990 60
rect 5060 140 5080 150
rect 5060 50 5080 60
rect 5150 140 5170 150
rect 5150 50 5170 60
rect 5240 140 5260 150
rect 5240 50 5260 60
rect 5330 140 5350 150
rect 5330 50 5350 60
rect 5420 140 5440 150
rect 5420 50 5440 60
rect 5510 140 5530 150
rect 5510 50 5530 60
rect 5600 140 5620 150
rect 5600 50 5620 60
rect 5690 140 5710 150
rect 5690 50 5710 60
rect 5780 140 5800 150
rect 5780 50 5800 60
rect 5870 140 5890 150
rect 5870 50 5890 60
rect 5960 140 5980 150
rect 5960 50 5980 60
rect 6050 140 6070 150
rect 6050 50 6070 60
rect 6140 140 6160 150
rect 6140 50 6160 60
rect 6230 140 6250 150
rect 6230 50 6250 60
rect 6320 140 6340 150
rect 6320 50 6340 60
rect 6410 140 6430 150
rect 6410 50 6430 60
rect 6500 140 6520 150
rect 6500 50 6520 60
rect 6590 140 6610 150
rect 6590 50 6610 60
rect 6680 140 6700 150
rect 6680 50 6700 60
rect 6770 140 6790 150
rect 6770 50 6790 60
rect 6860 140 6880 150
rect 6860 50 6880 60
rect 6950 140 6970 150
rect 6950 50 6970 60
rect 7040 140 7060 150
rect 7040 50 7060 60
rect 7130 140 7150 150
rect 7130 50 7150 60
rect 7220 140 7240 150
rect 7220 50 7240 60
rect 7310 140 7330 150
rect 7310 50 7330 60
rect 7400 140 7420 150
rect 7400 50 7420 60
rect 7490 140 7510 150
rect 7490 50 7510 60
rect 7580 140 7600 150
rect 7580 50 7600 60
rect 7670 140 7690 150
rect 7670 50 7690 60
rect 7760 140 7780 150
rect 7760 50 7780 60
rect 7855 140 7875 150
rect 7855 50 7875 60
rect 7945 140 7965 150
rect 7945 50 7965 60
rect 8035 140 8055 150
rect 8035 50 8055 60
rect 8125 140 8145 150
rect 8125 50 8145 60
rect 8215 140 8235 150
rect 8215 50 8235 60
rect 8305 140 8325 150
rect 8305 50 8325 60
rect 8395 140 8415 150
rect 8395 50 8415 60
rect 8485 140 8505 150
rect 8485 50 8505 60
rect 8575 140 8595 150
rect 8575 50 8595 60
rect 8665 140 8685 150
rect 8665 50 8685 60
rect 8755 140 8775 150
rect 8755 50 8775 60
rect 8845 140 8865 150
rect 8845 50 8865 60
rect 8935 140 8955 150
rect 8935 50 8955 60
rect 9025 140 9045 150
rect 9025 50 9045 60
rect 9115 140 9135 150
rect 9115 50 9135 60
rect 9205 140 9225 150
rect 9205 50 9225 60
rect 9295 140 9315 150
rect 9295 50 9315 60
rect 9385 140 9405 150
rect 9385 50 9405 60
rect 9475 140 9495 150
rect 9475 50 9495 60
rect 9565 140 9585 150
rect 9565 50 9585 60
rect 9655 140 9675 150
rect 9655 50 9675 60
rect 9745 140 9765 150
rect 9745 50 9765 60
rect 9835 140 9855 150
rect 9835 50 9855 60
rect 9925 140 9945 150
rect 9925 50 9945 60
rect 10015 140 10035 150
rect 10015 50 10035 60
rect 10105 140 10125 150
rect 10105 50 10125 60
rect 10195 140 10215 150
rect 10195 50 10215 60
rect 10285 140 10305 150
rect 10285 50 10305 60
rect 10375 140 10395 150
rect 10375 50 10395 60
rect 10465 140 10485 150
rect 10465 50 10485 60
rect 10555 140 10575 150
rect 10555 50 10575 60
rect 10645 140 10665 150
rect 10645 50 10665 60
rect 10735 140 10755 150
rect 10735 50 10755 60
rect 10825 140 10845 150
rect 10825 50 10845 60
rect 10915 140 10935 175
rect 10915 50 10935 60
rect 11005 140 11025 150
rect 11005 50 11025 60
rect 11095 140 11115 150
rect 11095 50 11115 60
rect 11185 140 11205 150
rect 11185 50 11205 60
rect 11320 20 11340 220
rect -485 0 -475 20
rect -455 0 -340 20
rect -320 0 -295 20
rect -275 0 -205 20
rect -185 0 -115 20
rect -95 0 -25 20
rect -5 0 65 20
rect 85 0 155 20
rect 175 0 200 20
rect 220 0 245 20
rect 265 0 335 20
rect 355 0 380 20
rect 400 0 425 20
rect 445 0 515 20
rect 535 0 560 20
rect 580 0 605 20
rect 625 0 695 20
rect 715 0 740 20
rect 760 0 785 20
rect 805 0 875 20
rect 895 0 920 20
rect 940 0 965 20
rect 985 0 1055 20
rect 1075 0 1100 20
rect 1120 0 1145 20
rect 1165 0 1235 20
rect 1255 0 1280 20
rect 1300 0 1325 20
rect 1345 0 1415 20
rect 1435 0 1460 20
rect 1480 0 1505 20
rect 1525 0 1595 20
rect 1615 0 1640 20
rect 1660 0 1685 20
rect 1705 0 1775 20
rect 1795 0 1820 20
rect 1840 0 1865 20
rect 1885 0 1955 20
rect 1975 0 2000 20
rect 2020 0 2045 20
rect 2065 0 2135 20
rect 2155 0 2180 20
rect 2200 0 2225 20
rect 2245 0 2315 20
rect 2335 0 2360 20
rect 2380 0 2405 20
rect 2425 0 2495 20
rect 2515 0 2540 20
rect 2560 0 2585 20
rect 2605 0 2675 20
rect 2695 0 2720 20
rect 2740 0 2765 20
rect 2785 0 2855 20
rect 2875 0 2900 20
rect 2920 0 2945 20
rect 2965 0 3035 20
rect 3055 0 3080 20
rect 3100 0 3125 20
rect 3145 0 3215 20
rect 3235 0 3260 20
rect 3280 0 3305 20
rect 3325 0 3395 20
rect 3415 0 3440 20
rect 3460 0 3485 20
rect 3505 0 3575 20
rect 3595 0 3620 20
rect 3640 0 3665 20
rect 3685 0 3755 20
rect 3775 0 3800 20
rect 3820 0 3845 20
rect 3865 0 3935 20
rect 3955 0 3980 20
rect 4000 0 4025 20
rect 4045 0 4115 20
rect 4135 0 4160 20
rect 4180 0 4205 20
rect 4225 0 4295 20
rect 4315 0 4340 20
rect 4360 0 4385 20
rect 4405 0 4475 20
rect 4495 0 4520 20
rect 4540 0 4565 20
rect 4585 0 4655 20
rect 4675 0 4700 20
rect 4720 0 4745 20
rect 4765 0 4835 20
rect 4855 0 4880 20
rect 4900 0 4925 20
rect 4945 0 5015 20
rect 5035 0 5060 20
rect 5080 0 5105 20
rect 5125 0 5195 20
rect 5215 0 5240 20
rect 5260 0 5285 20
rect 5305 0 5375 20
rect 5395 0 5420 20
rect 5440 0 5465 20
rect 5485 0 5555 20
rect 5575 0 5600 20
rect 5620 0 5645 20
rect 5665 0 5735 20
rect 5755 0 5780 20
rect 5800 0 5825 20
rect 5845 0 5915 20
rect 5935 0 5960 20
rect 5980 0 6005 20
rect 6025 0 6095 20
rect 6115 0 6140 20
rect 6160 0 6185 20
rect 6205 0 6275 20
rect 6295 0 6320 20
rect 6340 0 6365 20
rect 6385 0 6455 20
rect 6475 0 6500 20
rect 6520 0 6545 20
rect 6565 0 6635 20
rect 6655 0 6680 20
rect 6700 0 6725 20
rect 6745 0 6815 20
rect 6835 0 6860 20
rect 6880 0 6905 20
rect 6925 0 6995 20
rect 7015 0 7040 20
rect 7060 0 7085 20
rect 7105 0 7175 20
rect 7195 0 7220 20
rect 7240 0 7265 20
rect 7285 0 7355 20
rect 7375 0 7400 20
rect 7420 0 7445 20
rect 7465 0 7535 20
rect 7555 0 7580 20
rect 7600 0 7625 20
rect 7645 0 7715 20
rect 7735 0 7760 20
rect 7780 0 7810 20
rect 7830 0 7900 20
rect 7920 0 7945 20
rect 7965 0 7990 20
rect 8010 0 8080 20
rect 8100 0 8125 20
rect 8145 0 8170 20
rect 8190 0 8260 20
rect 8280 0 8305 20
rect 8325 0 8350 20
rect 8370 0 8440 20
rect 8460 0 8485 20
rect 8505 0 8530 20
rect 8550 0 8620 20
rect 8640 0 8665 20
rect 8685 0 8710 20
rect 8730 0 8800 20
rect 8820 0 8845 20
rect 8865 0 8890 20
rect 8910 0 8980 20
rect 9000 0 9025 20
rect 9045 0 9070 20
rect 9090 0 9160 20
rect 9180 0 9205 20
rect 9225 0 9250 20
rect 9270 0 9340 20
rect 9360 0 9385 20
rect 9405 0 9430 20
rect 9450 0 9520 20
rect 9540 0 9565 20
rect 9585 0 9610 20
rect 9630 0 9700 20
rect 9720 0 9745 20
rect 9765 0 9790 20
rect 9810 0 9880 20
rect 9900 0 9925 20
rect 9945 0 9970 20
rect 9990 0 10060 20
rect 10080 0 10105 20
rect 10125 0 10150 20
rect 10170 0 10240 20
rect 10260 0 10285 20
rect 10305 0 10330 20
rect 10350 0 10420 20
rect 10440 0 10465 20
rect 10485 0 10510 20
rect 10530 0 10600 20
rect 10620 0 10645 20
rect 10665 0 10690 20
rect 10710 0 10780 20
rect 10800 0 10870 20
rect 10890 0 10960 20
rect 10980 0 11050 20
rect 11070 0 11140 20
rect 11160 0 11185 20
rect 11205 0 11320 20
rect 11340 0 11350 20
<< viali >>
rect -475 1820 -455 1840
rect -340 1820 -320 1840
rect 200 1820 220 1840
rect 380 1820 400 1840
rect 560 1820 580 1840
rect 740 1820 760 1840
rect 920 1820 940 1840
rect 1100 1820 1120 1840
rect 1280 1820 1300 1840
rect 1460 1820 1480 1840
rect 1640 1820 1660 1840
rect 1820 1820 1840 1840
rect 2000 1820 2020 1840
rect 2180 1820 2200 1840
rect 2360 1820 2380 1840
rect 2540 1820 2560 1840
rect 2720 1820 2740 1840
rect 2900 1820 2920 1840
rect 3085 1820 3105 1840
rect 3265 1820 3285 1840
rect 3445 1820 3465 1840
rect 3625 1820 3645 1840
rect 3805 1820 3825 1840
rect 3985 1820 4005 1840
rect 4165 1820 4185 1840
rect 4345 1820 4365 1840
rect 4525 1820 4545 1840
rect 4705 1820 4725 1840
rect 4885 1820 4905 1840
rect 5065 1820 5085 1840
rect 5245 1820 5265 1840
rect 5425 1820 5445 1840
rect 5605 1820 5625 1840
rect 5785 1820 5805 1840
rect 5965 1820 5985 1840
rect 6145 1820 6165 1840
rect 6325 1820 6345 1840
rect 6505 1820 6525 1840
rect 6685 1820 6705 1840
rect 6865 1820 6885 1840
rect 7045 1820 7065 1840
rect 7225 1820 7245 1840
rect 7405 1820 7425 1840
rect 7585 1820 7605 1840
rect 7765 1820 7785 1840
rect 7945 1820 7965 1840
rect 8125 1820 8145 1840
rect 8305 1820 8325 1840
rect 8485 1820 8505 1840
rect 8665 1820 8685 1840
rect 8845 1820 8865 1840
rect 9025 1820 9045 1840
rect 9205 1820 9225 1840
rect 9385 1820 9405 1840
rect 9565 1820 9585 1840
rect 9745 1820 9765 1840
rect 9925 1820 9945 1840
rect 10105 1820 10125 1840
rect 10285 1820 10305 1840
rect 10465 1820 10485 1840
rect 10645 1820 10665 1840
rect 11185 1820 11205 1840
rect 11320 1820 11340 1840
rect -340 1700 -320 1780
rect 200 1700 220 1780
rect 290 1700 310 1780
rect 380 1700 400 1780
rect 470 1700 490 1780
rect 560 1700 580 1780
rect 650 1700 670 1780
rect 740 1700 760 1780
rect 830 1700 850 1780
rect 920 1700 940 1780
rect 1010 1700 1030 1780
rect 1100 1700 1120 1780
rect 1190 1700 1210 1780
rect 1280 1700 1300 1780
rect 1370 1700 1390 1780
rect 1460 1700 1480 1780
rect 1550 1700 1570 1780
rect 1640 1700 1660 1780
rect 1730 1700 1750 1780
rect 1820 1700 1840 1780
rect 1910 1700 1930 1780
rect 2000 1700 2020 1780
rect 2090 1700 2110 1780
rect 2180 1700 2200 1780
rect 2270 1700 2290 1780
rect 2360 1700 2380 1780
rect 2450 1700 2470 1780
rect 2540 1700 2560 1780
rect 2630 1700 2650 1780
rect 2720 1700 2740 1780
rect 2810 1700 2830 1780
rect 2900 1700 2920 1780
rect 2990 1700 3010 1780
rect 3085 1700 3105 1780
rect 3175 1700 3195 1780
rect 3265 1700 3285 1780
rect 3355 1700 3375 1780
rect 3445 1700 3465 1780
rect 3535 1700 3555 1780
rect 3625 1700 3645 1780
rect 3715 1700 3735 1780
rect 3805 1700 3825 1780
rect 3895 1700 3915 1780
rect 3985 1700 4005 1780
rect 4075 1700 4095 1780
rect 4165 1700 4185 1780
rect 4255 1700 4275 1780
rect 4345 1700 4365 1780
rect 4435 1700 4455 1780
rect 4525 1700 4545 1780
rect 4615 1700 4635 1780
rect 4705 1700 4725 1780
rect 4795 1700 4815 1780
rect 4885 1700 4905 1780
rect 4975 1700 4995 1780
rect 5065 1700 5085 1780
rect 5155 1700 5175 1780
rect 5245 1700 5265 1780
rect 5335 1700 5355 1780
rect 5425 1700 5445 1780
rect 5515 1700 5535 1780
rect 5605 1700 5625 1780
rect 5695 1700 5715 1780
rect 5785 1700 5805 1780
rect 5875 1700 5895 1780
rect 5965 1700 5985 1780
rect 6055 1700 6075 1780
rect 6145 1700 6165 1780
rect 6235 1700 6255 1780
rect 6325 1700 6345 1780
rect 6415 1700 6435 1780
rect 6505 1700 6525 1780
rect 6595 1700 6615 1780
rect 6685 1700 6705 1780
rect 6775 1700 6795 1780
rect 6865 1700 6885 1780
rect 6955 1700 6975 1780
rect 7045 1700 7065 1780
rect 7135 1700 7155 1780
rect 7225 1700 7245 1780
rect 7315 1700 7335 1780
rect 7405 1700 7425 1780
rect 7495 1700 7515 1780
rect 7585 1700 7605 1780
rect 7675 1700 7695 1780
rect 7765 1700 7785 1780
rect 7855 1700 7875 1780
rect 7945 1700 7965 1780
rect 8035 1700 8055 1780
rect 8125 1700 8145 1780
rect 8215 1700 8235 1780
rect 8305 1700 8325 1780
rect 8395 1700 8415 1780
rect 8485 1700 8505 1780
rect 8575 1700 8595 1780
rect 8665 1700 8685 1780
rect 8755 1700 8775 1780
rect 8845 1700 8865 1780
rect 8935 1700 8955 1780
rect 9025 1700 9045 1780
rect 9115 1700 9135 1780
rect 9205 1700 9225 1780
rect 9295 1700 9315 1780
rect 9385 1700 9405 1780
rect 9475 1700 9495 1780
rect 9565 1700 9585 1780
rect 9655 1700 9675 1780
rect 9745 1700 9765 1780
rect 9835 1700 9855 1780
rect 9925 1700 9945 1780
rect 10015 1700 10035 1780
rect 10105 1700 10125 1780
rect 10195 1700 10215 1780
rect 10285 1700 10305 1780
rect 10375 1700 10395 1780
rect 10465 1700 10485 1780
rect 10555 1700 10575 1780
rect 10645 1700 10665 1780
rect 11185 1700 11205 1780
rect 335 1645 355 1665
rect 515 1645 535 1665
rect 695 1645 715 1665
rect 875 1645 895 1665
rect 1055 1645 1075 1665
rect 1235 1645 1255 1665
rect 1415 1645 1435 1665
rect 1595 1645 1615 1665
rect 1775 1645 1795 1665
rect 1955 1645 1975 1665
rect 2135 1645 2155 1665
rect 2315 1645 2335 1665
rect 2495 1645 2515 1665
rect 2675 1645 2695 1665
rect 2855 1645 2875 1665
rect 3035 1645 3055 1665
rect 3220 1645 3240 1665
rect 3400 1645 3420 1665
rect 3580 1645 3600 1665
rect 3760 1645 3780 1665
rect 3940 1645 3960 1665
rect 4120 1645 4140 1665
rect 4300 1645 4320 1665
rect 4480 1645 4500 1665
rect 4660 1645 4680 1665
rect 4840 1645 4860 1665
rect 5020 1645 5040 1665
rect 5200 1645 5220 1665
rect 5380 1645 5400 1665
rect 5560 1645 5580 1665
rect 5740 1645 5760 1665
rect 5920 1645 5940 1665
rect 6100 1645 6120 1665
rect 6280 1645 6300 1665
rect 6460 1645 6480 1665
rect 6640 1645 6660 1665
rect 6820 1645 6840 1665
rect 7000 1645 7020 1665
rect 7180 1645 7200 1665
rect 7360 1645 7380 1665
rect 7540 1645 7560 1665
rect 7720 1645 7740 1665
rect 7900 1645 7920 1665
rect 8080 1645 8100 1665
rect 8260 1645 8280 1665
rect 8440 1645 8460 1665
rect 8620 1645 8640 1665
rect 8800 1645 8820 1665
rect 8980 1645 9000 1665
rect 9160 1645 9180 1665
rect 9340 1645 9360 1665
rect 9520 1645 9540 1665
rect 9700 1645 9720 1665
rect 9880 1645 9900 1665
rect 10060 1645 10080 1665
rect 10240 1645 10260 1665
rect 10420 1645 10440 1665
rect 10600 1645 10620 1665
rect 110 1560 130 1580
rect 6820 1560 6840 1580
rect 10510 1560 10530 1580
rect 10555 1560 10575 1580
rect 20 1520 40 1540
rect 335 1520 355 1540
rect 515 1520 535 1540
rect 695 1520 715 1540
rect 875 1520 895 1540
rect 1055 1520 1075 1540
rect 1235 1520 1255 1540
rect 1415 1520 1435 1540
rect 1595 1520 1615 1540
rect 7945 1520 7965 1540
rect 8665 1520 8685 1540
rect 9385 1520 9405 1540
rect 10105 1520 10125 1540
rect -70 1480 -50 1500
rect 4660 1480 4680 1500
rect 4840 1480 4860 1500
rect 5020 1480 5040 1500
rect 5200 1480 5220 1500
rect 5380 1480 5400 1500
rect 5560 1480 5580 1500
rect 5740 1480 5760 1500
rect 5920 1480 5940 1500
rect 8080 1480 8100 1500
rect 8260 1480 8280 1500
rect 8305 1480 8325 1500
rect 8440 1480 8460 1500
rect 8620 1480 8640 1500
rect -160 1440 -140 1460
rect 7720 1440 7740 1460
rect 7900 1440 7920 1460
rect 8800 1440 8820 1460
rect 8980 1440 9000 1460
rect 9160 1440 9180 1460
rect 9340 1440 9360 1460
rect 9385 1440 9405 1460
rect 9520 1440 9540 1460
rect 9700 1440 9720 1460
rect 9745 1440 9765 1460
rect 9880 1440 9900 1460
rect 10060 1440 10080 1460
rect 10105 1440 10125 1460
rect 10240 1440 10260 1460
rect 10420 1440 10440 1460
rect -250 1400 -230 1420
rect 1775 1400 1795 1420
rect 1955 1400 1975 1420
rect 2135 1400 2155 1420
rect 2315 1400 2335 1420
rect 2495 1400 2515 1420
rect 2675 1400 2695 1420
rect 2855 1400 2875 1420
rect 3035 1400 3055 1420
rect 3220 1400 3240 1420
rect 3400 1400 3420 1420
rect 3580 1400 3600 1420
rect 3760 1400 3780 1420
rect 3940 1400 3960 1420
rect 4120 1400 4140 1420
rect 4300 1400 4320 1420
rect 4480 1400 4500 1420
rect 6100 1400 6120 1420
rect 6280 1400 6300 1420
rect 6460 1400 6480 1420
rect 6640 1400 6660 1420
rect 6685 1400 6705 1420
rect 6730 1400 6750 1420
rect 6865 1400 6885 1420
rect 7000 1400 7020 1420
rect 7180 1400 7200 1420
rect 7360 1400 7380 1420
rect 7540 1400 7560 1420
rect 10600 1400 10620 1420
rect 920 1360 940 1380
rect 11005 1360 11025 1380
rect 605 1320 625 1340
rect 785 1320 805 1340
rect 965 1320 985 1340
rect 1145 1320 1165 1340
rect 1685 1320 1705 1340
rect 1865 1320 1885 1340
rect 2000 1320 2020 1340
rect 2045 1320 2065 1340
rect 2225 1320 2245 1340
rect 2360 1320 2380 1340
rect 2405 1320 2425 1340
rect 2585 1320 2605 1340
rect 2720 1320 2740 1340
rect 2765 1320 2785 1340
rect 2945 1320 2965 1340
rect 3490 1320 3510 1340
rect 3670 1320 3690 1340
rect 3850 1320 3870 1340
rect 4030 1320 4050 1340
rect 4930 1320 4950 1340
rect 5110 1320 5130 1340
rect 5290 1320 5310 1340
rect 5470 1320 5490 1340
rect 6370 1320 6390 1340
rect 6550 1320 6570 1340
rect 6910 1320 6930 1340
rect 7090 1320 7110 1340
rect 7990 1320 8010 1340
rect 8170 1320 8190 1340
rect 8350 1320 8370 1340
rect 8530 1320 8550 1340
rect 9250 1320 9270 1340
rect 9430 1320 9450 1340
rect 9970 1320 9990 1340
rect 10150 1320 10170 1340
rect 10915 1320 10935 1340
rect 245 1280 265 1300
rect 425 1280 445 1300
rect 1325 1280 1345 1300
rect 1505 1280 1525 1300
rect 3805 1280 3825 1300
rect 6010 1280 6030 1300
rect 6190 1280 6210 1300
rect 6775 1280 6795 1300
rect 7270 1280 7290 1300
rect 7450 1280 7470 1300
rect 7630 1280 7650 1300
rect 7810 1280 7830 1300
rect 8710 1280 8730 1300
rect 8890 1280 8910 1300
rect 9070 1280 9090 1300
rect 9610 1280 9630 1300
rect 9790 1280 9810 1300
rect 10330 1280 10350 1300
rect 10825 1280 10845 1300
rect 3130 1200 3150 1220
rect 3310 1200 3330 1220
rect 4210 1200 4230 1220
rect 4390 1200 4410 1220
rect 4570 1200 4590 1220
rect 4750 1200 4770 1220
rect 5245 1200 5265 1220
rect 5650 1200 5670 1220
rect 5830 1200 5850 1220
rect 10735 1200 10755 1220
rect 245 1115 265 1135
rect 425 1115 445 1135
rect 605 1115 625 1135
rect 785 1115 805 1135
rect 965 1115 985 1135
rect 1145 1115 1165 1135
rect 1325 1115 1345 1135
rect 1505 1115 1525 1135
rect 1685 1115 1705 1135
rect 1865 1115 1885 1135
rect 2045 1115 2065 1135
rect 2225 1115 2245 1135
rect 2405 1115 2425 1135
rect 2585 1115 2605 1135
rect 2765 1115 2785 1135
rect 2945 1115 2965 1135
rect 3130 1115 3150 1135
rect 3310 1115 3330 1135
rect 3490 1115 3510 1135
rect 3670 1115 3690 1135
rect 3850 1115 3870 1135
rect 4030 1115 4050 1135
rect 4210 1115 4230 1135
rect 4390 1115 4410 1135
rect 4570 1115 4590 1135
rect 4750 1115 4770 1135
rect 4930 1115 4950 1135
rect 5110 1115 5130 1135
rect 5290 1115 5310 1135
rect 5470 1115 5490 1135
rect 5650 1115 5670 1135
rect 5830 1115 5850 1135
rect 6010 1115 6030 1135
rect 6190 1115 6210 1135
rect 6370 1115 6390 1135
rect 6550 1115 6570 1135
rect 6730 1115 6750 1135
rect 6910 1115 6930 1135
rect 7090 1115 7110 1135
rect 7270 1115 7290 1135
rect 7450 1115 7470 1135
rect 7630 1115 7650 1135
rect 7810 1115 7830 1135
rect 7990 1115 8010 1135
rect 8170 1115 8190 1135
rect 8350 1115 8370 1135
rect 8530 1115 8550 1135
rect 8710 1115 8730 1135
rect 8890 1115 8910 1135
rect 9070 1115 9090 1135
rect 9250 1115 9270 1135
rect 9430 1115 9450 1135
rect 9610 1115 9630 1135
rect 9790 1115 9810 1135
rect 9970 1115 9990 1135
rect 10150 1115 10170 1135
rect 10330 1115 10350 1135
rect 10510 1115 10530 1135
rect -340 1000 -320 1080
rect 200 1000 220 1080
rect 290 1000 310 1080
rect 380 1000 400 1080
rect 470 1000 490 1080
rect 560 1000 580 1080
rect 650 1000 670 1080
rect 740 1000 760 1080
rect 830 1000 850 1080
rect 920 1000 940 1080
rect 1010 1000 1030 1080
rect 1100 1000 1120 1080
rect 1190 1000 1210 1080
rect 1280 1000 1300 1080
rect 1370 1000 1390 1080
rect 1460 1000 1480 1080
rect 1550 1000 1570 1080
rect 1640 1000 1660 1080
rect 1730 1000 1750 1080
rect 1820 1000 1840 1080
rect 1910 1000 1930 1080
rect 2000 1000 2020 1080
rect 2090 1000 2110 1080
rect 2180 1000 2200 1080
rect 2270 1000 2290 1080
rect 2360 1000 2380 1080
rect 2450 1000 2470 1080
rect 2540 1000 2560 1080
rect 2630 1000 2650 1080
rect 2720 1000 2740 1080
rect 2810 1000 2830 1080
rect 2900 1000 2920 1080
rect 2990 1000 3010 1080
rect 3085 1000 3105 1080
rect 3175 1000 3195 1080
rect 3265 1000 3285 1080
rect 3355 1000 3375 1080
rect 3445 1000 3465 1080
rect 3535 1000 3555 1080
rect 3625 1000 3645 1080
rect 3715 1000 3735 1080
rect 3805 1000 3825 1080
rect 3895 1000 3915 1080
rect 3985 1000 4005 1080
rect 4075 1000 4095 1080
rect 4165 1000 4185 1080
rect 4255 1000 4275 1080
rect 4345 1000 4365 1080
rect 4435 1000 4455 1080
rect 4525 1000 4545 1080
rect 4615 1000 4635 1080
rect 4705 1000 4725 1080
rect 4795 1000 4815 1080
rect 4885 1000 4905 1080
rect 4975 1000 4995 1080
rect 5065 1000 5085 1080
rect 5155 1000 5175 1080
rect 5245 1000 5265 1080
rect 5335 1000 5355 1080
rect 5425 1000 5445 1080
rect 5515 1000 5535 1080
rect 5605 1000 5625 1080
rect 5695 1000 5715 1080
rect 5785 1000 5805 1080
rect 5875 1000 5895 1080
rect 5965 1000 5985 1080
rect 6055 1000 6075 1080
rect 6145 1000 6165 1080
rect 6235 1000 6255 1080
rect 6325 1000 6345 1080
rect 6415 1000 6435 1080
rect 6505 1000 6525 1080
rect 6595 1000 6615 1080
rect 6685 1000 6705 1080
rect 6775 1000 6795 1080
rect 6865 1000 6885 1080
rect 6955 1000 6975 1080
rect 7045 1000 7065 1080
rect 7135 1000 7155 1080
rect 7225 1000 7245 1080
rect 7315 1000 7335 1080
rect 7405 1000 7425 1080
rect 7495 1000 7515 1080
rect 7585 1000 7605 1080
rect 7675 1000 7695 1080
rect 7765 1000 7785 1080
rect 7855 1000 7875 1080
rect 7945 1000 7965 1080
rect 8035 1000 8055 1080
rect 8125 1000 8145 1080
rect 8215 1000 8235 1080
rect 8305 1000 8325 1080
rect 8395 1000 8415 1080
rect 8485 1000 8505 1080
rect 8575 1000 8595 1080
rect 8665 1000 8685 1080
rect 8755 1000 8775 1080
rect 8845 1000 8865 1080
rect 8935 1000 8955 1080
rect 9025 1000 9045 1080
rect 9115 1000 9135 1080
rect 9205 1000 9225 1080
rect 9295 1000 9315 1080
rect 9385 1000 9405 1080
rect 9475 1000 9495 1080
rect 9565 1000 9585 1080
rect 9655 1000 9675 1080
rect 9745 1000 9765 1080
rect 9835 1000 9855 1080
rect 9925 1000 9945 1080
rect 10015 1000 10035 1080
rect 10105 1000 10125 1080
rect 10195 1000 10215 1080
rect 10285 1000 10305 1080
rect 10375 1000 10395 1080
rect 10465 1000 10485 1080
rect 10555 1000 10575 1080
rect 10645 1000 10665 1080
rect 11185 1000 11205 1080
rect -340 940 -320 960
rect 200 940 220 960
rect 380 940 400 960
rect 560 940 580 960
rect 740 940 760 960
rect 920 940 940 960
rect 1100 940 1120 960
rect 1280 940 1300 960
rect 1460 940 1480 960
rect 1640 940 1660 960
rect 1820 940 1840 960
rect 2000 940 2020 960
rect 2180 940 2200 960
rect 2360 940 2380 960
rect 2540 940 2560 960
rect 2720 940 2740 960
rect 2900 940 2920 960
rect 3085 940 3105 960
rect 3265 940 3285 960
rect 3445 940 3465 960
rect 3625 940 3645 960
rect 3805 940 3825 960
rect 3985 940 4005 960
rect 4165 940 4185 960
rect 4345 940 4365 960
rect 4525 940 4545 960
rect 4705 940 4725 960
rect 4885 940 4905 960
rect 5065 940 5085 960
rect 5245 940 5265 960
rect 5425 940 5445 960
rect 5605 940 5625 960
rect 5785 940 5805 960
rect 5965 940 5985 960
rect 6145 940 6165 960
rect 6325 940 6345 960
rect 6505 940 6525 960
rect 6685 940 6705 960
rect 6865 940 6885 960
rect 7045 940 7065 960
rect 7225 940 7245 960
rect 7405 940 7425 960
rect 7585 940 7605 960
rect 7765 940 7785 960
rect 7945 940 7965 960
rect 8125 940 8145 960
rect 8305 940 8325 960
rect 8485 940 8505 960
rect 8665 940 8685 960
rect 8845 940 8865 960
rect 9025 940 9045 960
rect 9205 940 9225 960
rect 9385 940 9405 960
rect 9565 940 9585 960
rect 9745 940 9765 960
rect 9925 940 9945 960
rect 10105 940 10125 960
rect 10285 940 10305 960
rect 10465 940 10485 960
rect 10645 940 10665 960
rect 11185 940 11205 960
rect -340 880 -320 900
rect 200 880 220 900
rect 380 880 400 900
rect 560 880 580 900
rect 740 880 760 900
rect 920 880 940 900
rect 1100 880 1120 900
rect 1280 880 1300 900
rect 1460 880 1480 900
rect 1640 880 1660 900
rect 1820 880 1840 900
rect 2000 880 2020 900
rect 2180 880 2200 900
rect 2360 880 2380 900
rect 2540 880 2560 900
rect 2720 880 2740 900
rect 2900 880 2920 900
rect 3080 880 3100 900
rect 3260 880 3280 900
rect 3440 880 3460 900
rect 3620 880 3640 900
rect 3800 880 3820 900
rect 3980 880 4000 900
rect 4160 880 4180 900
rect 4340 880 4360 900
rect 4520 880 4540 900
rect 4700 880 4720 900
rect 4880 880 4900 900
rect 5060 880 5080 900
rect 5240 880 5260 900
rect 5420 880 5440 900
rect 5600 880 5620 900
rect 5780 880 5800 900
rect 5960 880 5980 900
rect 6140 880 6160 900
rect 6320 880 6340 900
rect 6500 880 6520 900
rect 6680 880 6700 900
rect 6860 880 6880 900
rect 7040 880 7060 900
rect 7220 880 7240 900
rect 7400 880 7420 900
rect 7580 880 7600 900
rect 7760 880 7780 900
rect 7945 880 7965 900
rect 8125 880 8145 900
rect 8305 880 8325 900
rect 8485 880 8505 900
rect 8665 880 8685 900
rect 8845 880 8865 900
rect 9025 880 9045 900
rect 9205 880 9225 900
rect 9385 880 9405 900
rect 9565 880 9585 900
rect 9745 880 9765 900
rect 9925 880 9945 900
rect 10105 880 10125 900
rect 10285 880 10305 900
rect 10465 880 10485 900
rect 10645 880 10665 900
rect 11185 880 11205 900
rect -340 760 -320 840
rect 200 760 220 840
rect 290 760 310 840
rect 380 760 400 840
rect 470 760 490 840
rect 560 760 580 840
rect 650 760 670 840
rect 740 760 760 840
rect 830 760 850 840
rect 920 760 940 840
rect 1010 760 1030 840
rect 1100 760 1120 840
rect 1190 760 1210 840
rect 1280 760 1300 840
rect 1370 760 1390 840
rect 1460 760 1480 840
rect 1550 760 1570 840
rect 1640 760 1660 840
rect 1730 760 1750 840
rect 1820 760 1840 840
rect 1910 760 1930 840
rect 2000 760 2020 840
rect 2090 760 2110 840
rect 2180 760 2200 840
rect 2270 760 2290 840
rect 2360 760 2380 840
rect 2450 760 2470 840
rect 2540 760 2560 840
rect 2630 760 2650 840
rect 2720 760 2740 840
rect 2810 760 2830 840
rect 2900 760 2920 840
rect 2990 760 3010 840
rect 3080 760 3100 840
rect 3170 760 3190 840
rect 3260 760 3280 840
rect 3350 760 3370 840
rect 3440 760 3460 840
rect 3530 760 3550 840
rect 3620 760 3640 840
rect 3710 760 3730 840
rect 3800 760 3820 840
rect 3890 760 3910 840
rect 3980 760 4000 840
rect 4070 760 4090 840
rect 4160 760 4180 840
rect 4250 760 4270 840
rect 4340 760 4360 840
rect 4430 760 4450 840
rect 4520 760 4540 840
rect 4610 760 4630 840
rect 4700 760 4720 840
rect 4790 760 4810 840
rect 4880 760 4900 840
rect 4970 760 4990 840
rect 5060 760 5080 840
rect 5150 760 5170 840
rect 5240 760 5260 840
rect 5330 760 5350 840
rect 5420 760 5440 840
rect 5510 760 5530 840
rect 5600 760 5620 840
rect 5690 760 5710 840
rect 5780 760 5800 840
rect 5870 760 5890 840
rect 5960 760 5980 840
rect 6050 760 6070 840
rect 6140 760 6160 840
rect 6230 760 6250 840
rect 6320 760 6340 840
rect 6410 760 6430 840
rect 6500 760 6520 840
rect 6590 760 6610 840
rect 6680 760 6700 840
rect 6770 760 6790 840
rect 6860 760 6880 840
rect 6950 760 6970 840
rect 7040 760 7060 840
rect 7130 760 7150 840
rect 7220 760 7240 840
rect 7310 760 7330 840
rect 7400 760 7420 840
rect 7490 760 7510 840
rect 7580 760 7600 840
rect 7670 760 7690 840
rect 7760 760 7780 840
rect 7855 760 7875 840
rect 7945 760 7965 840
rect 8035 760 8055 840
rect 8125 760 8145 840
rect 8215 760 8235 840
rect 8305 760 8325 840
rect 8395 760 8415 840
rect 8485 760 8505 840
rect 8575 760 8595 840
rect 8665 760 8685 840
rect 8755 760 8775 840
rect 8845 760 8865 840
rect 8935 760 8955 840
rect 9025 760 9045 840
rect 9115 760 9135 840
rect 9205 760 9225 840
rect 9295 760 9315 840
rect 9385 760 9405 840
rect 9475 760 9495 840
rect 9565 760 9585 840
rect 9655 760 9675 840
rect 9745 760 9765 840
rect 9835 760 9855 840
rect 9925 760 9945 840
rect 10015 760 10035 840
rect 10105 760 10125 840
rect 10195 760 10215 840
rect 10285 760 10305 840
rect 10375 760 10395 840
rect 10465 760 10485 840
rect 10555 760 10575 840
rect 10645 760 10665 840
rect 11185 760 11205 840
rect 335 705 355 725
rect 515 705 535 725
rect 695 705 715 725
rect 875 705 895 725
rect 1055 705 1075 725
rect 1235 705 1255 725
rect 1415 705 1435 725
rect 1595 705 1615 725
rect 1775 705 1795 725
rect 1955 705 1975 725
rect 2135 705 2155 725
rect 2315 705 2335 725
rect 2495 705 2515 725
rect 2675 705 2695 725
rect 2855 705 2875 725
rect 3035 705 3055 725
rect 3215 705 3235 725
rect 3395 705 3415 725
rect 3575 705 3595 725
rect 3755 705 3775 725
rect 3935 705 3955 725
rect 4115 705 4135 725
rect 4295 705 4315 725
rect 4475 705 4495 725
rect 4655 705 4675 725
rect 4835 705 4855 725
rect 5015 705 5035 725
rect 5195 705 5215 725
rect 5375 705 5395 725
rect 5555 705 5575 725
rect 5735 705 5755 725
rect 5915 705 5935 725
rect 6095 705 6115 725
rect 6275 705 6295 725
rect 6455 705 6475 725
rect 6635 705 6655 725
rect 6815 705 6835 725
rect 6995 705 7015 725
rect 7175 705 7195 725
rect 7355 705 7375 725
rect 7535 705 7555 725
rect 7715 705 7735 725
rect 7900 705 7920 725
rect 8080 705 8100 725
rect 8260 705 8280 725
rect 8440 705 8460 725
rect 8620 705 8640 725
rect 8800 705 8820 725
rect 8980 705 9000 725
rect 9160 705 9180 725
rect 9340 705 9360 725
rect 9520 705 9540 725
rect 9700 705 9720 725
rect 9880 705 9900 725
rect 10060 705 10080 725
rect 10240 705 10260 725
rect 10420 705 10440 725
rect 10600 705 10620 725
rect 5015 620 5035 640
rect 5195 620 5215 640
rect 5600 620 5620 640
rect 6095 620 6115 640
rect 6275 620 6295 640
rect 6455 620 6475 640
rect 6635 620 6655 640
rect 7535 620 7555 640
rect 7715 620 7735 640
rect 10735 620 10755 640
rect 515 540 535 560
rect 1055 540 1075 560
rect 1235 540 1255 560
rect 1775 540 1795 560
rect 1955 540 1975 560
rect 2135 540 2155 560
rect 3035 540 3055 560
rect 3215 540 3235 560
rect 3395 540 3415 560
rect 3575 540 3595 560
rect 4070 540 4090 560
rect 4655 540 4675 560
rect 4835 540 4855 560
rect 7040 540 7060 560
rect 9340 540 9360 560
rect 9520 540 9540 560
rect 10420 540 10440 560
rect 10600 540 10620 560
rect 10825 540 10845 560
rect 695 500 715 520
rect 875 500 895 520
rect 1415 500 1435 520
rect 1595 500 1615 520
rect 2315 500 2335 520
rect 2495 500 2515 520
rect 2675 500 2695 520
rect 2855 500 2875 520
rect 3755 500 3775 520
rect 3935 500 3955 520
rect 4295 500 4315 520
rect 4475 500 4495 520
rect 5375 500 5395 520
rect 5555 500 5575 520
rect 5735 500 5755 520
rect 5915 500 5935 520
rect 6815 500 6835 520
rect 6995 500 7015 520
rect 7175 500 7195 520
rect 7355 500 7375 520
rect 7900 500 7920 520
rect 8080 500 8100 520
rect 8125 500 8145 520
rect 8260 500 8280 520
rect 8440 500 8460 520
rect 8485 500 8505 520
rect 8620 500 8640 520
rect 8800 500 8820 520
rect 8845 500 8865 520
rect 8980 500 9000 520
rect 9160 500 9180 520
rect 9700 500 9720 520
rect 9880 500 9900 520
rect 10060 500 10080 520
rect 10240 500 10260 520
rect 10915 500 10935 520
rect 9925 460 9945 480
rect 11005 460 11025 480
rect -250 420 -230 440
rect 245 420 265 440
rect 3305 420 3325 440
rect 3485 420 3505 440
rect 3665 420 3685 440
rect 3845 420 3865 440
rect 3980 420 4000 440
rect 4115 420 4135 440
rect 4160 420 4180 440
rect 4205 420 4225 440
rect 4385 420 4405 440
rect 4565 420 4585 440
rect 4745 420 4765 440
rect 6365 420 6385 440
rect 6545 420 6565 440
rect 6725 420 6745 440
rect 6905 420 6925 440
rect 7085 420 7105 440
rect 7265 420 7285 440
rect 7445 420 7465 440
rect 7625 420 7645 440
rect 7810 420 7830 440
rect 7990 420 8010 440
rect 8170 420 8190 440
rect 8350 420 8370 440
rect 8530 420 8550 440
rect 8710 420 8730 440
rect 8890 420 8910 440
rect 9070 420 9090 440
rect -160 380 -140 400
rect 425 380 445 400
rect 605 380 625 400
rect 740 380 760 400
rect 785 380 805 400
rect 965 380 985 400
rect 1100 380 1120 400
rect 1145 380 1165 400
rect 1325 380 1345 400
rect 1460 380 1480 400
rect 1505 380 1525 400
rect 1685 380 1705 400
rect 1865 380 1885 400
rect 2045 380 2065 400
rect 2945 380 2965 400
rect 3125 380 3145 400
rect -70 340 -50 360
rect 2225 340 2245 360
rect 2405 340 2425 360
rect 2540 340 2560 360
rect 2585 340 2605 360
rect 2765 340 2785 360
rect 4925 340 4945 360
rect 5105 340 5125 360
rect 5285 340 5305 360
rect 5465 340 5485 360
rect 5645 340 5665 360
rect 5825 340 5845 360
rect 6005 340 6025 360
rect 6185 340 6205 360
rect 20 300 40 320
rect 740 300 760 320
rect 1460 300 1480 320
rect 2180 300 2200 320
rect 2900 300 2920 320
rect 9250 300 9270 320
rect 9430 300 9450 320
rect 9610 300 9630 320
rect 9790 300 9810 320
rect 9970 300 9990 320
rect 10150 300 10170 320
rect 10330 300 10350 320
rect 10510 300 10530 320
rect 110 260 130 280
rect 290 260 310 280
rect 335 260 355 280
rect 4025 260 4045 280
rect 245 175 265 195
rect 425 175 445 195
rect 605 175 625 195
rect 785 175 805 195
rect 965 175 985 195
rect 1145 175 1165 195
rect 1325 175 1345 195
rect 1505 175 1525 195
rect 1685 175 1705 195
rect 1865 175 1885 195
rect 2045 175 2065 195
rect 2225 175 2245 195
rect 2405 175 2425 195
rect 2585 175 2605 195
rect 2765 175 2785 195
rect 2945 175 2965 195
rect 3125 175 3145 195
rect 3305 175 3325 195
rect 3485 175 3505 195
rect 3665 175 3685 195
rect 3845 175 3865 195
rect 4025 175 4045 195
rect 4205 175 4225 195
rect 4385 175 4405 195
rect 4565 175 4585 195
rect 4745 175 4765 195
rect 4925 175 4945 195
rect 5105 175 5125 195
rect 5285 175 5305 195
rect 5465 175 5485 195
rect 5645 175 5665 195
rect 5825 175 5845 195
rect 6005 175 6025 195
rect 6185 175 6205 195
rect 6365 175 6385 195
rect 6545 175 6565 195
rect 6725 175 6745 195
rect 6905 175 6925 195
rect 7085 175 7105 195
rect 7265 175 7285 195
rect 7445 175 7465 195
rect 7625 175 7645 195
rect 7810 175 7830 195
rect 7990 175 8010 195
rect 8170 175 8190 195
rect 8350 175 8370 195
rect 8530 175 8550 195
rect 8710 175 8730 195
rect 8890 175 8910 195
rect 9070 175 9090 195
rect 9250 175 9270 195
rect 9430 175 9450 195
rect 9610 175 9630 195
rect 9790 175 9810 195
rect 9970 175 9990 195
rect 10150 175 10170 195
rect 10330 175 10350 195
rect 10510 175 10530 195
rect -340 60 -320 140
rect 200 60 220 140
rect 290 60 310 140
rect 380 60 400 140
rect 470 60 490 140
rect 560 60 580 140
rect 650 60 670 140
rect 740 60 760 140
rect 830 60 850 140
rect 920 60 940 140
rect 1010 60 1030 140
rect 1100 60 1120 140
rect 1190 60 1210 140
rect 1280 60 1300 140
rect 1370 60 1390 140
rect 1460 60 1480 140
rect 1550 60 1570 140
rect 1640 60 1660 140
rect 1730 60 1750 140
rect 1820 60 1840 140
rect 1910 60 1930 140
rect 2000 60 2020 140
rect 2090 60 2110 140
rect 2180 60 2200 140
rect 2270 60 2290 140
rect 2360 60 2380 140
rect 2450 60 2470 140
rect 2540 60 2560 140
rect 2630 60 2650 140
rect 2720 60 2740 140
rect 2810 60 2830 140
rect 2900 60 2920 140
rect 2990 60 3010 140
rect 3080 60 3100 140
rect 3170 60 3190 140
rect 3260 60 3280 140
rect 3350 60 3370 140
rect 3440 60 3460 140
rect 3530 60 3550 140
rect 3620 60 3640 140
rect 3710 60 3730 140
rect 3800 60 3820 140
rect 3890 60 3910 140
rect 3980 60 4000 140
rect 4070 60 4090 140
rect 4160 60 4180 140
rect 4250 60 4270 140
rect 4340 60 4360 140
rect 4430 60 4450 140
rect 4520 60 4540 140
rect 4610 60 4630 140
rect 4700 60 4720 140
rect 4790 60 4810 140
rect 4880 60 4900 140
rect 4970 60 4990 140
rect 5060 60 5080 140
rect 5150 60 5170 140
rect 5240 60 5260 140
rect 5330 60 5350 140
rect 5420 60 5440 140
rect 5510 60 5530 140
rect 5600 60 5620 140
rect 5690 60 5710 140
rect 5780 60 5800 140
rect 5870 60 5890 140
rect 5960 60 5980 140
rect 6050 60 6070 140
rect 6140 60 6160 140
rect 6230 60 6250 140
rect 6320 60 6340 140
rect 6410 60 6430 140
rect 6500 60 6520 140
rect 6590 60 6610 140
rect 6680 60 6700 140
rect 6770 60 6790 140
rect 6860 60 6880 140
rect 6950 60 6970 140
rect 7040 60 7060 140
rect 7130 60 7150 140
rect 7220 60 7240 140
rect 7310 60 7330 140
rect 7400 60 7420 140
rect 7490 60 7510 140
rect 7580 60 7600 140
rect 7670 60 7690 140
rect 7760 60 7780 140
rect 7855 60 7875 140
rect 7945 60 7965 140
rect 8035 60 8055 140
rect 8125 60 8145 140
rect 8215 60 8235 140
rect 8305 60 8325 140
rect 8395 60 8415 140
rect 8485 60 8505 140
rect 8575 60 8595 140
rect 8665 60 8685 140
rect 8755 60 8775 140
rect 8845 60 8865 140
rect 8935 60 8955 140
rect 9025 60 9045 140
rect 9115 60 9135 140
rect 9205 60 9225 140
rect 9295 60 9315 140
rect 9385 60 9405 140
rect 9475 60 9495 140
rect 9565 60 9585 140
rect 9655 60 9675 140
rect 9745 60 9765 140
rect 9835 60 9855 140
rect 9925 60 9945 140
rect 10015 60 10035 140
rect 10105 60 10125 140
rect 10195 60 10215 140
rect 10285 60 10305 140
rect 10375 60 10395 140
rect 10465 60 10485 140
rect 10555 60 10575 140
rect 10645 60 10665 140
rect 11185 60 11205 140
rect -475 0 -455 20
rect -340 0 -320 20
rect 200 0 220 20
rect 380 0 400 20
rect 560 0 580 20
rect 740 0 760 20
rect 920 0 940 20
rect 1100 0 1120 20
rect 1280 0 1300 20
rect 1460 0 1480 20
rect 1640 0 1660 20
rect 1820 0 1840 20
rect 2000 0 2020 20
rect 2180 0 2200 20
rect 2360 0 2380 20
rect 2540 0 2560 20
rect 2720 0 2740 20
rect 2900 0 2920 20
rect 3080 0 3100 20
rect 3260 0 3280 20
rect 3440 0 3460 20
rect 3620 0 3640 20
rect 3800 0 3820 20
rect 3980 0 4000 20
rect 4160 0 4180 20
rect 4340 0 4360 20
rect 4520 0 4540 20
rect 4700 0 4720 20
rect 4880 0 4900 20
rect 5060 0 5080 20
rect 5240 0 5260 20
rect 5420 0 5440 20
rect 5600 0 5620 20
rect 5780 0 5800 20
rect 5960 0 5980 20
rect 6140 0 6160 20
rect 6320 0 6340 20
rect 6500 0 6520 20
rect 6680 0 6700 20
rect 6860 0 6880 20
rect 7040 0 7060 20
rect 7220 0 7240 20
rect 7400 0 7420 20
rect 7580 0 7600 20
rect 7760 0 7780 20
rect 7945 0 7965 20
rect 8125 0 8145 20
rect 8305 0 8325 20
rect 8485 0 8505 20
rect 8665 0 8685 20
rect 8845 0 8865 20
rect 9025 0 9045 20
rect 9205 0 9225 20
rect 9385 0 9405 20
rect 9565 0 9585 20
rect 9745 0 9765 20
rect 9925 0 9945 20
rect 10105 0 10125 20
rect 10285 0 10305 20
rect 10465 0 10485 20
rect 10645 0 10665 20
rect 11185 0 11205 20
rect 11320 0 11340 20
<< metal1 >>
rect -485 1845 -445 1850
rect -485 1815 -480 1845
rect -450 1815 -445 1845
rect -485 25 -445 1815
rect -350 1845 -315 1850
rect -350 1815 -345 1845
rect 190 1845 230 1850
rect -315 1815 -310 1840
rect -350 1810 -310 1815
rect 190 1815 195 1845
rect 225 1815 230 1845
rect 190 1810 230 1815
rect 370 1845 410 1850
rect 370 1815 375 1845
rect 405 1815 410 1845
rect 370 1810 410 1815
rect 550 1845 590 1850
rect 550 1815 555 1845
rect 585 1815 590 1845
rect 550 1810 590 1815
rect 730 1845 770 1850
rect 730 1815 735 1845
rect 765 1815 770 1845
rect 730 1810 770 1815
rect 910 1845 950 1850
rect 910 1815 915 1845
rect 945 1815 950 1845
rect 910 1810 950 1815
rect 1090 1845 1130 1850
rect 1090 1815 1095 1845
rect 1125 1815 1130 1845
rect 1090 1810 1130 1815
rect 1270 1845 1310 1850
rect 1270 1815 1275 1845
rect 1305 1815 1310 1845
rect 1270 1810 1310 1815
rect 1450 1845 1490 1850
rect 1450 1815 1455 1845
rect 1485 1815 1490 1845
rect 1450 1810 1490 1815
rect 1630 1845 1670 1850
rect 1630 1815 1635 1845
rect 1665 1815 1670 1845
rect 1630 1810 1670 1815
rect 1810 1845 1850 1850
rect 1810 1815 1815 1845
rect 1845 1815 1850 1845
rect 1810 1810 1850 1815
rect 1990 1845 2030 1850
rect 1990 1815 1995 1845
rect 2025 1815 2030 1845
rect 1990 1810 2030 1815
rect 2170 1845 2210 1850
rect 2170 1815 2175 1845
rect 2205 1815 2210 1845
rect 2170 1810 2210 1815
rect 2350 1845 2390 1850
rect 2350 1815 2355 1845
rect 2385 1815 2390 1845
rect 2350 1810 2390 1815
rect 2530 1845 2570 1850
rect 2530 1815 2535 1845
rect 2565 1815 2570 1845
rect 2530 1810 2570 1815
rect 2710 1845 2750 1850
rect 2710 1815 2715 1845
rect 2745 1815 2750 1845
rect 2710 1810 2750 1815
rect 2890 1845 2930 1850
rect 2890 1815 2895 1845
rect 2925 1815 2930 1845
rect 2890 1810 2930 1815
rect 3070 1845 3115 1850
rect 3070 1815 3080 1845
rect 3110 1815 3115 1845
rect 3070 1810 3115 1815
rect 3255 1845 3295 1850
rect 3255 1815 3260 1845
rect 3290 1815 3295 1845
rect 3255 1810 3295 1815
rect 3435 1845 3475 1850
rect 3435 1815 3440 1845
rect 3470 1815 3475 1845
rect 3435 1810 3475 1815
rect 3615 1845 3655 1850
rect 3615 1815 3620 1845
rect 3650 1815 3655 1845
rect 3615 1810 3655 1815
rect 3795 1845 3835 1850
rect 3795 1815 3800 1845
rect 3830 1815 3835 1845
rect 3795 1810 3835 1815
rect 3975 1845 4015 1850
rect 3975 1815 3980 1845
rect 4010 1815 4015 1845
rect 3975 1810 4015 1815
rect 4155 1845 4195 1850
rect 4155 1815 4160 1845
rect 4190 1815 4195 1845
rect 4155 1810 4195 1815
rect 4335 1845 4375 1850
rect 4335 1815 4340 1845
rect 4370 1815 4375 1845
rect 4335 1810 4375 1815
rect 4515 1845 4555 1850
rect 4515 1815 4520 1845
rect 4550 1815 4555 1845
rect 4515 1810 4555 1815
rect 4695 1845 4735 1850
rect 4695 1815 4700 1845
rect 4730 1815 4735 1845
rect 4695 1810 4735 1815
rect 4875 1845 4915 1850
rect 4875 1815 4880 1845
rect 4910 1815 4915 1845
rect 4875 1810 4915 1815
rect 5055 1845 5095 1850
rect 5055 1815 5060 1845
rect 5090 1815 5095 1845
rect 5055 1810 5095 1815
rect 5235 1845 5275 1850
rect 5235 1815 5240 1845
rect 5270 1815 5275 1845
rect 5235 1810 5275 1815
rect 5415 1845 5455 1850
rect 5415 1815 5420 1845
rect 5450 1815 5455 1845
rect 5415 1810 5455 1815
rect 5595 1845 5635 1850
rect 5595 1815 5600 1845
rect 5630 1815 5635 1845
rect 5595 1810 5635 1815
rect 5775 1845 5815 1850
rect 5775 1815 5780 1845
rect 5810 1815 5815 1845
rect 5775 1810 5815 1815
rect 5955 1845 5995 1850
rect 5955 1815 5960 1845
rect 5990 1815 5995 1845
rect 5955 1810 5995 1815
rect 6135 1845 6175 1850
rect 6135 1815 6140 1845
rect 6170 1815 6175 1845
rect 6135 1810 6175 1815
rect 6315 1845 6355 1850
rect 6315 1815 6320 1845
rect 6350 1815 6355 1845
rect 6315 1810 6355 1815
rect 6495 1845 6535 1850
rect 6495 1815 6500 1845
rect 6530 1815 6535 1845
rect 6495 1810 6535 1815
rect 6675 1845 6715 1850
rect 6675 1815 6680 1845
rect 6710 1815 6715 1845
rect 6675 1810 6715 1815
rect 6855 1845 6895 1850
rect 6855 1815 6860 1845
rect 6890 1815 6895 1845
rect 6855 1810 6895 1815
rect 7035 1845 7075 1850
rect 7035 1815 7040 1845
rect 7070 1815 7075 1845
rect 7035 1810 7075 1815
rect 7215 1845 7255 1850
rect 7215 1815 7220 1845
rect 7250 1815 7255 1845
rect 7215 1810 7255 1815
rect 7395 1845 7435 1850
rect 7395 1815 7400 1845
rect 7430 1815 7435 1845
rect 7395 1810 7435 1815
rect 7575 1845 7615 1850
rect 7575 1815 7580 1845
rect 7610 1815 7615 1845
rect 7575 1810 7615 1815
rect 7755 1845 7795 1850
rect 7755 1815 7760 1845
rect 7790 1815 7795 1845
rect 7755 1810 7795 1815
rect 7935 1845 7975 1850
rect 7935 1815 7940 1845
rect 7970 1815 7975 1845
rect 7935 1810 7975 1815
rect 8115 1845 8155 1850
rect 8115 1815 8120 1845
rect 8150 1815 8155 1845
rect 8115 1810 8155 1815
rect 8295 1845 8335 1850
rect 8295 1815 8300 1845
rect 8330 1815 8335 1845
rect 8295 1810 8335 1815
rect 8475 1845 8515 1850
rect 8475 1815 8480 1845
rect 8510 1815 8515 1845
rect 8475 1810 8515 1815
rect 8655 1845 8695 1850
rect 8655 1815 8660 1845
rect 8690 1815 8695 1845
rect 8655 1810 8695 1815
rect 8835 1845 8875 1850
rect 8835 1815 8840 1845
rect 8870 1815 8875 1845
rect 8835 1810 8875 1815
rect 9015 1845 9055 1850
rect 9015 1815 9020 1845
rect 9050 1815 9055 1845
rect 9015 1810 9055 1815
rect 9195 1845 9235 1850
rect 9195 1815 9200 1845
rect 9230 1815 9235 1845
rect 9195 1810 9235 1815
rect 9375 1845 9415 1850
rect 9375 1815 9380 1845
rect 9410 1815 9415 1845
rect 9375 1810 9415 1815
rect 9555 1845 9595 1850
rect 9555 1815 9560 1845
rect 9590 1815 9595 1845
rect 9555 1810 9595 1815
rect 9735 1845 9775 1850
rect 9735 1815 9740 1845
rect 9770 1815 9775 1845
rect 9735 1810 9775 1815
rect 9915 1845 9955 1850
rect 9915 1815 9920 1845
rect 9950 1815 9955 1845
rect 9915 1810 9955 1815
rect 10095 1845 10135 1850
rect 10095 1815 10100 1845
rect 10130 1815 10135 1845
rect 10095 1810 10135 1815
rect 10275 1845 10315 1850
rect 10275 1815 10280 1845
rect 10310 1815 10315 1845
rect 10275 1810 10315 1815
rect 10455 1845 10495 1850
rect 10455 1815 10460 1845
rect 10490 1815 10495 1845
rect 10640 1845 10675 1850
rect 10455 1810 10495 1815
rect 10635 1815 10640 1840
rect 10670 1815 10675 1845
rect 11180 1845 11350 1850
rect 10635 1810 10675 1815
rect 11175 1815 11180 1840
rect 11210 1815 11315 1845
rect 11345 1815 11350 1845
rect 11175 1810 11350 1815
rect -340 1790 -320 1810
rect 200 1790 220 1810
rect 920 1790 940 1810
rect 1640 1790 1660 1810
rect 3085 1790 3105 1810
rect 4525 1790 4545 1810
rect 5965 1790 5985 1810
rect 6145 1790 6165 1810
rect 7585 1790 7605 1810
rect 9025 1790 9045 1810
rect 10465 1790 10485 1810
rect 10645 1790 10665 1810
rect 11185 1790 11205 1810
rect -345 1780 -315 1790
rect -345 1700 -340 1780
rect -320 1700 -315 1780
rect -345 1690 -315 1700
rect -255 1690 -225 1790
rect -165 1690 -135 1790
rect -75 1690 -45 1790
rect 15 1690 45 1790
rect 105 1690 135 1790
rect 195 1780 225 1790
rect 195 1700 200 1780
rect 220 1700 225 1780
rect 195 1690 225 1700
rect 285 1780 315 1790
rect 285 1700 290 1780
rect 310 1700 315 1780
rect 285 1690 315 1700
rect 375 1780 405 1790
rect 375 1700 380 1780
rect 400 1700 405 1780
rect 375 1690 405 1700
rect 465 1780 495 1790
rect 465 1700 470 1780
rect 490 1700 495 1780
rect 465 1690 495 1700
rect 555 1780 585 1790
rect 555 1700 560 1780
rect 580 1700 585 1780
rect 555 1690 585 1700
rect 645 1780 675 1790
rect 645 1700 650 1780
rect 670 1700 675 1780
rect 645 1690 675 1700
rect 735 1780 765 1790
rect 735 1700 740 1780
rect 760 1700 765 1780
rect 735 1690 765 1700
rect 825 1780 855 1790
rect 825 1700 830 1780
rect 850 1700 855 1780
rect 825 1690 855 1700
rect 915 1780 945 1790
rect 915 1700 920 1780
rect 940 1700 945 1780
rect 915 1690 945 1700
rect 1005 1780 1035 1790
rect 1005 1700 1010 1780
rect 1030 1700 1035 1780
rect 1005 1690 1035 1700
rect 1095 1780 1125 1790
rect 1095 1700 1100 1780
rect 1120 1700 1125 1780
rect 1095 1690 1125 1700
rect 1185 1780 1215 1790
rect 1185 1700 1190 1780
rect 1210 1700 1215 1780
rect 1185 1690 1215 1700
rect 1275 1780 1305 1790
rect 1275 1700 1280 1780
rect 1300 1700 1305 1780
rect 1275 1690 1305 1700
rect 1365 1780 1395 1790
rect 1365 1700 1370 1780
rect 1390 1700 1395 1780
rect 1365 1690 1395 1700
rect 1455 1780 1485 1790
rect 1455 1700 1460 1780
rect 1480 1700 1485 1780
rect 1455 1690 1485 1700
rect 1545 1780 1575 1790
rect 1545 1700 1550 1780
rect 1570 1700 1575 1780
rect 1545 1690 1575 1700
rect 1635 1780 1665 1790
rect 1635 1700 1640 1780
rect 1660 1700 1665 1780
rect 1635 1690 1665 1700
rect 1725 1780 1755 1790
rect 1725 1700 1730 1780
rect 1750 1700 1755 1780
rect 1725 1690 1755 1700
rect 1815 1780 1845 1790
rect 1815 1700 1820 1780
rect 1840 1700 1845 1780
rect 1815 1690 1845 1700
rect 1905 1780 1935 1790
rect 1905 1700 1910 1780
rect 1930 1700 1935 1780
rect 1905 1690 1935 1700
rect 1995 1780 2025 1790
rect 1995 1700 2000 1780
rect 2020 1700 2025 1780
rect 1995 1690 2025 1700
rect 2085 1780 2115 1790
rect 2085 1700 2090 1780
rect 2110 1700 2115 1780
rect 2085 1690 2115 1700
rect 2175 1780 2205 1790
rect 2175 1700 2180 1780
rect 2200 1700 2205 1780
rect 2175 1690 2205 1700
rect 2265 1780 2295 1790
rect 2265 1700 2270 1780
rect 2290 1700 2295 1780
rect 2265 1690 2295 1700
rect 2355 1780 2385 1790
rect 2355 1700 2360 1780
rect 2380 1700 2385 1780
rect 2355 1690 2385 1700
rect 2445 1780 2475 1790
rect 2445 1700 2450 1780
rect 2470 1700 2475 1780
rect 2445 1690 2475 1700
rect 2535 1780 2565 1790
rect 2535 1700 2540 1780
rect 2560 1700 2565 1780
rect 2535 1690 2565 1700
rect 2625 1780 2655 1790
rect 2625 1700 2630 1780
rect 2650 1700 2655 1780
rect 2625 1690 2655 1700
rect 2715 1780 2745 1790
rect 2715 1700 2720 1780
rect 2740 1700 2745 1780
rect 2715 1690 2745 1700
rect 2805 1780 2835 1790
rect 2805 1700 2810 1780
rect 2830 1700 2835 1780
rect 2805 1690 2835 1700
rect 2895 1780 2925 1790
rect 2895 1700 2900 1780
rect 2920 1700 2925 1780
rect 2895 1690 2925 1700
rect 2985 1780 3015 1790
rect 2985 1700 2990 1780
rect 3010 1700 3015 1780
rect 2985 1690 3015 1700
rect 3080 1780 3110 1790
rect 3080 1700 3085 1780
rect 3105 1700 3110 1780
rect 3080 1690 3110 1700
rect 3170 1780 3200 1790
rect 3170 1700 3175 1780
rect 3195 1700 3200 1780
rect 3170 1690 3200 1700
rect 3260 1780 3290 1790
rect 3260 1700 3265 1780
rect 3285 1700 3290 1780
rect 3260 1690 3290 1700
rect 3350 1780 3380 1790
rect 3350 1700 3355 1780
rect 3375 1700 3380 1780
rect 3350 1690 3380 1700
rect 3440 1780 3470 1790
rect 3440 1700 3445 1780
rect 3465 1700 3470 1780
rect 3440 1690 3470 1700
rect 3530 1780 3560 1790
rect 3530 1700 3535 1780
rect 3555 1700 3560 1780
rect 3530 1690 3560 1700
rect 3620 1780 3650 1790
rect 3620 1700 3625 1780
rect 3645 1700 3650 1780
rect 3620 1690 3650 1700
rect 3710 1780 3740 1790
rect 3710 1700 3715 1780
rect 3735 1700 3740 1780
rect 3710 1690 3740 1700
rect 3800 1780 3830 1790
rect 3800 1700 3805 1780
rect 3825 1700 3830 1780
rect 3800 1690 3830 1700
rect 3890 1780 3920 1790
rect 3890 1700 3895 1780
rect 3915 1700 3920 1780
rect 3890 1690 3920 1700
rect 3980 1780 4010 1790
rect 3980 1700 3985 1780
rect 4005 1700 4010 1780
rect 3980 1690 4010 1700
rect 4070 1780 4100 1790
rect 4070 1700 4075 1780
rect 4095 1700 4100 1780
rect 4070 1690 4100 1700
rect 4160 1780 4190 1790
rect 4160 1700 4165 1780
rect 4185 1700 4190 1780
rect 4160 1690 4190 1700
rect 4250 1780 4280 1790
rect 4250 1700 4255 1780
rect 4275 1700 4280 1780
rect 4250 1690 4280 1700
rect 4340 1780 4370 1790
rect 4340 1700 4345 1780
rect 4365 1700 4370 1780
rect 4340 1690 4370 1700
rect 4430 1780 4460 1790
rect 4430 1700 4435 1780
rect 4455 1700 4460 1780
rect 4430 1690 4460 1700
rect 4520 1780 4550 1790
rect 4520 1700 4525 1780
rect 4545 1700 4550 1780
rect 4520 1690 4550 1700
rect 4610 1780 4640 1790
rect 4610 1700 4615 1780
rect 4635 1700 4640 1780
rect 4610 1690 4640 1700
rect 4700 1780 4730 1790
rect 4700 1700 4705 1780
rect 4725 1700 4730 1780
rect 4700 1690 4730 1700
rect 4790 1780 4820 1790
rect 4790 1700 4795 1780
rect 4815 1700 4820 1780
rect 4790 1690 4820 1700
rect 4880 1780 4910 1790
rect 4880 1700 4885 1780
rect 4905 1700 4910 1780
rect 4880 1690 4910 1700
rect 4970 1780 5000 1790
rect 4970 1700 4975 1780
rect 4995 1700 5000 1780
rect 4970 1690 5000 1700
rect 5060 1780 5090 1790
rect 5060 1700 5065 1780
rect 5085 1700 5090 1780
rect 5060 1690 5090 1700
rect 5150 1780 5180 1790
rect 5150 1700 5155 1780
rect 5175 1700 5180 1780
rect 5150 1690 5180 1700
rect 5240 1780 5270 1790
rect 5240 1700 5245 1780
rect 5265 1700 5270 1780
rect 5240 1690 5270 1700
rect 5330 1780 5360 1790
rect 5330 1700 5335 1780
rect 5355 1700 5360 1780
rect 5330 1690 5360 1700
rect 5420 1780 5450 1790
rect 5420 1700 5425 1780
rect 5445 1700 5450 1780
rect 5420 1690 5450 1700
rect 5510 1780 5540 1790
rect 5510 1700 5515 1780
rect 5535 1700 5540 1780
rect 5510 1690 5540 1700
rect 5600 1780 5630 1790
rect 5600 1700 5605 1780
rect 5625 1700 5630 1780
rect 5600 1690 5630 1700
rect 5690 1780 5720 1790
rect 5690 1700 5695 1780
rect 5715 1700 5720 1780
rect 5690 1690 5720 1700
rect 5780 1780 5810 1790
rect 5780 1700 5785 1780
rect 5805 1700 5810 1780
rect 5780 1690 5810 1700
rect 5870 1780 5900 1790
rect 5870 1700 5875 1780
rect 5895 1700 5900 1780
rect 5870 1690 5900 1700
rect 5960 1780 5990 1790
rect 5960 1700 5965 1780
rect 5985 1700 5990 1780
rect 5960 1690 5990 1700
rect 6050 1780 6080 1790
rect 6050 1700 6055 1780
rect 6075 1700 6080 1780
rect 6050 1690 6080 1700
rect 6140 1780 6170 1790
rect 6140 1700 6145 1780
rect 6165 1700 6170 1780
rect 6140 1690 6170 1700
rect 6230 1780 6260 1790
rect 6230 1700 6235 1780
rect 6255 1700 6260 1780
rect 6230 1690 6260 1700
rect 6320 1780 6350 1790
rect 6320 1700 6325 1780
rect 6345 1700 6350 1780
rect 6320 1690 6350 1700
rect 6410 1780 6440 1790
rect 6410 1700 6415 1780
rect 6435 1700 6440 1780
rect 6410 1690 6440 1700
rect 6500 1780 6530 1790
rect 6500 1700 6505 1780
rect 6525 1700 6530 1780
rect 6500 1690 6530 1700
rect 6590 1780 6620 1790
rect 6590 1700 6595 1780
rect 6615 1700 6620 1780
rect 6590 1690 6620 1700
rect 6680 1780 6710 1790
rect 6680 1700 6685 1780
rect 6705 1700 6710 1780
rect 6680 1690 6710 1700
rect 6770 1780 6800 1790
rect 6770 1700 6775 1780
rect 6795 1700 6800 1780
rect 6770 1690 6800 1700
rect 6860 1780 6890 1790
rect 6860 1700 6865 1780
rect 6885 1700 6890 1780
rect 6860 1690 6890 1700
rect 6950 1780 6980 1790
rect 6950 1700 6955 1780
rect 6975 1700 6980 1780
rect 6950 1690 6980 1700
rect 7040 1780 7070 1790
rect 7040 1700 7045 1780
rect 7065 1700 7070 1780
rect 7040 1690 7070 1700
rect 7130 1780 7160 1790
rect 7130 1700 7135 1780
rect 7155 1700 7160 1780
rect 7130 1690 7160 1700
rect 7220 1780 7250 1790
rect 7220 1700 7225 1780
rect 7245 1700 7250 1780
rect 7220 1690 7250 1700
rect 7310 1780 7340 1790
rect 7310 1700 7315 1780
rect 7335 1700 7340 1780
rect 7310 1690 7340 1700
rect 7400 1780 7430 1790
rect 7400 1700 7405 1780
rect 7425 1700 7430 1780
rect 7400 1690 7430 1700
rect 7490 1780 7520 1790
rect 7490 1700 7495 1780
rect 7515 1700 7520 1780
rect 7490 1690 7520 1700
rect 7580 1780 7610 1790
rect 7580 1700 7585 1780
rect 7605 1700 7610 1780
rect 7580 1690 7610 1700
rect 7670 1780 7700 1790
rect 7670 1700 7675 1780
rect 7695 1700 7700 1780
rect 7670 1690 7700 1700
rect 7760 1780 7790 1790
rect 7760 1700 7765 1780
rect 7785 1700 7790 1780
rect 7760 1690 7790 1700
rect 7850 1780 7880 1790
rect 7850 1700 7855 1780
rect 7875 1700 7880 1780
rect 7850 1690 7880 1700
rect 7940 1780 7970 1790
rect 7940 1700 7945 1780
rect 7965 1700 7970 1780
rect 7940 1690 7970 1700
rect 8030 1780 8060 1790
rect 8030 1700 8035 1780
rect 8055 1700 8060 1780
rect 8030 1690 8060 1700
rect 8120 1780 8150 1790
rect 8120 1700 8125 1780
rect 8145 1700 8150 1780
rect 8120 1690 8150 1700
rect 8210 1780 8240 1790
rect 8210 1700 8215 1780
rect 8235 1700 8240 1780
rect 8210 1690 8240 1700
rect 8300 1780 8330 1790
rect 8300 1700 8305 1780
rect 8325 1700 8330 1780
rect 8300 1690 8330 1700
rect 8390 1780 8420 1790
rect 8390 1700 8395 1780
rect 8415 1700 8420 1780
rect 8390 1690 8420 1700
rect 8480 1780 8510 1790
rect 8480 1700 8485 1780
rect 8505 1700 8510 1780
rect 8480 1690 8510 1700
rect 8570 1780 8600 1790
rect 8570 1700 8575 1780
rect 8595 1700 8600 1780
rect 8570 1690 8600 1700
rect 8660 1780 8690 1790
rect 8660 1700 8665 1780
rect 8685 1700 8690 1780
rect 8660 1690 8690 1700
rect 8750 1780 8780 1790
rect 8750 1700 8755 1780
rect 8775 1700 8780 1780
rect 8750 1690 8780 1700
rect 8840 1780 8870 1790
rect 8840 1700 8845 1780
rect 8865 1700 8870 1780
rect 8840 1690 8870 1700
rect 8930 1780 8960 1790
rect 8930 1700 8935 1780
rect 8955 1700 8960 1780
rect 8930 1690 8960 1700
rect 9020 1780 9050 1790
rect 9020 1700 9025 1780
rect 9045 1700 9050 1780
rect 9020 1690 9050 1700
rect 9110 1780 9140 1790
rect 9110 1700 9115 1780
rect 9135 1700 9140 1780
rect 9110 1690 9140 1700
rect 9200 1780 9230 1790
rect 9200 1700 9205 1780
rect 9225 1700 9230 1780
rect 9200 1690 9230 1700
rect 9290 1780 9320 1790
rect 9290 1700 9295 1780
rect 9315 1700 9320 1780
rect 9290 1690 9320 1700
rect 9380 1780 9410 1790
rect 9380 1700 9385 1780
rect 9405 1700 9410 1780
rect 9380 1690 9410 1700
rect 9470 1780 9500 1790
rect 9470 1700 9475 1780
rect 9495 1700 9500 1780
rect 9470 1690 9500 1700
rect 9560 1780 9590 1790
rect 9560 1700 9565 1780
rect 9585 1700 9590 1780
rect 9560 1690 9590 1700
rect 9650 1780 9680 1790
rect 9650 1700 9655 1780
rect 9675 1700 9680 1780
rect 9650 1690 9680 1700
rect 9740 1780 9770 1790
rect 9740 1700 9745 1780
rect 9765 1700 9770 1780
rect 9740 1690 9770 1700
rect 9830 1780 9860 1790
rect 9830 1700 9835 1780
rect 9855 1700 9860 1780
rect 9830 1690 9860 1700
rect 9920 1780 9950 1790
rect 9920 1700 9925 1780
rect 9945 1700 9950 1780
rect 9920 1690 9950 1700
rect 10010 1780 10040 1790
rect 10010 1700 10015 1780
rect 10035 1700 10040 1780
rect 10010 1690 10040 1700
rect 10100 1780 10130 1790
rect 10100 1700 10105 1780
rect 10125 1700 10130 1780
rect 10100 1690 10130 1700
rect 10190 1780 10220 1790
rect 10190 1700 10195 1780
rect 10215 1700 10220 1780
rect 10190 1690 10220 1700
rect 10280 1780 10310 1790
rect 10280 1700 10285 1780
rect 10305 1700 10310 1780
rect 10280 1690 10310 1700
rect 10370 1780 10400 1790
rect 10370 1700 10375 1780
rect 10395 1700 10400 1780
rect 10370 1690 10400 1700
rect 10460 1780 10490 1790
rect 10460 1700 10465 1780
rect 10485 1700 10490 1780
rect 10460 1690 10490 1700
rect 10550 1780 10580 1790
rect 10550 1700 10555 1780
rect 10575 1700 10580 1780
rect 10550 1690 10580 1700
rect 10640 1780 10670 1790
rect 10640 1700 10645 1780
rect 10665 1700 10670 1780
rect 10640 1690 10670 1700
rect 10730 1690 10760 1790
rect 10820 1690 10850 1790
rect 10910 1690 10940 1790
rect 11000 1690 11030 1790
rect 11090 1690 11120 1790
rect 11180 1780 11210 1790
rect 11180 1700 11185 1780
rect 11205 1700 11210 1780
rect 11180 1690 11210 1700
rect -250 1425 -230 1690
rect -160 1465 -140 1690
rect -70 1505 -50 1690
rect 20 1545 40 1690
rect 110 1585 130 1690
rect 335 1670 355 1675
rect 515 1670 535 1675
rect 695 1670 715 1675
rect 875 1670 895 1675
rect 1055 1670 1075 1675
rect 1235 1670 1255 1675
rect 1415 1670 1435 1675
rect 1595 1670 1615 1675
rect 1775 1670 1795 1675
rect 1955 1670 1975 1675
rect 330 1665 360 1670
rect 330 1645 335 1665
rect 355 1645 360 1665
rect 330 1640 360 1645
rect 510 1665 540 1670
rect 510 1645 515 1665
rect 535 1645 540 1665
rect 510 1640 540 1645
rect 690 1665 720 1670
rect 690 1645 695 1665
rect 715 1645 720 1665
rect 690 1640 720 1645
rect 870 1665 900 1670
rect 870 1645 875 1665
rect 895 1645 900 1665
rect 870 1640 900 1645
rect 1050 1665 1080 1670
rect 1050 1645 1055 1665
rect 1075 1645 1080 1665
rect 1050 1640 1080 1645
rect 1230 1665 1260 1670
rect 1230 1645 1235 1665
rect 1255 1645 1260 1665
rect 1230 1640 1260 1645
rect 1410 1665 1440 1670
rect 1410 1645 1415 1665
rect 1435 1645 1440 1665
rect 1410 1640 1440 1645
rect 1590 1665 1620 1670
rect 1590 1645 1595 1665
rect 1615 1645 1620 1665
rect 1590 1640 1620 1645
rect 1770 1665 1800 1670
rect 1770 1645 1775 1665
rect 1795 1645 1800 1665
rect 1770 1640 1800 1645
rect 1950 1665 1980 1670
rect 1950 1645 1955 1665
rect 1975 1645 1980 1665
rect 1950 1640 1980 1645
rect 105 1580 135 1585
rect 105 1560 110 1580
rect 130 1560 135 1580
rect 105 1555 135 1560
rect 15 1540 45 1545
rect 15 1520 20 1540
rect 40 1520 45 1540
rect 15 1515 45 1520
rect -75 1500 -45 1505
rect -75 1480 -70 1500
rect -50 1480 -45 1500
rect -75 1475 -45 1480
rect -165 1460 -135 1465
rect -165 1440 -160 1460
rect -140 1440 -135 1460
rect -165 1435 -135 1440
rect -255 1420 -225 1425
rect -255 1400 -250 1420
rect -230 1400 -225 1420
rect -255 1395 -225 1400
rect -250 1090 -230 1395
rect -160 1090 -140 1435
rect -70 1090 -50 1475
rect 20 1090 40 1515
rect 110 1090 130 1555
rect 335 1545 355 1640
rect 515 1545 535 1640
rect 695 1545 715 1640
rect 875 1545 895 1640
rect 1055 1545 1075 1640
rect 1235 1545 1255 1640
rect 1415 1545 1435 1640
rect 1595 1545 1615 1640
rect 330 1540 360 1545
rect 330 1520 335 1540
rect 355 1520 360 1540
rect 330 1515 360 1520
rect 510 1540 540 1545
rect 510 1520 515 1540
rect 535 1520 540 1540
rect 510 1515 540 1520
rect 690 1540 720 1545
rect 690 1520 695 1540
rect 715 1520 720 1540
rect 690 1515 720 1520
rect 870 1540 900 1545
rect 870 1520 875 1540
rect 895 1520 900 1540
rect 870 1515 900 1520
rect 1050 1540 1080 1545
rect 1050 1520 1055 1540
rect 1075 1520 1080 1540
rect 1050 1515 1080 1520
rect 1230 1540 1260 1545
rect 1230 1520 1235 1540
rect 1255 1520 1260 1540
rect 1230 1515 1260 1520
rect 1410 1540 1440 1545
rect 1410 1520 1415 1540
rect 1435 1520 1440 1540
rect 1410 1515 1440 1520
rect 1590 1540 1620 1545
rect 1590 1520 1595 1540
rect 1615 1520 1620 1540
rect 1590 1515 1620 1520
rect 335 1510 355 1515
rect 515 1510 535 1515
rect 695 1510 715 1515
rect 875 1510 895 1515
rect 1055 1510 1075 1515
rect 1235 1510 1255 1515
rect 1415 1510 1435 1515
rect 1595 1510 1615 1515
rect 1775 1425 1795 1640
rect 1955 1425 1975 1640
rect 1770 1420 1800 1425
rect 1770 1400 1775 1420
rect 1795 1400 1800 1420
rect 1770 1395 1800 1400
rect 1950 1420 1980 1425
rect 1950 1400 1955 1420
rect 1975 1400 1980 1420
rect 1950 1395 1980 1400
rect 1775 1390 1795 1395
rect 1955 1390 1975 1395
rect 920 1385 940 1390
rect 915 1380 945 1385
rect 915 1360 920 1380
rect 940 1360 945 1380
rect 915 1355 945 1360
rect 605 1345 625 1350
rect 785 1345 805 1350
rect 600 1340 630 1345
rect 600 1320 605 1340
rect 625 1320 630 1340
rect 600 1315 630 1320
rect 780 1340 810 1345
rect 780 1320 785 1340
rect 805 1320 810 1340
rect 780 1315 810 1320
rect 245 1305 265 1310
rect 425 1305 445 1310
rect 240 1300 270 1305
rect 240 1280 245 1300
rect 265 1280 270 1300
rect 240 1275 270 1280
rect 420 1300 450 1305
rect 420 1280 425 1300
rect 445 1280 450 1300
rect 420 1275 450 1280
rect 245 1140 265 1275
rect 425 1140 445 1275
rect 605 1140 625 1315
rect 785 1140 805 1315
rect 240 1135 270 1140
rect 240 1115 245 1135
rect 265 1115 270 1135
rect 240 1110 270 1115
rect 420 1135 450 1140
rect 420 1115 425 1135
rect 445 1115 450 1135
rect 420 1110 450 1115
rect 600 1135 630 1140
rect 600 1115 605 1135
rect 625 1115 630 1135
rect 600 1110 630 1115
rect 780 1135 810 1140
rect 780 1115 785 1135
rect 805 1115 810 1135
rect 780 1110 810 1115
rect 245 1105 265 1110
rect 425 1105 445 1110
rect 605 1105 625 1110
rect 785 1105 805 1110
rect 920 1090 940 1355
rect 965 1345 985 1350
rect 1145 1345 1165 1350
rect 1685 1345 1705 1350
rect 1865 1345 1885 1350
rect 2000 1345 2020 1690
rect 2135 1670 2155 1675
rect 2315 1670 2335 1675
rect 2495 1670 2515 1675
rect 2675 1670 2695 1675
rect 2130 1665 2160 1670
rect 2130 1645 2135 1665
rect 2155 1645 2160 1665
rect 2130 1640 2160 1645
rect 2310 1665 2340 1670
rect 2310 1645 2315 1665
rect 2335 1645 2340 1665
rect 2310 1640 2340 1645
rect 2490 1665 2520 1670
rect 2490 1645 2495 1665
rect 2515 1645 2520 1665
rect 2490 1640 2520 1645
rect 2670 1665 2700 1670
rect 2670 1645 2675 1665
rect 2695 1645 2700 1665
rect 2670 1640 2700 1645
rect 2135 1425 2155 1640
rect 2315 1425 2335 1640
rect 2495 1425 2515 1640
rect 2675 1425 2695 1640
rect 2130 1420 2160 1425
rect 2130 1400 2135 1420
rect 2155 1400 2160 1420
rect 2130 1395 2160 1400
rect 2310 1420 2340 1425
rect 2310 1400 2315 1420
rect 2335 1400 2340 1420
rect 2310 1395 2340 1400
rect 2490 1420 2520 1425
rect 2490 1400 2495 1420
rect 2515 1400 2520 1420
rect 2490 1395 2520 1400
rect 2670 1420 2700 1425
rect 2670 1400 2675 1420
rect 2695 1400 2700 1420
rect 2670 1395 2700 1400
rect 2135 1390 2155 1395
rect 2315 1390 2335 1395
rect 2495 1390 2515 1395
rect 2675 1390 2695 1395
rect 2045 1345 2065 1350
rect 2225 1345 2245 1350
rect 2360 1345 2380 1350
rect 2405 1345 2425 1350
rect 2585 1345 2605 1350
rect 2720 1345 2740 1690
rect 2855 1670 2875 1675
rect 3035 1670 3055 1675
rect 3220 1670 3240 1675
rect 3400 1670 3420 1675
rect 3580 1670 3600 1675
rect 3760 1670 3780 1675
rect 2850 1665 2880 1670
rect 2850 1645 2855 1665
rect 2875 1645 2880 1665
rect 2850 1640 2880 1645
rect 3030 1665 3060 1670
rect 3030 1645 3035 1665
rect 3055 1645 3060 1665
rect 3030 1640 3060 1645
rect 3215 1665 3245 1670
rect 3215 1645 3220 1665
rect 3240 1645 3245 1665
rect 3215 1640 3245 1645
rect 3395 1665 3425 1670
rect 3395 1645 3400 1665
rect 3420 1645 3425 1665
rect 3395 1640 3425 1645
rect 3575 1665 3605 1670
rect 3575 1645 3580 1665
rect 3600 1645 3605 1665
rect 3575 1640 3605 1645
rect 3755 1665 3785 1670
rect 3755 1645 3760 1665
rect 3780 1645 3785 1665
rect 3755 1640 3785 1645
rect 2855 1425 2875 1640
rect 3035 1425 3055 1640
rect 3220 1425 3240 1640
rect 3400 1425 3420 1640
rect 3580 1425 3600 1640
rect 3760 1425 3780 1640
rect 2850 1420 2880 1425
rect 2850 1400 2855 1420
rect 2875 1400 2880 1420
rect 2850 1395 2880 1400
rect 3030 1420 3060 1425
rect 3030 1400 3035 1420
rect 3055 1400 3060 1420
rect 3030 1395 3060 1400
rect 3215 1420 3245 1425
rect 3215 1400 3220 1420
rect 3240 1400 3245 1420
rect 3215 1395 3245 1400
rect 3395 1420 3425 1425
rect 3395 1400 3400 1420
rect 3420 1400 3425 1420
rect 3395 1395 3425 1400
rect 3575 1420 3605 1425
rect 3575 1400 3580 1420
rect 3600 1400 3605 1420
rect 3575 1395 3605 1400
rect 3755 1420 3785 1425
rect 3755 1400 3760 1420
rect 3780 1400 3785 1420
rect 3755 1395 3785 1400
rect 2855 1390 2875 1395
rect 3035 1390 3055 1395
rect 3220 1390 3240 1395
rect 3400 1390 3420 1395
rect 3580 1390 3600 1395
rect 3760 1390 3780 1395
rect 2765 1345 2785 1350
rect 2945 1345 2965 1350
rect 3490 1345 3510 1350
rect 3670 1345 3690 1350
rect 960 1340 990 1345
rect 960 1320 965 1340
rect 985 1320 990 1340
rect 960 1315 990 1320
rect 1140 1340 1170 1345
rect 1140 1320 1145 1340
rect 1165 1320 1170 1340
rect 1140 1315 1170 1320
rect 1680 1340 1710 1345
rect 1680 1320 1685 1340
rect 1705 1320 1710 1340
rect 1680 1315 1710 1320
rect 1860 1340 1890 1345
rect 1860 1320 1865 1340
rect 1885 1320 1890 1340
rect 1860 1315 1890 1320
rect 1995 1340 2025 1345
rect 1995 1320 2000 1340
rect 2020 1320 2025 1340
rect 1995 1315 2025 1320
rect 2040 1340 2070 1345
rect 2040 1320 2045 1340
rect 2065 1320 2070 1340
rect 2040 1315 2070 1320
rect 2220 1340 2250 1345
rect 2220 1320 2225 1340
rect 2245 1320 2250 1340
rect 2220 1315 2250 1320
rect 2355 1340 2385 1345
rect 2355 1320 2360 1340
rect 2380 1320 2385 1340
rect 2355 1315 2385 1320
rect 2400 1340 2430 1345
rect 2400 1320 2405 1340
rect 2425 1320 2430 1340
rect 2400 1315 2430 1320
rect 2580 1340 2610 1345
rect 2580 1320 2585 1340
rect 2605 1320 2610 1340
rect 2580 1315 2610 1320
rect 2715 1340 2745 1345
rect 2715 1320 2720 1340
rect 2740 1320 2745 1340
rect 2715 1315 2745 1320
rect 2760 1340 2790 1345
rect 2760 1320 2765 1340
rect 2785 1320 2790 1340
rect 2760 1315 2790 1320
rect 2940 1340 2970 1345
rect 2940 1320 2945 1340
rect 2965 1320 2970 1340
rect 2940 1315 2970 1320
rect 3485 1340 3515 1345
rect 3485 1320 3490 1340
rect 3510 1320 3515 1340
rect 3485 1315 3515 1320
rect 3665 1340 3695 1345
rect 3665 1320 3670 1340
rect 3690 1320 3695 1340
rect 3665 1315 3695 1320
rect 965 1140 985 1315
rect 1145 1140 1165 1315
rect 1325 1305 1345 1310
rect 1505 1305 1525 1310
rect 1320 1300 1350 1305
rect 1320 1280 1325 1300
rect 1345 1280 1350 1300
rect 1320 1275 1350 1280
rect 1500 1300 1530 1305
rect 1500 1280 1505 1300
rect 1525 1280 1530 1300
rect 1500 1275 1530 1280
rect 1325 1140 1345 1275
rect 1505 1140 1525 1275
rect 1685 1140 1705 1315
rect 1865 1140 1885 1315
rect 2000 1310 2020 1315
rect 2045 1140 2065 1315
rect 2225 1140 2245 1315
rect 960 1135 990 1140
rect 960 1115 965 1135
rect 985 1115 990 1135
rect 960 1110 990 1115
rect 1140 1135 1170 1140
rect 1140 1115 1145 1135
rect 1165 1115 1170 1135
rect 1140 1110 1170 1115
rect 1320 1135 1350 1140
rect 1320 1115 1325 1135
rect 1345 1115 1350 1135
rect 1320 1110 1350 1115
rect 1500 1135 1530 1140
rect 1500 1115 1505 1135
rect 1525 1115 1530 1135
rect 1500 1110 1530 1115
rect 1680 1135 1710 1140
rect 1680 1115 1685 1135
rect 1705 1115 1710 1135
rect 1680 1110 1710 1115
rect 1860 1135 1890 1140
rect 1860 1115 1865 1135
rect 1885 1115 1890 1135
rect 1860 1110 1890 1115
rect 2040 1135 2070 1140
rect 2040 1115 2045 1135
rect 2065 1115 2070 1135
rect 2040 1110 2070 1115
rect 2220 1135 2250 1140
rect 2220 1115 2225 1135
rect 2245 1115 2250 1135
rect 2220 1110 2250 1115
rect 965 1105 985 1110
rect 1145 1105 1165 1110
rect 1325 1105 1345 1110
rect 1505 1105 1525 1110
rect 1685 1105 1705 1110
rect 1865 1105 1885 1110
rect 2045 1105 2065 1110
rect 2225 1105 2245 1110
rect 2360 1090 2380 1315
rect 2405 1140 2425 1315
rect 2585 1140 2605 1315
rect 2720 1310 2740 1315
rect 2765 1140 2785 1315
rect 2945 1140 2965 1315
rect 3130 1225 3150 1230
rect 3310 1225 3330 1230
rect 3125 1220 3155 1225
rect 3125 1200 3130 1220
rect 3150 1200 3155 1220
rect 3125 1195 3155 1200
rect 3305 1220 3335 1225
rect 3305 1200 3310 1220
rect 3330 1200 3335 1220
rect 3305 1195 3335 1200
rect 3130 1140 3150 1195
rect 3310 1140 3330 1195
rect 3490 1140 3510 1315
rect 3670 1140 3690 1315
rect 3805 1305 3825 1690
rect 3940 1670 3960 1675
rect 4120 1670 4140 1675
rect 4300 1670 4320 1675
rect 4480 1670 4500 1675
rect 4660 1670 4680 1675
rect 4840 1670 4860 1675
rect 5020 1670 5040 1675
rect 5200 1670 5220 1675
rect 3935 1665 3965 1670
rect 3935 1645 3940 1665
rect 3960 1645 3965 1665
rect 3935 1640 3965 1645
rect 4115 1665 4145 1670
rect 4115 1645 4120 1665
rect 4140 1645 4145 1665
rect 4115 1640 4145 1645
rect 4295 1665 4325 1670
rect 4295 1645 4300 1665
rect 4320 1645 4325 1665
rect 4295 1640 4325 1645
rect 4475 1665 4505 1670
rect 4475 1645 4480 1665
rect 4500 1645 4505 1665
rect 4475 1640 4505 1645
rect 4655 1665 4685 1670
rect 4655 1645 4660 1665
rect 4680 1645 4685 1665
rect 4655 1640 4685 1645
rect 4835 1665 4865 1670
rect 4835 1645 4840 1665
rect 4860 1645 4865 1665
rect 4835 1640 4865 1645
rect 5015 1665 5045 1670
rect 5015 1645 5020 1665
rect 5040 1645 5045 1665
rect 5015 1640 5045 1645
rect 5195 1665 5225 1670
rect 5195 1645 5200 1665
rect 5220 1645 5225 1665
rect 5195 1640 5225 1645
rect 3940 1425 3960 1640
rect 4120 1425 4140 1640
rect 4300 1425 4320 1640
rect 4480 1425 4500 1640
rect 4660 1505 4680 1640
rect 4840 1505 4860 1640
rect 5020 1505 5040 1640
rect 5200 1505 5220 1640
rect 4655 1500 4685 1505
rect 4655 1480 4660 1500
rect 4680 1480 4685 1500
rect 4655 1475 4685 1480
rect 4835 1500 4865 1505
rect 4835 1480 4840 1500
rect 4860 1480 4865 1500
rect 4835 1475 4865 1480
rect 5015 1500 5045 1505
rect 5015 1480 5020 1500
rect 5040 1480 5045 1500
rect 5015 1475 5045 1480
rect 5195 1500 5225 1505
rect 5195 1480 5200 1500
rect 5220 1480 5225 1500
rect 5195 1475 5225 1480
rect 4660 1470 4680 1475
rect 4840 1470 4860 1475
rect 5020 1470 5040 1475
rect 5200 1470 5220 1475
rect 3935 1420 3965 1425
rect 3935 1400 3940 1420
rect 3960 1400 3965 1420
rect 3935 1395 3965 1400
rect 4115 1420 4145 1425
rect 4115 1400 4120 1420
rect 4140 1400 4145 1420
rect 4115 1395 4145 1400
rect 4295 1420 4325 1425
rect 4295 1400 4300 1420
rect 4320 1400 4325 1420
rect 4295 1395 4325 1400
rect 4475 1420 4505 1425
rect 4475 1400 4480 1420
rect 4500 1400 4505 1420
rect 4475 1395 4505 1400
rect 3940 1390 3960 1395
rect 4120 1390 4140 1395
rect 4300 1390 4320 1395
rect 4480 1390 4500 1395
rect 3850 1345 3870 1350
rect 4030 1345 4050 1350
rect 4930 1345 4950 1350
rect 5110 1345 5130 1350
rect 3845 1340 3875 1345
rect 3845 1320 3850 1340
rect 3870 1320 3875 1340
rect 3845 1315 3875 1320
rect 4025 1340 4055 1345
rect 4025 1320 4030 1340
rect 4050 1320 4055 1340
rect 4025 1315 4055 1320
rect 4925 1340 4955 1345
rect 4925 1320 4930 1340
rect 4950 1320 4955 1340
rect 4925 1315 4955 1320
rect 5105 1340 5135 1345
rect 5105 1320 5110 1340
rect 5130 1320 5135 1340
rect 5105 1315 5135 1320
rect 3800 1300 3830 1305
rect 3800 1280 3805 1300
rect 3825 1280 3830 1300
rect 3800 1275 3830 1280
rect 2400 1135 2430 1140
rect 2400 1115 2405 1135
rect 2425 1115 2430 1135
rect 2400 1110 2430 1115
rect 2580 1135 2610 1140
rect 2580 1115 2585 1135
rect 2605 1115 2610 1135
rect 2580 1110 2610 1115
rect 2760 1135 2790 1140
rect 2760 1115 2765 1135
rect 2785 1115 2790 1135
rect 2760 1110 2790 1115
rect 2940 1135 2970 1140
rect 2940 1115 2945 1135
rect 2965 1115 2970 1135
rect 2940 1110 2970 1115
rect 3125 1135 3155 1140
rect 3125 1115 3130 1135
rect 3150 1115 3155 1135
rect 3125 1110 3155 1115
rect 3305 1135 3335 1140
rect 3305 1115 3310 1135
rect 3330 1115 3335 1135
rect 3305 1110 3335 1115
rect 3485 1135 3515 1140
rect 3485 1115 3490 1135
rect 3510 1115 3515 1135
rect 3485 1110 3515 1115
rect 3665 1135 3695 1140
rect 3665 1115 3670 1135
rect 3690 1115 3695 1135
rect 3665 1110 3695 1115
rect 2405 1105 2425 1110
rect 2585 1105 2605 1110
rect 2765 1105 2785 1110
rect 2945 1105 2965 1110
rect 3130 1105 3150 1110
rect 3310 1105 3330 1110
rect 3490 1105 3510 1110
rect 3670 1105 3690 1110
rect 3805 1090 3825 1275
rect 3850 1140 3870 1315
rect 4030 1140 4050 1315
rect 4210 1225 4230 1230
rect 4390 1225 4410 1230
rect 4570 1225 4590 1230
rect 4750 1225 4770 1230
rect 4205 1220 4235 1225
rect 4205 1200 4210 1220
rect 4230 1200 4235 1220
rect 4205 1195 4235 1200
rect 4385 1220 4415 1225
rect 4385 1200 4390 1220
rect 4410 1200 4415 1220
rect 4385 1195 4415 1200
rect 4565 1220 4595 1225
rect 4565 1200 4570 1220
rect 4590 1200 4595 1220
rect 4565 1195 4595 1200
rect 4745 1220 4775 1225
rect 4745 1200 4750 1220
rect 4770 1200 4775 1220
rect 4745 1195 4775 1200
rect 4210 1140 4230 1195
rect 4390 1140 4410 1195
rect 4570 1140 4590 1195
rect 4750 1140 4770 1195
rect 4930 1140 4950 1315
rect 5110 1140 5130 1315
rect 5245 1225 5265 1690
rect 5380 1670 5400 1675
rect 5560 1670 5580 1675
rect 5740 1670 5760 1675
rect 5920 1670 5940 1675
rect 6100 1670 6120 1675
rect 6280 1670 6300 1675
rect 6460 1670 6480 1675
rect 6640 1670 6660 1675
rect 5375 1665 5405 1670
rect 5375 1645 5380 1665
rect 5400 1645 5405 1665
rect 5375 1640 5405 1645
rect 5555 1665 5585 1670
rect 5555 1645 5560 1665
rect 5580 1645 5585 1665
rect 5555 1640 5585 1645
rect 5735 1665 5765 1670
rect 5735 1645 5740 1665
rect 5760 1645 5765 1665
rect 5735 1640 5765 1645
rect 5915 1665 5945 1670
rect 5915 1645 5920 1665
rect 5940 1645 5945 1665
rect 5915 1640 5945 1645
rect 6095 1665 6125 1670
rect 6095 1645 6100 1665
rect 6120 1645 6125 1665
rect 6095 1640 6125 1645
rect 6275 1665 6305 1670
rect 6275 1645 6280 1665
rect 6300 1645 6305 1665
rect 6275 1640 6305 1645
rect 6455 1665 6485 1670
rect 6455 1645 6460 1665
rect 6480 1645 6485 1665
rect 6455 1640 6485 1645
rect 6635 1665 6665 1670
rect 6635 1645 6640 1665
rect 6660 1645 6665 1665
rect 6635 1640 6665 1645
rect 5380 1505 5400 1640
rect 5560 1505 5580 1640
rect 5740 1505 5760 1640
rect 5920 1505 5940 1640
rect 5375 1500 5405 1505
rect 5375 1480 5380 1500
rect 5400 1480 5405 1500
rect 5375 1475 5405 1480
rect 5555 1500 5585 1505
rect 5555 1480 5560 1500
rect 5580 1480 5585 1500
rect 5555 1475 5585 1480
rect 5735 1500 5765 1505
rect 5735 1480 5740 1500
rect 5760 1480 5765 1500
rect 5735 1475 5765 1480
rect 5915 1500 5945 1505
rect 5915 1480 5920 1500
rect 5940 1480 5945 1500
rect 5915 1475 5945 1480
rect 5380 1470 5400 1475
rect 5560 1470 5580 1475
rect 5740 1470 5760 1475
rect 5920 1470 5940 1475
rect 6100 1425 6120 1640
rect 6280 1425 6300 1640
rect 6460 1425 6480 1640
rect 6640 1425 6660 1640
rect 6685 1425 6705 1690
rect 6730 1425 6750 1430
rect 6095 1420 6125 1425
rect 6095 1400 6100 1420
rect 6120 1400 6125 1420
rect 6095 1395 6125 1400
rect 6275 1420 6305 1425
rect 6275 1400 6280 1420
rect 6300 1400 6305 1420
rect 6275 1395 6305 1400
rect 6455 1420 6485 1425
rect 6455 1400 6460 1420
rect 6480 1400 6485 1420
rect 6455 1395 6485 1400
rect 6635 1420 6665 1425
rect 6635 1400 6640 1420
rect 6660 1400 6665 1420
rect 6635 1395 6665 1400
rect 6680 1420 6710 1425
rect 6680 1400 6685 1420
rect 6705 1400 6710 1420
rect 6680 1395 6710 1400
rect 6725 1420 6755 1425
rect 6725 1400 6730 1420
rect 6750 1400 6755 1420
rect 6725 1395 6755 1400
rect 6100 1390 6120 1395
rect 6280 1390 6300 1395
rect 6460 1390 6480 1395
rect 6640 1390 6660 1395
rect 5290 1345 5310 1350
rect 5470 1345 5490 1350
rect 6370 1345 6390 1350
rect 6550 1345 6570 1350
rect 5285 1340 5315 1345
rect 5285 1320 5290 1340
rect 5310 1320 5315 1340
rect 5285 1315 5315 1320
rect 5465 1340 5495 1345
rect 5465 1320 5470 1340
rect 5490 1320 5495 1340
rect 5465 1315 5495 1320
rect 6365 1340 6395 1345
rect 6365 1320 6370 1340
rect 6390 1320 6395 1340
rect 6365 1315 6395 1320
rect 6545 1340 6575 1345
rect 6545 1320 6550 1340
rect 6570 1320 6575 1340
rect 6545 1315 6575 1320
rect 5240 1220 5270 1225
rect 5240 1200 5245 1220
rect 5265 1200 5270 1220
rect 5240 1195 5270 1200
rect 3845 1135 3875 1140
rect 3845 1115 3850 1135
rect 3870 1115 3875 1135
rect 3845 1110 3875 1115
rect 4025 1135 4055 1140
rect 4025 1115 4030 1135
rect 4050 1115 4055 1135
rect 4025 1110 4055 1115
rect 4205 1135 4235 1140
rect 4205 1115 4210 1135
rect 4230 1115 4235 1135
rect 4205 1110 4235 1115
rect 4385 1135 4415 1140
rect 4385 1115 4390 1135
rect 4410 1115 4415 1135
rect 4385 1110 4415 1115
rect 4565 1135 4595 1140
rect 4565 1115 4570 1135
rect 4590 1115 4595 1135
rect 4565 1110 4595 1115
rect 4745 1135 4775 1140
rect 4745 1115 4750 1135
rect 4770 1115 4775 1135
rect 4745 1110 4775 1115
rect 4925 1135 4955 1140
rect 4925 1115 4930 1135
rect 4950 1115 4955 1135
rect 4925 1110 4955 1115
rect 5105 1135 5135 1140
rect 5105 1115 5110 1135
rect 5130 1115 5135 1135
rect 5105 1110 5135 1115
rect 3850 1105 3870 1110
rect 4030 1105 4050 1110
rect 4210 1105 4230 1110
rect 4390 1105 4410 1110
rect 4570 1105 4590 1110
rect 4750 1105 4770 1110
rect 4930 1105 4950 1110
rect 5110 1105 5130 1110
rect 5245 1090 5265 1195
rect 5290 1140 5310 1315
rect 5470 1140 5490 1315
rect 6010 1305 6030 1310
rect 6190 1305 6210 1310
rect 6005 1300 6035 1305
rect 6005 1280 6010 1300
rect 6030 1280 6035 1300
rect 6005 1275 6035 1280
rect 6185 1300 6215 1305
rect 6185 1280 6190 1300
rect 6210 1280 6215 1300
rect 6185 1275 6215 1280
rect 5650 1225 5670 1230
rect 5830 1225 5850 1230
rect 5645 1220 5675 1225
rect 5645 1200 5650 1220
rect 5670 1200 5675 1220
rect 5645 1195 5675 1200
rect 5825 1220 5855 1225
rect 5825 1200 5830 1220
rect 5850 1200 5855 1220
rect 5825 1195 5855 1200
rect 5650 1140 5670 1195
rect 5830 1140 5850 1195
rect 6010 1140 6030 1275
rect 6190 1140 6210 1275
rect 6370 1140 6390 1315
rect 6550 1140 6570 1315
rect 5285 1135 5315 1140
rect 5285 1115 5290 1135
rect 5310 1115 5315 1135
rect 5285 1110 5315 1115
rect 5465 1135 5495 1140
rect 5465 1115 5470 1135
rect 5490 1115 5495 1135
rect 5465 1110 5495 1115
rect 5645 1135 5675 1140
rect 5645 1115 5650 1135
rect 5670 1115 5675 1135
rect 5645 1110 5675 1115
rect 5825 1135 5855 1140
rect 5825 1115 5830 1135
rect 5850 1115 5855 1135
rect 5825 1110 5855 1115
rect 6005 1135 6035 1140
rect 6005 1115 6010 1135
rect 6030 1115 6035 1135
rect 6005 1110 6035 1115
rect 6185 1135 6215 1140
rect 6185 1115 6190 1135
rect 6210 1115 6215 1135
rect 6185 1110 6215 1115
rect 6365 1135 6395 1140
rect 6365 1115 6370 1135
rect 6390 1115 6395 1135
rect 6365 1110 6395 1115
rect 6545 1135 6575 1140
rect 6545 1115 6550 1135
rect 6570 1115 6575 1135
rect 6545 1110 6575 1115
rect 5290 1105 5310 1110
rect 5470 1105 5490 1110
rect 5650 1105 5670 1110
rect 5830 1105 5850 1110
rect 6010 1105 6030 1110
rect 6190 1105 6210 1110
rect 6370 1105 6390 1110
rect 6550 1105 6570 1110
rect 6685 1090 6705 1395
rect 6730 1140 6750 1395
rect 6775 1305 6795 1690
rect 6820 1670 6840 1675
rect 6815 1665 6845 1670
rect 6815 1645 6820 1665
rect 6840 1645 6845 1665
rect 6815 1640 6845 1645
rect 6820 1585 6840 1640
rect 6815 1580 6845 1585
rect 6815 1560 6820 1580
rect 6840 1560 6845 1580
rect 6815 1555 6845 1560
rect 6820 1550 6840 1555
rect 6865 1425 6885 1690
rect 7000 1670 7020 1675
rect 7180 1670 7200 1675
rect 7360 1670 7380 1675
rect 7540 1670 7560 1675
rect 7720 1670 7740 1675
rect 7900 1670 7920 1675
rect 6995 1665 7025 1670
rect 6995 1645 7000 1665
rect 7020 1645 7025 1665
rect 6995 1640 7025 1645
rect 7175 1665 7205 1670
rect 7175 1645 7180 1665
rect 7200 1645 7205 1665
rect 7175 1640 7205 1645
rect 7355 1665 7385 1670
rect 7355 1645 7360 1665
rect 7380 1645 7385 1665
rect 7355 1640 7385 1645
rect 7535 1665 7565 1670
rect 7535 1645 7540 1665
rect 7560 1645 7565 1665
rect 7535 1640 7565 1645
rect 7715 1665 7745 1670
rect 7715 1645 7720 1665
rect 7740 1645 7745 1665
rect 7715 1640 7745 1645
rect 7895 1665 7925 1670
rect 7895 1645 7900 1665
rect 7920 1645 7925 1665
rect 7895 1640 7925 1645
rect 7000 1425 7020 1640
rect 7180 1425 7200 1640
rect 7360 1425 7380 1640
rect 7540 1425 7560 1640
rect 7720 1465 7740 1640
rect 7900 1465 7920 1640
rect 7945 1545 7965 1690
rect 8080 1670 8100 1675
rect 8260 1670 8280 1675
rect 8075 1665 8105 1670
rect 8075 1645 8080 1665
rect 8100 1645 8105 1665
rect 8075 1640 8105 1645
rect 8255 1665 8285 1670
rect 8255 1645 8260 1665
rect 8280 1645 8285 1665
rect 8255 1640 8285 1645
rect 7940 1540 7970 1545
rect 7940 1520 7945 1540
rect 7965 1520 7970 1540
rect 7940 1515 7970 1520
rect 7945 1510 7965 1515
rect 8080 1505 8100 1640
rect 8260 1505 8280 1640
rect 8305 1505 8325 1690
rect 8440 1670 8460 1675
rect 8620 1670 8640 1675
rect 8435 1665 8465 1670
rect 8435 1645 8440 1665
rect 8460 1645 8465 1665
rect 8435 1640 8465 1645
rect 8615 1665 8645 1670
rect 8615 1645 8620 1665
rect 8640 1645 8645 1665
rect 8615 1640 8645 1645
rect 8440 1505 8460 1640
rect 8620 1505 8640 1640
rect 8665 1545 8685 1690
rect 8800 1670 8820 1675
rect 8980 1670 9000 1675
rect 9160 1670 9180 1675
rect 9340 1670 9360 1675
rect 8795 1665 8825 1670
rect 8795 1645 8800 1665
rect 8820 1645 8825 1665
rect 8795 1640 8825 1645
rect 8975 1665 9005 1670
rect 8975 1645 8980 1665
rect 9000 1645 9005 1665
rect 8975 1640 9005 1645
rect 9155 1665 9185 1670
rect 9155 1645 9160 1665
rect 9180 1645 9185 1665
rect 9155 1640 9185 1645
rect 9335 1665 9365 1670
rect 9335 1645 9340 1665
rect 9360 1645 9365 1665
rect 9335 1640 9365 1645
rect 8660 1540 8690 1545
rect 8660 1520 8665 1540
rect 8685 1520 8690 1540
rect 8660 1515 8690 1520
rect 8665 1510 8685 1515
rect 8075 1500 8105 1505
rect 8075 1480 8080 1500
rect 8100 1480 8105 1500
rect 8075 1475 8105 1480
rect 8255 1500 8285 1505
rect 8255 1480 8260 1500
rect 8280 1480 8285 1500
rect 8255 1475 8285 1480
rect 8300 1500 8330 1505
rect 8300 1480 8305 1500
rect 8325 1480 8330 1500
rect 8300 1475 8330 1480
rect 8435 1500 8465 1505
rect 8435 1480 8440 1500
rect 8460 1480 8465 1500
rect 8435 1475 8465 1480
rect 8615 1500 8645 1505
rect 8615 1480 8620 1500
rect 8640 1480 8645 1500
rect 8615 1475 8645 1480
rect 8080 1470 8100 1475
rect 8260 1470 8280 1475
rect 7715 1460 7745 1465
rect 7715 1440 7720 1460
rect 7740 1440 7745 1460
rect 7715 1435 7745 1440
rect 7895 1460 7925 1465
rect 7895 1440 7900 1460
rect 7920 1440 7925 1460
rect 7895 1435 7925 1440
rect 7720 1430 7740 1435
rect 7900 1430 7920 1435
rect 6860 1420 6890 1425
rect 6860 1400 6865 1420
rect 6885 1400 6890 1420
rect 6860 1395 6890 1400
rect 6995 1420 7025 1425
rect 6995 1400 7000 1420
rect 7020 1400 7025 1420
rect 6995 1395 7025 1400
rect 7175 1420 7205 1425
rect 7175 1400 7180 1420
rect 7200 1400 7205 1420
rect 7175 1395 7205 1400
rect 7355 1420 7385 1425
rect 7355 1400 7360 1420
rect 7380 1400 7385 1420
rect 7355 1395 7385 1400
rect 7535 1420 7565 1425
rect 7535 1400 7540 1420
rect 7560 1400 7565 1420
rect 7535 1395 7565 1400
rect 6770 1300 6800 1305
rect 6770 1280 6775 1300
rect 6795 1280 6800 1300
rect 6770 1275 6800 1280
rect 6775 1270 6795 1275
rect 6725 1135 6755 1140
rect 6725 1115 6730 1135
rect 6750 1115 6755 1135
rect 6725 1110 6755 1115
rect 6730 1105 6750 1110
rect 6865 1090 6885 1395
rect 7000 1390 7020 1395
rect 7180 1390 7200 1395
rect 7360 1390 7380 1395
rect 7540 1390 7560 1395
rect 6910 1345 6930 1350
rect 7090 1345 7110 1350
rect 7990 1345 8010 1350
rect 8170 1345 8190 1350
rect 6905 1340 6935 1345
rect 6905 1320 6910 1340
rect 6930 1320 6935 1340
rect 6905 1315 6935 1320
rect 7085 1340 7115 1345
rect 7085 1320 7090 1340
rect 7110 1320 7115 1340
rect 7085 1315 7115 1320
rect 7985 1340 8015 1345
rect 7985 1320 7990 1340
rect 8010 1320 8015 1340
rect 7985 1315 8015 1320
rect 8165 1340 8195 1345
rect 8165 1320 8170 1340
rect 8190 1320 8195 1340
rect 8165 1315 8195 1320
rect 6910 1140 6930 1315
rect 7090 1140 7110 1315
rect 7270 1305 7290 1310
rect 7450 1305 7470 1310
rect 7630 1305 7650 1310
rect 7810 1305 7830 1310
rect 7265 1300 7295 1305
rect 7265 1280 7270 1300
rect 7290 1280 7295 1300
rect 7265 1275 7295 1280
rect 7445 1300 7475 1305
rect 7445 1280 7450 1300
rect 7470 1280 7475 1300
rect 7445 1275 7475 1280
rect 7625 1300 7655 1305
rect 7625 1280 7630 1300
rect 7650 1280 7655 1300
rect 7625 1275 7655 1280
rect 7805 1300 7835 1305
rect 7805 1280 7810 1300
rect 7830 1280 7835 1300
rect 7805 1275 7835 1280
rect 7270 1140 7290 1275
rect 7450 1140 7470 1275
rect 7630 1140 7650 1275
rect 7810 1140 7830 1275
rect 7990 1140 8010 1315
rect 8170 1140 8190 1315
rect 6905 1135 6935 1140
rect 6905 1115 6910 1135
rect 6930 1115 6935 1135
rect 6905 1110 6935 1115
rect 7085 1135 7115 1140
rect 7085 1115 7090 1135
rect 7110 1115 7115 1135
rect 7085 1110 7115 1115
rect 7265 1135 7295 1140
rect 7265 1115 7270 1135
rect 7290 1115 7295 1135
rect 7265 1110 7295 1115
rect 7445 1135 7475 1140
rect 7445 1115 7450 1135
rect 7470 1115 7475 1135
rect 7445 1110 7475 1115
rect 7625 1135 7655 1140
rect 7625 1115 7630 1135
rect 7650 1115 7655 1135
rect 7625 1110 7655 1115
rect 7805 1135 7835 1140
rect 7805 1115 7810 1135
rect 7830 1115 7835 1135
rect 7805 1110 7835 1115
rect 7985 1135 8015 1140
rect 7985 1115 7990 1135
rect 8010 1115 8015 1135
rect 7985 1110 8015 1115
rect 8165 1135 8195 1140
rect 8165 1115 8170 1135
rect 8190 1115 8195 1135
rect 8165 1110 8195 1115
rect 6910 1105 6930 1110
rect 7090 1105 7110 1110
rect 7270 1105 7290 1110
rect 7450 1105 7470 1110
rect 7630 1105 7650 1110
rect 7810 1105 7830 1110
rect 7990 1105 8010 1110
rect 8170 1105 8190 1110
rect 8305 1090 8325 1475
rect 8440 1470 8460 1475
rect 8620 1470 8640 1475
rect 8800 1465 8820 1640
rect 8980 1465 9000 1640
rect 9160 1465 9180 1640
rect 9340 1465 9360 1640
rect 9385 1545 9405 1690
rect 9520 1670 9540 1675
rect 9700 1670 9720 1675
rect 9515 1665 9545 1670
rect 9515 1645 9520 1665
rect 9540 1645 9545 1665
rect 9515 1640 9545 1645
rect 9695 1665 9725 1670
rect 9695 1645 9700 1665
rect 9720 1645 9725 1665
rect 9695 1640 9725 1645
rect 9380 1540 9410 1545
rect 9380 1520 9385 1540
rect 9405 1520 9410 1540
rect 9380 1515 9410 1520
rect 9385 1510 9405 1515
rect 9385 1465 9405 1470
rect 9520 1465 9540 1640
rect 9700 1465 9720 1640
rect 9745 1465 9765 1690
rect 9880 1670 9900 1675
rect 10060 1670 10080 1675
rect 9875 1665 9905 1670
rect 9875 1645 9880 1665
rect 9900 1645 9905 1665
rect 9875 1640 9905 1645
rect 10055 1665 10085 1670
rect 10055 1645 10060 1665
rect 10080 1645 10085 1665
rect 10055 1640 10085 1645
rect 9880 1465 9900 1640
rect 10060 1465 10080 1640
rect 10105 1545 10125 1690
rect 10240 1670 10260 1675
rect 10420 1670 10440 1675
rect 10235 1665 10265 1670
rect 10235 1645 10240 1665
rect 10260 1645 10265 1665
rect 10235 1640 10265 1645
rect 10415 1665 10445 1670
rect 10415 1645 10420 1665
rect 10440 1645 10445 1665
rect 10415 1640 10445 1645
rect 10100 1540 10130 1545
rect 10100 1520 10105 1540
rect 10125 1520 10130 1540
rect 10100 1515 10130 1520
rect 10105 1510 10125 1515
rect 10105 1465 10125 1470
rect 10240 1465 10260 1640
rect 10420 1465 10440 1640
rect 10510 1585 10530 1590
rect 10555 1585 10575 1690
rect 10600 1670 10620 1675
rect 10595 1665 10625 1670
rect 10595 1645 10600 1665
rect 10620 1645 10625 1665
rect 10595 1640 10625 1645
rect 10505 1580 10535 1585
rect 10505 1560 10510 1580
rect 10530 1560 10535 1580
rect 10505 1555 10535 1560
rect 10550 1580 10580 1585
rect 10550 1560 10555 1580
rect 10575 1560 10580 1580
rect 10550 1555 10580 1560
rect 8795 1460 8825 1465
rect 8795 1440 8800 1460
rect 8820 1440 8825 1460
rect 8795 1435 8825 1440
rect 8975 1460 9005 1465
rect 8975 1440 8980 1460
rect 9000 1440 9005 1460
rect 8975 1435 9005 1440
rect 9155 1460 9185 1465
rect 9155 1440 9160 1460
rect 9180 1440 9185 1460
rect 9155 1435 9185 1440
rect 9335 1460 9365 1465
rect 9335 1440 9340 1460
rect 9360 1440 9365 1460
rect 9335 1435 9365 1440
rect 9380 1460 9410 1465
rect 9380 1440 9385 1460
rect 9405 1440 9410 1460
rect 9380 1435 9410 1440
rect 9515 1460 9545 1465
rect 9515 1440 9520 1460
rect 9540 1440 9545 1460
rect 9515 1435 9545 1440
rect 9695 1460 9725 1465
rect 9695 1440 9700 1460
rect 9720 1440 9725 1460
rect 9695 1435 9725 1440
rect 9740 1460 9770 1465
rect 9740 1440 9745 1460
rect 9765 1440 9770 1460
rect 9740 1435 9770 1440
rect 9875 1460 9905 1465
rect 9875 1440 9880 1460
rect 9900 1440 9905 1460
rect 9875 1435 9905 1440
rect 10055 1460 10085 1465
rect 10055 1440 10060 1460
rect 10080 1440 10085 1460
rect 10055 1435 10085 1440
rect 10100 1460 10130 1465
rect 10100 1440 10105 1460
rect 10125 1440 10130 1460
rect 10100 1435 10130 1440
rect 10235 1460 10265 1465
rect 10235 1440 10240 1460
rect 10260 1440 10265 1460
rect 10235 1435 10265 1440
rect 10415 1460 10445 1465
rect 10415 1440 10420 1460
rect 10440 1440 10445 1460
rect 10415 1435 10445 1440
rect 8800 1430 8820 1435
rect 8980 1430 9000 1435
rect 9160 1430 9180 1435
rect 9340 1430 9360 1435
rect 8350 1345 8370 1350
rect 8530 1345 8550 1350
rect 9250 1345 9270 1350
rect 8345 1340 8375 1345
rect 8345 1320 8350 1340
rect 8370 1320 8375 1340
rect 8345 1315 8375 1320
rect 8525 1340 8555 1345
rect 8525 1320 8530 1340
rect 8550 1320 8555 1340
rect 8525 1315 8555 1320
rect 9245 1340 9275 1345
rect 9245 1320 9250 1340
rect 9270 1320 9275 1340
rect 9245 1315 9275 1320
rect 8350 1140 8370 1315
rect 8530 1140 8550 1315
rect 8710 1305 8730 1310
rect 8890 1305 8910 1310
rect 9070 1305 9090 1310
rect 8705 1300 8735 1305
rect 8705 1280 8710 1300
rect 8730 1280 8735 1300
rect 8705 1275 8735 1280
rect 8885 1300 8915 1305
rect 8885 1280 8890 1300
rect 8910 1280 8915 1300
rect 8885 1275 8915 1280
rect 9065 1300 9095 1305
rect 9065 1280 9070 1300
rect 9090 1280 9095 1300
rect 9065 1275 9095 1280
rect 8710 1140 8730 1275
rect 8890 1140 8910 1275
rect 9070 1140 9090 1275
rect 9250 1140 9270 1315
rect 8345 1135 8375 1140
rect 8345 1115 8350 1135
rect 8370 1115 8375 1135
rect 8345 1110 8375 1115
rect 8525 1135 8555 1140
rect 8525 1115 8530 1135
rect 8550 1115 8555 1135
rect 8525 1110 8555 1115
rect 8705 1135 8735 1140
rect 8705 1115 8710 1135
rect 8730 1115 8735 1135
rect 8705 1110 8735 1115
rect 8885 1135 8915 1140
rect 8885 1115 8890 1135
rect 8910 1115 8915 1135
rect 8885 1110 8915 1115
rect 9065 1135 9095 1140
rect 9065 1115 9070 1135
rect 9090 1115 9095 1135
rect 9065 1110 9095 1115
rect 9245 1135 9275 1140
rect 9245 1115 9250 1135
rect 9270 1115 9275 1135
rect 9245 1110 9275 1115
rect 8350 1105 8370 1110
rect 8530 1105 8550 1110
rect 8710 1105 8730 1110
rect 8890 1105 8910 1110
rect 9070 1105 9090 1110
rect 9250 1105 9270 1110
rect 9385 1090 9405 1435
rect 9520 1430 9540 1435
rect 9700 1430 9720 1435
rect 9745 1430 9765 1435
rect 9880 1430 9900 1435
rect 10060 1430 10080 1435
rect 9430 1345 9450 1350
rect 9970 1345 9990 1350
rect 9425 1340 9455 1345
rect 9425 1320 9430 1340
rect 9450 1320 9455 1340
rect 9425 1315 9455 1320
rect 9965 1340 9995 1345
rect 9965 1320 9970 1340
rect 9990 1320 9995 1340
rect 9965 1315 9995 1320
rect 9430 1140 9450 1315
rect 9610 1305 9630 1310
rect 9790 1305 9810 1310
rect 9605 1300 9635 1305
rect 9605 1280 9610 1300
rect 9630 1280 9635 1300
rect 9605 1275 9635 1280
rect 9785 1300 9815 1305
rect 9785 1280 9790 1300
rect 9810 1280 9815 1300
rect 9785 1275 9815 1280
rect 9610 1140 9630 1275
rect 9790 1140 9810 1275
rect 9970 1140 9990 1315
rect 9425 1135 9455 1140
rect 9425 1115 9430 1135
rect 9450 1115 9455 1135
rect 9425 1110 9455 1115
rect 9605 1135 9635 1140
rect 9605 1115 9610 1135
rect 9630 1115 9635 1135
rect 9605 1110 9635 1115
rect 9785 1135 9815 1140
rect 9785 1115 9790 1135
rect 9810 1115 9815 1135
rect 9785 1110 9815 1115
rect 9965 1135 9995 1140
rect 9965 1115 9970 1135
rect 9990 1115 9995 1135
rect 9965 1110 9995 1115
rect 9430 1105 9450 1110
rect 9610 1105 9630 1110
rect 9790 1105 9810 1110
rect 9970 1105 9990 1110
rect 10105 1090 10125 1435
rect 10240 1430 10260 1435
rect 10420 1430 10440 1435
rect 10150 1345 10170 1350
rect 10145 1340 10175 1345
rect 10145 1320 10150 1340
rect 10170 1320 10175 1340
rect 10145 1315 10175 1320
rect 10150 1140 10170 1315
rect 10330 1305 10350 1310
rect 10325 1300 10355 1305
rect 10325 1280 10330 1300
rect 10350 1280 10355 1300
rect 10325 1275 10355 1280
rect 10330 1140 10350 1275
rect 10510 1140 10530 1555
rect 10555 1550 10575 1555
rect 10600 1425 10620 1640
rect 10595 1420 10625 1425
rect 10595 1400 10600 1420
rect 10620 1400 10625 1420
rect 10595 1395 10625 1400
rect 10600 1390 10620 1395
rect 10735 1225 10755 1690
rect 10825 1305 10845 1690
rect 10915 1345 10935 1690
rect 11005 1385 11025 1690
rect 11000 1380 11030 1385
rect 11000 1360 11005 1380
rect 11025 1360 11030 1380
rect 11000 1355 11030 1360
rect 10910 1340 10940 1345
rect 10910 1320 10915 1340
rect 10935 1320 10940 1340
rect 10910 1315 10940 1320
rect 10820 1300 10850 1305
rect 10820 1280 10825 1300
rect 10845 1280 10850 1300
rect 10820 1275 10850 1280
rect 10730 1220 10760 1225
rect 10730 1200 10735 1220
rect 10755 1200 10760 1220
rect 10730 1195 10760 1200
rect 10145 1135 10175 1140
rect 10145 1115 10150 1135
rect 10170 1115 10175 1135
rect 10145 1110 10175 1115
rect 10325 1135 10355 1140
rect 10325 1115 10330 1135
rect 10350 1115 10355 1135
rect 10325 1110 10355 1115
rect 10505 1135 10535 1140
rect 10505 1115 10510 1135
rect 10530 1115 10535 1135
rect 10505 1110 10535 1115
rect 10150 1105 10170 1110
rect 10330 1105 10350 1110
rect 10510 1105 10530 1110
rect 10735 1090 10755 1195
rect 10825 1090 10845 1275
rect 10915 1090 10935 1315
rect 11005 1090 11025 1355
rect 11095 1090 11115 1690
rect -345 1080 -315 1090
rect -345 1000 -340 1080
rect -320 1000 -315 1080
rect -345 990 -315 1000
rect -255 990 -225 1090
rect -165 990 -135 1090
rect -75 990 -45 1090
rect 15 990 45 1090
rect 105 990 135 1090
rect 195 1080 225 1090
rect 195 1000 200 1080
rect 220 1000 225 1080
rect 195 990 225 1000
rect 285 1080 315 1090
rect 285 1000 290 1080
rect 310 1000 315 1080
rect 285 990 315 1000
rect 375 1080 405 1090
rect 375 1000 380 1080
rect 400 1000 405 1080
rect 375 990 405 1000
rect 465 1080 495 1090
rect 465 1000 470 1080
rect 490 1000 495 1080
rect 465 990 495 1000
rect 555 1080 585 1090
rect 555 1000 560 1080
rect 580 1000 585 1080
rect 555 990 585 1000
rect 645 1080 675 1090
rect 645 1000 650 1080
rect 670 1000 675 1080
rect 645 990 675 1000
rect 735 1080 765 1090
rect 735 1000 740 1080
rect 760 1000 765 1080
rect 735 990 765 1000
rect 825 1080 855 1090
rect 825 1000 830 1080
rect 850 1000 855 1080
rect 825 990 855 1000
rect 915 1080 945 1090
rect 915 1000 920 1080
rect 940 1000 945 1080
rect 915 990 945 1000
rect 1005 1080 1035 1090
rect 1005 1000 1010 1080
rect 1030 1000 1035 1080
rect 1005 990 1035 1000
rect 1095 1080 1125 1090
rect 1095 1000 1100 1080
rect 1120 1000 1125 1080
rect 1095 990 1125 1000
rect 1185 1080 1215 1090
rect 1185 1000 1190 1080
rect 1210 1000 1215 1080
rect 1185 990 1215 1000
rect 1275 1080 1305 1090
rect 1275 1000 1280 1080
rect 1300 1000 1305 1080
rect 1275 990 1305 1000
rect 1365 1080 1395 1090
rect 1365 1000 1370 1080
rect 1390 1000 1395 1080
rect 1365 990 1395 1000
rect 1455 1080 1485 1090
rect 1455 1000 1460 1080
rect 1480 1000 1485 1080
rect 1455 990 1485 1000
rect 1545 1080 1575 1090
rect 1545 1000 1550 1080
rect 1570 1000 1575 1080
rect 1545 990 1575 1000
rect 1635 1080 1665 1090
rect 1635 1000 1640 1080
rect 1660 1000 1665 1080
rect 1635 990 1665 1000
rect 1725 1080 1755 1090
rect 1725 1000 1730 1080
rect 1750 1000 1755 1080
rect 1725 990 1755 1000
rect 1815 1080 1845 1090
rect 1815 1000 1820 1080
rect 1840 1000 1845 1080
rect 1815 990 1845 1000
rect 1905 1080 1935 1090
rect 1905 1000 1910 1080
rect 1930 1000 1935 1080
rect 1905 990 1935 1000
rect 1995 1080 2025 1090
rect 1995 1000 2000 1080
rect 2020 1000 2025 1080
rect 1995 990 2025 1000
rect 2085 1080 2115 1090
rect 2085 1000 2090 1080
rect 2110 1000 2115 1080
rect 2085 990 2115 1000
rect 2175 1080 2205 1090
rect 2175 1000 2180 1080
rect 2200 1000 2205 1080
rect 2175 990 2205 1000
rect 2265 1080 2295 1090
rect 2265 1000 2270 1080
rect 2290 1000 2295 1080
rect 2265 990 2295 1000
rect 2355 1080 2385 1090
rect 2355 1000 2360 1080
rect 2380 1000 2385 1080
rect 2355 990 2385 1000
rect 2445 1080 2475 1090
rect 2445 1000 2450 1080
rect 2470 1000 2475 1080
rect 2445 990 2475 1000
rect 2535 1080 2565 1090
rect 2535 1000 2540 1080
rect 2560 1000 2565 1080
rect 2535 990 2565 1000
rect 2625 1080 2655 1090
rect 2625 1000 2630 1080
rect 2650 1000 2655 1080
rect 2625 990 2655 1000
rect 2715 1080 2745 1090
rect 2715 1000 2720 1080
rect 2740 1000 2745 1080
rect 2715 990 2745 1000
rect 2805 1080 2835 1090
rect 2805 1000 2810 1080
rect 2830 1000 2835 1080
rect 2805 990 2835 1000
rect 2895 1080 2925 1090
rect 2895 1000 2900 1080
rect 2920 1000 2925 1080
rect 2895 990 2925 1000
rect 2985 1080 3015 1090
rect 2985 1000 2990 1080
rect 3010 1000 3015 1080
rect 2985 990 3015 1000
rect 3080 1080 3110 1090
rect 3080 1000 3085 1080
rect 3105 1000 3110 1080
rect 3080 990 3110 1000
rect 3170 1080 3200 1090
rect 3170 1000 3175 1080
rect 3195 1000 3200 1080
rect 3170 990 3200 1000
rect 3260 1080 3290 1090
rect 3260 1000 3265 1080
rect 3285 1000 3290 1080
rect 3260 990 3290 1000
rect 3350 1080 3380 1090
rect 3350 1000 3355 1080
rect 3375 1000 3380 1080
rect 3350 990 3380 1000
rect 3440 1080 3470 1090
rect 3440 1000 3445 1080
rect 3465 1000 3470 1080
rect 3440 990 3470 1000
rect 3530 1080 3560 1090
rect 3530 1000 3535 1080
rect 3555 1000 3560 1080
rect 3530 990 3560 1000
rect 3620 1080 3650 1090
rect 3620 1000 3625 1080
rect 3645 1000 3650 1080
rect 3620 990 3650 1000
rect 3710 1080 3740 1090
rect 3710 1000 3715 1080
rect 3735 1000 3740 1080
rect 3710 990 3740 1000
rect 3800 1080 3830 1090
rect 3800 1000 3805 1080
rect 3825 1000 3830 1080
rect 3800 990 3830 1000
rect 3890 1080 3920 1090
rect 3890 1000 3895 1080
rect 3915 1000 3920 1080
rect 3890 990 3920 1000
rect 3980 1080 4010 1090
rect 3980 1000 3985 1080
rect 4005 1000 4010 1080
rect 3980 990 4010 1000
rect 4070 1080 4100 1090
rect 4070 1000 4075 1080
rect 4095 1000 4100 1080
rect 4070 990 4100 1000
rect 4160 1080 4190 1090
rect 4160 1000 4165 1080
rect 4185 1000 4190 1080
rect 4160 990 4190 1000
rect 4250 1080 4280 1090
rect 4250 1000 4255 1080
rect 4275 1000 4280 1080
rect 4250 990 4280 1000
rect 4340 1080 4370 1090
rect 4340 1000 4345 1080
rect 4365 1000 4370 1080
rect 4340 990 4370 1000
rect 4430 1080 4460 1090
rect 4430 1000 4435 1080
rect 4455 1000 4460 1080
rect 4430 990 4460 1000
rect 4520 1080 4550 1090
rect 4520 1000 4525 1080
rect 4545 1000 4550 1080
rect 4520 990 4550 1000
rect 4610 1080 4640 1090
rect 4610 1000 4615 1080
rect 4635 1000 4640 1080
rect 4610 990 4640 1000
rect 4700 1080 4730 1090
rect 4700 1000 4705 1080
rect 4725 1000 4730 1080
rect 4700 990 4730 1000
rect 4790 1080 4820 1090
rect 4790 1000 4795 1080
rect 4815 1000 4820 1080
rect 4790 990 4820 1000
rect 4880 1080 4910 1090
rect 4880 1000 4885 1080
rect 4905 1000 4910 1080
rect 4880 990 4910 1000
rect 4970 1080 5000 1090
rect 4970 1000 4975 1080
rect 4995 1000 5000 1080
rect 4970 990 5000 1000
rect 5060 1080 5090 1090
rect 5060 1000 5065 1080
rect 5085 1000 5090 1080
rect 5060 990 5090 1000
rect 5150 1080 5180 1090
rect 5150 1000 5155 1080
rect 5175 1000 5180 1080
rect 5150 990 5180 1000
rect 5240 1080 5270 1090
rect 5240 1000 5245 1080
rect 5265 1000 5270 1080
rect 5240 990 5270 1000
rect 5330 1080 5360 1090
rect 5330 1000 5335 1080
rect 5355 1000 5360 1080
rect 5330 990 5360 1000
rect 5420 1080 5450 1090
rect 5420 1000 5425 1080
rect 5445 1000 5450 1080
rect 5420 990 5450 1000
rect 5510 1080 5540 1090
rect 5510 1000 5515 1080
rect 5535 1000 5540 1080
rect 5510 990 5540 1000
rect 5600 1080 5630 1090
rect 5600 1000 5605 1080
rect 5625 1000 5630 1080
rect 5600 990 5630 1000
rect 5690 1080 5720 1090
rect 5690 1000 5695 1080
rect 5715 1000 5720 1080
rect 5690 990 5720 1000
rect 5780 1080 5810 1090
rect 5780 1000 5785 1080
rect 5805 1000 5810 1080
rect 5780 990 5810 1000
rect 5870 1080 5900 1090
rect 5870 1000 5875 1080
rect 5895 1000 5900 1080
rect 5870 990 5900 1000
rect 5960 1080 5990 1090
rect 5960 1000 5965 1080
rect 5985 1000 5990 1080
rect 5960 990 5990 1000
rect 6050 1080 6080 1090
rect 6050 1000 6055 1080
rect 6075 1000 6080 1080
rect 6050 990 6080 1000
rect 6140 1080 6170 1090
rect 6140 1000 6145 1080
rect 6165 1000 6170 1080
rect 6140 990 6170 1000
rect 6230 1080 6260 1090
rect 6230 1000 6235 1080
rect 6255 1000 6260 1080
rect 6230 990 6260 1000
rect 6320 1080 6350 1090
rect 6320 1000 6325 1080
rect 6345 1000 6350 1080
rect 6320 990 6350 1000
rect 6410 1080 6440 1090
rect 6410 1000 6415 1080
rect 6435 1000 6440 1080
rect 6410 990 6440 1000
rect 6500 1080 6530 1090
rect 6500 1000 6505 1080
rect 6525 1000 6530 1080
rect 6500 990 6530 1000
rect 6590 1080 6620 1090
rect 6590 1000 6595 1080
rect 6615 1000 6620 1080
rect 6590 990 6620 1000
rect 6680 1080 6710 1090
rect 6680 1000 6685 1080
rect 6705 1000 6710 1080
rect 6680 990 6710 1000
rect 6770 1080 6800 1090
rect 6770 1000 6775 1080
rect 6795 1000 6800 1080
rect 6770 990 6800 1000
rect 6860 1080 6890 1090
rect 6860 1000 6865 1080
rect 6885 1000 6890 1080
rect 6860 990 6890 1000
rect 6950 1080 6980 1090
rect 6950 1000 6955 1080
rect 6975 1000 6980 1080
rect 6950 990 6980 1000
rect 7040 1080 7070 1090
rect 7040 1000 7045 1080
rect 7065 1000 7070 1080
rect 7040 990 7070 1000
rect 7130 1080 7160 1090
rect 7130 1000 7135 1080
rect 7155 1000 7160 1080
rect 7130 990 7160 1000
rect 7220 1080 7250 1090
rect 7220 1000 7225 1080
rect 7245 1000 7250 1080
rect 7220 990 7250 1000
rect 7310 1080 7340 1090
rect 7310 1000 7315 1080
rect 7335 1000 7340 1080
rect 7310 990 7340 1000
rect 7400 1080 7430 1090
rect 7400 1000 7405 1080
rect 7425 1000 7430 1080
rect 7400 990 7430 1000
rect 7490 1080 7520 1090
rect 7490 1000 7495 1080
rect 7515 1000 7520 1080
rect 7490 990 7520 1000
rect 7580 1080 7610 1090
rect 7580 1000 7585 1080
rect 7605 1000 7610 1080
rect 7580 990 7610 1000
rect 7670 1080 7700 1090
rect 7670 1000 7675 1080
rect 7695 1000 7700 1080
rect 7670 990 7700 1000
rect 7760 1080 7790 1090
rect 7760 1000 7765 1080
rect 7785 1000 7790 1080
rect 7760 990 7790 1000
rect 7850 1080 7880 1090
rect 7850 1000 7855 1080
rect 7875 1000 7880 1080
rect 7850 990 7880 1000
rect 7940 1080 7970 1090
rect 7940 1000 7945 1080
rect 7965 1000 7970 1080
rect 7940 990 7970 1000
rect 8030 1080 8060 1090
rect 8030 1000 8035 1080
rect 8055 1000 8060 1080
rect 8030 990 8060 1000
rect 8120 1080 8150 1090
rect 8120 1000 8125 1080
rect 8145 1000 8150 1080
rect 8120 990 8150 1000
rect 8210 1080 8240 1090
rect 8210 1000 8215 1080
rect 8235 1000 8240 1080
rect 8210 990 8240 1000
rect 8300 1080 8330 1090
rect 8300 1000 8305 1080
rect 8325 1000 8330 1080
rect 8300 990 8330 1000
rect 8390 1080 8420 1090
rect 8390 1000 8395 1080
rect 8415 1000 8420 1080
rect 8390 990 8420 1000
rect 8480 1080 8510 1090
rect 8480 1000 8485 1080
rect 8505 1000 8510 1080
rect 8480 990 8510 1000
rect 8570 1080 8600 1090
rect 8570 1000 8575 1080
rect 8595 1000 8600 1080
rect 8570 990 8600 1000
rect 8660 1080 8690 1090
rect 8660 1000 8665 1080
rect 8685 1000 8690 1080
rect 8660 990 8690 1000
rect 8750 1080 8780 1090
rect 8750 1000 8755 1080
rect 8775 1000 8780 1080
rect 8750 990 8780 1000
rect 8840 1080 8870 1090
rect 8840 1000 8845 1080
rect 8865 1000 8870 1080
rect 8840 990 8870 1000
rect 8930 1080 8960 1090
rect 8930 1000 8935 1080
rect 8955 1000 8960 1080
rect 8930 990 8960 1000
rect 9020 1080 9050 1090
rect 9020 1000 9025 1080
rect 9045 1000 9050 1080
rect 9020 990 9050 1000
rect 9110 1080 9140 1090
rect 9110 1000 9115 1080
rect 9135 1000 9140 1080
rect 9110 990 9140 1000
rect 9200 1080 9230 1090
rect 9200 1000 9205 1080
rect 9225 1000 9230 1080
rect 9200 990 9230 1000
rect 9290 1080 9320 1090
rect 9290 1000 9295 1080
rect 9315 1000 9320 1080
rect 9290 990 9320 1000
rect 9380 1080 9410 1090
rect 9380 1000 9385 1080
rect 9405 1000 9410 1080
rect 9380 990 9410 1000
rect 9470 1080 9500 1090
rect 9470 1000 9475 1080
rect 9495 1000 9500 1080
rect 9470 990 9500 1000
rect 9560 1080 9590 1090
rect 9560 1000 9565 1080
rect 9585 1000 9590 1080
rect 9560 990 9590 1000
rect 9650 1080 9680 1090
rect 9650 1000 9655 1080
rect 9675 1000 9680 1080
rect 9650 990 9680 1000
rect 9740 1080 9770 1090
rect 9740 1000 9745 1080
rect 9765 1000 9770 1080
rect 9740 990 9770 1000
rect 9830 1080 9860 1090
rect 9830 1000 9835 1080
rect 9855 1000 9860 1080
rect 9830 990 9860 1000
rect 9920 1080 9950 1090
rect 9920 1000 9925 1080
rect 9945 1000 9950 1080
rect 9920 990 9950 1000
rect 10010 1080 10040 1090
rect 10010 1000 10015 1080
rect 10035 1000 10040 1080
rect 10010 990 10040 1000
rect 10100 1080 10130 1090
rect 10100 1000 10105 1080
rect 10125 1000 10130 1080
rect 10100 990 10130 1000
rect 10190 1080 10220 1090
rect 10190 1000 10195 1080
rect 10215 1000 10220 1080
rect 10190 990 10220 1000
rect 10280 1080 10310 1090
rect 10280 1000 10285 1080
rect 10305 1000 10310 1080
rect 10280 990 10310 1000
rect 10370 1080 10400 1090
rect 10370 1000 10375 1080
rect 10395 1000 10400 1080
rect 10370 990 10400 1000
rect 10460 1080 10490 1090
rect 10460 1000 10465 1080
rect 10485 1000 10490 1080
rect 10460 990 10490 1000
rect 10550 1080 10580 1090
rect 10550 1000 10555 1080
rect 10575 1000 10580 1080
rect 10550 990 10580 1000
rect 10640 1080 10670 1090
rect 10640 1000 10645 1080
rect 10665 1000 10670 1080
rect 10640 990 10670 1000
rect 10730 990 10760 1090
rect 10820 990 10850 1090
rect 10910 990 10940 1090
rect 11000 990 11030 1090
rect 11090 990 11120 1090
rect 11180 1080 11210 1090
rect 11180 1000 11185 1080
rect 11205 1000 11210 1080
rect 11180 990 11210 1000
rect -340 970 -320 990
rect -350 965 -310 970
rect -350 935 -345 965
rect -315 935 -310 965
rect -350 930 -310 935
rect -350 905 -310 910
rect -350 875 -345 905
rect -315 875 -310 905
rect -350 870 -310 875
rect -340 850 -320 870
rect -250 850 -230 990
rect -160 850 -140 990
rect -70 850 -50 990
rect 20 850 40 990
rect 110 850 130 990
rect 200 970 220 990
rect 1640 970 1660 990
rect 3085 970 3105 990
rect 4525 970 4545 990
rect 5965 970 5985 990
rect 7585 970 7605 990
rect 9025 970 9045 990
rect 9745 970 9765 990
rect 10465 970 10485 990
rect 10645 970 10665 990
rect 190 965 230 970
rect 190 935 195 965
rect 225 935 230 965
rect 190 930 230 935
rect 370 965 410 970
rect 370 935 375 965
rect 405 935 410 965
rect 370 930 410 935
rect 550 965 590 970
rect 550 935 555 965
rect 585 935 590 965
rect 550 930 590 935
rect 730 965 770 970
rect 730 935 735 965
rect 765 935 770 965
rect 730 930 770 935
rect 910 965 950 970
rect 910 935 915 965
rect 945 935 950 965
rect 910 930 950 935
rect 1090 965 1130 970
rect 1090 935 1095 965
rect 1125 935 1130 965
rect 1090 930 1130 935
rect 1270 965 1310 970
rect 1270 935 1275 965
rect 1305 935 1310 965
rect 1270 930 1310 935
rect 1450 965 1490 970
rect 1450 935 1455 965
rect 1485 935 1490 965
rect 1450 930 1490 935
rect 1630 965 1670 970
rect 1630 935 1635 965
rect 1665 935 1670 965
rect 1630 930 1670 935
rect 1810 965 1850 970
rect 1810 935 1815 965
rect 1845 935 1850 965
rect 1810 930 1850 935
rect 1990 965 2030 970
rect 1990 935 1995 965
rect 2025 935 2030 965
rect 1990 930 2030 935
rect 2170 965 2210 970
rect 2170 935 2175 965
rect 2205 935 2210 965
rect 2170 930 2210 935
rect 2350 965 2390 970
rect 2350 935 2355 965
rect 2385 935 2390 965
rect 2350 930 2390 935
rect 2530 965 2570 970
rect 2530 935 2535 965
rect 2565 935 2570 965
rect 2530 930 2570 935
rect 2710 965 2750 970
rect 2710 935 2715 965
rect 2745 935 2750 965
rect 2710 930 2750 935
rect 2890 965 2930 970
rect 2890 935 2895 965
rect 2925 935 2930 965
rect 2890 930 2930 935
rect 3070 965 3115 970
rect 3070 935 3080 965
rect 3110 935 3115 965
rect 3070 930 3115 935
rect 3255 965 3295 970
rect 3255 935 3260 965
rect 3290 935 3295 965
rect 3255 930 3295 935
rect 3435 965 3475 970
rect 3435 935 3440 965
rect 3470 935 3475 965
rect 3435 930 3475 935
rect 3615 965 3655 970
rect 3615 935 3620 965
rect 3650 935 3655 965
rect 3615 930 3655 935
rect 3795 965 3835 970
rect 3795 935 3800 965
rect 3830 935 3835 965
rect 3795 930 3835 935
rect 3975 965 4015 970
rect 3975 935 3980 965
rect 4010 935 4015 965
rect 3975 930 4015 935
rect 4155 965 4195 970
rect 4155 935 4160 965
rect 4190 935 4195 965
rect 4155 930 4195 935
rect 4335 965 4375 970
rect 4335 935 4340 965
rect 4370 935 4375 965
rect 4335 930 4375 935
rect 4515 965 4555 970
rect 4515 935 4520 965
rect 4550 935 4555 965
rect 4515 930 4555 935
rect 4695 965 4735 970
rect 4695 935 4700 965
rect 4730 935 4735 965
rect 4695 930 4735 935
rect 4875 965 4915 970
rect 4875 935 4880 965
rect 4910 935 4915 965
rect 4875 930 4915 935
rect 5055 965 5095 970
rect 5055 935 5060 965
rect 5090 935 5095 965
rect 5055 930 5095 935
rect 5235 965 5275 970
rect 5235 935 5240 965
rect 5270 935 5275 965
rect 5235 930 5275 935
rect 5415 965 5455 970
rect 5415 935 5420 965
rect 5450 935 5455 965
rect 5415 930 5455 935
rect 5595 965 5635 970
rect 5595 935 5600 965
rect 5630 935 5635 965
rect 5595 930 5635 935
rect 5775 965 5815 970
rect 5775 935 5780 965
rect 5810 935 5815 965
rect 5775 930 5815 935
rect 5955 965 5995 970
rect 5955 935 5960 965
rect 5990 935 5995 965
rect 5955 930 5995 935
rect 6135 965 6175 970
rect 6135 935 6140 965
rect 6170 935 6175 965
rect 6135 930 6175 935
rect 6315 965 6355 970
rect 6315 935 6320 965
rect 6350 935 6355 965
rect 6315 930 6355 935
rect 6495 965 6535 970
rect 6495 935 6500 965
rect 6530 935 6535 965
rect 6495 930 6535 935
rect 6675 965 6715 970
rect 6675 935 6680 965
rect 6710 935 6715 965
rect 6675 930 6715 935
rect 6855 965 6895 970
rect 6855 935 6860 965
rect 6890 935 6895 965
rect 6855 930 6895 935
rect 7035 965 7075 970
rect 7035 935 7040 965
rect 7070 935 7075 965
rect 7035 930 7075 935
rect 7215 965 7255 970
rect 7215 935 7220 965
rect 7250 935 7255 965
rect 7215 930 7255 935
rect 7395 965 7435 970
rect 7395 935 7400 965
rect 7430 935 7435 965
rect 7395 930 7435 935
rect 7575 965 7615 970
rect 7575 935 7580 965
rect 7610 935 7615 965
rect 7575 930 7615 935
rect 7755 965 7795 970
rect 7755 935 7760 965
rect 7790 935 7795 965
rect 7755 930 7795 935
rect 7935 965 7975 970
rect 7935 935 7940 965
rect 7970 935 7975 965
rect 7935 930 7975 935
rect 8115 965 8155 970
rect 8115 935 8120 965
rect 8150 935 8155 965
rect 8115 930 8155 935
rect 8295 965 8335 970
rect 8295 935 8300 965
rect 8330 935 8335 965
rect 8295 930 8335 935
rect 8475 965 8515 970
rect 8475 935 8480 965
rect 8510 935 8515 965
rect 8475 930 8515 935
rect 8655 965 8695 970
rect 8655 935 8660 965
rect 8690 935 8695 965
rect 8655 930 8695 935
rect 8835 965 8875 970
rect 8835 935 8840 965
rect 8870 935 8875 965
rect 8835 930 8875 935
rect 9015 965 9055 970
rect 9015 935 9020 965
rect 9050 935 9055 965
rect 9015 930 9055 935
rect 9195 965 9235 970
rect 9195 935 9200 965
rect 9230 935 9235 965
rect 9195 930 9235 935
rect 9375 965 9415 970
rect 9375 935 9380 965
rect 9410 935 9415 965
rect 9375 930 9415 935
rect 9555 965 9595 970
rect 9555 935 9560 965
rect 9590 935 9595 965
rect 9555 930 9595 935
rect 9735 965 9775 970
rect 9735 935 9740 965
rect 9770 935 9775 965
rect 9735 930 9775 935
rect 9915 965 9955 970
rect 9915 935 9920 965
rect 9950 935 9955 965
rect 9915 930 9955 935
rect 10095 965 10135 970
rect 10095 935 10100 965
rect 10130 935 10135 965
rect 10095 930 10135 935
rect 10275 965 10315 970
rect 10275 935 10280 965
rect 10310 935 10315 965
rect 10275 930 10315 935
rect 10455 965 10495 970
rect 10455 935 10460 965
rect 10490 935 10495 965
rect 10455 930 10495 935
rect 10635 965 10675 970
rect 10635 935 10640 965
rect 10670 935 10675 965
rect 10635 930 10675 935
rect 190 905 230 910
rect 190 875 195 905
rect 225 875 230 905
rect 190 870 230 875
rect 370 905 410 910
rect 370 875 375 905
rect 405 875 410 905
rect 370 870 410 875
rect 550 905 590 910
rect 550 875 555 905
rect 585 875 590 905
rect 550 870 590 875
rect 730 905 770 910
rect 730 875 735 905
rect 765 875 770 905
rect 730 870 770 875
rect 910 905 950 910
rect 910 875 915 905
rect 945 875 950 905
rect 910 870 950 875
rect 1090 905 1130 910
rect 1090 875 1095 905
rect 1125 875 1130 905
rect 1090 870 1130 875
rect 1270 905 1310 910
rect 1270 875 1275 905
rect 1305 875 1310 905
rect 1270 870 1310 875
rect 1450 905 1490 910
rect 1450 875 1455 905
rect 1485 875 1490 905
rect 1450 870 1490 875
rect 1630 905 1670 910
rect 1630 875 1635 905
rect 1665 875 1670 905
rect 1630 870 1670 875
rect 1810 905 1850 910
rect 1810 875 1815 905
rect 1845 875 1850 905
rect 1810 870 1850 875
rect 1990 905 2030 910
rect 1990 875 1995 905
rect 2025 875 2030 905
rect 1990 870 2030 875
rect 2170 905 2210 910
rect 2170 875 2175 905
rect 2205 875 2210 905
rect 2170 870 2210 875
rect 2350 905 2390 910
rect 2350 875 2355 905
rect 2385 875 2390 905
rect 2350 870 2390 875
rect 2530 905 2570 910
rect 2530 875 2535 905
rect 2565 875 2570 905
rect 2530 870 2570 875
rect 2710 905 2750 910
rect 2710 875 2715 905
rect 2745 875 2750 905
rect 2710 870 2750 875
rect 2890 905 2930 910
rect 2890 875 2895 905
rect 2925 875 2930 905
rect 2890 870 2930 875
rect 3070 905 3110 910
rect 3070 875 3075 905
rect 3105 875 3110 905
rect 3070 870 3110 875
rect 3250 905 3290 910
rect 3250 875 3255 905
rect 3285 875 3290 905
rect 3250 870 3290 875
rect 3430 905 3470 910
rect 3430 875 3435 905
rect 3465 875 3470 905
rect 3430 870 3470 875
rect 3610 905 3650 910
rect 3610 875 3615 905
rect 3645 875 3650 905
rect 3610 870 3650 875
rect 3790 905 3830 910
rect 3790 875 3795 905
rect 3825 875 3830 905
rect 3790 870 3830 875
rect 3970 905 4010 910
rect 3970 875 3975 905
rect 4005 875 4010 905
rect 3970 870 4010 875
rect 4150 905 4190 910
rect 4150 875 4155 905
rect 4185 875 4190 905
rect 4150 870 4190 875
rect 4330 905 4370 910
rect 4330 875 4335 905
rect 4365 875 4370 905
rect 4330 870 4370 875
rect 4510 905 4550 910
rect 4510 875 4515 905
rect 4545 875 4550 905
rect 4510 870 4550 875
rect 4690 905 4730 910
rect 4690 875 4695 905
rect 4725 875 4730 905
rect 4690 870 4730 875
rect 4870 905 4910 910
rect 4870 875 4875 905
rect 4905 875 4910 905
rect 4870 870 4910 875
rect 5050 905 5090 910
rect 5050 875 5055 905
rect 5085 875 5090 905
rect 5050 870 5090 875
rect 5230 905 5270 910
rect 5230 875 5235 905
rect 5265 875 5270 905
rect 5230 870 5270 875
rect 5410 905 5450 910
rect 5410 875 5415 905
rect 5445 875 5450 905
rect 5410 870 5450 875
rect 5590 905 5630 910
rect 5590 875 5595 905
rect 5625 875 5630 905
rect 5590 870 5630 875
rect 5770 905 5810 910
rect 5770 875 5775 905
rect 5805 875 5810 905
rect 5770 870 5810 875
rect 5950 905 5990 910
rect 5950 875 5955 905
rect 5985 875 5990 905
rect 5950 870 5990 875
rect 6130 905 6170 910
rect 6130 875 6135 905
rect 6165 875 6170 905
rect 6130 870 6170 875
rect 6310 905 6350 910
rect 6310 875 6315 905
rect 6345 875 6350 905
rect 6310 870 6350 875
rect 6490 905 6530 910
rect 6490 875 6495 905
rect 6525 875 6530 905
rect 6490 870 6530 875
rect 6670 905 6710 910
rect 6670 875 6675 905
rect 6705 875 6710 905
rect 6670 870 6710 875
rect 6850 905 6890 910
rect 6850 875 6855 905
rect 6885 875 6890 905
rect 6850 870 6890 875
rect 7030 905 7070 910
rect 7030 875 7035 905
rect 7065 875 7070 905
rect 7030 870 7070 875
rect 7210 905 7250 910
rect 7210 875 7215 905
rect 7245 875 7250 905
rect 7210 870 7250 875
rect 7390 905 7430 910
rect 7390 875 7395 905
rect 7425 875 7430 905
rect 7390 870 7430 875
rect 7570 905 7610 910
rect 7570 875 7575 905
rect 7605 875 7610 905
rect 7570 870 7610 875
rect 7750 905 7795 910
rect 7750 875 7755 905
rect 7785 875 7795 905
rect 7750 870 7795 875
rect 7935 905 7975 910
rect 7935 875 7940 905
rect 7970 875 7975 905
rect 7935 870 7975 875
rect 8115 905 8155 910
rect 8115 875 8120 905
rect 8150 875 8155 905
rect 8115 870 8155 875
rect 8295 905 8335 910
rect 8295 875 8300 905
rect 8330 875 8335 905
rect 8295 870 8335 875
rect 8475 905 8515 910
rect 8475 875 8480 905
rect 8510 875 8515 905
rect 8475 870 8515 875
rect 8655 905 8695 910
rect 8655 875 8660 905
rect 8690 875 8695 905
rect 8655 870 8695 875
rect 8835 905 8875 910
rect 8835 875 8840 905
rect 8870 875 8875 905
rect 8835 870 8875 875
rect 9015 905 9055 910
rect 9015 875 9020 905
rect 9050 875 9055 905
rect 9015 870 9055 875
rect 9195 905 9235 910
rect 9195 875 9200 905
rect 9230 875 9235 905
rect 9195 870 9235 875
rect 9375 905 9415 910
rect 9375 875 9380 905
rect 9410 875 9415 905
rect 9375 870 9415 875
rect 9555 905 9595 910
rect 9555 875 9560 905
rect 9590 875 9595 905
rect 9555 870 9595 875
rect 9735 905 9775 910
rect 9735 875 9740 905
rect 9770 875 9775 905
rect 9735 870 9775 875
rect 9915 905 9955 910
rect 9915 875 9920 905
rect 9950 875 9955 905
rect 9915 870 9955 875
rect 10095 905 10135 910
rect 10095 875 10100 905
rect 10130 875 10135 905
rect 10095 870 10135 875
rect 10275 905 10315 910
rect 10275 875 10280 905
rect 10310 875 10315 905
rect 10275 870 10315 875
rect 10455 905 10495 910
rect 10455 875 10460 905
rect 10490 875 10495 905
rect 10455 870 10495 875
rect 10635 905 10675 910
rect 10635 875 10640 905
rect 10670 875 10675 905
rect 10635 870 10675 875
rect 200 850 220 870
rect 380 850 400 870
rect 1100 850 1120 870
rect 1820 850 1840 870
rect 3260 850 3280 870
rect 4880 850 4900 870
rect 6320 850 6340 870
rect 7760 850 7780 870
rect 9205 850 9225 870
rect 10645 850 10665 870
rect 10735 850 10755 990
rect 10825 850 10845 990
rect 10915 850 10935 990
rect 11005 850 11025 990
rect 11095 850 11115 990
rect 11185 970 11205 990
rect 11175 965 11215 970
rect 11175 935 11180 965
rect 11210 935 11215 965
rect 11175 930 11215 935
rect 11175 905 11215 910
rect 11175 875 11180 905
rect 11210 875 11215 905
rect 11175 870 11215 875
rect 11185 850 11205 870
rect -345 840 -315 850
rect -345 760 -340 840
rect -320 760 -315 840
rect -345 750 -315 760
rect -255 750 -225 850
rect -165 750 -135 850
rect -75 750 -45 850
rect 15 750 45 850
rect 105 750 135 850
rect 195 840 225 850
rect 195 760 200 840
rect 220 760 225 840
rect 195 750 225 760
rect 285 840 315 850
rect 285 760 290 840
rect 310 760 315 840
rect 285 750 315 760
rect 375 840 405 850
rect 375 760 380 840
rect 400 760 405 840
rect 375 750 405 760
rect 465 840 495 850
rect 465 760 470 840
rect 490 760 495 840
rect 465 750 495 760
rect 555 840 585 850
rect 555 760 560 840
rect 580 760 585 840
rect 555 750 585 760
rect 645 840 675 850
rect 645 760 650 840
rect 670 760 675 840
rect 645 750 675 760
rect 735 840 765 850
rect 735 760 740 840
rect 760 760 765 840
rect 735 750 765 760
rect 825 840 855 850
rect 825 760 830 840
rect 850 760 855 840
rect 825 750 855 760
rect 915 840 945 850
rect 915 760 920 840
rect 940 760 945 840
rect 915 750 945 760
rect 1005 840 1035 850
rect 1005 760 1010 840
rect 1030 760 1035 840
rect 1005 750 1035 760
rect 1095 840 1125 850
rect 1095 760 1100 840
rect 1120 760 1125 840
rect 1095 750 1125 760
rect 1185 840 1215 850
rect 1185 760 1190 840
rect 1210 760 1215 840
rect 1185 750 1215 760
rect 1275 840 1305 850
rect 1275 760 1280 840
rect 1300 760 1305 840
rect 1275 750 1305 760
rect 1365 840 1395 850
rect 1365 760 1370 840
rect 1390 760 1395 840
rect 1365 750 1395 760
rect 1455 840 1485 850
rect 1455 760 1460 840
rect 1480 760 1485 840
rect 1455 750 1485 760
rect 1545 840 1575 850
rect 1545 760 1550 840
rect 1570 760 1575 840
rect 1545 750 1575 760
rect 1635 840 1665 850
rect 1635 760 1640 840
rect 1660 760 1665 840
rect 1635 750 1665 760
rect 1725 840 1755 850
rect 1725 760 1730 840
rect 1750 760 1755 840
rect 1725 750 1755 760
rect 1815 840 1845 850
rect 1815 760 1820 840
rect 1840 760 1845 840
rect 1815 750 1845 760
rect 1905 840 1935 850
rect 1905 760 1910 840
rect 1930 760 1935 840
rect 1905 750 1935 760
rect 1995 840 2025 850
rect 1995 760 2000 840
rect 2020 760 2025 840
rect 1995 750 2025 760
rect 2085 840 2115 850
rect 2085 760 2090 840
rect 2110 760 2115 840
rect 2085 750 2115 760
rect 2175 840 2205 850
rect 2175 760 2180 840
rect 2200 760 2205 840
rect 2175 750 2205 760
rect 2265 840 2295 850
rect 2265 760 2270 840
rect 2290 760 2295 840
rect 2265 750 2295 760
rect 2355 840 2385 850
rect 2355 760 2360 840
rect 2380 760 2385 840
rect 2355 750 2385 760
rect 2445 840 2475 850
rect 2445 760 2450 840
rect 2470 760 2475 840
rect 2445 750 2475 760
rect 2535 840 2565 850
rect 2535 760 2540 840
rect 2560 760 2565 840
rect 2535 750 2565 760
rect 2625 840 2655 850
rect 2625 760 2630 840
rect 2650 760 2655 840
rect 2625 750 2655 760
rect 2715 840 2745 850
rect 2715 760 2720 840
rect 2740 760 2745 840
rect 2715 750 2745 760
rect 2805 840 2835 850
rect 2805 760 2810 840
rect 2830 760 2835 840
rect 2805 750 2835 760
rect 2895 840 2925 850
rect 2895 760 2900 840
rect 2920 760 2925 840
rect 2895 750 2925 760
rect 2985 840 3015 850
rect 2985 760 2990 840
rect 3010 760 3015 840
rect 2985 750 3015 760
rect 3075 840 3105 850
rect 3075 760 3080 840
rect 3100 760 3105 840
rect 3075 750 3105 760
rect 3165 840 3195 850
rect 3165 760 3170 840
rect 3190 760 3195 840
rect 3165 750 3195 760
rect 3255 840 3285 850
rect 3255 760 3260 840
rect 3280 760 3285 840
rect 3255 750 3285 760
rect 3345 840 3375 850
rect 3345 760 3350 840
rect 3370 760 3375 840
rect 3345 750 3375 760
rect 3435 840 3465 850
rect 3435 760 3440 840
rect 3460 760 3465 840
rect 3435 750 3465 760
rect 3525 840 3555 850
rect 3525 760 3530 840
rect 3550 760 3555 840
rect 3525 750 3555 760
rect 3615 840 3645 850
rect 3615 760 3620 840
rect 3640 760 3645 840
rect 3615 750 3645 760
rect 3705 840 3735 850
rect 3705 760 3710 840
rect 3730 760 3735 840
rect 3705 750 3735 760
rect 3795 840 3825 850
rect 3795 760 3800 840
rect 3820 760 3825 840
rect 3795 750 3825 760
rect 3885 840 3915 850
rect 3885 760 3890 840
rect 3910 760 3915 840
rect 3885 750 3915 760
rect 3975 840 4005 850
rect 3975 760 3980 840
rect 4000 760 4005 840
rect 3975 750 4005 760
rect 4065 840 4095 850
rect 4065 760 4070 840
rect 4090 760 4095 840
rect 4065 750 4095 760
rect 4155 840 4185 850
rect 4155 760 4160 840
rect 4180 760 4185 840
rect 4155 750 4185 760
rect 4245 840 4275 850
rect 4245 760 4250 840
rect 4270 760 4275 840
rect 4245 750 4275 760
rect 4335 840 4365 850
rect 4335 760 4340 840
rect 4360 760 4365 840
rect 4335 750 4365 760
rect 4425 840 4455 850
rect 4425 760 4430 840
rect 4450 760 4455 840
rect 4425 750 4455 760
rect 4515 840 4545 850
rect 4515 760 4520 840
rect 4540 760 4545 840
rect 4515 750 4545 760
rect 4605 840 4635 850
rect 4605 760 4610 840
rect 4630 760 4635 840
rect 4605 750 4635 760
rect 4695 840 4725 850
rect 4695 760 4700 840
rect 4720 760 4725 840
rect 4695 750 4725 760
rect 4785 840 4815 850
rect 4785 760 4790 840
rect 4810 760 4815 840
rect 4785 750 4815 760
rect 4875 840 4905 850
rect 4875 760 4880 840
rect 4900 760 4905 840
rect 4875 750 4905 760
rect 4965 840 4995 850
rect 4965 760 4970 840
rect 4990 760 4995 840
rect 4965 750 4995 760
rect 5055 840 5085 850
rect 5055 760 5060 840
rect 5080 760 5085 840
rect 5055 750 5085 760
rect 5145 840 5175 850
rect 5145 760 5150 840
rect 5170 760 5175 840
rect 5145 750 5175 760
rect 5235 840 5265 850
rect 5235 760 5240 840
rect 5260 760 5265 840
rect 5235 750 5265 760
rect 5325 840 5355 850
rect 5325 760 5330 840
rect 5350 760 5355 840
rect 5325 750 5355 760
rect 5415 840 5445 850
rect 5415 760 5420 840
rect 5440 760 5445 840
rect 5415 750 5445 760
rect 5505 840 5535 850
rect 5505 760 5510 840
rect 5530 760 5535 840
rect 5505 750 5535 760
rect 5595 840 5625 850
rect 5595 760 5600 840
rect 5620 760 5625 840
rect 5595 750 5625 760
rect 5685 840 5715 850
rect 5685 760 5690 840
rect 5710 760 5715 840
rect 5685 750 5715 760
rect 5775 840 5805 850
rect 5775 760 5780 840
rect 5800 760 5805 840
rect 5775 750 5805 760
rect 5865 840 5895 850
rect 5865 760 5870 840
rect 5890 760 5895 840
rect 5865 750 5895 760
rect 5955 840 5985 850
rect 5955 760 5960 840
rect 5980 760 5985 840
rect 5955 750 5985 760
rect 6045 840 6075 850
rect 6045 760 6050 840
rect 6070 760 6075 840
rect 6045 750 6075 760
rect 6135 840 6165 850
rect 6135 760 6140 840
rect 6160 760 6165 840
rect 6135 750 6165 760
rect 6225 840 6255 850
rect 6225 760 6230 840
rect 6250 760 6255 840
rect 6225 750 6255 760
rect 6315 840 6345 850
rect 6315 760 6320 840
rect 6340 760 6345 840
rect 6315 750 6345 760
rect 6405 840 6435 850
rect 6405 760 6410 840
rect 6430 760 6435 840
rect 6405 750 6435 760
rect 6495 840 6525 850
rect 6495 760 6500 840
rect 6520 760 6525 840
rect 6495 750 6525 760
rect 6585 840 6615 850
rect 6585 760 6590 840
rect 6610 760 6615 840
rect 6585 750 6615 760
rect 6675 840 6705 850
rect 6675 760 6680 840
rect 6700 760 6705 840
rect 6675 750 6705 760
rect 6765 840 6795 850
rect 6765 760 6770 840
rect 6790 760 6795 840
rect 6765 750 6795 760
rect 6855 840 6885 850
rect 6855 760 6860 840
rect 6880 760 6885 840
rect 6855 750 6885 760
rect 6945 840 6975 850
rect 6945 760 6950 840
rect 6970 760 6975 840
rect 6945 750 6975 760
rect 7035 840 7065 850
rect 7035 760 7040 840
rect 7060 760 7065 840
rect 7035 750 7065 760
rect 7125 840 7155 850
rect 7125 760 7130 840
rect 7150 760 7155 840
rect 7125 750 7155 760
rect 7215 840 7245 850
rect 7215 760 7220 840
rect 7240 760 7245 840
rect 7215 750 7245 760
rect 7305 840 7335 850
rect 7305 760 7310 840
rect 7330 760 7335 840
rect 7305 750 7335 760
rect 7395 840 7425 850
rect 7395 760 7400 840
rect 7420 760 7425 840
rect 7395 750 7425 760
rect 7485 840 7515 850
rect 7485 760 7490 840
rect 7510 760 7515 840
rect 7485 750 7515 760
rect 7575 840 7605 850
rect 7575 760 7580 840
rect 7600 760 7605 840
rect 7575 750 7605 760
rect 7665 840 7695 850
rect 7665 760 7670 840
rect 7690 760 7695 840
rect 7665 750 7695 760
rect 7755 840 7785 850
rect 7755 760 7760 840
rect 7780 760 7785 840
rect 7755 750 7785 760
rect 7850 840 7880 850
rect 7850 760 7855 840
rect 7875 760 7880 840
rect 7850 750 7880 760
rect 7940 840 7970 850
rect 7940 760 7945 840
rect 7965 760 7970 840
rect 7940 750 7970 760
rect 8030 840 8060 850
rect 8030 760 8035 840
rect 8055 760 8060 840
rect 8030 750 8060 760
rect 8120 840 8150 850
rect 8120 760 8125 840
rect 8145 760 8150 840
rect 8120 750 8150 760
rect 8210 840 8240 850
rect 8210 760 8215 840
rect 8235 760 8240 840
rect 8210 750 8240 760
rect 8300 840 8330 850
rect 8300 760 8305 840
rect 8325 760 8330 840
rect 8300 750 8330 760
rect 8390 840 8420 850
rect 8390 760 8395 840
rect 8415 760 8420 840
rect 8390 750 8420 760
rect 8480 840 8510 850
rect 8480 760 8485 840
rect 8505 760 8510 840
rect 8480 750 8510 760
rect 8570 840 8600 850
rect 8570 760 8575 840
rect 8595 760 8600 840
rect 8570 750 8600 760
rect 8660 840 8690 850
rect 8660 760 8665 840
rect 8685 760 8690 840
rect 8660 750 8690 760
rect 8750 840 8780 850
rect 8750 760 8755 840
rect 8775 760 8780 840
rect 8750 750 8780 760
rect 8840 840 8870 850
rect 8840 760 8845 840
rect 8865 760 8870 840
rect 8840 750 8870 760
rect 8930 840 8960 850
rect 8930 760 8935 840
rect 8955 760 8960 840
rect 8930 750 8960 760
rect 9020 840 9050 850
rect 9020 760 9025 840
rect 9045 760 9050 840
rect 9020 750 9050 760
rect 9110 840 9140 850
rect 9110 760 9115 840
rect 9135 760 9140 840
rect 9110 750 9140 760
rect 9200 840 9230 850
rect 9200 760 9205 840
rect 9225 760 9230 840
rect 9200 750 9230 760
rect 9290 840 9320 850
rect 9290 760 9295 840
rect 9315 760 9320 840
rect 9290 750 9320 760
rect 9380 840 9410 850
rect 9380 760 9385 840
rect 9405 760 9410 840
rect 9380 750 9410 760
rect 9470 840 9500 850
rect 9470 760 9475 840
rect 9495 760 9500 840
rect 9470 750 9500 760
rect 9560 840 9590 850
rect 9560 760 9565 840
rect 9585 760 9590 840
rect 9560 750 9590 760
rect 9650 840 9680 850
rect 9650 760 9655 840
rect 9675 760 9680 840
rect 9650 750 9680 760
rect 9740 840 9770 850
rect 9740 760 9745 840
rect 9765 760 9770 840
rect 9740 750 9770 760
rect 9830 840 9860 850
rect 9830 760 9835 840
rect 9855 760 9860 840
rect 9830 750 9860 760
rect 9920 840 9950 850
rect 9920 760 9925 840
rect 9945 760 9950 840
rect 9920 750 9950 760
rect 10010 840 10040 850
rect 10010 760 10015 840
rect 10035 760 10040 840
rect 10010 750 10040 760
rect 10100 840 10130 850
rect 10100 760 10105 840
rect 10125 760 10130 840
rect 10100 750 10130 760
rect 10190 840 10220 850
rect 10190 760 10195 840
rect 10215 760 10220 840
rect 10190 750 10220 760
rect 10280 840 10310 850
rect 10280 760 10285 840
rect 10305 760 10310 840
rect 10280 750 10310 760
rect 10370 840 10400 850
rect 10370 760 10375 840
rect 10395 760 10400 840
rect 10370 750 10400 760
rect 10460 840 10490 850
rect 10460 760 10465 840
rect 10485 760 10490 840
rect 10460 750 10490 760
rect 10550 840 10580 850
rect 10550 760 10555 840
rect 10575 760 10580 840
rect 10550 750 10580 760
rect 10640 840 10670 850
rect 10640 760 10645 840
rect 10665 760 10670 840
rect 10640 750 10670 760
rect 10730 750 10760 850
rect 10820 750 10850 850
rect 10910 750 10940 850
rect 11000 750 11030 850
rect 11090 750 11120 850
rect 11180 840 11210 850
rect 11180 760 11185 840
rect 11205 760 11210 840
rect 11180 750 11210 760
rect -250 445 -230 750
rect -255 440 -225 445
rect -255 420 -250 440
rect -230 420 -225 440
rect -255 415 -225 420
rect -250 150 -230 415
rect -160 405 -140 750
rect -165 400 -135 405
rect -165 380 -160 400
rect -140 380 -135 400
rect -165 375 -135 380
rect -160 150 -140 375
rect -70 365 -50 750
rect -75 360 -45 365
rect -75 340 -70 360
rect -50 340 -45 360
rect -75 335 -45 340
rect -70 150 -50 335
rect 20 325 40 750
rect 15 320 45 325
rect 15 300 20 320
rect 40 300 45 320
rect 15 295 45 300
rect 20 150 40 295
rect 110 285 130 750
rect 335 730 355 735
rect 515 730 535 735
rect 695 730 715 735
rect 330 725 360 730
rect 330 705 335 725
rect 355 705 360 725
rect 330 700 360 705
rect 510 725 540 730
rect 510 705 515 725
rect 535 705 540 725
rect 510 700 540 705
rect 690 725 720 730
rect 690 705 695 725
rect 715 705 720 725
rect 690 700 720 705
rect 245 445 265 450
rect 240 440 270 445
rect 240 420 245 440
rect 265 420 270 440
rect 240 415 270 420
rect 105 280 135 285
rect 105 260 110 280
rect 130 260 135 280
rect 105 255 135 260
rect 110 150 130 255
rect 245 200 265 415
rect 290 285 310 290
rect 335 285 355 700
rect 515 565 535 700
rect 510 560 540 565
rect 510 540 515 560
rect 535 540 540 560
rect 510 535 540 540
rect 515 530 535 535
rect 695 525 715 700
rect 690 520 720 525
rect 690 500 695 520
rect 715 500 720 520
rect 690 495 720 500
rect 695 490 715 495
rect 425 405 445 410
rect 605 405 625 410
rect 740 405 760 750
rect 875 730 895 735
rect 1055 730 1075 735
rect 1235 730 1255 735
rect 1415 730 1435 735
rect 870 725 900 730
rect 870 705 875 725
rect 895 705 900 725
rect 870 700 900 705
rect 1050 725 1080 730
rect 1050 705 1055 725
rect 1075 705 1080 725
rect 1050 700 1080 705
rect 1230 725 1260 730
rect 1230 705 1235 725
rect 1255 705 1260 725
rect 1230 700 1260 705
rect 1410 725 1440 730
rect 1410 705 1415 725
rect 1435 705 1440 725
rect 1410 700 1440 705
rect 875 525 895 700
rect 1055 565 1075 700
rect 1235 565 1255 700
rect 1050 560 1080 565
rect 1050 540 1055 560
rect 1075 540 1080 560
rect 1050 535 1080 540
rect 1230 560 1260 565
rect 1230 540 1235 560
rect 1255 540 1260 560
rect 1230 535 1260 540
rect 1055 530 1075 535
rect 1235 530 1255 535
rect 1415 525 1435 700
rect 870 520 900 525
rect 870 500 875 520
rect 895 500 900 520
rect 870 495 900 500
rect 1410 520 1440 525
rect 1410 500 1415 520
rect 1435 500 1440 520
rect 1410 495 1440 500
rect 875 490 895 495
rect 1415 490 1435 495
rect 785 405 805 410
rect 965 405 985 410
rect 1100 405 1120 410
rect 1145 405 1165 410
rect 1325 405 1345 410
rect 1460 405 1480 750
rect 1595 730 1615 735
rect 1775 730 1795 735
rect 1955 730 1975 735
rect 2135 730 2155 735
rect 2315 730 2335 735
rect 2495 730 2515 735
rect 1590 725 1620 730
rect 1590 705 1595 725
rect 1615 705 1620 725
rect 1590 700 1620 705
rect 1770 725 1800 730
rect 1770 705 1775 725
rect 1795 705 1800 725
rect 1770 700 1800 705
rect 1950 725 1980 730
rect 1950 705 1955 725
rect 1975 705 1980 725
rect 1950 700 1980 705
rect 2130 725 2160 730
rect 2130 705 2135 725
rect 2155 705 2160 725
rect 2130 700 2160 705
rect 2310 725 2340 730
rect 2310 705 2315 725
rect 2335 705 2340 725
rect 2310 700 2340 705
rect 2490 725 2520 730
rect 2490 705 2495 725
rect 2515 705 2520 725
rect 2490 700 2520 705
rect 1595 525 1615 700
rect 1775 565 1795 700
rect 1955 565 1975 700
rect 2135 565 2155 700
rect 1770 560 1800 565
rect 1770 540 1775 560
rect 1795 540 1800 560
rect 1770 535 1800 540
rect 1950 560 1980 565
rect 1950 540 1955 560
rect 1975 540 1980 560
rect 1950 535 1980 540
rect 2130 560 2160 565
rect 2130 540 2135 560
rect 2155 540 2160 560
rect 2130 535 2160 540
rect 1775 530 1795 535
rect 1955 530 1975 535
rect 2135 530 2155 535
rect 2315 525 2335 700
rect 2495 525 2515 700
rect 1590 520 1620 525
rect 1590 500 1595 520
rect 1615 500 1620 520
rect 1590 495 1620 500
rect 2310 520 2340 525
rect 2310 500 2315 520
rect 2335 500 2340 520
rect 2310 495 2340 500
rect 2490 520 2520 525
rect 2490 500 2495 520
rect 2515 500 2520 520
rect 2490 495 2520 500
rect 1595 490 1615 495
rect 2315 490 2335 495
rect 2495 490 2515 495
rect 1505 405 1525 410
rect 1685 405 1705 410
rect 1865 405 1885 410
rect 2045 405 2065 410
rect 420 400 450 405
rect 420 380 425 400
rect 445 380 450 400
rect 420 375 450 380
rect 600 400 630 405
rect 600 380 605 400
rect 625 380 630 400
rect 600 375 630 380
rect 735 400 765 405
rect 735 380 740 400
rect 760 380 765 400
rect 735 375 765 380
rect 780 400 810 405
rect 780 380 785 400
rect 805 380 810 400
rect 780 375 810 380
rect 960 400 990 405
rect 960 380 965 400
rect 985 380 990 400
rect 960 375 990 380
rect 1095 400 1125 405
rect 1095 380 1100 400
rect 1120 380 1125 400
rect 1095 375 1125 380
rect 1140 400 1170 405
rect 1140 380 1145 400
rect 1165 380 1170 400
rect 1140 375 1170 380
rect 1320 400 1350 405
rect 1320 380 1325 400
rect 1345 380 1350 400
rect 1320 375 1350 380
rect 1455 400 1485 405
rect 1455 380 1460 400
rect 1480 380 1485 400
rect 1455 375 1485 380
rect 1500 400 1530 405
rect 1500 380 1505 400
rect 1525 380 1530 400
rect 1500 375 1530 380
rect 1680 400 1710 405
rect 1680 380 1685 400
rect 1705 380 1710 400
rect 1680 375 1710 380
rect 1860 400 1890 405
rect 1860 380 1865 400
rect 1885 380 1890 400
rect 1860 375 1890 380
rect 2040 400 2070 405
rect 2040 380 2045 400
rect 2065 380 2070 400
rect 2040 375 2070 380
rect 285 280 315 285
rect 285 260 290 280
rect 310 260 315 280
rect 285 255 315 260
rect 330 280 360 285
rect 330 260 335 280
rect 355 260 360 280
rect 330 255 360 260
rect 240 195 270 200
rect 240 175 245 195
rect 265 175 270 195
rect 240 170 270 175
rect 245 165 265 170
rect 290 150 310 255
rect 335 250 355 255
rect 425 200 445 375
rect 605 200 625 375
rect 740 370 760 375
rect 740 325 760 330
rect 735 320 765 325
rect 735 300 740 320
rect 760 300 765 320
rect 735 295 765 300
rect 420 195 450 200
rect 420 175 425 195
rect 445 175 450 195
rect 420 170 450 175
rect 600 195 630 200
rect 600 175 605 195
rect 625 175 630 195
rect 600 170 630 175
rect 425 165 445 170
rect 605 165 625 170
rect 740 150 760 295
rect 785 200 805 375
rect 965 200 985 375
rect 780 195 810 200
rect 780 175 785 195
rect 805 175 810 195
rect 780 170 810 175
rect 960 195 990 200
rect 960 175 965 195
rect 985 175 990 195
rect 960 170 990 175
rect 785 165 805 170
rect 965 165 985 170
rect 1100 150 1120 375
rect 1145 200 1165 375
rect 1325 200 1345 375
rect 1460 370 1480 375
rect 1460 325 1480 330
rect 1455 320 1485 325
rect 1455 300 1460 320
rect 1480 300 1485 320
rect 1455 295 1485 300
rect 1140 195 1170 200
rect 1140 175 1145 195
rect 1165 175 1170 195
rect 1140 170 1170 175
rect 1320 195 1350 200
rect 1320 175 1325 195
rect 1345 175 1350 195
rect 1320 170 1350 175
rect 1145 165 1165 170
rect 1325 165 1345 170
rect 1460 150 1480 295
rect 1505 200 1525 375
rect 1685 200 1705 375
rect 1865 200 1885 375
rect 2045 200 2065 375
rect 2225 365 2245 370
rect 2405 365 2425 370
rect 2540 365 2560 750
rect 2675 730 2695 735
rect 2855 730 2875 735
rect 3035 730 3055 735
rect 3215 730 3235 735
rect 3395 730 3415 735
rect 3575 730 3595 735
rect 3755 730 3775 735
rect 3935 730 3955 735
rect 2670 725 2700 730
rect 2670 705 2675 725
rect 2695 705 2700 725
rect 2670 700 2700 705
rect 2850 725 2880 730
rect 2850 705 2855 725
rect 2875 705 2880 725
rect 2850 700 2880 705
rect 3030 725 3060 730
rect 3030 705 3035 725
rect 3055 705 3060 725
rect 3030 700 3060 705
rect 3210 725 3240 730
rect 3210 705 3215 725
rect 3235 705 3240 725
rect 3210 700 3240 705
rect 3390 725 3420 730
rect 3390 705 3395 725
rect 3415 705 3420 725
rect 3390 700 3420 705
rect 3570 725 3600 730
rect 3570 705 3575 725
rect 3595 705 3600 725
rect 3570 700 3600 705
rect 3750 725 3780 730
rect 3750 705 3755 725
rect 3775 705 3780 725
rect 3750 700 3780 705
rect 3930 725 3960 730
rect 3930 705 3935 725
rect 3955 705 3960 725
rect 3930 700 3960 705
rect 2675 525 2695 700
rect 2855 525 2875 700
rect 3035 565 3055 700
rect 3215 565 3235 700
rect 3395 565 3415 700
rect 3575 565 3595 700
rect 3030 560 3060 565
rect 3030 540 3035 560
rect 3055 540 3060 560
rect 3030 535 3060 540
rect 3210 560 3240 565
rect 3210 540 3215 560
rect 3235 540 3240 560
rect 3210 535 3240 540
rect 3390 560 3420 565
rect 3390 540 3395 560
rect 3415 540 3420 560
rect 3390 535 3420 540
rect 3570 560 3600 565
rect 3570 540 3575 560
rect 3595 540 3600 560
rect 3570 535 3600 540
rect 3035 530 3055 535
rect 3215 530 3235 535
rect 3395 530 3415 535
rect 3575 530 3595 535
rect 3755 525 3775 700
rect 3935 525 3955 700
rect 2670 520 2700 525
rect 2670 500 2675 520
rect 2695 500 2700 520
rect 2670 495 2700 500
rect 2850 520 2880 525
rect 2850 500 2855 520
rect 2875 500 2880 520
rect 2850 495 2880 500
rect 3750 520 3780 525
rect 3750 500 3755 520
rect 3775 500 3780 520
rect 3750 495 3780 500
rect 3930 520 3960 525
rect 3930 500 3935 520
rect 3955 500 3960 520
rect 3930 495 3960 500
rect 2675 490 2695 495
rect 2855 490 2875 495
rect 3755 490 3775 495
rect 3935 490 3955 495
rect 3305 445 3325 450
rect 3485 445 3505 450
rect 3665 445 3685 450
rect 3845 445 3865 450
rect 3980 445 4000 750
rect 4115 730 4135 735
rect 4110 725 4140 730
rect 4110 705 4115 725
rect 4135 705 4140 725
rect 4110 700 4140 705
rect 4070 565 4090 570
rect 4065 560 4095 565
rect 4065 540 4070 560
rect 4090 540 4095 560
rect 4065 535 4095 540
rect 3300 440 3330 445
rect 3300 420 3305 440
rect 3325 420 3330 440
rect 3300 415 3330 420
rect 3480 440 3510 445
rect 3480 420 3485 440
rect 3505 420 3510 440
rect 3480 415 3510 420
rect 3660 440 3690 445
rect 3660 420 3665 440
rect 3685 420 3690 440
rect 3660 415 3690 420
rect 3840 440 3870 445
rect 3840 420 3845 440
rect 3865 420 3870 440
rect 3840 415 3870 420
rect 3975 440 4005 445
rect 3975 420 3980 440
rect 4000 420 4005 440
rect 3975 415 4005 420
rect 2945 405 2965 410
rect 3125 405 3145 410
rect 2940 400 2970 405
rect 2940 380 2945 400
rect 2965 380 2970 400
rect 2940 375 2970 380
rect 3120 400 3150 405
rect 3120 380 3125 400
rect 3145 380 3150 400
rect 3120 375 3150 380
rect 2585 365 2605 370
rect 2765 365 2785 370
rect 2220 360 2250 365
rect 2220 340 2225 360
rect 2245 340 2250 360
rect 2220 335 2250 340
rect 2400 360 2430 365
rect 2400 340 2405 360
rect 2425 340 2430 360
rect 2400 335 2430 340
rect 2535 360 2565 365
rect 2535 340 2540 360
rect 2560 340 2565 360
rect 2535 335 2565 340
rect 2580 360 2610 365
rect 2580 340 2585 360
rect 2605 340 2610 360
rect 2580 335 2610 340
rect 2760 360 2790 365
rect 2760 340 2765 360
rect 2785 340 2790 360
rect 2760 335 2790 340
rect 2180 325 2200 330
rect 2175 320 2205 325
rect 2175 300 2180 320
rect 2200 300 2205 320
rect 2175 295 2205 300
rect 1500 195 1530 200
rect 1500 175 1505 195
rect 1525 175 1530 195
rect 1500 170 1530 175
rect 1680 195 1710 200
rect 1680 175 1685 195
rect 1705 175 1710 195
rect 1680 170 1710 175
rect 1860 195 1890 200
rect 1860 175 1865 195
rect 1885 175 1890 195
rect 1860 170 1890 175
rect 2040 195 2070 200
rect 2040 175 2045 195
rect 2065 175 2070 195
rect 2040 170 2070 175
rect 1505 165 1525 170
rect 1685 165 1705 170
rect 1865 165 1885 170
rect 2045 165 2065 170
rect 2180 150 2200 295
rect 2225 200 2245 335
rect 2405 200 2425 335
rect 2220 195 2250 200
rect 2220 175 2225 195
rect 2245 175 2250 195
rect 2220 170 2250 175
rect 2400 195 2430 200
rect 2400 175 2405 195
rect 2425 175 2430 195
rect 2400 170 2430 175
rect 2225 165 2245 170
rect 2405 165 2425 170
rect 2540 150 2560 335
rect 2585 200 2605 335
rect 2765 200 2785 335
rect 2900 325 2920 330
rect 2895 320 2925 325
rect 2895 300 2900 320
rect 2920 300 2925 320
rect 2895 295 2925 300
rect 2580 195 2610 200
rect 2580 175 2585 195
rect 2605 175 2610 195
rect 2580 170 2610 175
rect 2760 195 2790 200
rect 2760 175 2765 195
rect 2785 175 2790 195
rect 2760 170 2790 175
rect 2585 165 2605 170
rect 2765 165 2785 170
rect 2900 150 2920 295
rect 2945 200 2965 375
rect 3125 200 3145 375
rect 3305 200 3325 415
rect 3485 200 3505 415
rect 3665 200 3685 415
rect 3845 200 3865 415
rect 2940 195 2970 200
rect 2940 175 2945 195
rect 2965 175 2970 195
rect 2940 170 2970 175
rect 3120 195 3150 200
rect 3120 175 3125 195
rect 3145 175 3150 195
rect 3120 170 3150 175
rect 3300 195 3330 200
rect 3300 175 3305 195
rect 3325 175 3330 195
rect 3300 170 3330 175
rect 3480 195 3510 200
rect 3480 175 3485 195
rect 3505 175 3510 195
rect 3480 170 3510 175
rect 3660 195 3690 200
rect 3660 175 3665 195
rect 3685 175 3690 195
rect 3660 170 3690 175
rect 3840 195 3870 200
rect 3840 175 3845 195
rect 3865 175 3870 195
rect 3840 170 3870 175
rect 2945 165 2965 170
rect 3125 165 3145 170
rect 3305 165 3325 170
rect 3485 165 3505 170
rect 3665 165 3685 170
rect 3845 165 3865 170
rect 3980 150 4000 415
rect 4025 285 4045 290
rect 4020 280 4050 285
rect 4020 260 4025 280
rect 4045 260 4050 280
rect 4020 255 4050 260
rect 4025 200 4045 255
rect 4020 195 4050 200
rect 4020 175 4025 195
rect 4045 175 4050 195
rect 4020 170 4050 175
rect 4025 165 4045 170
rect 4070 150 4090 535
rect 4115 445 4135 700
rect 4160 445 4180 750
rect 4295 730 4315 735
rect 4475 730 4495 735
rect 4655 730 4675 735
rect 4835 730 4855 735
rect 5015 730 5035 735
rect 5195 730 5215 735
rect 5375 730 5395 735
rect 5555 730 5575 735
rect 4290 725 4320 730
rect 4290 705 4295 725
rect 4315 705 4320 725
rect 4290 700 4320 705
rect 4470 725 4500 730
rect 4470 705 4475 725
rect 4495 705 4500 725
rect 4470 700 4500 705
rect 4650 725 4680 730
rect 4650 705 4655 725
rect 4675 705 4680 725
rect 4650 700 4680 705
rect 4830 725 4860 730
rect 4830 705 4835 725
rect 4855 705 4860 725
rect 4830 700 4860 705
rect 5010 725 5040 730
rect 5010 705 5015 725
rect 5035 705 5040 725
rect 5010 700 5040 705
rect 5190 725 5220 730
rect 5190 705 5195 725
rect 5215 705 5220 725
rect 5190 700 5220 705
rect 5370 725 5400 730
rect 5370 705 5375 725
rect 5395 705 5400 725
rect 5370 700 5400 705
rect 5550 725 5580 730
rect 5550 705 5555 725
rect 5575 705 5580 725
rect 5550 700 5580 705
rect 4295 525 4315 700
rect 4475 525 4495 700
rect 4655 565 4675 700
rect 4835 565 4855 700
rect 5015 645 5035 700
rect 5195 645 5215 700
rect 5010 640 5040 645
rect 5010 620 5015 640
rect 5035 620 5040 640
rect 5010 615 5040 620
rect 5190 640 5220 645
rect 5190 620 5195 640
rect 5215 620 5220 640
rect 5190 615 5220 620
rect 5015 610 5035 615
rect 5195 610 5215 615
rect 4650 560 4680 565
rect 4650 540 4655 560
rect 4675 540 4680 560
rect 4650 535 4680 540
rect 4830 560 4860 565
rect 4830 540 4835 560
rect 4855 540 4860 560
rect 4830 535 4860 540
rect 4655 530 4675 535
rect 4835 530 4855 535
rect 5375 525 5395 700
rect 5555 525 5575 700
rect 5600 645 5620 750
rect 5735 730 5755 735
rect 5915 730 5935 735
rect 6095 730 6115 735
rect 6275 730 6295 735
rect 6455 730 6475 735
rect 6635 730 6655 735
rect 6815 730 6835 735
rect 6995 730 7015 735
rect 5730 725 5760 730
rect 5730 705 5735 725
rect 5755 705 5760 725
rect 5730 700 5760 705
rect 5910 725 5940 730
rect 5910 705 5915 725
rect 5935 705 5940 725
rect 5910 700 5940 705
rect 6090 725 6120 730
rect 6090 705 6095 725
rect 6115 705 6120 725
rect 6090 700 6120 705
rect 6270 725 6300 730
rect 6270 705 6275 725
rect 6295 705 6300 725
rect 6270 700 6300 705
rect 6450 725 6480 730
rect 6450 705 6455 725
rect 6475 705 6480 725
rect 6450 700 6480 705
rect 6630 725 6660 730
rect 6630 705 6635 725
rect 6655 705 6660 725
rect 6630 700 6660 705
rect 6810 725 6840 730
rect 6810 705 6815 725
rect 6835 705 6840 725
rect 6810 700 6840 705
rect 6990 725 7020 730
rect 6990 705 6995 725
rect 7015 705 7020 725
rect 6990 700 7020 705
rect 5595 640 5625 645
rect 5595 620 5600 640
rect 5620 620 5625 640
rect 5595 615 5625 620
rect 4290 520 4320 525
rect 4290 500 4295 520
rect 4315 500 4320 520
rect 4290 495 4320 500
rect 4470 520 4500 525
rect 4470 500 4475 520
rect 4495 500 4500 520
rect 4470 495 4500 500
rect 5370 520 5400 525
rect 5370 500 5375 520
rect 5395 500 5400 520
rect 5370 495 5400 500
rect 5550 520 5580 525
rect 5550 500 5555 520
rect 5575 500 5580 520
rect 5550 495 5580 500
rect 4295 490 4315 495
rect 4475 490 4495 495
rect 5375 490 5395 495
rect 5555 490 5575 495
rect 4205 445 4225 450
rect 4385 445 4405 450
rect 4565 445 4585 450
rect 4745 445 4765 450
rect 4110 440 4140 445
rect 4110 420 4115 440
rect 4135 420 4140 440
rect 4110 415 4140 420
rect 4155 440 4185 445
rect 4155 420 4160 440
rect 4180 420 4185 440
rect 4155 415 4185 420
rect 4200 440 4230 445
rect 4200 420 4205 440
rect 4225 420 4230 440
rect 4200 415 4230 420
rect 4380 440 4410 445
rect 4380 420 4385 440
rect 4405 420 4410 440
rect 4380 415 4410 420
rect 4560 440 4590 445
rect 4560 420 4565 440
rect 4585 420 4590 440
rect 4560 415 4590 420
rect 4740 440 4770 445
rect 4740 420 4745 440
rect 4765 420 4770 440
rect 4740 415 4770 420
rect 4115 410 4135 415
rect 4160 150 4180 415
rect 4205 200 4225 415
rect 4385 200 4405 415
rect 4565 200 4585 415
rect 4745 200 4765 415
rect 4925 365 4945 370
rect 5105 365 5125 370
rect 5285 365 5305 370
rect 5465 365 5485 370
rect 4920 360 4950 365
rect 4920 340 4925 360
rect 4945 340 4950 360
rect 4920 335 4950 340
rect 5100 360 5130 365
rect 5100 340 5105 360
rect 5125 340 5130 360
rect 5100 335 5130 340
rect 5280 360 5310 365
rect 5280 340 5285 360
rect 5305 340 5310 360
rect 5280 335 5310 340
rect 5460 360 5490 365
rect 5460 340 5465 360
rect 5485 340 5490 360
rect 5460 335 5490 340
rect 4925 200 4945 335
rect 5105 200 5125 335
rect 5285 200 5305 335
rect 5465 200 5485 335
rect 4200 195 4230 200
rect 4200 175 4205 195
rect 4225 175 4230 195
rect 4200 170 4230 175
rect 4380 195 4410 200
rect 4380 175 4385 195
rect 4405 175 4410 195
rect 4380 170 4410 175
rect 4560 195 4590 200
rect 4560 175 4565 195
rect 4585 175 4590 195
rect 4560 170 4590 175
rect 4740 195 4770 200
rect 4740 175 4745 195
rect 4765 175 4770 195
rect 4740 170 4770 175
rect 4920 195 4950 200
rect 4920 175 4925 195
rect 4945 175 4950 195
rect 4920 170 4950 175
rect 5100 195 5130 200
rect 5100 175 5105 195
rect 5125 175 5130 195
rect 5100 170 5130 175
rect 5280 195 5310 200
rect 5280 175 5285 195
rect 5305 175 5310 195
rect 5280 170 5310 175
rect 5460 195 5490 200
rect 5460 175 5465 195
rect 5485 175 5490 195
rect 5460 170 5490 175
rect 4205 165 4225 170
rect 4385 165 4405 170
rect 4565 165 4585 170
rect 4745 165 4765 170
rect 4925 165 4945 170
rect 5105 165 5125 170
rect 5285 165 5305 170
rect 5465 165 5485 170
rect 5600 150 5620 615
rect 5735 525 5755 700
rect 5915 525 5935 700
rect 6095 645 6115 700
rect 6275 645 6295 700
rect 6455 645 6475 700
rect 6635 645 6655 700
rect 6090 640 6120 645
rect 6090 620 6095 640
rect 6115 620 6120 640
rect 6090 615 6120 620
rect 6270 640 6300 645
rect 6270 620 6275 640
rect 6295 620 6300 640
rect 6270 615 6300 620
rect 6450 640 6480 645
rect 6450 620 6455 640
rect 6475 620 6480 640
rect 6450 615 6480 620
rect 6630 640 6660 645
rect 6630 620 6635 640
rect 6655 620 6660 640
rect 6630 615 6660 620
rect 6095 610 6115 615
rect 6275 610 6295 615
rect 6455 610 6475 615
rect 6635 610 6655 615
rect 6815 525 6835 700
rect 6995 525 7015 700
rect 7040 565 7060 750
rect 7175 730 7195 735
rect 7355 730 7375 735
rect 7535 730 7555 735
rect 7715 730 7735 735
rect 7900 730 7920 735
rect 8080 730 8100 735
rect 8260 730 8280 735
rect 8440 730 8460 735
rect 7170 725 7200 730
rect 7170 705 7175 725
rect 7195 705 7200 725
rect 7170 700 7200 705
rect 7350 725 7380 730
rect 7350 705 7355 725
rect 7375 705 7380 725
rect 7350 700 7380 705
rect 7530 725 7560 730
rect 7530 705 7535 725
rect 7555 705 7560 725
rect 7530 700 7560 705
rect 7710 725 7740 730
rect 7710 705 7715 725
rect 7735 705 7740 725
rect 7710 700 7740 705
rect 7895 725 7925 730
rect 7895 705 7900 725
rect 7920 705 7925 725
rect 7895 700 7925 705
rect 8075 725 8105 730
rect 8075 705 8080 725
rect 8100 705 8105 725
rect 8075 700 8105 705
rect 8255 725 8285 730
rect 8255 705 8260 725
rect 8280 705 8285 725
rect 8255 700 8285 705
rect 8435 725 8465 730
rect 8435 705 8440 725
rect 8460 705 8465 725
rect 8435 700 8465 705
rect 7035 560 7065 565
rect 7035 540 7040 560
rect 7060 540 7065 560
rect 7035 535 7065 540
rect 5730 520 5760 525
rect 5730 500 5735 520
rect 5755 500 5760 520
rect 5730 495 5760 500
rect 5910 520 5940 525
rect 5910 500 5915 520
rect 5935 500 5940 520
rect 5910 495 5940 500
rect 6810 520 6840 525
rect 6810 500 6815 520
rect 6835 500 6840 520
rect 6810 495 6840 500
rect 6990 520 7020 525
rect 6990 500 6995 520
rect 7015 500 7020 520
rect 6990 495 7020 500
rect 5735 490 5755 495
rect 5915 490 5935 495
rect 6815 490 6835 495
rect 6995 490 7015 495
rect 6365 445 6385 450
rect 6545 445 6565 450
rect 6725 445 6745 450
rect 6905 445 6925 450
rect 6360 440 6390 445
rect 6360 420 6365 440
rect 6385 420 6390 440
rect 6360 415 6390 420
rect 6540 440 6570 445
rect 6540 420 6545 440
rect 6565 420 6570 440
rect 6540 415 6570 420
rect 6720 440 6750 445
rect 6720 420 6725 440
rect 6745 420 6750 440
rect 6720 415 6750 420
rect 6900 440 6930 445
rect 6900 420 6905 440
rect 6925 420 6930 440
rect 6900 415 6930 420
rect 5645 365 5665 370
rect 5825 365 5845 370
rect 6005 365 6025 370
rect 6185 365 6205 370
rect 5640 360 5670 365
rect 5640 340 5645 360
rect 5665 340 5670 360
rect 5640 335 5670 340
rect 5820 360 5850 365
rect 5820 340 5825 360
rect 5845 340 5850 360
rect 5820 335 5850 340
rect 6000 360 6030 365
rect 6000 340 6005 360
rect 6025 340 6030 360
rect 6000 335 6030 340
rect 6180 360 6210 365
rect 6180 340 6185 360
rect 6205 340 6210 360
rect 6180 335 6210 340
rect 5645 200 5665 335
rect 5825 200 5845 335
rect 6005 200 6025 335
rect 6185 200 6205 335
rect 6365 200 6385 415
rect 6545 200 6565 415
rect 6725 200 6745 415
rect 6905 200 6925 415
rect 5640 195 5670 200
rect 5640 175 5645 195
rect 5665 175 5670 195
rect 5640 170 5670 175
rect 5820 195 5850 200
rect 5820 175 5825 195
rect 5845 175 5850 195
rect 5820 170 5850 175
rect 6000 195 6030 200
rect 6000 175 6005 195
rect 6025 175 6030 195
rect 6000 170 6030 175
rect 6180 195 6210 200
rect 6180 175 6185 195
rect 6205 175 6210 195
rect 6180 170 6210 175
rect 6360 195 6390 200
rect 6360 175 6365 195
rect 6385 175 6390 195
rect 6360 170 6390 175
rect 6540 195 6570 200
rect 6540 175 6545 195
rect 6565 175 6570 195
rect 6540 170 6570 175
rect 6720 195 6750 200
rect 6720 175 6725 195
rect 6745 175 6750 195
rect 6720 170 6750 175
rect 6900 195 6930 200
rect 6900 175 6905 195
rect 6925 175 6930 195
rect 6900 170 6930 175
rect 5645 165 5665 170
rect 5825 165 5845 170
rect 6005 165 6025 170
rect 6185 165 6205 170
rect 6365 165 6385 170
rect 6545 165 6565 170
rect 6725 165 6745 170
rect 6905 165 6925 170
rect 7040 150 7060 535
rect 7175 525 7195 700
rect 7355 525 7375 700
rect 7535 645 7555 700
rect 7715 645 7735 700
rect 7530 640 7560 645
rect 7530 620 7535 640
rect 7555 620 7560 640
rect 7530 615 7560 620
rect 7710 640 7740 645
rect 7710 620 7715 640
rect 7735 620 7740 640
rect 7710 615 7740 620
rect 7535 610 7555 615
rect 7715 610 7735 615
rect 7900 525 7920 700
rect 8080 525 8100 700
rect 8125 525 8145 530
rect 8260 525 8280 700
rect 8440 525 8460 700
rect 8485 525 8505 750
rect 8620 730 8640 735
rect 8800 730 8820 735
rect 8980 730 9000 735
rect 9160 730 9180 735
rect 9340 730 9360 735
rect 9520 730 9540 735
rect 9700 730 9720 735
rect 9880 730 9900 735
rect 8615 725 8645 730
rect 8615 705 8620 725
rect 8640 705 8645 725
rect 8615 700 8645 705
rect 8795 725 8825 730
rect 8795 705 8800 725
rect 8820 705 8825 725
rect 8795 700 8825 705
rect 8975 725 9005 730
rect 8975 705 8980 725
rect 9000 705 9005 725
rect 8975 700 9005 705
rect 9155 725 9185 730
rect 9155 705 9160 725
rect 9180 705 9185 725
rect 9155 700 9185 705
rect 9335 725 9365 730
rect 9335 705 9340 725
rect 9360 705 9365 725
rect 9335 700 9365 705
rect 9515 725 9545 730
rect 9515 705 9520 725
rect 9540 705 9545 725
rect 9515 700 9545 705
rect 9695 725 9725 730
rect 9695 705 9700 725
rect 9720 705 9725 725
rect 9695 700 9725 705
rect 9875 725 9905 730
rect 9875 705 9880 725
rect 9900 705 9905 725
rect 9875 700 9905 705
rect 8620 525 8640 700
rect 8800 525 8820 700
rect 8845 525 8865 530
rect 8980 525 9000 700
rect 9160 525 9180 700
rect 9340 565 9360 700
rect 9520 565 9540 700
rect 9335 560 9365 565
rect 9335 540 9340 560
rect 9360 540 9365 560
rect 9335 535 9365 540
rect 9515 560 9545 565
rect 9515 540 9520 560
rect 9540 540 9545 560
rect 9515 535 9545 540
rect 9340 530 9360 535
rect 9520 530 9540 535
rect 9700 525 9720 700
rect 9880 525 9900 700
rect 7170 520 7200 525
rect 7170 500 7175 520
rect 7195 500 7200 520
rect 7170 495 7200 500
rect 7350 520 7380 525
rect 7350 500 7355 520
rect 7375 500 7380 520
rect 7350 495 7380 500
rect 7895 520 7925 525
rect 7895 500 7900 520
rect 7920 500 7925 520
rect 7895 495 7925 500
rect 8075 520 8105 525
rect 8075 500 8080 520
rect 8100 500 8105 520
rect 8075 495 8105 500
rect 8120 520 8150 525
rect 8120 500 8125 520
rect 8145 500 8150 520
rect 8120 495 8150 500
rect 8255 520 8285 525
rect 8255 500 8260 520
rect 8280 500 8285 520
rect 8255 495 8285 500
rect 8435 520 8465 525
rect 8435 500 8440 520
rect 8460 500 8465 520
rect 8435 495 8465 500
rect 8480 520 8510 525
rect 8480 500 8485 520
rect 8505 500 8510 520
rect 8480 495 8510 500
rect 8615 520 8645 525
rect 8615 500 8620 520
rect 8640 500 8645 520
rect 8615 495 8645 500
rect 8795 520 8825 525
rect 8795 500 8800 520
rect 8820 500 8825 520
rect 8795 495 8825 500
rect 8840 520 8870 525
rect 8840 500 8845 520
rect 8865 500 8870 520
rect 8840 495 8870 500
rect 8975 520 9005 525
rect 8975 500 8980 520
rect 9000 500 9005 520
rect 8975 495 9005 500
rect 9155 520 9185 525
rect 9155 500 9160 520
rect 9180 500 9185 520
rect 9155 495 9185 500
rect 9695 520 9725 525
rect 9695 500 9700 520
rect 9720 500 9725 520
rect 9695 495 9725 500
rect 9875 520 9905 525
rect 9875 500 9880 520
rect 9900 500 9905 520
rect 9875 495 9905 500
rect 7175 490 7195 495
rect 7355 490 7375 495
rect 7900 490 7920 495
rect 8080 490 8100 495
rect 7085 445 7105 450
rect 7265 445 7285 450
rect 7445 445 7465 450
rect 7625 445 7645 450
rect 7810 445 7830 450
rect 7990 445 8010 450
rect 7080 440 7110 445
rect 7080 420 7085 440
rect 7105 420 7110 440
rect 7080 415 7110 420
rect 7260 440 7290 445
rect 7260 420 7265 440
rect 7285 420 7290 440
rect 7260 415 7290 420
rect 7440 440 7470 445
rect 7440 420 7445 440
rect 7465 420 7470 440
rect 7440 415 7470 420
rect 7620 440 7650 445
rect 7620 420 7625 440
rect 7645 420 7650 440
rect 7620 415 7650 420
rect 7805 440 7835 445
rect 7805 420 7810 440
rect 7830 420 7835 440
rect 7805 415 7835 420
rect 7985 440 8015 445
rect 7985 420 7990 440
rect 8010 420 8015 440
rect 7985 415 8015 420
rect 7085 200 7105 415
rect 7265 200 7285 415
rect 7445 200 7465 415
rect 7625 200 7645 415
rect 7810 200 7830 415
rect 7990 200 8010 415
rect 7080 195 7110 200
rect 7080 175 7085 195
rect 7105 175 7110 195
rect 7080 170 7110 175
rect 7260 195 7290 200
rect 7260 175 7265 195
rect 7285 175 7290 195
rect 7260 170 7290 175
rect 7440 195 7470 200
rect 7440 175 7445 195
rect 7465 175 7470 195
rect 7440 170 7470 175
rect 7620 195 7650 200
rect 7620 175 7625 195
rect 7645 175 7650 195
rect 7620 170 7650 175
rect 7805 195 7835 200
rect 7805 175 7810 195
rect 7830 175 7835 195
rect 7805 170 7835 175
rect 7985 195 8015 200
rect 7985 175 7990 195
rect 8010 175 8015 195
rect 7985 170 8015 175
rect 7085 165 7105 170
rect 7265 165 7285 170
rect 7445 165 7465 170
rect 7625 165 7645 170
rect 7810 165 7830 170
rect 7990 165 8010 170
rect 8125 150 8145 495
rect 8260 490 8280 495
rect 8440 490 8460 495
rect 8485 490 8505 495
rect 8620 490 8640 495
rect 8800 490 8820 495
rect 8170 445 8190 450
rect 8350 445 8370 450
rect 8530 445 8550 450
rect 8710 445 8730 450
rect 8165 440 8195 445
rect 8165 420 8170 440
rect 8190 420 8195 440
rect 8165 415 8195 420
rect 8345 440 8375 445
rect 8345 420 8350 440
rect 8370 420 8375 440
rect 8345 415 8375 420
rect 8525 440 8555 445
rect 8525 420 8530 440
rect 8550 420 8555 440
rect 8525 415 8555 420
rect 8705 440 8735 445
rect 8705 420 8710 440
rect 8730 420 8735 440
rect 8705 415 8735 420
rect 8170 200 8190 415
rect 8350 200 8370 415
rect 8530 200 8550 415
rect 8710 200 8730 415
rect 8165 195 8195 200
rect 8165 175 8170 195
rect 8190 175 8195 195
rect 8165 170 8195 175
rect 8345 195 8375 200
rect 8345 175 8350 195
rect 8370 175 8375 195
rect 8345 170 8375 175
rect 8525 195 8555 200
rect 8525 175 8530 195
rect 8550 175 8555 195
rect 8525 170 8555 175
rect 8705 195 8735 200
rect 8705 175 8710 195
rect 8730 175 8735 195
rect 8705 170 8735 175
rect 8170 165 8190 170
rect 8350 165 8370 170
rect 8530 165 8550 170
rect 8710 165 8730 170
rect 8845 150 8865 495
rect 8980 490 9000 495
rect 9160 490 9180 495
rect 9700 490 9720 495
rect 9880 490 9900 495
rect 9925 485 9945 750
rect 10060 730 10080 735
rect 10240 730 10260 735
rect 10420 730 10440 735
rect 10600 730 10620 735
rect 10055 725 10085 730
rect 10055 705 10060 725
rect 10080 705 10085 725
rect 10055 700 10085 705
rect 10235 725 10265 730
rect 10235 705 10240 725
rect 10260 705 10265 725
rect 10235 700 10265 705
rect 10415 725 10445 730
rect 10415 705 10420 725
rect 10440 705 10445 725
rect 10415 700 10445 705
rect 10595 725 10625 730
rect 10595 705 10600 725
rect 10620 705 10625 725
rect 10595 700 10625 705
rect 10060 525 10080 700
rect 10240 525 10260 700
rect 10420 565 10440 700
rect 10600 565 10620 700
rect 10735 645 10755 750
rect 10730 640 10760 645
rect 10730 620 10735 640
rect 10755 620 10760 640
rect 10730 615 10760 620
rect 10415 560 10445 565
rect 10415 540 10420 560
rect 10440 540 10445 560
rect 10415 535 10445 540
rect 10595 560 10625 565
rect 10595 540 10600 560
rect 10620 540 10625 560
rect 10595 535 10625 540
rect 10420 530 10440 535
rect 10600 530 10620 535
rect 10055 520 10085 525
rect 10055 500 10060 520
rect 10080 500 10085 520
rect 10055 495 10085 500
rect 10235 520 10265 525
rect 10235 500 10240 520
rect 10260 500 10265 520
rect 10235 495 10265 500
rect 10060 490 10080 495
rect 10240 490 10260 495
rect 9920 480 9950 485
rect 9920 460 9925 480
rect 9945 460 9950 480
rect 9920 455 9950 460
rect 9925 450 9945 455
rect 8890 445 8910 450
rect 9070 445 9090 450
rect 8885 440 8915 445
rect 8885 420 8890 440
rect 8910 420 8915 440
rect 8885 415 8915 420
rect 9065 440 9095 445
rect 9065 420 9070 440
rect 9090 420 9095 440
rect 9065 415 9095 420
rect 8890 200 8910 415
rect 9070 200 9090 415
rect 9250 325 9270 330
rect 9430 325 9450 330
rect 9610 325 9630 330
rect 9790 325 9810 330
rect 9970 325 9990 330
rect 10150 325 10170 330
rect 10330 325 10350 330
rect 10510 325 10530 330
rect 9245 320 9275 325
rect 9245 300 9250 320
rect 9270 300 9275 320
rect 9245 295 9275 300
rect 9425 320 9455 325
rect 9425 300 9430 320
rect 9450 300 9455 320
rect 9425 295 9455 300
rect 9605 320 9635 325
rect 9605 300 9610 320
rect 9630 300 9635 320
rect 9605 295 9635 300
rect 9785 320 9815 325
rect 9785 300 9790 320
rect 9810 300 9815 320
rect 9785 295 9815 300
rect 9965 320 9995 325
rect 9965 300 9970 320
rect 9990 300 9995 320
rect 9965 295 9995 300
rect 10145 320 10175 325
rect 10145 300 10150 320
rect 10170 300 10175 320
rect 10145 295 10175 300
rect 10325 320 10355 325
rect 10325 300 10330 320
rect 10350 300 10355 320
rect 10325 295 10355 300
rect 10505 320 10535 325
rect 10505 300 10510 320
rect 10530 300 10535 320
rect 10505 295 10535 300
rect 9250 200 9270 295
rect 9430 200 9450 295
rect 9610 200 9630 295
rect 9790 200 9810 295
rect 9970 200 9990 295
rect 10150 200 10170 295
rect 10330 200 10350 295
rect 10510 200 10530 295
rect 8885 195 8915 200
rect 8885 175 8890 195
rect 8910 175 8915 195
rect 8885 170 8915 175
rect 9065 195 9095 200
rect 9065 175 9070 195
rect 9090 175 9095 195
rect 9065 170 9095 175
rect 9245 195 9275 200
rect 9245 175 9250 195
rect 9270 175 9275 195
rect 9245 170 9275 175
rect 9425 195 9455 200
rect 9425 175 9430 195
rect 9450 175 9455 195
rect 9425 170 9455 175
rect 9605 195 9635 200
rect 9605 175 9610 195
rect 9630 175 9635 195
rect 9605 170 9635 175
rect 9785 195 9815 200
rect 9785 175 9790 195
rect 9810 175 9815 195
rect 9785 170 9815 175
rect 9965 195 9995 200
rect 9965 175 9970 195
rect 9990 175 9995 195
rect 9965 170 9995 175
rect 10145 195 10175 200
rect 10145 175 10150 195
rect 10170 175 10175 195
rect 10145 170 10175 175
rect 10325 195 10355 200
rect 10325 175 10330 195
rect 10350 175 10355 195
rect 10325 170 10355 175
rect 10505 195 10535 200
rect 10505 175 10510 195
rect 10530 175 10535 195
rect 10505 170 10535 175
rect 8890 165 8910 170
rect 9070 165 9090 170
rect 9250 165 9270 170
rect 9430 165 9450 170
rect 9610 165 9630 170
rect 9790 165 9810 170
rect 9970 165 9990 170
rect 10150 165 10170 170
rect 10330 165 10350 170
rect 10510 165 10530 170
rect 10735 150 10755 615
rect 10825 565 10845 750
rect 10820 560 10850 565
rect 10820 540 10825 560
rect 10845 540 10850 560
rect 10820 535 10850 540
rect 10825 150 10845 535
rect 10915 525 10935 750
rect 10910 520 10940 525
rect 10910 500 10915 520
rect 10935 500 10940 520
rect 10910 495 10940 500
rect 10915 150 10935 495
rect 11005 485 11025 750
rect 11000 480 11030 485
rect 11000 460 11005 480
rect 11025 460 11030 480
rect 11000 455 11030 460
rect 11005 150 11025 455
rect 11095 150 11115 750
rect -345 140 -315 150
rect -345 60 -340 140
rect -320 60 -315 140
rect -345 50 -315 60
rect -255 50 -225 150
rect -165 50 -135 150
rect -75 50 -45 150
rect 15 50 45 150
rect 105 50 135 150
rect 195 140 225 150
rect 195 60 200 140
rect 220 60 225 140
rect 195 50 225 60
rect 285 140 315 150
rect 285 60 290 140
rect 310 60 315 140
rect 285 50 315 60
rect 375 140 405 150
rect 375 60 380 140
rect 400 60 405 140
rect 375 50 405 60
rect 465 140 495 150
rect 465 60 470 140
rect 490 60 495 140
rect 465 50 495 60
rect 555 140 585 150
rect 555 60 560 140
rect 580 60 585 140
rect 555 50 585 60
rect 645 140 675 150
rect 645 60 650 140
rect 670 60 675 140
rect 645 50 675 60
rect 735 140 765 150
rect 735 60 740 140
rect 760 60 765 140
rect 735 50 765 60
rect 825 140 855 150
rect 825 60 830 140
rect 850 60 855 140
rect 825 50 855 60
rect 915 140 945 150
rect 915 60 920 140
rect 940 60 945 140
rect 915 50 945 60
rect 1005 140 1035 150
rect 1005 60 1010 140
rect 1030 60 1035 140
rect 1005 50 1035 60
rect 1095 140 1125 150
rect 1095 60 1100 140
rect 1120 60 1125 140
rect 1095 50 1125 60
rect 1185 140 1215 150
rect 1185 60 1190 140
rect 1210 60 1215 140
rect 1185 50 1215 60
rect 1275 140 1305 150
rect 1275 60 1280 140
rect 1300 60 1305 140
rect 1275 50 1305 60
rect 1365 140 1395 150
rect 1365 60 1370 140
rect 1390 60 1395 140
rect 1365 50 1395 60
rect 1455 140 1485 150
rect 1455 60 1460 140
rect 1480 60 1485 140
rect 1455 50 1485 60
rect 1545 140 1575 150
rect 1545 60 1550 140
rect 1570 60 1575 140
rect 1545 50 1575 60
rect 1635 140 1665 150
rect 1635 60 1640 140
rect 1660 60 1665 140
rect 1635 50 1665 60
rect 1725 140 1755 150
rect 1725 60 1730 140
rect 1750 60 1755 140
rect 1725 50 1755 60
rect 1815 140 1845 150
rect 1815 60 1820 140
rect 1840 60 1845 140
rect 1815 50 1845 60
rect 1905 140 1935 150
rect 1905 60 1910 140
rect 1930 60 1935 140
rect 1905 50 1935 60
rect 1995 140 2025 150
rect 1995 60 2000 140
rect 2020 60 2025 140
rect 1995 50 2025 60
rect 2085 140 2115 150
rect 2085 60 2090 140
rect 2110 60 2115 140
rect 2085 50 2115 60
rect 2175 140 2205 150
rect 2175 60 2180 140
rect 2200 60 2205 140
rect 2175 50 2205 60
rect 2265 140 2295 150
rect 2265 60 2270 140
rect 2290 60 2295 140
rect 2265 50 2295 60
rect 2355 140 2385 150
rect 2355 60 2360 140
rect 2380 60 2385 140
rect 2355 50 2385 60
rect 2445 140 2475 150
rect 2445 60 2450 140
rect 2470 60 2475 140
rect 2445 50 2475 60
rect 2535 140 2565 150
rect 2535 60 2540 140
rect 2560 60 2565 140
rect 2535 50 2565 60
rect 2625 140 2655 150
rect 2625 60 2630 140
rect 2650 60 2655 140
rect 2625 50 2655 60
rect 2715 140 2745 150
rect 2715 60 2720 140
rect 2740 60 2745 140
rect 2715 50 2745 60
rect 2805 140 2835 150
rect 2805 60 2810 140
rect 2830 60 2835 140
rect 2805 50 2835 60
rect 2895 140 2925 150
rect 2895 60 2900 140
rect 2920 60 2925 140
rect 2895 50 2925 60
rect 2985 140 3015 150
rect 2985 60 2990 140
rect 3010 60 3015 140
rect 2985 50 3015 60
rect 3075 140 3105 150
rect 3075 60 3080 140
rect 3100 60 3105 140
rect 3075 50 3105 60
rect 3165 140 3195 150
rect 3165 60 3170 140
rect 3190 60 3195 140
rect 3165 50 3195 60
rect 3255 140 3285 150
rect 3255 60 3260 140
rect 3280 60 3285 140
rect 3255 50 3285 60
rect 3345 140 3375 150
rect 3345 60 3350 140
rect 3370 60 3375 140
rect 3345 50 3375 60
rect 3435 140 3465 150
rect 3435 60 3440 140
rect 3460 60 3465 140
rect 3435 50 3465 60
rect 3525 140 3555 150
rect 3525 60 3530 140
rect 3550 60 3555 140
rect 3525 50 3555 60
rect 3615 140 3645 150
rect 3615 60 3620 140
rect 3640 60 3645 140
rect 3615 50 3645 60
rect 3705 140 3735 150
rect 3705 60 3710 140
rect 3730 60 3735 140
rect 3705 50 3735 60
rect 3795 140 3825 150
rect 3795 60 3800 140
rect 3820 60 3825 140
rect 3795 50 3825 60
rect 3885 140 3915 150
rect 3885 60 3890 140
rect 3910 60 3915 140
rect 3885 50 3915 60
rect 3975 140 4005 150
rect 3975 60 3980 140
rect 4000 60 4005 140
rect 3975 50 4005 60
rect 4065 140 4095 150
rect 4065 60 4070 140
rect 4090 60 4095 140
rect 4065 50 4095 60
rect 4155 140 4185 150
rect 4155 60 4160 140
rect 4180 60 4185 140
rect 4155 50 4185 60
rect 4245 140 4275 150
rect 4245 60 4250 140
rect 4270 60 4275 140
rect 4245 50 4275 60
rect 4335 140 4365 150
rect 4335 60 4340 140
rect 4360 60 4365 140
rect 4335 50 4365 60
rect 4425 140 4455 150
rect 4425 60 4430 140
rect 4450 60 4455 140
rect 4425 50 4455 60
rect 4515 140 4545 150
rect 4515 60 4520 140
rect 4540 60 4545 140
rect 4515 50 4545 60
rect 4605 140 4635 150
rect 4605 60 4610 140
rect 4630 60 4635 140
rect 4605 50 4635 60
rect 4695 140 4725 150
rect 4695 60 4700 140
rect 4720 60 4725 140
rect 4695 50 4725 60
rect 4785 140 4815 150
rect 4785 60 4790 140
rect 4810 60 4815 140
rect 4785 50 4815 60
rect 4875 140 4905 150
rect 4875 60 4880 140
rect 4900 60 4905 140
rect 4875 50 4905 60
rect 4965 140 4995 150
rect 4965 60 4970 140
rect 4990 60 4995 140
rect 4965 50 4995 60
rect 5055 140 5085 150
rect 5055 60 5060 140
rect 5080 60 5085 140
rect 5055 50 5085 60
rect 5145 140 5175 150
rect 5145 60 5150 140
rect 5170 60 5175 140
rect 5145 50 5175 60
rect 5235 140 5265 150
rect 5235 60 5240 140
rect 5260 60 5265 140
rect 5235 50 5265 60
rect 5325 140 5355 150
rect 5325 60 5330 140
rect 5350 60 5355 140
rect 5325 50 5355 60
rect 5415 140 5445 150
rect 5415 60 5420 140
rect 5440 60 5445 140
rect 5415 50 5445 60
rect 5505 140 5535 150
rect 5505 60 5510 140
rect 5530 60 5535 140
rect 5505 50 5535 60
rect 5595 140 5625 150
rect 5595 60 5600 140
rect 5620 60 5625 140
rect 5595 50 5625 60
rect 5685 140 5715 150
rect 5685 60 5690 140
rect 5710 60 5715 140
rect 5685 50 5715 60
rect 5775 140 5805 150
rect 5775 60 5780 140
rect 5800 60 5805 140
rect 5775 50 5805 60
rect 5865 140 5895 150
rect 5865 60 5870 140
rect 5890 60 5895 140
rect 5865 50 5895 60
rect 5955 140 5985 150
rect 5955 60 5960 140
rect 5980 60 5985 140
rect 5955 50 5985 60
rect 6045 140 6075 150
rect 6045 60 6050 140
rect 6070 60 6075 140
rect 6045 50 6075 60
rect 6135 140 6165 150
rect 6135 60 6140 140
rect 6160 60 6165 140
rect 6135 50 6165 60
rect 6225 140 6255 150
rect 6225 60 6230 140
rect 6250 60 6255 140
rect 6225 50 6255 60
rect 6315 140 6345 150
rect 6315 60 6320 140
rect 6340 60 6345 140
rect 6315 50 6345 60
rect 6405 140 6435 150
rect 6405 60 6410 140
rect 6430 60 6435 140
rect 6405 50 6435 60
rect 6495 140 6525 150
rect 6495 60 6500 140
rect 6520 60 6525 140
rect 6495 50 6525 60
rect 6585 140 6615 150
rect 6585 60 6590 140
rect 6610 60 6615 140
rect 6585 50 6615 60
rect 6675 140 6705 150
rect 6675 60 6680 140
rect 6700 60 6705 140
rect 6675 50 6705 60
rect 6765 140 6795 150
rect 6765 60 6770 140
rect 6790 60 6795 140
rect 6765 50 6795 60
rect 6855 140 6885 150
rect 6855 60 6860 140
rect 6880 60 6885 140
rect 6855 50 6885 60
rect 6945 140 6975 150
rect 6945 60 6950 140
rect 6970 60 6975 140
rect 6945 50 6975 60
rect 7035 140 7065 150
rect 7035 60 7040 140
rect 7060 60 7065 140
rect 7035 50 7065 60
rect 7125 140 7155 150
rect 7125 60 7130 140
rect 7150 60 7155 140
rect 7125 50 7155 60
rect 7215 140 7245 150
rect 7215 60 7220 140
rect 7240 60 7245 140
rect 7215 50 7245 60
rect 7305 140 7335 150
rect 7305 60 7310 140
rect 7330 60 7335 140
rect 7305 50 7335 60
rect 7395 140 7425 150
rect 7395 60 7400 140
rect 7420 60 7425 140
rect 7395 50 7425 60
rect 7485 140 7515 150
rect 7485 60 7490 140
rect 7510 60 7515 140
rect 7485 50 7515 60
rect 7575 140 7605 150
rect 7575 60 7580 140
rect 7600 60 7605 140
rect 7575 50 7605 60
rect 7665 140 7695 150
rect 7665 60 7670 140
rect 7690 60 7695 140
rect 7665 50 7695 60
rect 7755 140 7785 150
rect 7755 60 7760 140
rect 7780 60 7785 140
rect 7755 50 7785 60
rect 7850 140 7880 150
rect 7850 60 7855 140
rect 7875 60 7880 140
rect 7850 50 7880 60
rect 7940 140 7970 150
rect 7940 60 7945 140
rect 7965 60 7970 140
rect 7940 50 7970 60
rect 8030 140 8060 150
rect 8030 60 8035 140
rect 8055 60 8060 140
rect 8030 50 8060 60
rect 8120 140 8150 150
rect 8120 60 8125 140
rect 8145 60 8150 140
rect 8120 50 8150 60
rect 8210 140 8240 150
rect 8210 60 8215 140
rect 8235 60 8240 140
rect 8210 50 8240 60
rect 8300 140 8330 150
rect 8300 60 8305 140
rect 8325 60 8330 140
rect 8300 50 8330 60
rect 8390 140 8420 150
rect 8390 60 8395 140
rect 8415 60 8420 140
rect 8390 50 8420 60
rect 8480 140 8510 150
rect 8480 60 8485 140
rect 8505 60 8510 140
rect 8480 50 8510 60
rect 8570 140 8600 150
rect 8570 60 8575 140
rect 8595 60 8600 140
rect 8570 50 8600 60
rect 8660 140 8690 150
rect 8660 60 8665 140
rect 8685 60 8690 140
rect 8660 50 8690 60
rect 8750 140 8780 150
rect 8750 60 8755 140
rect 8775 60 8780 140
rect 8750 50 8780 60
rect 8840 140 8870 150
rect 8840 60 8845 140
rect 8865 60 8870 140
rect 8840 50 8870 60
rect 8930 140 8960 150
rect 8930 60 8935 140
rect 8955 60 8960 140
rect 8930 50 8960 60
rect 9020 140 9050 150
rect 9020 60 9025 140
rect 9045 60 9050 140
rect 9020 50 9050 60
rect 9110 140 9140 150
rect 9110 60 9115 140
rect 9135 60 9140 140
rect 9110 50 9140 60
rect 9200 140 9230 150
rect 9200 60 9205 140
rect 9225 60 9230 140
rect 9200 50 9230 60
rect 9290 140 9320 150
rect 9290 60 9295 140
rect 9315 60 9320 140
rect 9290 50 9320 60
rect 9380 140 9410 150
rect 9380 60 9385 140
rect 9405 60 9410 140
rect 9380 50 9410 60
rect 9470 140 9500 150
rect 9470 60 9475 140
rect 9495 60 9500 140
rect 9470 50 9500 60
rect 9560 140 9590 150
rect 9560 60 9565 140
rect 9585 60 9590 140
rect 9560 50 9590 60
rect 9650 140 9680 150
rect 9650 60 9655 140
rect 9675 60 9680 140
rect 9650 50 9680 60
rect 9740 140 9770 150
rect 9740 60 9745 140
rect 9765 60 9770 140
rect 9740 50 9770 60
rect 9830 140 9860 150
rect 9830 60 9835 140
rect 9855 60 9860 140
rect 9830 50 9860 60
rect 9920 140 9950 150
rect 9920 60 9925 140
rect 9945 60 9950 140
rect 9920 50 9950 60
rect 10010 140 10040 150
rect 10010 60 10015 140
rect 10035 60 10040 140
rect 10010 50 10040 60
rect 10100 140 10130 150
rect 10100 60 10105 140
rect 10125 60 10130 140
rect 10100 50 10130 60
rect 10190 140 10220 150
rect 10190 60 10195 140
rect 10215 60 10220 140
rect 10190 50 10220 60
rect 10280 140 10310 150
rect 10280 60 10285 140
rect 10305 60 10310 140
rect 10280 50 10310 60
rect 10370 140 10400 150
rect 10370 60 10375 140
rect 10395 60 10400 140
rect 10370 50 10400 60
rect 10460 140 10490 150
rect 10460 60 10465 140
rect 10485 60 10490 140
rect 10460 50 10490 60
rect 10550 140 10580 150
rect 10550 60 10555 140
rect 10575 60 10580 140
rect 10550 50 10580 60
rect 10640 140 10670 150
rect 10640 60 10645 140
rect 10665 60 10670 140
rect 10640 50 10670 60
rect 10730 50 10760 150
rect 10820 50 10850 150
rect 10910 50 10940 150
rect 11000 50 11030 150
rect 11090 50 11120 150
rect 11180 140 11210 150
rect 11180 60 11185 140
rect 11205 60 11210 140
rect 11180 50 11210 60
rect -340 30 -320 50
rect 200 30 220 50
rect 380 30 400 50
rect 1820 30 1840 50
rect 3260 30 3280 50
rect 4700 30 4720 50
rect 4880 30 4900 50
rect 6320 30 6340 50
rect 7760 30 7780 50
rect 9205 30 9225 50
rect 9925 30 9945 50
rect 10645 30 10665 50
rect 11185 30 11205 50
rect -485 -5 -480 25
rect -450 -5 -445 25
rect -485 -10 -445 -5
rect -350 25 -310 30
rect -350 -5 -345 25
rect -315 0 -310 25
rect 190 25 230 30
rect -350 -10 -315 -5
rect 190 -5 195 25
rect 225 0 230 25
rect 370 25 410 30
rect 190 -10 225 -5
rect 370 -5 375 25
rect 405 -5 410 25
rect 370 -10 410 -5
rect 550 25 590 30
rect 550 -5 555 25
rect 585 -5 590 25
rect 550 -10 590 -5
rect 730 25 770 30
rect 730 -5 735 25
rect 765 -5 770 25
rect 730 -10 770 -5
rect 910 25 950 30
rect 910 -5 915 25
rect 945 -5 950 25
rect 910 -10 950 -5
rect 1090 25 1130 30
rect 1090 -5 1095 25
rect 1125 -5 1130 25
rect 1090 -10 1130 -5
rect 1270 25 1310 30
rect 1270 -5 1275 25
rect 1305 -5 1310 25
rect 1270 -10 1310 -5
rect 1450 25 1490 30
rect 1450 -5 1455 25
rect 1485 -5 1490 25
rect 1450 -10 1490 -5
rect 1630 25 1670 30
rect 1630 -5 1635 25
rect 1665 -5 1670 25
rect 1630 -10 1670 -5
rect 1810 25 1850 30
rect 1810 -5 1815 25
rect 1845 -5 1850 25
rect 1810 -10 1850 -5
rect 1990 25 2030 30
rect 1990 -5 1995 25
rect 2025 -5 2030 25
rect 1990 -10 2030 -5
rect 2170 25 2210 30
rect 2170 -5 2175 25
rect 2205 -5 2210 25
rect 2170 -10 2210 -5
rect 2350 25 2390 30
rect 2350 -5 2355 25
rect 2385 -5 2390 25
rect 2350 -10 2390 -5
rect 2530 25 2570 30
rect 2530 -5 2535 25
rect 2565 -5 2570 25
rect 2530 -10 2570 -5
rect 2710 25 2750 30
rect 2710 -5 2715 25
rect 2745 -5 2750 25
rect 2710 -10 2750 -5
rect 2890 25 2930 30
rect 2890 -5 2895 25
rect 2925 -5 2930 25
rect 2890 -10 2930 -5
rect 3070 25 3110 30
rect 3070 -5 3075 25
rect 3105 -5 3110 25
rect 3070 -10 3110 -5
rect 3250 25 3290 30
rect 3250 -5 3255 25
rect 3285 -5 3290 25
rect 3250 -10 3290 -5
rect 3430 25 3470 30
rect 3430 -5 3435 25
rect 3465 -5 3470 25
rect 3430 -10 3470 -5
rect 3610 25 3650 30
rect 3610 -5 3615 25
rect 3645 -5 3650 25
rect 3610 -10 3650 -5
rect 3790 25 3830 30
rect 3790 -5 3795 25
rect 3825 -5 3830 25
rect 3790 -10 3830 -5
rect 3970 25 4010 30
rect 3970 -5 3975 25
rect 4005 -5 4010 25
rect 3970 -10 4010 -5
rect 4150 25 4190 30
rect 4150 -5 4155 25
rect 4185 -5 4190 25
rect 4150 -10 4190 -5
rect 4330 25 4370 30
rect 4330 -5 4335 25
rect 4365 -5 4370 25
rect 4330 -10 4370 -5
rect 4510 25 4550 30
rect 4510 -5 4515 25
rect 4545 -5 4550 25
rect 4510 -10 4550 -5
rect 4690 25 4730 30
rect 4690 -5 4695 25
rect 4725 -5 4730 25
rect 4690 -10 4730 -5
rect 4870 25 4910 30
rect 4870 -5 4875 25
rect 4905 -5 4910 25
rect 4870 -10 4910 -5
rect 5050 25 5090 30
rect 5050 -5 5055 25
rect 5085 -5 5090 25
rect 5050 -10 5090 -5
rect 5230 25 5270 30
rect 5230 -5 5235 25
rect 5265 -5 5270 25
rect 5230 -10 5270 -5
rect 5410 25 5450 30
rect 5410 -5 5415 25
rect 5445 -5 5450 25
rect 5410 -10 5450 -5
rect 5590 25 5630 30
rect 5590 -5 5595 25
rect 5625 -5 5630 25
rect 5590 -10 5630 -5
rect 5770 25 5810 30
rect 5770 -5 5775 25
rect 5805 -5 5810 25
rect 5770 -10 5810 -5
rect 5950 25 5990 30
rect 5950 -5 5955 25
rect 5985 -5 5990 25
rect 5950 -10 5990 -5
rect 6130 25 6170 30
rect 6130 -5 6135 25
rect 6165 -5 6170 25
rect 6130 -10 6170 -5
rect 6310 25 6350 30
rect 6310 -5 6315 25
rect 6345 -5 6350 25
rect 6310 -10 6350 -5
rect 6490 25 6530 30
rect 6490 -5 6495 25
rect 6525 -5 6530 25
rect 6490 -10 6530 -5
rect 6670 25 6710 30
rect 6670 -5 6675 25
rect 6705 -5 6710 25
rect 6670 -10 6710 -5
rect 6850 25 6890 30
rect 6850 -5 6855 25
rect 6885 -5 6890 25
rect 6850 -10 6890 -5
rect 7030 25 7070 30
rect 7030 -5 7035 25
rect 7065 -5 7070 25
rect 7030 -10 7070 -5
rect 7210 25 7250 30
rect 7210 -5 7215 25
rect 7245 -5 7250 25
rect 7210 -10 7250 -5
rect 7390 25 7430 30
rect 7390 -5 7395 25
rect 7425 -5 7430 25
rect 7390 -10 7430 -5
rect 7570 25 7610 30
rect 7570 -5 7575 25
rect 7605 -5 7610 25
rect 7570 -10 7610 -5
rect 7750 25 7795 30
rect 7750 -5 7755 25
rect 7785 -5 7795 25
rect 7750 -10 7795 -5
rect 7935 25 7975 30
rect 7935 -5 7940 25
rect 7970 -5 7975 25
rect 7935 -10 7975 -5
rect 8115 25 8155 30
rect 8115 -5 8120 25
rect 8150 -5 8155 25
rect 8115 -10 8155 -5
rect 8295 25 8335 30
rect 8295 -5 8300 25
rect 8330 -5 8335 25
rect 8295 -10 8335 -5
rect 8475 25 8515 30
rect 8475 -5 8480 25
rect 8510 -5 8515 25
rect 8475 -10 8515 -5
rect 8655 25 8695 30
rect 8655 -5 8660 25
rect 8690 -5 8695 25
rect 8655 -10 8695 -5
rect 8835 25 8875 30
rect 8835 -5 8840 25
rect 8870 -5 8875 25
rect 8835 -10 8875 -5
rect 9015 25 9055 30
rect 9015 -5 9020 25
rect 9050 -5 9055 25
rect 9015 -10 9055 -5
rect 9195 25 9235 30
rect 9195 -5 9200 25
rect 9230 -5 9235 25
rect 9195 -10 9235 -5
rect 9375 25 9415 30
rect 9375 -5 9380 25
rect 9410 -5 9415 25
rect 9375 -10 9415 -5
rect 9555 25 9595 30
rect 9555 -5 9560 25
rect 9590 -5 9595 25
rect 9555 -10 9595 -5
rect 9735 25 9775 30
rect 9735 -5 9740 25
rect 9770 -5 9775 25
rect 9735 -10 9775 -5
rect 9915 25 9955 30
rect 9915 -5 9920 25
rect 9950 -5 9955 25
rect 9915 -10 9955 -5
rect 10095 25 10135 30
rect 10095 -5 10100 25
rect 10130 -5 10135 25
rect 10095 -10 10135 -5
rect 10275 25 10315 30
rect 10275 -5 10280 25
rect 10310 -5 10315 25
rect 10275 -10 10315 -5
rect 10455 25 10495 30
rect 10455 -5 10460 25
rect 10490 -5 10495 25
rect 10455 -10 10495 -5
rect 10635 25 10675 30
rect 10635 -5 10640 25
rect 10670 -5 10675 25
rect 10635 -10 10675 -5
rect 11175 25 11215 30
rect 11175 -5 11180 25
rect 11210 -5 11215 25
rect 11175 -10 11215 -5
rect 11310 25 11350 1810
rect 11310 -5 11315 25
rect 11345 -5 11350 25
rect 11310 -10 11350 -5
<< via1 >>
rect -480 1840 -450 1845
rect -480 1820 -475 1840
rect -475 1820 -455 1840
rect -455 1820 -450 1840
rect -480 1815 -450 1820
rect -345 1840 -315 1845
rect -345 1820 -340 1840
rect -340 1820 -320 1840
rect -320 1820 -315 1840
rect -345 1815 -315 1820
rect 195 1840 225 1845
rect 195 1820 200 1840
rect 200 1820 220 1840
rect 220 1820 225 1840
rect 195 1815 225 1820
rect 375 1840 405 1845
rect 375 1820 380 1840
rect 380 1820 400 1840
rect 400 1820 405 1840
rect 375 1815 405 1820
rect 555 1840 585 1845
rect 555 1820 560 1840
rect 560 1820 580 1840
rect 580 1820 585 1840
rect 555 1815 585 1820
rect 735 1840 765 1845
rect 735 1820 740 1840
rect 740 1820 760 1840
rect 760 1820 765 1840
rect 735 1815 765 1820
rect 915 1840 945 1845
rect 915 1820 920 1840
rect 920 1820 940 1840
rect 940 1820 945 1840
rect 915 1815 945 1820
rect 1095 1840 1125 1845
rect 1095 1820 1100 1840
rect 1100 1820 1120 1840
rect 1120 1820 1125 1840
rect 1095 1815 1125 1820
rect 1275 1840 1305 1845
rect 1275 1820 1280 1840
rect 1280 1820 1300 1840
rect 1300 1820 1305 1840
rect 1275 1815 1305 1820
rect 1455 1840 1485 1845
rect 1455 1820 1460 1840
rect 1460 1820 1480 1840
rect 1480 1820 1485 1840
rect 1455 1815 1485 1820
rect 1635 1840 1665 1845
rect 1635 1820 1640 1840
rect 1640 1820 1660 1840
rect 1660 1820 1665 1840
rect 1635 1815 1665 1820
rect 1815 1840 1845 1845
rect 1815 1820 1820 1840
rect 1820 1820 1840 1840
rect 1840 1820 1845 1840
rect 1815 1815 1845 1820
rect 1995 1840 2025 1845
rect 1995 1820 2000 1840
rect 2000 1820 2020 1840
rect 2020 1820 2025 1840
rect 1995 1815 2025 1820
rect 2175 1840 2205 1845
rect 2175 1820 2180 1840
rect 2180 1820 2200 1840
rect 2200 1820 2205 1840
rect 2175 1815 2205 1820
rect 2355 1840 2385 1845
rect 2355 1820 2360 1840
rect 2360 1820 2380 1840
rect 2380 1820 2385 1840
rect 2355 1815 2385 1820
rect 2535 1840 2565 1845
rect 2535 1820 2540 1840
rect 2540 1820 2560 1840
rect 2560 1820 2565 1840
rect 2535 1815 2565 1820
rect 2715 1840 2745 1845
rect 2715 1820 2720 1840
rect 2720 1820 2740 1840
rect 2740 1820 2745 1840
rect 2715 1815 2745 1820
rect 2895 1840 2925 1845
rect 2895 1820 2900 1840
rect 2900 1820 2920 1840
rect 2920 1820 2925 1840
rect 2895 1815 2925 1820
rect 3080 1840 3110 1845
rect 3080 1820 3085 1840
rect 3085 1820 3105 1840
rect 3105 1820 3110 1840
rect 3080 1815 3110 1820
rect 3260 1840 3290 1845
rect 3260 1820 3265 1840
rect 3265 1820 3285 1840
rect 3285 1820 3290 1840
rect 3260 1815 3290 1820
rect 3440 1840 3470 1845
rect 3440 1820 3445 1840
rect 3445 1820 3465 1840
rect 3465 1820 3470 1840
rect 3440 1815 3470 1820
rect 3620 1840 3650 1845
rect 3620 1820 3625 1840
rect 3625 1820 3645 1840
rect 3645 1820 3650 1840
rect 3620 1815 3650 1820
rect 3800 1840 3830 1845
rect 3800 1820 3805 1840
rect 3805 1820 3825 1840
rect 3825 1820 3830 1840
rect 3800 1815 3830 1820
rect 3980 1840 4010 1845
rect 3980 1820 3985 1840
rect 3985 1820 4005 1840
rect 4005 1820 4010 1840
rect 3980 1815 4010 1820
rect 4160 1840 4190 1845
rect 4160 1820 4165 1840
rect 4165 1820 4185 1840
rect 4185 1820 4190 1840
rect 4160 1815 4190 1820
rect 4340 1840 4370 1845
rect 4340 1820 4345 1840
rect 4345 1820 4365 1840
rect 4365 1820 4370 1840
rect 4340 1815 4370 1820
rect 4520 1840 4550 1845
rect 4520 1820 4525 1840
rect 4525 1820 4545 1840
rect 4545 1820 4550 1840
rect 4520 1815 4550 1820
rect 4700 1840 4730 1845
rect 4700 1820 4705 1840
rect 4705 1820 4725 1840
rect 4725 1820 4730 1840
rect 4700 1815 4730 1820
rect 4880 1840 4910 1845
rect 4880 1820 4885 1840
rect 4885 1820 4905 1840
rect 4905 1820 4910 1840
rect 4880 1815 4910 1820
rect 5060 1840 5090 1845
rect 5060 1820 5065 1840
rect 5065 1820 5085 1840
rect 5085 1820 5090 1840
rect 5060 1815 5090 1820
rect 5240 1840 5270 1845
rect 5240 1820 5245 1840
rect 5245 1820 5265 1840
rect 5265 1820 5270 1840
rect 5240 1815 5270 1820
rect 5420 1840 5450 1845
rect 5420 1820 5425 1840
rect 5425 1820 5445 1840
rect 5445 1820 5450 1840
rect 5420 1815 5450 1820
rect 5600 1840 5630 1845
rect 5600 1820 5605 1840
rect 5605 1820 5625 1840
rect 5625 1820 5630 1840
rect 5600 1815 5630 1820
rect 5780 1840 5810 1845
rect 5780 1820 5785 1840
rect 5785 1820 5805 1840
rect 5805 1820 5810 1840
rect 5780 1815 5810 1820
rect 5960 1840 5990 1845
rect 5960 1820 5965 1840
rect 5965 1820 5985 1840
rect 5985 1820 5990 1840
rect 5960 1815 5990 1820
rect 6140 1840 6170 1845
rect 6140 1820 6145 1840
rect 6145 1820 6165 1840
rect 6165 1820 6170 1840
rect 6140 1815 6170 1820
rect 6320 1840 6350 1845
rect 6320 1820 6325 1840
rect 6325 1820 6345 1840
rect 6345 1820 6350 1840
rect 6320 1815 6350 1820
rect 6500 1840 6530 1845
rect 6500 1820 6505 1840
rect 6505 1820 6525 1840
rect 6525 1820 6530 1840
rect 6500 1815 6530 1820
rect 6680 1840 6710 1845
rect 6680 1820 6685 1840
rect 6685 1820 6705 1840
rect 6705 1820 6710 1840
rect 6680 1815 6710 1820
rect 6860 1840 6890 1845
rect 6860 1820 6865 1840
rect 6865 1820 6885 1840
rect 6885 1820 6890 1840
rect 6860 1815 6890 1820
rect 7040 1840 7070 1845
rect 7040 1820 7045 1840
rect 7045 1820 7065 1840
rect 7065 1820 7070 1840
rect 7040 1815 7070 1820
rect 7220 1840 7250 1845
rect 7220 1820 7225 1840
rect 7225 1820 7245 1840
rect 7245 1820 7250 1840
rect 7220 1815 7250 1820
rect 7400 1840 7430 1845
rect 7400 1820 7405 1840
rect 7405 1820 7425 1840
rect 7425 1820 7430 1840
rect 7400 1815 7430 1820
rect 7580 1840 7610 1845
rect 7580 1820 7585 1840
rect 7585 1820 7605 1840
rect 7605 1820 7610 1840
rect 7580 1815 7610 1820
rect 7760 1840 7790 1845
rect 7760 1820 7765 1840
rect 7765 1820 7785 1840
rect 7785 1820 7790 1840
rect 7760 1815 7790 1820
rect 7940 1840 7970 1845
rect 7940 1820 7945 1840
rect 7945 1820 7965 1840
rect 7965 1820 7970 1840
rect 7940 1815 7970 1820
rect 8120 1840 8150 1845
rect 8120 1820 8125 1840
rect 8125 1820 8145 1840
rect 8145 1820 8150 1840
rect 8120 1815 8150 1820
rect 8300 1840 8330 1845
rect 8300 1820 8305 1840
rect 8305 1820 8325 1840
rect 8325 1820 8330 1840
rect 8300 1815 8330 1820
rect 8480 1840 8510 1845
rect 8480 1820 8485 1840
rect 8485 1820 8505 1840
rect 8505 1820 8510 1840
rect 8480 1815 8510 1820
rect 8660 1840 8690 1845
rect 8660 1820 8665 1840
rect 8665 1820 8685 1840
rect 8685 1820 8690 1840
rect 8660 1815 8690 1820
rect 8840 1840 8870 1845
rect 8840 1820 8845 1840
rect 8845 1820 8865 1840
rect 8865 1820 8870 1840
rect 8840 1815 8870 1820
rect 9020 1840 9050 1845
rect 9020 1820 9025 1840
rect 9025 1820 9045 1840
rect 9045 1820 9050 1840
rect 9020 1815 9050 1820
rect 9200 1840 9230 1845
rect 9200 1820 9205 1840
rect 9205 1820 9225 1840
rect 9225 1820 9230 1840
rect 9200 1815 9230 1820
rect 9380 1840 9410 1845
rect 9380 1820 9385 1840
rect 9385 1820 9405 1840
rect 9405 1820 9410 1840
rect 9380 1815 9410 1820
rect 9560 1840 9590 1845
rect 9560 1820 9565 1840
rect 9565 1820 9585 1840
rect 9585 1820 9590 1840
rect 9560 1815 9590 1820
rect 9740 1840 9770 1845
rect 9740 1820 9745 1840
rect 9745 1820 9765 1840
rect 9765 1820 9770 1840
rect 9740 1815 9770 1820
rect 9920 1840 9950 1845
rect 9920 1820 9925 1840
rect 9925 1820 9945 1840
rect 9945 1820 9950 1840
rect 9920 1815 9950 1820
rect 10100 1840 10130 1845
rect 10100 1820 10105 1840
rect 10105 1820 10125 1840
rect 10125 1820 10130 1840
rect 10100 1815 10130 1820
rect 10280 1840 10310 1845
rect 10280 1820 10285 1840
rect 10285 1820 10305 1840
rect 10305 1820 10310 1840
rect 10280 1815 10310 1820
rect 10460 1840 10490 1845
rect 10460 1820 10465 1840
rect 10465 1820 10485 1840
rect 10485 1820 10490 1840
rect 10460 1815 10490 1820
rect 10640 1840 10670 1845
rect 10640 1820 10645 1840
rect 10645 1820 10665 1840
rect 10665 1820 10670 1840
rect 10640 1815 10670 1820
rect 11180 1840 11210 1845
rect 11180 1820 11185 1840
rect 11185 1820 11205 1840
rect 11205 1820 11210 1840
rect 11180 1815 11210 1820
rect 11315 1840 11345 1845
rect 11315 1820 11320 1840
rect 11320 1820 11340 1840
rect 11340 1820 11345 1840
rect 11315 1815 11345 1820
rect -345 960 -315 965
rect -345 940 -340 960
rect -340 940 -320 960
rect -320 940 -315 960
rect -345 935 -315 940
rect -345 900 -315 905
rect -345 880 -340 900
rect -340 880 -320 900
rect -320 880 -315 900
rect -345 875 -315 880
rect 195 960 225 965
rect 195 940 200 960
rect 200 940 220 960
rect 220 940 225 960
rect 195 935 225 940
rect 375 960 405 965
rect 375 940 380 960
rect 380 940 400 960
rect 400 940 405 960
rect 375 935 405 940
rect 555 960 585 965
rect 555 940 560 960
rect 560 940 580 960
rect 580 940 585 960
rect 555 935 585 940
rect 735 960 765 965
rect 735 940 740 960
rect 740 940 760 960
rect 760 940 765 960
rect 735 935 765 940
rect 915 960 945 965
rect 915 940 920 960
rect 920 940 940 960
rect 940 940 945 960
rect 915 935 945 940
rect 1095 960 1125 965
rect 1095 940 1100 960
rect 1100 940 1120 960
rect 1120 940 1125 960
rect 1095 935 1125 940
rect 1275 960 1305 965
rect 1275 940 1280 960
rect 1280 940 1300 960
rect 1300 940 1305 960
rect 1275 935 1305 940
rect 1455 960 1485 965
rect 1455 940 1460 960
rect 1460 940 1480 960
rect 1480 940 1485 960
rect 1455 935 1485 940
rect 1635 960 1665 965
rect 1635 940 1640 960
rect 1640 940 1660 960
rect 1660 940 1665 960
rect 1635 935 1665 940
rect 1815 960 1845 965
rect 1815 940 1820 960
rect 1820 940 1840 960
rect 1840 940 1845 960
rect 1815 935 1845 940
rect 1995 960 2025 965
rect 1995 940 2000 960
rect 2000 940 2020 960
rect 2020 940 2025 960
rect 1995 935 2025 940
rect 2175 960 2205 965
rect 2175 940 2180 960
rect 2180 940 2200 960
rect 2200 940 2205 960
rect 2175 935 2205 940
rect 2355 960 2385 965
rect 2355 940 2360 960
rect 2360 940 2380 960
rect 2380 940 2385 960
rect 2355 935 2385 940
rect 2535 960 2565 965
rect 2535 940 2540 960
rect 2540 940 2560 960
rect 2560 940 2565 960
rect 2535 935 2565 940
rect 2715 960 2745 965
rect 2715 940 2720 960
rect 2720 940 2740 960
rect 2740 940 2745 960
rect 2715 935 2745 940
rect 2895 960 2925 965
rect 2895 940 2900 960
rect 2900 940 2920 960
rect 2920 940 2925 960
rect 2895 935 2925 940
rect 3080 960 3110 965
rect 3080 940 3085 960
rect 3085 940 3105 960
rect 3105 940 3110 960
rect 3080 935 3110 940
rect 3260 960 3290 965
rect 3260 940 3265 960
rect 3265 940 3285 960
rect 3285 940 3290 960
rect 3260 935 3290 940
rect 3440 960 3470 965
rect 3440 940 3445 960
rect 3445 940 3465 960
rect 3465 940 3470 960
rect 3440 935 3470 940
rect 3620 960 3650 965
rect 3620 940 3625 960
rect 3625 940 3645 960
rect 3645 940 3650 960
rect 3620 935 3650 940
rect 3800 960 3830 965
rect 3800 940 3805 960
rect 3805 940 3825 960
rect 3825 940 3830 960
rect 3800 935 3830 940
rect 3980 960 4010 965
rect 3980 940 3985 960
rect 3985 940 4005 960
rect 4005 940 4010 960
rect 3980 935 4010 940
rect 4160 960 4190 965
rect 4160 940 4165 960
rect 4165 940 4185 960
rect 4185 940 4190 960
rect 4160 935 4190 940
rect 4340 960 4370 965
rect 4340 940 4345 960
rect 4345 940 4365 960
rect 4365 940 4370 960
rect 4340 935 4370 940
rect 4520 960 4550 965
rect 4520 940 4525 960
rect 4525 940 4545 960
rect 4545 940 4550 960
rect 4520 935 4550 940
rect 4700 960 4730 965
rect 4700 940 4705 960
rect 4705 940 4725 960
rect 4725 940 4730 960
rect 4700 935 4730 940
rect 4880 960 4910 965
rect 4880 940 4885 960
rect 4885 940 4905 960
rect 4905 940 4910 960
rect 4880 935 4910 940
rect 5060 960 5090 965
rect 5060 940 5065 960
rect 5065 940 5085 960
rect 5085 940 5090 960
rect 5060 935 5090 940
rect 5240 960 5270 965
rect 5240 940 5245 960
rect 5245 940 5265 960
rect 5265 940 5270 960
rect 5240 935 5270 940
rect 5420 960 5450 965
rect 5420 940 5425 960
rect 5425 940 5445 960
rect 5445 940 5450 960
rect 5420 935 5450 940
rect 5600 960 5630 965
rect 5600 940 5605 960
rect 5605 940 5625 960
rect 5625 940 5630 960
rect 5600 935 5630 940
rect 5780 960 5810 965
rect 5780 940 5785 960
rect 5785 940 5805 960
rect 5805 940 5810 960
rect 5780 935 5810 940
rect 5960 960 5990 965
rect 5960 940 5965 960
rect 5965 940 5985 960
rect 5985 940 5990 960
rect 5960 935 5990 940
rect 6140 960 6170 965
rect 6140 940 6145 960
rect 6145 940 6165 960
rect 6165 940 6170 960
rect 6140 935 6170 940
rect 6320 960 6350 965
rect 6320 940 6325 960
rect 6325 940 6345 960
rect 6345 940 6350 960
rect 6320 935 6350 940
rect 6500 960 6530 965
rect 6500 940 6505 960
rect 6505 940 6525 960
rect 6525 940 6530 960
rect 6500 935 6530 940
rect 6680 960 6710 965
rect 6680 940 6685 960
rect 6685 940 6705 960
rect 6705 940 6710 960
rect 6680 935 6710 940
rect 6860 960 6890 965
rect 6860 940 6865 960
rect 6865 940 6885 960
rect 6885 940 6890 960
rect 6860 935 6890 940
rect 7040 960 7070 965
rect 7040 940 7045 960
rect 7045 940 7065 960
rect 7065 940 7070 960
rect 7040 935 7070 940
rect 7220 960 7250 965
rect 7220 940 7225 960
rect 7225 940 7245 960
rect 7245 940 7250 960
rect 7220 935 7250 940
rect 7400 960 7430 965
rect 7400 940 7405 960
rect 7405 940 7425 960
rect 7425 940 7430 960
rect 7400 935 7430 940
rect 7580 960 7610 965
rect 7580 940 7585 960
rect 7585 940 7605 960
rect 7605 940 7610 960
rect 7580 935 7610 940
rect 7760 960 7790 965
rect 7760 940 7765 960
rect 7765 940 7785 960
rect 7785 940 7790 960
rect 7760 935 7790 940
rect 7940 960 7970 965
rect 7940 940 7945 960
rect 7945 940 7965 960
rect 7965 940 7970 960
rect 7940 935 7970 940
rect 8120 960 8150 965
rect 8120 940 8125 960
rect 8125 940 8145 960
rect 8145 940 8150 960
rect 8120 935 8150 940
rect 8300 960 8330 965
rect 8300 940 8305 960
rect 8305 940 8325 960
rect 8325 940 8330 960
rect 8300 935 8330 940
rect 8480 960 8510 965
rect 8480 940 8485 960
rect 8485 940 8505 960
rect 8505 940 8510 960
rect 8480 935 8510 940
rect 8660 960 8690 965
rect 8660 940 8665 960
rect 8665 940 8685 960
rect 8685 940 8690 960
rect 8660 935 8690 940
rect 8840 960 8870 965
rect 8840 940 8845 960
rect 8845 940 8865 960
rect 8865 940 8870 960
rect 8840 935 8870 940
rect 9020 960 9050 965
rect 9020 940 9025 960
rect 9025 940 9045 960
rect 9045 940 9050 960
rect 9020 935 9050 940
rect 9200 960 9230 965
rect 9200 940 9205 960
rect 9205 940 9225 960
rect 9225 940 9230 960
rect 9200 935 9230 940
rect 9380 960 9410 965
rect 9380 940 9385 960
rect 9385 940 9405 960
rect 9405 940 9410 960
rect 9380 935 9410 940
rect 9560 960 9590 965
rect 9560 940 9565 960
rect 9565 940 9585 960
rect 9585 940 9590 960
rect 9560 935 9590 940
rect 9740 960 9770 965
rect 9740 940 9745 960
rect 9745 940 9765 960
rect 9765 940 9770 960
rect 9740 935 9770 940
rect 9920 960 9950 965
rect 9920 940 9925 960
rect 9925 940 9945 960
rect 9945 940 9950 960
rect 9920 935 9950 940
rect 10100 960 10130 965
rect 10100 940 10105 960
rect 10105 940 10125 960
rect 10125 940 10130 960
rect 10100 935 10130 940
rect 10280 960 10310 965
rect 10280 940 10285 960
rect 10285 940 10305 960
rect 10305 940 10310 960
rect 10280 935 10310 940
rect 10460 960 10490 965
rect 10460 940 10465 960
rect 10465 940 10485 960
rect 10485 940 10490 960
rect 10460 935 10490 940
rect 10640 960 10670 965
rect 10640 940 10645 960
rect 10645 940 10665 960
rect 10665 940 10670 960
rect 10640 935 10670 940
rect 195 900 225 905
rect 195 880 200 900
rect 200 880 220 900
rect 220 880 225 900
rect 195 875 225 880
rect 375 900 405 905
rect 375 880 380 900
rect 380 880 400 900
rect 400 880 405 900
rect 375 875 405 880
rect 555 900 585 905
rect 555 880 560 900
rect 560 880 580 900
rect 580 880 585 900
rect 555 875 585 880
rect 735 900 765 905
rect 735 880 740 900
rect 740 880 760 900
rect 760 880 765 900
rect 735 875 765 880
rect 915 900 945 905
rect 915 880 920 900
rect 920 880 940 900
rect 940 880 945 900
rect 915 875 945 880
rect 1095 900 1125 905
rect 1095 880 1100 900
rect 1100 880 1120 900
rect 1120 880 1125 900
rect 1095 875 1125 880
rect 1275 900 1305 905
rect 1275 880 1280 900
rect 1280 880 1300 900
rect 1300 880 1305 900
rect 1275 875 1305 880
rect 1455 900 1485 905
rect 1455 880 1460 900
rect 1460 880 1480 900
rect 1480 880 1485 900
rect 1455 875 1485 880
rect 1635 900 1665 905
rect 1635 880 1640 900
rect 1640 880 1660 900
rect 1660 880 1665 900
rect 1635 875 1665 880
rect 1815 900 1845 905
rect 1815 880 1820 900
rect 1820 880 1840 900
rect 1840 880 1845 900
rect 1815 875 1845 880
rect 1995 900 2025 905
rect 1995 880 2000 900
rect 2000 880 2020 900
rect 2020 880 2025 900
rect 1995 875 2025 880
rect 2175 900 2205 905
rect 2175 880 2180 900
rect 2180 880 2200 900
rect 2200 880 2205 900
rect 2175 875 2205 880
rect 2355 900 2385 905
rect 2355 880 2360 900
rect 2360 880 2380 900
rect 2380 880 2385 900
rect 2355 875 2385 880
rect 2535 900 2565 905
rect 2535 880 2540 900
rect 2540 880 2560 900
rect 2560 880 2565 900
rect 2535 875 2565 880
rect 2715 900 2745 905
rect 2715 880 2720 900
rect 2720 880 2740 900
rect 2740 880 2745 900
rect 2715 875 2745 880
rect 2895 900 2925 905
rect 2895 880 2900 900
rect 2900 880 2920 900
rect 2920 880 2925 900
rect 2895 875 2925 880
rect 3075 900 3105 905
rect 3075 880 3080 900
rect 3080 880 3100 900
rect 3100 880 3105 900
rect 3075 875 3105 880
rect 3255 900 3285 905
rect 3255 880 3260 900
rect 3260 880 3280 900
rect 3280 880 3285 900
rect 3255 875 3285 880
rect 3435 900 3465 905
rect 3435 880 3440 900
rect 3440 880 3460 900
rect 3460 880 3465 900
rect 3435 875 3465 880
rect 3615 900 3645 905
rect 3615 880 3620 900
rect 3620 880 3640 900
rect 3640 880 3645 900
rect 3615 875 3645 880
rect 3795 900 3825 905
rect 3795 880 3800 900
rect 3800 880 3820 900
rect 3820 880 3825 900
rect 3795 875 3825 880
rect 3975 900 4005 905
rect 3975 880 3980 900
rect 3980 880 4000 900
rect 4000 880 4005 900
rect 3975 875 4005 880
rect 4155 900 4185 905
rect 4155 880 4160 900
rect 4160 880 4180 900
rect 4180 880 4185 900
rect 4155 875 4185 880
rect 4335 900 4365 905
rect 4335 880 4340 900
rect 4340 880 4360 900
rect 4360 880 4365 900
rect 4335 875 4365 880
rect 4515 900 4545 905
rect 4515 880 4520 900
rect 4520 880 4540 900
rect 4540 880 4545 900
rect 4515 875 4545 880
rect 4695 900 4725 905
rect 4695 880 4700 900
rect 4700 880 4720 900
rect 4720 880 4725 900
rect 4695 875 4725 880
rect 4875 900 4905 905
rect 4875 880 4880 900
rect 4880 880 4900 900
rect 4900 880 4905 900
rect 4875 875 4905 880
rect 5055 900 5085 905
rect 5055 880 5060 900
rect 5060 880 5080 900
rect 5080 880 5085 900
rect 5055 875 5085 880
rect 5235 900 5265 905
rect 5235 880 5240 900
rect 5240 880 5260 900
rect 5260 880 5265 900
rect 5235 875 5265 880
rect 5415 900 5445 905
rect 5415 880 5420 900
rect 5420 880 5440 900
rect 5440 880 5445 900
rect 5415 875 5445 880
rect 5595 900 5625 905
rect 5595 880 5600 900
rect 5600 880 5620 900
rect 5620 880 5625 900
rect 5595 875 5625 880
rect 5775 900 5805 905
rect 5775 880 5780 900
rect 5780 880 5800 900
rect 5800 880 5805 900
rect 5775 875 5805 880
rect 5955 900 5985 905
rect 5955 880 5960 900
rect 5960 880 5980 900
rect 5980 880 5985 900
rect 5955 875 5985 880
rect 6135 900 6165 905
rect 6135 880 6140 900
rect 6140 880 6160 900
rect 6160 880 6165 900
rect 6135 875 6165 880
rect 6315 900 6345 905
rect 6315 880 6320 900
rect 6320 880 6340 900
rect 6340 880 6345 900
rect 6315 875 6345 880
rect 6495 900 6525 905
rect 6495 880 6500 900
rect 6500 880 6520 900
rect 6520 880 6525 900
rect 6495 875 6525 880
rect 6675 900 6705 905
rect 6675 880 6680 900
rect 6680 880 6700 900
rect 6700 880 6705 900
rect 6675 875 6705 880
rect 6855 900 6885 905
rect 6855 880 6860 900
rect 6860 880 6880 900
rect 6880 880 6885 900
rect 6855 875 6885 880
rect 7035 900 7065 905
rect 7035 880 7040 900
rect 7040 880 7060 900
rect 7060 880 7065 900
rect 7035 875 7065 880
rect 7215 900 7245 905
rect 7215 880 7220 900
rect 7220 880 7240 900
rect 7240 880 7245 900
rect 7215 875 7245 880
rect 7395 900 7425 905
rect 7395 880 7400 900
rect 7400 880 7420 900
rect 7420 880 7425 900
rect 7395 875 7425 880
rect 7575 900 7605 905
rect 7575 880 7580 900
rect 7580 880 7600 900
rect 7600 880 7605 900
rect 7575 875 7605 880
rect 7755 900 7785 905
rect 7755 880 7760 900
rect 7760 880 7780 900
rect 7780 880 7785 900
rect 7755 875 7785 880
rect 7940 900 7970 905
rect 7940 880 7945 900
rect 7945 880 7965 900
rect 7965 880 7970 900
rect 7940 875 7970 880
rect 8120 900 8150 905
rect 8120 880 8125 900
rect 8125 880 8145 900
rect 8145 880 8150 900
rect 8120 875 8150 880
rect 8300 900 8330 905
rect 8300 880 8305 900
rect 8305 880 8325 900
rect 8325 880 8330 900
rect 8300 875 8330 880
rect 8480 900 8510 905
rect 8480 880 8485 900
rect 8485 880 8505 900
rect 8505 880 8510 900
rect 8480 875 8510 880
rect 8660 900 8690 905
rect 8660 880 8665 900
rect 8665 880 8685 900
rect 8685 880 8690 900
rect 8660 875 8690 880
rect 8840 900 8870 905
rect 8840 880 8845 900
rect 8845 880 8865 900
rect 8865 880 8870 900
rect 8840 875 8870 880
rect 9020 900 9050 905
rect 9020 880 9025 900
rect 9025 880 9045 900
rect 9045 880 9050 900
rect 9020 875 9050 880
rect 9200 900 9230 905
rect 9200 880 9205 900
rect 9205 880 9225 900
rect 9225 880 9230 900
rect 9200 875 9230 880
rect 9380 900 9410 905
rect 9380 880 9385 900
rect 9385 880 9405 900
rect 9405 880 9410 900
rect 9380 875 9410 880
rect 9560 900 9590 905
rect 9560 880 9565 900
rect 9565 880 9585 900
rect 9585 880 9590 900
rect 9560 875 9590 880
rect 9740 900 9770 905
rect 9740 880 9745 900
rect 9745 880 9765 900
rect 9765 880 9770 900
rect 9740 875 9770 880
rect 9920 900 9950 905
rect 9920 880 9925 900
rect 9925 880 9945 900
rect 9945 880 9950 900
rect 9920 875 9950 880
rect 10100 900 10130 905
rect 10100 880 10105 900
rect 10105 880 10125 900
rect 10125 880 10130 900
rect 10100 875 10130 880
rect 10280 900 10310 905
rect 10280 880 10285 900
rect 10285 880 10305 900
rect 10305 880 10310 900
rect 10280 875 10310 880
rect 10460 900 10490 905
rect 10460 880 10465 900
rect 10465 880 10485 900
rect 10485 880 10490 900
rect 10460 875 10490 880
rect 10640 900 10670 905
rect 10640 880 10645 900
rect 10645 880 10665 900
rect 10665 880 10670 900
rect 10640 875 10670 880
rect 11180 960 11210 965
rect 11180 940 11185 960
rect 11185 940 11205 960
rect 11205 940 11210 960
rect 11180 935 11210 940
rect 11180 900 11210 905
rect 11180 880 11185 900
rect 11185 880 11205 900
rect 11205 880 11210 900
rect 11180 875 11210 880
rect -480 20 -450 25
rect -480 0 -475 20
rect -475 0 -455 20
rect -455 0 -450 20
rect -480 -5 -450 0
rect -345 20 -315 25
rect -345 0 -340 20
rect -340 0 -320 20
rect -320 0 -315 20
rect -345 -5 -315 0
rect 195 20 225 25
rect 195 0 200 20
rect 200 0 220 20
rect 220 0 225 20
rect 195 -5 225 0
rect 375 20 405 25
rect 375 0 380 20
rect 380 0 400 20
rect 400 0 405 20
rect 375 -5 405 0
rect 555 20 585 25
rect 555 0 560 20
rect 560 0 580 20
rect 580 0 585 20
rect 555 -5 585 0
rect 735 20 765 25
rect 735 0 740 20
rect 740 0 760 20
rect 760 0 765 20
rect 735 -5 765 0
rect 915 20 945 25
rect 915 0 920 20
rect 920 0 940 20
rect 940 0 945 20
rect 915 -5 945 0
rect 1095 20 1125 25
rect 1095 0 1100 20
rect 1100 0 1120 20
rect 1120 0 1125 20
rect 1095 -5 1125 0
rect 1275 20 1305 25
rect 1275 0 1280 20
rect 1280 0 1300 20
rect 1300 0 1305 20
rect 1275 -5 1305 0
rect 1455 20 1485 25
rect 1455 0 1460 20
rect 1460 0 1480 20
rect 1480 0 1485 20
rect 1455 -5 1485 0
rect 1635 20 1665 25
rect 1635 0 1640 20
rect 1640 0 1660 20
rect 1660 0 1665 20
rect 1635 -5 1665 0
rect 1815 20 1845 25
rect 1815 0 1820 20
rect 1820 0 1840 20
rect 1840 0 1845 20
rect 1815 -5 1845 0
rect 1995 20 2025 25
rect 1995 0 2000 20
rect 2000 0 2020 20
rect 2020 0 2025 20
rect 1995 -5 2025 0
rect 2175 20 2205 25
rect 2175 0 2180 20
rect 2180 0 2200 20
rect 2200 0 2205 20
rect 2175 -5 2205 0
rect 2355 20 2385 25
rect 2355 0 2360 20
rect 2360 0 2380 20
rect 2380 0 2385 20
rect 2355 -5 2385 0
rect 2535 20 2565 25
rect 2535 0 2540 20
rect 2540 0 2560 20
rect 2560 0 2565 20
rect 2535 -5 2565 0
rect 2715 20 2745 25
rect 2715 0 2720 20
rect 2720 0 2740 20
rect 2740 0 2745 20
rect 2715 -5 2745 0
rect 2895 20 2925 25
rect 2895 0 2900 20
rect 2900 0 2920 20
rect 2920 0 2925 20
rect 2895 -5 2925 0
rect 3075 20 3105 25
rect 3075 0 3080 20
rect 3080 0 3100 20
rect 3100 0 3105 20
rect 3075 -5 3105 0
rect 3255 20 3285 25
rect 3255 0 3260 20
rect 3260 0 3280 20
rect 3280 0 3285 20
rect 3255 -5 3285 0
rect 3435 20 3465 25
rect 3435 0 3440 20
rect 3440 0 3460 20
rect 3460 0 3465 20
rect 3435 -5 3465 0
rect 3615 20 3645 25
rect 3615 0 3620 20
rect 3620 0 3640 20
rect 3640 0 3645 20
rect 3615 -5 3645 0
rect 3795 20 3825 25
rect 3795 0 3800 20
rect 3800 0 3820 20
rect 3820 0 3825 20
rect 3795 -5 3825 0
rect 3975 20 4005 25
rect 3975 0 3980 20
rect 3980 0 4000 20
rect 4000 0 4005 20
rect 3975 -5 4005 0
rect 4155 20 4185 25
rect 4155 0 4160 20
rect 4160 0 4180 20
rect 4180 0 4185 20
rect 4155 -5 4185 0
rect 4335 20 4365 25
rect 4335 0 4340 20
rect 4340 0 4360 20
rect 4360 0 4365 20
rect 4335 -5 4365 0
rect 4515 20 4545 25
rect 4515 0 4520 20
rect 4520 0 4540 20
rect 4540 0 4545 20
rect 4515 -5 4545 0
rect 4695 20 4725 25
rect 4695 0 4700 20
rect 4700 0 4720 20
rect 4720 0 4725 20
rect 4695 -5 4725 0
rect 4875 20 4905 25
rect 4875 0 4880 20
rect 4880 0 4900 20
rect 4900 0 4905 20
rect 4875 -5 4905 0
rect 5055 20 5085 25
rect 5055 0 5060 20
rect 5060 0 5080 20
rect 5080 0 5085 20
rect 5055 -5 5085 0
rect 5235 20 5265 25
rect 5235 0 5240 20
rect 5240 0 5260 20
rect 5260 0 5265 20
rect 5235 -5 5265 0
rect 5415 20 5445 25
rect 5415 0 5420 20
rect 5420 0 5440 20
rect 5440 0 5445 20
rect 5415 -5 5445 0
rect 5595 20 5625 25
rect 5595 0 5600 20
rect 5600 0 5620 20
rect 5620 0 5625 20
rect 5595 -5 5625 0
rect 5775 20 5805 25
rect 5775 0 5780 20
rect 5780 0 5800 20
rect 5800 0 5805 20
rect 5775 -5 5805 0
rect 5955 20 5985 25
rect 5955 0 5960 20
rect 5960 0 5980 20
rect 5980 0 5985 20
rect 5955 -5 5985 0
rect 6135 20 6165 25
rect 6135 0 6140 20
rect 6140 0 6160 20
rect 6160 0 6165 20
rect 6135 -5 6165 0
rect 6315 20 6345 25
rect 6315 0 6320 20
rect 6320 0 6340 20
rect 6340 0 6345 20
rect 6315 -5 6345 0
rect 6495 20 6525 25
rect 6495 0 6500 20
rect 6500 0 6520 20
rect 6520 0 6525 20
rect 6495 -5 6525 0
rect 6675 20 6705 25
rect 6675 0 6680 20
rect 6680 0 6700 20
rect 6700 0 6705 20
rect 6675 -5 6705 0
rect 6855 20 6885 25
rect 6855 0 6860 20
rect 6860 0 6880 20
rect 6880 0 6885 20
rect 6855 -5 6885 0
rect 7035 20 7065 25
rect 7035 0 7040 20
rect 7040 0 7060 20
rect 7060 0 7065 20
rect 7035 -5 7065 0
rect 7215 20 7245 25
rect 7215 0 7220 20
rect 7220 0 7240 20
rect 7240 0 7245 20
rect 7215 -5 7245 0
rect 7395 20 7425 25
rect 7395 0 7400 20
rect 7400 0 7420 20
rect 7420 0 7425 20
rect 7395 -5 7425 0
rect 7575 20 7605 25
rect 7575 0 7580 20
rect 7580 0 7600 20
rect 7600 0 7605 20
rect 7575 -5 7605 0
rect 7755 20 7785 25
rect 7755 0 7760 20
rect 7760 0 7780 20
rect 7780 0 7785 20
rect 7755 -5 7785 0
rect 7940 20 7970 25
rect 7940 0 7945 20
rect 7945 0 7965 20
rect 7965 0 7970 20
rect 7940 -5 7970 0
rect 8120 20 8150 25
rect 8120 0 8125 20
rect 8125 0 8145 20
rect 8145 0 8150 20
rect 8120 -5 8150 0
rect 8300 20 8330 25
rect 8300 0 8305 20
rect 8305 0 8325 20
rect 8325 0 8330 20
rect 8300 -5 8330 0
rect 8480 20 8510 25
rect 8480 0 8485 20
rect 8485 0 8505 20
rect 8505 0 8510 20
rect 8480 -5 8510 0
rect 8660 20 8690 25
rect 8660 0 8665 20
rect 8665 0 8685 20
rect 8685 0 8690 20
rect 8660 -5 8690 0
rect 8840 20 8870 25
rect 8840 0 8845 20
rect 8845 0 8865 20
rect 8865 0 8870 20
rect 8840 -5 8870 0
rect 9020 20 9050 25
rect 9020 0 9025 20
rect 9025 0 9045 20
rect 9045 0 9050 20
rect 9020 -5 9050 0
rect 9200 20 9230 25
rect 9200 0 9205 20
rect 9205 0 9225 20
rect 9225 0 9230 20
rect 9200 -5 9230 0
rect 9380 20 9410 25
rect 9380 0 9385 20
rect 9385 0 9405 20
rect 9405 0 9410 20
rect 9380 -5 9410 0
rect 9560 20 9590 25
rect 9560 0 9565 20
rect 9565 0 9585 20
rect 9585 0 9590 20
rect 9560 -5 9590 0
rect 9740 20 9770 25
rect 9740 0 9745 20
rect 9745 0 9765 20
rect 9765 0 9770 20
rect 9740 -5 9770 0
rect 9920 20 9950 25
rect 9920 0 9925 20
rect 9925 0 9945 20
rect 9945 0 9950 20
rect 9920 -5 9950 0
rect 10100 20 10130 25
rect 10100 0 10105 20
rect 10105 0 10125 20
rect 10125 0 10130 20
rect 10100 -5 10130 0
rect 10280 20 10310 25
rect 10280 0 10285 20
rect 10285 0 10305 20
rect 10305 0 10310 20
rect 10280 -5 10310 0
rect 10460 20 10490 25
rect 10460 0 10465 20
rect 10465 0 10485 20
rect 10485 0 10490 20
rect 10460 -5 10490 0
rect 10640 20 10670 25
rect 10640 0 10645 20
rect 10645 0 10665 20
rect 10665 0 10670 20
rect 10640 -5 10670 0
rect 11180 20 11210 25
rect 11180 0 11185 20
rect 11185 0 11205 20
rect 11205 0 11210 20
rect 11180 -5 11210 0
rect 11315 20 11345 25
rect 11315 0 11320 20
rect 11320 0 11340 20
rect 11340 0 11345 20
rect 11315 -5 11345 0
<< metal2 >>
rect -485 1845 11350 1850
rect -485 1815 -480 1845
rect -450 1815 -345 1845
rect -315 1815 195 1845
rect 225 1815 375 1845
rect 405 1815 555 1845
rect 585 1815 735 1845
rect 765 1815 915 1845
rect 945 1815 1095 1845
rect 1125 1815 1275 1845
rect 1305 1815 1455 1845
rect 1485 1815 1635 1845
rect 1665 1815 1815 1845
rect 1845 1815 1995 1845
rect 2025 1815 2175 1845
rect 2205 1815 2355 1845
rect 2385 1815 2535 1845
rect 2565 1815 2715 1845
rect 2745 1815 2895 1845
rect 2925 1815 3080 1845
rect 3110 1815 3260 1845
rect 3290 1815 3440 1845
rect 3470 1815 3620 1845
rect 3650 1815 3800 1845
rect 3830 1815 3980 1845
rect 4010 1815 4160 1845
rect 4190 1815 4340 1845
rect 4370 1815 4520 1845
rect 4550 1815 4700 1845
rect 4730 1815 4880 1845
rect 4910 1815 5060 1845
rect 5090 1815 5240 1845
rect 5270 1815 5420 1845
rect 5450 1815 5600 1845
rect 5630 1815 5780 1845
rect 5810 1815 5960 1845
rect 5990 1815 6140 1845
rect 6170 1815 6320 1845
rect 6350 1815 6500 1845
rect 6530 1815 6680 1845
rect 6710 1815 6860 1845
rect 6890 1815 7040 1845
rect 7070 1815 7220 1845
rect 7250 1815 7400 1845
rect 7430 1815 7580 1845
rect 7610 1815 7760 1845
rect 7790 1815 7940 1845
rect 7970 1815 8120 1845
rect 8150 1815 8300 1845
rect 8330 1815 8480 1845
rect 8510 1815 8660 1845
rect 8690 1815 8840 1845
rect 8870 1815 9020 1845
rect 9050 1815 9200 1845
rect 9230 1815 9380 1845
rect 9410 1815 9560 1845
rect 9590 1815 9740 1845
rect 9770 1815 9920 1845
rect 9950 1815 10100 1845
rect 10130 1815 10280 1845
rect 10310 1815 10460 1845
rect 10490 1815 10640 1845
rect 10670 1815 11180 1845
rect 11210 1815 11315 1845
rect 11345 1815 11350 1845
rect -485 1810 11350 1815
rect -350 965 11215 970
rect -350 935 -345 965
rect -315 935 195 965
rect 225 935 375 965
rect 405 935 555 965
rect 585 935 735 965
rect 765 935 915 965
rect 945 935 1095 965
rect 1125 935 1275 965
rect 1305 935 1455 965
rect 1485 935 1635 965
rect 1665 935 1815 965
rect 1845 935 1995 965
rect 2025 935 2175 965
rect 2205 935 2355 965
rect 2385 935 2535 965
rect 2565 935 2715 965
rect 2745 935 2895 965
rect 2925 935 3080 965
rect 3110 935 3260 965
rect 3290 935 3440 965
rect 3470 935 3620 965
rect 3650 935 3800 965
rect 3830 935 3980 965
rect 4010 935 4160 965
rect 4190 935 4340 965
rect 4370 935 4520 965
rect 4550 935 4700 965
rect 4730 935 4880 965
rect 4910 935 5060 965
rect 5090 935 5240 965
rect 5270 935 5420 965
rect 5450 935 5600 965
rect 5630 935 5780 965
rect 5810 935 5960 965
rect 5990 935 6140 965
rect 6170 935 6320 965
rect 6350 935 6500 965
rect 6530 935 6680 965
rect 6710 935 6860 965
rect 6890 935 7040 965
rect 7070 935 7220 965
rect 7250 935 7400 965
rect 7430 935 7580 965
rect 7610 935 7760 965
rect 7790 935 7940 965
rect 7970 935 8120 965
rect 8150 935 8300 965
rect 8330 935 8480 965
rect 8510 935 8660 965
rect 8690 935 8840 965
rect 8870 935 9020 965
rect 9050 935 9200 965
rect 9230 935 9380 965
rect 9410 935 9560 965
rect 9590 935 9740 965
rect 9770 935 9920 965
rect 9950 935 10100 965
rect 10130 935 10280 965
rect 10310 935 10460 965
rect 10490 935 10640 965
rect 10670 935 11180 965
rect 11210 935 11215 965
rect -350 930 11215 935
rect -350 905 11215 910
rect -350 875 -345 905
rect -315 875 195 905
rect 225 875 375 905
rect 405 875 555 905
rect 585 875 735 905
rect 765 875 915 905
rect 945 875 1095 905
rect 1125 875 1275 905
rect 1305 875 1455 905
rect 1485 875 1635 905
rect 1665 875 1815 905
rect 1845 875 1995 905
rect 2025 875 2175 905
rect 2205 875 2355 905
rect 2385 875 2535 905
rect 2565 875 2715 905
rect 2745 875 2895 905
rect 2925 875 3075 905
rect 3105 875 3255 905
rect 3285 875 3435 905
rect 3465 875 3615 905
rect 3645 875 3795 905
rect 3825 875 3975 905
rect 4005 875 4155 905
rect 4185 875 4335 905
rect 4365 875 4515 905
rect 4545 875 4695 905
rect 4725 875 4875 905
rect 4905 875 5055 905
rect 5085 875 5235 905
rect 5265 875 5415 905
rect 5445 875 5595 905
rect 5625 875 5775 905
rect 5805 875 5955 905
rect 5985 875 6135 905
rect 6165 875 6315 905
rect 6345 875 6495 905
rect 6525 875 6675 905
rect 6705 875 6855 905
rect 6885 875 7035 905
rect 7065 875 7215 905
rect 7245 875 7395 905
rect 7425 875 7575 905
rect 7605 875 7755 905
rect 7785 875 7940 905
rect 7970 875 8120 905
rect 8150 875 8300 905
rect 8330 875 8480 905
rect 8510 875 8660 905
rect 8690 875 8840 905
rect 8870 875 9020 905
rect 9050 875 9200 905
rect 9230 875 9380 905
rect 9410 875 9560 905
rect 9590 875 9740 905
rect 9770 875 9920 905
rect 9950 875 10100 905
rect 10130 875 10280 905
rect 10310 875 10460 905
rect 10490 875 10640 905
rect 10670 875 11180 905
rect 11210 875 11215 905
rect -350 870 11215 875
rect -485 25 11350 30
rect -485 -5 -480 25
rect -450 -5 -345 25
rect -315 -5 195 25
rect 225 -5 375 25
rect 405 -5 555 25
rect 585 -5 735 25
rect 765 -5 915 25
rect 945 -5 1095 25
rect 1125 -5 1275 25
rect 1305 -5 1455 25
rect 1485 -5 1635 25
rect 1665 -5 1815 25
rect 1845 -5 1995 25
rect 2025 -5 2175 25
rect 2205 -5 2355 25
rect 2385 -5 2535 25
rect 2565 -5 2715 25
rect 2745 -5 2895 25
rect 2925 -5 3075 25
rect 3105 -5 3255 25
rect 3285 -5 3435 25
rect 3465 -5 3615 25
rect 3645 -5 3795 25
rect 3825 -5 3975 25
rect 4005 -5 4155 25
rect 4185 -5 4335 25
rect 4365 -5 4515 25
rect 4545 -5 4695 25
rect 4725 -5 4875 25
rect 4905 -5 5055 25
rect 5085 -5 5235 25
rect 5265 -5 5415 25
rect 5445 -5 5595 25
rect 5625 -5 5775 25
rect 5805 -5 5955 25
rect 5985 -5 6135 25
rect 6165 -5 6315 25
rect 6345 -5 6495 25
rect 6525 -5 6675 25
rect 6705 -5 6855 25
rect 6885 -5 7035 25
rect 7065 -5 7215 25
rect 7245 -5 7395 25
rect 7425 -5 7575 25
rect 7605 -5 7755 25
rect 7785 -5 7940 25
rect 7970 -5 8120 25
rect 8150 -5 8300 25
rect 8330 -5 8480 25
rect 8510 -5 8660 25
rect 8690 -5 8840 25
rect 8870 -5 9020 25
rect 9050 -5 9200 25
rect 9230 -5 9380 25
rect 9410 -5 9560 25
rect 9590 -5 9740 25
rect 9770 -5 9920 25
rect 9950 -5 10100 25
rect 10130 -5 10280 25
rect 10310 -5 10460 25
rect 10490 -5 10640 25
rect 10670 -5 11180 25
rect 11210 -5 11315 25
rect 11345 -5 11350 25
rect -485 -10 11350 -5
<< labels >>
rlabel locali 200 270 200 270 1 LO
rlabel locali 200 430 200 430 1 N
rlabel metal2 195 10 195 10 1 VSSA
port 2 n
rlabel metal2 195 890 195 890 1 VDDA
port 1 n
rlabel locali 195 550 195 550 1 P1
rlabel locali 195 470 195 470 1 DP
port 3 n
rlabel locali 195 510 195 510 1 P2
rlabel locali 195 390 195 390 1 X
rlabel locali 195 350 195 350 1 Y
rlabel locali 195 310 195 310 1 Z
rlabel locali 200 630 200 630 1 P0
<< end >>
