* NGSPICE file created from res.ext - technology: sky130A

.subckt res A B C gnd
X0 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X1 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X2 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X3 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X4 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X5 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X6 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X7 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X8 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X9 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X10 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X11 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X12 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X13 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X14 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X15 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X16 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X17 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X18 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X19 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X20 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X21 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X22 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X23 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X24 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X25 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X26 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X27 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X28 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X29 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X30 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X31 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X32 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X33 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X34 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X35 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X36 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X37 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X38 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X39 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X40 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X41 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X42 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X43 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X44 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X45 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X46 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X47 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X48 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X49 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X50 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X51 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X52 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X53 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X54 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X55 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X56 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X57 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X58 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X59 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X60 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X61 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X62 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X63 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X64 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X65 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X66 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X67 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X68 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X69 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X70 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X71 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X72 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X73 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X74 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X75 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X76 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X77 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X78 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X79 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X80 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X81 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X82 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X83 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X84 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X85 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X86 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X87 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X88 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X89 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X90 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X91 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X92 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X93 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X94 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X95 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X96 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X97 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X98 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X99 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X100 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X101 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X102 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X103 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X104 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X105 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X106 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X107 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X108 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X109 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X110 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X111 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X112 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X113 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X114 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X115 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X116 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X117 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X118 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X119 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X120 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X121 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X122 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X123 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X124 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X125 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X126 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X127 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X128 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X129 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X130 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X131 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X132 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X133 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X134 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X135 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X136 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X137 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X138 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X139 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X140 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X141 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X142 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X143 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X144 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X145 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X146 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X147 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X148 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X149 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X150 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X151 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X152 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X153 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X154 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X155 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X156 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X157 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X158 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X159 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X160 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X161 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X162 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X163 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X164 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X165 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X166 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X167 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X168 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X169 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X170 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X171 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X172 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X173 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X174 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X175 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X176 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X177 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X178 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X179 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X180 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X181 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X182 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X183 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X184 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X185 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X186 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X187 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X188 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X189 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X190 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X191 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X192 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X193 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X194 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X195 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X196 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X197 C B gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X198 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
X199 B A gnd sky130_fd_pr__res_xhigh_po w=350000u l=3.5e+07u
.ends

