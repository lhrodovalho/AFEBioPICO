magic
tech sky130A
timestamp 1634675472
<< metal3 >>
rect -220 -170 820 920
rect -220 -260 -200 -170
rect 800 -260 820 -170
rect -220 -1350 820 -260
<< via3 >>
rect -200 -260 800 -170
<< mimcap >>
rect -200 800 800 900
rect -200 0 -100 800
rect 700 0 800 800
rect -200 -100 800 0
rect -200 -430 800 -330
rect -200 -1230 -100 -430
rect 700 -1230 800 -430
rect -200 -1330 800 -1230
<< mimcapcontact >>
rect -100 0 700 800
rect -100 -1230 700 -430
<< metal4 >>
rect -250 1140 850 1250
rect -250 920 850 1030
rect -220 800 820 920
rect -220 0 -100 800
rect 700 0 820 800
rect -220 -120 820 0
rect -250 -170 820 -160
rect -250 -260 -200 -170
rect 800 -260 820 -170
rect -250 -270 820 -260
rect -220 -430 820 -310
rect -220 -1230 -100 -430
rect 700 -1230 820 -430
rect -220 -1350 820 -1230
rect -250 -1460 850 -1350
rect -250 -1680 850 -1570
<< end >>
