magic
tech sky130A
timestamp 1633742592
<< dnwell >>
rect -180 -130 2150 2020
<< nwell >>
rect -290 1980 2260 2130
rect -290 1260 -140 1980
rect 940 1260 1030 1980
rect 2110 1260 2260 1980
rect -290 630 2260 1260
rect -290 -90 -140 630
rect 940 -90 1030 630
rect 2110 -90 2260 630
rect -290 -240 2260 -90
<< mvnmos >>
rect 0 1790 800 1890
rect 0 1660 800 1760
rect 0 1530 800 1630
rect 0 1400 800 1500
rect 0 390 800 490
rect 0 260 800 360
rect 0 130 800 230
rect 0 0 800 100
rect 1170 1790 1970 1890
rect 1170 1660 1970 1760
rect 1170 1530 1970 1630
rect 1170 1400 1970 1500
rect 1170 390 1970 490
rect 1170 260 1970 360
rect 1170 130 1970 230
rect 1170 0 1970 100
<< mvndiff >>
rect -50 1870 0 1890
rect -50 1810 -40 1870
rect -10 1810 0 1870
rect -50 1790 0 1810
rect 800 1870 850 1890
rect 800 1810 810 1870
rect 840 1810 850 1870
rect 800 1790 850 1810
rect -50 1740 0 1760
rect -50 1680 -40 1740
rect -10 1680 0 1740
rect -50 1660 0 1680
rect 800 1740 850 1760
rect 800 1680 810 1740
rect 840 1680 850 1740
rect 800 1660 850 1680
rect -50 1610 0 1630
rect -50 1550 -40 1610
rect -10 1550 0 1610
rect -50 1530 0 1550
rect 800 1610 850 1630
rect 800 1550 810 1610
rect 840 1550 850 1610
rect 800 1530 850 1550
rect -50 1480 0 1500
rect -50 1420 -40 1480
rect -10 1420 0 1480
rect -50 1400 0 1420
rect 800 1480 850 1500
rect 800 1420 810 1480
rect 840 1420 850 1480
rect 800 1400 850 1420
rect -50 470 0 490
rect -50 410 -40 470
rect -10 410 0 470
rect -50 390 0 410
rect 800 470 850 490
rect 800 410 810 470
rect 840 410 850 470
rect 800 390 850 410
rect -50 340 0 360
rect -50 280 -40 340
rect -10 280 0 340
rect -50 260 0 280
rect 800 340 850 360
rect 800 280 810 340
rect 840 280 850 340
rect 800 260 850 280
rect -50 210 0 230
rect -50 150 -40 210
rect -10 150 0 210
rect -50 130 0 150
rect 800 210 850 230
rect 800 150 810 210
rect 840 150 850 210
rect 800 130 850 150
rect -50 80 0 100
rect -50 20 -40 80
rect -10 20 0 80
rect -50 0 0 20
rect 800 80 850 100
rect 800 20 810 80
rect 840 20 850 80
rect 800 0 850 20
rect 1120 1870 1170 1890
rect 1120 1810 1130 1870
rect 1160 1810 1170 1870
rect 1120 1790 1170 1810
rect 1970 1870 2020 1890
rect 1970 1810 1980 1870
rect 2010 1810 2020 1870
rect 1970 1790 2020 1810
rect 1120 1740 1170 1760
rect 1120 1680 1130 1740
rect 1160 1680 1170 1740
rect 1120 1660 1170 1680
rect 1970 1740 2020 1760
rect 1970 1680 1980 1740
rect 2010 1680 2020 1740
rect 1970 1660 2020 1680
rect 1120 1610 1170 1630
rect 1120 1550 1130 1610
rect 1160 1550 1170 1610
rect 1120 1530 1170 1550
rect 1970 1610 2020 1630
rect 1970 1550 1980 1610
rect 2010 1550 2020 1610
rect 1970 1530 2020 1550
rect 1120 1480 1170 1500
rect 1120 1420 1130 1480
rect 1160 1420 1170 1480
rect 1120 1400 1170 1420
rect 1970 1480 2020 1500
rect 1970 1420 1980 1480
rect 2010 1420 2020 1480
rect 1970 1400 2020 1420
rect 1120 470 1170 490
rect 1120 410 1130 470
rect 1160 410 1170 470
rect 1120 390 1170 410
rect 1970 470 2020 490
rect 1970 410 1980 470
rect 2010 410 2020 470
rect 1970 390 2020 410
rect 1120 340 1170 360
rect 1120 280 1130 340
rect 1160 280 1170 340
rect 1120 260 1170 280
rect 1970 340 2020 360
rect 1970 280 1980 340
rect 2010 280 2020 340
rect 1970 260 2020 280
rect 1120 210 1170 230
rect 1120 150 1130 210
rect 1160 150 1170 210
rect 1120 130 1170 150
rect 1970 210 2020 230
rect 1970 150 1980 210
rect 2010 150 2020 210
rect 1970 130 2020 150
rect 1120 80 1170 100
rect 1120 20 1130 80
rect 1160 20 1170 80
rect 1120 0 1170 20
rect 1970 80 2020 100
rect 1970 20 1980 80
rect 2010 20 2020 80
rect 1970 0 2020 20
<< mvndiffc >>
rect -40 1810 -10 1870
rect 810 1810 840 1870
rect -40 1680 -10 1740
rect 810 1680 840 1740
rect -40 1550 -10 1610
rect 810 1550 840 1610
rect -40 1420 -10 1480
rect 810 1420 840 1480
rect -40 410 -10 470
rect 810 410 840 470
rect -40 280 -10 340
rect 810 280 840 340
rect -40 150 -10 210
rect 810 150 840 210
rect -40 20 -10 80
rect 810 20 840 80
rect 1130 1810 1160 1870
rect 1980 1810 2010 1870
rect 1130 1680 1160 1740
rect 1980 1680 2010 1740
rect 1130 1550 1160 1610
rect 1980 1550 2010 1610
rect 1130 1420 1160 1480
rect 1980 1420 2010 1480
rect 1130 410 1160 470
rect 1980 410 2010 470
rect 1130 280 1160 340
rect 1980 280 2010 340
rect 1130 150 1160 210
rect 1980 150 2010 210
rect 1130 20 1160 80
rect 1980 20 2010 80
<< psubdiff >>
rect -360 2170 -310 2200
rect 2280 2170 2330 2200
rect -360 2150 -330 2170
rect 2300 2150 2330 2170
rect -360 -280 -330 -260
rect 2300 -280 2330 -260
rect -360 -310 -310 -280
rect 2280 -310 2330 -280
<< nsubdiff >>
rect -210 2020 -140 2050
rect 940 2020 1030 2050
rect 2110 2020 2180 2050
rect -210 1980 -180 2020
rect -180 930 -160 960
rect 950 930 970 960
rect -210 -130 -180 -90
rect 2150 1980 2180 2020
rect 1000 930 1020 960
rect 2130 930 2150 960
rect 2150 -130 2180 -90
rect -210 -160 -140 -130
rect 940 -160 1030 -130
rect 2110 -160 2180 -130
<< mvpsubdiff >>
rect -120 1930 -70 1960
rect 870 1930 920 1960
rect -120 1910 -90 1930
rect 890 1910 920 1930
rect -120 1310 -90 1330
rect 890 1310 920 1330
rect -120 1280 -70 1310
rect 870 1280 920 1310
rect -120 580 -70 610
rect 870 580 920 610
rect -120 560 -90 580
rect 890 560 920 580
rect -120 -40 -90 -20
rect 890 -40 920 -20
rect -120 -70 -70 -40
rect 870 -70 920 -40
rect 1050 1930 1100 1960
rect 2040 1930 2090 1960
rect 1050 1910 1080 1930
rect 2060 1910 2090 1930
rect 1050 1310 1080 1330
rect 2060 1310 2090 1330
rect 1050 1280 1100 1310
rect 2040 1280 2090 1310
rect 1050 580 1100 610
rect 2040 580 2090 610
rect 1050 560 1080 580
rect 2060 560 2090 580
rect 1050 -40 1080 -20
rect 2060 -40 2090 -20
rect 1050 -70 1100 -40
rect 2040 -70 2090 -40
<< psubdiffcont >>
rect -310 2170 2280 2200
rect -360 -260 -330 2150
rect 2300 -260 2330 2150
rect -310 -310 2280 -280
<< nsubdiffcont >>
rect -140 2020 940 2050
rect 1030 2020 2110 2050
rect -210 -90 -180 1980
rect -160 930 950 960
rect 970 -130 1000 2020
rect 1020 930 2130 960
rect 2150 -90 2180 1980
rect -140 -160 940 -130
rect 1030 -160 2110 -130
<< mvpsubdiffcont >>
rect -70 1930 870 1960
rect -120 1330 -90 1910
rect 890 1330 920 1910
rect -70 1280 870 1310
rect -70 580 870 610
rect -120 -20 -90 560
rect 890 -20 920 560
rect -70 -70 870 -40
rect 1100 1930 2040 1960
rect 1050 1330 1080 1910
rect 2060 1330 2090 1910
rect 1100 1280 2040 1310
rect 1100 580 2040 610
rect 1050 -20 1080 560
rect 2060 -20 2090 560
rect 1100 -70 2040 -40
<< poly >>
rect 0 1890 800 1910
rect 0 1760 800 1790
rect 0 1630 800 1660
rect 0 1500 800 1530
rect 0 1370 800 1400
rect 0 1340 20 1370
rect 780 1340 800 1370
rect 0 1330 800 1340
rect 0 550 800 560
rect 0 520 20 550
rect 780 520 800 550
rect 0 490 800 520
rect 0 360 800 390
rect 0 230 800 260
rect 0 100 800 130
rect 0 -20 800 0
rect 1170 1890 1970 1910
rect 1170 1760 1970 1790
rect 1170 1630 1970 1660
rect 1170 1500 1970 1530
rect 1170 1370 1970 1400
rect 1170 1340 1190 1370
rect 1950 1340 1970 1370
rect 1170 1330 1970 1340
rect 1170 550 1970 560
rect 1170 520 1190 550
rect 1950 520 1970 550
rect 1170 490 1970 520
rect 1170 360 1970 390
rect 1170 230 1970 260
rect 1170 100 1970 130
rect 1170 -20 1970 0
<< polycont >>
rect 20 1340 780 1370
rect 20 520 780 550
rect 1190 1340 1950 1370
rect 1190 520 1950 550
<< locali >>
rect -360 2170 -310 2200
rect 2280 2170 2330 2200
rect -360 2150 -330 2170
rect 2300 2150 2330 2170
rect -180 2020 -140 2050
rect 940 2020 1030 2050
rect 2110 2020 2180 2050
rect -210 1980 -180 2020
rect -120 1930 -70 1960
rect 870 1930 920 1960
rect -120 1910 -90 1930
rect -40 1870 -10 1930
rect 890 1910 920 1930
rect -40 1790 -10 1810
rect 810 1870 840 1890
rect -40 1740 -10 1760
rect -40 1610 -10 1680
rect 810 1740 840 1810
rect 810 1660 840 1680
rect -40 1530 -10 1550
rect 810 1610 840 1630
rect -40 1480 -10 1500
rect -40 1400 -10 1420
rect 810 1480 840 1550
rect 810 1400 840 1420
rect 10 1340 20 1370
rect 780 1340 790 1370
rect -120 1310 -90 1330
rect 890 1310 920 1330
rect -120 1280 -70 1310
rect 870 1280 920 1310
rect -180 930 -160 960
rect 950 930 970 960
rect -120 580 -70 610
rect 870 580 920 610
rect -120 560 -90 580
rect 890 560 920 580
rect 10 520 20 550
rect 780 520 790 550
rect -40 470 -10 490
rect -40 390 -10 410
rect 810 470 840 490
rect -40 340 -10 360
rect -40 210 -10 280
rect 810 340 840 410
rect 810 260 840 280
rect -40 130 -10 150
rect 810 210 840 230
rect -120 -40 -90 -20
rect -40 80 -10 100
rect -40 -40 -10 20
rect 810 80 840 150
rect 810 0 840 20
rect 890 -40 920 -20
rect -120 -70 -70 -40
rect 870 -70 920 -40
rect -210 -130 -180 -90
rect 2150 1980 2180 2020
rect 1050 1930 1100 1960
rect 2040 1930 2090 1960
rect 1050 1910 1080 1930
rect 1130 1870 1160 1890
rect 1130 1740 1160 1810
rect 1980 1870 2010 1930
rect 1980 1790 2010 1810
rect 2060 1910 2090 1930
rect 1130 1660 1160 1680
rect 1980 1740 2010 1760
rect 1130 1610 1160 1630
rect 1130 1480 1160 1550
rect 1980 1610 2010 1680
rect 1980 1530 2010 1550
rect 1130 1400 1160 1420
rect 1980 1480 2010 1500
rect 1980 1400 2010 1420
rect 1180 1340 1190 1370
rect 1950 1340 1960 1370
rect 1050 1310 1080 1330
rect 2060 1310 2090 1330
rect 1050 1280 1100 1310
rect 2040 1280 2090 1310
rect 1000 930 1020 960
rect 2130 930 2150 960
rect 1050 580 1100 610
rect 2040 580 2090 610
rect 1050 560 1080 580
rect 2060 560 2090 580
rect 1180 520 1190 550
rect 1950 520 1960 550
rect 1130 470 1160 490
rect 1130 340 1160 410
rect 1980 470 2010 490
rect 1980 390 2010 410
rect 1130 260 1160 280
rect 1980 340 2010 360
rect 1130 210 1160 230
rect 1130 80 1160 150
rect 1980 210 2010 280
rect 1980 130 2010 150
rect 1130 0 1160 20
rect 1980 80 2010 100
rect 1050 -40 1080 -20
rect 1980 -40 2010 20
rect 2060 -40 2090 -20
rect 1050 -70 1100 -40
rect 2040 -70 2090 -40
rect 2150 -130 2180 -90
rect -180 -160 -140 -130
rect 940 -160 1030 -130
rect 2110 -160 2180 -130
rect -360 -280 -330 -260
rect 2300 -280 2330 -260
rect -360 -310 -310 -280
rect 2280 -310 2330 -280
<< viali >>
rect -210 2020 -180 2050
rect -40 1810 -10 1870
rect -40 1420 -10 1480
rect 750 1340 780 1370
rect -210 1230 -180 1260
rect -210 1130 -180 1160
rect -210 1030 -180 1060
rect -210 930 -180 960
rect -210 830 -180 860
rect -210 730 -180 760
rect -210 630 -180 660
rect 750 520 780 550
rect -40 410 -10 470
rect -40 20 -10 80
rect 1980 1810 2010 1870
rect 1980 1420 2010 1480
rect 1190 1340 1220 1370
rect 1190 520 1220 550
rect 1980 410 2010 470
rect 1980 20 2010 80
rect -210 -160 -180 -130
<< metal1 >>
rect -40 2100 -10 2110
rect -220 2050 -170 2060
rect -220 2020 -210 2050
rect -180 2020 -170 2050
rect -220 2010 -170 2020
rect -40 1890 -10 2070
rect 1980 2000 2010 2110
rect 1980 1890 2010 1970
rect -50 1870 0 1890
rect -50 1810 -40 1870
rect -10 1810 0 1870
rect -50 1790 0 1810
rect 1970 1870 2020 1890
rect 1970 1810 1980 1870
rect 2010 1810 2020 1870
rect 1970 1790 2020 1810
rect -50 1480 0 1500
rect -50 1420 -40 1480
rect -10 1420 0 1480
rect -50 1400 0 1420
rect 1970 1480 2020 1500
rect 1970 1420 1980 1480
rect 2010 1420 2020 1480
rect 1970 1400 2020 1420
rect -220 1260 -170 1270
rect -220 1230 -210 1260
rect -180 1230 -170 1260
rect -220 1160 -170 1230
rect -220 1130 -210 1160
rect -180 1130 -170 1160
rect -220 1060 -170 1130
rect -220 1030 -210 1060
rect -180 1030 -170 1060
rect -220 960 -170 1030
rect -40 1010 -10 1400
rect 740 1370 790 1380
rect 740 1340 750 1370
rect 780 1340 790 1370
rect 740 1330 790 1340
rect 1180 1370 1230 1380
rect 1180 1340 1190 1370
rect 1220 1340 1230 1370
rect 1180 1330 1230 1340
rect -40 970 -10 980
rect 20 1260 50 1270
rect -220 930 -210 960
rect -180 930 -170 960
rect -220 860 -170 930
rect -220 830 -210 860
rect -180 830 -170 860
rect -220 760 -170 830
rect -220 730 -210 760
rect -180 730 -170 760
rect -220 660 -170 730
rect -220 630 -210 660
rect -180 630 -170 660
rect -220 620 -170 630
rect -40 810 -10 820
rect -40 490 -10 780
rect 20 660 50 1230
rect 80 1110 110 1120
rect 80 810 110 1080
rect 750 910 780 1330
rect 750 870 780 880
rect 810 1260 840 1270
rect 80 770 110 780
rect 20 620 50 630
rect 750 710 780 720
rect 750 560 780 680
rect 810 660 840 1230
rect 870 1210 900 1220
rect 870 710 900 1180
rect 1190 1210 1220 1330
rect 1190 1170 1220 1180
rect 1980 1110 2010 1400
rect 1980 1070 2010 1080
rect 1980 1010 2010 1020
rect 870 670 900 680
rect 1190 910 1220 920
rect 810 620 840 630
rect 1190 560 1220 880
rect 740 550 790 560
rect 740 520 750 550
rect 780 520 790 550
rect 740 510 790 520
rect 1180 550 1230 560
rect 1180 520 1190 550
rect 1220 520 1230 550
rect 1180 510 1230 520
rect 1980 490 2010 980
rect -50 470 0 490
rect -50 410 -40 470
rect -10 410 0 470
rect -50 390 0 410
rect 1970 470 2020 490
rect 1970 410 1980 470
rect 2010 410 2020 470
rect 1970 390 2020 410
rect -50 80 0 100
rect -50 20 -40 80
rect -10 20 0 80
rect -50 0 0 20
rect 1970 80 2020 100
rect 1970 20 1980 80
rect 2010 20 2020 80
rect 1970 0 2020 20
rect -40 -80 -10 0
rect -220 -130 -170 -120
rect -220 -160 -210 -130
rect -180 -160 -170 -130
rect -220 -170 -170 -160
rect -40 -220 -10 -110
rect 1980 -180 2010 0
rect 1980 -220 2010 -210
<< via1 >>
rect -40 2070 -10 2100
rect -210 2020 -180 2050
rect 1980 1970 2010 2000
rect -40 980 -10 1010
rect 20 1230 50 1260
rect -40 780 -10 810
rect 80 1080 110 1110
rect 750 880 780 910
rect 810 1230 840 1260
rect 80 780 110 810
rect 20 630 50 660
rect 750 680 780 710
rect 870 1180 900 1210
rect 1190 1180 1220 1210
rect 1980 1080 2010 1110
rect 1980 980 2010 1010
rect 870 680 900 710
rect 1190 880 1220 910
rect 810 630 840 660
rect -40 -110 -10 -80
rect -210 -160 -180 -130
rect 1980 -210 2010 -180
<< metal2 >>
rect -370 2070 -40 2100
rect -10 2070 2340 2100
rect -370 2020 -210 2050
rect -180 2020 2340 2050
rect -370 1970 1980 2000
rect 2010 1970 2340 2000
rect -370 1230 20 1260
rect 50 1230 810 1260
rect 840 1230 2340 1260
rect -370 1180 870 1210
rect 900 1180 1190 1210
rect 1220 1180 2340 1210
rect -370 1130 2340 1160
rect -370 1080 80 1110
rect 110 1080 1980 1110
rect 2010 1080 2340 1110
rect -370 1030 2340 1060
rect -370 980 -40 1010
rect -10 980 1980 1010
rect 2010 980 2340 1010
rect -370 930 2340 960
rect -370 880 750 910
rect 780 880 1190 910
rect 1220 880 2340 910
rect -370 830 2340 860
rect -370 780 -40 810
rect -10 780 80 810
rect 110 780 2340 810
rect -370 730 2340 760
rect -370 680 750 710
rect 780 680 870 710
rect 900 680 2340 710
rect -370 630 20 660
rect 50 630 810 660
rect 840 630 2340 660
rect -370 -110 -40 -80
rect -10 -110 2340 -80
rect -370 -160 -210 -130
rect -180 -160 2340 -130
rect -370 -210 1980 -180
rect 2010 -210 2340 -180
<< labels >>
rlabel metal2 -370 1180 -360 1210 3 ga
port 1 e
rlabel metal2 -370 1080 -360 1110 3 da
port 2 e
rlabel metal2 -370 -110 -360 -80 3 pa
port 3 e
rlabel metal2 2330 1970 2340 2000 7 ma
port 4 w
rlabel metal2 -370 880 -360 910 3 gb
port 5 e
rlabel metal2 -370 980 -360 1010 3 db
port 6 e
rlabel metal2 -370 2070 -360 2100 3 pb
port 7 e
rlabel metal2 2330 -210 2340 -180 7 mb
port 8 w
rlabel metal2 -370 630 -360 660 3 cm
port 9 e
rlabel locali -360 -310 -330 -280 1 gnd
port 10 n
rlabel locali 820 110 830 120 1 a1
rlabel locali -30 240 -20 250 1 a2
rlabel locali 820 370 830 380 1 a3
rlabel locali 1140 1510 1150 1520 1 a4
rlabel locali 1990 1640 2000 1650 1 a5
rlabel locali 1140 1770 1150 1780 1 a6
rlabel locali 820 1770 830 1780 1 b1
rlabel locali -30 1640 -20 1650 1 b2
rlabel locali 820 1510 830 1520 1 b3
rlabel locali 1140 370 1150 380 1 b4
rlabel locali 1990 240 2000 250 1 b5
rlabel locali 1140 110 1150 120 1 b6
<< end >>
