* NGSPICE file created from iref.ext - technology: sky130A

.subckt iref VDDA VSSA DP
X0 a_6585_1690# N a_6495_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X1 a_4425_1690# N a_4335_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X2 a_10995_50# a_10675_35# a_10675_35# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X3 a_10005_750# P2 DP VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X4 a_4060_750# N N VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=1.6e+12p ps=1.12e+07u w=1e+06u l=500000u
X5 a_n170_990# a_n310_975# a_n260_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X6 a_8475_1690# Y a_8385_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X7 a_3520_750# P1 a_3430_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X8 a_6315_1690# N a_6225_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X9 a_9195_990# P1 a_9105_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X10 a_5770_750# P2 a_5680_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X11 a_1360_750# P2 a_1270_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X12 VSSA X a_10365_1690# VSSA sky130_fd_pr__nfet_01v8 ad=1.05e+13p pd=7.3e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X13 N LO P1 VSSA sky130_fd_pr__nfet_01v8 ad=1.6e+12p pd=1.12e+07u as=1.6e+12p ps=1.12e+07u w=1e+06u l=500000u
X14 a_1990_50# X a_1900_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X15 a_4245_990# P0 a_4155_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X16 a_8205_1690# Y a_8115_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X17 a_8475_50# N a_8385_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X18 a_6495_990# P2 a_6405_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X19 a_5680_50# Y P0 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X20 VDDA LO a_280_750# VDDA sky130_fd_pr__pfet_01v8 ad=9.7e+12p pd=6.74e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X21 a_10005_1690# X a_9915_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X22 a_10185_1690# X Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=3.2e+12p ps=2.24e+07u w=1e+06u l=500000u
X23 a_10275_750# P2 a_10185_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X24 a_10005_50# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X25 a_7845_1690# X a_7755_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X26 P1 P2 a_3705_990# VDDA sky130_fd_pr__pfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X27 a_2260_990# P2 a_2170_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X28 a_4420_50# N a_4330_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X29 P2 P2 a_8385_750# VDDA sky130_fd_pr__pfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X30 VSSA N LO VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X31 a_1720_990# P2 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X32 X X a_9645_1690# VSSA sky130_fd_pr__nfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X33 a_8745_50# N a_8655_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X34 a_370_1690# Z a_280_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X35 a_2350_1690# N a_2260_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X36 a_6400_750# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X37 a_7935_750# P2 a_7845_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X38 VDDA a_10675_975# a_11085_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X39 a_730_990# P2 a_640_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X40 P2 N a_1900_1690# VSSA sky130_fd_pr__nfet_01v8 ad=1.6e+12p pd=1.12e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X41 a_2080_1690# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X42 VDDA LO a_10545_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X43 a_7125_990# P2 a_7035_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X44 a_3700_750# P2 a_3610_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X45 a_2260_50# Y Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X46 X P2 a_9285_990# VDDA sky130_fd_pr__pfet_01v8 ad=1.6e+12p pd=1.12e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X47 a_640_50# X a_550_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X48 a_5950_750# P2 a_5860_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X49 a_n310_700# a_n310_700# a_n170_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X50 a_8835_990# P1 a_8745_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X51 a_1720_1690# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X52 a_3790_50# N a_3700_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X53 a_4425_990# P0 a_4335_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X54 a_9105_750# P2 a_9015_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X55 N P2 a_6585_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X56 a_10_1690# a_n310_1640# a_n310_1640# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X57 a_7480_50# N a_7390_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X58 a_550_750# P1 a_460_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X59 a_10455_750# P1 a_10365_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X60 Y Y a_2440_50# VSSA sky130_fd_pr__nfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X61 a_3975_1690# N a_3885_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X62 a_10_990# a_n310_975# a_n310_975# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X63 a_4065_1690# N a_3975_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X64 a_3975_990# P2 a_3885_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X65 a_6220_50# Y a_6130_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X66 a_8655_750# P2 a_8565_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X67 a_4330_750# P2 a_4240_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X68 a_1900_990# P2 a_1810_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X69 a_5865_1690# Y a_5775_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X70 a_10675_35# a_10675_35# a_10815_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X71 a_6580_750# P0 a_6490_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X72 a_3705_1690# N a_3615_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X73 a_2170_750# P1 a_2080_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X74 a_6040_750# P0 a_5950_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X75 DP P2 a_820_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X76 a_1630_750# P2 a_1540_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X77 a_7755_1690# X a_7665_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X78 a_5595_1690# Y a_5505_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X79 a_6850_50# N a_6760_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X80 a_10815_990# a_10675_975# a_10725_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X81 a_7305_990# P1 a_7215_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X82 a_3880_750# P2 a_3790_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X83 a_3435_1690# N a_3345_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X84 P1 LO N VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X85 a_9555_990# P2 a_9465_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X86 a_1900_50# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X87 a_100_50# a_n310_35# a_10_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X88 a_11085_750# a_10675_700# a_10995_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X89 a_640_750# P2 a_550_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X90 a_7485_1690# N a_7395_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X91 a_8385_50# N a_8295_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X92 a_n260_750# a_n310_700# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X93 VDDA P1 a_8925_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X94 P0 Y a_5500_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X95 a_10545_750# P1 a_10455_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X96 VDDA P2 a_2980_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X97 a_5325_1690# Y P0 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X98 a_10_50# a_n310_35# a_n310_35# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X99 a_4605_990# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X100 a_9285_750# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X101 N N a_6765_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X102 VSSA Z a_9825_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X103 a_2530_990# P2 a_2440_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X104 Z X a_9285_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X105 a_7210_750# P2 a_7120_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X106 a_8745_750# P2 a_8655_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X107 a_7215_1690# N a_7125_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X108 a_4330_50# N a_4240_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X109 LO N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X110 a_5050_750# P0 a_4960_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X111 VSSA a_10675_35# a_11085_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X112 VSSA X a_8925_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X113 a_9105_1690# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X114 a_4510_750# P2 a_4420_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X115 a_6760_750# P2 a_6670_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X116 a_10995_1690# a_10675_1640# a_10675_1640# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X117 a_2350_750# P2 a_2260_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X118 a_n170_1690# a_n310_1640# a_n260_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X119 a_11085_1690# a_10675_1640# a_10995_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X120 a_4960_50# Y VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X121 a_9645_990# P1 a_9555_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X122 a_1360_1690# Z a_1270_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X123 a_8745_1690# X Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X124 P0 P2 a_5145_990# VDDA sky130_fd_pr__pfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X125 Z X a_2080_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X126 VDDA P1 a_1720_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X127 a_10995_990# a_10675_975# a_10675_975# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X128 a_7485_990# P1 a_7395_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X129 a_10725_1690# a_10675_1640# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X130 a_3700_50# N a_3610_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X131 a_820_750# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X132 a_6945_990# P2 N VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X133 a_n260_50# a_n310_35# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X134 a_1090_1690# Z a_1000_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X135 a_8025_50# N a_7935_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X136 a_7390_50# N a_7300_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X137 a_10725_750# a_10675_700# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X138 a_4785_990# P0 a_4695_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X139 a_9465_750# P1 a_9375_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X140 a_5140_750# P0 a_5050_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X141 a_2890_1690# N a_2800_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X142 a_2440_50# Y a_2350_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X143 a_2710_990# P2 a_2620_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X144 VSSA Z a_820_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X145 a_7390_750# P2 a_7300_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X146 a_8925_750# P2 a_8835_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X147 a_6130_50# Y a_6040_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X148 a_10815_50# a_10675_35# a_10725_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X149 a_2440_750# P2 a_2350_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X150 a_640_1690# Z a_550_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X151 a_2620_1690# N a_2530_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X152 a_8115_990# P2 a_8025_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X153 a_4690_750# P1 a_4600_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X154 a_9555_50# Z a_9465_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X155 a_6760_50# N a_6670_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X156 a_9825_990# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X157 a_100_1690# a_n310_1640# a_10_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X158 a_4875_1690# Y a_4785_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X159 a_5415_990# P2 a_5325_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X160 a_1990_750# P1 a_1900_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X161 VSSA X a_1720_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X162 a_7665_990# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X163 a_3255_990# P0 a_3165_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X164 a_8295_50# N a_8205_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X165 P1 LO N VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X166 a_5500_50# Y a_5410_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X167 a_1000_750# P1 a_910_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X168 a_1180_990# P2 a_1090_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X169 a_4605_1690# Y VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X170 a_9825_50# Z a_9735_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X171 a_10675_700# a_10675_700# a_10815_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X172 a_4965_990# P2 a_4875_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X173 P1 N a_6940_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X174 a_100_750# a_n310_700# a_10_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X175 a_5320_750# P2 a_5230_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X176 VDDA a_n310_975# a_100_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X177 Z Y a_8565_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X178 a_4240_50# N N VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X179 a_2890_990# P2 a_2800_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X180 a_6495_1690# N a_6405_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X181 VSSA a_n310_35# a_100_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X182 a_7570_750# P0 a_7480_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X183 a_4335_1690# N a_4245_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X184 a_11085_50# a_10675_35# a_10995_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X185 X P2 a_10005_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X186 a_3160_750# P1 a_3070_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X187 P1 P2 a_6940_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X188 a_8385_1690# Y Y VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X189 a_2620_750# P2 Y VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X190 a_6225_1690# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X191 Y P2 a_8205_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X192 VDDA P1 a_4780_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X193 VSSA N a_4780_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X194 a_10365_1690# X a_10275_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X195 a_3345_990# P0 a_3255_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X196 a_8025_1690# Y Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X197 a_2080_50# X a_1990_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X198 a_8115_1690# Y a_8025_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X199 a_10005_990# P2 a_9915_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X200 a_5595_990# P2 a_5505_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X201 a_3610_50# N a_3520_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X202 a_n170_50# a_n310_35# a_n260_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X203 a_9915_1690# X a_9825_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X204 Z X a_10005_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X205 a_550_1690# Z a_460_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X206 a_10455_50# Z a_10365_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X207 a_7935_50# N a_7845_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X208 a_9735_750# P2 a_9645_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X209 a_7300_50# N a_7210_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X210 a_1360_990# P1 a_1270_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X211 a_2260_1690# N a_2170_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X212 a_9645_1690# X a_9555_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X213 a_280_1690# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X214 a_5500_750# P2 a_5410_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X215 a_370_990# P1 a_280_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X216 VDDA P1 a_1000_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X217 VDDA P0 a_7660_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X218 Z X a_1360_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X219 a_10275_990# P2 a_10185_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X220 a_10725_50# a_10675_35# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X221 a_1900_1690# N a_1810_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X222 a_6225_990# P1 a_6135_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X223 a_2980_50# X Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X224 a_2800_750# P2 a_2710_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X225 a_8475_990# P2 a_8385_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X226 a_9465_50# Z a_9375_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X227 a_4065_990# P2 a_3975_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X228 a_6670_50# N a_6580_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X229 a_7935_990# P1 a_7845_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X230 VSSA Z a_1540_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X231 a_3525_990# P2 a_3435_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X232 a_1720_50# X a_1630_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X233 a_8205_750# P2 a_8115_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X234 a_5775_990# P0 a_5685_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X235 a_8205_50# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X236 a_5410_50# Y a_5320_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X237 a_6130_750# P0 a_6040_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X238 a_3885_1690# N P1 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X239 a_9735_50# Z a_9645_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X240 DP P2 a_9825_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X241 a_6940_50# N a_6850_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X242 a_n310_975# a_n310_975# a_n170_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X243 a_3430_750# P1 a_3340_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X244 a_5775_1690# Y a_5685_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X245 a_9105_990# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X246 a_5680_750# P2 P0 VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X247 a_550_990# P1 a_460_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X248 a_3615_1690# N a_3525_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X249 a_1270_750# P1 a_1180_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X250 VSSA X a_3160_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X251 VDDA P1 a_10365_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X252 a_7665_1690# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X253 a_5505_1690# Y a_5415_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X254 a_6405_990# P2 a_6315_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X255 a_4780_50# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X256 a_2980_750# P1 a_2890_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X257 a_280_750# LO VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X258 a_3345_1690# N a_3255_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X259 a_8655_990# P2 a_8565_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X260 a_10185_750# P2 a_10095_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X261 a_9555_1690# X a_9465_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X262 a_7395_1690# N a_7305_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X263 a_3705_990# P2 a_3615_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X264 a_2170_990# P2 a_2080_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X265 P0 Y a_5145_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X266 a_3520_50# N a_3430_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X267 a_n310_35# a_n310_35# a_n170_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X268 a_8385_750# P2 a_8295_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X269 VDDA P0 a_5865_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X270 a_10365_50# Z a_10275_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X271 VDDA P1 a_1540_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X272 a_7845_50# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X273 a_9285_1690# X a_9195_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X274 a_7210_50# N a_7120_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X275 VDDA P0 a_6220_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X276 a_7035_1690# N a_6945_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X277 a_7845_750# P2 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X278 a_7125_1690# N a_7035_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X279 a_1000_50# X a_910_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X280 a_11085_990# a_10675_975# a_10995_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X281 N N a_4060_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X282 a_640_990# P2 a_550_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X283 a_n260_990# a_n310_975# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X284 a_8925_1690# X a_8835_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X285 a_10545_990# LO VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X286 a_3610_750# P1 a_3520_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X287 a_1360_50# X a_1270_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X288 a_9285_990# P2 a_9195_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X289 a_5860_750# P2 a_5770_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X290 VSSA Z a_10545_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X291 a_10675_1640# a_10675_1640# a_10815_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X292 X P2 a_1360_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X293 a_n310_1640# a_n310_1640# a_n170_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X294 a_5050_50# Y a_4960_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X295 a_8745_990# P1 a_8655_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X296 Z Y a_2800_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X297 a_4335_990# P0 a_4245_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X298 a_1270_1690# Z a_1180_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X299 a_9375_50# Z a_9285_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X300 a_6585_990# P2 a_6495_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X301 a_6580_50# N a_6490_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X302 a_460_750# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X303 VSSA N LO VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X304 a_6045_990# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X305 a_10365_750# P1 a_10275_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X306 a_1630_50# X a_1540_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X307 P2 N a_8025_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X308 P2 P2 a_2260_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X309 a_3885_990# P2 P1 VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X310 a_5320_50# Y a_5230_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X311 a_8565_750# P2 P2 VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X312 a_4240_750# P2 N VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X313 a_2800_1690# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X314 a_1810_990# P2 a_1720_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X315 a_820_1690# Z a_730_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X316 a_9645_50# Z a_9555_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X317 a_6490_750# P0 a_6400_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X318 a_8025_750# P2 a_7935_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X319 a_2080_750# P1 a_1990_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X320 a_3255_1690# N a_3165_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X321 a_820_990# P2 a_730_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X322 a_1540_750# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X323 a_2530_1690# N a_2440_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X324 a_5950_50# Y a_5860_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X325 a_10725_990# a_10675_975# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X326 a_7215_990# P2 a_7125_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X327 a_3790_750# P2 a_3700_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X328 a_3160_50# X a_3070_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X329 a_9465_990# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X330 a_5055_990# P2 a_4965_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X331 a_n170_750# a_n310_700# a_n260_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X332 a_8925_990# P1 a_8835_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X333 VSSA N a_4600_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X334 VDDA P0 a_4425_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X335 a_4785_1690# Y a_4695_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X336 VDDA P2 a_9105_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X337 a_6765_990# N N VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X338 a_9015_50# N a_8925_50# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X339 a_2440_990# P2 P2 VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X340 a_7120_750# P2 P1 VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X341 N N a_6585_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X342 a_3430_50# N a_3340_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X343 VSSA N a_4425_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X344 a_10275_50# Z a_10185_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X345 a_7120_50# N P1 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X346 a_8565_1690# Y a_8475_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X347 a_4420_750# P2 a_4330_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X348 a_910_50# X a_820_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X349 a_1990_990# P2 a_1900_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X350 a_6405_1690# N a_6315_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X351 a_6670_750# P0 a_6580_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X352 a_4245_1690# N a_4155_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X353 a_2260_750# P2 a_2170_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X354 a_5145_990# P2 a_5055_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X355 a_1000_990# P2 DP VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X356 a_6045_1690# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X357 Y Y a_8205_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X358 a_1270_50# X a_1180_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X359 a_1720_750# P1 a_1630_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X360 VSSA N a_6045_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X361 VSSA N a_7660_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X362 a_10545_50# Z a_10455_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X363 a_10675_975# a_10675_975# a_10815_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X364 a_7395_990# P1 a_7305_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X365 N P2 a_3880_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X366 a_100_990# a_n310_975# a_10_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X367 a_2800_50# Y a_2710_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X368 a_10275_1690# X a_10185_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X369 VDDA a_10675_700# a_11085_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X370 X P2 a_640_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X371 Z X a_7845_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X372 a_9285_50# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X373 VDDA P1 a_10545_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X374 a_6490_50# N a_6400_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X375 a_4695_990# P0 a_4605_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X376 a_9375_750# P1 a_9285_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X377 a_1540_50# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X378 a_2620_990# P2 a_2530_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X379 a_9825_1690# X X VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X380 a_460_1690# Z a_370_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X381 a_7300_750# P2 a_7210_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X382 a_8835_750# P2 a_8745_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X383 a_5230_50# Y a_5140_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X384 a_2170_1690# N a_2080_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X385 VSSA a_n310_1640# a_100_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X386 a_4600_750# P1 a_4510_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X387 a_6850_750# P2 a_6760_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X388 a_10_750# a_n310_700# a_n310_700# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X389 a_8655_50# N a_8565_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X390 a_5860_50# Y a_5770_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X391 VDDA P1 a_9645_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X392 a_1810_1690# N a_1720_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X393 a_5325_990# P2 P0 VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X394 a_1900_750# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X395 a_3070_50# X a_2980_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X396 VDDA P1 a_7485_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X397 a_3165_990# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X398 a_4600_50# N a_4510_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X399 a_7035_990# P2 a_6945_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X400 a_1540_1690# Z a_1450_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X401 a_910_750# P2 a_820_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X402 a_1090_990# P2 a_1000_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X403 a_550_50# X a_460_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X404 a_4155_1690# N a_4065_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X405 a_8925_50# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X406 a_10815_750# a_10675_700# a_10725_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X407 a_4875_990# P0 a_4785_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X408 a_9555_750# P1 a_9465_750# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X409 a_5230_750# P0 a_5140_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X410 a_3340_50# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X411 a_2800_990# P2 a_2710_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X412 VSSA Y a_5865_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X413 a_7480_750# P0 a_7390_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X414 P1 N a_3705_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X415 a_10185_50# Z a_10095_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X416 a_9015_750# P2 a_8925_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X417 a_3070_750# P1 a_2980_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X418 a_6940_750# P2 a_6850_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X419 a_820_50# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X420 Y P2 a_2440_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X421 a_5685_1690# Y a_5595_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X422 a_8205_990# P2 a_8115_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X423 a_4780_750# P1 a_4690_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X424 a_3525_1690# N a_3435_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X425 N N a_3880_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X426 a_1180_50# X X VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X427 VSSA N a_7485_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X428 a_7660_50# N a_7570_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X429 a_9915_990# P1 a_9825_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X430 a_5415_1690# Y a_5325_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X431 a_5505_990# P2 a_5415_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X432 a_2710_50# Y a_2620_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X433 a_7755_990# P1 a_7665_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X434 VSSA N a_9105_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X435 a_9465_1690# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X436 a_9645_750# P2 a_9555_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X437 a_7305_1690# N a_7215_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X438 a_6400_50# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X439 a_1270_990# P2 a_1180_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X440 a_5145_1690# Y a_5055_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X441 a_10995_750# a_10675_700# a_10675_700# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X442 a_6945_1690# N N VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X443 a_9195_1690# X a_9105_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X444 a_5410_750# P2 a_5320_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X445 a_280_990# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X446 a_5140_50# Y a_5050_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X447 a_2980_990# P2 a_2890_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X448 a_7660_750# P0 a_7570_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X449 a_10185_990# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X450 VDDA P1 a_3160_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X451 a_n260_1690# a_n310_1640# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X452 VSSA a_10675_1640# a_11085_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X453 a_1450_1690# Z a_1360_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X454 a_8835_1690# X a_8745_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X455 a_6135_990# P1 a_6045_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X456 a_2710_750# P2 a_2620_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X457 a_8385_990# P2 Y VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X458 a_4960_750# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X459 a_8565_50# N a_8475_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X460 a_10815_1690# a_10675_1640# a_10725_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X461 a_5770_50# Y a_5680_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X462 a_7845_990# P1 a_7755_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X463 a_3435_990# P0 a_3345_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X464 a_1180_1690# Z a_1090_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X465 a_8115_750# P2 a_8025_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X466 a_5685_990# P0 a_5595_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X467 LO N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X468 a_4510_50# N a_4420_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X469 a_2980_1690# N a_2890_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X470 a_1000_1690# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X471 VSSA N a_2980_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X472 a_460_50# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X473 P2 N a_8745_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X474 a_9825_750# P2 a_9735_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X475 a_6040_50# Y a_5950_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X476 a_1450_990# P1 a_1360_990# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X477 a_3340_750# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X478 P2 N a_2620_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X479 a_730_1690# Z a_640_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X480 a_10095_50# Z a_10005_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X481 P0 P2 a_5500_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X482 a_460_990# P1 a_370_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X483 a_1180_750# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X484 a_3165_1690# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X485 a_2350_50# Y a_2260_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X486 a_10365_990# P1 a_10275_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X487 Z X a_640_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X488 a_2440_1690# N a_2350_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X489 a_4965_1690# Y a_4875_1690# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X490 a_6315_990# P1 a_6225_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X491 a_3880_50# N a_3790_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X492 a_2890_750# P2 a_2800_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X493 VDDA a_n310_700# a_100_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X494 a_5055_1690# Y a_4965_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X495 a_8565_990# P2 a_8475_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X496 X X a_1000_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X497 a_10095_750# P2 a_10005_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X498 a_4155_990# P2 a_4065_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X499 a_7570_50# N a_7480_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X500 N LO P1 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X501 a_8025_990# P2 a_7935_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X502 a_3615_990# P2 a_3525_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X503 a_2080_990# P2 a_1990_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X504 a_4695_1690# Y a_4605_1690# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X505 a_2620_50# Y Y VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X506 a_8295_750# P2 a_8205_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X507 a_5865_990# P0 a_5775_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X508 a_9105_50# N a_9015_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X509 a_1540_990# P1 a_1450_990# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X510 VSSA Y a_6220_50# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X511 a_6220_750# P0 a_6130_750# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
.ends

