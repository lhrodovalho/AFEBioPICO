magic
tech sky130A
timestamp 1634082498
<< nwell >>
rect -1220 -6310 15650 2540
rect -1220 -12540 15650 -9710
<< pwell >>
rect -1270 -280 -1240 -230
rect -1270 -370 -1240 -360
rect -1270 -500 -1240 -490
rect -1270 -540 -1240 -530
rect -1270 -3300 -1240 -3250
rect -1270 -3420 -1240 -3370
rect -1270 -3540 -1240 -3490
rect -1270 -7900 -1240 -6250
rect 15670 -280 15700 -230
rect 15670 -370 15700 -360
rect 15670 -500 15700 -490
rect 15670 -540 15700 -530
rect 15670 -3300 15700 -3250
rect 15670 -3420 15700 -3370
rect 15670 -3540 15700 -3490
rect -340 -6740 -310 -6670
rect 590 -6740 620 -6670
rect 730 -6740 760 -6700
rect 2510 -6740 2540 -6700
rect 4450 -6740 4480 -6700
rect 6230 -6740 6260 -6700
rect 8170 -6740 8200 -6700
rect 9950 -6740 9980 -6700
rect 11890 -6740 11920 -6700
rect 13670 -6740 13700 -6700
rect -1140 -6770 1620 -6740
rect 1630 -6770 1640 -6740
rect 1650 -6770 5340 -6740
rect 5350 -6770 5360 -6740
rect 5370 -6770 9060 -6740
rect 9070 -6770 9080 -6740
rect 9090 -6770 12780 -6740
rect 12790 -6770 12800 -6740
rect 12810 -6770 15570 -6740
rect -1270 -7930 -1090 -7900
rect -1130 -7950 -1100 -7930
rect -1130 -8090 -1100 -8070
rect -1270 -8120 -1090 -8090
rect -1270 -9770 -1240 -8120
rect -340 -9250 -310 -6770
rect 590 -7900 620 -6770
rect 15670 -7900 15700 -6250
rect -290 -7930 1620 -7900
rect 1630 -7930 1640 -7900
rect 1650 -7930 5340 -7900
rect 5350 -7930 5360 -7900
rect 5370 -7930 9060 -7900
rect 9070 -7930 9080 -7900
rect 9090 -7930 12780 -7900
rect 12790 -7930 12800 -7900
rect 12810 -7930 14720 -7900
rect 15520 -7930 15700 -7900
rect 590 -8090 620 -7930
rect 15530 -7950 15560 -7930
rect 15530 -8090 15560 -8070
rect -290 -8120 1620 -8090
rect 1630 -8120 1640 -8090
rect 1650 -8120 5340 -8090
rect 5350 -8120 5360 -8090
rect 5370 -8120 9060 -8090
rect 9070 -8120 9080 -8090
rect 9090 -8120 12780 -8090
rect 12790 -8120 12800 -8090
rect 12810 -8120 14720 -8090
rect 15520 -8120 15700 -8090
rect 590 -9240 620 -8120
rect -1140 -9280 1620 -9250
rect 1630 -9280 1640 -9250
rect 1650 -9280 5340 -9250
rect 5350 -9280 5360 -9250
rect 5370 -9280 9060 -9250
rect 9070 -9280 9080 -9250
rect 9090 -9280 12780 -9250
rect 12790 -9280 12800 -9250
rect 12810 -9280 15570 -9250
rect -340 -9350 -310 -9280
rect 590 -9350 620 -9300
rect 730 -9590 760 -9280
rect 1520 -9470 1550 -9290
rect 1720 -9470 1750 -9290
rect 2510 -9590 2540 -9280
rect 4310 -9350 4340 -9300
rect 4450 -9590 4480 -9280
rect 5240 -9470 5270 -9300
rect 5440 -9470 5470 -9300
rect 6230 -9590 6260 -9280
rect 8030 -9350 8060 -9300
rect 8170 -9590 8200 -9280
rect 8960 -9470 8990 -9300
rect 9160 -9470 9190 -9300
rect 9950 -9590 9980 -9280
rect 11750 -9350 11780 -9300
rect 11890 -9590 11920 -9280
rect 12680 -9470 12710 -9300
rect 12880 -9470 12910 -9300
rect 13670 -9590 13700 -9280
rect 15670 -9770 15700 -8120
rect 15670 -12530 15700 -12480
<< psubdiff >>
rect -1270 2570 -1220 2600
rect 15650 2570 15700 2600
rect -1270 2540 -1240 2570
rect 15670 2540 15700 2570
rect -1240 -6770 -1220 -6740
rect 15650 -6770 15670 -6740
rect -1270 -7900 -1240 -7880
rect 15670 -7900 15700 -7880
rect -1270 -7930 15700 -7900
rect -1270 -8120 15700 -8090
rect -1270 -8140 -1240 -8120
rect 15670 -8140 15700 -8120
rect -1240 -9280 -1220 -9250
rect 15650 -9280 15670 -9250
rect -1270 -12560 -1240 -12530
rect 15700 -9280 15710 -9250
rect 15670 -12560 15700 -12530
rect -1270 -12590 -1220 -12560
rect 15650 -12590 15700 -12560
<< nsubdiff >>
rect -1200 2490 15630 2520
rect -1200 2470 -1170 2490
rect 15600 2470 15630 2490
rect -1170 -270 -1150 -240
rect 15580 -270 15600 -240
rect -1170 -530 15600 -500
rect 15600 -3260 15630 -3240
rect -1170 -3290 -1150 -3260
rect 15580 -3290 15630 -3260
rect -1200 -3500 -1170 -3290
rect 15600 -3500 15630 -3290
rect -1170 -3530 15630 -3500
rect -1200 -6260 -1170 -6240
rect 15600 -3550 15630 -3530
rect 15600 -6260 15630 -6240
rect -1200 -6290 -1150 -6260
rect 15580 -6290 15630 -6260
rect -1200 -9760 -1150 -9730
rect 15580 -9760 15630 -9730
rect -1200 -9780 -1170 -9760
rect 15600 -9780 15630 -9760
rect 15600 -12490 15630 -12470
rect -1200 -12520 15630 -12490
<< psubdiffcont >>
rect -1220 2570 15650 2600
rect -1270 -7880 -1240 2540
rect -1220 -6770 15650 -6740
rect 15670 -7880 15700 2540
rect -1270 -12530 -1240 -8140
rect -1220 -9280 15650 -9250
rect 15670 -12530 15700 -8140
rect -1220 -12590 15650 -12560
<< nsubdiffcont >>
rect -1200 -3290 -1170 2470
rect -1150 -270 15580 -240
rect 15600 -3240 15630 2470
rect -1150 -3290 15580 -3260
rect -1200 -6240 -1170 -3500
rect 15600 -6240 15630 -3550
rect -1150 -6290 15580 -6260
rect -1150 -9760 15580 -9730
rect -1200 -12490 -1170 -9780
rect 15600 -12470 15630 -9780
<< locali >>
rect -1270 2570 -1220 2600
rect 15650 2570 15700 2600
rect -1270 2540 -1240 2570
rect -1280 -3300 -1270 -3250
rect 15670 2540 15700 2570
rect -1200 2490 -280 2520
rect -250 2490 14680 2520
rect 14710 2490 15630 2520
rect -1200 2470 -1170 2490
rect 15600 2470 15630 2490
rect -1170 -270 -1150 -240
rect 15580 -270 15600 -240
rect -1280 -3420 -1270 -3370
rect -1240 -3300 -1230 -3250
rect 640 -370 690 -360
rect 640 -470 650 -370
rect 680 -470 690 -370
rect 640 -480 690 -470
rect 2580 -370 2630 -360
rect 2580 -470 2590 -370
rect 2620 -470 2630 -370
rect 2580 -480 2630 -470
rect 4360 -370 4410 -360
rect 4360 -470 4370 -370
rect 4400 -470 4410 -370
rect 4360 -480 4410 -470
rect 6300 -370 6350 -360
rect 6300 -470 6310 -370
rect 6340 -470 6350 -370
rect 6300 -480 6350 -470
rect 8080 -370 8130 -360
rect 8080 -470 8090 -370
rect 8120 -470 8130 -370
rect 8080 -480 8130 -470
rect 10020 -370 10070 -360
rect 10020 -470 10030 -370
rect 10060 -470 10070 -370
rect 10020 -480 10070 -470
rect 11800 -370 11850 -360
rect 11800 -470 11810 -370
rect 11840 -470 11850 -370
rect 11800 -480 11850 -470
rect 13740 -370 13790 -360
rect 13740 -470 13750 -370
rect 13780 -470 13790 -370
rect 13740 -480 13790 -470
rect 650 -500 680 -480
rect 2590 -500 2620 -480
rect 4370 -500 4400 -480
rect 6310 -500 6340 -480
rect 8090 -500 8120 -480
rect 10030 -500 10060 -480
rect 11810 -500 11840 -480
rect 13750 -500 13780 -480
rect -1170 -530 15600 -500
rect 15600 -3260 15630 -3240
rect -1170 -3290 -1150 -3260
rect 15580 -3290 15630 -3260
rect -1280 -3540 -1270 -3490
rect -1240 -3420 -1230 -3370
rect -1240 -3540 -1230 -3490
rect -1200 -3500 -1170 -3290
rect 15660 -3300 15670 -3250
rect -1150 -3470 15670 -3320
rect 15700 -3300 15710 -3250
rect -1170 -3530 15630 -3500
rect -1200 -6260 -1170 -6240
rect 15600 -3550 15630 -3530
rect 15660 -3540 15670 -3490
rect 15700 -3420 15710 -3370
rect 15600 -6260 15630 -6240
rect -1200 -6290 -1150 -6260
rect 15580 -6290 15630 -6260
rect 15700 -3540 15710 -3490
rect -1280 -6710 -1270 -6320
rect -1240 -6710 15670 -6320
rect 15700 -6710 15710 -6320
rect -1240 -6770 -1220 -6740
rect 15650 -6770 15670 -6740
rect -1270 -7900 -1240 -7880
rect 15670 -7900 15700 -7880
rect -1270 -7930 15700 -7900
rect -1130 -7950 -1100 -7930
rect 15530 -7950 15560 -7930
rect -1140 -7960 -1090 -7950
rect -1140 -8060 -1130 -7960
rect -1100 -8060 -1090 -7960
rect -1140 -8070 -1090 -8060
rect 15520 -7960 15570 -7950
rect 15520 -8060 15530 -7960
rect 15560 -8060 15570 -7960
rect 15520 -8070 15570 -8060
rect -1130 -8090 -1100 -8070
rect 15530 -8090 15560 -8070
rect -1270 -8120 15700 -8090
rect -1270 -8140 -1240 -8120
rect -1280 -9290 -1270 -9240
rect 15670 -8140 15700 -8120
rect -1240 -9280 -1220 -9250
rect 15650 -9280 15670 -9250
rect 15700 -9280 15710 -9250
rect -1280 -9410 -1270 -9360
rect -1280 -9530 -1270 -9480
rect -1280 -9650 -1270 -9600
rect -1280 -9770 -1270 -9720
rect -1240 -9700 15670 -9310
rect 15700 -9410 15710 -9360
rect 15700 -9530 15710 -9480
rect 15700 -9650 15710 -9600
rect -1200 -9760 -1150 -9730
rect 15580 -9760 15630 -9730
rect -1200 -9780 -1170 -9760
rect 15600 -9780 15630 -9760
rect -290 -12490 -240 -12480
rect 15600 -12490 15630 -12470
rect -1200 -12520 -280 -12490
rect -250 -12520 15630 -12490
rect -290 -12530 -240 -12520
rect 15660 -12530 15670 -12480
rect 15700 -9770 15710 -9720
rect 15700 -12530 15710 -12480
rect -1270 -12560 -1240 -12530
rect 15670 -12560 15700 -12530
rect -1270 -12590 -1220 -12560
rect 15650 -12590 15700 -12560
<< viali >>
rect -280 2490 -250 2520
rect 14680 2490 14710 2520
rect -1200 -270 -1170 -240
rect 15600 -270 15630 -240
rect -1270 -3290 -1240 -3260
rect 650 -470 680 -370
rect 2590 -470 2620 -370
rect 4370 -470 4400 -370
rect 6310 -470 6340 -370
rect 8090 -470 8120 -370
rect 10030 -470 10060 -370
rect 11810 -470 11840 -370
rect 13750 -470 13780 -370
rect -1270 -3410 -1240 -3380
rect -1270 -3530 -1240 -3500
rect 15670 -3290 15700 -3260
rect 15670 -3410 15700 -3380
rect -1270 -6290 -1240 -6260
rect 15670 -3530 15700 -3500
rect 15670 -6290 15700 -6260
rect -1270 -6410 -1240 -6380
rect -1270 -6530 -1240 -6500
rect -1270 -6650 -1240 -6620
rect 15670 -6410 15700 -6380
rect 15670 -6530 15700 -6500
rect 15670 -6650 15700 -6620
rect -1270 -6770 -1240 -6740
rect 15670 -6770 15700 -6740
rect -1130 -8060 -1100 -7960
rect 15530 -8060 15560 -7960
rect -1270 -9280 -1240 -9250
rect 15670 -9280 15700 -9250
rect -1270 -9400 -1240 -9370
rect -1270 -9520 -1240 -9490
rect -1270 -9640 -1240 -9610
rect 15670 -9400 15700 -9370
rect 15670 -9520 15700 -9490
rect 15670 -9640 15700 -9610
rect -1270 -9760 -1240 -9730
rect 15670 -9760 15700 -9730
rect -280 -12520 -250 -12490
rect 15670 -12520 15700 -12490
<< metal1 >>
rect -280 2530 -250 2540
rect 14680 2530 14710 2540
rect -290 2520 -240 2530
rect 14670 2520 14720 2530
rect -290 2490 -280 2520
rect -250 2490 -240 2520
rect 650 2490 13780 2520
rect 14670 2490 14680 2520
rect 14710 2490 14720 2520
rect -290 2480 -240 2490
rect 14670 2480 14720 2490
rect -1210 -240 -1160 -230
rect -1210 -270 -1200 -240
rect -1170 -270 -1160 -240
rect -1210 -280 -1160 -270
rect -1070 -300 -1040 -170
rect -1280 -3260 -1230 -3250
rect -1280 -3290 -1270 -3260
rect -1240 -3290 -1230 -3260
rect -1280 -3300 -1230 -3290
rect -1280 -3380 -1230 -3370
rect -1280 -3410 -1270 -3380
rect -1240 -3410 -1230 -3380
rect -1280 -3420 -1230 -3410
rect -1280 -3500 -1230 -3490
rect -1280 -3530 -1270 -3500
rect -1240 -3530 -1230 -3500
rect -1280 -3540 -1230 -3530
rect -1280 -6260 -1230 -6250
rect -1280 -6290 -1270 -6260
rect -1240 -6290 -1230 -6260
rect -1280 -6300 -1230 -6290
rect -1070 -6310 -1040 -330
rect -400 -300 -370 -290
rect -400 -3320 -370 -330
rect -400 -3360 -370 -3350
rect -280 -6310 -250 2480
rect -140 -300 -110 -240
rect -140 -340 -110 -330
rect 650 -300 680 -240
rect 650 -340 680 -330
rect 640 -370 690 -360
rect 640 -470 650 -370
rect 680 -470 690 -370
rect 640 -480 690 -470
rect 730 -370 760 -240
rect 1520 -300 1550 -240
rect 1520 -340 1550 -330
rect 1720 -300 1750 -240
rect 1720 -340 1750 -330
rect 730 -480 760 -470
rect 1580 -370 1610 -360
rect 1580 -480 1610 -470
rect 1660 -370 1690 -360
rect 1660 -480 1690 -470
rect 2510 -370 2540 -240
rect 2590 -300 2620 -240
rect 2590 -340 2620 -330
rect 3380 -300 3410 -240
rect 3380 -340 3410 -330
rect 3580 -300 3610 -240
rect 3580 -340 3610 -330
rect 4370 -300 4400 -240
rect 4370 -340 4400 -330
rect 2510 -480 2540 -470
rect 2580 -370 2630 -360
rect 2580 -470 2590 -370
rect 2620 -470 2630 -370
rect 2580 -480 2630 -470
rect 4360 -370 4410 -360
rect 4360 -470 4370 -370
rect 4400 -470 4410 -370
rect 4360 -480 4410 -470
rect 4450 -370 4480 -240
rect 5240 -300 5270 -240
rect 5240 -340 5270 -330
rect 5440 -300 5470 -240
rect 5440 -340 5470 -330
rect 4450 -480 4480 -470
rect 5300 -370 5330 -360
rect 5300 -480 5330 -470
rect 5380 -370 5410 -360
rect 5380 -480 5410 -470
rect 6230 -370 6260 -240
rect 6310 -300 6340 -240
rect 6310 -340 6340 -330
rect 7100 -300 7130 -240
rect 7100 -340 7130 -330
rect 7300 -300 7330 -240
rect 7300 -340 7330 -330
rect 8090 -300 8120 -240
rect 8090 -340 8120 -330
rect 6230 -480 6260 -470
rect 6300 -370 6350 -360
rect 6300 -470 6310 -370
rect 6340 -470 6350 -370
rect 6300 -480 6350 -470
rect 8080 -370 8130 -360
rect 8080 -470 8090 -370
rect 8120 -470 8130 -370
rect 8080 -480 8130 -470
rect 8170 -370 8200 -240
rect 8960 -300 8990 -240
rect 8960 -340 8990 -330
rect 9160 -300 9190 -240
rect 9160 -340 9190 -330
rect 8170 -480 8200 -470
rect 9020 -370 9050 -360
rect 9020 -480 9050 -470
rect 9100 -370 9130 -360
rect 9100 -480 9130 -470
rect 9950 -370 9980 -240
rect 10030 -300 10060 -240
rect 10030 -340 10060 -330
rect 10820 -300 10850 -240
rect 10820 -340 10850 -330
rect 11020 -300 11050 -240
rect 11020 -340 11050 -330
rect 11810 -300 11840 -240
rect 11810 -340 11840 -330
rect 9950 -480 9980 -470
rect 10020 -370 10070 -360
rect 10020 -470 10030 -370
rect 10060 -470 10070 -370
rect 10020 -480 10070 -470
rect 11800 -370 11850 -360
rect 11800 -470 11810 -370
rect 11840 -470 11850 -370
rect 11800 -480 11850 -470
rect 11890 -370 11920 -240
rect 12680 -300 12710 -240
rect 12680 -340 12710 -330
rect 12880 -300 12910 -240
rect 12880 -340 12910 -330
rect 11890 -480 11920 -470
rect 12740 -370 12770 -360
rect 12740 -480 12770 -470
rect 12820 -370 12850 -360
rect 12820 -480 12850 -470
rect 13670 -370 13700 -240
rect 13750 -300 13780 -240
rect 13750 -340 13780 -330
rect 14540 -300 14570 -240
rect 14540 -340 14570 -330
rect 13670 -480 13700 -470
rect 13740 -370 13790 -360
rect 13740 -470 13750 -370
rect 13780 -470 13790 -370
rect 13740 -480 13790 -470
rect 650 -530 680 -480
rect 2590 -530 2620 -480
rect 4370 -530 4400 -480
rect 6310 -530 6340 -480
rect 8090 -530 8120 -480
rect 10030 -530 10060 -480
rect 11810 -530 11840 -480
rect 13750 -530 13780 -480
rect -140 -3320 -110 -3260
rect -140 -3360 -110 -3350
rect 650 -3440 680 -3260
rect 790 -3320 820 -3260
rect 790 -3360 820 -3350
rect 650 -3500 680 -3470
rect 1580 -3440 1610 -3260
rect 1580 -3500 1610 -3470
rect 1660 -3440 1690 -3260
rect 2450 -3320 2480 -3260
rect 2450 -3360 2480 -3350
rect 1660 -3500 1690 -3470
rect 2590 -3440 2620 -3260
rect 3380 -3320 3410 -3260
rect 3380 -3360 3410 -3350
rect 3580 -3320 3610 -3260
rect 3580 -3360 3610 -3350
rect 2590 -3500 2620 -3470
rect 4370 -3440 4400 -3260
rect 4510 -3320 4540 -3260
rect 4510 -3360 4540 -3350
rect 4370 -3500 4400 -3470
rect 5300 -3440 5330 -3260
rect 5300 -3500 5330 -3470
rect 5380 -3440 5410 -3260
rect 6170 -3320 6200 -3260
rect 6170 -3360 6200 -3350
rect 5380 -3500 5410 -3470
rect 6310 -3440 6340 -3260
rect 7100 -3320 7130 -3260
rect 7100 -3360 7130 -3350
rect 7300 -3320 7330 -3260
rect 7300 -3360 7330 -3350
rect 6310 -3500 6340 -3470
rect 8090 -3440 8120 -3260
rect 8230 -3320 8260 -3260
rect 8230 -3360 8260 -3350
rect 8090 -3500 8120 -3470
rect 9020 -3440 9050 -3260
rect 9020 -3500 9050 -3470
rect 9100 -3440 9130 -3260
rect 9890 -3320 9920 -3260
rect 9890 -3360 9920 -3350
rect 9100 -3500 9130 -3470
rect 10030 -3440 10060 -3260
rect 10820 -3320 10850 -3260
rect 10820 -3360 10850 -3350
rect 11020 -3320 11050 -3260
rect 11020 -3360 11050 -3350
rect 10030 -3500 10060 -3470
rect 11810 -3440 11840 -3260
rect 11950 -3320 11980 -3260
rect 11950 -3360 11980 -3350
rect 11810 -3500 11840 -3470
rect 12740 -3440 12770 -3260
rect 12740 -3500 12770 -3470
rect 12820 -3440 12850 -3260
rect 13610 -3320 13640 -3260
rect 13610 -3360 13640 -3350
rect 12820 -3500 12850 -3470
rect 13750 -3440 13780 -3260
rect 14540 -3320 14570 -3260
rect 14540 -3360 14570 -3350
rect 13750 -3500 13780 -3470
rect -140 -6320 -110 -6260
rect -140 -6360 -110 -6350
rect -1280 -6380 -1230 -6370
rect -1280 -6410 -1270 -6380
rect -1240 -6410 -1230 -6380
rect -1280 -6420 -1230 -6410
rect -1280 -6500 -1230 -6490
rect -1280 -6530 -1270 -6500
rect -1240 -6530 -1230 -6500
rect -1280 -6540 -1230 -6530
rect -200 -6560 -170 -6550
rect -1280 -6620 -1230 -6610
rect -1280 -6650 -1270 -6620
rect -1240 -6650 -1230 -6620
rect -1280 -6660 -1230 -6650
rect -340 -6680 -310 -6670
rect -1280 -6740 -1230 -6730
rect -1280 -6770 -1270 -6740
rect -1240 -6770 -1230 -6740
rect -1280 -6780 -1230 -6770
rect -1130 -7950 -1100 -6730
rect -1140 -7960 -1090 -7950
rect -1140 -8060 -1130 -7960
rect -1100 -8060 -1090 -7960
rect -1140 -8070 -1090 -8060
rect -1280 -9250 -1230 -9240
rect -1280 -9280 -1270 -9250
rect -1240 -9280 -1230 -9250
rect -1280 -9290 -1230 -9280
rect -1130 -9290 -1100 -8070
rect -340 -9310 -310 -6710
rect -200 -6770 -170 -6590
rect 650 -6560 680 -6260
rect 790 -6440 820 -6260
rect 790 -6480 820 -6470
rect 650 -6600 680 -6590
rect 590 -6680 620 -6670
rect -200 -7960 -170 -7900
rect -200 -8120 -170 -8060
rect 590 -9240 620 -6710
rect 730 -6680 760 -6670
rect 730 -6770 760 -6710
rect 1520 -6680 1550 -6670
rect 1520 -6830 1550 -6710
rect 1580 -6680 1610 -6260
rect 1580 -6720 1610 -6710
rect 1660 -6680 1690 -6260
rect 2450 -6440 2480 -6260
rect 2450 -6480 2480 -6470
rect 2590 -6560 2620 -6260
rect 3380 -6320 3410 -6260
rect 3380 -6360 3410 -6350
rect 3580 -6320 3610 -6260
rect 3580 -6360 3610 -6350
rect 2590 -6600 2620 -6590
rect 2650 -6560 2680 -6550
rect 1660 -6720 1690 -6710
rect 1720 -6680 1750 -6670
rect 1720 -6830 1750 -6710
rect 2510 -6680 2540 -6670
rect 2510 -6770 2540 -6710
rect 2650 -6770 2680 -6590
rect 3440 -6560 3470 -6550
rect 3440 -6770 3470 -6590
rect 3520 -6560 3550 -6550
rect 3520 -6770 3550 -6590
rect 4310 -6560 4340 -6550
rect 4310 -6770 4340 -6590
rect 4370 -6560 4400 -6260
rect 4510 -6440 4540 -6260
rect 4510 -6480 4540 -6470
rect 4370 -6600 4400 -6590
rect 4450 -6680 4480 -6670
rect 4450 -6770 4480 -6710
rect 5240 -6680 5270 -6670
rect 5240 -6830 5270 -6710
rect 5300 -6680 5330 -6260
rect 5300 -6720 5330 -6710
rect 5380 -6680 5410 -6260
rect 6170 -6440 6200 -6260
rect 6170 -6480 6200 -6470
rect 6310 -6560 6340 -6260
rect 7100 -6320 7130 -6260
rect 7100 -6360 7130 -6350
rect 7300 -6320 7330 -6260
rect 7300 -6360 7330 -6350
rect 6310 -6600 6340 -6590
rect 6370 -6560 6400 -6550
rect 5380 -6720 5410 -6710
rect 5440 -6680 5470 -6670
rect 5440 -6830 5470 -6710
rect 6230 -6680 6260 -6670
rect 6230 -6770 6260 -6710
rect 6370 -6770 6400 -6590
rect 7160 -6560 7190 -6550
rect 7160 -6770 7190 -6590
rect 7240 -6560 7270 -6550
rect 7240 -6770 7270 -6590
rect 8030 -6560 8060 -6550
rect 8030 -6770 8060 -6590
rect 8090 -6560 8120 -6260
rect 8230 -6440 8260 -6260
rect 8230 -6480 8260 -6470
rect 8090 -6600 8120 -6590
rect 8170 -6680 8200 -6670
rect 8170 -6770 8200 -6710
rect 8960 -6680 8990 -6670
rect 8960 -6830 8990 -6710
rect 9020 -6680 9050 -6260
rect 9020 -6720 9050 -6710
rect 9100 -6680 9130 -6260
rect 9890 -6440 9920 -6260
rect 9890 -6480 9920 -6470
rect 10030 -6560 10060 -6260
rect 10820 -6320 10850 -6260
rect 10820 -6360 10850 -6350
rect 11020 -6320 11050 -6260
rect 11020 -6360 11050 -6350
rect 10030 -6600 10060 -6590
rect 10090 -6560 10120 -6550
rect 9100 -6720 9130 -6710
rect 9160 -6680 9190 -6670
rect 9160 -6830 9190 -6710
rect 9950 -6680 9980 -6670
rect 9950 -6770 9980 -6710
rect 10090 -6770 10120 -6590
rect 10880 -6560 10910 -6550
rect 10880 -6770 10910 -6590
rect 10960 -6560 10990 -6550
rect 10960 -6770 10990 -6590
rect 11750 -6560 11780 -6550
rect 11750 -6770 11780 -6590
rect 11810 -6560 11840 -6260
rect 11950 -6440 11980 -6260
rect 11950 -6480 11980 -6470
rect 11810 -6600 11840 -6590
rect 11890 -6680 11920 -6670
rect 11890 -6770 11920 -6710
rect 12680 -6680 12710 -6670
rect 12680 -6830 12710 -6710
rect 12740 -6680 12770 -6260
rect 12740 -6720 12770 -6710
rect 12820 -6680 12850 -6260
rect 13610 -6440 13640 -6260
rect 13610 -6480 13640 -6470
rect 13750 -6560 13780 -6260
rect 14540 -6320 14570 -6260
rect 14680 -6310 14710 2480
rect 14800 -300 14830 -290
rect 14800 -3320 14830 -330
rect 14800 -3360 14830 -3350
rect 15470 -300 15500 -170
rect 15590 -240 15640 -230
rect 15590 -270 15600 -240
rect 15630 -270 15640 -240
rect 15590 -280 15640 -270
rect 15470 -6310 15500 -330
rect 15660 -3260 15710 -3250
rect 15660 -3290 15670 -3260
rect 15700 -3290 15710 -3260
rect 15660 -3300 15710 -3290
rect 15660 -3380 15710 -3370
rect 15660 -3410 15670 -3380
rect 15700 -3410 15710 -3380
rect 15660 -3420 15710 -3410
rect 15660 -3500 15710 -3490
rect 15660 -3530 15670 -3500
rect 15700 -3530 15710 -3500
rect 15660 -3540 15710 -3530
rect 15660 -6260 15710 -6250
rect 15660 -6290 15670 -6260
rect 15700 -6290 15710 -6260
rect 15660 -6300 15710 -6290
rect 14540 -6360 14570 -6350
rect 15660 -6380 15710 -6370
rect 15660 -6410 15670 -6380
rect 15700 -6410 15710 -6380
rect 15660 -6420 15710 -6410
rect 15660 -6500 15710 -6490
rect 15660 -6530 15670 -6500
rect 15700 -6530 15710 -6500
rect 15660 -6540 15710 -6530
rect 13750 -6600 13780 -6590
rect 13810 -6560 13840 -6550
rect 12820 -6720 12850 -6710
rect 12880 -6680 12910 -6670
rect 12880 -6830 12910 -6710
rect 13670 -6680 13700 -6670
rect 13670 -6770 13700 -6710
rect 13810 -6770 13840 -6590
rect 14600 -6560 14630 -6550
rect 14600 -6770 14630 -6590
rect 14740 -6560 14770 -6550
rect 730 -7960 760 -7900
rect 730 -8120 760 -8060
rect 2510 -7960 2540 -7900
rect 2510 -8120 2540 -8060
rect 3440 -7960 3470 -7900
rect 3440 -8120 3470 -8060
rect 3520 -7960 3550 -7900
rect 3520 -8120 3550 -8060
rect 4450 -7960 4480 -7900
rect 4450 -8120 4480 -8060
rect 6230 -7960 6260 -7900
rect 6230 -8120 6260 -8060
rect 7160 -7960 7190 -7900
rect 7160 -8120 7190 -8060
rect 7240 -7960 7270 -7900
rect 7240 -8120 7270 -8060
rect 8170 -7960 8200 -7900
rect 8170 -8120 8200 -8060
rect 9950 -7960 9980 -7900
rect 9950 -8120 9980 -8060
rect 10880 -7960 10910 -7900
rect 10880 -8120 10910 -8060
rect 10960 -7960 10990 -7900
rect 10960 -8120 10990 -8060
rect 11890 -7960 11920 -7900
rect 11890 -8120 11920 -8060
rect 13670 -7960 13700 -7900
rect 13670 -8120 13700 -8060
rect 14600 -7960 14630 -7900
rect 14600 -8120 14630 -8060
rect -340 -9350 -310 -9340
rect -1280 -9370 -1230 -9360
rect -1280 -9400 -1270 -9370
rect -1240 -9400 -1230 -9370
rect -1280 -9410 -1230 -9400
rect -1280 -9490 -1230 -9480
rect -1280 -9520 -1270 -9490
rect -1240 -9520 -1230 -9490
rect -1280 -9530 -1230 -9520
rect -1280 -9610 -1230 -9600
rect -1280 -9640 -1270 -9610
rect -1240 -9640 -1230 -9610
rect -1280 -9650 -1230 -9640
rect -1070 -9670 -1040 -9660
rect -1280 -9730 -1230 -9720
rect -1280 -9760 -1270 -9730
rect -1240 -9760 -1230 -9730
rect -1070 -9760 -1040 -9700
rect -200 -9670 -170 -9250
rect 590 -9310 620 -9250
rect 590 -9350 620 -9340
rect 730 -9550 760 -9250
rect 1520 -9430 1550 -9190
rect 1520 -9470 1550 -9460
rect 1720 -9430 1750 -9190
rect 1720 -9470 1750 -9460
rect 730 -9590 760 -9580
rect 1580 -9550 1610 -9540
rect -200 -9710 -170 -9700
rect -140 -9670 -110 -9660
rect -1280 -9770 -1230 -9760
rect -280 -12480 -250 -9710
rect -140 -9760 -110 -9700
rect 650 -9670 680 -9660
rect 650 -9760 680 -9700
rect 790 -9670 820 -9660
rect 790 -9760 820 -9700
rect 1580 -9760 1610 -9580
rect 1660 -9550 1690 -9540
rect 1660 -9760 1690 -9580
rect 2510 -9550 2540 -9250
rect 2650 -9310 2680 -9250
rect 2650 -9350 2680 -9340
rect 2510 -9590 2540 -9580
rect 2450 -9670 2480 -9660
rect 2450 -9760 2480 -9700
rect 2590 -9670 2620 -9660
rect 2590 -9760 2620 -9700
rect 3380 -9670 3410 -9660
rect 3380 -9760 3410 -9700
rect 3440 -9670 3470 -9250
rect 3440 -9710 3470 -9700
rect 3520 -9670 3550 -9250
rect 4310 -9310 4340 -9250
rect 4310 -9350 4340 -9340
rect 4450 -9550 4480 -9250
rect 5240 -9430 5270 -9190
rect 5240 -9470 5270 -9460
rect 5440 -9430 5470 -9190
rect 5440 -9470 5470 -9460
rect 4450 -9590 4480 -9580
rect 5300 -9550 5330 -9540
rect 3520 -9710 3550 -9700
rect 3580 -9670 3610 -9660
rect 3580 -9760 3610 -9700
rect 4370 -9670 4400 -9660
rect 4370 -9760 4400 -9700
rect 4510 -9670 4540 -9660
rect 4510 -9760 4540 -9700
rect 5300 -9760 5330 -9580
rect 5380 -9550 5410 -9540
rect 5380 -9760 5410 -9580
rect 6230 -9550 6260 -9250
rect 6370 -9310 6400 -9250
rect 6370 -9350 6400 -9340
rect 6230 -9590 6260 -9580
rect 6170 -9670 6200 -9660
rect 6170 -9760 6200 -9700
rect 6310 -9670 6340 -9660
rect 6310 -9760 6340 -9700
rect 7100 -9670 7130 -9660
rect 7100 -9760 7130 -9700
rect 7160 -9670 7190 -9250
rect 7160 -9710 7190 -9700
rect 7240 -9670 7270 -9250
rect 8030 -9310 8060 -9250
rect 8030 -9350 8060 -9340
rect 8170 -9550 8200 -9250
rect 8960 -9430 8990 -9190
rect 8960 -9470 8990 -9460
rect 9160 -9430 9190 -9190
rect 9160 -9470 9190 -9460
rect 8170 -9590 8200 -9580
rect 9020 -9550 9050 -9540
rect 7240 -9710 7270 -9700
rect 7300 -9670 7330 -9660
rect 7300 -9760 7330 -9700
rect 8090 -9670 8120 -9660
rect 8090 -9760 8120 -9700
rect 8230 -9670 8260 -9660
rect 8230 -9760 8260 -9700
rect 9020 -9760 9050 -9580
rect 9100 -9550 9130 -9540
rect 9100 -9760 9130 -9580
rect 9950 -9550 9980 -9250
rect 10090 -9310 10120 -9250
rect 10090 -9350 10120 -9340
rect 9950 -9590 9980 -9580
rect 9890 -9670 9920 -9660
rect 9890 -9760 9920 -9700
rect 10030 -9670 10060 -9660
rect 10030 -9760 10060 -9700
rect 10820 -9670 10850 -9660
rect 10820 -9760 10850 -9700
rect 10880 -9670 10910 -9250
rect 10880 -9710 10910 -9700
rect 10960 -9670 10990 -9250
rect 11750 -9310 11780 -9250
rect 11750 -9350 11780 -9340
rect 11890 -9550 11920 -9250
rect 12680 -9430 12710 -9190
rect 12680 -9470 12710 -9460
rect 12880 -9430 12910 -9190
rect 12880 -9470 12910 -9460
rect 11890 -9590 11920 -9580
rect 12740 -9550 12770 -9540
rect 10960 -9710 10990 -9700
rect 11020 -9670 11050 -9660
rect 11020 -9760 11050 -9700
rect 11810 -9670 11840 -9660
rect 11810 -9760 11840 -9700
rect 11950 -9670 11980 -9660
rect 11950 -9760 11980 -9700
rect 12740 -9760 12770 -9580
rect 12820 -9550 12850 -9540
rect 12820 -9760 12850 -9580
rect 13670 -9550 13700 -9250
rect 13810 -9310 13840 -9250
rect 13810 -9350 13840 -9340
rect 13670 -9590 13700 -9580
rect 13610 -9670 13640 -9660
rect 13610 -9760 13640 -9700
rect 13750 -9670 13780 -9660
rect 13750 -9760 13780 -9700
rect 14540 -9670 14570 -9660
rect 14540 -9760 14570 -9700
rect 14600 -9670 14630 -9250
rect 14740 -9430 14770 -6590
rect 15660 -6620 15710 -6610
rect 15660 -6650 15670 -6620
rect 15700 -6650 15710 -6620
rect 15660 -6660 15710 -6650
rect 15530 -7950 15560 -6730
rect 15660 -6740 15710 -6730
rect 15660 -6770 15670 -6740
rect 15700 -6770 15710 -6740
rect 15660 -6780 15710 -6770
rect 15520 -7960 15570 -7950
rect 15520 -8060 15530 -7960
rect 15560 -8060 15570 -7960
rect 15520 -8070 15570 -8060
rect 15530 -9290 15560 -8070
rect 15660 -9250 15710 -9240
rect 15660 -9280 15670 -9250
rect 15700 -9280 15710 -9250
rect 15660 -9290 15710 -9280
rect 15660 -9370 15710 -9360
rect 15660 -9400 15670 -9370
rect 15700 -9400 15710 -9370
rect 15660 -9410 15710 -9400
rect 14740 -9470 14770 -9460
rect 15660 -9490 15710 -9480
rect 15660 -9520 15670 -9490
rect 15700 -9520 15710 -9490
rect 15660 -9530 15710 -9520
rect 15660 -9610 15710 -9600
rect 15660 -9640 15670 -9610
rect 15700 -9640 15710 -9610
rect 15660 -9650 15710 -9640
rect 14600 -9710 14630 -9700
rect -290 -12490 -240 -12480
rect -290 -12520 -280 -12490
rect -250 -12520 -240 -12490
rect 14680 -12520 14710 -9710
rect -290 -12530 -240 -12520
rect -280 -12560 -250 -12530
rect -280 -12650 -250 -12640
rect 650 -12560 680 -12540
rect 650 -12650 680 -12640
rect 1580 -12560 1610 -12540
rect 1580 -12650 1610 -12640
rect 1660 -12560 1690 -12540
rect 1660 -12650 1690 -12640
rect 2590 -12560 2620 -12540
rect 2590 -12650 2620 -12640
rect 4370 -12560 4400 -12540
rect 4370 -12650 4400 -12640
rect 5300 -12560 5330 -12540
rect 5300 -12650 5330 -12640
rect 5380 -12560 5410 -12540
rect 5380 -12650 5410 -12640
rect 6310 -12560 6340 -12540
rect 6310 -12650 6340 -12640
rect 8090 -12560 8120 -12540
rect 8090 -12650 8120 -12640
rect 9020 -12560 9050 -12540
rect 9020 -12650 9050 -12640
rect 9100 -12560 9130 -12540
rect 9100 -12650 9130 -12640
rect 10030 -12560 10060 -12540
rect 10030 -12650 10060 -12640
rect 11810 -12560 11840 -12540
rect 11810 -12650 11840 -12640
rect 12740 -12560 12770 -12540
rect 12740 -12650 12770 -12640
rect 12820 -12560 12850 -12540
rect 12820 -12650 12850 -12640
rect 13750 -12560 13780 -12540
rect 13750 -12650 13780 -12640
rect 14680 -12560 14710 -12540
rect 14680 -12650 14710 -12640
rect 15470 -12560 15500 -9710
rect 15660 -9730 15710 -9720
rect 15660 -9760 15670 -9730
rect 15700 -9760 15710 -9730
rect 15660 -9770 15710 -9760
rect 15660 -12490 15710 -12480
rect 15660 -12520 15670 -12490
rect 15700 -12520 15710 -12490
rect 15660 -12530 15710 -12520
rect 15470 -12650 15500 -12640
<< via1 >>
rect -1200 -270 -1170 -240
rect -1070 -330 -1040 -300
rect -1270 -3290 -1240 -3260
rect -1270 -3410 -1240 -3380
rect -1270 -3530 -1240 -3500
rect -1270 -6290 -1240 -6260
rect -400 -330 -370 -300
rect -400 -3350 -370 -3320
rect -140 -330 -110 -300
rect 650 -330 680 -300
rect 650 -470 680 -370
rect 1520 -330 1550 -300
rect 1720 -330 1750 -300
rect 730 -470 760 -370
rect 1580 -470 1610 -370
rect 1660 -470 1690 -370
rect 2590 -330 2620 -300
rect 3380 -330 3410 -300
rect 3580 -330 3610 -300
rect 4370 -330 4400 -300
rect 2510 -470 2540 -370
rect 2590 -470 2620 -370
rect 4370 -470 4400 -370
rect 5240 -330 5270 -300
rect 5440 -330 5470 -300
rect 4450 -470 4480 -370
rect 5300 -470 5330 -370
rect 5380 -470 5410 -370
rect 6310 -330 6340 -300
rect 7100 -330 7130 -300
rect 7300 -330 7330 -300
rect 8090 -330 8120 -300
rect 6230 -470 6260 -370
rect 6310 -470 6340 -370
rect 8090 -470 8120 -370
rect 8960 -330 8990 -300
rect 9160 -330 9190 -300
rect 8170 -470 8200 -370
rect 9020 -470 9050 -370
rect 9100 -470 9130 -370
rect 10030 -330 10060 -300
rect 10820 -330 10850 -300
rect 11020 -330 11050 -300
rect 11810 -330 11840 -300
rect 9950 -470 9980 -370
rect 10030 -470 10060 -370
rect 11810 -470 11840 -370
rect 12680 -330 12710 -300
rect 12880 -330 12910 -300
rect 11890 -470 11920 -370
rect 12740 -470 12770 -370
rect 12820 -470 12850 -370
rect 13750 -330 13780 -300
rect 14540 -330 14570 -300
rect 13670 -470 13700 -370
rect 13750 -470 13780 -370
rect -140 -3350 -110 -3320
rect 790 -3350 820 -3320
rect 650 -3470 680 -3440
rect 1580 -3470 1610 -3440
rect 2450 -3350 2480 -3320
rect 1660 -3470 1690 -3440
rect 3380 -3350 3410 -3320
rect 3580 -3350 3610 -3320
rect 2590 -3470 2620 -3440
rect 4510 -3350 4540 -3320
rect 4370 -3470 4400 -3440
rect 5300 -3470 5330 -3440
rect 6170 -3350 6200 -3320
rect 5380 -3470 5410 -3440
rect 7100 -3350 7130 -3320
rect 7300 -3350 7330 -3320
rect 6310 -3470 6340 -3440
rect 8230 -3350 8260 -3320
rect 8090 -3470 8120 -3440
rect 9020 -3470 9050 -3440
rect 9890 -3350 9920 -3320
rect 9100 -3470 9130 -3440
rect 10820 -3350 10850 -3320
rect 11020 -3350 11050 -3320
rect 10030 -3470 10060 -3440
rect 11950 -3350 11980 -3320
rect 11810 -3470 11840 -3440
rect 12740 -3470 12770 -3440
rect 13610 -3350 13640 -3320
rect 12820 -3470 12850 -3440
rect 14540 -3350 14570 -3320
rect 13750 -3470 13780 -3440
rect -140 -6350 -110 -6320
rect -1270 -6410 -1240 -6380
rect -1270 -6530 -1240 -6500
rect -200 -6590 -170 -6560
rect -1270 -6650 -1240 -6620
rect -340 -6710 -310 -6680
rect -1270 -6770 -1240 -6740
rect -1130 -8060 -1100 -7960
rect -1270 -9280 -1240 -9250
rect 790 -6470 820 -6440
rect 650 -6590 680 -6560
rect 590 -6710 620 -6680
rect -200 -8060 -170 -7960
rect 730 -6710 760 -6680
rect 1520 -6710 1550 -6680
rect 1580 -6710 1610 -6680
rect 2450 -6470 2480 -6440
rect 3380 -6350 3410 -6320
rect 3580 -6350 3610 -6320
rect 2590 -6590 2620 -6560
rect 2650 -6590 2680 -6560
rect 1660 -6710 1690 -6680
rect 1720 -6710 1750 -6680
rect 2510 -6710 2540 -6680
rect 3440 -6590 3470 -6560
rect 3520 -6590 3550 -6560
rect 4310 -6590 4340 -6560
rect 4510 -6470 4540 -6440
rect 4370 -6590 4400 -6560
rect 4450 -6710 4480 -6680
rect 5240 -6710 5270 -6680
rect 5300 -6710 5330 -6680
rect 6170 -6470 6200 -6440
rect 7100 -6350 7130 -6320
rect 7300 -6350 7330 -6320
rect 6310 -6590 6340 -6560
rect 6370 -6590 6400 -6560
rect 5380 -6710 5410 -6680
rect 5440 -6710 5470 -6680
rect 6230 -6710 6260 -6680
rect 7160 -6590 7190 -6560
rect 7240 -6590 7270 -6560
rect 8030 -6590 8060 -6560
rect 8230 -6470 8260 -6440
rect 8090 -6590 8120 -6560
rect 8170 -6710 8200 -6680
rect 8960 -6710 8990 -6680
rect 9020 -6710 9050 -6680
rect 9890 -6470 9920 -6440
rect 10820 -6350 10850 -6320
rect 11020 -6350 11050 -6320
rect 10030 -6590 10060 -6560
rect 10090 -6590 10120 -6560
rect 9100 -6710 9130 -6680
rect 9160 -6710 9190 -6680
rect 9950 -6710 9980 -6680
rect 10880 -6590 10910 -6560
rect 10960 -6590 10990 -6560
rect 11750 -6590 11780 -6560
rect 11950 -6470 11980 -6440
rect 11810 -6590 11840 -6560
rect 11890 -6710 11920 -6680
rect 12680 -6710 12710 -6680
rect 12740 -6710 12770 -6680
rect 13610 -6470 13640 -6440
rect 14800 -330 14830 -300
rect 14800 -3350 14830 -3320
rect 15600 -270 15630 -240
rect 15470 -330 15500 -300
rect 15670 -3290 15700 -3260
rect 15670 -3410 15700 -3380
rect 15670 -3530 15700 -3500
rect 15670 -6290 15700 -6260
rect 14540 -6350 14570 -6320
rect 15670 -6410 15700 -6380
rect 15670 -6530 15700 -6500
rect 13750 -6590 13780 -6560
rect 13810 -6590 13840 -6560
rect 12820 -6710 12850 -6680
rect 12880 -6710 12910 -6680
rect 13670 -6710 13700 -6680
rect 14600 -6590 14630 -6560
rect 14740 -6590 14770 -6560
rect 730 -8060 760 -7960
rect 2510 -8060 2540 -7960
rect 3440 -8060 3470 -7960
rect 3520 -8060 3550 -7960
rect 4450 -8060 4480 -7960
rect 6230 -8060 6260 -7960
rect 7160 -8060 7190 -7960
rect 7240 -8060 7270 -7960
rect 8170 -8060 8200 -7960
rect 9950 -8060 9980 -7960
rect 10880 -8060 10910 -7960
rect 10960 -8060 10990 -7960
rect 11890 -8060 11920 -7960
rect 13670 -8060 13700 -7960
rect 14600 -8060 14630 -7960
rect -340 -9340 -310 -9310
rect -1270 -9400 -1240 -9370
rect -1270 -9520 -1240 -9490
rect -1270 -9640 -1240 -9610
rect -1070 -9700 -1040 -9670
rect -1270 -9760 -1240 -9730
rect 590 -9340 620 -9310
rect 1520 -9460 1550 -9430
rect 1720 -9460 1750 -9430
rect 730 -9580 760 -9550
rect 1580 -9580 1610 -9550
rect -200 -9700 -170 -9670
rect -140 -9700 -110 -9670
rect 650 -9700 680 -9670
rect 790 -9700 820 -9670
rect 1660 -9580 1690 -9550
rect 2650 -9340 2680 -9310
rect 2510 -9580 2540 -9550
rect 2450 -9700 2480 -9670
rect 2590 -9700 2620 -9670
rect 3380 -9700 3410 -9670
rect 3440 -9700 3470 -9670
rect 4310 -9340 4340 -9310
rect 5240 -9460 5270 -9430
rect 5440 -9460 5470 -9430
rect 4450 -9580 4480 -9550
rect 5300 -9580 5330 -9550
rect 3520 -9700 3550 -9670
rect 3580 -9700 3610 -9670
rect 4370 -9700 4400 -9670
rect 4510 -9700 4540 -9670
rect 5380 -9580 5410 -9550
rect 6370 -9340 6400 -9310
rect 6230 -9580 6260 -9550
rect 6170 -9700 6200 -9670
rect 6310 -9700 6340 -9670
rect 7100 -9700 7130 -9670
rect 7160 -9700 7190 -9670
rect 8030 -9340 8060 -9310
rect 8960 -9460 8990 -9430
rect 9160 -9460 9190 -9430
rect 8170 -9580 8200 -9550
rect 9020 -9580 9050 -9550
rect 7240 -9700 7270 -9670
rect 7300 -9700 7330 -9670
rect 8090 -9700 8120 -9670
rect 8230 -9700 8260 -9670
rect 9100 -9580 9130 -9550
rect 10090 -9340 10120 -9310
rect 9950 -9580 9980 -9550
rect 9890 -9700 9920 -9670
rect 10030 -9700 10060 -9670
rect 10820 -9700 10850 -9670
rect 10880 -9700 10910 -9670
rect 11750 -9340 11780 -9310
rect 12680 -9460 12710 -9430
rect 12880 -9460 12910 -9430
rect 11890 -9580 11920 -9550
rect 12740 -9580 12770 -9550
rect 10960 -9700 10990 -9670
rect 11020 -9700 11050 -9670
rect 11810 -9700 11840 -9670
rect 11950 -9700 11980 -9670
rect 12820 -9580 12850 -9550
rect 13810 -9340 13840 -9310
rect 13670 -9580 13700 -9550
rect 13610 -9700 13640 -9670
rect 13750 -9700 13780 -9670
rect 14540 -9700 14570 -9670
rect 15670 -6650 15700 -6620
rect 15670 -6770 15700 -6740
rect 15530 -8060 15560 -7960
rect 15670 -9280 15700 -9250
rect 15670 -9400 15700 -9370
rect 14740 -9460 14770 -9430
rect 15670 -9520 15700 -9490
rect 15670 -9640 15700 -9610
rect 14600 -9700 14630 -9670
rect -280 -12640 -250 -12560
rect 650 -12640 680 -12560
rect 1580 -12640 1610 -12560
rect 1660 -12640 1690 -12560
rect 2590 -12640 2620 -12560
rect 4370 -12640 4400 -12560
rect 5300 -12640 5330 -12560
rect 5380 -12640 5410 -12560
rect 6310 -12640 6340 -12560
rect 8090 -12640 8120 -12560
rect 9020 -12640 9050 -12560
rect 9100 -12640 9130 -12560
rect 10030 -12640 10060 -12560
rect 11810 -12640 11840 -12560
rect 12740 -12640 12770 -12560
rect 12820 -12640 12850 -12560
rect 13750 -12640 13780 -12560
rect 14680 -12640 14710 -12560
rect 15670 -9760 15700 -9730
rect 15670 -12520 15700 -12490
rect 15470 -12640 15500 -12560
<< metal2 >>
rect -1270 -270 -1200 -240
rect -1170 -270 15600 -240
rect 15630 -270 15700 -240
rect -1280 -330 -1070 -300
rect -1040 -330 -400 -300
rect -370 -330 -140 -300
rect -110 -330 650 -300
rect 680 -330 1520 -300
rect 1550 -330 1720 -300
rect 1750 -330 2590 -300
rect 2620 -330 3380 -300
rect 3410 -330 3580 -300
rect 3610 -330 4370 -300
rect 4400 -330 5240 -300
rect 5270 -330 5440 -300
rect 5470 -330 6310 -300
rect 6340 -330 7100 -300
rect 7130 -330 7300 -300
rect 7330 -330 8090 -300
rect 8120 -330 8960 -300
rect 8990 -330 9160 -300
rect 9190 -330 10030 -300
rect 10060 -330 10820 -300
rect 10850 -330 11020 -300
rect 11050 -330 11810 -300
rect 11840 -330 12680 -300
rect 12710 -330 12880 -300
rect 12910 -330 13750 -300
rect 13780 -330 14540 -300
rect 14570 -330 14800 -300
rect 14830 -330 15470 -300
rect 15500 -330 15710 -300
rect -1380 -380 650 -370
rect -1380 -460 -1370 -380
rect -1290 -460 650 -380
rect -1380 -470 650 -460
rect 680 -470 730 -370
rect 760 -470 1580 -370
rect 1610 -470 1660 -370
rect 1690 -470 2510 -370
rect 2540 -470 2590 -370
rect 2620 -470 4370 -370
rect 4400 -470 4450 -370
rect 4480 -470 5300 -370
rect 5330 -470 5380 -370
rect 5410 -470 6230 -370
rect 6260 -470 6310 -370
rect 6340 -470 8090 -370
rect 8120 -470 8170 -370
rect 8200 -470 9020 -370
rect 9050 -470 9100 -370
rect 9130 -470 9950 -370
rect 9980 -470 10030 -370
rect 10060 -470 11810 -370
rect 11840 -470 11890 -370
rect 11920 -470 12740 -370
rect 12770 -470 12820 -370
rect 12850 -470 13670 -370
rect 13700 -470 13750 -370
rect 13780 -470 15710 -370
rect -1280 -3290 -1270 -3260
rect -1240 -3290 15670 -3260
rect 15700 -3290 15710 -3260
rect -1270 -3350 -400 -3320
rect -370 -3350 -140 -3320
rect -110 -3350 790 -3320
rect 820 -3350 2450 -3320
rect 2480 -3350 3380 -3320
rect 3410 -3350 3580 -3320
rect 3610 -3350 4510 -3320
rect 4540 -3350 6170 -3320
rect 6200 -3350 7100 -3320
rect 7130 -3350 7300 -3320
rect 7330 -3350 8230 -3320
rect 8260 -3350 9890 -3320
rect 9920 -3350 10820 -3320
rect 10850 -3350 11020 -3320
rect 11050 -3350 11950 -3320
rect 11980 -3350 13610 -3320
rect 13640 -3350 14540 -3320
rect 14570 -3350 14800 -3320
rect 14830 -3350 15700 -3320
rect -1280 -3410 -1270 -3380
rect -1240 -3410 15670 -3380
rect 15700 -3410 15710 -3380
rect -1270 -3470 650 -3440
rect 680 -3470 1580 -3440
rect 1610 -3470 1660 -3440
rect 1690 -3470 2590 -3440
rect 2620 -3470 4370 -3440
rect 4400 -3470 5300 -3440
rect 5330 -3470 5380 -3440
rect 5410 -3470 6310 -3440
rect 6340 -3470 8090 -3440
rect 8120 -3470 9020 -3440
rect 9050 -3470 9100 -3440
rect 9130 -3470 10030 -3440
rect 10060 -3470 11810 -3440
rect 11840 -3470 12740 -3440
rect 12770 -3470 12820 -3440
rect 12850 -3470 13750 -3440
rect 13780 -3470 15700 -3440
rect -1280 -3530 -1270 -3500
rect -1240 -3530 15670 -3500
rect 15700 -3530 15710 -3500
rect -1280 -6290 -1270 -6260
rect -1240 -6290 15670 -6260
rect 15700 -6290 15710 -6260
rect -1280 -6350 -140 -6320
rect -110 -6350 3380 -6320
rect 3410 -6350 3580 -6320
rect 3610 -6350 7100 -6320
rect 7130 -6350 7300 -6320
rect 7330 -6350 10820 -6320
rect 10850 -6350 11020 -6320
rect 11050 -6350 14540 -6320
rect 14570 -6350 15710 -6320
rect -1280 -6410 -1270 -6380
rect -1240 -6410 15670 -6380
rect 15700 -6410 15710 -6380
rect -1280 -6470 790 -6440
rect 820 -6470 2450 -6440
rect 2480 -6470 4510 -6440
rect 4540 -6470 6170 -6440
rect 6200 -6470 8230 -6440
rect 8260 -6470 9890 -6440
rect 9920 -6470 11950 -6440
rect 11980 -6470 13610 -6440
rect 13640 -6470 15710 -6440
rect -1280 -6530 -1270 -6500
rect -1240 -6530 15670 -6500
rect 15700 -6530 15710 -6500
rect -1280 -6590 -200 -6560
rect -170 -6590 650 -6560
rect 680 -6590 2590 -6560
rect 2620 -6590 2650 -6560
rect 2680 -6590 3440 -6560
rect 3470 -6590 3520 -6560
rect 3550 -6590 4310 -6560
rect 4340 -6590 4370 -6560
rect 4400 -6590 6310 -6560
rect 6340 -6590 6370 -6560
rect 6400 -6590 7160 -6560
rect 7190 -6590 7240 -6560
rect 7270 -6590 8030 -6560
rect 8060 -6590 8090 -6560
rect 8120 -6590 10030 -6560
rect 10060 -6590 10090 -6560
rect 10120 -6590 10880 -6560
rect 10910 -6590 10960 -6560
rect 10990 -6590 11750 -6560
rect 11780 -6590 11810 -6560
rect 11840 -6590 13750 -6560
rect 13780 -6590 13810 -6560
rect 13840 -6590 14600 -6560
rect 14630 -6590 14740 -6560
rect 14770 -6590 15710 -6560
rect -1280 -6650 -1270 -6620
rect -1240 -6650 15670 -6620
rect 15700 -6650 15710 -6620
rect -1280 -6710 -340 -6680
rect -310 -6710 590 -6680
rect 620 -6710 730 -6680
rect 760 -6710 1520 -6680
rect 1550 -6710 1580 -6680
rect 1610 -6710 1660 -6680
rect 1690 -6710 1720 -6680
rect 1750 -6710 2510 -6680
rect 2540 -6710 4450 -6680
rect 4480 -6710 5240 -6680
rect 5270 -6710 5300 -6680
rect 5330 -6710 5380 -6680
rect 5410 -6710 5440 -6680
rect 5470 -6710 6230 -6680
rect 6260 -6710 8170 -6680
rect 8200 -6710 8960 -6680
rect 8990 -6710 9020 -6680
rect 9050 -6710 9100 -6680
rect 9130 -6710 9160 -6680
rect 9190 -6710 9950 -6680
rect 9980 -6710 11890 -6680
rect 11920 -6710 12680 -6680
rect 12710 -6710 12740 -6680
rect 12770 -6710 12820 -6680
rect 12850 -6710 12880 -6680
rect 12910 -6710 13670 -6680
rect 13700 -6710 15710 -6680
rect -1280 -6770 -1270 -6740
rect -1240 -6770 15670 -6740
rect 15700 -6770 15710 -6740
rect -1280 -8060 -1130 -7960
rect -1100 -8060 -200 -7960
rect -170 -8060 730 -7960
rect 760 -8060 2510 -7960
rect 2540 -8060 3440 -7960
rect 3470 -8060 3520 -7960
rect 3550 -8060 4450 -7960
rect 4480 -8060 6230 -7960
rect 6260 -8060 7160 -7960
rect 7190 -8060 7240 -7960
rect 7270 -8060 8170 -7960
rect 8200 -8060 9950 -7960
rect 9980 -8060 10880 -7960
rect 10910 -8060 10960 -7960
rect 10990 -8060 11890 -7960
rect 11920 -8060 13670 -7960
rect 13700 -8060 14600 -7960
rect 14630 -8060 15530 -7960
rect 15560 -7970 15810 -7960
rect 15560 -8050 15720 -7970
rect 15800 -8050 15810 -7970
rect 15560 -8060 15810 -8050
rect -1280 -9280 -1270 -9250
rect -1240 -9280 15670 -9250
rect 15700 -9280 15710 -9250
rect -1270 -9340 -340 -9310
rect -310 -9340 590 -9310
rect 620 -9340 2650 -9310
rect 2680 -9340 4310 -9310
rect 4340 -9340 6370 -9310
rect 6400 -9340 8030 -9310
rect 8060 -9340 10090 -9310
rect 10120 -9340 11750 -9310
rect 11780 -9340 13810 -9310
rect 13840 -9340 15700 -9310
rect -1280 -9400 -1270 -9370
rect -1240 -9400 15670 -9370
rect 15700 -9400 15710 -9370
rect -1270 -9460 1520 -9430
rect 1550 -9460 1720 -9430
rect 1750 -9460 5240 -9430
rect 5270 -9460 5440 -9430
rect 5470 -9460 8960 -9430
rect 8990 -9460 9160 -9430
rect 9190 -9460 12680 -9430
rect 12710 -9460 12880 -9430
rect 12910 -9460 14740 -9430
rect 14770 -9460 15700 -9430
rect -1280 -9520 -1270 -9490
rect -1240 -9520 15670 -9490
rect 15700 -9520 15710 -9490
rect -1280 -9580 730 -9550
rect 760 -9580 1580 -9550
rect 1610 -9580 1660 -9550
rect 1690 -9580 2510 -9550
rect 2540 -9580 4450 -9550
rect 4480 -9580 5300 -9550
rect 5330 -9580 5380 -9550
rect 5410 -9580 6230 -9550
rect 6260 -9580 8170 -9550
rect 8200 -9580 9020 -9550
rect 9050 -9580 9100 -9550
rect 9130 -9580 9950 -9550
rect 9980 -9580 11890 -9550
rect 11920 -9580 12740 -9550
rect 12770 -9580 12820 -9550
rect 12850 -9580 13670 -9550
rect 13700 -9580 15700 -9550
rect -1280 -9640 -1270 -9610
rect -1240 -9640 15670 -9610
rect 15700 -9640 15710 -9610
rect -1270 -9700 -1070 -9670
rect -1040 -9700 -200 -9670
rect -170 -9700 -140 -9670
rect -110 -9700 650 -9670
rect 680 -9700 790 -9670
rect 820 -9700 2450 -9670
rect 2480 -9700 2590 -9670
rect 2620 -9700 3380 -9670
rect 3410 -9700 3440 -9670
rect 3470 -9700 3520 -9670
rect 3550 -9700 3580 -9670
rect 3610 -9700 4370 -9670
rect 4400 -9700 4510 -9670
rect 4540 -9700 6170 -9670
rect 6200 -9700 6310 -9670
rect 6340 -9700 7100 -9670
rect 7130 -9700 7160 -9670
rect 7190 -9700 7240 -9670
rect 7270 -9700 7300 -9670
rect 7330 -9700 8090 -9670
rect 8120 -9700 8230 -9670
rect 8260 -9700 9890 -9670
rect 9920 -9700 10030 -9670
rect 10060 -9700 10820 -9670
rect 10850 -9700 10880 -9670
rect 10910 -9700 10960 -9670
rect 10990 -9700 11020 -9670
rect 11050 -9700 11810 -9670
rect 11840 -9700 11950 -9670
rect 11980 -9700 13610 -9670
rect 13640 -9700 13750 -9670
rect 13780 -9700 14540 -9670
rect 14570 -9700 14600 -9670
rect 14630 -9700 15700 -9670
rect -1280 -9760 -1270 -9730
rect -1240 -9760 15670 -9730
rect 15700 -9760 15710 -9730
rect -1230 -12520 -1200 -12490
rect -1170 -12520 15670 -12490
rect 15700 -12520 15710 -12490
rect -1380 -12560 15710 -12550
rect -1380 -12640 -1370 -12560
rect -1290 -12640 -280 -12560
rect -250 -12640 650 -12560
rect 680 -12640 1580 -12560
rect 1610 -12640 1660 -12560
rect 1690 -12640 2590 -12560
rect 2620 -12640 4370 -12560
rect 4400 -12640 5300 -12560
rect 5330 -12640 5380 -12560
rect 5410 -12640 6310 -12560
rect 6340 -12640 8090 -12560
rect 8120 -12640 9020 -12560
rect 9050 -12640 9100 -12560
rect 9130 -12640 10030 -12560
rect 10060 -12640 11810 -12560
rect 11840 -12640 12740 -12560
rect 12770 -12640 12820 -12560
rect 12850 -12640 13750 -12560
rect 13780 -12640 14680 -12560
rect 14710 -12640 15470 -12560
rect 15500 -12640 15710 -12560
rect -1380 -12650 15710 -12640
<< via2 >>
rect -1370 -460 -1290 -380
rect 15720 -8050 15800 -7970
rect -1370 -12640 -1290 -12560
<< metal3 >>
rect -1380 -380 -1280 2700
rect -1380 -460 -1370 -380
rect -1290 -460 -1280 -380
rect -1380 -12560 -1280 -460
rect -1380 -12640 -1370 -12560
rect -1290 -12640 -1280 -12560
rect -1380 -12650 -1280 -12640
rect 15710 -7970 15810 2600
rect 15710 -8050 15720 -7970
rect 15800 -8050 15810 -7970
rect 15710 -12650 15810 -8050
use p1_8  p1_8_54
timestamp 1633696558
transform 1 0 -790 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_55
timestamp 1633696558
transform 1 0 140 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_56
timestamp 1633696558
transform 1 0 1070 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_67
timestamp 1633696558
transform -1 0 2200 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_68
timestamp 1633696558
transform -1 0 3130 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_69
timestamp 1633696558
transform 1 0 3860 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_70
timestamp 1633696558
transform 1 0 4790 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_71
timestamp 1633696558
transform -1 0 5920 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_62
timestamp 1633696558
transform -1 0 6850 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_63
timestamp 1633696558
transform 1 0 7580 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_64
timestamp 1633696558
transform 1 0 8510 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_65
timestamp 1633696558
transform -1 0 9640 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_66
timestamp 1633696558
transform -1 0 10570 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_57
timestamp 1633696558
transform 1 0 11300 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_58
timestamp 1633696558
transform 1 0 12230 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_59
timestamp 1633696558
transform -1 0 13360 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_60
timestamp 1633696558
transform -1 0 14290 0 -1 -9850
box -370 -140 570 2690
use p1_8  p1_8_61
timestamp 1633696558
transform -1 0 15220 0 -1 -9850
box -370 -140 570 2690
use n1_8  n1_8_0
timestamp 1634082396
transform 1 0 -5360 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_16
timestamp 1634082396
transform 1 0 -6290 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_19
timestamp 1634082396
transform 1 0 -5360 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_18
timestamp 1634082396
transform 1 0 -6290 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_1
timestamp 1634082396
transform 1 0 -4430 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_20
timestamp 1634082396
transform 1 0 -4430 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_3
timestamp 1634082396
transform -1 0 7700 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_31
timestamp 1634082396
transform -1 0 7700 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_2
timestamp 1634082396
transform -1 0 8630 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_32
timestamp 1634082396
transform -1 0 8630 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_5
timestamp 1634082396
transform 1 0 -1640 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_33
timestamp 1634082396
transform 1 0 -1640 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_4
timestamp 1634082396
transform 1 0 -710 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_34
timestamp 1634082396
transform 1 0 -710 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_6
timestamp 1634082396
transform -1 0 11420 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_35
timestamp 1634082396
transform -1 0 11420 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_7
timestamp 1634082396
transform -1 0 12350 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_26
timestamp 1634082396
transform -1 0 12350 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_10
timestamp 1634082396
transform 1 0 2080 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_27
timestamp 1634082396
transform 1 0 2080 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_8
timestamp 1634082396
transform 1 0 3010 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_28
timestamp 1634082396
transform 1 0 3010 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_9
timestamp 1634082396
transform -1 0 15140 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_29
timestamp 1634082396
transform -1 0 15140 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_13
timestamp 1634082396
transform -1 0 16070 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_30
timestamp 1634082396
transform -1 0 16070 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_14
timestamp 1634082396
transform 1 0 5800 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_21
timestamp 1634082396
transform 1 0 5800 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_11
timestamp 1634082396
transform 1 0 6730 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_22
timestamp 1634082396
transform 1 0 6730 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_12
timestamp 1634082396
transform -1 0 18860 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_23
timestamp 1634082396
transform -1 0 18860 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_15
timestamp 1634082396
transform -1 0 19790 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_24
timestamp 1634082396
transform -1 0 19790 0 -1 -1350
box 5130 6720 6070 7950
use n1_8  n1_8_17
timestamp 1634082396
transform -1 0 20720 0 1 -14670
box 5130 6720 6070 7950
use n1_8  n1_8_25
timestamp 1634082396
transform -1 0 20720 0 -1 -1350
box 5130 6720 6070 7950
use p1_8  p1_8_48
timestamp 1633696558
transform 1 0 -790 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_5
timestamp 1633696558
transform 1 0 140 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_4
timestamp 1633696558
transform 1 0 1070 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_7
timestamp 1633696558
transform -1 0 2200 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_6
timestamp 1633696558
transform -1 0 3130 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_13
timestamp 1633696558
transform 1 0 3860 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_12
timestamp 1633696558
transform 1 0 4790 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_14
timestamp 1633696558
transform -1 0 5920 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_15
timestamp 1633696558
transform -1 0 6850 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_26
timestamp 1633696558
transform 1 0 7580 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_24
timestamp 1633696558
transform 1 0 8510 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_25
timestamp 1633696558
transform -1 0 9640 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_29
timestamp 1633696558
transform -1 0 10570 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_30
timestamp 1633696558
transform 1 0 11300 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_27
timestamp 1633696558
transform 1 0 12230 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_28
timestamp 1633696558
transform -1 0 13360 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_31
timestamp 1633696558
transform -1 0 14290 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_51
timestamp 1633696558
transform -1 0 15220 0 1 -6170
box -370 -140 570 2690
use p1_8  p1_8_49
timestamp 1633696558
transform 1 0 -790 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_2
timestamp 1633696558
transform 1 0 140 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_3
timestamp 1633696558
transform 1 0 1070 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_9
timestamp 1633696558
transform -1 0 2200 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_8
timestamp 1633696558
transform -1 0 3130 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_17
timestamp 1633696558
transform 1 0 3860 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_16
timestamp 1633696558
transform 1 0 4790 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_18
timestamp 1633696558
transform -1 0 5920 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_19
timestamp 1633696558
transform -1 0 6850 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_34
timestamp 1633696558
transform 1 0 7580 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_32
timestamp 1633696558
transform 1 0 8510 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_33
timestamp 1633696558
transform -1 0 9640 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_37
timestamp 1633696558
transform -1 0 10570 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_38
timestamp 1633696558
transform 1 0 11300 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_35
timestamp 1633696558
transform 1 0 12230 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_36
timestamp 1633696558
transform -1 0 13360 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_39
timestamp 1633696558
transform -1 0 14290 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_52
timestamp 1633696558
transform -1 0 15220 0 1 -3170
box -370 -140 570 2690
use p1_8  p1_8_50
timestamp 1633696558
transform 1 0 -790 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_0
timestamp 1633696558
transform 1 0 140 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_1
timestamp 1633696558
transform -1 0 1270 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_10
timestamp 1633696558
transform 1 0 2000 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_11
timestamp 1633696558
transform -1 0 3130 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_20
timestamp 1633696558
transform 1 0 3860 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_21
timestamp 1633696558
transform -1 0 4990 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_22
timestamp 1633696558
transform 1 0 5720 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_23
timestamp 1633696558
transform -1 0 6850 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_42
timestamp 1633696558
transform 1 0 7580 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_41
timestamp 1633696558
transform -1 0 8710 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_40
timestamp 1633696558
transform 1 0 9440 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_46
timestamp 1633696558
transform -1 0 10570 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_45
timestamp 1633696558
transform 1 0 11300 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_43
timestamp 1633696558
transform -1 0 12430 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_44
timestamp 1633696558
transform 1 0 13160 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_47
timestamp 1633696558
transform -1 0 14290 0 1 -150
box -370 -140 570 2690
use p1_8  p1_8_53
timestamp 1633696558
transform -1 0 15220 0 1 -150
box -370 -140 570 2690
<< labels >>
rlabel metal2 -1270 -3470 -1240 -3440 1 x
rlabel metal2 -1280 -6590 -1270 -6560 3 ym
rlabel metal2 -1280 -6710 -1270 -6680 3 yp
rlabel metal2 -1270 -9700 -1240 -9670 1 z
rlabel metal2 -1280 -6470 -1270 -6440 1 inm
port 1 n
rlabel metal2 -1280 -6350 -1270 -6320 1 inp
port 2 n
rlabel metal2 -1280 -9580 -1270 -9550 1 out
port 3 n
rlabel metal2 -1280 -330 -1270 -300 1 ibias
port 4 n
rlabel metal2 -1280 -470 -1270 -370 1 vdda
port 5 n
rlabel metal2 -1280 -8060 -1270 -7960 1 gnd
port 6 n
rlabel metal1 650 2490 13780 2520 1 a
<< end >>
