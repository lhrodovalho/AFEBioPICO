magic
tech sky130A
magscale 1 2
timestamp 1638148091
<< pwell >>
rect 1094 934 1226 1066
<< psubdiff >>
rect 1120 960 1200 1040
<< locali >>
rect 1120 1017 1200 31920
rect 1120 983 1143 1017
rect 1177 983 1200 1017
rect 1120 960 1200 983
rect 28800 1017 28880 31920
rect 28800 983 28823 1017
rect 28857 983 28880 1017
rect 28800 960 28880 983
<< viali >>
rect 1143 983 1177 1017
rect 28823 983 28857 1017
<< metal1 >>
rect 1120 1026 1200 1040
rect 1120 974 1134 1026
rect 1186 974 1200 1026
rect 1120 960 1200 974
rect 28800 1026 28880 1040
rect 28800 974 28814 1026
rect 28866 974 28880 1026
rect 28800 960 28880 974
<< via1 >>
rect 1134 1017 1186 1026
rect 1134 983 1143 1017
rect 1143 983 1177 1017
rect 1177 983 1186 1017
rect 1134 974 1186 983
rect 28814 1017 28866 1026
rect 28814 983 28823 1017
rect 28823 983 28857 1017
rect 28857 983 28866 1017
rect 28814 974 28866 983
<< metal2 >>
rect 0 31908 1040 31920
rect 0 31852 12 31908
rect 68 31852 332 31908
rect 388 31852 652 31908
rect 708 31852 972 31908
rect 1028 31852 1040 31908
rect 0 31840 1040 31852
rect 28960 31908 30000 31920
rect 28960 31852 28972 31908
rect 29028 31852 29292 31908
rect 29348 31852 29612 31908
rect 29668 31852 29932 31908
rect 29988 31852 30000 31908
rect 28960 31840 30000 31852
rect 0 31748 1040 31760
rect 0 31692 12 31748
rect 68 31692 332 31748
rect 388 31692 652 31748
rect 708 31692 972 31748
rect 1028 31692 1040 31748
rect 0 31680 1040 31692
rect 28960 31748 30000 31760
rect 28960 31692 28972 31748
rect 29028 31692 29292 31748
rect 29348 31692 29612 31748
rect 29668 31692 29932 31748
rect 29988 31692 30000 31748
rect 28960 31680 30000 31692
rect 0 31588 1040 31600
rect 0 31532 12 31588
rect 68 31532 332 31588
rect 388 31532 652 31588
rect 708 31532 972 31588
rect 1028 31532 1040 31588
rect 0 31520 1040 31532
rect 28960 31588 30000 31600
rect 28960 31532 28972 31588
rect 29028 31532 29292 31588
rect 29348 31532 29612 31588
rect 29668 31532 29932 31588
rect 29988 31532 30000 31588
rect 28960 31520 30000 31532
rect 0 31428 1040 31440
rect 0 31372 12 31428
rect 68 31372 332 31428
rect 388 31372 652 31428
rect 708 31372 972 31428
rect 1028 31372 1040 31428
rect 0 31360 1040 31372
rect 28960 31428 30000 31440
rect 28960 31372 28972 31428
rect 29028 31372 29292 31428
rect 29348 31372 29612 31428
rect 29668 31372 29932 31428
rect 29988 31372 30000 31428
rect 28960 31360 30000 31372
rect 0 31268 1040 31280
rect 0 31212 12 31268
rect 68 31212 332 31268
rect 388 31212 652 31268
rect 708 31212 972 31268
rect 1028 31212 1040 31268
rect 0 31200 1040 31212
rect 28960 31268 30000 31280
rect 28960 31212 28972 31268
rect 29028 31212 29292 31268
rect 29348 31212 29612 31268
rect 29668 31212 29932 31268
rect 29988 31212 30000 31268
rect 28960 31200 30000 31212
rect 0 31108 1040 31120
rect 0 31052 12 31108
rect 68 31052 332 31108
rect 388 31052 652 31108
rect 708 31052 972 31108
rect 1028 31052 1040 31108
rect 0 31040 1040 31052
rect 28960 31108 30000 31120
rect 28960 31052 28972 31108
rect 29028 31052 29292 31108
rect 29348 31052 29612 31108
rect 29668 31052 29932 31108
rect 29988 31052 30000 31108
rect 28960 31040 30000 31052
rect 0 30948 1040 30960
rect 0 30892 12 30948
rect 68 30892 332 30948
rect 388 30892 652 30948
rect 708 30892 972 30948
rect 1028 30892 1040 30948
rect 0 30880 1040 30892
rect 28960 30948 30000 30960
rect 28960 30892 28972 30948
rect 29028 30892 29292 30948
rect 29348 30892 29612 30948
rect 29668 30892 29932 30948
rect 29988 30892 30000 30948
rect 28960 30880 30000 30892
rect 0 30788 1040 30800
rect 0 30732 12 30788
rect 68 30732 332 30788
rect 388 30732 652 30788
rect 708 30732 972 30788
rect 1028 30732 1040 30788
rect 0 30720 1040 30732
rect 28960 30788 30000 30800
rect 28960 30732 28972 30788
rect 29028 30732 29292 30788
rect 29348 30732 29612 30788
rect 29668 30732 29932 30788
rect 29988 30732 30000 30788
rect 28960 30720 30000 30732
rect 0 30628 1040 30640
rect 0 30572 12 30628
rect 68 30572 332 30628
rect 388 30572 652 30628
rect 708 30572 972 30628
rect 1028 30572 1040 30628
rect 0 30560 1040 30572
rect 28960 30628 30000 30640
rect 28960 30572 28972 30628
rect 29028 30572 29292 30628
rect 29348 30572 29612 30628
rect 29668 30572 29932 30628
rect 29988 30572 30000 30628
rect 28960 30560 30000 30572
rect 0 30468 1040 30480
rect 0 30412 12 30468
rect 68 30412 332 30468
rect 388 30412 652 30468
rect 708 30412 972 30468
rect 1028 30412 1040 30468
rect 0 30400 1040 30412
rect 28960 30468 30000 30480
rect 28960 30412 28972 30468
rect 29028 30412 29292 30468
rect 29348 30412 29612 30468
rect 29668 30412 29932 30468
rect 29988 30412 30000 30468
rect 28960 30400 30000 30412
rect 0 30308 1040 30320
rect 0 30252 12 30308
rect 68 30252 332 30308
rect 388 30252 652 30308
rect 708 30252 972 30308
rect 1028 30252 1040 30308
rect 0 30240 1040 30252
rect 28960 30308 30000 30320
rect 28960 30252 28972 30308
rect 29028 30252 29292 30308
rect 29348 30252 29612 30308
rect 29668 30252 29932 30308
rect 29988 30252 30000 30308
rect 28960 30240 30000 30252
rect 0 30148 1040 30160
rect 0 30092 12 30148
rect 68 30092 332 30148
rect 388 30092 652 30148
rect 708 30092 972 30148
rect 1028 30092 1040 30148
rect 0 30080 1040 30092
rect 28960 30148 30000 30160
rect 28960 30092 28972 30148
rect 29028 30092 29292 30148
rect 29348 30092 29612 30148
rect 29668 30092 29932 30148
rect 29988 30092 30000 30148
rect 28960 30080 30000 30092
rect 0 29988 1040 30000
rect 0 29932 12 29988
rect 68 29932 332 29988
rect 388 29932 652 29988
rect 708 29932 972 29988
rect 1028 29932 1040 29988
rect 0 29920 1040 29932
rect 28960 29988 30000 30000
rect 28960 29932 28972 29988
rect 29028 29932 29292 29988
rect 29348 29932 29612 29988
rect 29668 29932 29932 29988
rect 29988 29932 30000 29988
rect 28960 29920 30000 29932
rect 0 29828 1040 29840
rect 0 29772 12 29828
rect 68 29772 332 29828
rect 388 29772 652 29828
rect 708 29772 972 29828
rect 1028 29772 1040 29828
rect 0 29760 1040 29772
rect 28960 29828 30000 29840
rect 28960 29772 28972 29828
rect 29028 29772 29292 29828
rect 29348 29772 29612 29828
rect 29668 29772 29932 29828
rect 29988 29772 30000 29828
rect 28960 29760 30000 29772
rect 0 29668 1040 29680
rect 0 29612 12 29668
rect 68 29612 332 29668
rect 388 29612 652 29668
rect 708 29612 972 29668
rect 1028 29612 1040 29668
rect 0 29600 1040 29612
rect 28960 29668 30000 29680
rect 28960 29612 28972 29668
rect 29028 29612 29292 29668
rect 29348 29612 29612 29668
rect 29668 29612 29932 29668
rect 29988 29612 30000 29668
rect 28960 29600 30000 29612
rect 0 29508 1040 29520
rect 0 29452 12 29508
rect 68 29452 332 29508
rect 388 29452 652 29508
rect 708 29452 972 29508
rect 1028 29452 1040 29508
rect 0 29440 1040 29452
rect 28960 29508 30000 29520
rect 28960 29452 28972 29508
rect 29028 29452 29292 29508
rect 29348 29452 29612 29508
rect 29668 29452 29932 29508
rect 29988 29452 30000 29508
rect 28960 29440 30000 29452
rect 0 29348 1040 29360
rect 0 29292 12 29348
rect 68 29292 332 29348
rect 388 29292 652 29348
rect 708 29292 972 29348
rect 1028 29292 1040 29348
rect 0 29280 1040 29292
rect 28960 29348 30000 29360
rect 28960 29292 28972 29348
rect 29028 29292 29292 29348
rect 29348 29292 29612 29348
rect 29668 29292 29932 29348
rect 29988 29292 30000 29348
rect 28960 29280 30000 29292
rect 0 29188 1040 29200
rect 0 29132 12 29188
rect 68 29132 332 29188
rect 388 29132 652 29188
rect 708 29132 972 29188
rect 1028 29132 1040 29188
rect 0 29120 1040 29132
rect 0 29028 1040 29040
rect 0 28972 12 29028
rect 68 28972 332 29028
rect 388 28972 652 29028
rect 708 28972 972 29028
rect 1028 28972 1040 29028
rect 0 28960 1040 28972
rect 28960 29028 30000 29040
rect 28960 28972 28972 29028
rect 29028 28972 29292 29028
rect 29348 28972 29612 29028
rect 29668 28972 29932 29028
rect 29988 28972 30000 29028
rect 28960 28960 30000 28972
rect 0 28868 1040 28880
rect 0 28812 12 28868
rect 68 28812 332 28868
rect 388 28812 652 28868
rect 708 28812 972 28868
rect 1028 28812 1040 28868
rect 0 28800 1040 28812
rect 29600 28868 30000 28880
rect 29600 28812 29612 28868
rect 29668 28812 29932 28868
rect 29988 28812 30000 28868
rect 29600 28800 30000 28812
rect 0 28708 1040 28720
rect 0 28652 12 28708
rect 68 28652 332 28708
rect 388 28652 652 28708
rect 708 28652 972 28708
rect 1028 28652 1040 28708
rect 0 28640 1040 28652
rect 28960 28708 30000 28720
rect 28960 28652 28972 28708
rect 29028 28652 29292 28708
rect 29348 28652 29612 28708
rect 29668 28652 29932 28708
rect 29988 28652 30000 28708
rect 28960 28640 30000 28652
rect 0 28548 1040 28560
rect 0 28492 12 28548
rect 68 28492 332 28548
rect 388 28492 652 28548
rect 708 28492 972 28548
rect 1028 28492 1040 28548
rect 0 28480 1040 28492
rect 28960 28548 30000 28560
rect 28960 28492 28972 28548
rect 29028 28492 29292 28548
rect 29348 28492 29612 28548
rect 29668 28492 29932 28548
rect 29988 28492 30000 28548
rect 28960 28480 30000 28492
rect 0 28388 1040 28400
rect 0 28332 12 28388
rect 68 28332 332 28388
rect 388 28332 652 28388
rect 708 28332 972 28388
rect 1028 28332 1040 28388
rect 0 28320 1040 28332
rect 28960 28388 30000 28400
rect 28960 28332 28972 28388
rect 29028 28332 29292 28388
rect 29348 28332 29612 28388
rect 29668 28332 29932 28388
rect 29988 28332 30000 28388
rect 28960 28320 30000 28332
rect 0 28228 1040 28240
rect 0 28172 12 28228
rect 68 28172 332 28228
rect 388 28172 652 28228
rect 708 28172 972 28228
rect 1028 28172 1040 28228
rect 0 28160 1040 28172
rect 28960 28228 30000 28240
rect 28960 28172 28972 28228
rect 29028 28172 29292 28228
rect 29348 28172 29612 28228
rect 29668 28172 29932 28228
rect 29988 28172 30000 28228
rect 28960 28160 30000 28172
rect 0 28068 1040 28080
rect 0 28012 12 28068
rect 68 28012 332 28068
rect 388 28012 652 28068
rect 708 28012 972 28068
rect 1028 28012 1040 28068
rect 0 28000 1040 28012
rect 28960 28068 30000 28080
rect 28960 28012 28972 28068
rect 29028 28012 29292 28068
rect 29348 28012 29612 28068
rect 29668 28012 29932 28068
rect 29988 28012 30000 28068
rect 28960 28000 30000 28012
rect 0 27908 1040 27920
rect 0 27852 12 27908
rect 68 27852 332 27908
rect 388 27852 652 27908
rect 708 27852 972 27908
rect 1028 27852 1040 27908
rect 0 27840 1040 27852
rect 28960 27908 30000 27920
rect 28960 27852 28972 27908
rect 29028 27852 29292 27908
rect 29348 27852 29612 27908
rect 29668 27852 29932 27908
rect 29988 27852 30000 27908
rect 28960 27840 30000 27852
rect 0 27748 1040 27760
rect 0 27692 12 27748
rect 68 27692 332 27748
rect 388 27692 652 27748
rect 708 27692 972 27748
rect 1028 27692 1040 27748
rect 0 27680 1040 27692
rect 28960 27748 30000 27760
rect 28960 27692 28972 27748
rect 29028 27692 29292 27748
rect 29348 27692 29612 27748
rect 29668 27692 29932 27748
rect 29988 27692 30000 27748
rect 28960 27680 30000 27692
rect 0 27588 1040 27600
rect 0 27532 12 27588
rect 68 27532 332 27588
rect 388 27532 652 27588
rect 708 27532 972 27588
rect 1028 27532 1040 27588
rect 0 27520 1040 27532
rect 28960 27588 30000 27600
rect 28960 27532 28972 27588
rect 29028 27532 29292 27588
rect 29348 27532 29612 27588
rect 29668 27532 29932 27588
rect 29988 27532 30000 27588
rect 28960 27520 30000 27532
rect 0 27428 1040 27440
rect 0 27372 12 27428
rect 68 27372 332 27428
rect 388 27372 652 27428
rect 708 27372 972 27428
rect 1028 27372 1040 27428
rect 0 27360 1040 27372
rect 28960 27428 30000 27440
rect 28960 27372 28972 27428
rect 29028 27372 29292 27428
rect 29348 27372 29612 27428
rect 29668 27372 29932 27428
rect 29988 27372 30000 27428
rect 28960 27360 30000 27372
rect 0 27268 1040 27280
rect 0 27212 12 27268
rect 68 27212 332 27268
rect 388 27212 652 27268
rect 708 27212 972 27268
rect 1028 27212 1040 27268
rect 0 27200 1040 27212
rect 28960 27268 30000 27280
rect 28960 27212 28972 27268
rect 29028 27212 29292 27268
rect 29348 27212 29612 27268
rect 29668 27212 29932 27268
rect 29988 27212 30000 27268
rect 28960 27200 30000 27212
rect 0 27108 1040 27120
rect 0 27052 12 27108
rect 68 27052 332 27108
rect 388 27052 652 27108
rect 708 27052 972 27108
rect 1028 27052 1040 27108
rect 0 27040 1040 27052
rect 28960 27108 30000 27120
rect 28960 27052 28972 27108
rect 29028 27052 29292 27108
rect 29348 27052 29612 27108
rect 29668 27052 29932 27108
rect 29988 27052 30000 27108
rect 28960 27040 30000 27052
rect 0 26948 1040 26960
rect 0 26892 12 26948
rect 68 26892 332 26948
rect 388 26892 652 26948
rect 708 26892 972 26948
rect 1028 26892 1040 26948
rect 0 26880 1040 26892
rect 28960 26948 30000 26960
rect 28960 26892 28972 26948
rect 29028 26892 29292 26948
rect 29348 26892 29612 26948
rect 29668 26892 29932 26948
rect 29988 26892 30000 26948
rect 28960 26880 30000 26892
rect 0 26788 1040 26800
rect 0 26732 12 26788
rect 68 26732 332 26788
rect 388 26732 652 26788
rect 708 26732 972 26788
rect 1028 26732 1040 26788
rect 0 26720 1040 26732
rect 28960 26788 30000 26800
rect 28960 26732 28972 26788
rect 29028 26732 29292 26788
rect 29348 26732 29612 26788
rect 29668 26732 29932 26788
rect 29988 26732 30000 26788
rect 28960 26720 30000 26732
rect 0 26628 1040 26640
rect 0 26572 12 26628
rect 68 26572 332 26628
rect 388 26572 652 26628
rect 708 26572 972 26628
rect 1028 26572 1040 26628
rect 0 26560 1040 26572
rect 28960 26628 30000 26640
rect 28960 26572 28972 26628
rect 29028 26572 29292 26628
rect 29348 26572 29612 26628
rect 29668 26572 29932 26628
rect 29988 26572 30000 26628
rect 28960 26560 30000 26572
rect 0 26468 1040 26480
rect 0 26412 12 26468
rect 68 26412 332 26468
rect 388 26412 652 26468
rect 708 26412 972 26468
rect 1028 26412 1040 26468
rect 0 26400 1040 26412
rect 28960 26468 30000 26480
rect 28960 26412 28972 26468
rect 29028 26412 29292 26468
rect 29348 26412 29612 26468
rect 29668 26412 29932 26468
rect 29988 26412 30000 26468
rect 28960 26400 30000 26412
rect 0 26308 1040 26320
rect 0 26252 12 26308
rect 68 26252 332 26308
rect 388 26252 652 26308
rect 708 26252 972 26308
rect 1028 26252 1040 26308
rect 0 26240 1040 26252
rect 29280 26308 30000 26320
rect 29280 26252 29292 26308
rect 29348 26252 29612 26308
rect 29668 26252 29932 26308
rect 29988 26252 30000 26308
rect 29280 26240 30000 26252
rect 0 26148 1040 26160
rect 0 26092 12 26148
rect 68 26092 332 26148
rect 388 26092 652 26148
rect 708 26092 972 26148
rect 1028 26092 1040 26148
rect 0 26080 1040 26092
rect 28960 26148 30000 26160
rect 28960 26092 28972 26148
rect 29028 26092 29292 26148
rect 29348 26092 29612 26148
rect 29668 26092 29932 26148
rect 29988 26092 30000 26148
rect 28960 26080 30000 26092
rect 0 25988 1040 26000
rect 0 25932 12 25988
rect 68 25932 332 25988
rect 388 25932 652 25988
rect 708 25932 972 25988
rect 1028 25932 1040 25988
rect 0 25920 1040 25932
rect 28960 25988 30000 26000
rect 28960 25932 28972 25988
rect 29028 25932 29292 25988
rect 29348 25932 29612 25988
rect 29668 25932 29932 25988
rect 29988 25932 30000 25988
rect 28960 25920 30000 25932
rect 0 25828 1040 25840
rect 0 25772 12 25828
rect 68 25772 332 25828
rect 388 25772 652 25828
rect 708 25772 972 25828
rect 1028 25772 1040 25828
rect 0 25760 1040 25772
rect 28960 25828 30000 25840
rect 28960 25772 28972 25828
rect 29028 25772 29292 25828
rect 29348 25772 29612 25828
rect 29668 25772 29932 25828
rect 29988 25772 30000 25828
rect 28960 25760 30000 25772
rect 0 25668 1040 25680
rect 0 25612 12 25668
rect 68 25612 332 25668
rect 388 25612 652 25668
rect 708 25612 972 25668
rect 1028 25612 1040 25668
rect 0 25600 1040 25612
rect 28960 25668 30000 25680
rect 28960 25612 28972 25668
rect 29028 25612 29292 25668
rect 29348 25612 29612 25668
rect 29668 25612 29932 25668
rect 29988 25612 30000 25668
rect 28960 25600 30000 25612
rect 0 25508 1040 25520
rect 0 25452 12 25508
rect 68 25452 332 25508
rect 388 25452 652 25508
rect 708 25452 972 25508
rect 1028 25452 1040 25508
rect 0 25440 1040 25452
rect 28960 25508 30000 25520
rect 28960 25452 28972 25508
rect 29028 25452 29292 25508
rect 29348 25452 29612 25508
rect 29668 25452 29932 25508
rect 29988 25452 30000 25508
rect 28960 25440 30000 25452
rect 0 25348 1040 25360
rect 0 25292 12 25348
rect 68 25292 332 25348
rect 388 25292 652 25348
rect 708 25292 972 25348
rect 1028 25292 1040 25348
rect 0 25280 1040 25292
rect 28960 25348 30000 25360
rect 28960 25292 28972 25348
rect 29028 25292 29292 25348
rect 29348 25292 29612 25348
rect 29668 25292 29932 25348
rect 29988 25292 30000 25348
rect 28960 25280 30000 25292
rect 0 25188 1040 25200
rect 0 25132 12 25188
rect 68 25132 332 25188
rect 388 25132 652 25188
rect 708 25132 972 25188
rect 1028 25132 1040 25188
rect 0 25120 1040 25132
rect 28960 25188 30000 25200
rect 28960 25132 28972 25188
rect 29028 25132 29292 25188
rect 29348 25132 29612 25188
rect 29668 25132 29932 25188
rect 29988 25132 30000 25188
rect 28960 25120 30000 25132
rect 0 25028 1040 25040
rect 0 24972 12 25028
rect 68 24972 332 25028
rect 388 24972 652 25028
rect 708 24972 972 25028
rect 1028 24972 1040 25028
rect 0 24960 1040 24972
rect 28960 25028 30000 25040
rect 28960 24972 28972 25028
rect 29028 24972 29292 25028
rect 29348 24972 29612 25028
rect 29668 24972 29932 25028
rect 29988 24972 30000 25028
rect 28960 24960 30000 24972
rect 0 24868 1040 24880
rect 0 24812 12 24868
rect 68 24812 332 24868
rect 388 24812 652 24868
rect 708 24812 972 24868
rect 1028 24812 1040 24868
rect 0 24800 1040 24812
rect 28960 24868 30000 24880
rect 28960 24812 28972 24868
rect 29028 24812 29292 24868
rect 29348 24812 29612 24868
rect 29668 24812 29932 24868
rect 29988 24812 30000 24868
rect 28960 24800 30000 24812
rect 0 24708 1040 24720
rect 0 24652 12 24708
rect 68 24652 332 24708
rect 388 24652 652 24708
rect 708 24652 972 24708
rect 1028 24652 1040 24708
rect 0 24640 1040 24652
rect 28960 24708 30000 24720
rect 28960 24652 28972 24708
rect 29028 24652 29292 24708
rect 29348 24652 29612 24708
rect 29668 24652 29932 24708
rect 29988 24652 30000 24708
rect 28960 24640 30000 24652
rect 0 24548 1040 24560
rect 0 24492 12 24548
rect 68 24492 332 24548
rect 388 24492 652 24548
rect 708 24492 972 24548
rect 1028 24492 1040 24548
rect 0 24480 1040 24492
rect 28960 24548 30000 24560
rect 28960 24492 28972 24548
rect 29028 24492 29292 24548
rect 29348 24492 29612 24548
rect 29668 24492 29932 24548
rect 29988 24492 30000 24548
rect 28960 24480 30000 24492
rect 0 24388 1040 24400
rect 0 24332 12 24388
rect 68 24332 332 24388
rect 388 24332 652 24388
rect 708 24332 972 24388
rect 1028 24332 1040 24388
rect 0 24320 1040 24332
rect 28960 24388 30000 24400
rect 28960 24332 28972 24388
rect 29028 24332 29292 24388
rect 29348 24332 29612 24388
rect 29668 24332 29932 24388
rect 29988 24332 30000 24388
rect 28960 24320 30000 24332
rect 0 24228 1040 24240
rect 0 24172 12 24228
rect 68 24172 332 24228
rect 388 24172 652 24228
rect 708 24172 972 24228
rect 1028 24172 1040 24228
rect 0 24160 1040 24172
rect 28960 24228 30000 24240
rect 28960 24172 28972 24228
rect 29028 24172 29292 24228
rect 29348 24172 29612 24228
rect 29668 24172 29932 24228
rect 29988 24172 30000 24228
rect 28960 24160 30000 24172
rect 0 24068 1040 24080
rect 0 24012 12 24068
rect 68 24012 332 24068
rect 388 24012 652 24068
rect 708 24012 972 24068
rect 1028 24012 1040 24068
rect 0 24000 1040 24012
rect 28960 24068 30000 24080
rect 28960 24012 28972 24068
rect 29028 24012 29292 24068
rect 29348 24012 29612 24068
rect 29668 24012 29932 24068
rect 29988 24012 30000 24068
rect 28960 24000 30000 24012
rect 0 23908 1040 23920
rect 0 23852 12 23908
rect 68 23852 332 23908
rect 388 23852 652 23908
rect 708 23852 972 23908
rect 1028 23852 1040 23908
rect 0 23840 1040 23852
rect 28960 23908 30000 23920
rect 28960 23852 28972 23908
rect 29028 23852 29292 23908
rect 29348 23852 29612 23908
rect 29668 23852 29932 23908
rect 29988 23852 30000 23908
rect 28960 23840 30000 23852
rect 0 23748 1040 23760
rect 0 23692 12 23748
rect 68 23692 332 23748
rect 388 23692 652 23748
rect 708 23692 972 23748
rect 1028 23692 1040 23748
rect 0 23680 1040 23692
rect 29600 23748 30000 23760
rect 29600 23692 29612 23748
rect 29668 23692 29932 23748
rect 29988 23692 30000 23748
rect 29600 23680 30000 23692
rect 0 23588 1040 23600
rect 0 23532 12 23588
rect 68 23532 332 23588
rect 388 23532 652 23588
rect 708 23532 972 23588
rect 1028 23532 1040 23588
rect 0 23520 1040 23532
rect 28960 23588 30000 23600
rect 28960 23532 28972 23588
rect 29028 23532 29292 23588
rect 29348 23532 29612 23588
rect 29668 23532 29932 23588
rect 29988 23532 30000 23588
rect 28960 23520 30000 23532
rect 0 23428 1040 23440
rect 0 23372 12 23428
rect 68 23372 332 23428
rect 388 23372 652 23428
rect 708 23372 972 23428
rect 1028 23372 1040 23428
rect 0 23360 1040 23372
rect 0 23268 1040 23280
rect 0 23212 12 23268
rect 68 23212 332 23268
rect 388 23212 652 23268
rect 708 23212 972 23268
rect 1028 23212 1040 23268
rect 0 23200 1040 23212
rect 28960 23268 30000 23280
rect 28960 23212 28972 23268
rect 29028 23212 29292 23268
rect 29348 23212 29612 23268
rect 29668 23212 29932 23268
rect 29988 23212 30000 23268
rect 28960 23200 30000 23212
rect 0 23108 1040 23120
rect 0 23052 12 23108
rect 68 23052 332 23108
rect 388 23052 652 23108
rect 708 23052 972 23108
rect 1028 23052 1040 23108
rect 0 23040 1040 23052
rect 28960 23108 30000 23120
rect 28960 23052 28972 23108
rect 29028 23052 29292 23108
rect 29348 23052 29612 23108
rect 29668 23052 29932 23108
rect 29988 23052 30000 23108
rect 28960 23040 30000 23052
rect 0 22948 1040 22960
rect 0 22892 12 22948
rect 68 22892 332 22948
rect 388 22892 652 22948
rect 708 22892 972 22948
rect 1028 22892 1040 22948
rect 0 22880 1040 22892
rect 28960 22948 30000 22960
rect 28960 22892 28972 22948
rect 29028 22892 29292 22948
rect 29348 22892 29612 22948
rect 29668 22892 29932 22948
rect 29988 22892 30000 22948
rect 28960 22880 30000 22892
rect 0 22788 1040 22800
rect 0 22732 12 22788
rect 68 22732 332 22788
rect 388 22732 652 22788
rect 708 22732 972 22788
rect 1028 22732 1040 22788
rect 0 22720 1040 22732
rect 28960 22788 30000 22800
rect 28960 22732 28972 22788
rect 29028 22732 29292 22788
rect 29348 22732 29612 22788
rect 29668 22732 29932 22788
rect 29988 22732 30000 22788
rect 28960 22720 30000 22732
rect 28960 22628 30000 22640
rect 28960 22572 28972 22628
rect 29028 22572 29292 22628
rect 29348 22572 29612 22628
rect 29668 22572 29932 22628
rect 29988 22572 30000 22628
rect 28960 22560 30000 22572
rect 0 22468 1040 22480
rect 0 22412 12 22468
rect 68 22412 332 22468
rect 388 22412 652 22468
rect 708 22412 972 22468
rect 1028 22412 1040 22468
rect 0 22400 1040 22412
rect 28960 22468 30000 22480
rect 28960 22412 28972 22468
rect 29028 22412 29292 22468
rect 29348 22412 29612 22468
rect 29668 22412 29932 22468
rect 29988 22412 30000 22468
rect 28960 22400 30000 22412
rect 0 22308 400 22320
rect 0 22252 12 22308
rect 68 22252 332 22308
rect 388 22252 400 22308
rect 0 22240 400 22252
rect 28960 22308 30000 22320
rect 28960 22252 28972 22308
rect 29028 22252 29292 22308
rect 29348 22252 29612 22308
rect 29668 22252 29932 22308
rect 29988 22252 30000 22308
rect 28960 22240 30000 22252
rect 0 22148 1040 22160
rect 0 22092 12 22148
rect 68 22092 332 22148
rect 388 22092 652 22148
rect 708 22092 972 22148
rect 1028 22092 1040 22148
rect 0 22080 1040 22092
rect 28960 22148 30000 22160
rect 28960 22092 28972 22148
rect 29028 22092 29292 22148
rect 29348 22092 29612 22148
rect 29668 22092 29932 22148
rect 29988 22092 30000 22148
rect 28960 22080 30000 22092
rect 0 21988 1040 22000
rect 0 21932 12 21988
rect 68 21932 332 21988
rect 388 21932 652 21988
rect 708 21932 972 21988
rect 1028 21932 1040 21988
rect 0 21920 1040 21932
rect 28960 21988 30000 22000
rect 28960 21932 28972 21988
rect 29028 21932 29292 21988
rect 29348 21932 29612 21988
rect 29668 21932 29932 21988
rect 29988 21932 30000 21988
rect 28960 21920 30000 21932
rect 0 21828 1040 21840
rect 0 21772 12 21828
rect 68 21772 332 21828
rect 388 21772 652 21828
rect 708 21772 972 21828
rect 1028 21772 1040 21828
rect 0 21760 1040 21772
rect 28960 21828 30000 21840
rect 28960 21772 28972 21828
rect 29028 21772 29292 21828
rect 29348 21772 29612 21828
rect 29668 21772 29932 21828
rect 29988 21772 30000 21828
rect 28960 21760 30000 21772
rect 0 21668 1040 21680
rect 0 21612 12 21668
rect 68 21612 332 21668
rect 388 21612 652 21668
rect 708 21612 972 21668
rect 1028 21612 1040 21668
rect 0 21600 1040 21612
rect 28960 21668 30000 21680
rect 28960 21612 28972 21668
rect 29028 21612 29292 21668
rect 29348 21612 29612 21668
rect 29668 21612 29932 21668
rect 29988 21612 30000 21668
rect 28960 21600 30000 21612
rect 0 21508 1040 21520
rect 0 21452 12 21508
rect 68 21452 332 21508
rect 388 21452 652 21508
rect 708 21452 972 21508
rect 1028 21452 1040 21508
rect 0 21440 1040 21452
rect 28960 21508 30000 21520
rect 28960 21452 28972 21508
rect 29028 21452 29292 21508
rect 29348 21452 29612 21508
rect 29668 21452 29932 21508
rect 29988 21452 30000 21508
rect 28960 21440 30000 21452
rect 0 21348 1040 21360
rect 0 21292 12 21348
rect 68 21292 332 21348
rect 388 21292 652 21348
rect 708 21292 972 21348
rect 1028 21292 1040 21348
rect 0 21280 1040 21292
rect 28960 21348 30000 21360
rect 28960 21292 28972 21348
rect 29028 21292 29292 21348
rect 29348 21292 29612 21348
rect 29668 21292 29932 21348
rect 29988 21292 30000 21348
rect 28960 21280 30000 21292
rect 0 21188 1040 21200
rect 0 21132 12 21188
rect 68 21132 332 21188
rect 388 21132 652 21188
rect 708 21132 972 21188
rect 1028 21132 1040 21188
rect 0 21120 1040 21132
rect 28960 21188 30000 21200
rect 28960 21132 28972 21188
rect 29028 21132 29292 21188
rect 29348 21132 29612 21188
rect 29668 21132 29932 21188
rect 29988 21132 30000 21188
rect 28960 21120 30000 21132
rect 0 21028 1040 21040
rect 0 20972 12 21028
rect 68 20972 332 21028
rect 388 20972 652 21028
rect 708 20972 972 21028
rect 1028 20972 1040 21028
rect 0 20960 1040 20972
rect 28960 21028 30000 21040
rect 28960 20972 28972 21028
rect 29028 20972 29292 21028
rect 29348 20972 29612 21028
rect 29668 20972 29932 21028
rect 29988 20972 30000 21028
rect 28960 20960 30000 20972
rect 0 20868 1040 20880
rect 0 20812 12 20868
rect 68 20812 332 20868
rect 388 20812 652 20868
rect 708 20812 972 20868
rect 1028 20812 1040 20868
rect 0 20800 1040 20812
rect 28960 20868 30000 20880
rect 28960 20812 28972 20868
rect 29028 20812 29292 20868
rect 29348 20812 29612 20868
rect 29668 20812 29932 20868
rect 29988 20812 30000 20868
rect 28960 20800 30000 20812
rect 0 20708 1040 20720
rect 0 20652 12 20708
rect 68 20652 332 20708
rect 388 20652 652 20708
rect 708 20652 972 20708
rect 1028 20652 1040 20708
rect 0 20640 1040 20652
rect 28960 20708 30000 20720
rect 28960 20652 28972 20708
rect 29028 20652 29292 20708
rect 29348 20652 29612 20708
rect 29668 20652 29932 20708
rect 29988 20652 30000 20708
rect 28960 20640 30000 20652
rect 0 20548 1040 20560
rect 0 20492 12 20548
rect 68 20492 332 20548
rect 388 20492 652 20548
rect 708 20492 972 20548
rect 1028 20492 1040 20548
rect 0 20480 1040 20492
rect 28960 20548 30000 20560
rect 28960 20492 28972 20548
rect 29028 20492 29292 20548
rect 29348 20492 29612 20548
rect 29668 20492 29932 20548
rect 29988 20492 30000 20548
rect 28960 20480 30000 20492
rect 0 20388 1040 20400
rect 0 20332 12 20388
rect 68 20332 332 20388
rect 388 20332 652 20388
rect 708 20332 972 20388
rect 1028 20332 1040 20388
rect 0 20320 1040 20332
rect 28960 20388 30000 20400
rect 28960 20332 28972 20388
rect 29028 20332 29292 20388
rect 29348 20332 29612 20388
rect 29668 20332 29932 20388
rect 29988 20332 30000 20388
rect 28960 20320 30000 20332
rect 0 20228 1040 20240
rect 0 20172 12 20228
rect 68 20172 332 20228
rect 388 20172 652 20228
rect 708 20172 972 20228
rect 1028 20172 1040 20228
rect 0 20160 1040 20172
rect 28960 20228 30000 20240
rect 28960 20172 28972 20228
rect 29028 20172 29292 20228
rect 29348 20172 29612 20228
rect 29668 20172 29932 20228
rect 29988 20172 30000 20228
rect 28960 20160 30000 20172
rect 0 20068 1040 20080
rect 0 20012 12 20068
rect 68 20012 332 20068
rect 388 20012 652 20068
rect 708 20012 972 20068
rect 1028 20012 1040 20068
rect 0 20000 1040 20012
rect 28960 20068 30000 20080
rect 28960 20012 28972 20068
rect 29028 20012 29292 20068
rect 29348 20012 29612 20068
rect 29668 20012 29932 20068
rect 29988 20012 30000 20068
rect 28960 20000 30000 20012
rect 0 19908 1040 19920
rect 0 19852 12 19908
rect 68 19852 332 19908
rect 388 19852 652 19908
rect 708 19852 972 19908
rect 1028 19852 1040 19908
rect 0 19840 1040 19852
rect 28960 19908 30000 19920
rect 28960 19852 28972 19908
rect 29028 19852 29292 19908
rect 29348 19852 29612 19908
rect 29668 19852 29932 19908
rect 29988 19852 30000 19908
rect 28960 19840 30000 19852
rect 0 19748 720 19760
rect 0 19692 12 19748
rect 68 19692 332 19748
rect 388 19692 652 19748
rect 708 19692 720 19748
rect 0 19680 720 19692
rect 28960 19748 30000 19760
rect 28960 19692 28972 19748
rect 29028 19692 29292 19748
rect 29348 19692 29612 19748
rect 29668 19692 29932 19748
rect 29988 19692 30000 19748
rect 28960 19680 30000 19692
rect 0 19588 1040 19600
rect 0 19532 12 19588
rect 68 19532 332 19588
rect 388 19532 652 19588
rect 708 19532 972 19588
rect 1028 19532 1040 19588
rect 0 19520 1040 19532
rect 28960 19588 30000 19600
rect 28960 19532 28972 19588
rect 29028 19532 29292 19588
rect 29348 19532 29612 19588
rect 29668 19532 29932 19588
rect 29988 19532 30000 19588
rect 28960 19520 30000 19532
rect 0 19428 1040 19440
rect 0 19372 12 19428
rect 68 19372 332 19428
rect 388 19372 652 19428
rect 708 19372 972 19428
rect 1028 19372 1040 19428
rect 0 19360 1040 19372
rect 28960 19428 30000 19440
rect 28960 19372 28972 19428
rect 29028 19372 29292 19428
rect 29348 19372 29612 19428
rect 29668 19372 29932 19428
rect 29988 19372 30000 19428
rect 28960 19360 30000 19372
rect 0 19268 1040 19280
rect 0 19212 12 19268
rect 68 19212 332 19268
rect 388 19212 652 19268
rect 708 19212 972 19268
rect 1028 19212 1040 19268
rect 0 19200 1040 19212
rect 28960 19268 30000 19280
rect 28960 19212 28972 19268
rect 29028 19212 29292 19268
rect 29348 19212 29612 19268
rect 29668 19212 29932 19268
rect 29988 19212 30000 19268
rect 28960 19200 30000 19212
rect 0 19108 1040 19120
rect 0 19052 12 19108
rect 68 19052 332 19108
rect 388 19052 652 19108
rect 708 19052 972 19108
rect 1028 19052 1040 19108
rect 0 19040 1040 19052
rect 28960 19108 30000 19120
rect 28960 19052 28972 19108
rect 29028 19052 29292 19108
rect 29348 19052 29612 19108
rect 29668 19052 29932 19108
rect 29988 19052 30000 19108
rect 28960 19040 30000 19052
rect 0 18948 1040 18960
rect 0 18892 12 18948
rect 68 18892 332 18948
rect 388 18892 652 18948
rect 708 18892 972 18948
rect 1028 18892 1040 18948
rect 0 18880 1040 18892
rect 28960 18948 30000 18960
rect 28960 18892 28972 18948
rect 29028 18892 29292 18948
rect 29348 18892 29612 18948
rect 29668 18892 29932 18948
rect 29988 18892 30000 18948
rect 28960 18880 30000 18892
rect 0 18788 1040 18800
rect 0 18732 12 18788
rect 68 18732 332 18788
rect 388 18732 652 18788
rect 708 18732 972 18788
rect 1028 18732 1040 18788
rect 0 18720 1040 18732
rect 28960 18788 30000 18800
rect 28960 18732 28972 18788
rect 29028 18732 29292 18788
rect 29348 18732 29612 18788
rect 29668 18732 29932 18788
rect 29988 18732 30000 18788
rect 28960 18720 30000 18732
rect 0 18628 1040 18640
rect 0 18572 12 18628
rect 68 18572 332 18628
rect 388 18572 652 18628
rect 708 18572 972 18628
rect 1028 18572 1040 18628
rect 0 18560 1040 18572
rect 28960 18628 30000 18640
rect 28960 18572 28972 18628
rect 29028 18572 29292 18628
rect 29348 18572 29612 18628
rect 29668 18572 29932 18628
rect 29988 18572 30000 18628
rect 28960 18560 30000 18572
rect 0 18468 1040 18480
rect 0 18412 12 18468
rect 68 18412 332 18468
rect 388 18412 652 18468
rect 708 18412 972 18468
rect 1028 18412 1040 18468
rect 0 18400 1040 18412
rect 28960 18468 30000 18480
rect 28960 18412 28972 18468
rect 29028 18412 29292 18468
rect 29348 18412 29612 18468
rect 29668 18412 29932 18468
rect 29988 18412 30000 18468
rect 28960 18400 30000 18412
rect 0 18308 1040 18320
rect 0 18252 12 18308
rect 68 18252 332 18308
rect 388 18252 652 18308
rect 708 18252 972 18308
rect 1028 18252 1040 18308
rect 0 18240 1040 18252
rect 28960 18308 30000 18320
rect 28960 18252 28972 18308
rect 29028 18252 29292 18308
rect 29348 18252 29612 18308
rect 29668 18252 29932 18308
rect 29988 18252 30000 18308
rect 28960 18240 30000 18252
rect 0 18148 1040 18160
rect 0 18092 12 18148
rect 68 18092 332 18148
rect 388 18092 652 18148
rect 708 18092 972 18148
rect 1028 18092 1040 18148
rect 0 18080 1040 18092
rect 28960 18148 30000 18160
rect 28960 18092 28972 18148
rect 29028 18092 29292 18148
rect 29348 18092 29612 18148
rect 29668 18092 29932 18148
rect 29988 18092 30000 18148
rect 28960 18080 30000 18092
rect 0 17988 1040 18000
rect 0 17932 12 17988
rect 68 17932 332 17988
rect 388 17932 652 17988
rect 708 17932 972 17988
rect 1028 17932 1040 17988
rect 0 17920 1040 17932
rect 28960 17988 30000 18000
rect 28960 17932 28972 17988
rect 29028 17932 29292 17988
rect 29348 17932 29612 17988
rect 29668 17932 29932 17988
rect 29988 17932 30000 17988
rect 28960 17920 30000 17932
rect 0 17828 1040 17840
rect 0 17772 12 17828
rect 68 17772 332 17828
rect 388 17772 652 17828
rect 708 17772 972 17828
rect 1028 17772 1040 17828
rect 0 17760 1040 17772
rect 28960 17828 30000 17840
rect 28960 17772 28972 17828
rect 29028 17772 29292 17828
rect 29348 17772 29612 17828
rect 29668 17772 29932 17828
rect 29988 17772 30000 17828
rect 28960 17760 30000 17772
rect 0 17668 1040 17680
rect 0 17612 12 17668
rect 68 17612 332 17668
rect 388 17612 652 17668
rect 708 17612 972 17668
rect 1028 17612 1040 17668
rect 0 17600 1040 17612
rect 28960 17668 30000 17680
rect 28960 17612 28972 17668
rect 29028 17612 29292 17668
rect 29348 17612 29612 17668
rect 29668 17612 29932 17668
rect 29988 17612 30000 17668
rect 28960 17600 30000 17612
rect 0 17508 1040 17520
rect 0 17452 12 17508
rect 68 17452 332 17508
rect 388 17452 652 17508
rect 708 17452 972 17508
rect 1028 17452 1040 17508
rect 0 17440 1040 17452
rect 28960 17508 30000 17520
rect 28960 17452 28972 17508
rect 29028 17452 29292 17508
rect 29348 17452 29612 17508
rect 29668 17452 29932 17508
rect 29988 17452 30000 17508
rect 28960 17440 30000 17452
rect 0 17348 1040 17360
rect 0 17292 12 17348
rect 68 17292 332 17348
rect 388 17292 652 17348
rect 708 17292 972 17348
rect 1028 17292 1040 17348
rect 0 17280 1040 17292
rect 28960 17348 30000 17360
rect 28960 17292 28972 17348
rect 29028 17292 29292 17348
rect 29348 17292 29612 17348
rect 29668 17292 29932 17348
rect 29988 17292 30000 17348
rect 28960 17280 30000 17292
rect 0 17188 400 17200
rect 0 17132 12 17188
rect 68 17132 332 17188
rect 388 17132 400 17188
rect 0 17120 400 17132
rect 28960 17188 30000 17200
rect 28960 17132 28972 17188
rect 29028 17132 29292 17188
rect 29348 17132 29612 17188
rect 29668 17132 29932 17188
rect 29988 17132 30000 17188
rect 28960 17120 30000 17132
rect 0 17028 1040 17040
rect 0 16972 12 17028
rect 68 16972 332 17028
rect 388 16972 652 17028
rect 708 16972 972 17028
rect 1028 16972 1040 17028
rect 0 16960 1040 16972
rect 28960 17028 30000 17040
rect 28960 16972 28972 17028
rect 29028 16972 29292 17028
rect 29348 16972 29612 17028
rect 29668 16972 29932 17028
rect 29988 16972 30000 17028
rect 28960 16960 30000 16972
rect 28960 16868 30000 16880
rect 28960 16812 28972 16868
rect 29028 16812 29292 16868
rect 29348 16812 29612 16868
rect 29668 16812 29932 16868
rect 29988 16812 30000 16868
rect 28960 16800 30000 16812
rect 0 16708 1040 16720
rect 0 16652 12 16708
rect 68 16652 332 16708
rect 388 16652 652 16708
rect 708 16652 972 16708
rect 1028 16652 1040 16708
rect 0 16640 1040 16652
rect 28960 16708 30000 16720
rect 28960 16652 28972 16708
rect 29028 16652 29292 16708
rect 29348 16652 29612 16708
rect 29668 16652 29932 16708
rect 29988 16652 30000 16708
rect 28960 16640 30000 16652
rect 0 16548 1040 16560
rect 0 16492 12 16548
rect 68 16492 332 16548
rect 388 16492 652 16548
rect 708 16492 972 16548
rect 1028 16492 1040 16548
rect 0 16480 1040 16492
rect 28960 16548 30000 16560
rect 28960 16492 28972 16548
rect 29028 16492 29292 16548
rect 29348 16492 29612 16548
rect 29668 16492 29932 16548
rect 29988 16492 30000 16548
rect 28960 16480 30000 16492
rect 0 16388 1040 16400
rect 0 16332 12 16388
rect 68 16332 332 16388
rect 388 16332 652 16388
rect 708 16332 972 16388
rect 1028 16332 1040 16388
rect 0 16320 1040 16332
rect 28960 16388 30000 16400
rect 28960 16332 28972 16388
rect 29028 16332 29292 16388
rect 29348 16332 29612 16388
rect 29668 16332 29932 16388
rect 29988 16332 30000 16388
rect 28960 16320 30000 16332
rect 0 16228 1040 16240
rect 0 16172 12 16228
rect 68 16172 332 16228
rect 388 16172 652 16228
rect 708 16172 972 16228
rect 1028 16172 1040 16228
rect 0 16160 1040 16172
rect 28960 16228 30000 16240
rect 28960 16172 28972 16228
rect 29028 16172 29292 16228
rect 29348 16172 29612 16228
rect 29668 16172 29932 16228
rect 29988 16172 30000 16228
rect 28960 16160 30000 16172
rect 28960 16068 30000 16080
rect 28960 16012 28972 16068
rect 29028 16012 29292 16068
rect 29348 16012 29612 16068
rect 29668 16012 29932 16068
rect 29988 16012 30000 16068
rect 28960 16000 30000 16012
rect 0 15908 1040 15920
rect 0 15852 12 15908
rect 68 15852 332 15908
rect 388 15852 652 15908
rect 708 15852 972 15908
rect 1028 15852 1040 15908
rect 0 15840 1040 15852
rect 28960 15908 30000 15920
rect 28960 15852 28972 15908
rect 29028 15852 29292 15908
rect 29348 15852 29612 15908
rect 29668 15852 29932 15908
rect 29988 15852 30000 15908
rect 28960 15840 30000 15852
rect 0 15748 400 15760
rect 0 15692 12 15748
rect 68 15692 332 15748
rect 388 15692 400 15748
rect 0 15680 400 15692
rect 28960 15748 30000 15760
rect 28960 15692 28972 15748
rect 29028 15692 29292 15748
rect 29348 15692 29612 15748
rect 29668 15692 29932 15748
rect 29988 15692 30000 15748
rect 28960 15680 30000 15692
rect 0 15588 1040 15600
rect 0 15532 12 15588
rect 68 15532 332 15588
rect 388 15532 652 15588
rect 708 15532 972 15588
rect 1028 15532 1040 15588
rect 0 15520 1040 15532
rect 28960 15588 30000 15600
rect 28960 15532 28972 15588
rect 29028 15532 29292 15588
rect 29348 15532 29612 15588
rect 29668 15532 29932 15588
rect 29988 15532 30000 15588
rect 28960 15520 30000 15532
rect 0 15428 1040 15440
rect 0 15372 12 15428
rect 68 15372 332 15428
rect 388 15372 652 15428
rect 708 15372 972 15428
rect 1028 15372 1040 15428
rect 0 15360 1040 15372
rect 28960 15428 30000 15440
rect 28960 15372 28972 15428
rect 29028 15372 29292 15428
rect 29348 15372 29612 15428
rect 29668 15372 29932 15428
rect 29988 15372 30000 15428
rect 28960 15360 30000 15372
rect 0 15268 1040 15280
rect 0 15212 12 15268
rect 68 15212 332 15268
rect 388 15212 652 15268
rect 708 15212 972 15268
rect 1028 15212 1040 15268
rect 0 15200 1040 15212
rect 28960 15268 30000 15280
rect 28960 15212 28972 15268
rect 29028 15212 29292 15268
rect 29348 15212 29612 15268
rect 29668 15212 29932 15268
rect 29988 15212 30000 15268
rect 28960 15200 30000 15212
rect 0 15108 1040 15120
rect 0 15052 12 15108
rect 68 15052 332 15108
rect 388 15052 652 15108
rect 708 15052 972 15108
rect 1028 15052 1040 15108
rect 0 15040 1040 15052
rect 28960 15108 30000 15120
rect 28960 15052 28972 15108
rect 29028 15052 29292 15108
rect 29348 15052 29612 15108
rect 29668 15052 29932 15108
rect 29988 15052 30000 15108
rect 28960 15040 30000 15052
rect 0 14948 1040 14960
rect 0 14892 12 14948
rect 68 14892 332 14948
rect 388 14892 652 14948
rect 708 14892 972 14948
rect 1028 14892 1040 14948
rect 0 14880 1040 14892
rect 28960 14948 30000 14960
rect 28960 14892 28972 14948
rect 29028 14892 29292 14948
rect 29348 14892 29612 14948
rect 29668 14892 29932 14948
rect 29988 14892 30000 14948
rect 28960 14880 30000 14892
rect 0 14788 1040 14800
rect 0 14732 12 14788
rect 68 14732 332 14788
rect 388 14732 652 14788
rect 708 14732 972 14788
rect 1028 14732 1040 14788
rect 0 14720 1040 14732
rect 28960 14788 30000 14800
rect 28960 14732 28972 14788
rect 29028 14732 29292 14788
rect 29348 14732 29612 14788
rect 29668 14732 29932 14788
rect 29988 14732 30000 14788
rect 28960 14720 30000 14732
rect 0 14628 1040 14640
rect 0 14572 12 14628
rect 68 14572 332 14628
rect 388 14572 652 14628
rect 708 14572 972 14628
rect 1028 14572 1040 14628
rect 0 14560 1040 14572
rect 28960 14628 30000 14640
rect 28960 14572 28972 14628
rect 29028 14572 29292 14628
rect 29348 14572 29612 14628
rect 29668 14572 29932 14628
rect 29988 14572 30000 14628
rect 28960 14560 30000 14572
rect 0 14468 1040 14480
rect 0 14412 12 14468
rect 68 14412 332 14468
rect 388 14412 652 14468
rect 708 14412 972 14468
rect 1028 14412 1040 14468
rect 0 14400 1040 14412
rect 28960 14468 30000 14480
rect 28960 14412 28972 14468
rect 29028 14412 29292 14468
rect 29348 14412 29612 14468
rect 29668 14412 29932 14468
rect 29988 14412 30000 14468
rect 28960 14400 30000 14412
rect 0 14308 1040 14320
rect 0 14252 12 14308
rect 68 14252 332 14308
rect 388 14252 652 14308
rect 708 14252 972 14308
rect 1028 14252 1040 14308
rect 0 14240 1040 14252
rect 28960 14308 30000 14320
rect 28960 14252 28972 14308
rect 29028 14252 29292 14308
rect 29348 14252 29612 14308
rect 29668 14252 29932 14308
rect 29988 14252 30000 14308
rect 28960 14240 30000 14252
rect 0 14148 1040 14160
rect 0 14092 12 14148
rect 68 14092 332 14148
rect 388 14092 652 14148
rect 708 14092 972 14148
rect 1028 14092 1040 14148
rect 0 14080 1040 14092
rect 28960 14148 30000 14160
rect 28960 14092 28972 14148
rect 29028 14092 29292 14148
rect 29348 14092 29612 14148
rect 29668 14092 29932 14148
rect 29988 14092 30000 14148
rect 28960 14080 30000 14092
rect 0 13988 1040 14000
rect 0 13932 12 13988
rect 68 13932 332 13988
rect 388 13932 652 13988
rect 708 13932 972 13988
rect 1028 13932 1040 13988
rect 0 13920 1040 13932
rect 28960 13988 30000 14000
rect 28960 13932 28972 13988
rect 29028 13932 29292 13988
rect 29348 13932 29612 13988
rect 29668 13932 29932 13988
rect 29988 13932 30000 13988
rect 28960 13920 30000 13932
rect 0 13828 1040 13840
rect 0 13772 12 13828
rect 68 13772 332 13828
rect 388 13772 652 13828
rect 708 13772 972 13828
rect 1028 13772 1040 13828
rect 0 13760 1040 13772
rect 28960 13828 30000 13840
rect 28960 13772 28972 13828
rect 29028 13772 29292 13828
rect 29348 13772 29612 13828
rect 29668 13772 29932 13828
rect 29988 13772 30000 13828
rect 28960 13760 30000 13772
rect 0 13668 1040 13680
rect 0 13612 12 13668
rect 68 13612 332 13668
rect 388 13612 652 13668
rect 708 13612 972 13668
rect 1028 13612 1040 13668
rect 0 13600 1040 13612
rect 28960 13668 30000 13680
rect 28960 13612 28972 13668
rect 29028 13612 29292 13668
rect 29348 13612 29612 13668
rect 29668 13612 29932 13668
rect 29988 13612 30000 13668
rect 28960 13600 30000 13612
rect 0 13508 1040 13520
rect 0 13452 12 13508
rect 68 13452 332 13508
rect 388 13452 652 13508
rect 708 13452 972 13508
rect 1028 13452 1040 13508
rect 0 13440 1040 13452
rect 28960 13508 30000 13520
rect 28960 13452 28972 13508
rect 29028 13452 29292 13508
rect 29348 13452 29612 13508
rect 29668 13452 29932 13508
rect 29988 13452 30000 13508
rect 28960 13440 30000 13452
rect 0 13348 1040 13360
rect 0 13292 12 13348
rect 68 13292 332 13348
rect 388 13292 652 13348
rect 708 13292 972 13348
rect 1028 13292 1040 13348
rect 0 13280 1040 13292
rect 28960 13348 30000 13360
rect 28960 13292 28972 13348
rect 29028 13292 29292 13348
rect 29348 13292 29612 13348
rect 29668 13292 29932 13348
rect 29988 13292 30000 13348
rect 28960 13280 30000 13292
rect 0 13188 720 13200
rect 0 13132 12 13188
rect 68 13132 332 13188
rect 388 13132 652 13188
rect 708 13132 720 13188
rect 0 13120 720 13132
rect 28960 13188 30000 13200
rect 28960 13132 28972 13188
rect 29028 13132 29292 13188
rect 29348 13132 29612 13188
rect 29668 13132 29932 13188
rect 29988 13132 30000 13188
rect 28960 13120 30000 13132
rect 0 13028 1040 13040
rect 0 12972 12 13028
rect 68 12972 332 13028
rect 388 12972 652 13028
rect 708 12972 972 13028
rect 1028 12972 1040 13028
rect 0 12960 1040 12972
rect 28960 13028 30000 13040
rect 28960 12972 28972 13028
rect 29028 12972 29292 13028
rect 29348 12972 29612 13028
rect 29668 12972 29932 13028
rect 29988 12972 30000 13028
rect 28960 12960 30000 12972
rect 0 12868 1040 12880
rect 0 12812 12 12868
rect 68 12812 332 12868
rect 388 12812 652 12868
rect 708 12812 972 12868
rect 1028 12812 1040 12868
rect 0 12800 1040 12812
rect 28960 12868 30000 12880
rect 28960 12812 28972 12868
rect 29028 12812 29292 12868
rect 29348 12812 29612 12868
rect 29668 12812 29932 12868
rect 29988 12812 30000 12868
rect 28960 12800 30000 12812
rect 0 12708 1040 12720
rect 0 12652 12 12708
rect 68 12652 332 12708
rect 388 12652 652 12708
rect 708 12652 972 12708
rect 1028 12652 1040 12708
rect 0 12640 1040 12652
rect 28960 12708 30000 12720
rect 28960 12652 28972 12708
rect 29028 12652 29292 12708
rect 29348 12652 29612 12708
rect 29668 12652 29932 12708
rect 29988 12652 30000 12708
rect 28960 12640 30000 12652
rect 0 12548 1040 12560
rect 0 12492 12 12548
rect 68 12492 332 12548
rect 388 12492 652 12548
rect 708 12492 972 12548
rect 1028 12492 1040 12548
rect 0 12480 1040 12492
rect 28960 12548 30000 12560
rect 28960 12492 28972 12548
rect 29028 12492 29292 12548
rect 29348 12492 29612 12548
rect 29668 12492 29932 12548
rect 29988 12492 30000 12548
rect 28960 12480 30000 12492
rect 0 12388 1040 12400
rect 0 12332 12 12388
rect 68 12332 332 12388
rect 388 12332 652 12388
rect 708 12332 972 12388
rect 1028 12332 1040 12388
rect 0 12320 1040 12332
rect 28960 12388 30000 12400
rect 28960 12332 28972 12388
rect 29028 12332 29292 12388
rect 29348 12332 29612 12388
rect 29668 12332 29932 12388
rect 29988 12332 30000 12388
rect 28960 12320 30000 12332
rect 0 12228 1040 12240
rect 0 12172 12 12228
rect 68 12172 332 12228
rect 388 12172 652 12228
rect 708 12172 972 12228
rect 1028 12172 1040 12228
rect 0 12160 1040 12172
rect 28960 12228 30000 12240
rect 28960 12172 28972 12228
rect 29028 12172 29292 12228
rect 29348 12172 29612 12228
rect 29668 12172 29932 12228
rect 29988 12172 30000 12228
rect 28960 12160 30000 12172
rect 0 12068 1040 12080
rect 0 12012 12 12068
rect 68 12012 332 12068
rect 388 12012 652 12068
rect 708 12012 972 12068
rect 1028 12012 1040 12068
rect 0 12000 1040 12012
rect 28960 12068 30000 12080
rect 28960 12012 28972 12068
rect 29028 12012 29292 12068
rect 29348 12012 29612 12068
rect 29668 12012 29932 12068
rect 29988 12012 30000 12068
rect 28960 12000 30000 12012
rect 0 11908 1040 11920
rect 0 11852 12 11908
rect 68 11852 332 11908
rect 388 11852 652 11908
rect 708 11852 972 11908
rect 1028 11852 1040 11908
rect 0 11840 1040 11852
rect 28960 11908 30000 11920
rect 28960 11852 28972 11908
rect 29028 11852 29292 11908
rect 29348 11852 29612 11908
rect 29668 11852 29932 11908
rect 29988 11852 30000 11908
rect 28960 11840 30000 11852
rect 0 11748 1040 11760
rect 0 11692 12 11748
rect 68 11692 332 11748
rect 388 11692 652 11748
rect 708 11692 972 11748
rect 1028 11692 1040 11748
rect 0 11680 1040 11692
rect 28960 11748 30000 11760
rect 28960 11692 28972 11748
rect 29028 11692 29292 11748
rect 29348 11692 29612 11748
rect 29668 11692 29932 11748
rect 29988 11692 30000 11748
rect 28960 11680 30000 11692
rect 0 11588 1040 11600
rect 0 11532 12 11588
rect 68 11532 332 11588
rect 388 11532 652 11588
rect 708 11532 972 11588
rect 1028 11532 1040 11588
rect 0 11520 1040 11532
rect 28960 11588 30000 11600
rect 28960 11532 28972 11588
rect 29028 11532 29292 11588
rect 29348 11532 29612 11588
rect 29668 11532 29932 11588
rect 29988 11532 30000 11588
rect 28960 11520 30000 11532
rect 0 11428 1040 11440
rect 0 11372 12 11428
rect 68 11372 332 11428
rect 388 11372 652 11428
rect 708 11372 972 11428
rect 1028 11372 1040 11428
rect 0 11360 1040 11372
rect 28960 11428 30000 11440
rect 28960 11372 28972 11428
rect 29028 11372 29292 11428
rect 29348 11372 29612 11428
rect 29668 11372 29932 11428
rect 29988 11372 30000 11428
rect 28960 11360 30000 11372
rect 0 11268 1040 11280
rect 0 11212 12 11268
rect 68 11212 332 11268
rect 388 11212 652 11268
rect 708 11212 972 11268
rect 1028 11212 1040 11268
rect 0 11200 1040 11212
rect 28960 11268 30000 11280
rect 28960 11212 28972 11268
rect 29028 11212 29292 11268
rect 29348 11212 29612 11268
rect 29668 11212 29932 11268
rect 29988 11212 30000 11268
rect 28960 11200 30000 11212
rect 0 11108 1040 11120
rect 0 11052 12 11108
rect 68 11052 332 11108
rect 388 11052 652 11108
rect 708 11052 972 11108
rect 1028 11052 1040 11108
rect 0 11040 1040 11052
rect 28960 11108 30000 11120
rect 28960 11052 28972 11108
rect 29028 11052 29292 11108
rect 29348 11052 29612 11108
rect 29668 11052 29932 11108
rect 29988 11052 30000 11108
rect 28960 11040 30000 11052
rect 0 10948 1040 10960
rect 0 10892 12 10948
rect 68 10892 332 10948
rect 388 10892 652 10948
rect 708 10892 972 10948
rect 1028 10892 1040 10948
rect 0 10880 1040 10892
rect 28960 10948 30000 10960
rect 28960 10892 28972 10948
rect 29028 10892 29292 10948
rect 29348 10892 29612 10948
rect 29668 10892 29932 10948
rect 29988 10892 30000 10948
rect 28960 10880 30000 10892
rect 0 10788 1040 10800
rect 0 10732 12 10788
rect 68 10732 332 10788
rect 388 10732 652 10788
rect 708 10732 972 10788
rect 1028 10732 1040 10788
rect 0 10720 1040 10732
rect 28960 10788 30000 10800
rect 28960 10732 28972 10788
rect 29028 10732 29292 10788
rect 29348 10732 29612 10788
rect 29668 10732 29932 10788
rect 29988 10732 30000 10788
rect 28960 10720 30000 10732
rect 0 10628 400 10640
rect 0 10572 12 10628
rect 68 10572 332 10628
rect 388 10572 400 10628
rect 0 10560 400 10572
rect 28960 10628 30000 10640
rect 28960 10572 28972 10628
rect 29028 10572 29292 10628
rect 29348 10572 29612 10628
rect 29668 10572 29932 10628
rect 29988 10572 30000 10628
rect 28960 10560 30000 10572
rect 0 10468 1040 10480
rect 0 10412 12 10468
rect 68 10412 332 10468
rect 388 10412 652 10468
rect 708 10412 972 10468
rect 1028 10412 1040 10468
rect 0 10400 1040 10412
rect 28960 10468 30000 10480
rect 28960 10412 28972 10468
rect 29028 10412 29292 10468
rect 29348 10412 29612 10468
rect 29668 10412 29932 10468
rect 29988 10412 30000 10468
rect 28960 10400 30000 10412
rect 28960 10308 30000 10320
rect 28960 10252 28972 10308
rect 29028 10252 29292 10308
rect 29348 10252 29612 10308
rect 29668 10252 29932 10308
rect 29988 10252 30000 10308
rect 28960 10240 30000 10252
rect 0 10148 1040 10160
rect 0 10092 12 10148
rect 68 10092 332 10148
rect 388 10092 652 10148
rect 708 10092 972 10148
rect 1028 10092 1040 10148
rect 0 10080 1040 10092
rect 28960 10148 30000 10160
rect 28960 10092 28972 10148
rect 29028 10092 29292 10148
rect 29348 10092 29612 10148
rect 29668 10092 29932 10148
rect 29988 10092 30000 10148
rect 28960 10080 30000 10092
rect 0 9988 1040 10000
rect 0 9932 12 9988
rect 68 9932 332 9988
rect 388 9932 652 9988
rect 708 9932 972 9988
rect 1028 9932 1040 9988
rect 0 9920 1040 9932
rect 28960 9988 30000 10000
rect 28960 9932 28972 9988
rect 29028 9932 29292 9988
rect 29348 9932 29612 9988
rect 29668 9932 29932 9988
rect 29988 9932 30000 9988
rect 28960 9920 30000 9932
rect 0 9828 1040 9840
rect 0 9772 12 9828
rect 68 9772 332 9828
rect 388 9772 652 9828
rect 708 9772 972 9828
rect 1028 9772 1040 9828
rect 0 9760 1040 9772
rect 28960 9828 30000 9840
rect 28960 9772 28972 9828
rect 29028 9772 29292 9828
rect 29348 9772 29612 9828
rect 29668 9772 29932 9828
rect 29988 9772 30000 9828
rect 28960 9760 30000 9772
rect 0 9668 1040 9680
rect 0 9612 12 9668
rect 68 9612 332 9668
rect 388 9612 652 9668
rect 708 9612 972 9668
rect 1028 9612 1040 9668
rect 0 9600 1040 9612
rect 28960 9668 30000 9680
rect 28960 9612 28972 9668
rect 29028 9612 29292 9668
rect 29348 9612 29612 9668
rect 29668 9612 29932 9668
rect 29988 9612 30000 9668
rect 28960 9600 30000 9612
rect 0 9508 1040 9520
rect 0 9452 12 9508
rect 68 9452 332 9508
rect 388 9452 652 9508
rect 708 9452 972 9508
rect 1028 9452 1040 9508
rect 0 9440 1040 9452
rect 0 9348 1040 9360
rect 0 9292 12 9348
rect 68 9292 332 9348
rect 388 9292 652 9348
rect 708 9292 972 9348
rect 1028 9292 1040 9348
rect 0 9280 1040 9292
rect 28960 9348 30000 9360
rect 28960 9292 28972 9348
rect 29028 9292 29292 9348
rect 29348 9292 29612 9348
rect 29668 9292 29932 9348
rect 29988 9292 30000 9348
rect 28960 9280 30000 9292
rect 0 9188 1040 9200
rect 0 9132 12 9188
rect 68 9132 332 9188
rect 388 9132 652 9188
rect 708 9132 972 9188
rect 1028 9132 1040 9188
rect 0 9120 1040 9132
rect 29600 9188 30000 9200
rect 29600 9132 29612 9188
rect 29668 9132 29932 9188
rect 29988 9132 30000 9188
rect 29600 9120 30000 9132
rect 0 9028 1040 9040
rect 0 8972 12 9028
rect 68 8972 332 9028
rect 388 8972 652 9028
rect 708 8972 972 9028
rect 1028 8972 1040 9028
rect 0 8960 1040 8972
rect 28960 9028 30000 9040
rect 28960 8972 28972 9028
rect 29028 8972 29292 9028
rect 29348 8972 29612 9028
rect 29668 8972 29932 9028
rect 29988 8972 30000 9028
rect 28960 8960 30000 8972
rect 0 8868 1040 8880
rect 0 8812 12 8868
rect 68 8812 332 8868
rect 388 8812 652 8868
rect 708 8812 972 8868
rect 1028 8812 1040 8868
rect 0 8800 1040 8812
rect 28960 8868 30000 8880
rect 28960 8812 28972 8868
rect 29028 8812 29292 8868
rect 29348 8812 29612 8868
rect 29668 8812 29932 8868
rect 29988 8812 30000 8868
rect 28960 8800 30000 8812
rect 0 8708 1040 8720
rect 0 8652 12 8708
rect 68 8652 332 8708
rect 388 8652 652 8708
rect 708 8652 972 8708
rect 1028 8652 1040 8708
rect 0 8640 1040 8652
rect 28960 8708 30000 8720
rect 28960 8652 28972 8708
rect 29028 8652 29292 8708
rect 29348 8652 29612 8708
rect 29668 8652 29932 8708
rect 29988 8652 30000 8708
rect 28960 8640 30000 8652
rect 0 8548 1040 8560
rect 0 8492 12 8548
rect 68 8492 332 8548
rect 388 8492 652 8548
rect 708 8492 972 8548
rect 1028 8492 1040 8548
rect 0 8480 1040 8492
rect 28960 8548 30000 8560
rect 28960 8492 28972 8548
rect 29028 8492 29292 8548
rect 29348 8492 29612 8548
rect 29668 8492 29932 8548
rect 29988 8492 30000 8548
rect 28960 8480 30000 8492
rect 0 8388 1040 8400
rect 0 8332 12 8388
rect 68 8332 332 8388
rect 388 8332 652 8388
rect 708 8332 972 8388
rect 1028 8332 1040 8388
rect 0 8320 1040 8332
rect 28960 8388 30000 8400
rect 28960 8332 28972 8388
rect 29028 8332 29292 8388
rect 29348 8332 29612 8388
rect 29668 8332 29932 8388
rect 29988 8332 30000 8388
rect 28960 8320 30000 8332
rect 0 8228 1040 8240
rect 0 8172 12 8228
rect 68 8172 332 8228
rect 388 8172 652 8228
rect 708 8172 972 8228
rect 1028 8172 1040 8228
rect 0 8160 1040 8172
rect 28960 8228 30000 8240
rect 28960 8172 28972 8228
rect 29028 8172 29292 8228
rect 29348 8172 29612 8228
rect 29668 8172 29932 8228
rect 29988 8172 30000 8228
rect 28960 8160 30000 8172
rect 0 8068 1040 8080
rect 0 8012 12 8068
rect 68 8012 332 8068
rect 388 8012 652 8068
rect 708 8012 972 8068
rect 1028 8012 1040 8068
rect 0 8000 1040 8012
rect 28960 8068 30000 8080
rect 28960 8012 28972 8068
rect 29028 8012 29292 8068
rect 29348 8012 29612 8068
rect 29668 8012 29932 8068
rect 29988 8012 30000 8068
rect 28960 8000 30000 8012
rect 0 7908 1040 7920
rect 0 7852 12 7908
rect 68 7852 332 7908
rect 388 7852 652 7908
rect 708 7852 972 7908
rect 1028 7852 1040 7908
rect 0 7840 1040 7852
rect 28960 7908 30000 7920
rect 28960 7852 28972 7908
rect 29028 7852 29292 7908
rect 29348 7852 29612 7908
rect 29668 7852 29932 7908
rect 29988 7852 30000 7908
rect 28960 7840 30000 7852
rect 0 7748 1040 7760
rect 0 7692 12 7748
rect 68 7692 332 7748
rect 388 7692 652 7748
rect 708 7692 972 7748
rect 1028 7692 1040 7748
rect 0 7680 1040 7692
rect 28960 7748 30000 7760
rect 28960 7692 28972 7748
rect 29028 7692 29292 7748
rect 29348 7692 29612 7748
rect 29668 7692 29932 7748
rect 29988 7692 30000 7748
rect 28960 7680 30000 7692
rect 0 7588 1040 7600
rect 0 7532 12 7588
rect 68 7532 332 7588
rect 388 7532 652 7588
rect 708 7532 972 7588
rect 1028 7532 1040 7588
rect 0 7520 1040 7532
rect 28960 7588 30000 7600
rect 28960 7532 28972 7588
rect 29028 7532 29292 7588
rect 29348 7532 29612 7588
rect 29668 7532 29932 7588
rect 29988 7532 30000 7588
rect 28960 7520 30000 7532
rect 0 7428 1040 7440
rect 0 7372 12 7428
rect 68 7372 332 7428
rect 388 7372 652 7428
rect 708 7372 972 7428
rect 1028 7372 1040 7428
rect 0 7360 1040 7372
rect 28960 7428 30000 7440
rect 28960 7372 28972 7428
rect 29028 7372 29292 7428
rect 29348 7372 29612 7428
rect 29668 7372 29932 7428
rect 29988 7372 30000 7428
rect 28960 7360 30000 7372
rect 0 7268 1040 7280
rect 0 7212 12 7268
rect 68 7212 332 7268
rect 388 7212 652 7268
rect 708 7212 972 7268
rect 1028 7212 1040 7268
rect 0 7200 1040 7212
rect 28960 7268 30000 7280
rect 28960 7212 28972 7268
rect 29028 7212 29292 7268
rect 29348 7212 29612 7268
rect 29668 7212 29932 7268
rect 29988 7212 30000 7268
rect 28960 7200 30000 7212
rect 0 7108 1040 7120
rect 0 7052 12 7108
rect 68 7052 332 7108
rect 388 7052 652 7108
rect 708 7052 972 7108
rect 1028 7052 1040 7108
rect 0 7040 1040 7052
rect 28960 7108 30000 7120
rect 28960 7052 28972 7108
rect 29028 7052 29292 7108
rect 29348 7052 29612 7108
rect 29668 7052 29932 7108
rect 29988 7052 30000 7108
rect 28960 7040 30000 7052
rect 0 6948 1040 6960
rect 0 6892 12 6948
rect 68 6892 332 6948
rect 388 6892 652 6948
rect 708 6892 972 6948
rect 1028 6892 1040 6948
rect 0 6880 1040 6892
rect 28960 6948 30000 6960
rect 28960 6892 28972 6948
rect 29028 6892 29292 6948
rect 29348 6892 29612 6948
rect 29668 6892 29932 6948
rect 29988 6892 30000 6948
rect 28960 6880 30000 6892
rect 0 6788 1040 6800
rect 0 6732 12 6788
rect 68 6732 332 6788
rect 388 6732 652 6788
rect 708 6732 972 6788
rect 1028 6732 1040 6788
rect 0 6720 1040 6732
rect 28960 6788 30000 6800
rect 28960 6732 28972 6788
rect 29028 6732 29292 6788
rect 29348 6732 29612 6788
rect 29668 6732 29932 6788
rect 29988 6732 30000 6788
rect 28960 6720 30000 6732
rect 0 6628 1040 6640
rect 0 6572 12 6628
rect 68 6572 332 6628
rect 388 6572 652 6628
rect 708 6572 972 6628
rect 1028 6572 1040 6628
rect 0 6560 1040 6572
rect 29280 6628 30000 6640
rect 29280 6572 29292 6628
rect 29348 6572 29612 6628
rect 29668 6572 29932 6628
rect 29988 6572 30000 6628
rect 29280 6560 30000 6572
rect 0 6468 1040 6480
rect 0 6412 12 6468
rect 68 6412 332 6468
rect 388 6412 652 6468
rect 708 6412 972 6468
rect 1028 6412 1040 6468
rect 0 6400 1040 6412
rect 28960 6468 30000 6480
rect 28960 6412 28972 6468
rect 29028 6412 29292 6468
rect 29348 6412 29612 6468
rect 29668 6412 29932 6468
rect 29988 6412 30000 6468
rect 28960 6400 30000 6412
rect 0 6308 1040 6320
rect 0 6252 12 6308
rect 68 6252 332 6308
rect 388 6252 652 6308
rect 708 6252 972 6308
rect 1028 6252 1040 6308
rect 0 6240 1040 6252
rect 28960 6308 30000 6320
rect 28960 6252 28972 6308
rect 29028 6252 29292 6308
rect 29348 6252 29612 6308
rect 29668 6252 29932 6308
rect 29988 6252 30000 6308
rect 28960 6240 30000 6252
rect 0 6148 1040 6160
rect 0 6092 12 6148
rect 68 6092 332 6148
rect 388 6092 652 6148
rect 708 6092 972 6148
rect 1028 6092 1040 6148
rect 0 6080 1040 6092
rect 28960 6148 30000 6160
rect 28960 6092 28972 6148
rect 29028 6092 29292 6148
rect 29348 6092 29612 6148
rect 29668 6092 29932 6148
rect 29988 6092 30000 6148
rect 28960 6080 30000 6092
rect 0 5988 1040 6000
rect 0 5932 12 5988
rect 68 5932 332 5988
rect 388 5932 652 5988
rect 708 5932 972 5988
rect 1028 5932 1040 5988
rect 0 5920 1040 5932
rect 28960 5988 30000 6000
rect 28960 5932 28972 5988
rect 29028 5932 29292 5988
rect 29348 5932 29612 5988
rect 29668 5932 29932 5988
rect 29988 5932 30000 5988
rect 28960 5920 30000 5932
rect 0 5828 1040 5840
rect 0 5772 12 5828
rect 68 5772 332 5828
rect 388 5772 652 5828
rect 708 5772 972 5828
rect 1028 5772 1040 5828
rect 0 5760 1040 5772
rect 28960 5828 30000 5840
rect 28960 5772 28972 5828
rect 29028 5772 29292 5828
rect 29348 5772 29612 5828
rect 29668 5772 29932 5828
rect 29988 5772 30000 5828
rect 28960 5760 30000 5772
rect 0 5668 1040 5680
rect 0 5612 12 5668
rect 68 5612 332 5668
rect 388 5612 652 5668
rect 708 5612 972 5668
rect 1028 5612 1040 5668
rect 0 5600 1040 5612
rect 28960 5668 30000 5680
rect 28960 5612 28972 5668
rect 29028 5612 29292 5668
rect 29348 5612 29612 5668
rect 29668 5612 29932 5668
rect 29988 5612 30000 5668
rect 28960 5600 30000 5612
rect 0 5508 1040 5520
rect 0 5452 12 5508
rect 68 5452 332 5508
rect 388 5452 652 5508
rect 708 5452 972 5508
rect 1028 5452 1040 5508
rect 0 5440 1040 5452
rect 28960 5508 30000 5520
rect 28960 5452 28972 5508
rect 29028 5452 29292 5508
rect 29348 5452 29612 5508
rect 29668 5452 29932 5508
rect 29988 5452 30000 5508
rect 28960 5440 30000 5452
rect 0 5348 1040 5360
rect 0 5292 12 5348
rect 68 5292 332 5348
rect 388 5292 652 5348
rect 708 5292 972 5348
rect 1028 5292 1040 5348
rect 0 5280 1040 5292
rect 28960 5348 30000 5360
rect 28960 5292 28972 5348
rect 29028 5292 29292 5348
rect 29348 5292 29612 5348
rect 29668 5292 29932 5348
rect 29988 5292 30000 5348
rect 28960 5280 30000 5292
rect 0 5188 1040 5200
rect 0 5132 12 5188
rect 68 5132 332 5188
rect 388 5132 652 5188
rect 708 5132 972 5188
rect 1028 5132 1040 5188
rect 0 5120 1040 5132
rect 28960 5188 30000 5200
rect 28960 5132 28972 5188
rect 29028 5132 29292 5188
rect 29348 5132 29612 5188
rect 29668 5132 29932 5188
rect 29988 5132 30000 5188
rect 28960 5120 30000 5132
rect 0 5028 1040 5040
rect 0 4972 12 5028
rect 68 4972 332 5028
rect 388 4972 652 5028
rect 708 4972 972 5028
rect 1028 4972 1040 5028
rect 0 4960 1040 4972
rect 28960 5028 30000 5040
rect 28960 4972 28972 5028
rect 29028 4972 29292 5028
rect 29348 4972 29612 5028
rect 29668 4972 29932 5028
rect 29988 4972 30000 5028
rect 28960 4960 30000 4972
rect 0 4868 1040 4880
rect 0 4812 12 4868
rect 68 4812 332 4868
rect 388 4812 652 4868
rect 708 4812 972 4868
rect 1028 4812 1040 4868
rect 0 4800 1040 4812
rect 28960 4868 30000 4880
rect 28960 4812 28972 4868
rect 29028 4812 29292 4868
rect 29348 4812 29612 4868
rect 29668 4812 29932 4868
rect 29988 4812 30000 4868
rect 28960 4800 30000 4812
rect 0 4708 1040 4720
rect 0 4652 12 4708
rect 68 4652 332 4708
rect 388 4652 652 4708
rect 708 4652 972 4708
rect 1028 4652 1040 4708
rect 0 4640 1040 4652
rect 28960 4708 30000 4720
rect 28960 4652 28972 4708
rect 29028 4652 29292 4708
rect 29348 4652 29612 4708
rect 29668 4652 29932 4708
rect 29988 4652 30000 4708
rect 28960 4640 30000 4652
rect 0 4548 1040 4560
rect 0 4492 12 4548
rect 68 4492 332 4548
rect 388 4492 652 4548
rect 708 4492 972 4548
rect 1028 4492 1040 4548
rect 0 4480 1040 4492
rect 28960 4548 30000 4560
rect 28960 4492 28972 4548
rect 29028 4492 29292 4548
rect 29348 4492 29612 4548
rect 29668 4492 29932 4548
rect 29988 4492 30000 4548
rect 28960 4480 30000 4492
rect 0 4388 1040 4400
rect 0 4332 12 4388
rect 68 4332 332 4388
rect 388 4332 652 4388
rect 708 4332 972 4388
rect 1028 4332 1040 4388
rect 0 4320 1040 4332
rect 28960 4388 30000 4400
rect 28960 4332 28972 4388
rect 29028 4332 29292 4388
rect 29348 4332 29612 4388
rect 29668 4332 29932 4388
rect 29988 4332 30000 4388
rect 28960 4320 30000 4332
rect 0 4228 1040 4240
rect 0 4172 12 4228
rect 68 4172 332 4228
rect 388 4172 652 4228
rect 708 4172 972 4228
rect 1028 4172 1040 4228
rect 0 4160 1040 4172
rect 28960 4228 30000 4240
rect 28960 4172 28972 4228
rect 29028 4172 29292 4228
rect 29348 4172 29612 4228
rect 29668 4172 29932 4228
rect 29988 4172 30000 4228
rect 28960 4160 30000 4172
rect 0 4068 1040 4080
rect 0 4012 12 4068
rect 68 4012 332 4068
rect 388 4012 652 4068
rect 708 4012 972 4068
rect 1028 4012 1040 4068
rect 0 4000 1040 4012
rect 29600 4068 30000 4080
rect 29600 4012 29612 4068
rect 29668 4012 29932 4068
rect 29988 4012 30000 4068
rect 29600 4000 30000 4012
rect 0 3908 1040 3920
rect 0 3852 12 3908
rect 68 3852 332 3908
rect 388 3852 652 3908
rect 708 3852 972 3908
rect 1028 3852 1040 3908
rect 0 3840 1040 3852
rect 28960 3908 30000 3920
rect 28960 3852 28972 3908
rect 29028 3852 29292 3908
rect 29348 3852 29612 3908
rect 29668 3852 29932 3908
rect 29988 3852 30000 3908
rect 28960 3840 30000 3852
rect 0 3748 1040 3760
rect 0 3692 12 3748
rect 68 3692 332 3748
rect 388 3692 652 3748
rect 708 3692 972 3748
rect 1028 3692 1040 3748
rect 0 3680 1040 3692
rect 0 3588 1040 3600
rect 0 3532 12 3588
rect 68 3532 332 3588
rect 388 3532 652 3588
rect 708 3532 972 3588
rect 1028 3532 1040 3588
rect 0 3520 1040 3532
rect 28960 3588 30000 3600
rect 28960 3532 28972 3588
rect 29028 3532 29292 3588
rect 29348 3532 29612 3588
rect 29668 3532 29932 3588
rect 29988 3532 30000 3588
rect 28960 3520 30000 3532
rect 0 3428 1040 3440
rect 0 3372 12 3428
rect 68 3372 332 3428
rect 388 3372 652 3428
rect 708 3372 972 3428
rect 1028 3372 1040 3428
rect 0 3360 1040 3372
rect 28960 3428 30000 3440
rect 28960 3372 28972 3428
rect 29028 3372 29292 3428
rect 29348 3372 29612 3428
rect 29668 3372 29932 3428
rect 29988 3372 30000 3428
rect 28960 3360 30000 3372
rect 0 3268 1040 3280
rect 0 3212 12 3268
rect 68 3212 332 3268
rect 388 3212 652 3268
rect 708 3212 972 3268
rect 1028 3212 1040 3268
rect 0 3200 1040 3212
rect 28960 3268 30000 3280
rect 28960 3212 28972 3268
rect 29028 3212 29292 3268
rect 29348 3212 29612 3268
rect 29668 3212 29932 3268
rect 29988 3212 30000 3268
rect 28960 3200 30000 3212
rect 0 3108 1040 3120
rect 0 3052 12 3108
rect 68 3052 332 3108
rect 388 3052 652 3108
rect 708 3052 972 3108
rect 1028 3052 1040 3108
rect 0 3040 1040 3052
rect 28960 3108 30000 3120
rect 28960 3052 28972 3108
rect 29028 3052 29292 3108
rect 29348 3052 29612 3108
rect 29668 3052 29932 3108
rect 29988 3052 30000 3108
rect 28960 3040 30000 3052
rect 0 2948 1040 2960
rect 0 2892 12 2948
rect 68 2892 332 2948
rect 388 2892 652 2948
rect 708 2892 972 2948
rect 1028 2892 1040 2948
rect 0 2880 1040 2892
rect 28960 2948 30000 2960
rect 28960 2892 28972 2948
rect 29028 2892 29292 2948
rect 29348 2892 29612 2948
rect 29668 2892 29932 2948
rect 29988 2892 30000 2948
rect 28960 2880 30000 2892
rect 0 2788 1040 2800
rect 0 2732 12 2788
rect 68 2732 332 2788
rect 388 2732 652 2788
rect 708 2732 972 2788
rect 1028 2732 1040 2788
rect 0 2720 1040 2732
rect 28960 2788 30000 2800
rect 28960 2732 28972 2788
rect 29028 2732 29292 2788
rect 29348 2732 29612 2788
rect 29668 2732 29932 2788
rect 29988 2732 30000 2788
rect 28960 2720 30000 2732
rect 0 2628 1040 2640
rect 0 2572 12 2628
rect 68 2572 332 2628
rect 388 2572 652 2628
rect 708 2572 972 2628
rect 1028 2572 1040 2628
rect 0 2560 1040 2572
rect 28960 2628 30000 2640
rect 28960 2572 28972 2628
rect 29028 2572 29292 2628
rect 29348 2572 29612 2628
rect 29668 2572 29932 2628
rect 29988 2572 30000 2628
rect 28960 2560 30000 2572
rect 0 2468 1040 2480
rect 0 2412 12 2468
rect 68 2412 332 2468
rect 388 2412 652 2468
rect 708 2412 972 2468
rect 1028 2412 1040 2468
rect 0 2400 1040 2412
rect 28960 2468 30000 2480
rect 28960 2412 28972 2468
rect 29028 2412 29292 2468
rect 29348 2412 29612 2468
rect 29668 2412 29932 2468
rect 29988 2412 30000 2468
rect 28960 2400 30000 2412
rect 0 2308 1040 2320
rect 0 2252 12 2308
rect 68 2252 332 2308
rect 388 2252 652 2308
rect 708 2252 972 2308
rect 1028 2252 1040 2308
rect 0 2240 1040 2252
rect 28960 2308 30000 2320
rect 28960 2252 28972 2308
rect 29028 2252 29292 2308
rect 29348 2252 29612 2308
rect 29668 2252 29932 2308
rect 29988 2252 30000 2308
rect 28960 2240 30000 2252
rect 0 2148 1040 2160
rect 0 2092 12 2148
rect 68 2092 332 2148
rect 388 2092 652 2148
rect 708 2092 972 2148
rect 1028 2092 1040 2148
rect 0 2080 1040 2092
rect 28960 2148 30000 2160
rect 28960 2092 28972 2148
rect 29028 2092 29292 2148
rect 29348 2092 29612 2148
rect 29668 2092 29932 2148
rect 29988 2092 30000 2148
rect 28960 2080 30000 2092
rect 0 1988 1040 2000
rect 0 1932 12 1988
rect 68 1932 332 1988
rect 388 1932 652 1988
rect 708 1932 972 1988
rect 1028 1932 1040 1988
rect 0 1920 1040 1932
rect 28960 1988 30000 2000
rect 28960 1932 28972 1988
rect 29028 1932 29292 1988
rect 29348 1932 29612 1988
rect 29668 1932 29932 1988
rect 29988 1932 30000 1988
rect 28960 1920 30000 1932
rect 0 1828 1040 1840
rect 0 1772 12 1828
rect 68 1772 332 1828
rect 388 1772 652 1828
rect 708 1772 972 1828
rect 1028 1772 1040 1828
rect 0 1760 1040 1772
rect 28960 1828 30000 1840
rect 28960 1772 28972 1828
rect 29028 1772 29292 1828
rect 29348 1772 29612 1828
rect 29668 1772 29932 1828
rect 29988 1772 30000 1828
rect 28960 1760 30000 1772
rect 0 1668 1040 1680
rect 0 1612 12 1668
rect 68 1612 332 1668
rect 388 1612 652 1668
rect 708 1612 972 1668
rect 1028 1612 1040 1668
rect 0 1600 1040 1612
rect 28960 1668 30000 1680
rect 28960 1612 28972 1668
rect 29028 1612 29292 1668
rect 29348 1612 29612 1668
rect 29668 1612 29932 1668
rect 29988 1612 30000 1668
rect 28960 1600 30000 1612
rect 0 1508 1040 1520
rect 0 1452 12 1508
rect 68 1452 332 1508
rect 388 1452 652 1508
rect 708 1452 972 1508
rect 1028 1452 1040 1508
rect 0 1440 1040 1452
rect 28960 1508 30000 1520
rect 28960 1452 28972 1508
rect 29028 1452 29292 1508
rect 29348 1452 29612 1508
rect 29668 1452 29932 1508
rect 29988 1452 30000 1508
rect 28960 1440 30000 1452
rect 0 1348 1040 1360
rect 0 1292 12 1348
rect 68 1292 332 1348
rect 388 1292 652 1348
rect 708 1292 972 1348
rect 1028 1292 1040 1348
rect 0 1280 1040 1292
rect 28960 1348 30000 1360
rect 28960 1292 28972 1348
rect 29028 1292 29292 1348
rect 29348 1292 29612 1348
rect 29668 1292 29932 1348
rect 29988 1292 30000 1348
rect 28960 1280 30000 1292
rect 0 1188 1040 1200
rect 0 1132 12 1188
rect 68 1132 332 1188
rect 388 1132 652 1188
rect 708 1132 972 1188
rect 1028 1132 1040 1188
rect 0 1120 1040 1132
rect 28960 1188 30000 1200
rect 28960 1132 28972 1188
rect 29028 1132 29292 1188
rect 29348 1132 29612 1188
rect 29668 1132 29932 1188
rect 29988 1132 30000 1188
rect 28960 1120 30000 1132
rect 0 1028 1040 1040
rect 0 972 12 1028
rect 68 972 332 1028
rect 388 972 652 1028
rect 708 972 972 1028
rect 1028 972 1040 1028
rect 0 960 1040 972
rect 1120 1028 1200 1040
rect 1120 972 1132 1028
rect 1188 972 1200 1028
rect 1120 960 1200 972
rect 28800 1028 28880 1040
rect 28800 972 28812 1028
rect 28868 972 28880 1028
rect 28800 960 28880 972
rect 28960 1028 30000 1040
rect 28960 972 28972 1028
rect 29028 972 29292 1028
rect 29348 972 29612 1028
rect 29668 972 29932 1028
rect 29988 972 30000 1028
rect 28960 960 30000 972
<< via2 >>
rect 12 31852 68 31908
rect 332 31852 388 31908
rect 652 31852 708 31908
rect 972 31852 1028 31908
rect 28972 31852 29028 31908
rect 29292 31852 29348 31908
rect 29612 31852 29668 31908
rect 29932 31852 29988 31908
rect 12 31692 68 31748
rect 332 31692 388 31748
rect 652 31692 708 31748
rect 972 31692 1028 31748
rect 28972 31692 29028 31748
rect 29292 31692 29348 31748
rect 29612 31692 29668 31748
rect 29932 31692 29988 31748
rect 12 31532 68 31588
rect 332 31532 388 31588
rect 652 31532 708 31588
rect 972 31532 1028 31588
rect 28972 31532 29028 31588
rect 29292 31532 29348 31588
rect 29612 31532 29668 31588
rect 29932 31532 29988 31588
rect 12 31372 68 31428
rect 332 31372 388 31428
rect 652 31372 708 31428
rect 972 31372 1028 31428
rect 28972 31372 29028 31428
rect 29292 31372 29348 31428
rect 29612 31372 29668 31428
rect 29932 31372 29988 31428
rect 12 31212 68 31268
rect 332 31212 388 31268
rect 652 31212 708 31268
rect 972 31212 1028 31268
rect 28972 31212 29028 31268
rect 29292 31212 29348 31268
rect 29612 31212 29668 31268
rect 29932 31212 29988 31268
rect 12 31052 68 31108
rect 332 31052 388 31108
rect 652 31052 708 31108
rect 972 31052 1028 31108
rect 28972 31052 29028 31108
rect 29292 31052 29348 31108
rect 29612 31052 29668 31108
rect 29932 31052 29988 31108
rect 12 30892 68 30948
rect 332 30892 388 30948
rect 652 30892 708 30948
rect 972 30892 1028 30948
rect 28972 30892 29028 30948
rect 29292 30892 29348 30948
rect 29612 30892 29668 30948
rect 29932 30892 29988 30948
rect 12 30732 68 30788
rect 332 30732 388 30788
rect 652 30732 708 30788
rect 972 30732 1028 30788
rect 28972 30732 29028 30788
rect 29292 30732 29348 30788
rect 29612 30732 29668 30788
rect 29932 30732 29988 30788
rect 12 30572 68 30628
rect 332 30572 388 30628
rect 652 30572 708 30628
rect 972 30572 1028 30628
rect 28972 30572 29028 30628
rect 29292 30572 29348 30628
rect 29612 30572 29668 30628
rect 29932 30572 29988 30628
rect 12 30412 68 30468
rect 332 30412 388 30468
rect 652 30412 708 30468
rect 972 30412 1028 30468
rect 28972 30412 29028 30468
rect 29292 30412 29348 30468
rect 29612 30412 29668 30468
rect 29932 30412 29988 30468
rect 12 30252 68 30308
rect 332 30252 388 30308
rect 652 30252 708 30308
rect 972 30252 1028 30308
rect 28972 30252 29028 30308
rect 29292 30252 29348 30308
rect 29612 30252 29668 30308
rect 29932 30252 29988 30308
rect 12 30092 68 30148
rect 332 30092 388 30148
rect 652 30092 708 30148
rect 972 30092 1028 30148
rect 28972 30092 29028 30148
rect 29292 30092 29348 30148
rect 29612 30092 29668 30148
rect 29932 30092 29988 30148
rect 12 29932 68 29988
rect 332 29932 388 29988
rect 652 29932 708 29988
rect 972 29932 1028 29988
rect 28972 29932 29028 29988
rect 29292 29932 29348 29988
rect 29612 29932 29668 29988
rect 29932 29932 29988 29988
rect 12 29772 68 29828
rect 332 29772 388 29828
rect 652 29772 708 29828
rect 972 29772 1028 29828
rect 28972 29772 29028 29828
rect 29292 29772 29348 29828
rect 29612 29772 29668 29828
rect 29932 29772 29988 29828
rect 12 29612 68 29668
rect 332 29612 388 29668
rect 652 29612 708 29668
rect 972 29612 1028 29668
rect 28972 29612 29028 29668
rect 29292 29612 29348 29668
rect 29612 29612 29668 29668
rect 29932 29612 29988 29668
rect 12 29452 68 29508
rect 332 29452 388 29508
rect 652 29452 708 29508
rect 972 29452 1028 29508
rect 28972 29452 29028 29508
rect 29292 29452 29348 29508
rect 29612 29452 29668 29508
rect 29932 29452 29988 29508
rect 12 29292 68 29348
rect 332 29292 388 29348
rect 652 29292 708 29348
rect 972 29292 1028 29348
rect 28972 29292 29028 29348
rect 29292 29292 29348 29348
rect 29612 29292 29668 29348
rect 29932 29292 29988 29348
rect 12 29132 68 29188
rect 332 29132 388 29188
rect 652 29132 708 29188
rect 972 29132 1028 29188
rect 12 28972 68 29028
rect 332 28972 388 29028
rect 652 28972 708 29028
rect 972 28972 1028 29028
rect 28972 28972 29028 29028
rect 29292 28972 29348 29028
rect 29612 28972 29668 29028
rect 29932 28972 29988 29028
rect 12 28812 68 28868
rect 332 28812 388 28868
rect 652 28812 708 28868
rect 972 28812 1028 28868
rect 29612 28812 29668 28868
rect 29932 28812 29988 28868
rect 12 28652 68 28708
rect 332 28652 388 28708
rect 652 28652 708 28708
rect 972 28652 1028 28708
rect 28972 28652 29028 28708
rect 29292 28652 29348 28708
rect 29612 28652 29668 28708
rect 29932 28652 29988 28708
rect 12 28492 68 28548
rect 332 28492 388 28548
rect 652 28492 708 28548
rect 972 28492 1028 28548
rect 28972 28492 29028 28548
rect 29292 28492 29348 28548
rect 29612 28492 29668 28548
rect 29932 28492 29988 28548
rect 12 28332 68 28388
rect 332 28332 388 28388
rect 652 28332 708 28388
rect 972 28332 1028 28388
rect 28972 28332 29028 28388
rect 29292 28332 29348 28388
rect 29612 28332 29668 28388
rect 29932 28332 29988 28388
rect 12 28172 68 28228
rect 332 28172 388 28228
rect 652 28172 708 28228
rect 972 28172 1028 28228
rect 28972 28172 29028 28228
rect 29292 28172 29348 28228
rect 29612 28172 29668 28228
rect 29932 28172 29988 28228
rect 12 28012 68 28068
rect 332 28012 388 28068
rect 652 28012 708 28068
rect 972 28012 1028 28068
rect 28972 28012 29028 28068
rect 29292 28012 29348 28068
rect 29612 28012 29668 28068
rect 29932 28012 29988 28068
rect 12 27852 68 27908
rect 332 27852 388 27908
rect 652 27852 708 27908
rect 972 27852 1028 27908
rect 28972 27852 29028 27908
rect 29292 27852 29348 27908
rect 29612 27852 29668 27908
rect 29932 27852 29988 27908
rect 12 27692 68 27748
rect 332 27692 388 27748
rect 652 27692 708 27748
rect 972 27692 1028 27748
rect 28972 27692 29028 27748
rect 29292 27692 29348 27748
rect 29612 27692 29668 27748
rect 29932 27692 29988 27748
rect 12 27532 68 27588
rect 332 27532 388 27588
rect 652 27532 708 27588
rect 972 27532 1028 27588
rect 28972 27532 29028 27588
rect 29292 27532 29348 27588
rect 29612 27532 29668 27588
rect 29932 27532 29988 27588
rect 12 27372 68 27428
rect 332 27372 388 27428
rect 652 27372 708 27428
rect 972 27372 1028 27428
rect 28972 27372 29028 27428
rect 29292 27372 29348 27428
rect 29612 27372 29668 27428
rect 29932 27372 29988 27428
rect 12 27212 68 27268
rect 332 27212 388 27268
rect 652 27212 708 27268
rect 972 27212 1028 27268
rect 28972 27212 29028 27268
rect 29292 27212 29348 27268
rect 29612 27212 29668 27268
rect 29932 27212 29988 27268
rect 12 27052 68 27108
rect 332 27052 388 27108
rect 652 27052 708 27108
rect 972 27052 1028 27108
rect 28972 27052 29028 27108
rect 29292 27052 29348 27108
rect 29612 27052 29668 27108
rect 29932 27052 29988 27108
rect 12 26892 68 26948
rect 332 26892 388 26948
rect 652 26892 708 26948
rect 972 26892 1028 26948
rect 28972 26892 29028 26948
rect 29292 26892 29348 26948
rect 29612 26892 29668 26948
rect 29932 26892 29988 26948
rect 12 26732 68 26788
rect 332 26732 388 26788
rect 652 26732 708 26788
rect 972 26732 1028 26788
rect 28972 26732 29028 26788
rect 29292 26732 29348 26788
rect 29612 26732 29668 26788
rect 29932 26732 29988 26788
rect 12 26572 68 26628
rect 332 26572 388 26628
rect 652 26572 708 26628
rect 972 26572 1028 26628
rect 28972 26572 29028 26628
rect 29292 26572 29348 26628
rect 29612 26572 29668 26628
rect 29932 26572 29988 26628
rect 12 26412 68 26468
rect 332 26412 388 26468
rect 652 26412 708 26468
rect 972 26412 1028 26468
rect 28972 26412 29028 26468
rect 29292 26412 29348 26468
rect 29612 26412 29668 26468
rect 29932 26412 29988 26468
rect 12 26252 68 26308
rect 332 26252 388 26308
rect 652 26252 708 26308
rect 972 26252 1028 26308
rect 29292 26252 29348 26308
rect 29612 26252 29668 26308
rect 29932 26252 29988 26308
rect 12 26092 68 26148
rect 332 26092 388 26148
rect 652 26092 708 26148
rect 972 26092 1028 26148
rect 28972 26092 29028 26148
rect 29292 26092 29348 26148
rect 29612 26092 29668 26148
rect 29932 26092 29988 26148
rect 12 25932 68 25988
rect 332 25932 388 25988
rect 652 25932 708 25988
rect 972 25932 1028 25988
rect 28972 25932 29028 25988
rect 29292 25932 29348 25988
rect 29612 25932 29668 25988
rect 29932 25932 29988 25988
rect 12 25772 68 25828
rect 332 25772 388 25828
rect 652 25772 708 25828
rect 972 25772 1028 25828
rect 28972 25772 29028 25828
rect 29292 25772 29348 25828
rect 29612 25772 29668 25828
rect 29932 25772 29988 25828
rect 12 25612 68 25668
rect 332 25612 388 25668
rect 652 25612 708 25668
rect 972 25612 1028 25668
rect 28972 25612 29028 25668
rect 29292 25612 29348 25668
rect 29612 25612 29668 25668
rect 29932 25612 29988 25668
rect 12 25452 68 25508
rect 332 25452 388 25508
rect 652 25452 708 25508
rect 972 25452 1028 25508
rect 28972 25452 29028 25508
rect 29292 25452 29348 25508
rect 29612 25452 29668 25508
rect 29932 25452 29988 25508
rect 12 25292 68 25348
rect 332 25292 388 25348
rect 652 25292 708 25348
rect 972 25292 1028 25348
rect 28972 25292 29028 25348
rect 29292 25292 29348 25348
rect 29612 25292 29668 25348
rect 29932 25292 29988 25348
rect 12 25132 68 25188
rect 332 25132 388 25188
rect 652 25132 708 25188
rect 972 25132 1028 25188
rect 28972 25132 29028 25188
rect 29292 25132 29348 25188
rect 29612 25132 29668 25188
rect 29932 25132 29988 25188
rect 12 24972 68 25028
rect 332 24972 388 25028
rect 652 24972 708 25028
rect 972 24972 1028 25028
rect 28972 24972 29028 25028
rect 29292 24972 29348 25028
rect 29612 24972 29668 25028
rect 29932 24972 29988 25028
rect 12 24812 68 24868
rect 332 24812 388 24868
rect 652 24812 708 24868
rect 972 24812 1028 24868
rect 28972 24812 29028 24868
rect 29292 24812 29348 24868
rect 29612 24812 29668 24868
rect 29932 24812 29988 24868
rect 12 24652 68 24708
rect 332 24652 388 24708
rect 652 24652 708 24708
rect 972 24652 1028 24708
rect 28972 24652 29028 24708
rect 29292 24652 29348 24708
rect 29612 24652 29668 24708
rect 29932 24652 29988 24708
rect 12 24492 68 24548
rect 332 24492 388 24548
rect 652 24492 708 24548
rect 972 24492 1028 24548
rect 28972 24492 29028 24548
rect 29292 24492 29348 24548
rect 29612 24492 29668 24548
rect 29932 24492 29988 24548
rect 12 24332 68 24388
rect 332 24332 388 24388
rect 652 24332 708 24388
rect 972 24332 1028 24388
rect 28972 24332 29028 24388
rect 29292 24332 29348 24388
rect 29612 24332 29668 24388
rect 29932 24332 29988 24388
rect 12 24172 68 24228
rect 332 24172 388 24228
rect 652 24172 708 24228
rect 972 24172 1028 24228
rect 28972 24172 29028 24228
rect 29292 24172 29348 24228
rect 29612 24172 29668 24228
rect 29932 24172 29988 24228
rect 12 24012 68 24068
rect 332 24012 388 24068
rect 652 24012 708 24068
rect 972 24012 1028 24068
rect 28972 24012 29028 24068
rect 29292 24012 29348 24068
rect 29612 24012 29668 24068
rect 29932 24012 29988 24068
rect 12 23852 68 23908
rect 332 23852 388 23908
rect 652 23852 708 23908
rect 972 23852 1028 23908
rect 28972 23852 29028 23908
rect 29292 23852 29348 23908
rect 29612 23852 29668 23908
rect 29932 23852 29988 23908
rect 12 23692 68 23748
rect 332 23692 388 23748
rect 652 23692 708 23748
rect 972 23692 1028 23748
rect 29612 23692 29668 23748
rect 29932 23692 29988 23748
rect 12 23532 68 23588
rect 332 23532 388 23588
rect 652 23532 708 23588
rect 972 23532 1028 23588
rect 28972 23532 29028 23588
rect 29292 23532 29348 23588
rect 29612 23532 29668 23588
rect 29932 23532 29988 23588
rect 12 23372 68 23428
rect 332 23372 388 23428
rect 652 23372 708 23428
rect 972 23372 1028 23428
rect 12 23212 68 23268
rect 332 23212 388 23268
rect 652 23212 708 23268
rect 972 23212 1028 23268
rect 28972 23212 29028 23268
rect 29292 23212 29348 23268
rect 29612 23212 29668 23268
rect 29932 23212 29988 23268
rect 12 23052 68 23108
rect 332 23052 388 23108
rect 652 23052 708 23108
rect 972 23052 1028 23108
rect 28972 23052 29028 23108
rect 29292 23052 29348 23108
rect 29612 23052 29668 23108
rect 29932 23052 29988 23108
rect 12 22892 68 22948
rect 332 22892 388 22948
rect 652 22892 708 22948
rect 972 22892 1028 22948
rect 28972 22892 29028 22948
rect 29292 22892 29348 22948
rect 29612 22892 29668 22948
rect 29932 22892 29988 22948
rect 12 22732 68 22788
rect 332 22732 388 22788
rect 652 22732 708 22788
rect 972 22732 1028 22788
rect 28972 22732 29028 22788
rect 29292 22732 29348 22788
rect 29612 22732 29668 22788
rect 29932 22732 29988 22788
rect 28972 22572 29028 22628
rect 29292 22572 29348 22628
rect 29612 22572 29668 22628
rect 29932 22572 29988 22628
rect 12 22412 68 22468
rect 332 22412 388 22468
rect 652 22412 708 22468
rect 972 22412 1028 22468
rect 28972 22412 29028 22468
rect 29292 22412 29348 22468
rect 29612 22412 29668 22468
rect 29932 22412 29988 22468
rect 12 22252 68 22308
rect 332 22252 388 22308
rect 28972 22252 29028 22308
rect 29292 22252 29348 22308
rect 29612 22252 29668 22308
rect 29932 22252 29988 22308
rect 12 22092 68 22148
rect 332 22092 388 22148
rect 652 22092 708 22148
rect 972 22092 1028 22148
rect 28972 22092 29028 22148
rect 29292 22092 29348 22148
rect 29612 22092 29668 22148
rect 29932 22092 29988 22148
rect 12 21932 68 21988
rect 332 21932 388 21988
rect 652 21932 708 21988
rect 972 21932 1028 21988
rect 28972 21932 29028 21988
rect 29292 21932 29348 21988
rect 29612 21932 29668 21988
rect 29932 21932 29988 21988
rect 12 21772 68 21828
rect 332 21772 388 21828
rect 652 21772 708 21828
rect 972 21772 1028 21828
rect 28972 21772 29028 21828
rect 29292 21772 29348 21828
rect 29612 21772 29668 21828
rect 29932 21772 29988 21828
rect 12 21612 68 21668
rect 332 21612 388 21668
rect 652 21612 708 21668
rect 972 21612 1028 21668
rect 28972 21612 29028 21668
rect 29292 21612 29348 21668
rect 29612 21612 29668 21668
rect 29932 21612 29988 21668
rect 12 21452 68 21508
rect 332 21452 388 21508
rect 652 21452 708 21508
rect 972 21452 1028 21508
rect 28972 21452 29028 21508
rect 29292 21452 29348 21508
rect 29612 21452 29668 21508
rect 29932 21452 29988 21508
rect 12 21292 68 21348
rect 332 21292 388 21348
rect 652 21292 708 21348
rect 972 21292 1028 21348
rect 28972 21292 29028 21348
rect 29292 21292 29348 21348
rect 29612 21292 29668 21348
rect 29932 21292 29988 21348
rect 12 21132 68 21188
rect 332 21132 388 21188
rect 652 21132 708 21188
rect 972 21132 1028 21188
rect 28972 21132 29028 21188
rect 29292 21132 29348 21188
rect 29612 21132 29668 21188
rect 29932 21132 29988 21188
rect 12 20972 68 21028
rect 332 20972 388 21028
rect 652 20972 708 21028
rect 972 20972 1028 21028
rect 28972 20972 29028 21028
rect 29292 20972 29348 21028
rect 29612 20972 29668 21028
rect 29932 20972 29988 21028
rect 12 20812 68 20868
rect 332 20812 388 20868
rect 652 20812 708 20868
rect 972 20812 1028 20868
rect 28972 20812 29028 20868
rect 29292 20812 29348 20868
rect 29612 20812 29668 20868
rect 29932 20812 29988 20868
rect 12 20652 68 20708
rect 332 20652 388 20708
rect 652 20652 708 20708
rect 972 20652 1028 20708
rect 28972 20652 29028 20708
rect 29292 20652 29348 20708
rect 29612 20652 29668 20708
rect 29932 20652 29988 20708
rect 12 20492 68 20548
rect 332 20492 388 20548
rect 652 20492 708 20548
rect 972 20492 1028 20548
rect 28972 20492 29028 20548
rect 29292 20492 29348 20548
rect 29612 20492 29668 20548
rect 29932 20492 29988 20548
rect 12 20332 68 20388
rect 332 20332 388 20388
rect 652 20332 708 20388
rect 972 20332 1028 20388
rect 28972 20332 29028 20388
rect 29292 20332 29348 20388
rect 29612 20332 29668 20388
rect 29932 20332 29988 20388
rect 12 20172 68 20228
rect 332 20172 388 20228
rect 652 20172 708 20228
rect 972 20172 1028 20228
rect 28972 20172 29028 20228
rect 29292 20172 29348 20228
rect 29612 20172 29668 20228
rect 29932 20172 29988 20228
rect 12 20012 68 20068
rect 332 20012 388 20068
rect 652 20012 708 20068
rect 972 20012 1028 20068
rect 28972 20012 29028 20068
rect 29292 20012 29348 20068
rect 29612 20012 29668 20068
rect 29932 20012 29988 20068
rect 12 19852 68 19908
rect 332 19852 388 19908
rect 652 19852 708 19908
rect 972 19852 1028 19908
rect 28972 19852 29028 19908
rect 29292 19852 29348 19908
rect 29612 19852 29668 19908
rect 29932 19852 29988 19908
rect 12 19692 68 19748
rect 332 19692 388 19748
rect 652 19692 708 19748
rect 28972 19692 29028 19748
rect 29292 19692 29348 19748
rect 29612 19692 29668 19748
rect 29932 19692 29988 19748
rect 12 19532 68 19588
rect 332 19532 388 19588
rect 652 19532 708 19588
rect 972 19532 1028 19588
rect 28972 19532 29028 19588
rect 29292 19532 29348 19588
rect 29612 19532 29668 19588
rect 29932 19532 29988 19588
rect 12 19372 68 19428
rect 332 19372 388 19428
rect 652 19372 708 19428
rect 972 19372 1028 19428
rect 28972 19372 29028 19428
rect 29292 19372 29348 19428
rect 29612 19372 29668 19428
rect 29932 19372 29988 19428
rect 12 19212 68 19268
rect 332 19212 388 19268
rect 652 19212 708 19268
rect 972 19212 1028 19268
rect 28972 19212 29028 19268
rect 29292 19212 29348 19268
rect 29612 19212 29668 19268
rect 29932 19212 29988 19268
rect 12 19052 68 19108
rect 332 19052 388 19108
rect 652 19052 708 19108
rect 972 19052 1028 19108
rect 28972 19052 29028 19108
rect 29292 19052 29348 19108
rect 29612 19052 29668 19108
rect 29932 19052 29988 19108
rect 12 18892 68 18948
rect 332 18892 388 18948
rect 652 18892 708 18948
rect 972 18892 1028 18948
rect 28972 18892 29028 18948
rect 29292 18892 29348 18948
rect 29612 18892 29668 18948
rect 29932 18892 29988 18948
rect 12 18732 68 18788
rect 332 18732 388 18788
rect 652 18732 708 18788
rect 972 18732 1028 18788
rect 28972 18732 29028 18788
rect 29292 18732 29348 18788
rect 29612 18732 29668 18788
rect 29932 18732 29988 18788
rect 12 18572 68 18628
rect 332 18572 388 18628
rect 652 18572 708 18628
rect 972 18572 1028 18628
rect 28972 18572 29028 18628
rect 29292 18572 29348 18628
rect 29612 18572 29668 18628
rect 29932 18572 29988 18628
rect 12 18412 68 18468
rect 332 18412 388 18468
rect 652 18412 708 18468
rect 972 18412 1028 18468
rect 28972 18412 29028 18468
rect 29292 18412 29348 18468
rect 29612 18412 29668 18468
rect 29932 18412 29988 18468
rect 12 18252 68 18308
rect 332 18252 388 18308
rect 652 18252 708 18308
rect 972 18252 1028 18308
rect 28972 18252 29028 18308
rect 29292 18252 29348 18308
rect 29612 18252 29668 18308
rect 29932 18252 29988 18308
rect 12 18092 68 18148
rect 332 18092 388 18148
rect 652 18092 708 18148
rect 972 18092 1028 18148
rect 28972 18092 29028 18148
rect 29292 18092 29348 18148
rect 29612 18092 29668 18148
rect 29932 18092 29988 18148
rect 12 17932 68 17988
rect 332 17932 388 17988
rect 652 17932 708 17988
rect 972 17932 1028 17988
rect 28972 17932 29028 17988
rect 29292 17932 29348 17988
rect 29612 17932 29668 17988
rect 29932 17932 29988 17988
rect 12 17772 68 17828
rect 332 17772 388 17828
rect 652 17772 708 17828
rect 972 17772 1028 17828
rect 28972 17772 29028 17828
rect 29292 17772 29348 17828
rect 29612 17772 29668 17828
rect 29932 17772 29988 17828
rect 12 17612 68 17668
rect 332 17612 388 17668
rect 652 17612 708 17668
rect 972 17612 1028 17668
rect 28972 17612 29028 17668
rect 29292 17612 29348 17668
rect 29612 17612 29668 17668
rect 29932 17612 29988 17668
rect 12 17452 68 17508
rect 332 17452 388 17508
rect 652 17452 708 17508
rect 972 17452 1028 17508
rect 28972 17452 29028 17508
rect 29292 17452 29348 17508
rect 29612 17452 29668 17508
rect 29932 17452 29988 17508
rect 12 17292 68 17348
rect 332 17292 388 17348
rect 652 17292 708 17348
rect 972 17292 1028 17348
rect 28972 17292 29028 17348
rect 29292 17292 29348 17348
rect 29612 17292 29668 17348
rect 29932 17292 29988 17348
rect 12 17132 68 17188
rect 332 17132 388 17188
rect 28972 17132 29028 17188
rect 29292 17132 29348 17188
rect 29612 17132 29668 17188
rect 29932 17132 29988 17188
rect 12 16972 68 17028
rect 332 16972 388 17028
rect 652 16972 708 17028
rect 972 16972 1028 17028
rect 28972 16972 29028 17028
rect 29292 16972 29348 17028
rect 29612 16972 29668 17028
rect 29932 16972 29988 17028
rect 28972 16812 29028 16868
rect 29292 16812 29348 16868
rect 29612 16812 29668 16868
rect 29932 16812 29988 16868
rect 12 16652 68 16708
rect 332 16652 388 16708
rect 652 16652 708 16708
rect 972 16652 1028 16708
rect 28972 16652 29028 16708
rect 29292 16652 29348 16708
rect 29612 16652 29668 16708
rect 29932 16652 29988 16708
rect 12 16492 68 16548
rect 332 16492 388 16548
rect 652 16492 708 16548
rect 972 16492 1028 16548
rect 28972 16492 29028 16548
rect 29292 16492 29348 16548
rect 29612 16492 29668 16548
rect 29932 16492 29988 16548
rect 12 16332 68 16388
rect 332 16332 388 16388
rect 652 16332 708 16388
rect 972 16332 1028 16388
rect 28972 16332 29028 16388
rect 29292 16332 29348 16388
rect 29612 16332 29668 16388
rect 29932 16332 29988 16388
rect 12 16172 68 16228
rect 332 16172 388 16228
rect 652 16172 708 16228
rect 972 16172 1028 16228
rect 28972 16172 29028 16228
rect 29292 16172 29348 16228
rect 29612 16172 29668 16228
rect 29932 16172 29988 16228
rect 28972 16012 29028 16068
rect 29292 16012 29348 16068
rect 29612 16012 29668 16068
rect 29932 16012 29988 16068
rect 12 15852 68 15908
rect 332 15852 388 15908
rect 652 15852 708 15908
rect 972 15852 1028 15908
rect 28972 15852 29028 15908
rect 29292 15852 29348 15908
rect 29612 15852 29668 15908
rect 29932 15852 29988 15908
rect 12 15692 68 15748
rect 332 15692 388 15748
rect 28972 15692 29028 15748
rect 29292 15692 29348 15748
rect 29612 15692 29668 15748
rect 29932 15692 29988 15748
rect 12 15532 68 15588
rect 332 15532 388 15588
rect 652 15532 708 15588
rect 972 15532 1028 15588
rect 28972 15532 29028 15588
rect 29292 15532 29348 15588
rect 29612 15532 29668 15588
rect 29932 15532 29988 15588
rect 12 15372 68 15428
rect 332 15372 388 15428
rect 652 15372 708 15428
rect 972 15372 1028 15428
rect 28972 15372 29028 15428
rect 29292 15372 29348 15428
rect 29612 15372 29668 15428
rect 29932 15372 29988 15428
rect 12 15212 68 15268
rect 332 15212 388 15268
rect 652 15212 708 15268
rect 972 15212 1028 15268
rect 28972 15212 29028 15268
rect 29292 15212 29348 15268
rect 29612 15212 29668 15268
rect 29932 15212 29988 15268
rect 12 15052 68 15108
rect 332 15052 388 15108
rect 652 15052 708 15108
rect 972 15052 1028 15108
rect 28972 15052 29028 15108
rect 29292 15052 29348 15108
rect 29612 15052 29668 15108
rect 29932 15052 29988 15108
rect 12 14892 68 14948
rect 332 14892 388 14948
rect 652 14892 708 14948
rect 972 14892 1028 14948
rect 28972 14892 29028 14948
rect 29292 14892 29348 14948
rect 29612 14892 29668 14948
rect 29932 14892 29988 14948
rect 12 14732 68 14788
rect 332 14732 388 14788
rect 652 14732 708 14788
rect 972 14732 1028 14788
rect 28972 14732 29028 14788
rect 29292 14732 29348 14788
rect 29612 14732 29668 14788
rect 29932 14732 29988 14788
rect 12 14572 68 14628
rect 332 14572 388 14628
rect 652 14572 708 14628
rect 972 14572 1028 14628
rect 28972 14572 29028 14628
rect 29292 14572 29348 14628
rect 29612 14572 29668 14628
rect 29932 14572 29988 14628
rect 12 14412 68 14468
rect 332 14412 388 14468
rect 652 14412 708 14468
rect 972 14412 1028 14468
rect 28972 14412 29028 14468
rect 29292 14412 29348 14468
rect 29612 14412 29668 14468
rect 29932 14412 29988 14468
rect 12 14252 68 14308
rect 332 14252 388 14308
rect 652 14252 708 14308
rect 972 14252 1028 14308
rect 28972 14252 29028 14308
rect 29292 14252 29348 14308
rect 29612 14252 29668 14308
rect 29932 14252 29988 14308
rect 12 14092 68 14148
rect 332 14092 388 14148
rect 652 14092 708 14148
rect 972 14092 1028 14148
rect 28972 14092 29028 14148
rect 29292 14092 29348 14148
rect 29612 14092 29668 14148
rect 29932 14092 29988 14148
rect 12 13932 68 13988
rect 332 13932 388 13988
rect 652 13932 708 13988
rect 972 13932 1028 13988
rect 28972 13932 29028 13988
rect 29292 13932 29348 13988
rect 29612 13932 29668 13988
rect 29932 13932 29988 13988
rect 12 13772 68 13828
rect 332 13772 388 13828
rect 652 13772 708 13828
rect 972 13772 1028 13828
rect 28972 13772 29028 13828
rect 29292 13772 29348 13828
rect 29612 13772 29668 13828
rect 29932 13772 29988 13828
rect 12 13612 68 13668
rect 332 13612 388 13668
rect 652 13612 708 13668
rect 972 13612 1028 13668
rect 28972 13612 29028 13668
rect 29292 13612 29348 13668
rect 29612 13612 29668 13668
rect 29932 13612 29988 13668
rect 12 13452 68 13508
rect 332 13452 388 13508
rect 652 13452 708 13508
rect 972 13452 1028 13508
rect 28972 13452 29028 13508
rect 29292 13452 29348 13508
rect 29612 13452 29668 13508
rect 29932 13452 29988 13508
rect 12 13292 68 13348
rect 332 13292 388 13348
rect 652 13292 708 13348
rect 972 13292 1028 13348
rect 28972 13292 29028 13348
rect 29292 13292 29348 13348
rect 29612 13292 29668 13348
rect 29932 13292 29988 13348
rect 12 13132 68 13188
rect 332 13132 388 13188
rect 652 13132 708 13188
rect 28972 13132 29028 13188
rect 29292 13132 29348 13188
rect 29612 13132 29668 13188
rect 29932 13132 29988 13188
rect 12 12972 68 13028
rect 332 12972 388 13028
rect 652 12972 708 13028
rect 972 12972 1028 13028
rect 28972 12972 29028 13028
rect 29292 12972 29348 13028
rect 29612 12972 29668 13028
rect 29932 12972 29988 13028
rect 12 12812 68 12868
rect 332 12812 388 12868
rect 652 12812 708 12868
rect 972 12812 1028 12868
rect 28972 12812 29028 12868
rect 29292 12812 29348 12868
rect 29612 12812 29668 12868
rect 29932 12812 29988 12868
rect 12 12652 68 12708
rect 332 12652 388 12708
rect 652 12652 708 12708
rect 972 12652 1028 12708
rect 28972 12652 29028 12708
rect 29292 12652 29348 12708
rect 29612 12652 29668 12708
rect 29932 12652 29988 12708
rect 12 12492 68 12548
rect 332 12492 388 12548
rect 652 12492 708 12548
rect 972 12492 1028 12548
rect 28972 12492 29028 12548
rect 29292 12492 29348 12548
rect 29612 12492 29668 12548
rect 29932 12492 29988 12548
rect 12 12332 68 12388
rect 332 12332 388 12388
rect 652 12332 708 12388
rect 972 12332 1028 12388
rect 28972 12332 29028 12388
rect 29292 12332 29348 12388
rect 29612 12332 29668 12388
rect 29932 12332 29988 12388
rect 12 12172 68 12228
rect 332 12172 388 12228
rect 652 12172 708 12228
rect 972 12172 1028 12228
rect 28972 12172 29028 12228
rect 29292 12172 29348 12228
rect 29612 12172 29668 12228
rect 29932 12172 29988 12228
rect 12 12012 68 12068
rect 332 12012 388 12068
rect 652 12012 708 12068
rect 972 12012 1028 12068
rect 28972 12012 29028 12068
rect 29292 12012 29348 12068
rect 29612 12012 29668 12068
rect 29932 12012 29988 12068
rect 12 11852 68 11908
rect 332 11852 388 11908
rect 652 11852 708 11908
rect 972 11852 1028 11908
rect 28972 11852 29028 11908
rect 29292 11852 29348 11908
rect 29612 11852 29668 11908
rect 29932 11852 29988 11908
rect 12 11692 68 11748
rect 332 11692 388 11748
rect 652 11692 708 11748
rect 972 11692 1028 11748
rect 28972 11692 29028 11748
rect 29292 11692 29348 11748
rect 29612 11692 29668 11748
rect 29932 11692 29988 11748
rect 12 11532 68 11588
rect 332 11532 388 11588
rect 652 11532 708 11588
rect 972 11532 1028 11588
rect 28972 11532 29028 11588
rect 29292 11532 29348 11588
rect 29612 11532 29668 11588
rect 29932 11532 29988 11588
rect 12 11372 68 11428
rect 332 11372 388 11428
rect 652 11372 708 11428
rect 972 11372 1028 11428
rect 28972 11372 29028 11428
rect 29292 11372 29348 11428
rect 29612 11372 29668 11428
rect 29932 11372 29988 11428
rect 12 11212 68 11268
rect 332 11212 388 11268
rect 652 11212 708 11268
rect 972 11212 1028 11268
rect 28972 11212 29028 11268
rect 29292 11212 29348 11268
rect 29612 11212 29668 11268
rect 29932 11212 29988 11268
rect 12 11052 68 11108
rect 332 11052 388 11108
rect 652 11052 708 11108
rect 972 11052 1028 11108
rect 28972 11052 29028 11108
rect 29292 11052 29348 11108
rect 29612 11052 29668 11108
rect 29932 11052 29988 11108
rect 12 10892 68 10948
rect 332 10892 388 10948
rect 652 10892 708 10948
rect 972 10892 1028 10948
rect 28972 10892 29028 10948
rect 29292 10892 29348 10948
rect 29612 10892 29668 10948
rect 29932 10892 29988 10948
rect 12 10732 68 10788
rect 332 10732 388 10788
rect 652 10732 708 10788
rect 972 10732 1028 10788
rect 28972 10732 29028 10788
rect 29292 10732 29348 10788
rect 29612 10732 29668 10788
rect 29932 10732 29988 10788
rect 12 10572 68 10628
rect 332 10572 388 10628
rect 28972 10572 29028 10628
rect 29292 10572 29348 10628
rect 29612 10572 29668 10628
rect 29932 10572 29988 10628
rect 12 10412 68 10468
rect 332 10412 388 10468
rect 652 10412 708 10468
rect 972 10412 1028 10468
rect 28972 10412 29028 10468
rect 29292 10412 29348 10468
rect 29612 10412 29668 10468
rect 29932 10412 29988 10468
rect 28972 10252 29028 10308
rect 29292 10252 29348 10308
rect 29612 10252 29668 10308
rect 29932 10252 29988 10308
rect 12 10092 68 10148
rect 332 10092 388 10148
rect 652 10092 708 10148
rect 972 10092 1028 10148
rect 28972 10092 29028 10148
rect 29292 10092 29348 10148
rect 29612 10092 29668 10148
rect 29932 10092 29988 10148
rect 12 9932 68 9988
rect 332 9932 388 9988
rect 652 9932 708 9988
rect 972 9932 1028 9988
rect 28972 9932 29028 9988
rect 29292 9932 29348 9988
rect 29612 9932 29668 9988
rect 29932 9932 29988 9988
rect 12 9772 68 9828
rect 332 9772 388 9828
rect 652 9772 708 9828
rect 972 9772 1028 9828
rect 28972 9772 29028 9828
rect 29292 9772 29348 9828
rect 29612 9772 29668 9828
rect 29932 9772 29988 9828
rect 12 9612 68 9668
rect 332 9612 388 9668
rect 652 9612 708 9668
rect 972 9612 1028 9668
rect 28972 9612 29028 9668
rect 29292 9612 29348 9668
rect 29612 9612 29668 9668
rect 29932 9612 29988 9668
rect 12 9452 68 9508
rect 332 9452 388 9508
rect 652 9452 708 9508
rect 972 9452 1028 9508
rect 12 9292 68 9348
rect 332 9292 388 9348
rect 652 9292 708 9348
rect 972 9292 1028 9348
rect 28972 9292 29028 9348
rect 29292 9292 29348 9348
rect 29612 9292 29668 9348
rect 29932 9292 29988 9348
rect 12 9132 68 9188
rect 332 9132 388 9188
rect 652 9132 708 9188
rect 972 9132 1028 9188
rect 29612 9132 29668 9188
rect 29932 9132 29988 9188
rect 12 8972 68 9028
rect 332 8972 388 9028
rect 652 8972 708 9028
rect 972 8972 1028 9028
rect 28972 8972 29028 9028
rect 29292 8972 29348 9028
rect 29612 8972 29668 9028
rect 29932 8972 29988 9028
rect 12 8812 68 8868
rect 332 8812 388 8868
rect 652 8812 708 8868
rect 972 8812 1028 8868
rect 28972 8812 29028 8868
rect 29292 8812 29348 8868
rect 29612 8812 29668 8868
rect 29932 8812 29988 8868
rect 12 8652 68 8708
rect 332 8652 388 8708
rect 652 8652 708 8708
rect 972 8652 1028 8708
rect 28972 8652 29028 8708
rect 29292 8652 29348 8708
rect 29612 8652 29668 8708
rect 29932 8652 29988 8708
rect 12 8492 68 8548
rect 332 8492 388 8548
rect 652 8492 708 8548
rect 972 8492 1028 8548
rect 28972 8492 29028 8548
rect 29292 8492 29348 8548
rect 29612 8492 29668 8548
rect 29932 8492 29988 8548
rect 12 8332 68 8388
rect 332 8332 388 8388
rect 652 8332 708 8388
rect 972 8332 1028 8388
rect 28972 8332 29028 8388
rect 29292 8332 29348 8388
rect 29612 8332 29668 8388
rect 29932 8332 29988 8388
rect 12 8172 68 8228
rect 332 8172 388 8228
rect 652 8172 708 8228
rect 972 8172 1028 8228
rect 28972 8172 29028 8228
rect 29292 8172 29348 8228
rect 29612 8172 29668 8228
rect 29932 8172 29988 8228
rect 12 8012 68 8068
rect 332 8012 388 8068
rect 652 8012 708 8068
rect 972 8012 1028 8068
rect 28972 8012 29028 8068
rect 29292 8012 29348 8068
rect 29612 8012 29668 8068
rect 29932 8012 29988 8068
rect 12 7852 68 7908
rect 332 7852 388 7908
rect 652 7852 708 7908
rect 972 7852 1028 7908
rect 28972 7852 29028 7908
rect 29292 7852 29348 7908
rect 29612 7852 29668 7908
rect 29932 7852 29988 7908
rect 12 7692 68 7748
rect 332 7692 388 7748
rect 652 7692 708 7748
rect 972 7692 1028 7748
rect 28972 7692 29028 7748
rect 29292 7692 29348 7748
rect 29612 7692 29668 7748
rect 29932 7692 29988 7748
rect 12 7532 68 7588
rect 332 7532 388 7588
rect 652 7532 708 7588
rect 972 7532 1028 7588
rect 28972 7532 29028 7588
rect 29292 7532 29348 7588
rect 29612 7532 29668 7588
rect 29932 7532 29988 7588
rect 12 7372 68 7428
rect 332 7372 388 7428
rect 652 7372 708 7428
rect 972 7372 1028 7428
rect 28972 7372 29028 7428
rect 29292 7372 29348 7428
rect 29612 7372 29668 7428
rect 29932 7372 29988 7428
rect 12 7212 68 7268
rect 332 7212 388 7268
rect 652 7212 708 7268
rect 972 7212 1028 7268
rect 28972 7212 29028 7268
rect 29292 7212 29348 7268
rect 29612 7212 29668 7268
rect 29932 7212 29988 7268
rect 12 7052 68 7108
rect 332 7052 388 7108
rect 652 7052 708 7108
rect 972 7052 1028 7108
rect 28972 7052 29028 7108
rect 29292 7052 29348 7108
rect 29612 7052 29668 7108
rect 29932 7052 29988 7108
rect 12 6892 68 6948
rect 332 6892 388 6948
rect 652 6892 708 6948
rect 972 6892 1028 6948
rect 28972 6892 29028 6948
rect 29292 6892 29348 6948
rect 29612 6892 29668 6948
rect 29932 6892 29988 6948
rect 12 6732 68 6788
rect 332 6732 388 6788
rect 652 6732 708 6788
rect 972 6732 1028 6788
rect 28972 6732 29028 6788
rect 29292 6732 29348 6788
rect 29612 6732 29668 6788
rect 29932 6732 29988 6788
rect 12 6572 68 6628
rect 332 6572 388 6628
rect 652 6572 708 6628
rect 972 6572 1028 6628
rect 29292 6572 29348 6628
rect 29612 6572 29668 6628
rect 29932 6572 29988 6628
rect 12 6412 68 6468
rect 332 6412 388 6468
rect 652 6412 708 6468
rect 972 6412 1028 6468
rect 28972 6412 29028 6468
rect 29292 6412 29348 6468
rect 29612 6412 29668 6468
rect 29932 6412 29988 6468
rect 12 6252 68 6308
rect 332 6252 388 6308
rect 652 6252 708 6308
rect 972 6252 1028 6308
rect 28972 6252 29028 6308
rect 29292 6252 29348 6308
rect 29612 6252 29668 6308
rect 29932 6252 29988 6308
rect 12 6092 68 6148
rect 332 6092 388 6148
rect 652 6092 708 6148
rect 972 6092 1028 6148
rect 28972 6092 29028 6148
rect 29292 6092 29348 6148
rect 29612 6092 29668 6148
rect 29932 6092 29988 6148
rect 12 5932 68 5988
rect 332 5932 388 5988
rect 652 5932 708 5988
rect 972 5932 1028 5988
rect 28972 5932 29028 5988
rect 29292 5932 29348 5988
rect 29612 5932 29668 5988
rect 29932 5932 29988 5988
rect 12 5772 68 5828
rect 332 5772 388 5828
rect 652 5772 708 5828
rect 972 5772 1028 5828
rect 28972 5772 29028 5828
rect 29292 5772 29348 5828
rect 29612 5772 29668 5828
rect 29932 5772 29988 5828
rect 12 5612 68 5668
rect 332 5612 388 5668
rect 652 5612 708 5668
rect 972 5612 1028 5668
rect 28972 5612 29028 5668
rect 29292 5612 29348 5668
rect 29612 5612 29668 5668
rect 29932 5612 29988 5668
rect 12 5452 68 5508
rect 332 5452 388 5508
rect 652 5452 708 5508
rect 972 5452 1028 5508
rect 28972 5452 29028 5508
rect 29292 5452 29348 5508
rect 29612 5452 29668 5508
rect 29932 5452 29988 5508
rect 12 5292 68 5348
rect 332 5292 388 5348
rect 652 5292 708 5348
rect 972 5292 1028 5348
rect 28972 5292 29028 5348
rect 29292 5292 29348 5348
rect 29612 5292 29668 5348
rect 29932 5292 29988 5348
rect 12 5132 68 5188
rect 332 5132 388 5188
rect 652 5132 708 5188
rect 972 5132 1028 5188
rect 28972 5132 29028 5188
rect 29292 5132 29348 5188
rect 29612 5132 29668 5188
rect 29932 5132 29988 5188
rect 12 4972 68 5028
rect 332 4972 388 5028
rect 652 4972 708 5028
rect 972 4972 1028 5028
rect 28972 4972 29028 5028
rect 29292 4972 29348 5028
rect 29612 4972 29668 5028
rect 29932 4972 29988 5028
rect 12 4812 68 4868
rect 332 4812 388 4868
rect 652 4812 708 4868
rect 972 4812 1028 4868
rect 28972 4812 29028 4868
rect 29292 4812 29348 4868
rect 29612 4812 29668 4868
rect 29932 4812 29988 4868
rect 12 4652 68 4708
rect 332 4652 388 4708
rect 652 4652 708 4708
rect 972 4652 1028 4708
rect 28972 4652 29028 4708
rect 29292 4652 29348 4708
rect 29612 4652 29668 4708
rect 29932 4652 29988 4708
rect 12 4492 68 4548
rect 332 4492 388 4548
rect 652 4492 708 4548
rect 972 4492 1028 4548
rect 28972 4492 29028 4548
rect 29292 4492 29348 4548
rect 29612 4492 29668 4548
rect 29932 4492 29988 4548
rect 12 4332 68 4388
rect 332 4332 388 4388
rect 652 4332 708 4388
rect 972 4332 1028 4388
rect 28972 4332 29028 4388
rect 29292 4332 29348 4388
rect 29612 4332 29668 4388
rect 29932 4332 29988 4388
rect 12 4172 68 4228
rect 332 4172 388 4228
rect 652 4172 708 4228
rect 972 4172 1028 4228
rect 28972 4172 29028 4228
rect 29292 4172 29348 4228
rect 29612 4172 29668 4228
rect 29932 4172 29988 4228
rect 12 4012 68 4068
rect 332 4012 388 4068
rect 652 4012 708 4068
rect 972 4012 1028 4068
rect 29612 4012 29668 4068
rect 29932 4012 29988 4068
rect 12 3852 68 3908
rect 332 3852 388 3908
rect 652 3852 708 3908
rect 972 3852 1028 3908
rect 28972 3852 29028 3908
rect 29292 3852 29348 3908
rect 29612 3852 29668 3908
rect 29932 3852 29988 3908
rect 12 3692 68 3748
rect 332 3692 388 3748
rect 652 3692 708 3748
rect 972 3692 1028 3748
rect 12 3532 68 3588
rect 332 3532 388 3588
rect 652 3532 708 3588
rect 972 3532 1028 3588
rect 28972 3532 29028 3588
rect 29292 3532 29348 3588
rect 29612 3532 29668 3588
rect 29932 3532 29988 3588
rect 12 3372 68 3428
rect 332 3372 388 3428
rect 652 3372 708 3428
rect 972 3372 1028 3428
rect 28972 3372 29028 3428
rect 29292 3372 29348 3428
rect 29612 3372 29668 3428
rect 29932 3372 29988 3428
rect 12 3212 68 3268
rect 332 3212 388 3268
rect 652 3212 708 3268
rect 972 3212 1028 3268
rect 28972 3212 29028 3268
rect 29292 3212 29348 3268
rect 29612 3212 29668 3268
rect 29932 3212 29988 3268
rect 12 3052 68 3108
rect 332 3052 388 3108
rect 652 3052 708 3108
rect 972 3052 1028 3108
rect 28972 3052 29028 3108
rect 29292 3052 29348 3108
rect 29612 3052 29668 3108
rect 29932 3052 29988 3108
rect 12 2892 68 2948
rect 332 2892 388 2948
rect 652 2892 708 2948
rect 972 2892 1028 2948
rect 28972 2892 29028 2948
rect 29292 2892 29348 2948
rect 29612 2892 29668 2948
rect 29932 2892 29988 2948
rect 12 2732 68 2788
rect 332 2732 388 2788
rect 652 2732 708 2788
rect 972 2732 1028 2788
rect 28972 2732 29028 2788
rect 29292 2732 29348 2788
rect 29612 2732 29668 2788
rect 29932 2732 29988 2788
rect 12 2572 68 2628
rect 332 2572 388 2628
rect 652 2572 708 2628
rect 972 2572 1028 2628
rect 28972 2572 29028 2628
rect 29292 2572 29348 2628
rect 29612 2572 29668 2628
rect 29932 2572 29988 2628
rect 12 2412 68 2468
rect 332 2412 388 2468
rect 652 2412 708 2468
rect 972 2412 1028 2468
rect 28972 2412 29028 2468
rect 29292 2412 29348 2468
rect 29612 2412 29668 2468
rect 29932 2412 29988 2468
rect 12 2252 68 2308
rect 332 2252 388 2308
rect 652 2252 708 2308
rect 972 2252 1028 2308
rect 28972 2252 29028 2308
rect 29292 2252 29348 2308
rect 29612 2252 29668 2308
rect 29932 2252 29988 2308
rect 12 2092 68 2148
rect 332 2092 388 2148
rect 652 2092 708 2148
rect 972 2092 1028 2148
rect 28972 2092 29028 2148
rect 29292 2092 29348 2148
rect 29612 2092 29668 2148
rect 29932 2092 29988 2148
rect 12 1932 68 1988
rect 332 1932 388 1988
rect 652 1932 708 1988
rect 972 1932 1028 1988
rect 28972 1932 29028 1988
rect 29292 1932 29348 1988
rect 29612 1932 29668 1988
rect 29932 1932 29988 1988
rect 12 1772 68 1828
rect 332 1772 388 1828
rect 652 1772 708 1828
rect 972 1772 1028 1828
rect 28972 1772 29028 1828
rect 29292 1772 29348 1828
rect 29612 1772 29668 1828
rect 29932 1772 29988 1828
rect 12 1612 68 1668
rect 332 1612 388 1668
rect 652 1612 708 1668
rect 972 1612 1028 1668
rect 28972 1612 29028 1668
rect 29292 1612 29348 1668
rect 29612 1612 29668 1668
rect 29932 1612 29988 1668
rect 12 1452 68 1508
rect 332 1452 388 1508
rect 652 1452 708 1508
rect 972 1452 1028 1508
rect 28972 1452 29028 1508
rect 29292 1452 29348 1508
rect 29612 1452 29668 1508
rect 29932 1452 29988 1508
rect 12 1292 68 1348
rect 332 1292 388 1348
rect 652 1292 708 1348
rect 972 1292 1028 1348
rect 28972 1292 29028 1348
rect 29292 1292 29348 1348
rect 29612 1292 29668 1348
rect 29932 1292 29988 1348
rect 12 1132 68 1188
rect 332 1132 388 1188
rect 652 1132 708 1188
rect 972 1132 1028 1188
rect 28972 1132 29028 1188
rect 29292 1132 29348 1188
rect 29612 1132 29668 1188
rect 29932 1132 29988 1188
rect 12 972 68 1028
rect 332 972 388 1028
rect 652 972 708 1028
rect 972 972 1028 1028
rect 1132 1026 1188 1028
rect 1132 974 1134 1026
rect 1134 974 1186 1026
rect 1186 974 1188 1026
rect 1132 972 1188 974
rect 28812 1026 28868 1028
rect 28812 974 28814 1026
rect 28814 974 28866 1026
rect 28866 974 28868 1026
rect 28812 972 28868 974
rect 28972 972 29028 1028
rect 29292 972 29348 1028
rect 29612 972 29668 1028
rect 29932 972 29988 1028
<< metal3 >>
rect 0 31912 80 31920
rect 0 31848 8 31912
rect 72 31848 80 31912
rect 0 31752 80 31848
rect 0 31688 8 31752
rect 72 31688 80 31752
rect 0 31592 80 31688
rect 0 31528 8 31592
rect 72 31528 80 31592
rect 0 31432 80 31528
rect 0 31368 8 31432
rect 72 31368 80 31432
rect 0 31272 80 31368
rect 0 31208 8 31272
rect 72 31208 80 31272
rect 0 31112 80 31208
rect 0 31048 8 31112
rect 72 31048 80 31112
rect 0 30952 80 31048
rect 0 30888 8 30952
rect 72 30888 80 30952
rect 0 30792 80 30888
rect 0 30728 8 30792
rect 72 30728 80 30792
rect 0 30632 80 30728
rect 0 30568 8 30632
rect 72 30568 80 30632
rect 0 30472 80 30568
rect 0 30408 8 30472
rect 72 30408 80 30472
rect 0 30312 80 30408
rect 0 30248 8 30312
rect 72 30248 80 30312
rect 0 30152 80 30248
rect 0 30088 8 30152
rect 72 30088 80 30152
rect 0 29992 80 30088
rect 0 29928 8 29992
rect 72 29928 80 29992
rect 0 29832 80 29928
rect 0 29768 8 29832
rect 72 29768 80 29832
rect 0 29672 80 29768
rect 0 29608 8 29672
rect 72 29608 80 29672
rect 0 29512 80 29608
rect 0 29448 8 29512
rect 72 29448 80 29512
rect 0 29352 80 29448
rect 0 29288 8 29352
rect 72 29288 80 29352
rect 0 29192 80 29288
rect 0 29128 8 29192
rect 72 29128 80 29192
rect 0 29032 80 29128
rect 0 28968 8 29032
rect 72 28968 80 29032
rect 0 28872 80 28968
rect 0 28808 8 28872
rect 72 28808 80 28872
rect 0 28712 80 28808
rect 0 28648 8 28712
rect 72 28648 80 28712
rect 0 28552 80 28648
rect 0 28488 8 28552
rect 72 28488 80 28552
rect 0 28392 80 28488
rect 0 28328 8 28392
rect 72 28328 80 28392
rect 0 28232 80 28328
rect 0 28168 8 28232
rect 72 28168 80 28232
rect 0 28072 80 28168
rect 0 28008 8 28072
rect 72 28008 80 28072
rect 0 27912 80 28008
rect 0 27848 8 27912
rect 72 27848 80 27912
rect 0 27752 80 27848
rect 0 27688 8 27752
rect 72 27688 80 27752
rect 0 27592 80 27688
rect 0 27528 8 27592
rect 72 27528 80 27592
rect 0 27432 80 27528
rect 0 27368 8 27432
rect 72 27368 80 27432
rect 0 27272 80 27368
rect 0 27208 8 27272
rect 72 27208 80 27272
rect 0 27112 80 27208
rect 0 27048 8 27112
rect 72 27048 80 27112
rect 0 26952 80 27048
rect 0 26888 8 26952
rect 72 26888 80 26952
rect 0 26792 80 26888
rect 0 26728 8 26792
rect 72 26728 80 26792
rect 0 26632 80 26728
rect 0 26568 8 26632
rect 72 26568 80 26632
rect 0 26472 80 26568
rect 0 26408 8 26472
rect 72 26408 80 26472
rect 0 26312 80 26408
rect 0 26248 8 26312
rect 72 26248 80 26312
rect 0 26152 80 26248
rect 0 26088 8 26152
rect 72 26088 80 26152
rect 0 25992 80 26088
rect 0 25928 8 25992
rect 72 25928 80 25992
rect 0 25832 80 25928
rect 0 25768 8 25832
rect 72 25768 80 25832
rect 0 25672 80 25768
rect 0 25608 8 25672
rect 72 25608 80 25672
rect 0 25512 80 25608
rect 0 25448 8 25512
rect 72 25448 80 25512
rect 0 25352 80 25448
rect 0 25288 8 25352
rect 72 25288 80 25352
rect 0 25192 80 25288
rect 0 25128 8 25192
rect 72 25128 80 25192
rect 0 25032 80 25128
rect 0 24968 8 25032
rect 72 24968 80 25032
rect 0 24872 80 24968
rect 0 24808 8 24872
rect 72 24808 80 24872
rect 0 24712 80 24808
rect 0 24648 8 24712
rect 72 24648 80 24712
rect 0 24552 80 24648
rect 0 24488 8 24552
rect 72 24488 80 24552
rect 0 24392 80 24488
rect 0 24328 8 24392
rect 72 24328 80 24392
rect 0 24232 80 24328
rect 0 24168 8 24232
rect 72 24168 80 24232
rect 0 24072 80 24168
rect 0 24008 8 24072
rect 72 24008 80 24072
rect 0 23912 80 24008
rect 0 23848 8 23912
rect 72 23848 80 23912
rect 0 23752 80 23848
rect 0 23688 8 23752
rect 72 23688 80 23752
rect 0 23592 80 23688
rect 0 23528 8 23592
rect 72 23528 80 23592
rect 0 23432 80 23528
rect 0 23368 8 23432
rect 72 23368 80 23432
rect 0 23272 80 23368
rect 0 23208 8 23272
rect 72 23208 80 23272
rect 0 23112 80 23208
rect 0 23048 8 23112
rect 72 23048 80 23112
rect 0 22952 80 23048
rect 0 22888 8 22952
rect 72 22888 80 22952
rect 0 22792 80 22888
rect 0 22728 8 22792
rect 72 22728 80 22792
rect 0 22472 80 22728
rect 0 22408 8 22472
rect 72 22408 80 22472
rect 0 22312 80 22408
rect 0 22248 8 22312
rect 72 22248 80 22312
rect 0 22152 80 22248
rect 0 22088 8 22152
rect 72 22088 80 22152
rect 0 21992 80 22088
rect 0 21928 8 21992
rect 72 21928 80 21992
rect 0 21832 80 21928
rect 0 21768 8 21832
rect 72 21768 80 21832
rect 0 21672 80 21768
rect 0 21608 8 21672
rect 72 21608 80 21672
rect 0 21512 80 21608
rect 0 21448 8 21512
rect 72 21448 80 21512
rect 0 21352 80 21448
rect 0 21288 8 21352
rect 72 21288 80 21352
rect 0 21192 80 21288
rect 0 21128 8 21192
rect 72 21128 80 21192
rect 0 21032 80 21128
rect 0 20968 8 21032
rect 72 20968 80 21032
rect 0 20872 80 20968
rect 0 20808 8 20872
rect 72 20808 80 20872
rect 0 20712 80 20808
rect 0 20648 8 20712
rect 72 20648 80 20712
rect 0 20552 80 20648
rect 0 20488 8 20552
rect 72 20488 80 20552
rect 0 20392 80 20488
rect 0 20328 8 20392
rect 72 20328 80 20392
rect 0 20232 80 20328
rect 0 20168 8 20232
rect 72 20168 80 20232
rect 0 20072 80 20168
rect 0 20008 8 20072
rect 72 20008 80 20072
rect 0 19912 80 20008
rect 0 19848 8 19912
rect 72 19848 80 19912
rect 0 19752 80 19848
rect 0 19688 8 19752
rect 72 19688 80 19752
rect 0 19592 80 19688
rect 0 19528 8 19592
rect 72 19528 80 19592
rect 0 19432 80 19528
rect 0 19368 8 19432
rect 72 19368 80 19432
rect 0 19272 80 19368
rect 0 19208 8 19272
rect 72 19208 80 19272
rect 0 19112 80 19208
rect 0 19048 8 19112
rect 72 19048 80 19112
rect 0 18952 80 19048
rect 0 18888 8 18952
rect 72 18888 80 18952
rect 0 18792 80 18888
rect 0 18728 8 18792
rect 72 18728 80 18792
rect 0 18632 80 18728
rect 0 18568 8 18632
rect 72 18568 80 18632
rect 0 18472 80 18568
rect 0 18408 8 18472
rect 72 18408 80 18472
rect 0 18312 80 18408
rect 0 18248 8 18312
rect 72 18248 80 18312
rect 0 18152 80 18248
rect 0 18088 8 18152
rect 72 18088 80 18152
rect 0 17992 80 18088
rect 0 17928 8 17992
rect 72 17928 80 17992
rect 0 17832 80 17928
rect 0 17768 8 17832
rect 72 17768 80 17832
rect 0 17672 80 17768
rect 0 17608 8 17672
rect 72 17608 80 17672
rect 0 17512 80 17608
rect 0 17448 8 17512
rect 72 17448 80 17512
rect 0 17352 80 17448
rect 0 17288 8 17352
rect 72 17288 80 17352
rect 0 17192 80 17288
rect 0 17128 8 17192
rect 72 17128 80 17192
rect 0 17032 80 17128
rect 0 16968 8 17032
rect 72 16968 80 17032
rect 0 16712 80 16968
rect 0 16648 8 16712
rect 72 16648 80 16712
rect 0 16552 80 16648
rect 0 16488 8 16552
rect 72 16488 80 16552
rect 0 16392 80 16488
rect 0 16328 8 16392
rect 72 16328 80 16392
rect 0 16232 80 16328
rect 0 16168 8 16232
rect 72 16168 80 16232
rect 0 15912 80 16168
rect 0 15848 8 15912
rect 72 15848 80 15912
rect 0 15752 80 15848
rect 0 15688 8 15752
rect 72 15688 80 15752
rect 0 15592 80 15688
rect 0 15528 8 15592
rect 72 15528 80 15592
rect 0 15432 80 15528
rect 0 15368 8 15432
rect 72 15368 80 15432
rect 0 15272 80 15368
rect 0 15208 8 15272
rect 72 15208 80 15272
rect 0 15112 80 15208
rect 0 15048 8 15112
rect 72 15048 80 15112
rect 0 14952 80 15048
rect 0 14888 8 14952
rect 72 14888 80 14952
rect 0 14792 80 14888
rect 0 14728 8 14792
rect 72 14728 80 14792
rect 0 14632 80 14728
rect 0 14568 8 14632
rect 72 14568 80 14632
rect 0 14472 80 14568
rect 0 14408 8 14472
rect 72 14408 80 14472
rect 0 14312 80 14408
rect 0 14248 8 14312
rect 72 14248 80 14312
rect 0 14152 80 14248
rect 0 14088 8 14152
rect 72 14088 80 14152
rect 0 13992 80 14088
rect 0 13928 8 13992
rect 72 13928 80 13992
rect 0 13832 80 13928
rect 0 13768 8 13832
rect 72 13768 80 13832
rect 0 13672 80 13768
rect 0 13608 8 13672
rect 72 13608 80 13672
rect 0 13512 80 13608
rect 0 13448 8 13512
rect 72 13448 80 13512
rect 0 13352 80 13448
rect 0 13288 8 13352
rect 72 13288 80 13352
rect 0 13192 80 13288
rect 0 13128 8 13192
rect 72 13128 80 13192
rect 0 13032 80 13128
rect 0 12968 8 13032
rect 72 12968 80 13032
rect 0 12872 80 12968
rect 0 12808 8 12872
rect 72 12808 80 12872
rect 0 12712 80 12808
rect 0 12648 8 12712
rect 72 12648 80 12712
rect 0 12552 80 12648
rect 0 12488 8 12552
rect 72 12488 80 12552
rect 0 12392 80 12488
rect 0 12328 8 12392
rect 72 12328 80 12392
rect 0 12232 80 12328
rect 0 12168 8 12232
rect 72 12168 80 12232
rect 0 12072 80 12168
rect 0 12008 8 12072
rect 72 12008 80 12072
rect 0 11912 80 12008
rect 0 11848 8 11912
rect 72 11848 80 11912
rect 0 11752 80 11848
rect 0 11688 8 11752
rect 72 11688 80 11752
rect 0 11592 80 11688
rect 0 11528 8 11592
rect 72 11528 80 11592
rect 0 11432 80 11528
rect 0 11368 8 11432
rect 72 11368 80 11432
rect 0 11272 80 11368
rect 0 11208 8 11272
rect 72 11208 80 11272
rect 0 11112 80 11208
rect 0 11048 8 11112
rect 72 11048 80 11112
rect 0 10952 80 11048
rect 0 10888 8 10952
rect 72 10888 80 10952
rect 0 10792 80 10888
rect 0 10728 8 10792
rect 72 10728 80 10792
rect 0 10632 80 10728
rect 0 10568 8 10632
rect 72 10568 80 10632
rect 0 10472 80 10568
rect 0 10408 8 10472
rect 72 10408 80 10472
rect 0 10152 80 10408
rect 0 10088 8 10152
rect 72 10088 80 10152
rect 0 9992 80 10088
rect 0 9928 8 9992
rect 72 9928 80 9992
rect 0 9832 80 9928
rect 0 9768 8 9832
rect 72 9768 80 9832
rect 0 9672 80 9768
rect 0 9608 8 9672
rect 72 9608 80 9672
rect 0 9512 80 9608
rect 0 9448 8 9512
rect 72 9448 80 9512
rect 0 9352 80 9448
rect 0 9288 8 9352
rect 72 9288 80 9352
rect 0 9192 80 9288
rect 0 9128 8 9192
rect 72 9128 80 9192
rect 0 9032 80 9128
rect 0 8968 8 9032
rect 72 8968 80 9032
rect 0 8872 80 8968
rect 0 8808 8 8872
rect 72 8808 80 8872
rect 0 8712 80 8808
rect 0 8648 8 8712
rect 72 8648 80 8712
rect 0 8552 80 8648
rect 0 8488 8 8552
rect 72 8488 80 8552
rect 0 8392 80 8488
rect 0 8328 8 8392
rect 72 8328 80 8392
rect 0 8232 80 8328
rect 0 8168 8 8232
rect 72 8168 80 8232
rect 0 8072 80 8168
rect 0 8008 8 8072
rect 72 8008 80 8072
rect 0 7912 80 8008
rect 0 7848 8 7912
rect 72 7848 80 7912
rect 0 7752 80 7848
rect 0 7688 8 7752
rect 72 7688 80 7752
rect 0 7592 80 7688
rect 0 7528 8 7592
rect 72 7528 80 7592
rect 0 7432 80 7528
rect 0 7368 8 7432
rect 72 7368 80 7432
rect 0 7272 80 7368
rect 0 7208 8 7272
rect 72 7208 80 7272
rect 0 7112 80 7208
rect 0 7048 8 7112
rect 72 7048 80 7112
rect 0 6952 80 7048
rect 0 6888 8 6952
rect 72 6888 80 6952
rect 0 6792 80 6888
rect 0 6728 8 6792
rect 72 6728 80 6792
rect 0 6632 80 6728
rect 0 6568 8 6632
rect 72 6568 80 6632
rect 0 6472 80 6568
rect 0 6408 8 6472
rect 72 6408 80 6472
rect 0 6312 80 6408
rect 0 6248 8 6312
rect 72 6248 80 6312
rect 0 6152 80 6248
rect 0 6088 8 6152
rect 72 6088 80 6152
rect 0 5992 80 6088
rect 0 5928 8 5992
rect 72 5928 80 5992
rect 0 5832 80 5928
rect 0 5768 8 5832
rect 72 5768 80 5832
rect 0 5672 80 5768
rect 0 5608 8 5672
rect 72 5608 80 5672
rect 0 5512 80 5608
rect 0 5448 8 5512
rect 72 5448 80 5512
rect 0 5352 80 5448
rect 0 5288 8 5352
rect 72 5288 80 5352
rect 0 5192 80 5288
rect 0 5128 8 5192
rect 72 5128 80 5192
rect 0 5032 80 5128
rect 0 4968 8 5032
rect 72 4968 80 5032
rect 0 4872 80 4968
rect 0 4808 8 4872
rect 72 4808 80 4872
rect 0 4712 80 4808
rect 0 4648 8 4712
rect 72 4648 80 4712
rect 0 4552 80 4648
rect 0 4488 8 4552
rect 72 4488 80 4552
rect 0 4392 80 4488
rect 0 4328 8 4392
rect 72 4328 80 4392
rect 0 4232 80 4328
rect 0 4168 8 4232
rect 72 4168 80 4232
rect 0 4072 80 4168
rect 0 4008 8 4072
rect 72 4008 80 4072
rect 0 3912 80 4008
rect 0 3848 8 3912
rect 72 3848 80 3912
rect 0 3752 80 3848
rect 0 3688 8 3752
rect 72 3688 80 3752
rect 0 3592 80 3688
rect 0 3528 8 3592
rect 72 3528 80 3592
rect 0 3432 80 3528
rect 0 3368 8 3432
rect 72 3368 80 3432
rect 0 3272 80 3368
rect 0 3208 8 3272
rect 72 3208 80 3272
rect 0 3112 80 3208
rect 0 3048 8 3112
rect 72 3048 80 3112
rect 0 2952 80 3048
rect 0 2888 8 2952
rect 72 2888 80 2952
rect 0 2792 80 2888
rect 0 2728 8 2792
rect 72 2728 80 2792
rect 0 2632 80 2728
rect 0 2568 8 2632
rect 72 2568 80 2632
rect 0 2472 80 2568
rect 0 2408 8 2472
rect 72 2408 80 2472
rect 0 2312 80 2408
rect 0 2248 8 2312
rect 72 2248 80 2312
rect 0 2152 80 2248
rect 0 2088 8 2152
rect 72 2088 80 2152
rect 0 1992 80 2088
rect 0 1928 8 1992
rect 72 1928 80 1992
rect 0 1832 80 1928
rect 0 1768 8 1832
rect 72 1768 80 1832
rect 0 1672 80 1768
rect 0 1608 8 1672
rect 72 1608 80 1672
rect 0 1512 80 1608
rect 0 1448 8 1512
rect 72 1448 80 1512
rect 0 1352 80 1448
rect 0 1288 8 1352
rect 72 1288 80 1352
rect 0 1192 80 1288
rect 0 1128 8 1192
rect 72 1128 80 1192
rect 0 1032 80 1128
rect 0 968 8 1032
rect 72 968 80 1032
rect 0 872 80 968
rect 160 22632 240 31920
rect 160 22568 168 22632
rect 232 22568 240 22632
rect 160 16872 240 22568
rect 160 16808 168 16872
rect 232 16808 240 16872
rect 160 16072 240 16808
rect 160 16008 168 16072
rect 232 16008 240 16072
rect 160 10312 240 16008
rect 160 10248 168 10312
rect 232 10248 240 10312
rect 160 960 240 10248
rect 320 31912 400 31920
rect 320 31848 328 31912
rect 392 31848 400 31912
rect 320 31752 400 31848
rect 320 31688 328 31752
rect 392 31688 400 31752
rect 320 31592 400 31688
rect 320 31528 328 31592
rect 392 31528 400 31592
rect 320 31432 400 31528
rect 320 31368 328 31432
rect 392 31368 400 31432
rect 320 31272 400 31368
rect 320 31208 328 31272
rect 392 31208 400 31272
rect 320 31112 400 31208
rect 320 31048 328 31112
rect 392 31048 400 31112
rect 320 30952 400 31048
rect 320 30888 328 30952
rect 392 30888 400 30952
rect 320 30792 400 30888
rect 320 30728 328 30792
rect 392 30728 400 30792
rect 320 30632 400 30728
rect 320 30568 328 30632
rect 392 30568 400 30632
rect 320 30472 400 30568
rect 320 30408 328 30472
rect 392 30408 400 30472
rect 320 30312 400 30408
rect 320 30248 328 30312
rect 392 30248 400 30312
rect 320 30152 400 30248
rect 320 30088 328 30152
rect 392 30088 400 30152
rect 320 29992 400 30088
rect 320 29928 328 29992
rect 392 29928 400 29992
rect 320 29832 400 29928
rect 320 29768 328 29832
rect 392 29768 400 29832
rect 320 29672 400 29768
rect 320 29608 328 29672
rect 392 29608 400 29672
rect 320 29512 400 29608
rect 320 29448 328 29512
rect 392 29448 400 29512
rect 320 29352 400 29448
rect 320 29288 328 29352
rect 392 29288 400 29352
rect 320 29192 400 29288
rect 320 29128 328 29192
rect 392 29128 400 29192
rect 320 29032 400 29128
rect 320 28968 328 29032
rect 392 28968 400 29032
rect 320 28872 400 28968
rect 320 28808 328 28872
rect 392 28808 400 28872
rect 320 28712 400 28808
rect 320 28648 328 28712
rect 392 28648 400 28712
rect 320 28552 400 28648
rect 320 28488 328 28552
rect 392 28488 400 28552
rect 320 28392 400 28488
rect 320 28328 328 28392
rect 392 28328 400 28392
rect 320 28232 400 28328
rect 320 28168 328 28232
rect 392 28168 400 28232
rect 320 28072 400 28168
rect 320 28008 328 28072
rect 392 28008 400 28072
rect 320 27912 400 28008
rect 320 27848 328 27912
rect 392 27848 400 27912
rect 320 27752 400 27848
rect 320 27688 328 27752
rect 392 27688 400 27752
rect 320 27592 400 27688
rect 320 27528 328 27592
rect 392 27528 400 27592
rect 320 27432 400 27528
rect 320 27368 328 27432
rect 392 27368 400 27432
rect 320 27272 400 27368
rect 320 27208 328 27272
rect 392 27208 400 27272
rect 320 27112 400 27208
rect 320 27048 328 27112
rect 392 27048 400 27112
rect 320 26952 400 27048
rect 320 26888 328 26952
rect 392 26888 400 26952
rect 320 26792 400 26888
rect 320 26728 328 26792
rect 392 26728 400 26792
rect 320 26632 400 26728
rect 320 26568 328 26632
rect 392 26568 400 26632
rect 320 26472 400 26568
rect 320 26408 328 26472
rect 392 26408 400 26472
rect 320 26312 400 26408
rect 320 26248 328 26312
rect 392 26248 400 26312
rect 320 26152 400 26248
rect 320 26088 328 26152
rect 392 26088 400 26152
rect 320 25992 400 26088
rect 320 25928 328 25992
rect 392 25928 400 25992
rect 320 25832 400 25928
rect 320 25768 328 25832
rect 392 25768 400 25832
rect 320 25672 400 25768
rect 320 25608 328 25672
rect 392 25608 400 25672
rect 320 25512 400 25608
rect 320 25448 328 25512
rect 392 25448 400 25512
rect 320 25352 400 25448
rect 320 25288 328 25352
rect 392 25288 400 25352
rect 320 25192 400 25288
rect 320 25128 328 25192
rect 392 25128 400 25192
rect 320 25032 400 25128
rect 320 24968 328 25032
rect 392 24968 400 25032
rect 320 24872 400 24968
rect 320 24808 328 24872
rect 392 24808 400 24872
rect 320 24712 400 24808
rect 320 24648 328 24712
rect 392 24648 400 24712
rect 320 24552 400 24648
rect 320 24488 328 24552
rect 392 24488 400 24552
rect 320 24392 400 24488
rect 320 24328 328 24392
rect 392 24328 400 24392
rect 320 24232 400 24328
rect 320 24168 328 24232
rect 392 24168 400 24232
rect 320 24072 400 24168
rect 320 24008 328 24072
rect 392 24008 400 24072
rect 320 23912 400 24008
rect 320 23848 328 23912
rect 392 23848 400 23912
rect 320 23752 400 23848
rect 320 23688 328 23752
rect 392 23688 400 23752
rect 320 23592 400 23688
rect 320 23528 328 23592
rect 392 23528 400 23592
rect 320 23432 400 23528
rect 320 23368 328 23432
rect 392 23368 400 23432
rect 320 23272 400 23368
rect 320 23208 328 23272
rect 392 23208 400 23272
rect 320 23112 400 23208
rect 320 23048 328 23112
rect 392 23048 400 23112
rect 320 22952 400 23048
rect 320 22888 328 22952
rect 392 22888 400 22952
rect 320 22792 400 22888
rect 320 22728 328 22792
rect 392 22728 400 22792
rect 320 22472 400 22728
rect 320 22408 328 22472
rect 392 22408 400 22472
rect 320 22312 400 22408
rect 320 22248 328 22312
rect 392 22248 400 22312
rect 320 22152 400 22248
rect 320 22088 328 22152
rect 392 22088 400 22152
rect 320 21992 400 22088
rect 320 21928 328 21992
rect 392 21928 400 21992
rect 320 21832 400 21928
rect 320 21768 328 21832
rect 392 21768 400 21832
rect 320 21672 400 21768
rect 320 21608 328 21672
rect 392 21608 400 21672
rect 320 21512 400 21608
rect 320 21448 328 21512
rect 392 21448 400 21512
rect 320 21352 400 21448
rect 320 21288 328 21352
rect 392 21288 400 21352
rect 320 21192 400 21288
rect 320 21128 328 21192
rect 392 21128 400 21192
rect 320 21032 400 21128
rect 320 20968 328 21032
rect 392 20968 400 21032
rect 320 20872 400 20968
rect 320 20808 328 20872
rect 392 20808 400 20872
rect 320 20712 400 20808
rect 320 20648 328 20712
rect 392 20648 400 20712
rect 320 20552 400 20648
rect 320 20488 328 20552
rect 392 20488 400 20552
rect 320 20392 400 20488
rect 320 20328 328 20392
rect 392 20328 400 20392
rect 320 20232 400 20328
rect 320 20168 328 20232
rect 392 20168 400 20232
rect 320 20072 400 20168
rect 320 20008 328 20072
rect 392 20008 400 20072
rect 320 19912 400 20008
rect 320 19848 328 19912
rect 392 19848 400 19912
rect 320 19752 400 19848
rect 320 19688 328 19752
rect 392 19688 400 19752
rect 320 19592 400 19688
rect 320 19528 328 19592
rect 392 19528 400 19592
rect 320 19432 400 19528
rect 320 19368 328 19432
rect 392 19368 400 19432
rect 320 19272 400 19368
rect 320 19208 328 19272
rect 392 19208 400 19272
rect 320 19112 400 19208
rect 320 19048 328 19112
rect 392 19048 400 19112
rect 320 18952 400 19048
rect 320 18888 328 18952
rect 392 18888 400 18952
rect 320 18792 400 18888
rect 320 18728 328 18792
rect 392 18728 400 18792
rect 320 18632 400 18728
rect 320 18568 328 18632
rect 392 18568 400 18632
rect 320 18472 400 18568
rect 320 18408 328 18472
rect 392 18408 400 18472
rect 320 18312 400 18408
rect 320 18248 328 18312
rect 392 18248 400 18312
rect 320 18152 400 18248
rect 320 18088 328 18152
rect 392 18088 400 18152
rect 320 17992 400 18088
rect 320 17928 328 17992
rect 392 17928 400 17992
rect 320 17832 400 17928
rect 320 17768 328 17832
rect 392 17768 400 17832
rect 320 17672 400 17768
rect 320 17608 328 17672
rect 392 17608 400 17672
rect 320 17512 400 17608
rect 320 17448 328 17512
rect 392 17448 400 17512
rect 320 17352 400 17448
rect 320 17288 328 17352
rect 392 17288 400 17352
rect 320 17192 400 17288
rect 320 17128 328 17192
rect 392 17128 400 17192
rect 320 17032 400 17128
rect 320 16968 328 17032
rect 392 16968 400 17032
rect 320 16712 400 16968
rect 320 16648 328 16712
rect 392 16648 400 16712
rect 320 16552 400 16648
rect 320 16488 328 16552
rect 392 16488 400 16552
rect 320 16392 400 16488
rect 320 16328 328 16392
rect 392 16328 400 16392
rect 320 16232 400 16328
rect 320 16168 328 16232
rect 392 16168 400 16232
rect 320 15912 400 16168
rect 320 15848 328 15912
rect 392 15848 400 15912
rect 320 15752 400 15848
rect 320 15688 328 15752
rect 392 15688 400 15752
rect 320 15592 400 15688
rect 320 15528 328 15592
rect 392 15528 400 15592
rect 320 15432 400 15528
rect 320 15368 328 15432
rect 392 15368 400 15432
rect 320 15272 400 15368
rect 320 15208 328 15272
rect 392 15208 400 15272
rect 320 15112 400 15208
rect 320 15048 328 15112
rect 392 15048 400 15112
rect 320 14952 400 15048
rect 320 14888 328 14952
rect 392 14888 400 14952
rect 320 14792 400 14888
rect 320 14728 328 14792
rect 392 14728 400 14792
rect 320 14632 400 14728
rect 320 14568 328 14632
rect 392 14568 400 14632
rect 320 14472 400 14568
rect 320 14408 328 14472
rect 392 14408 400 14472
rect 320 14312 400 14408
rect 320 14248 328 14312
rect 392 14248 400 14312
rect 320 14152 400 14248
rect 320 14088 328 14152
rect 392 14088 400 14152
rect 320 13992 400 14088
rect 320 13928 328 13992
rect 392 13928 400 13992
rect 320 13832 400 13928
rect 320 13768 328 13832
rect 392 13768 400 13832
rect 320 13672 400 13768
rect 320 13608 328 13672
rect 392 13608 400 13672
rect 320 13512 400 13608
rect 320 13448 328 13512
rect 392 13448 400 13512
rect 320 13352 400 13448
rect 320 13288 328 13352
rect 392 13288 400 13352
rect 320 13192 400 13288
rect 320 13128 328 13192
rect 392 13128 400 13192
rect 320 13032 400 13128
rect 320 12968 328 13032
rect 392 12968 400 13032
rect 320 12872 400 12968
rect 320 12808 328 12872
rect 392 12808 400 12872
rect 320 12712 400 12808
rect 320 12648 328 12712
rect 392 12648 400 12712
rect 320 12552 400 12648
rect 320 12488 328 12552
rect 392 12488 400 12552
rect 320 12392 400 12488
rect 320 12328 328 12392
rect 392 12328 400 12392
rect 320 12232 400 12328
rect 320 12168 328 12232
rect 392 12168 400 12232
rect 320 12072 400 12168
rect 320 12008 328 12072
rect 392 12008 400 12072
rect 320 11912 400 12008
rect 320 11848 328 11912
rect 392 11848 400 11912
rect 320 11752 400 11848
rect 320 11688 328 11752
rect 392 11688 400 11752
rect 320 11592 400 11688
rect 320 11528 328 11592
rect 392 11528 400 11592
rect 320 11432 400 11528
rect 320 11368 328 11432
rect 392 11368 400 11432
rect 320 11272 400 11368
rect 320 11208 328 11272
rect 392 11208 400 11272
rect 320 11112 400 11208
rect 320 11048 328 11112
rect 392 11048 400 11112
rect 320 10952 400 11048
rect 320 10888 328 10952
rect 392 10888 400 10952
rect 320 10792 400 10888
rect 320 10728 328 10792
rect 392 10728 400 10792
rect 320 10632 400 10728
rect 320 10568 328 10632
rect 392 10568 400 10632
rect 320 10472 400 10568
rect 320 10408 328 10472
rect 392 10408 400 10472
rect 320 10152 400 10408
rect 320 10088 328 10152
rect 392 10088 400 10152
rect 320 9992 400 10088
rect 320 9928 328 9992
rect 392 9928 400 9992
rect 320 9832 400 9928
rect 320 9768 328 9832
rect 392 9768 400 9832
rect 320 9672 400 9768
rect 320 9608 328 9672
rect 392 9608 400 9672
rect 320 9512 400 9608
rect 320 9448 328 9512
rect 392 9448 400 9512
rect 320 9352 400 9448
rect 320 9288 328 9352
rect 392 9288 400 9352
rect 320 9192 400 9288
rect 320 9128 328 9192
rect 392 9128 400 9192
rect 320 9032 400 9128
rect 320 8968 328 9032
rect 392 8968 400 9032
rect 320 8872 400 8968
rect 320 8808 328 8872
rect 392 8808 400 8872
rect 320 8712 400 8808
rect 320 8648 328 8712
rect 392 8648 400 8712
rect 320 8552 400 8648
rect 320 8488 328 8552
rect 392 8488 400 8552
rect 320 8392 400 8488
rect 320 8328 328 8392
rect 392 8328 400 8392
rect 320 8232 400 8328
rect 320 8168 328 8232
rect 392 8168 400 8232
rect 320 8072 400 8168
rect 320 8008 328 8072
rect 392 8008 400 8072
rect 320 7912 400 8008
rect 320 7848 328 7912
rect 392 7848 400 7912
rect 320 7752 400 7848
rect 320 7688 328 7752
rect 392 7688 400 7752
rect 320 7592 400 7688
rect 320 7528 328 7592
rect 392 7528 400 7592
rect 320 7432 400 7528
rect 320 7368 328 7432
rect 392 7368 400 7432
rect 320 7272 400 7368
rect 320 7208 328 7272
rect 392 7208 400 7272
rect 320 7112 400 7208
rect 320 7048 328 7112
rect 392 7048 400 7112
rect 320 6952 400 7048
rect 320 6888 328 6952
rect 392 6888 400 6952
rect 320 6792 400 6888
rect 320 6728 328 6792
rect 392 6728 400 6792
rect 320 6632 400 6728
rect 320 6568 328 6632
rect 392 6568 400 6632
rect 320 6472 400 6568
rect 320 6408 328 6472
rect 392 6408 400 6472
rect 320 6312 400 6408
rect 320 6248 328 6312
rect 392 6248 400 6312
rect 320 6152 400 6248
rect 320 6088 328 6152
rect 392 6088 400 6152
rect 320 5992 400 6088
rect 320 5928 328 5992
rect 392 5928 400 5992
rect 320 5832 400 5928
rect 320 5768 328 5832
rect 392 5768 400 5832
rect 320 5672 400 5768
rect 320 5608 328 5672
rect 392 5608 400 5672
rect 320 5512 400 5608
rect 320 5448 328 5512
rect 392 5448 400 5512
rect 320 5352 400 5448
rect 320 5288 328 5352
rect 392 5288 400 5352
rect 320 5192 400 5288
rect 320 5128 328 5192
rect 392 5128 400 5192
rect 320 5032 400 5128
rect 320 4968 328 5032
rect 392 4968 400 5032
rect 320 4872 400 4968
rect 320 4808 328 4872
rect 392 4808 400 4872
rect 320 4712 400 4808
rect 320 4648 328 4712
rect 392 4648 400 4712
rect 320 4552 400 4648
rect 320 4488 328 4552
rect 392 4488 400 4552
rect 320 4392 400 4488
rect 320 4328 328 4392
rect 392 4328 400 4392
rect 320 4232 400 4328
rect 320 4168 328 4232
rect 392 4168 400 4232
rect 320 4072 400 4168
rect 320 4008 328 4072
rect 392 4008 400 4072
rect 320 3912 400 4008
rect 320 3848 328 3912
rect 392 3848 400 3912
rect 320 3752 400 3848
rect 320 3688 328 3752
rect 392 3688 400 3752
rect 320 3592 400 3688
rect 320 3528 328 3592
rect 392 3528 400 3592
rect 320 3432 400 3528
rect 320 3368 328 3432
rect 392 3368 400 3432
rect 320 3272 400 3368
rect 320 3208 328 3272
rect 392 3208 400 3272
rect 320 3112 400 3208
rect 320 3048 328 3112
rect 392 3048 400 3112
rect 320 2952 400 3048
rect 320 2888 328 2952
rect 392 2888 400 2952
rect 320 2792 400 2888
rect 320 2728 328 2792
rect 392 2728 400 2792
rect 320 2632 400 2728
rect 320 2568 328 2632
rect 392 2568 400 2632
rect 320 2472 400 2568
rect 320 2408 328 2472
rect 392 2408 400 2472
rect 320 2312 400 2408
rect 320 2248 328 2312
rect 392 2248 400 2312
rect 320 2152 400 2248
rect 320 2088 328 2152
rect 392 2088 400 2152
rect 320 1992 400 2088
rect 320 1928 328 1992
rect 392 1928 400 1992
rect 320 1832 400 1928
rect 320 1768 328 1832
rect 392 1768 400 1832
rect 320 1672 400 1768
rect 320 1608 328 1672
rect 392 1608 400 1672
rect 320 1512 400 1608
rect 320 1448 328 1512
rect 392 1448 400 1512
rect 320 1352 400 1448
rect 320 1288 328 1352
rect 392 1288 400 1352
rect 320 1192 400 1288
rect 320 1128 328 1192
rect 392 1128 400 1192
rect 320 1032 400 1128
rect 320 968 328 1032
rect 392 968 400 1032
rect 0 808 8 872
rect 72 808 80 872
rect 0 792 80 808
rect 0 728 8 792
rect 72 728 80 792
rect 0 712 80 728
rect 0 648 8 712
rect 72 648 80 712
rect 0 632 80 648
rect 0 568 8 632
rect 72 568 80 632
rect 0 552 80 568
rect 0 488 8 552
rect 72 488 80 552
rect 0 480 80 488
rect 320 872 400 968
rect 480 22312 560 31920
rect 480 22248 488 22312
rect 552 22248 560 22312
rect 480 17192 560 22248
rect 480 17128 488 17192
rect 552 17128 560 17192
rect 480 15752 560 17128
rect 480 15688 488 15752
rect 552 15688 560 15752
rect 480 10632 560 15688
rect 480 10568 488 10632
rect 552 10568 560 10632
rect 480 960 560 10568
rect 640 31912 720 31920
rect 640 31848 648 31912
rect 712 31848 720 31912
rect 640 31752 720 31848
rect 640 31688 648 31752
rect 712 31688 720 31752
rect 640 31592 720 31688
rect 640 31528 648 31592
rect 712 31528 720 31592
rect 640 31432 720 31528
rect 640 31368 648 31432
rect 712 31368 720 31432
rect 640 31272 720 31368
rect 640 31208 648 31272
rect 712 31208 720 31272
rect 640 31112 720 31208
rect 640 31048 648 31112
rect 712 31048 720 31112
rect 640 30952 720 31048
rect 640 30888 648 30952
rect 712 30888 720 30952
rect 640 30792 720 30888
rect 640 30728 648 30792
rect 712 30728 720 30792
rect 640 30632 720 30728
rect 640 30568 648 30632
rect 712 30568 720 30632
rect 640 30472 720 30568
rect 640 30408 648 30472
rect 712 30408 720 30472
rect 640 30312 720 30408
rect 640 30248 648 30312
rect 712 30248 720 30312
rect 640 30152 720 30248
rect 640 30088 648 30152
rect 712 30088 720 30152
rect 640 29992 720 30088
rect 640 29928 648 29992
rect 712 29928 720 29992
rect 640 29832 720 29928
rect 640 29768 648 29832
rect 712 29768 720 29832
rect 640 29672 720 29768
rect 640 29608 648 29672
rect 712 29608 720 29672
rect 640 29512 720 29608
rect 640 29448 648 29512
rect 712 29448 720 29512
rect 640 29352 720 29448
rect 640 29288 648 29352
rect 712 29288 720 29352
rect 640 29192 720 29288
rect 640 29128 648 29192
rect 712 29128 720 29192
rect 640 29032 720 29128
rect 640 28968 648 29032
rect 712 28968 720 29032
rect 640 28872 720 28968
rect 640 28808 648 28872
rect 712 28808 720 28872
rect 640 28712 720 28808
rect 640 28648 648 28712
rect 712 28648 720 28712
rect 640 28552 720 28648
rect 640 28488 648 28552
rect 712 28488 720 28552
rect 640 28392 720 28488
rect 640 28328 648 28392
rect 712 28328 720 28392
rect 640 28232 720 28328
rect 640 28168 648 28232
rect 712 28168 720 28232
rect 640 28072 720 28168
rect 640 28008 648 28072
rect 712 28008 720 28072
rect 640 27912 720 28008
rect 640 27848 648 27912
rect 712 27848 720 27912
rect 640 27752 720 27848
rect 640 27688 648 27752
rect 712 27688 720 27752
rect 640 27592 720 27688
rect 640 27528 648 27592
rect 712 27528 720 27592
rect 640 27432 720 27528
rect 640 27368 648 27432
rect 712 27368 720 27432
rect 640 27272 720 27368
rect 640 27208 648 27272
rect 712 27208 720 27272
rect 640 27112 720 27208
rect 640 27048 648 27112
rect 712 27048 720 27112
rect 640 26952 720 27048
rect 640 26888 648 26952
rect 712 26888 720 26952
rect 640 26792 720 26888
rect 640 26728 648 26792
rect 712 26728 720 26792
rect 640 26632 720 26728
rect 640 26568 648 26632
rect 712 26568 720 26632
rect 640 26472 720 26568
rect 640 26408 648 26472
rect 712 26408 720 26472
rect 640 26312 720 26408
rect 640 26248 648 26312
rect 712 26248 720 26312
rect 640 26152 720 26248
rect 640 26088 648 26152
rect 712 26088 720 26152
rect 640 25992 720 26088
rect 640 25928 648 25992
rect 712 25928 720 25992
rect 640 25832 720 25928
rect 640 25768 648 25832
rect 712 25768 720 25832
rect 640 25672 720 25768
rect 640 25608 648 25672
rect 712 25608 720 25672
rect 640 25512 720 25608
rect 640 25448 648 25512
rect 712 25448 720 25512
rect 640 25352 720 25448
rect 640 25288 648 25352
rect 712 25288 720 25352
rect 640 25192 720 25288
rect 640 25128 648 25192
rect 712 25128 720 25192
rect 640 25032 720 25128
rect 640 24968 648 25032
rect 712 24968 720 25032
rect 640 24872 720 24968
rect 640 24808 648 24872
rect 712 24808 720 24872
rect 640 24712 720 24808
rect 640 24648 648 24712
rect 712 24648 720 24712
rect 640 24552 720 24648
rect 640 24488 648 24552
rect 712 24488 720 24552
rect 640 24392 720 24488
rect 640 24328 648 24392
rect 712 24328 720 24392
rect 640 24232 720 24328
rect 640 24168 648 24232
rect 712 24168 720 24232
rect 640 24072 720 24168
rect 640 24008 648 24072
rect 712 24008 720 24072
rect 640 23912 720 24008
rect 640 23848 648 23912
rect 712 23848 720 23912
rect 640 23752 720 23848
rect 640 23688 648 23752
rect 712 23688 720 23752
rect 640 23592 720 23688
rect 640 23528 648 23592
rect 712 23528 720 23592
rect 640 23432 720 23528
rect 640 23368 648 23432
rect 712 23368 720 23432
rect 640 23272 720 23368
rect 640 23208 648 23272
rect 712 23208 720 23272
rect 640 23112 720 23208
rect 640 23048 648 23112
rect 712 23048 720 23112
rect 640 22952 720 23048
rect 640 22888 648 22952
rect 712 22888 720 22952
rect 640 22792 720 22888
rect 640 22728 648 22792
rect 712 22728 720 22792
rect 640 22472 720 22728
rect 640 22408 648 22472
rect 712 22408 720 22472
rect 640 22152 720 22408
rect 640 22088 648 22152
rect 712 22088 720 22152
rect 640 21992 720 22088
rect 640 21928 648 21992
rect 712 21928 720 21992
rect 640 21832 720 21928
rect 640 21768 648 21832
rect 712 21768 720 21832
rect 640 21672 720 21768
rect 640 21608 648 21672
rect 712 21608 720 21672
rect 640 21512 720 21608
rect 640 21448 648 21512
rect 712 21448 720 21512
rect 640 21352 720 21448
rect 640 21288 648 21352
rect 712 21288 720 21352
rect 640 21192 720 21288
rect 640 21128 648 21192
rect 712 21128 720 21192
rect 640 21032 720 21128
rect 640 20968 648 21032
rect 712 20968 720 21032
rect 640 20872 720 20968
rect 640 20808 648 20872
rect 712 20808 720 20872
rect 640 20712 720 20808
rect 640 20648 648 20712
rect 712 20648 720 20712
rect 640 20552 720 20648
rect 640 20488 648 20552
rect 712 20488 720 20552
rect 640 20392 720 20488
rect 640 20328 648 20392
rect 712 20328 720 20392
rect 640 20232 720 20328
rect 640 20168 648 20232
rect 712 20168 720 20232
rect 640 20072 720 20168
rect 640 20008 648 20072
rect 712 20008 720 20072
rect 640 19912 720 20008
rect 640 19848 648 19912
rect 712 19848 720 19912
rect 640 19752 720 19848
rect 640 19688 648 19752
rect 712 19688 720 19752
rect 640 19592 720 19688
rect 640 19528 648 19592
rect 712 19528 720 19592
rect 640 19432 720 19528
rect 640 19368 648 19432
rect 712 19368 720 19432
rect 640 19272 720 19368
rect 640 19208 648 19272
rect 712 19208 720 19272
rect 640 19112 720 19208
rect 640 19048 648 19112
rect 712 19048 720 19112
rect 640 18952 720 19048
rect 640 18888 648 18952
rect 712 18888 720 18952
rect 640 18792 720 18888
rect 640 18728 648 18792
rect 712 18728 720 18792
rect 640 18632 720 18728
rect 640 18568 648 18632
rect 712 18568 720 18632
rect 640 18472 720 18568
rect 640 18408 648 18472
rect 712 18408 720 18472
rect 640 18312 720 18408
rect 640 18248 648 18312
rect 712 18248 720 18312
rect 640 18152 720 18248
rect 640 18088 648 18152
rect 712 18088 720 18152
rect 640 17992 720 18088
rect 640 17928 648 17992
rect 712 17928 720 17992
rect 640 17832 720 17928
rect 640 17768 648 17832
rect 712 17768 720 17832
rect 640 17672 720 17768
rect 640 17608 648 17672
rect 712 17608 720 17672
rect 640 17512 720 17608
rect 640 17448 648 17512
rect 712 17448 720 17512
rect 640 17352 720 17448
rect 640 17288 648 17352
rect 712 17288 720 17352
rect 640 17032 720 17288
rect 640 16968 648 17032
rect 712 16968 720 17032
rect 640 16712 720 16968
rect 640 16648 648 16712
rect 712 16648 720 16712
rect 640 16552 720 16648
rect 640 16488 648 16552
rect 712 16488 720 16552
rect 640 16392 720 16488
rect 640 16328 648 16392
rect 712 16328 720 16392
rect 640 16232 720 16328
rect 640 16168 648 16232
rect 712 16168 720 16232
rect 640 15912 720 16168
rect 640 15848 648 15912
rect 712 15848 720 15912
rect 640 15592 720 15848
rect 640 15528 648 15592
rect 712 15528 720 15592
rect 640 15432 720 15528
rect 640 15368 648 15432
rect 712 15368 720 15432
rect 640 15272 720 15368
rect 640 15208 648 15272
rect 712 15208 720 15272
rect 640 15112 720 15208
rect 640 15048 648 15112
rect 712 15048 720 15112
rect 640 14952 720 15048
rect 640 14888 648 14952
rect 712 14888 720 14952
rect 640 14792 720 14888
rect 640 14728 648 14792
rect 712 14728 720 14792
rect 640 14632 720 14728
rect 640 14568 648 14632
rect 712 14568 720 14632
rect 640 14472 720 14568
rect 640 14408 648 14472
rect 712 14408 720 14472
rect 640 14312 720 14408
rect 640 14248 648 14312
rect 712 14248 720 14312
rect 640 14152 720 14248
rect 640 14088 648 14152
rect 712 14088 720 14152
rect 640 13992 720 14088
rect 640 13928 648 13992
rect 712 13928 720 13992
rect 640 13832 720 13928
rect 640 13768 648 13832
rect 712 13768 720 13832
rect 640 13672 720 13768
rect 640 13608 648 13672
rect 712 13608 720 13672
rect 640 13512 720 13608
rect 640 13448 648 13512
rect 712 13448 720 13512
rect 640 13352 720 13448
rect 640 13288 648 13352
rect 712 13288 720 13352
rect 640 13192 720 13288
rect 640 13128 648 13192
rect 712 13128 720 13192
rect 640 13032 720 13128
rect 640 12968 648 13032
rect 712 12968 720 13032
rect 640 12872 720 12968
rect 640 12808 648 12872
rect 712 12808 720 12872
rect 640 12712 720 12808
rect 640 12648 648 12712
rect 712 12648 720 12712
rect 640 12552 720 12648
rect 640 12488 648 12552
rect 712 12488 720 12552
rect 640 12392 720 12488
rect 640 12328 648 12392
rect 712 12328 720 12392
rect 640 12232 720 12328
rect 640 12168 648 12232
rect 712 12168 720 12232
rect 640 12072 720 12168
rect 640 12008 648 12072
rect 712 12008 720 12072
rect 640 11912 720 12008
rect 640 11848 648 11912
rect 712 11848 720 11912
rect 640 11752 720 11848
rect 640 11688 648 11752
rect 712 11688 720 11752
rect 640 11592 720 11688
rect 640 11528 648 11592
rect 712 11528 720 11592
rect 640 11432 720 11528
rect 640 11368 648 11432
rect 712 11368 720 11432
rect 640 11272 720 11368
rect 640 11208 648 11272
rect 712 11208 720 11272
rect 640 11112 720 11208
rect 640 11048 648 11112
rect 712 11048 720 11112
rect 640 10952 720 11048
rect 640 10888 648 10952
rect 712 10888 720 10952
rect 640 10792 720 10888
rect 640 10728 648 10792
rect 712 10728 720 10792
rect 640 10472 720 10728
rect 640 10408 648 10472
rect 712 10408 720 10472
rect 640 10152 720 10408
rect 640 10088 648 10152
rect 712 10088 720 10152
rect 640 9992 720 10088
rect 640 9928 648 9992
rect 712 9928 720 9992
rect 640 9832 720 9928
rect 640 9768 648 9832
rect 712 9768 720 9832
rect 640 9672 720 9768
rect 640 9608 648 9672
rect 712 9608 720 9672
rect 640 9512 720 9608
rect 640 9448 648 9512
rect 712 9448 720 9512
rect 640 9352 720 9448
rect 640 9288 648 9352
rect 712 9288 720 9352
rect 640 9192 720 9288
rect 640 9128 648 9192
rect 712 9128 720 9192
rect 640 9032 720 9128
rect 640 8968 648 9032
rect 712 8968 720 9032
rect 640 8872 720 8968
rect 640 8808 648 8872
rect 712 8808 720 8872
rect 640 8712 720 8808
rect 640 8648 648 8712
rect 712 8648 720 8712
rect 640 8552 720 8648
rect 640 8488 648 8552
rect 712 8488 720 8552
rect 640 8392 720 8488
rect 640 8328 648 8392
rect 712 8328 720 8392
rect 640 8232 720 8328
rect 640 8168 648 8232
rect 712 8168 720 8232
rect 640 8072 720 8168
rect 640 8008 648 8072
rect 712 8008 720 8072
rect 640 7912 720 8008
rect 640 7848 648 7912
rect 712 7848 720 7912
rect 640 7752 720 7848
rect 640 7688 648 7752
rect 712 7688 720 7752
rect 640 7592 720 7688
rect 640 7528 648 7592
rect 712 7528 720 7592
rect 640 7432 720 7528
rect 640 7368 648 7432
rect 712 7368 720 7432
rect 640 7272 720 7368
rect 640 7208 648 7272
rect 712 7208 720 7272
rect 640 7112 720 7208
rect 640 7048 648 7112
rect 712 7048 720 7112
rect 640 6952 720 7048
rect 640 6888 648 6952
rect 712 6888 720 6952
rect 640 6792 720 6888
rect 640 6728 648 6792
rect 712 6728 720 6792
rect 640 6632 720 6728
rect 640 6568 648 6632
rect 712 6568 720 6632
rect 640 6472 720 6568
rect 640 6408 648 6472
rect 712 6408 720 6472
rect 640 6312 720 6408
rect 640 6248 648 6312
rect 712 6248 720 6312
rect 640 6152 720 6248
rect 640 6088 648 6152
rect 712 6088 720 6152
rect 640 5992 720 6088
rect 640 5928 648 5992
rect 712 5928 720 5992
rect 640 5832 720 5928
rect 640 5768 648 5832
rect 712 5768 720 5832
rect 640 5672 720 5768
rect 640 5608 648 5672
rect 712 5608 720 5672
rect 640 5512 720 5608
rect 640 5448 648 5512
rect 712 5448 720 5512
rect 640 5352 720 5448
rect 640 5288 648 5352
rect 712 5288 720 5352
rect 640 5192 720 5288
rect 640 5128 648 5192
rect 712 5128 720 5192
rect 640 5032 720 5128
rect 640 4968 648 5032
rect 712 4968 720 5032
rect 640 4872 720 4968
rect 640 4808 648 4872
rect 712 4808 720 4872
rect 640 4712 720 4808
rect 640 4648 648 4712
rect 712 4648 720 4712
rect 640 4552 720 4648
rect 640 4488 648 4552
rect 712 4488 720 4552
rect 640 4392 720 4488
rect 640 4328 648 4392
rect 712 4328 720 4392
rect 640 4232 720 4328
rect 640 4168 648 4232
rect 712 4168 720 4232
rect 640 4072 720 4168
rect 640 4008 648 4072
rect 712 4008 720 4072
rect 640 3912 720 4008
rect 640 3848 648 3912
rect 712 3848 720 3912
rect 640 3752 720 3848
rect 640 3688 648 3752
rect 712 3688 720 3752
rect 640 3592 720 3688
rect 640 3528 648 3592
rect 712 3528 720 3592
rect 640 3432 720 3528
rect 640 3368 648 3432
rect 712 3368 720 3432
rect 640 3272 720 3368
rect 640 3208 648 3272
rect 712 3208 720 3272
rect 640 3112 720 3208
rect 640 3048 648 3112
rect 712 3048 720 3112
rect 640 2952 720 3048
rect 640 2888 648 2952
rect 712 2888 720 2952
rect 640 2792 720 2888
rect 640 2728 648 2792
rect 712 2728 720 2792
rect 640 2632 720 2728
rect 640 2568 648 2632
rect 712 2568 720 2632
rect 640 2472 720 2568
rect 640 2408 648 2472
rect 712 2408 720 2472
rect 640 2312 720 2408
rect 640 2248 648 2312
rect 712 2248 720 2312
rect 640 2152 720 2248
rect 640 2088 648 2152
rect 712 2088 720 2152
rect 640 1992 720 2088
rect 640 1928 648 1992
rect 712 1928 720 1992
rect 640 1832 720 1928
rect 640 1768 648 1832
rect 712 1768 720 1832
rect 640 1672 720 1768
rect 640 1608 648 1672
rect 712 1608 720 1672
rect 640 1512 720 1608
rect 640 1448 648 1512
rect 712 1448 720 1512
rect 640 1352 720 1448
rect 640 1288 648 1352
rect 712 1288 720 1352
rect 640 1192 720 1288
rect 640 1128 648 1192
rect 712 1128 720 1192
rect 640 1032 720 1128
rect 640 968 648 1032
rect 712 968 720 1032
rect 320 808 328 872
rect 392 808 400 872
rect 320 792 400 808
rect 320 728 328 792
rect 392 728 400 792
rect 320 712 400 728
rect 320 648 328 712
rect 392 648 400 712
rect 320 632 400 648
rect 320 568 328 632
rect 392 568 400 632
rect 320 552 400 568
rect 320 488 328 552
rect 392 488 400 552
rect 320 480 400 488
rect 640 872 720 968
rect 800 19752 880 31920
rect 800 19688 808 19752
rect 872 19688 880 19752
rect 800 13192 880 19688
rect 800 13128 808 13192
rect 872 13128 880 13192
rect 800 960 880 13128
rect 960 31912 1040 31920
rect 960 31848 968 31912
rect 1032 31848 1040 31912
rect 960 31752 1040 31848
rect 960 31688 968 31752
rect 1032 31688 1040 31752
rect 960 31592 1040 31688
rect 960 31528 968 31592
rect 1032 31528 1040 31592
rect 960 31432 1040 31528
rect 960 31368 968 31432
rect 1032 31368 1040 31432
rect 960 31272 1040 31368
rect 960 31208 968 31272
rect 1032 31208 1040 31272
rect 960 31112 1040 31208
rect 960 31048 968 31112
rect 1032 31048 1040 31112
rect 960 30952 1040 31048
rect 960 30888 968 30952
rect 1032 30888 1040 30952
rect 960 30792 1040 30888
rect 960 30728 968 30792
rect 1032 30728 1040 30792
rect 960 30632 1040 30728
rect 960 30568 968 30632
rect 1032 30568 1040 30632
rect 960 30472 1040 30568
rect 960 30408 968 30472
rect 1032 30408 1040 30472
rect 960 30312 1040 30408
rect 960 30248 968 30312
rect 1032 30248 1040 30312
rect 960 30152 1040 30248
rect 960 30088 968 30152
rect 1032 30088 1040 30152
rect 960 29992 1040 30088
rect 960 29928 968 29992
rect 1032 29928 1040 29992
rect 960 29832 1040 29928
rect 960 29768 968 29832
rect 1032 29768 1040 29832
rect 960 29672 1040 29768
rect 960 29608 968 29672
rect 1032 29608 1040 29672
rect 960 29512 1040 29608
rect 960 29448 968 29512
rect 1032 29448 1040 29512
rect 960 29352 1040 29448
rect 960 29288 968 29352
rect 1032 29288 1040 29352
rect 960 29192 1040 29288
rect 960 29128 968 29192
rect 1032 29128 1040 29192
rect 960 29032 1040 29128
rect 960 28968 968 29032
rect 1032 28968 1040 29032
rect 960 28872 1040 28968
rect 960 28808 968 28872
rect 1032 28808 1040 28872
rect 960 28712 1040 28808
rect 960 28648 968 28712
rect 1032 28648 1040 28712
rect 960 28552 1040 28648
rect 960 28488 968 28552
rect 1032 28488 1040 28552
rect 960 28392 1040 28488
rect 960 28328 968 28392
rect 1032 28328 1040 28392
rect 960 28232 1040 28328
rect 960 28168 968 28232
rect 1032 28168 1040 28232
rect 960 28072 1040 28168
rect 960 28008 968 28072
rect 1032 28008 1040 28072
rect 960 27912 1040 28008
rect 960 27848 968 27912
rect 1032 27848 1040 27912
rect 960 27752 1040 27848
rect 960 27688 968 27752
rect 1032 27688 1040 27752
rect 960 27592 1040 27688
rect 960 27528 968 27592
rect 1032 27528 1040 27592
rect 960 27432 1040 27528
rect 960 27368 968 27432
rect 1032 27368 1040 27432
rect 960 27272 1040 27368
rect 960 27208 968 27272
rect 1032 27208 1040 27272
rect 960 27112 1040 27208
rect 960 27048 968 27112
rect 1032 27048 1040 27112
rect 960 26952 1040 27048
rect 960 26888 968 26952
rect 1032 26888 1040 26952
rect 960 26792 1040 26888
rect 960 26728 968 26792
rect 1032 26728 1040 26792
rect 960 26632 1040 26728
rect 960 26568 968 26632
rect 1032 26568 1040 26632
rect 960 26472 1040 26568
rect 960 26408 968 26472
rect 1032 26408 1040 26472
rect 960 26312 1040 26408
rect 960 26248 968 26312
rect 1032 26248 1040 26312
rect 960 26152 1040 26248
rect 960 26088 968 26152
rect 1032 26088 1040 26152
rect 960 25992 1040 26088
rect 960 25928 968 25992
rect 1032 25928 1040 25992
rect 960 25832 1040 25928
rect 960 25768 968 25832
rect 1032 25768 1040 25832
rect 960 25672 1040 25768
rect 960 25608 968 25672
rect 1032 25608 1040 25672
rect 960 25512 1040 25608
rect 960 25448 968 25512
rect 1032 25448 1040 25512
rect 960 25352 1040 25448
rect 960 25288 968 25352
rect 1032 25288 1040 25352
rect 960 25192 1040 25288
rect 960 25128 968 25192
rect 1032 25128 1040 25192
rect 960 25032 1040 25128
rect 960 24968 968 25032
rect 1032 24968 1040 25032
rect 960 24872 1040 24968
rect 960 24808 968 24872
rect 1032 24808 1040 24872
rect 960 24712 1040 24808
rect 960 24648 968 24712
rect 1032 24648 1040 24712
rect 960 24552 1040 24648
rect 960 24488 968 24552
rect 1032 24488 1040 24552
rect 960 24392 1040 24488
rect 960 24328 968 24392
rect 1032 24328 1040 24392
rect 960 24232 1040 24328
rect 960 24168 968 24232
rect 1032 24168 1040 24232
rect 960 24072 1040 24168
rect 960 24008 968 24072
rect 1032 24008 1040 24072
rect 960 23912 1040 24008
rect 960 23848 968 23912
rect 1032 23848 1040 23912
rect 960 23752 1040 23848
rect 960 23688 968 23752
rect 1032 23688 1040 23752
rect 960 23592 1040 23688
rect 960 23528 968 23592
rect 1032 23528 1040 23592
rect 960 23432 1040 23528
rect 960 23368 968 23432
rect 1032 23368 1040 23432
rect 960 23272 1040 23368
rect 960 23208 968 23272
rect 1032 23208 1040 23272
rect 960 23112 1040 23208
rect 960 23048 968 23112
rect 1032 23048 1040 23112
rect 960 22952 1040 23048
rect 960 22888 968 22952
rect 1032 22888 1040 22952
rect 960 22792 1040 22888
rect 960 22728 968 22792
rect 1032 22728 1040 22792
rect 960 22472 1040 22728
rect 960 22408 968 22472
rect 1032 22408 1040 22472
rect 960 22152 1040 22408
rect 960 22088 968 22152
rect 1032 22088 1040 22152
rect 960 21992 1040 22088
rect 960 21928 968 21992
rect 1032 21928 1040 21992
rect 960 21832 1040 21928
rect 960 21768 968 21832
rect 1032 21768 1040 21832
rect 960 21672 1040 21768
rect 960 21608 968 21672
rect 1032 21608 1040 21672
rect 960 21512 1040 21608
rect 960 21448 968 21512
rect 1032 21448 1040 21512
rect 960 21352 1040 21448
rect 960 21288 968 21352
rect 1032 21288 1040 21352
rect 960 21192 1040 21288
rect 960 21128 968 21192
rect 1032 21128 1040 21192
rect 960 21032 1040 21128
rect 960 20968 968 21032
rect 1032 20968 1040 21032
rect 960 20872 1040 20968
rect 960 20808 968 20872
rect 1032 20808 1040 20872
rect 960 20712 1040 20808
rect 960 20648 968 20712
rect 1032 20648 1040 20712
rect 960 20552 1040 20648
rect 960 20488 968 20552
rect 1032 20488 1040 20552
rect 960 20392 1040 20488
rect 960 20328 968 20392
rect 1032 20328 1040 20392
rect 960 20232 1040 20328
rect 960 20168 968 20232
rect 1032 20168 1040 20232
rect 960 20072 1040 20168
rect 960 20008 968 20072
rect 1032 20008 1040 20072
rect 960 19912 1040 20008
rect 960 19848 968 19912
rect 1032 19848 1040 19912
rect 960 19592 1040 19848
rect 960 19528 968 19592
rect 1032 19528 1040 19592
rect 960 19432 1040 19528
rect 960 19368 968 19432
rect 1032 19368 1040 19432
rect 960 19272 1040 19368
rect 960 19208 968 19272
rect 1032 19208 1040 19272
rect 960 19112 1040 19208
rect 960 19048 968 19112
rect 1032 19048 1040 19112
rect 960 18952 1040 19048
rect 960 18888 968 18952
rect 1032 18888 1040 18952
rect 960 18792 1040 18888
rect 960 18728 968 18792
rect 1032 18728 1040 18792
rect 960 18632 1040 18728
rect 960 18568 968 18632
rect 1032 18568 1040 18632
rect 960 18472 1040 18568
rect 960 18408 968 18472
rect 1032 18408 1040 18472
rect 960 18312 1040 18408
rect 960 18248 968 18312
rect 1032 18248 1040 18312
rect 960 18152 1040 18248
rect 960 18088 968 18152
rect 1032 18088 1040 18152
rect 960 17992 1040 18088
rect 960 17928 968 17992
rect 1032 17928 1040 17992
rect 960 17832 1040 17928
rect 960 17768 968 17832
rect 1032 17768 1040 17832
rect 960 17672 1040 17768
rect 960 17608 968 17672
rect 1032 17608 1040 17672
rect 960 17512 1040 17608
rect 960 17448 968 17512
rect 1032 17448 1040 17512
rect 960 17352 1040 17448
rect 960 17288 968 17352
rect 1032 17288 1040 17352
rect 960 17032 1040 17288
rect 960 16968 968 17032
rect 1032 16968 1040 17032
rect 960 16712 1040 16968
rect 960 16648 968 16712
rect 1032 16648 1040 16712
rect 960 16552 1040 16648
rect 960 16488 968 16552
rect 1032 16488 1040 16552
rect 960 16392 1040 16488
rect 960 16328 968 16392
rect 1032 16328 1040 16392
rect 960 16232 1040 16328
rect 960 16168 968 16232
rect 1032 16168 1040 16232
rect 960 15912 1040 16168
rect 960 15848 968 15912
rect 1032 15848 1040 15912
rect 960 15592 1040 15848
rect 960 15528 968 15592
rect 1032 15528 1040 15592
rect 960 15432 1040 15528
rect 960 15368 968 15432
rect 1032 15368 1040 15432
rect 960 15272 1040 15368
rect 960 15208 968 15272
rect 1032 15208 1040 15272
rect 960 15112 1040 15208
rect 960 15048 968 15112
rect 1032 15048 1040 15112
rect 960 14952 1040 15048
rect 960 14888 968 14952
rect 1032 14888 1040 14952
rect 960 14792 1040 14888
rect 960 14728 968 14792
rect 1032 14728 1040 14792
rect 960 14632 1040 14728
rect 960 14568 968 14632
rect 1032 14568 1040 14632
rect 960 14472 1040 14568
rect 960 14408 968 14472
rect 1032 14408 1040 14472
rect 960 14312 1040 14408
rect 960 14248 968 14312
rect 1032 14248 1040 14312
rect 960 14152 1040 14248
rect 960 14088 968 14152
rect 1032 14088 1040 14152
rect 960 13992 1040 14088
rect 960 13928 968 13992
rect 1032 13928 1040 13992
rect 960 13832 1040 13928
rect 960 13768 968 13832
rect 1032 13768 1040 13832
rect 960 13672 1040 13768
rect 960 13608 968 13672
rect 1032 13608 1040 13672
rect 960 13512 1040 13608
rect 960 13448 968 13512
rect 1032 13448 1040 13512
rect 960 13352 1040 13448
rect 960 13288 968 13352
rect 1032 13288 1040 13352
rect 960 13032 1040 13288
rect 960 12968 968 13032
rect 1032 12968 1040 13032
rect 960 12872 1040 12968
rect 960 12808 968 12872
rect 1032 12808 1040 12872
rect 960 12712 1040 12808
rect 960 12648 968 12712
rect 1032 12648 1040 12712
rect 960 12552 1040 12648
rect 960 12488 968 12552
rect 1032 12488 1040 12552
rect 960 12392 1040 12488
rect 960 12328 968 12392
rect 1032 12328 1040 12392
rect 960 12232 1040 12328
rect 960 12168 968 12232
rect 1032 12168 1040 12232
rect 960 12072 1040 12168
rect 960 12008 968 12072
rect 1032 12008 1040 12072
rect 960 11912 1040 12008
rect 960 11848 968 11912
rect 1032 11848 1040 11912
rect 960 11752 1040 11848
rect 960 11688 968 11752
rect 1032 11688 1040 11752
rect 960 11592 1040 11688
rect 960 11528 968 11592
rect 1032 11528 1040 11592
rect 960 11432 1040 11528
rect 960 11368 968 11432
rect 1032 11368 1040 11432
rect 960 11272 1040 11368
rect 960 11208 968 11272
rect 1032 11208 1040 11272
rect 960 11112 1040 11208
rect 960 11048 968 11112
rect 1032 11048 1040 11112
rect 960 10952 1040 11048
rect 960 10888 968 10952
rect 1032 10888 1040 10952
rect 960 10792 1040 10888
rect 960 10728 968 10792
rect 1032 10728 1040 10792
rect 960 10472 1040 10728
rect 960 10408 968 10472
rect 1032 10408 1040 10472
rect 960 10152 1040 10408
rect 960 10088 968 10152
rect 1032 10088 1040 10152
rect 960 9992 1040 10088
rect 960 9928 968 9992
rect 1032 9928 1040 9992
rect 960 9832 1040 9928
rect 960 9768 968 9832
rect 1032 9768 1040 9832
rect 960 9672 1040 9768
rect 960 9608 968 9672
rect 1032 9608 1040 9672
rect 960 9512 1040 9608
rect 960 9448 968 9512
rect 1032 9448 1040 9512
rect 960 9352 1040 9448
rect 960 9288 968 9352
rect 1032 9288 1040 9352
rect 960 9192 1040 9288
rect 960 9128 968 9192
rect 1032 9128 1040 9192
rect 960 9032 1040 9128
rect 960 8968 968 9032
rect 1032 8968 1040 9032
rect 960 8872 1040 8968
rect 960 8808 968 8872
rect 1032 8808 1040 8872
rect 960 8712 1040 8808
rect 960 8648 968 8712
rect 1032 8648 1040 8712
rect 960 8552 1040 8648
rect 960 8488 968 8552
rect 1032 8488 1040 8552
rect 960 8392 1040 8488
rect 960 8328 968 8392
rect 1032 8328 1040 8392
rect 960 8232 1040 8328
rect 960 8168 968 8232
rect 1032 8168 1040 8232
rect 960 8072 1040 8168
rect 960 8008 968 8072
rect 1032 8008 1040 8072
rect 960 7912 1040 8008
rect 960 7848 968 7912
rect 1032 7848 1040 7912
rect 960 7752 1040 7848
rect 960 7688 968 7752
rect 1032 7688 1040 7752
rect 960 7592 1040 7688
rect 960 7528 968 7592
rect 1032 7528 1040 7592
rect 960 7432 1040 7528
rect 960 7368 968 7432
rect 1032 7368 1040 7432
rect 960 7272 1040 7368
rect 960 7208 968 7272
rect 1032 7208 1040 7272
rect 960 7112 1040 7208
rect 960 7048 968 7112
rect 1032 7048 1040 7112
rect 960 6952 1040 7048
rect 960 6888 968 6952
rect 1032 6888 1040 6952
rect 960 6792 1040 6888
rect 960 6728 968 6792
rect 1032 6728 1040 6792
rect 960 6632 1040 6728
rect 960 6568 968 6632
rect 1032 6568 1040 6632
rect 960 6472 1040 6568
rect 960 6408 968 6472
rect 1032 6408 1040 6472
rect 960 6312 1040 6408
rect 960 6248 968 6312
rect 1032 6248 1040 6312
rect 960 6152 1040 6248
rect 960 6088 968 6152
rect 1032 6088 1040 6152
rect 960 5992 1040 6088
rect 960 5928 968 5992
rect 1032 5928 1040 5992
rect 960 5832 1040 5928
rect 960 5768 968 5832
rect 1032 5768 1040 5832
rect 960 5672 1040 5768
rect 960 5608 968 5672
rect 1032 5608 1040 5672
rect 960 5512 1040 5608
rect 960 5448 968 5512
rect 1032 5448 1040 5512
rect 960 5352 1040 5448
rect 960 5288 968 5352
rect 1032 5288 1040 5352
rect 960 5192 1040 5288
rect 960 5128 968 5192
rect 1032 5128 1040 5192
rect 960 5032 1040 5128
rect 960 4968 968 5032
rect 1032 4968 1040 5032
rect 960 4872 1040 4968
rect 960 4808 968 4872
rect 1032 4808 1040 4872
rect 960 4712 1040 4808
rect 960 4648 968 4712
rect 1032 4648 1040 4712
rect 960 4552 1040 4648
rect 960 4488 968 4552
rect 1032 4488 1040 4552
rect 960 4392 1040 4488
rect 960 4328 968 4392
rect 1032 4328 1040 4392
rect 960 4232 1040 4328
rect 960 4168 968 4232
rect 1032 4168 1040 4232
rect 960 4072 1040 4168
rect 960 4008 968 4072
rect 1032 4008 1040 4072
rect 960 3912 1040 4008
rect 960 3848 968 3912
rect 1032 3848 1040 3912
rect 960 3752 1040 3848
rect 960 3688 968 3752
rect 1032 3688 1040 3752
rect 960 3592 1040 3688
rect 960 3528 968 3592
rect 1032 3528 1040 3592
rect 960 3432 1040 3528
rect 960 3368 968 3432
rect 1032 3368 1040 3432
rect 960 3272 1040 3368
rect 960 3208 968 3272
rect 1032 3208 1040 3272
rect 960 3112 1040 3208
rect 960 3048 968 3112
rect 1032 3048 1040 3112
rect 960 2952 1040 3048
rect 960 2888 968 2952
rect 1032 2888 1040 2952
rect 960 2792 1040 2888
rect 960 2728 968 2792
rect 1032 2728 1040 2792
rect 960 2632 1040 2728
rect 960 2568 968 2632
rect 1032 2568 1040 2632
rect 960 2472 1040 2568
rect 960 2408 968 2472
rect 1032 2408 1040 2472
rect 960 2312 1040 2408
rect 960 2248 968 2312
rect 1032 2248 1040 2312
rect 960 2152 1040 2248
rect 960 2088 968 2152
rect 1032 2088 1040 2152
rect 960 1992 1040 2088
rect 960 1928 968 1992
rect 1032 1928 1040 1992
rect 960 1832 1040 1928
rect 960 1768 968 1832
rect 1032 1768 1040 1832
rect 960 1672 1040 1768
rect 960 1608 968 1672
rect 1032 1608 1040 1672
rect 960 1512 1040 1608
rect 960 1448 968 1512
rect 1032 1448 1040 1512
rect 960 1352 1040 1448
rect 960 1288 968 1352
rect 1032 1288 1040 1352
rect 960 1192 1040 1288
rect 960 1128 968 1192
rect 1032 1128 1040 1192
rect 960 1032 1040 1128
rect 28960 31912 29040 31920
rect 28960 31848 28968 31912
rect 29032 31848 29040 31912
rect 28960 31752 29040 31848
rect 28960 31688 28968 31752
rect 29032 31688 29040 31752
rect 28960 31592 29040 31688
rect 28960 31528 28968 31592
rect 29032 31528 29040 31592
rect 28960 31432 29040 31528
rect 28960 31368 28968 31432
rect 29032 31368 29040 31432
rect 28960 31272 29040 31368
rect 28960 31208 28968 31272
rect 29032 31208 29040 31272
rect 28960 31112 29040 31208
rect 28960 31048 28968 31112
rect 29032 31048 29040 31112
rect 28960 30952 29040 31048
rect 28960 30888 28968 30952
rect 29032 30888 29040 30952
rect 28960 30792 29040 30888
rect 28960 30728 28968 30792
rect 29032 30728 29040 30792
rect 28960 30632 29040 30728
rect 28960 30568 28968 30632
rect 29032 30568 29040 30632
rect 28960 30472 29040 30568
rect 28960 30408 28968 30472
rect 29032 30408 29040 30472
rect 28960 30312 29040 30408
rect 28960 30248 28968 30312
rect 29032 30248 29040 30312
rect 28960 30152 29040 30248
rect 28960 30088 28968 30152
rect 29032 30088 29040 30152
rect 28960 29992 29040 30088
rect 28960 29928 28968 29992
rect 29032 29928 29040 29992
rect 28960 29832 29040 29928
rect 28960 29768 28968 29832
rect 29032 29768 29040 29832
rect 28960 29672 29040 29768
rect 28960 29608 28968 29672
rect 29032 29608 29040 29672
rect 28960 29512 29040 29608
rect 28960 29448 28968 29512
rect 29032 29448 29040 29512
rect 28960 29352 29040 29448
rect 28960 29288 28968 29352
rect 29032 29288 29040 29352
rect 28960 29032 29040 29288
rect 28960 28968 28968 29032
rect 29032 28968 29040 29032
rect 28960 28712 29040 28968
rect 28960 28648 28968 28712
rect 29032 28648 29040 28712
rect 28960 28552 29040 28648
rect 28960 28488 28968 28552
rect 29032 28488 29040 28552
rect 28960 28392 29040 28488
rect 28960 28328 28968 28392
rect 29032 28328 29040 28392
rect 28960 28232 29040 28328
rect 28960 28168 28968 28232
rect 29032 28168 29040 28232
rect 28960 28072 29040 28168
rect 28960 28008 28968 28072
rect 29032 28008 29040 28072
rect 28960 27912 29040 28008
rect 28960 27848 28968 27912
rect 29032 27848 29040 27912
rect 28960 27752 29040 27848
rect 28960 27688 28968 27752
rect 29032 27688 29040 27752
rect 28960 27592 29040 27688
rect 28960 27528 28968 27592
rect 29032 27528 29040 27592
rect 28960 27432 29040 27528
rect 28960 27368 28968 27432
rect 29032 27368 29040 27432
rect 28960 27272 29040 27368
rect 28960 27208 28968 27272
rect 29032 27208 29040 27272
rect 28960 27112 29040 27208
rect 28960 27048 28968 27112
rect 29032 27048 29040 27112
rect 28960 26952 29040 27048
rect 28960 26888 28968 26952
rect 29032 26888 29040 26952
rect 28960 26792 29040 26888
rect 28960 26728 28968 26792
rect 29032 26728 29040 26792
rect 28960 26632 29040 26728
rect 28960 26568 28968 26632
rect 29032 26568 29040 26632
rect 28960 26472 29040 26568
rect 28960 26408 28968 26472
rect 29032 26408 29040 26472
rect 28960 26152 29040 26408
rect 28960 26088 28968 26152
rect 29032 26088 29040 26152
rect 28960 25992 29040 26088
rect 28960 25928 28968 25992
rect 29032 25928 29040 25992
rect 28960 25832 29040 25928
rect 28960 25768 28968 25832
rect 29032 25768 29040 25832
rect 28960 25672 29040 25768
rect 28960 25608 28968 25672
rect 29032 25608 29040 25672
rect 28960 25512 29040 25608
rect 28960 25448 28968 25512
rect 29032 25448 29040 25512
rect 28960 25352 29040 25448
rect 28960 25288 28968 25352
rect 29032 25288 29040 25352
rect 28960 25192 29040 25288
rect 28960 25128 28968 25192
rect 29032 25128 29040 25192
rect 28960 25032 29040 25128
rect 28960 24968 28968 25032
rect 29032 24968 29040 25032
rect 28960 24872 29040 24968
rect 28960 24808 28968 24872
rect 29032 24808 29040 24872
rect 28960 24712 29040 24808
rect 28960 24648 28968 24712
rect 29032 24648 29040 24712
rect 28960 24552 29040 24648
rect 28960 24488 28968 24552
rect 29032 24488 29040 24552
rect 28960 24392 29040 24488
rect 28960 24328 28968 24392
rect 29032 24328 29040 24392
rect 28960 24232 29040 24328
rect 28960 24168 28968 24232
rect 29032 24168 29040 24232
rect 28960 24072 29040 24168
rect 28960 24008 28968 24072
rect 29032 24008 29040 24072
rect 28960 23912 29040 24008
rect 28960 23848 28968 23912
rect 29032 23848 29040 23912
rect 28960 23592 29040 23848
rect 28960 23528 28968 23592
rect 29032 23528 29040 23592
rect 28960 23272 29040 23528
rect 28960 23208 28968 23272
rect 29032 23208 29040 23272
rect 28960 23112 29040 23208
rect 28960 23048 28968 23112
rect 29032 23048 29040 23112
rect 28960 22952 29040 23048
rect 28960 22888 28968 22952
rect 29032 22888 29040 22952
rect 28960 22792 29040 22888
rect 28960 22728 28968 22792
rect 29032 22728 29040 22792
rect 28960 22632 29040 22728
rect 28960 22568 28968 22632
rect 29032 22568 29040 22632
rect 28960 22472 29040 22568
rect 28960 22408 28968 22472
rect 29032 22408 29040 22472
rect 28960 22312 29040 22408
rect 28960 22248 28968 22312
rect 29032 22248 29040 22312
rect 28960 22152 29040 22248
rect 28960 22088 28968 22152
rect 29032 22088 29040 22152
rect 28960 21992 29040 22088
rect 28960 21928 28968 21992
rect 29032 21928 29040 21992
rect 28960 21832 29040 21928
rect 28960 21768 28968 21832
rect 29032 21768 29040 21832
rect 28960 21672 29040 21768
rect 28960 21608 28968 21672
rect 29032 21608 29040 21672
rect 28960 21512 29040 21608
rect 28960 21448 28968 21512
rect 29032 21448 29040 21512
rect 28960 21352 29040 21448
rect 28960 21288 28968 21352
rect 29032 21288 29040 21352
rect 28960 21192 29040 21288
rect 28960 21128 28968 21192
rect 29032 21128 29040 21192
rect 28960 21032 29040 21128
rect 28960 20968 28968 21032
rect 29032 20968 29040 21032
rect 28960 20872 29040 20968
rect 28960 20808 28968 20872
rect 29032 20808 29040 20872
rect 28960 20712 29040 20808
rect 28960 20648 28968 20712
rect 29032 20648 29040 20712
rect 28960 20552 29040 20648
rect 28960 20488 28968 20552
rect 29032 20488 29040 20552
rect 28960 20392 29040 20488
rect 28960 20328 28968 20392
rect 29032 20328 29040 20392
rect 28960 20232 29040 20328
rect 28960 20168 28968 20232
rect 29032 20168 29040 20232
rect 28960 20072 29040 20168
rect 28960 20008 28968 20072
rect 29032 20008 29040 20072
rect 28960 19912 29040 20008
rect 28960 19848 28968 19912
rect 29032 19848 29040 19912
rect 28960 19752 29040 19848
rect 28960 19688 28968 19752
rect 29032 19688 29040 19752
rect 28960 19592 29040 19688
rect 28960 19528 28968 19592
rect 29032 19528 29040 19592
rect 28960 19432 29040 19528
rect 28960 19368 28968 19432
rect 29032 19368 29040 19432
rect 28960 19272 29040 19368
rect 28960 19208 28968 19272
rect 29032 19208 29040 19272
rect 28960 19112 29040 19208
rect 28960 19048 28968 19112
rect 29032 19048 29040 19112
rect 28960 18952 29040 19048
rect 28960 18888 28968 18952
rect 29032 18888 29040 18952
rect 28960 18792 29040 18888
rect 28960 18728 28968 18792
rect 29032 18728 29040 18792
rect 28960 18632 29040 18728
rect 28960 18568 28968 18632
rect 29032 18568 29040 18632
rect 28960 18472 29040 18568
rect 28960 18408 28968 18472
rect 29032 18408 29040 18472
rect 28960 18312 29040 18408
rect 28960 18248 28968 18312
rect 29032 18248 29040 18312
rect 28960 18152 29040 18248
rect 28960 18088 28968 18152
rect 29032 18088 29040 18152
rect 28960 17992 29040 18088
rect 28960 17928 28968 17992
rect 29032 17928 29040 17992
rect 28960 17832 29040 17928
rect 28960 17768 28968 17832
rect 29032 17768 29040 17832
rect 28960 17672 29040 17768
rect 28960 17608 28968 17672
rect 29032 17608 29040 17672
rect 28960 17512 29040 17608
rect 28960 17448 28968 17512
rect 29032 17448 29040 17512
rect 28960 17352 29040 17448
rect 28960 17288 28968 17352
rect 29032 17288 29040 17352
rect 28960 17192 29040 17288
rect 28960 17128 28968 17192
rect 29032 17128 29040 17192
rect 28960 17032 29040 17128
rect 28960 16968 28968 17032
rect 29032 16968 29040 17032
rect 28960 16872 29040 16968
rect 28960 16808 28968 16872
rect 29032 16808 29040 16872
rect 28960 16712 29040 16808
rect 28960 16648 28968 16712
rect 29032 16648 29040 16712
rect 28960 16552 29040 16648
rect 28960 16488 28968 16552
rect 29032 16488 29040 16552
rect 28960 16392 29040 16488
rect 28960 16328 28968 16392
rect 29032 16328 29040 16392
rect 28960 16232 29040 16328
rect 28960 16168 28968 16232
rect 29032 16168 29040 16232
rect 28960 16072 29040 16168
rect 28960 16008 28968 16072
rect 29032 16008 29040 16072
rect 28960 15912 29040 16008
rect 28960 15848 28968 15912
rect 29032 15848 29040 15912
rect 28960 15752 29040 15848
rect 28960 15688 28968 15752
rect 29032 15688 29040 15752
rect 28960 15592 29040 15688
rect 28960 15528 28968 15592
rect 29032 15528 29040 15592
rect 28960 15432 29040 15528
rect 28960 15368 28968 15432
rect 29032 15368 29040 15432
rect 28960 15272 29040 15368
rect 28960 15208 28968 15272
rect 29032 15208 29040 15272
rect 28960 15112 29040 15208
rect 28960 15048 28968 15112
rect 29032 15048 29040 15112
rect 28960 14952 29040 15048
rect 28960 14888 28968 14952
rect 29032 14888 29040 14952
rect 28960 14792 29040 14888
rect 28960 14728 28968 14792
rect 29032 14728 29040 14792
rect 28960 14632 29040 14728
rect 28960 14568 28968 14632
rect 29032 14568 29040 14632
rect 28960 14472 29040 14568
rect 28960 14408 28968 14472
rect 29032 14408 29040 14472
rect 28960 14312 29040 14408
rect 28960 14248 28968 14312
rect 29032 14248 29040 14312
rect 28960 14152 29040 14248
rect 28960 14088 28968 14152
rect 29032 14088 29040 14152
rect 28960 13992 29040 14088
rect 28960 13928 28968 13992
rect 29032 13928 29040 13992
rect 28960 13832 29040 13928
rect 28960 13768 28968 13832
rect 29032 13768 29040 13832
rect 28960 13672 29040 13768
rect 28960 13608 28968 13672
rect 29032 13608 29040 13672
rect 28960 13512 29040 13608
rect 28960 13448 28968 13512
rect 29032 13448 29040 13512
rect 28960 13352 29040 13448
rect 28960 13288 28968 13352
rect 29032 13288 29040 13352
rect 28960 13192 29040 13288
rect 28960 13128 28968 13192
rect 29032 13128 29040 13192
rect 28960 13032 29040 13128
rect 28960 12968 28968 13032
rect 29032 12968 29040 13032
rect 28960 12872 29040 12968
rect 28960 12808 28968 12872
rect 29032 12808 29040 12872
rect 28960 12712 29040 12808
rect 28960 12648 28968 12712
rect 29032 12648 29040 12712
rect 28960 12552 29040 12648
rect 28960 12488 28968 12552
rect 29032 12488 29040 12552
rect 28960 12392 29040 12488
rect 28960 12328 28968 12392
rect 29032 12328 29040 12392
rect 28960 12232 29040 12328
rect 28960 12168 28968 12232
rect 29032 12168 29040 12232
rect 28960 12072 29040 12168
rect 28960 12008 28968 12072
rect 29032 12008 29040 12072
rect 28960 11912 29040 12008
rect 28960 11848 28968 11912
rect 29032 11848 29040 11912
rect 28960 11752 29040 11848
rect 28960 11688 28968 11752
rect 29032 11688 29040 11752
rect 28960 11592 29040 11688
rect 28960 11528 28968 11592
rect 29032 11528 29040 11592
rect 28960 11432 29040 11528
rect 28960 11368 28968 11432
rect 29032 11368 29040 11432
rect 28960 11272 29040 11368
rect 28960 11208 28968 11272
rect 29032 11208 29040 11272
rect 28960 11112 29040 11208
rect 28960 11048 28968 11112
rect 29032 11048 29040 11112
rect 28960 10952 29040 11048
rect 28960 10888 28968 10952
rect 29032 10888 29040 10952
rect 28960 10792 29040 10888
rect 28960 10728 28968 10792
rect 29032 10728 29040 10792
rect 28960 10632 29040 10728
rect 28960 10568 28968 10632
rect 29032 10568 29040 10632
rect 28960 10472 29040 10568
rect 28960 10408 28968 10472
rect 29032 10408 29040 10472
rect 28960 10312 29040 10408
rect 28960 10248 28968 10312
rect 29032 10248 29040 10312
rect 28960 10152 29040 10248
rect 28960 10088 28968 10152
rect 29032 10088 29040 10152
rect 28960 9992 29040 10088
rect 28960 9928 28968 9992
rect 29032 9928 29040 9992
rect 28960 9832 29040 9928
rect 28960 9768 28968 9832
rect 29032 9768 29040 9832
rect 28960 9672 29040 9768
rect 28960 9608 28968 9672
rect 29032 9608 29040 9672
rect 28960 9352 29040 9608
rect 28960 9288 28968 9352
rect 29032 9288 29040 9352
rect 28960 9032 29040 9288
rect 28960 8968 28968 9032
rect 29032 8968 29040 9032
rect 28960 8872 29040 8968
rect 28960 8808 28968 8872
rect 29032 8808 29040 8872
rect 28960 8712 29040 8808
rect 28960 8648 28968 8712
rect 29032 8648 29040 8712
rect 28960 8552 29040 8648
rect 28960 8488 28968 8552
rect 29032 8488 29040 8552
rect 28960 8392 29040 8488
rect 28960 8328 28968 8392
rect 29032 8328 29040 8392
rect 28960 8232 29040 8328
rect 28960 8168 28968 8232
rect 29032 8168 29040 8232
rect 28960 8072 29040 8168
rect 28960 8008 28968 8072
rect 29032 8008 29040 8072
rect 28960 7912 29040 8008
rect 28960 7848 28968 7912
rect 29032 7848 29040 7912
rect 28960 7752 29040 7848
rect 28960 7688 28968 7752
rect 29032 7688 29040 7752
rect 28960 7592 29040 7688
rect 28960 7528 28968 7592
rect 29032 7528 29040 7592
rect 28960 7432 29040 7528
rect 28960 7368 28968 7432
rect 29032 7368 29040 7432
rect 28960 7272 29040 7368
rect 28960 7208 28968 7272
rect 29032 7208 29040 7272
rect 28960 7112 29040 7208
rect 28960 7048 28968 7112
rect 29032 7048 29040 7112
rect 28960 6952 29040 7048
rect 28960 6888 28968 6952
rect 29032 6888 29040 6952
rect 28960 6792 29040 6888
rect 28960 6728 28968 6792
rect 29032 6728 29040 6792
rect 28960 6472 29040 6728
rect 28960 6408 28968 6472
rect 29032 6408 29040 6472
rect 28960 6312 29040 6408
rect 28960 6248 28968 6312
rect 29032 6248 29040 6312
rect 28960 6152 29040 6248
rect 28960 6088 28968 6152
rect 29032 6088 29040 6152
rect 28960 5992 29040 6088
rect 28960 5928 28968 5992
rect 29032 5928 29040 5992
rect 28960 5832 29040 5928
rect 28960 5768 28968 5832
rect 29032 5768 29040 5832
rect 28960 5672 29040 5768
rect 28960 5608 28968 5672
rect 29032 5608 29040 5672
rect 28960 5512 29040 5608
rect 28960 5448 28968 5512
rect 29032 5448 29040 5512
rect 28960 5352 29040 5448
rect 28960 5288 28968 5352
rect 29032 5288 29040 5352
rect 28960 5192 29040 5288
rect 28960 5128 28968 5192
rect 29032 5128 29040 5192
rect 28960 5032 29040 5128
rect 28960 4968 28968 5032
rect 29032 4968 29040 5032
rect 28960 4872 29040 4968
rect 28960 4808 28968 4872
rect 29032 4808 29040 4872
rect 28960 4712 29040 4808
rect 28960 4648 28968 4712
rect 29032 4648 29040 4712
rect 28960 4552 29040 4648
rect 28960 4488 28968 4552
rect 29032 4488 29040 4552
rect 28960 4392 29040 4488
rect 28960 4328 28968 4392
rect 29032 4328 29040 4392
rect 28960 4232 29040 4328
rect 28960 4168 28968 4232
rect 29032 4168 29040 4232
rect 28960 3912 29040 4168
rect 28960 3848 28968 3912
rect 29032 3848 29040 3912
rect 28960 3592 29040 3848
rect 28960 3528 28968 3592
rect 29032 3528 29040 3592
rect 28960 3432 29040 3528
rect 28960 3368 28968 3432
rect 29032 3368 29040 3432
rect 28960 3272 29040 3368
rect 28960 3208 28968 3272
rect 29032 3208 29040 3272
rect 28960 3112 29040 3208
rect 28960 3048 28968 3112
rect 29032 3048 29040 3112
rect 28960 2952 29040 3048
rect 28960 2888 28968 2952
rect 29032 2888 29040 2952
rect 28960 2792 29040 2888
rect 28960 2728 28968 2792
rect 29032 2728 29040 2792
rect 28960 2632 29040 2728
rect 28960 2568 28968 2632
rect 29032 2568 29040 2632
rect 28960 2472 29040 2568
rect 28960 2408 28968 2472
rect 29032 2408 29040 2472
rect 28960 2312 29040 2408
rect 28960 2248 28968 2312
rect 29032 2248 29040 2312
rect 28960 2152 29040 2248
rect 28960 2088 28968 2152
rect 29032 2088 29040 2152
rect 28960 1992 29040 2088
rect 28960 1928 28968 1992
rect 29032 1928 29040 1992
rect 28960 1832 29040 1928
rect 28960 1768 28968 1832
rect 29032 1768 29040 1832
rect 28960 1672 29040 1768
rect 28960 1608 28968 1672
rect 29032 1608 29040 1672
rect 28960 1512 29040 1608
rect 28960 1448 28968 1512
rect 29032 1448 29040 1512
rect 28960 1352 29040 1448
rect 28960 1288 28968 1352
rect 29032 1288 29040 1352
rect 28960 1192 29040 1288
rect 28960 1128 28968 1192
rect 29032 1128 29040 1192
rect 960 968 968 1032
rect 1032 968 1040 1032
rect 640 808 648 872
rect 712 808 720 872
rect 640 792 720 808
rect 640 728 648 792
rect 712 728 720 792
rect 640 712 720 728
rect 640 648 648 712
rect 712 648 720 712
rect 640 632 720 648
rect 640 568 648 632
rect 712 568 720 632
rect 640 552 720 568
rect 640 488 648 552
rect 712 488 720 552
rect 640 480 720 488
rect 960 872 1040 968
rect 960 808 968 872
rect 1032 808 1040 872
rect 960 792 1040 808
rect 960 728 968 792
rect 1032 728 1040 792
rect 960 712 1040 728
rect 960 648 968 712
rect 1032 648 1040 712
rect 960 632 1040 648
rect 960 568 968 632
rect 1032 568 1040 632
rect 960 552 1040 568
rect 960 488 968 552
rect 1032 488 1040 552
rect 960 480 1040 488
rect 1120 1028 1200 1040
rect 1120 972 1132 1028
rect 1188 972 1200 1028
rect 1120 392 1200 972
rect 1120 328 1128 392
rect 1192 328 1200 392
rect 1120 312 1200 328
rect 1120 248 1128 312
rect 1192 248 1200 312
rect 1120 232 1200 248
rect 1120 168 1128 232
rect 1192 168 1200 232
rect 1120 152 1200 168
rect 1120 88 1128 152
rect 1192 88 1200 152
rect 1120 72 1200 88
rect 1120 8 1128 72
rect 1192 8 1200 72
rect 1120 0 1200 8
rect 28800 1028 28880 1040
rect 28800 972 28812 1028
rect 28868 972 28880 1028
rect 28800 392 28880 972
rect 28960 1032 29040 1128
rect 28960 968 28968 1032
rect 29032 968 29040 1032
rect 28960 872 29040 968
rect 29120 26312 29200 31920
rect 29120 26248 29128 26312
rect 29192 26248 29200 26312
rect 29120 6632 29200 26248
rect 29120 6568 29128 6632
rect 29192 6568 29200 6632
rect 29120 960 29200 6568
rect 29280 31912 29360 31920
rect 29280 31848 29288 31912
rect 29352 31848 29360 31912
rect 29280 31752 29360 31848
rect 29280 31688 29288 31752
rect 29352 31688 29360 31752
rect 29280 31592 29360 31688
rect 29280 31528 29288 31592
rect 29352 31528 29360 31592
rect 29280 31432 29360 31528
rect 29280 31368 29288 31432
rect 29352 31368 29360 31432
rect 29280 31272 29360 31368
rect 29280 31208 29288 31272
rect 29352 31208 29360 31272
rect 29280 31112 29360 31208
rect 29280 31048 29288 31112
rect 29352 31048 29360 31112
rect 29280 30952 29360 31048
rect 29280 30888 29288 30952
rect 29352 30888 29360 30952
rect 29280 30792 29360 30888
rect 29280 30728 29288 30792
rect 29352 30728 29360 30792
rect 29280 30632 29360 30728
rect 29280 30568 29288 30632
rect 29352 30568 29360 30632
rect 29280 30472 29360 30568
rect 29280 30408 29288 30472
rect 29352 30408 29360 30472
rect 29280 30312 29360 30408
rect 29280 30248 29288 30312
rect 29352 30248 29360 30312
rect 29280 30152 29360 30248
rect 29280 30088 29288 30152
rect 29352 30088 29360 30152
rect 29280 29992 29360 30088
rect 29280 29928 29288 29992
rect 29352 29928 29360 29992
rect 29280 29832 29360 29928
rect 29280 29768 29288 29832
rect 29352 29768 29360 29832
rect 29280 29672 29360 29768
rect 29280 29608 29288 29672
rect 29352 29608 29360 29672
rect 29280 29512 29360 29608
rect 29280 29448 29288 29512
rect 29352 29448 29360 29512
rect 29280 29352 29360 29448
rect 29280 29288 29288 29352
rect 29352 29288 29360 29352
rect 29280 29032 29360 29288
rect 29280 28968 29288 29032
rect 29352 28968 29360 29032
rect 29280 28712 29360 28968
rect 29280 28648 29288 28712
rect 29352 28648 29360 28712
rect 29280 28552 29360 28648
rect 29280 28488 29288 28552
rect 29352 28488 29360 28552
rect 29280 28392 29360 28488
rect 29280 28328 29288 28392
rect 29352 28328 29360 28392
rect 29280 28232 29360 28328
rect 29280 28168 29288 28232
rect 29352 28168 29360 28232
rect 29280 28072 29360 28168
rect 29280 28008 29288 28072
rect 29352 28008 29360 28072
rect 29280 27912 29360 28008
rect 29280 27848 29288 27912
rect 29352 27848 29360 27912
rect 29280 27752 29360 27848
rect 29280 27688 29288 27752
rect 29352 27688 29360 27752
rect 29280 27592 29360 27688
rect 29280 27528 29288 27592
rect 29352 27528 29360 27592
rect 29280 27432 29360 27528
rect 29280 27368 29288 27432
rect 29352 27368 29360 27432
rect 29280 27272 29360 27368
rect 29280 27208 29288 27272
rect 29352 27208 29360 27272
rect 29280 27112 29360 27208
rect 29280 27048 29288 27112
rect 29352 27048 29360 27112
rect 29280 26952 29360 27048
rect 29280 26888 29288 26952
rect 29352 26888 29360 26952
rect 29280 26792 29360 26888
rect 29280 26728 29288 26792
rect 29352 26728 29360 26792
rect 29280 26632 29360 26728
rect 29280 26568 29288 26632
rect 29352 26568 29360 26632
rect 29280 26472 29360 26568
rect 29280 26408 29288 26472
rect 29352 26408 29360 26472
rect 29280 26312 29360 26408
rect 29280 26248 29288 26312
rect 29352 26248 29360 26312
rect 29280 26152 29360 26248
rect 29280 26088 29288 26152
rect 29352 26088 29360 26152
rect 29280 25992 29360 26088
rect 29280 25928 29288 25992
rect 29352 25928 29360 25992
rect 29280 25832 29360 25928
rect 29280 25768 29288 25832
rect 29352 25768 29360 25832
rect 29280 25672 29360 25768
rect 29280 25608 29288 25672
rect 29352 25608 29360 25672
rect 29280 25512 29360 25608
rect 29280 25448 29288 25512
rect 29352 25448 29360 25512
rect 29280 25352 29360 25448
rect 29280 25288 29288 25352
rect 29352 25288 29360 25352
rect 29280 25192 29360 25288
rect 29280 25128 29288 25192
rect 29352 25128 29360 25192
rect 29280 25032 29360 25128
rect 29280 24968 29288 25032
rect 29352 24968 29360 25032
rect 29280 24872 29360 24968
rect 29280 24808 29288 24872
rect 29352 24808 29360 24872
rect 29280 24712 29360 24808
rect 29280 24648 29288 24712
rect 29352 24648 29360 24712
rect 29280 24552 29360 24648
rect 29280 24488 29288 24552
rect 29352 24488 29360 24552
rect 29280 24392 29360 24488
rect 29280 24328 29288 24392
rect 29352 24328 29360 24392
rect 29280 24232 29360 24328
rect 29280 24168 29288 24232
rect 29352 24168 29360 24232
rect 29280 24072 29360 24168
rect 29280 24008 29288 24072
rect 29352 24008 29360 24072
rect 29280 23912 29360 24008
rect 29280 23848 29288 23912
rect 29352 23848 29360 23912
rect 29280 23592 29360 23848
rect 29280 23528 29288 23592
rect 29352 23528 29360 23592
rect 29280 23272 29360 23528
rect 29280 23208 29288 23272
rect 29352 23208 29360 23272
rect 29280 23112 29360 23208
rect 29280 23048 29288 23112
rect 29352 23048 29360 23112
rect 29280 22952 29360 23048
rect 29280 22888 29288 22952
rect 29352 22888 29360 22952
rect 29280 22792 29360 22888
rect 29280 22728 29288 22792
rect 29352 22728 29360 22792
rect 29280 22632 29360 22728
rect 29280 22568 29288 22632
rect 29352 22568 29360 22632
rect 29280 22472 29360 22568
rect 29280 22408 29288 22472
rect 29352 22408 29360 22472
rect 29280 22312 29360 22408
rect 29280 22248 29288 22312
rect 29352 22248 29360 22312
rect 29280 22152 29360 22248
rect 29280 22088 29288 22152
rect 29352 22088 29360 22152
rect 29280 21992 29360 22088
rect 29280 21928 29288 21992
rect 29352 21928 29360 21992
rect 29280 21832 29360 21928
rect 29280 21768 29288 21832
rect 29352 21768 29360 21832
rect 29280 21672 29360 21768
rect 29280 21608 29288 21672
rect 29352 21608 29360 21672
rect 29280 21512 29360 21608
rect 29280 21448 29288 21512
rect 29352 21448 29360 21512
rect 29280 21352 29360 21448
rect 29280 21288 29288 21352
rect 29352 21288 29360 21352
rect 29280 21192 29360 21288
rect 29280 21128 29288 21192
rect 29352 21128 29360 21192
rect 29280 21032 29360 21128
rect 29280 20968 29288 21032
rect 29352 20968 29360 21032
rect 29280 20872 29360 20968
rect 29280 20808 29288 20872
rect 29352 20808 29360 20872
rect 29280 20712 29360 20808
rect 29280 20648 29288 20712
rect 29352 20648 29360 20712
rect 29280 20552 29360 20648
rect 29280 20488 29288 20552
rect 29352 20488 29360 20552
rect 29280 20392 29360 20488
rect 29280 20328 29288 20392
rect 29352 20328 29360 20392
rect 29280 20232 29360 20328
rect 29280 20168 29288 20232
rect 29352 20168 29360 20232
rect 29280 20072 29360 20168
rect 29280 20008 29288 20072
rect 29352 20008 29360 20072
rect 29280 19912 29360 20008
rect 29280 19848 29288 19912
rect 29352 19848 29360 19912
rect 29280 19752 29360 19848
rect 29280 19688 29288 19752
rect 29352 19688 29360 19752
rect 29280 19592 29360 19688
rect 29280 19528 29288 19592
rect 29352 19528 29360 19592
rect 29280 19432 29360 19528
rect 29280 19368 29288 19432
rect 29352 19368 29360 19432
rect 29280 19272 29360 19368
rect 29280 19208 29288 19272
rect 29352 19208 29360 19272
rect 29280 19112 29360 19208
rect 29280 19048 29288 19112
rect 29352 19048 29360 19112
rect 29280 18952 29360 19048
rect 29280 18888 29288 18952
rect 29352 18888 29360 18952
rect 29280 18792 29360 18888
rect 29280 18728 29288 18792
rect 29352 18728 29360 18792
rect 29280 18632 29360 18728
rect 29280 18568 29288 18632
rect 29352 18568 29360 18632
rect 29280 18472 29360 18568
rect 29280 18408 29288 18472
rect 29352 18408 29360 18472
rect 29280 18312 29360 18408
rect 29280 18248 29288 18312
rect 29352 18248 29360 18312
rect 29280 18152 29360 18248
rect 29280 18088 29288 18152
rect 29352 18088 29360 18152
rect 29280 17992 29360 18088
rect 29280 17928 29288 17992
rect 29352 17928 29360 17992
rect 29280 17832 29360 17928
rect 29280 17768 29288 17832
rect 29352 17768 29360 17832
rect 29280 17672 29360 17768
rect 29280 17608 29288 17672
rect 29352 17608 29360 17672
rect 29280 17512 29360 17608
rect 29280 17448 29288 17512
rect 29352 17448 29360 17512
rect 29280 17352 29360 17448
rect 29280 17288 29288 17352
rect 29352 17288 29360 17352
rect 29280 17192 29360 17288
rect 29280 17128 29288 17192
rect 29352 17128 29360 17192
rect 29280 17032 29360 17128
rect 29280 16968 29288 17032
rect 29352 16968 29360 17032
rect 29280 16872 29360 16968
rect 29280 16808 29288 16872
rect 29352 16808 29360 16872
rect 29280 16712 29360 16808
rect 29280 16648 29288 16712
rect 29352 16648 29360 16712
rect 29280 16552 29360 16648
rect 29280 16488 29288 16552
rect 29352 16488 29360 16552
rect 29280 16392 29360 16488
rect 29280 16328 29288 16392
rect 29352 16328 29360 16392
rect 29280 16232 29360 16328
rect 29280 16168 29288 16232
rect 29352 16168 29360 16232
rect 29280 16072 29360 16168
rect 29280 16008 29288 16072
rect 29352 16008 29360 16072
rect 29280 15912 29360 16008
rect 29280 15848 29288 15912
rect 29352 15848 29360 15912
rect 29280 15752 29360 15848
rect 29280 15688 29288 15752
rect 29352 15688 29360 15752
rect 29280 15592 29360 15688
rect 29280 15528 29288 15592
rect 29352 15528 29360 15592
rect 29280 15432 29360 15528
rect 29280 15368 29288 15432
rect 29352 15368 29360 15432
rect 29280 15272 29360 15368
rect 29280 15208 29288 15272
rect 29352 15208 29360 15272
rect 29280 15112 29360 15208
rect 29280 15048 29288 15112
rect 29352 15048 29360 15112
rect 29280 14952 29360 15048
rect 29280 14888 29288 14952
rect 29352 14888 29360 14952
rect 29280 14792 29360 14888
rect 29280 14728 29288 14792
rect 29352 14728 29360 14792
rect 29280 14632 29360 14728
rect 29280 14568 29288 14632
rect 29352 14568 29360 14632
rect 29280 14472 29360 14568
rect 29280 14408 29288 14472
rect 29352 14408 29360 14472
rect 29280 14312 29360 14408
rect 29280 14248 29288 14312
rect 29352 14248 29360 14312
rect 29280 14152 29360 14248
rect 29280 14088 29288 14152
rect 29352 14088 29360 14152
rect 29280 13992 29360 14088
rect 29280 13928 29288 13992
rect 29352 13928 29360 13992
rect 29280 13832 29360 13928
rect 29280 13768 29288 13832
rect 29352 13768 29360 13832
rect 29280 13672 29360 13768
rect 29280 13608 29288 13672
rect 29352 13608 29360 13672
rect 29280 13512 29360 13608
rect 29280 13448 29288 13512
rect 29352 13448 29360 13512
rect 29280 13352 29360 13448
rect 29280 13288 29288 13352
rect 29352 13288 29360 13352
rect 29280 13192 29360 13288
rect 29280 13128 29288 13192
rect 29352 13128 29360 13192
rect 29280 13032 29360 13128
rect 29280 12968 29288 13032
rect 29352 12968 29360 13032
rect 29280 12872 29360 12968
rect 29280 12808 29288 12872
rect 29352 12808 29360 12872
rect 29280 12712 29360 12808
rect 29280 12648 29288 12712
rect 29352 12648 29360 12712
rect 29280 12552 29360 12648
rect 29280 12488 29288 12552
rect 29352 12488 29360 12552
rect 29280 12392 29360 12488
rect 29280 12328 29288 12392
rect 29352 12328 29360 12392
rect 29280 12232 29360 12328
rect 29280 12168 29288 12232
rect 29352 12168 29360 12232
rect 29280 12072 29360 12168
rect 29280 12008 29288 12072
rect 29352 12008 29360 12072
rect 29280 11912 29360 12008
rect 29280 11848 29288 11912
rect 29352 11848 29360 11912
rect 29280 11752 29360 11848
rect 29280 11688 29288 11752
rect 29352 11688 29360 11752
rect 29280 11592 29360 11688
rect 29280 11528 29288 11592
rect 29352 11528 29360 11592
rect 29280 11432 29360 11528
rect 29280 11368 29288 11432
rect 29352 11368 29360 11432
rect 29280 11272 29360 11368
rect 29280 11208 29288 11272
rect 29352 11208 29360 11272
rect 29280 11112 29360 11208
rect 29280 11048 29288 11112
rect 29352 11048 29360 11112
rect 29280 10952 29360 11048
rect 29280 10888 29288 10952
rect 29352 10888 29360 10952
rect 29280 10792 29360 10888
rect 29280 10728 29288 10792
rect 29352 10728 29360 10792
rect 29280 10632 29360 10728
rect 29280 10568 29288 10632
rect 29352 10568 29360 10632
rect 29280 10472 29360 10568
rect 29280 10408 29288 10472
rect 29352 10408 29360 10472
rect 29280 10312 29360 10408
rect 29280 10248 29288 10312
rect 29352 10248 29360 10312
rect 29280 10152 29360 10248
rect 29280 10088 29288 10152
rect 29352 10088 29360 10152
rect 29280 9992 29360 10088
rect 29280 9928 29288 9992
rect 29352 9928 29360 9992
rect 29280 9832 29360 9928
rect 29280 9768 29288 9832
rect 29352 9768 29360 9832
rect 29280 9672 29360 9768
rect 29280 9608 29288 9672
rect 29352 9608 29360 9672
rect 29280 9352 29360 9608
rect 29280 9288 29288 9352
rect 29352 9288 29360 9352
rect 29280 9032 29360 9288
rect 29280 8968 29288 9032
rect 29352 8968 29360 9032
rect 29280 8872 29360 8968
rect 29280 8808 29288 8872
rect 29352 8808 29360 8872
rect 29280 8712 29360 8808
rect 29280 8648 29288 8712
rect 29352 8648 29360 8712
rect 29280 8552 29360 8648
rect 29280 8488 29288 8552
rect 29352 8488 29360 8552
rect 29280 8392 29360 8488
rect 29280 8328 29288 8392
rect 29352 8328 29360 8392
rect 29280 8232 29360 8328
rect 29280 8168 29288 8232
rect 29352 8168 29360 8232
rect 29280 8072 29360 8168
rect 29280 8008 29288 8072
rect 29352 8008 29360 8072
rect 29280 7912 29360 8008
rect 29280 7848 29288 7912
rect 29352 7848 29360 7912
rect 29280 7752 29360 7848
rect 29280 7688 29288 7752
rect 29352 7688 29360 7752
rect 29280 7592 29360 7688
rect 29280 7528 29288 7592
rect 29352 7528 29360 7592
rect 29280 7432 29360 7528
rect 29280 7368 29288 7432
rect 29352 7368 29360 7432
rect 29280 7272 29360 7368
rect 29280 7208 29288 7272
rect 29352 7208 29360 7272
rect 29280 7112 29360 7208
rect 29280 7048 29288 7112
rect 29352 7048 29360 7112
rect 29280 6952 29360 7048
rect 29280 6888 29288 6952
rect 29352 6888 29360 6952
rect 29280 6792 29360 6888
rect 29280 6728 29288 6792
rect 29352 6728 29360 6792
rect 29280 6632 29360 6728
rect 29280 6568 29288 6632
rect 29352 6568 29360 6632
rect 29280 6472 29360 6568
rect 29280 6408 29288 6472
rect 29352 6408 29360 6472
rect 29280 6312 29360 6408
rect 29280 6248 29288 6312
rect 29352 6248 29360 6312
rect 29280 6152 29360 6248
rect 29280 6088 29288 6152
rect 29352 6088 29360 6152
rect 29280 5992 29360 6088
rect 29280 5928 29288 5992
rect 29352 5928 29360 5992
rect 29280 5832 29360 5928
rect 29280 5768 29288 5832
rect 29352 5768 29360 5832
rect 29280 5672 29360 5768
rect 29280 5608 29288 5672
rect 29352 5608 29360 5672
rect 29280 5512 29360 5608
rect 29280 5448 29288 5512
rect 29352 5448 29360 5512
rect 29280 5352 29360 5448
rect 29280 5288 29288 5352
rect 29352 5288 29360 5352
rect 29280 5192 29360 5288
rect 29280 5128 29288 5192
rect 29352 5128 29360 5192
rect 29280 5032 29360 5128
rect 29280 4968 29288 5032
rect 29352 4968 29360 5032
rect 29280 4872 29360 4968
rect 29280 4808 29288 4872
rect 29352 4808 29360 4872
rect 29280 4712 29360 4808
rect 29280 4648 29288 4712
rect 29352 4648 29360 4712
rect 29280 4552 29360 4648
rect 29280 4488 29288 4552
rect 29352 4488 29360 4552
rect 29280 4392 29360 4488
rect 29280 4328 29288 4392
rect 29352 4328 29360 4392
rect 29280 4232 29360 4328
rect 29280 4168 29288 4232
rect 29352 4168 29360 4232
rect 29280 3912 29360 4168
rect 29280 3848 29288 3912
rect 29352 3848 29360 3912
rect 29280 3592 29360 3848
rect 29280 3528 29288 3592
rect 29352 3528 29360 3592
rect 29280 3432 29360 3528
rect 29280 3368 29288 3432
rect 29352 3368 29360 3432
rect 29280 3272 29360 3368
rect 29280 3208 29288 3272
rect 29352 3208 29360 3272
rect 29280 3112 29360 3208
rect 29280 3048 29288 3112
rect 29352 3048 29360 3112
rect 29280 2952 29360 3048
rect 29280 2888 29288 2952
rect 29352 2888 29360 2952
rect 29280 2792 29360 2888
rect 29280 2728 29288 2792
rect 29352 2728 29360 2792
rect 29280 2632 29360 2728
rect 29280 2568 29288 2632
rect 29352 2568 29360 2632
rect 29280 2472 29360 2568
rect 29280 2408 29288 2472
rect 29352 2408 29360 2472
rect 29280 2312 29360 2408
rect 29280 2248 29288 2312
rect 29352 2248 29360 2312
rect 29280 2152 29360 2248
rect 29280 2088 29288 2152
rect 29352 2088 29360 2152
rect 29280 1992 29360 2088
rect 29280 1928 29288 1992
rect 29352 1928 29360 1992
rect 29280 1832 29360 1928
rect 29280 1768 29288 1832
rect 29352 1768 29360 1832
rect 29280 1672 29360 1768
rect 29280 1608 29288 1672
rect 29352 1608 29360 1672
rect 29280 1512 29360 1608
rect 29280 1448 29288 1512
rect 29352 1448 29360 1512
rect 29280 1352 29360 1448
rect 29280 1288 29288 1352
rect 29352 1288 29360 1352
rect 29280 1192 29360 1288
rect 29280 1128 29288 1192
rect 29352 1128 29360 1192
rect 29280 1032 29360 1128
rect 29280 968 29288 1032
rect 29352 968 29360 1032
rect 28960 808 28968 872
rect 29032 808 29040 872
rect 28960 792 29040 808
rect 28960 728 28968 792
rect 29032 728 29040 792
rect 28960 712 29040 728
rect 28960 648 28968 712
rect 29032 648 29040 712
rect 28960 632 29040 648
rect 28960 568 28968 632
rect 29032 568 29040 632
rect 28960 552 29040 568
rect 28960 488 28968 552
rect 29032 488 29040 552
rect 28960 480 29040 488
rect 29280 872 29360 968
rect 29440 28872 29520 31920
rect 29440 28808 29448 28872
rect 29512 28808 29520 28872
rect 29440 23752 29520 28808
rect 29440 23688 29448 23752
rect 29512 23688 29520 23752
rect 29440 9192 29520 23688
rect 29440 9128 29448 9192
rect 29512 9128 29520 9192
rect 29440 4072 29520 9128
rect 29440 4008 29448 4072
rect 29512 4008 29520 4072
rect 29440 960 29520 4008
rect 29600 31912 29680 31920
rect 29600 31848 29608 31912
rect 29672 31848 29680 31912
rect 29600 31752 29680 31848
rect 29600 31688 29608 31752
rect 29672 31688 29680 31752
rect 29600 31592 29680 31688
rect 29600 31528 29608 31592
rect 29672 31528 29680 31592
rect 29600 31432 29680 31528
rect 29600 31368 29608 31432
rect 29672 31368 29680 31432
rect 29600 31272 29680 31368
rect 29600 31208 29608 31272
rect 29672 31208 29680 31272
rect 29600 31112 29680 31208
rect 29600 31048 29608 31112
rect 29672 31048 29680 31112
rect 29600 30952 29680 31048
rect 29600 30888 29608 30952
rect 29672 30888 29680 30952
rect 29600 30792 29680 30888
rect 29600 30728 29608 30792
rect 29672 30728 29680 30792
rect 29600 30632 29680 30728
rect 29600 30568 29608 30632
rect 29672 30568 29680 30632
rect 29600 30472 29680 30568
rect 29600 30408 29608 30472
rect 29672 30408 29680 30472
rect 29600 30312 29680 30408
rect 29600 30248 29608 30312
rect 29672 30248 29680 30312
rect 29600 30152 29680 30248
rect 29600 30088 29608 30152
rect 29672 30088 29680 30152
rect 29600 29992 29680 30088
rect 29600 29928 29608 29992
rect 29672 29928 29680 29992
rect 29600 29832 29680 29928
rect 29600 29768 29608 29832
rect 29672 29768 29680 29832
rect 29600 29672 29680 29768
rect 29600 29608 29608 29672
rect 29672 29608 29680 29672
rect 29600 29512 29680 29608
rect 29600 29448 29608 29512
rect 29672 29448 29680 29512
rect 29600 29352 29680 29448
rect 29600 29288 29608 29352
rect 29672 29288 29680 29352
rect 29600 29032 29680 29288
rect 29600 28968 29608 29032
rect 29672 28968 29680 29032
rect 29600 28872 29680 28968
rect 29600 28808 29608 28872
rect 29672 28808 29680 28872
rect 29600 28712 29680 28808
rect 29600 28648 29608 28712
rect 29672 28648 29680 28712
rect 29600 28552 29680 28648
rect 29600 28488 29608 28552
rect 29672 28488 29680 28552
rect 29600 28392 29680 28488
rect 29600 28328 29608 28392
rect 29672 28328 29680 28392
rect 29600 28232 29680 28328
rect 29600 28168 29608 28232
rect 29672 28168 29680 28232
rect 29600 28072 29680 28168
rect 29600 28008 29608 28072
rect 29672 28008 29680 28072
rect 29600 27912 29680 28008
rect 29600 27848 29608 27912
rect 29672 27848 29680 27912
rect 29600 27752 29680 27848
rect 29600 27688 29608 27752
rect 29672 27688 29680 27752
rect 29600 27592 29680 27688
rect 29600 27528 29608 27592
rect 29672 27528 29680 27592
rect 29600 27432 29680 27528
rect 29600 27368 29608 27432
rect 29672 27368 29680 27432
rect 29600 27272 29680 27368
rect 29600 27208 29608 27272
rect 29672 27208 29680 27272
rect 29600 27112 29680 27208
rect 29600 27048 29608 27112
rect 29672 27048 29680 27112
rect 29600 26952 29680 27048
rect 29600 26888 29608 26952
rect 29672 26888 29680 26952
rect 29600 26792 29680 26888
rect 29600 26728 29608 26792
rect 29672 26728 29680 26792
rect 29600 26632 29680 26728
rect 29600 26568 29608 26632
rect 29672 26568 29680 26632
rect 29600 26472 29680 26568
rect 29600 26408 29608 26472
rect 29672 26408 29680 26472
rect 29600 26312 29680 26408
rect 29600 26248 29608 26312
rect 29672 26248 29680 26312
rect 29600 26152 29680 26248
rect 29600 26088 29608 26152
rect 29672 26088 29680 26152
rect 29600 25992 29680 26088
rect 29600 25928 29608 25992
rect 29672 25928 29680 25992
rect 29600 25832 29680 25928
rect 29600 25768 29608 25832
rect 29672 25768 29680 25832
rect 29600 25672 29680 25768
rect 29600 25608 29608 25672
rect 29672 25608 29680 25672
rect 29600 25512 29680 25608
rect 29600 25448 29608 25512
rect 29672 25448 29680 25512
rect 29600 25352 29680 25448
rect 29600 25288 29608 25352
rect 29672 25288 29680 25352
rect 29600 25192 29680 25288
rect 29600 25128 29608 25192
rect 29672 25128 29680 25192
rect 29600 25032 29680 25128
rect 29600 24968 29608 25032
rect 29672 24968 29680 25032
rect 29600 24872 29680 24968
rect 29600 24808 29608 24872
rect 29672 24808 29680 24872
rect 29600 24712 29680 24808
rect 29600 24648 29608 24712
rect 29672 24648 29680 24712
rect 29600 24552 29680 24648
rect 29600 24488 29608 24552
rect 29672 24488 29680 24552
rect 29600 24392 29680 24488
rect 29600 24328 29608 24392
rect 29672 24328 29680 24392
rect 29600 24232 29680 24328
rect 29600 24168 29608 24232
rect 29672 24168 29680 24232
rect 29600 24072 29680 24168
rect 29600 24008 29608 24072
rect 29672 24008 29680 24072
rect 29600 23912 29680 24008
rect 29600 23848 29608 23912
rect 29672 23848 29680 23912
rect 29600 23752 29680 23848
rect 29600 23688 29608 23752
rect 29672 23688 29680 23752
rect 29600 23592 29680 23688
rect 29600 23528 29608 23592
rect 29672 23528 29680 23592
rect 29600 23272 29680 23528
rect 29600 23208 29608 23272
rect 29672 23208 29680 23272
rect 29600 23112 29680 23208
rect 29600 23048 29608 23112
rect 29672 23048 29680 23112
rect 29600 22952 29680 23048
rect 29600 22888 29608 22952
rect 29672 22888 29680 22952
rect 29600 22792 29680 22888
rect 29600 22728 29608 22792
rect 29672 22728 29680 22792
rect 29600 22632 29680 22728
rect 29600 22568 29608 22632
rect 29672 22568 29680 22632
rect 29600 22472 29680 22568
rect 29600 22408 29608 22472
rect 29672 22408 29680 22472
rect 29600 22312 29680 22408
rect 29600 22248 29608 22312
rect 29672 22248 29680 22312
rect 29600 22152 29680 22248
rect 29600 22088 29608 22152
rect 29672 22088 29680 22152
rect 29600 21992 29680 22088
rect 29600 21928 29608 21992
rect 29672 21928 29680 21992
rect 29600 21832 29680 21928
rect 29600 21768 29608 21832
rect 29672 21768 29680 21832
rect 29600 21672 29680 21768
rect 29600 21608 29608 21672
rect 29672 21608 29680 21672
rect 29600 21512 29680 21608
rect 29600 21448 29608 21512
rect 29672 21448 29680 21512
rect 29600 21352 29680 21448
rect 29600 21288 29608 21352
rect 29672 21288 29680 21352
rect 29600 21192 29680 21288
rect 29600 21128 29608 21192
rect 29672 21128 29680 21192
rect 29600 21032 29680 21128
rect 29600 20968 29608 21032
rect 29672 20968 29680 21032
rect 29600 20872 29680 20968
rect 29600 20808 29608 20872
rect 29672 20808 29680 20872
rect 29600 20712 29680 20808
rect 29600 20648 29608 20712
rect 29672 20648 29680 20712
rect 29600 20552 29680 20648
rect 29600 20488 29608 20552
rect 29672 20488 29680 20552
rect 29600 20392 29680 20488
rect 29600 20328 29608 20392
rect 29672 20328 29680 20392
rect 29600 20232 29680 20328
rect 29600 20168 29608 20232
rect 29672 20168 29680 20232
rect 29600 20072 29680 20168
rect 29600 20008 29608 20072
rect 29672 20008 29680 20072
rect 29600 19912 29680 20008
rect 29600 19848 29608 19912
rect 29672 19848 29680 19912
rect 29600 19752 29680 19848
rect 29600 19688 29608 19752
rect 29672 19688 29680 19752
rect 29600 19592 29680 19688
rect 29600 19528 29608 19592
rect 29672 19528 29680 19592
rect 29600 19432 29680 19528
rect 29600 19368 29608 19432
rect 29672 19368 29680 19432
rect 29600 19272 29680 19368
rect 29600 19208 29608 19272
rect 29672 19208 29680 19272
rect 29600 19112 29680 19208
rect 29600 19048 29608 19112
rect 29672 19048 29680 19112
rect 29600 18952 29680 19048
rect 29600 18888 29608 18952
rect 29672 18888 29680 18952
rect 29600 18792 29680 18888
rect 29600 18728 29608 18792
rect 29672 18728 29680 18792
rect 29600 18632 29680 18728
rect 29600 18568 29608 18632
rect 29672 18568 29680 18632
rect 29600 18472 29680 18568
rect 29600 18408 29608 18472
rect 29672 18408 29680 18472
rect 29600 18312 29680 18408
rect 29600 18248 29608 18312
rect 29672 18248 29680 18312
rect 29600 18152 29680 18248
rect 29600 18088 29608 18152
rect 29672 18088 29680 18152
rect 29600 17992 29680 18088
rect 29600 17928 29608 17992
rect 29672 17928 29680 17992
rect 29600 17832 29680 17928
rect 29600 17768 29608 17832
rect 29672 17768 29680 17832
rect 29600 17672 29680 17768
rect 29600 17608 29608 17672
rect 29672 17608 29680 17672
rect 29600 17512 29680 17608
rect 29600 17448 29608 17512
rect 29672 17448 29680 17512
rect 29600 17352 29680 17448
rect 29600 17288 29608 17352
rect 29672 17288 29680 17352
rect 29600 17192 29680 17288
rect 29600 17128 29608 17192
rect 29672 17128 29680 17192
rect 29600 17032 29680 17128
rect 29600 16968 29608 17032
rect 29672 16968 29680 17032
rect 29600 16872 29680 16968
rect 29600 16808 29608 16872
rect 29672 16808 29680 16872
rect 29600 16712 29680 16808
rect 29600 16648 29608 16712
rect 29672 16648 29680 16712
rect 29600 16552 29680 16648
rect 29600 16488 29608 16552
rect 29672 16488 29680 16552
rect 29600 16392 29680 16488
rect 29600 16328 29608 16392
rect 29672 16328 29680 16392
rect 29600 16232 29680 16328
rect 29600 16168 29608 16232
rect 29672 16168 29680 16232
rect 29600 16072 29680 16168
rect 29600 16008 29608 16072
rect 29672 16008 29680 16072
rect 29600 15912 29680 16008
rect 29600 15848 29608 15912
rect 29672 15848 29680 15912
rect 29600 15752 29680 15848
rect 29600 15688 29608 15752
rect 29672 15688 29680 15752
rect 29600 15592 29680 15688
rect 29600 15528 29608 15592
rect 29672 15528 29680 15592
rect 29600 15432 29680 15528
rect 29600 15368 29608 15432
rect 29672 15368 29680 15432
rect 29600 15272 29680 15368
rect 29600 15208 29608 15272
rect 29672 15208 29680 15272
rect 29600 15112 29680 15208
rect 29600 15048 29608 15112
rect 29672 15048 29680 15112
rect 29600 14952 29680 15048
rect 29600 14888 29608 14952
rect 29672 14888 29680 14952
rect 29600 14792 29680 14888
rect 29600 14728 29608 14792
rect 29672 14728 29680 14792
rect 29600 14632 29680 14728
rect 29600 14568 29608 14632
rect 29672 14568 29680 14632
rect 29600 14472 29680 14568
rect 29600 14408 29608 14472
rect 29672 14408 29680 14472
rect 29600 14312 29680 14408
rect 29600 14248 29608 14312
rect 29672 14248 29680 14312
rect 29600 14152 29680 14248
rect 29600 14088 29608 14152
rect 29672 14088 29680 14152
rect 29600 13992 29680 14088
rect 29600 13928 29608 13992
rect 29672 13928 29680 13992
rect 29600 13832 29680 13928
rect 29600 13768 29608 13832
rect 29672 13768 29680 13832
rect 29600 13672 29680 13768
rect 29600 13608 29608 13672
rect 29672 13608 29680 13672
rect 29600 13512 29680 13608
rect 29600 13448 29608 13512
rect 29672 13448 29680 13512
rect 29600 13352 29680 13448
rect 29600 13288 29608 13352
rect 29672 13288 29680 13352
rect 29600 13192 29680 13288
rect 29600 13128 29608 13192
rect 29672 13128 29680 13192
rect 29600 13032 29680 13128
rect 29600 12968 29608 13032
rect 29672 12968 29680 13032
rect 29600 12872 29680 12968
rect 29600 12808 29608 12872
rect 29672 12808 29680 12872
rect 29600 12712 29680 12808
rect 29600 12648 29608 12712
rect 29672 12648 29680 12712
rect 29600 12552 29680 12648
rect 29600 12488 29608 12552
rect 29672 12488 29680 12552
rect 29600 12392 29680 12488
rect 29600 12328 29608 12392
rect 29672 12328 29680 12392
rect 29600 12232 29680 12328
rect 29600 12168 29608 12232
rect 29672 12168 29680 12232
rect 29600 12072 29680 12168
rect 29600 12008 29608 12072
rect 29672 12008 29680 12072
rect 29600 11912 29680 12008
rect 29600 11848 29608 11912
rect 29672 11848 29680 11912
rect 29600 11752 29680 11848
rect 29600 11688 29608 11752
rect 29672 11688 29680 11752
rect 29600 11592 29680 11688
rect 29600 11528 29608 11592
rect 29672 11528 29680 11592
rect 29600 11432 29680 11528
rect 29600 11368 29608 11432
rect 29672 11368 29680 11432
rect 29600 11272 29680 11368
rect 29600 11208 29608 11272
rect 29672 11208 29680 11272
rect 29600 11112 29680 11208
rect 29600 11048 29608 11112
rect 29672 11048 29680 11112
rect 29600 10952 29680 11048
rect 29600 10888 29608 10952
rect 29672 10888 29680 10952
rect 29600 10792 29680 10888
rect 29600 10728 29608 10792
rect 29672 10728 29680 10792
rect 29600 10632 29680 10728
rect 29600 10568 29608 10632
rect 29672 10568 29680 10632
rect 29600 10472 29680 10568
rect 29600 10408 29608 10472
rect 29672 10408 29680 10472
rect 29600 10312 29680 10408
rect 29600 10248 29608 10312
rect 29672 10248 29680 10312
rect 29600 10152 29680 10248
rect 29600 10088 29608 10152
rect 29672 10088 29680 10152
rect 29600 9992 29680 10088
rect 29600 9928 29608 9992
rect 29672 9928 29680 9992
rect 29600 9832 29680 9928
rect 29600 9768 29608 9832
rect 29672 9768 29680 9832
rect 29600 9672 29680 9768
rect 29600 9608 29608 9672
rect 29672 9608 29680 9672
rect 29600 9352 29680 9608
rect 29600 9288 29608 9352
rect 29672 9288 29680 9352
rect 29600 9192 29680 9288
rect 29600 9128 29608 9192
rect 29672 9128 29680 9192
rect 29600 9032 29680 9128
rect 29600 8968 29608 9032
rect 29672 8968 29680 9032
rect 29600 8872 29680 8968
rect 29600 8808 29608 8872
rect 29672 8808 29680 8872
rect 29600 8712 29680 8808
rect 29600 8648 29608 8712
rect 29672 8648 29680 8712
rect 29600 8552 29680 8648
rect 29600 8488 29608 8552
rect 29672 8488 29680 8552
rect 29600 8392 29680 8488
rect 29600 8328 29608 8392
rect 29672 8328 29680 8392
rect 29600 8232 29680 8328
rect 29600 8168 29608 8232
rect 29672 8168 29680 8232
rect 29600 8072 29680 8168
rect 29600 8008 29608 8072
rect 29672 8008 29680 8072
rect 29600 7912 29680 8008
rect 29600 7848 29608 7912
rect 29672 7848 29680 7912
rect 29600 7752 29680 7848
rect 29600 7688 29608 7752
rect 29672 7688 29680 7752
rect 29600 7592 29680 7688
rect 29600 7528 29608 7592
rect 29672 7528 29680 7592
rect 29600 7432 29680 7528
rect 29600 7368 29608 7432
rect 29672 7368 29680 7432
rect 29600 7272 29680 7368
rect 29600 7208 29608 7272
rect 29672 7208 29680 7272
rect 29600 7112 29680 7208
rect 29600 7048 29608 7112
rect 29672 7048 29680 7112
rect 29600 6952 29680 7048
rect 29600 6888 29608 6952
rect 29672 6888 29680 6952
rect 29600 6792 29680 6888
rect 29600 6728 29608 6792
rect 29672 6728 29680 6792
rect 29600 6632 29680 6728
rect 29600 6568 29608 6632
rect 29672 6568 29680 6632
rect 29600 6472 29680 6568
rect 29600 6408 29608 6472
rect 29672 6408 29680 6472
rect 29600 6312 29680 6408
rect 29600 6248 29608 6312
rect 29672 6248 29680 6312
rect 29600 6152 29680 6248
rect 29600 6088 29608 6152
rect 29672 6088 29680 6152
rect 29600 5992 29680 6088
rect 29600 5928 29608 5992
rect 29672 5928 29680 5992
rect 29600 5832 29680 5928
rect 29600 5768 29608 5832
rect 29672 5768 29680 5832
rect 29600 5672 29680 5768
rect 29600 5608 29608 5672
rect 29672 5608 29680 5672
rect 29600 5512 29680 5608
rect 29600 5448 29608 5512
rect 29672 5448 29680 5512
rect 29600 5352 29680 5448
rect 29600 5288 29608 5352
rect 29672 5288 29680 5352
rect 29600 5192 29680 5288
rect 29600 5128 29608 5192
rect 29672 5128 29680 5192
rect 29600 5032 29680 5128
rect 29600 4968 29608 5032
rect 29672 4968 29680 5032
rect 29600 4872 29680 4968
rect 29600 4808 29608 4872
rect 29672 4808 29680 4872
rect 29600 4712 29680 4808
rect 29600 4648 29608 4712
rect 29672 4648 29680 4712
rect 29600 4552 29680 4648
rect 29600 4488 29608 4552
rect 29672 4488 29680 4552
rect 29600 4392 29680 4488
rect 29600 4328 29608 4392
rect 29672 4328 29680 4392
rect 29600 4232 29680 4328
rect 29600 4168 29608 4232
rect 29672 4168 29680 4232
rect 29600 4072 29680 4168
rect 29600 4008 29608 4072
rect 29672 4008 29680 4072
rect 29600 3912 29680 4008
rect 29600 3848 29608 3912
rect 29672 3848 29680 3912
rect 29600 3592 29680 3848
rect 29600 3528 29608 3592
rect 29672 3528 29680 3592
rect 29600 3432 29680 3528
rect 29600 3368 29608 3432
rect 29672 3368 29680 3432
rect 29600 3272 29680 3368
rect 29600 3208 29608 3272
rect 29672 3208 29680 3272
rect 29600 3112 29680 3208
rect 29600 3048 29608 3112
rect 29672 3048 29680 3112
rect 29600 2952 29680 3048
rect 29600 2888 29608 2952
rect 29672 2888 29680 2952
rect 29600 2792 29680 2888
rect 29600 2728 29608 2792
rect 29672 2728 29680 2792
rect 29600 2632 29680 2728
rect 29600 2568 29608 2632
rect 29672 2568 29680 2632
rect 29600 2472 29680 2568
rect 29600 2408 29608 2472
rect 29672 2408 29680 2472
rect 29600 2312 29680 2408
rect 29600 2248 29608 2312
rect 29672 2248 29680 2312
rect 29600 2152 29680 2248
rect 29600 2088 29608 2152
rect 29672 2088 29680 2152
rect 29600 1992 29680 2088
rect 29600 1928 29608 1992
rect 29672 1928 29680 1992
rect 29600 1832 29680 1928
rect 29600 1768 29608 1832
rect 29672 1768 29680 1832
rect 29600 1672 29680 1768
rect 29600 1608 29608 1672
rect 29672 1608 29680 1672
rect 29600 1512 29680 1608
rect 29600 1448 29608 1512
rect 29672 1448 29680 1512
rect 29600 1352 29680 1448
rect 29600 1288 29608 1352
rect 29672 1288 29680 1352
rect 29600 1192 29680 1288
rect 29600 1128 29608 1192
rect 29672 1128 29680 1192
rect 29600 1032 29680 1128
rect 29600 968 29608 1032
rect 29672 968 29680 1032
rect 29280 808 29288 872
rect 29352 808 29360 872
rect 29280 792 29360 808
rect 29280 728 29288 792
rect 29352 728 29360 792
rect 29280 712 29360 728
rect 29280 648 29288 712
rect 29352 648 29360 712
rect 29280 632 29360 648
rect 29280 568 29288 632
rect 29352 568 29360 632
rect 29280 552 29360 568
rect 29280 488 29288 552
rect 29352 488 29360 552
rect 29280 480 29360 488
rect 29600 872 29680 968
rect 29760 29192 29840 31920
rect 29760 29128 29768 29192
rect 29832 29128 29840 29192
rect 29760 23432 29840 29128
rect 29760 23368 29768 23432
rect 29832 23368 29840 23432
rect 29760 9512 29840 23368
rect 29760 9448 29768 9512
rect 29832 9448 29840 9512
rect 29760 3752 29840 9448
rect 29760 3688 29768 3752
rect 29832 3688 29840 3752
rect 29760 960 29840 3688
rect 29920 31912 30000 31920
rect 29920 31848 29928 31912
rect 29992 31848 30000 31912
rect 29920 31752 30000 31848
rect 29920 31688 29928 31752
rect 29992 31688 30000 31752
rect 29920 31592 30000 31688
rect 29920 31528 29928 31592
rect 29992 31528 30000 31592
rect 29920 31432 30000 31528
rect 29920 31368 29928 31432
rect 29992 31368 30000 31432
rect 29920 31272 30000 31368
rect 29920 31208 29928 31272
rect 29992 31208 30000 31272
rect 29920 31112 30000 31208
rect 29920 31048 29928 31112
rect 29992 31048 30000 31112
rect 29920 30952 30000 31048
rect 29920 30888 29928 30952
rect 29992 30888 30000 30952
rect 29920 30792 30000 30888
rect 29920 30728 29928 30792
rect 29992 30728 30000 30792
rect 29920 30632 30000 30728
rect 29920 30568 29928 30632
rect 29992 30568 30000 30632
rect 29920 30472 30000 30568
rect 29920 30408 29928 30472
rect 29992 30408 30000 30472
rect 29920 30312 30000 30408
rect 29920 30248 29928 30312
rect 29992 30248 30000 30312
rect 29920 30152 30000 30248
rect 29920 30088 29928 30152
rect 29992 30088 30000 30152
rect 29920 29992 30000 30088
rect 29920 29928 29928 29992
rect 29992 29928 30000 29992
rect 29920 29832 30000 29928
rect 29920 29768 29928 29832
rect 29992 29768 30000 29832
rect 29920 29672 30000 29768
rect 29920 29608 29928 29672
rect 29992 29608 30000 29672
rect 29920 29512 30000 29608
rect 29920 29448 29928 29512
rect 29992 29448 30000 29512
rect 29920 29352 30000 29448
rect 29920 29288 29928 29352
rect 29992 29288 30000 29352
rect 29920 29032 30000 29288
rect 29920 28968 29928 29032
rect 29992 28968 30000 29032
rect 29920 28872 30000 28968
rect 29920 28808 29928 28872
rect 29992 28808 30000 28872
rect 29920 28712 30000 28808
rect 29920 28648 29928 28712
rect 29992 28648 30000 28712
rect 29920 28552 30000 28648
rect 29920 28488 29928 28552
rect 29992 28488 30000 28552
rect 29920 28392 30000 28488
rect 29920 28328 29928 28392
rect 29992 28328 30000 28392
rect 29920 28232 30000 28328
rect 29920 28168 29928 28232
rect 29992 28168 30000 28232
rect 29920 28072 30000 28168
rect 29920 28008 29928 28072
rect 29992 28008 30000 28072
rect 29920 27912 30000 28008
rect 29920 27848 29928 27912
rect 29992 27848 30000 27912
rect 29920 27752 30000 27848
rect 29920 27688 29928 27752
rect 29992 27688 30000 27752
rect 29920 27592 30000 27688
rect 29920 27528 29928 27592
rect 29992 27528 30000 27592
rect 29920 27432 30000 27528
rect 29920 27368 29928 27432
rect 29992 27368 30000 27432
rect 29920 27272 30000 27368
rect 29920 27208 29928 27272
rect 29992 27208 30000 27272
rect 29920 27112 30000 27208
rect 29920 27048 29928 27112
rect 29992 27048 30000 27112
rect 29920 26952 30000 27048
rect 29920 26888 29928 26952
rect 29992 26888 30000 26952
rect 29920 26792 30000 26888
rect 29920 26728 29928 26792
rect 29992 26728 30000 26792
rect 29920 26632 30000 26728
rect 29920 26568 29928 26632
rect 29992 26568 30000 26632
rect 29920 26472 30000 26568
rect 29920 26408 29928 26472
rect 29992 26408 30000 26472
rect 29920 26312 30000 26408
rect 29920 26248 29928 26312
rect 29992 26248 30000 26312
rect 29920 26152 30000 26248
rect 29920 26088 29928 26152
rect 29992 26088 30000 26152
rect 29920 25992 30000 26088
rect 29920 25928 29928 25992
rect 29992 25928 30000 25992
rect 29920 25832 30000 25928
rect 29920 25768 29928 25832
rect 29992 25768 30000 25832
rect 29920 25672 30000 25768
rect 29920 25608 29928 25672
rect 29992 25608 30000 25672
rect 29920 25512 30000 25608
rect 29920 25448 29928 25512
rect 29992 25448 30000 25512
rect 29920 25352 30000 25448
rect 29920 25288 29928 25352
rect 29992 25288 30000 25352
rect 29920 25192 30000 25288
rect 29920 25128 29928 25192
rect 29992 25128 30000 25192
rect 29920 25032 30000 25128
rect 29920 24968 29928 25032
rect 29992 24968 30000 25032
rect 29920 24872 30000 24968
rect 29920 24808 29928 24872
rect 29992 24808 30000 24872
rect 29920 24712 30000 24808
rect 29920 24648 29928 24712
rect 29992 24648 30000 24712
rect 29920 24552 30000 24648
rect 29920 24488 29928 24552
rect 29992 24488 30000 24552
rect 29920 24392 30000 24488
rect 29920 24328 29928 24392
rect 29992 24328 30000 24392
rect 29920 24232 30000 24328
rect 29920 24168 29928 24232
rect 29992 24168 30000 24232
rect 29920 24072 30000 24168
rect 29920 24008 29928 24072
rect 29992 24008 30000 24072
rect 29920 23912 30000 24008
rect 29920 23848 29928 23912
rect 29992 23848 30000 23912
rect 29920 23752 30000 23848
rect 29920 23688 29928 23752
rect 29992 23688 30000 23752
rect 29920 23592 30000 23688
rect 29920 23528 29928 23592
rect 29992 23528 30000 23592
rect 29920 23272 30000 23528
rect 29920 23208 29928 23272
rect 29992 23208 30000 23272
rect 29920 23112 30000 23208
rect 29920 23048 29928 23112
rect 29992 23048 30000 23112
rect 29920 22952 30000 23048
rect 29920 22888 29928 22952
rect 29992 22888 30000 22952
rect 29920 22792 30000 22888
rect 29920 22728 29928 22792
rect 29992 22728 30000 22792
rect 29920 22632 30000 22728
rect 29920 22568 29928 22632
rect 29992 22568 30000 22632
rect 29920 22472 30000 22568
rect 29920 22408 29928 22472
rect 29992 22408 30000 22472
rect 29920 22312 30000 22408
rect 29920 22248 29928 22312
rect 29992 22248 30000 22312
rect 29920 22152 30000 22248
rect 29920 22088 29928 22152
rect 29992 22088 30000 22152
rect 29920 21992 30000 22088
rect 29920 21928 29928 21992
rect 29992 21928 30000 21992
rect 29920 21832 30000 21928
rect 29920 21768 29928 21832
rect 29992 21768 30000 21832
rect 29920 21672 30000 21768
rect 29920 21608 29928 21672
rect 29992 21608 30000 21672
rect 29920 21512 30000 21608
rect 29920 21448 29928 21512
rect 29992 21448 30000 21512
rect 29920 21352 30000 21448
rect 29920 21288 29928 21352
rect 29992 21288 30000 21352
rect 29920 21192 30000 21288
rect 29920 21128 29928 21192
rect 29992 21128 30000 21192
rect 29920 21032 30000 21128
rect 29920 20968 29928 21032
rect 29992 20968 30000 21032
rect 29920 20872 30000 20968
rect 29920 20808 29928 20872
rect 29992 20808 30000 20872
rect 29920 20712 30000 20808
rect 29920 20648 29928 20712
rect 29992 20648 30000 20712
rect 29920 20552 30000 20648
rect 29920 20488 29928 20552
rect 29992 20488 30000 20552
rect 29920 20392 30000 20488
rect 29920 20328 29928 20392
rect 29992 20328 30000 20392
rect 29920 20232 30000 20328
rect 29920 20168 29928 20232
rect 29992 20168 30000 20232
rect 29920 20072 30000 20168
rect 29920 20008 29928 20072
rect 29992 20008 30000 20072
rect 29920 19912 30000 20008
rect 29920 19848 29928 19912
rect 29992 19848 30000 19912
rect 29920 19752 30000 19848
rect 29920 19688 29928 19752
rect 29992 19688 30000 19752
rect 29920 19592 30000 19688
rect 29920 19528 29928 19592
rect 29992 19528 30000 19592
rect 29920 19432 30000 19528
rect 29920 19368 29928 19432
rect 29992 19368 30000 19432
rect 29920 19272 30000 19368
rect 29920 19208 29928 19272
rect 29992 19208 30000 19272
rect 29920 19112 30000 19208
rect 29920 19048 29928 19112
rect 29992 19048 30000 19112
rect 29920 18952 30000 19048
rect 29920 18888 29928 18952
rect 29992 18888 30000 18952
rect 29920 18792 30000 18888
rect 29920 18728 29928 18792
rect 29992 18728 30000 18792
rect 29920 18632 30000 18728
rect 29920 18568 29928 18632
rect 29992 18568 30000 18632
rect 29920 18472 30000 18568
rect 29920 18408 29928 18472
rect 29992 18408 30000 18472
rect 29920 18312 30000 18408
rect 29920 18248 29928 18312
rect 29992 18248 30000 18312
rect 29920 18152 30000 18248
rect 29920 18088 29928 18152
rect 29992 18088 30000 18152
rect 29920 17992 30000 18088
rect 29920 17928 29928 17992
rect 29992 17928 30000 17992
rect 29920 17832 30000 17928
rect 29920 17768 29928 17832
rect 29992 17768 30000 17832
rect 29920 17672 30000 17768
rect 29920 17608 29928 17672
rect 29992 17608 30000 17672
rect 29920 17512 30000 17608
rect 29920 17448 29928 17512
rect 29992 17448 30000 17512
rect 29920 17352 30000 17448
rect 29920 17288 29928 17352
rect 29992 17288 30000 17352
rect 29920 17192 30000 17288
rect 29920 17128 29928 17192
rect 29992 17128 30000 17192
rect 29920 17032 30000 17128
rect 29920 16968 29928 17032
rect 29992 16968 30000 17032
rect 29920 16872 30000 16968
rect 29920 16808 29928 16872
rect 29992 16808 30000 16872
rect 29920 16712 30000 16808
rect 29920 16648 29928 16712
rect 29992 16648 30000 16712
rect 29920 16552 30000 16648
rect 29920 16488 29928 16552
rect 29992 16488 30000 16552
rect 29920 16392 30000 16488
rect 29920 16328 29928 16392
rect 29992 16328 30000 16392
rect 29920 16232 30000 16328
rect 29920 16168 29928 16232
rect 29992 16168 30000 16232
rect 29920 16072 30000 16168
rect 29920 16008 29928 16072
rect 29992 16008 30000 16072
rect 29920 15912 30000 16008
rect 29920 15848 29928 15912
rect 29992 15848 30000 15912
rect 29920 15752 30000 15848
rect 29920 15688 29928 15752
rect 29992 15688 30000 15752
rect 29920 15592 30000 15688
rect 29920 15528 29928 15592
rect 29992 15528 30000 15592
rect 29920 15432 30000 15528
rect 29920 15368 29928 15432
rect 29992 15368 30000 15432
rect 29920 15272 30000 15368
rect 29920 15208 29928 15272
rect 29992 15208 30000 15272
rect 29920 15112 30000 15208
rect 29920 15048 29928 15112
rect 29992 15048 30000 15112
rect 29920 14952 30000 15048
rect 29920 14888 29928 14952
rect 29992 14888 30000 14952
rect 29920 14792 30000 14888
rect 29920 14728 29928 14792
rect 29992 14728 30000 14792
rect 29920 14632 30000 14728
rect 29920 14568 29928 14632
rect 29992 14568 30000 14632
rect 29920 14472 30000 14568
rect 29920 14408 29928 14472
rect 29992 14408 30000 14472
rect 29920 14312 30000 14408
rect 29920 14248 29928 14312
rect 29992 14248 30000 14312
rect 29920 14152 30000 14248
rect 29920 14088 29928 14152
rect 29992 14088 30000 14152
rect 29920 13992 30000 14088
rect 29920 13928 29928 13992
rect 29992 13928 30000 13992
rect 29920 13832 30000 13928
rect 29920 13768 29928 13832
rect 29992 13768 30000 13832
rect 29920 13672 30000 13768
rect 29920 13608 29928 13672
rect 29992 13608 30000 13672
rect 29920 13512 30000 13608
rect 29920 13448 29928 13512
rect 29992 13448 30000 13512
rect 29920 13352 30000 13448
rect 29920 13288 29928 13352
rect 29992 13288 30000 13352
rect 29920 13192 30000 13288
rect 29920 13128 29928 13192
rect 29992 13128 30000 13192
rect 29920 13032 30000 13128
rect 29920 12968 29928 13032
rect 29992 12968 30000 13032
rect 29920 12872 30000 12968
rect 29920 12808 29928 12872
rect 29992 12808 30000 12872
rect 29920 12712 30000 12808
rect 29920 12648 29928 12712
rect 29992 12648 30000 12712
rect 29920 12552 30000 12648
rect 29920 12488 29928 12552
rect 29992 12488 30000 12552
rect 29920 12392 30000 12488
rect 29920 12328 29928 12392
rect 29992 12328 30000 12392
rect 29920 12232 30000 12328
rect 29920 12168 29928 12232
rect 29992 12168 30000 12232
rect 29920 12072 30000 12168
rect 29920 12008 29928 12072
rect 29992 12008 30000 12072
rect 29920 11912 30000 12008
rect 29920 11848 29928 11912
rect 29992 11848 30000 11912
rect 29920 11752 30000 11848
rect 29920 11688 29928 11752
rect 29992 11688 30000 11752
rect 29920 11592 30000 11688
rect 29920 11528 29928 11592
rect 29992 11528 30000 11592
rect 29920 11432 30000 11528
rect 29920 11368 29928 11432
rect 29992 11368 30000 11432
rect 29920 11272 30000 11368
rect 29920 11208 29928 11272
rect 29992 11208 30000 11272
rect 29920 11112 30000 11208
rect 29920 11048 29928 11112
rect 29992 11048 30000 11112
rect 29920 10952 30000 11048
rect 29920 10888 29928 10952
rect 29992 10888 30000 10952
rect 29920 10792 30000 10888
rect 29920 10728 29928 10792
rect 29992 10728 30000 10792
rect 29920 10632 30000 10728
rect 29920 10568 29928 10632
rect 29992 10568 30000 10632
rect 29920 10472 30000 10568
rect 29920 10408 29928 10472
rect 29992 10408 30000 10472
rect 29920 10312 30000 10408
rect 29920 10248 29928 10312
rect 29992 10248 30000 10312
rect 29920 10152 30000 10248
rect 29920 10088 29928 10152
rect 29992 10088 30000 10152
rect 29920 9992 30000 10088
rect 29920 9928 29928 9992
rect 29992 9928 30000 9992
rect 29920 9832 30000 9928
rect 29920 9768 29928 9832
rect 29992 9768 30000 9832
rect 29920 9672 30000 9768
rect 29920 9608 29928 9672
rect 29992 9608 30000 9672
rect 29920 9352 30000 9608
rect 29920 9288 29928 9352
rect 29992 9288 30000 9352
rect 29920 9192 30000 9288
rect 29920 9128 29928 9192
rect 29992 9128 30000 9192
rect 29920 9032 30000 9128
rect 29920 8968 29928 9032
rect 29992 8968 30000 9032
rect 29920 8872 30000 8968
rect 29920 8808 29928 8872
rect 29992 8808 30000 8872
rect 29920 8712 30000 8808
rect 29920 8648 29928 8712
rect 29992 8648 30000 8712
rect 29920 8552 30000 8648
rect 29920 8488 29928 8552
rect 29992 8488 30000 8552
rect 29920 8392 30000 8488
rect 29920 8328 29928 8392
rect 29992 8328 30000 8392
rect 29920 8232 30000 8328
rect 29920 8168 29928 8232
rect 29992 8168 30000 8232
rect 29920 8072 30000 8168
rect 29920 8008 29928 8072
rect 29992 8008 30000 8072
rect 29920 7912 30000 8008
rect 29920 7848 29928 7912
rect 29992 7848 30000 7912
rect 29920 7752 30000 7848
rect 29920 7688 29928 7752
rect 29992 7688 30000 7752
rect 29920 7592 30000 7688
rect 29920 7528 29928 7592
rect 29992 7528 30000 7592
rect 29920 7432 30000 7528
rect 29920 7368 29928 7432
rect 29992 7368 30000 7432
rect 29920 7272 30000 7368
rect 29920 7208 29928 7272
rect 29992 7208 30000 7272
rect 29920 7112 30000 7208
rect 29920 7048 29928 7112
rect 29992 7048 30000 7112
rect 29920 6952 30000 7048
rect 29920 6888 29928 6952
rect 29992 6888 30000 6952
rect 29920 6792 30000 6888
rect 29920 6728 29928 6792
rect 29992 6728 30000 6792
rect 29920 6632 30000 6728
rect 29920 6568 29928 6632
rect 29992 6568 30000 6632
rect 29920 6472 30000 6568
rect 29920 6408 29928 6472
rect 29992 6408 30000 6472
rect 29920 6312 30000 6408
rect 29920 6248 29928 6312
rect 29992 6248 30000 6312
rect 29920 6152 30000 6248
rect 29920 6088 29928 6152
rect 29992 6088 30000 6152
rect 29920 5992 30000 6088
rect 29920 5928 29928 5992
rect 29992 5928 30000 5992
rect 29920 5832 30000 5928
rect 29920 5768 29928 5832
rect 29992 5768 30000 5832
rect 29920 5672 30000 5768
rect 29920 5608 29928 5672
rect 29992 5608 30000 5672
rect 29920 5512 30000 5608
rect 29920 5448 29928 5512
rect 29992 5448 30000 5512
rect 29920 5352 30000 5448
rect 29920 5288 29928 5352
rect 29992 5288 30000 5352
rect 29920 5192 30000 5288
rect 29920 5128 29928 5192
rect 29992 5128 30000 5192
rect 29920 5032 30000 5128
rect 29920 4968 29928 5032
rect 29992 4968 30000 5032
rect 29920 4872 30000 4968
rect 29920 4808 29928 4872
rect 29992 4808 30000 4872
rect 29920 4712 30000 4808
rect 29920 4648 29928 4712
rect 29992 4648 30000 4712
rect 29920 4552 30000 4648
rect 29920 4488 29928 4552
rect 29992 4488 30000 4552
rect 29920 4392 30000 4488
rect 29920 4328 29928 4392
rect 29992 4328 30000 4392
rect 29920 4232 30000 4328
rect 29920 4168 29928 4232
rect 29992 4168 30000 4232
rect 29920 4072 30000 4168
rect 29920 4008 29928 4072
rect 29992 4008 30000 4072
rect 29920 3912 30000 4008
rect 29920 3848 29928 3912
rect 29992 3848 30000 3912
rect 29920 3592 30000 3848
rect 29920 3528 29928 3592
rect 29992 3528 30000 3592
rect 29920 3432 30000 3528
rect 29920 3368 29928 3432
rect 29992 3368 30000 3432
rect 29920 3272 30000 3368
rect 29920 3208 29928 3272
rect 29992 3208 30000 3272
rect 29920 3112 30000 3208
rect 29920 3048 29928 3112
rect 29992 3048 30000 3112
rect 29920 2952 30000 3048
rect 29920 2888 29928 2952
rect 29992 2888 30000 2952
rect 29920 2792 30000 2888
rect 29920 2728 29928 2792
rect 29992 2728 30000 2792
rect 29920 2632 30000 2728
rect 29920 2568 29928 2632
rect 29992 2568 30000 2632
rect 29920 2472 30000 2568
rect 29920 2408 29928 2472
rect 29992 2408 30000 2472
rect 29920 2312 30000 2408
rect 29920 2248 29928 2312
rect 29992 2248 30000 2312
rect 29920 2152 30000 2248
rect 29920 2088 29928 2152
rect 29992 2088 30000 2152
rect 29920 1992 30000 2088
rect 29920 1928 29928 1992
rect 29992 1928 30000 1992
rect 29920 1832 30000 1928
rect 29920 1768 29928 1832
rect 29992 1768 30000 1832
rect 29920 1672 30000 1768
rect 29920 1608 29928 1672
rect 29992 1608 30000 1672
rect 29920 1512 30000 1608
rect 29920 1448 29928 1512
rect 29992 1448 30000 1512
rect 29920 1352 30000 1448
rect 29920 1288 29928 1352
rect 29992 1288 30000 1352
rect 29920 1192 30000 1288
rect 29920 1128 29928 1192
rect 29992 1128 30000 1192
rect 29920 1032 30000 1128
rect 29920 968 29928 1032
rect 29992 968 30000 1032
rect 29600 808 29608 872
rect 29672 808 29680 872
rect 29600 792 29680 808
rect 29600 728 29608 792
rect 29672 728 29680 792
rect 29600 712 29680 728
rect 29600 648 29608 712
rect 29672 648 29680 712
rect 29600 632 29680 648
rect 29600 568 29608 632
rect 29672 568 29680 632
rect 29600 552 29680 568
rect 29600 488 29608 552
rect 29672 488 29680 552
rect 29600 480 29680 488
rect 29920 872 30000 968
rect 29920 808 29928 872
rect 29992 808 30000 872
rect 29920 792 30000 808
rect 29920 728 29928 792
rect 29992 728 30000 792
rect 29920 712 30000 728
rect 29920 648 29928 712
rect 29992 648 30000 712
rect 29920 632 30000 648
rect 29920 568 29928 632
rect 29992 568 30000 632
rect 29920 552 30000 568
rect 29920 488 29928 552
rect 29992 488 30000 552
rect 29920 480 30000 488
rect 28800 328 28808 392
rect 28872 328 28880 392
rect 28800 312 28880 328
rect 28800 248 28808 312
rect 28872 248 28880 312
rect 28800 232 28880 248
rect 28800 168 28808 232
rect 28872 168 28880 232
rect 28800 152 28880 168
rect 28800 88 28808 152
rect 28872 88 28880 152
rect 28800 72 28880 88
rect 28800 8 28808 72
rect 28872 8 28880 72
rect 28800 0 28880 8
<< via3 >>
rect 8 31908 72 31912
rect 8 31852 12 31908
rect 12 31852 68 31908
rect 68 31852 72 31908
rect 8 31848 72 31852
rect 8 31748 72 31752
rect 8 31692 12 31748
rect 12 31692 68 31748
rect 68 31692 72 31748
rect 8 31688 72 31692
rect 8 31588 72 31592
rect 8 31532 12 31588
rect 12 31532 68 31588
rect 68 31532 72 31588
rect 8 31528 72 31532
rect 8 31428 72 31432
rect 8 31372 12 31428
rect 12 31372 68 31428
rect 68 31372 72 31428
rect 8 31368 72 31372
rect 8 31268 72 31272
rect 8 31212 12 31268
rect 12 31212 68 31268
rect 68 31212 72 31268
rect 8 31208 72 31212
rect 8 31108 72 31112
rect 8 31052 12 31108
rect 12 31052 68 31108
rect 68 31052 72 31108
rect 8 31048 72 31052
rect 8 30948 72 30952
rect 8 30892 12 30948
rect 12 30892 68 30948
rect 68 30892 72 30948
rect 8 30888 72 30892
rect 8 30788 72 30792
rect 8 30732 12 30788
rect 12 30732 68 30788
rect 68 30732 72 30788
rect 8 30728 72 30732
rect 8 30628 72 30632
rect 8 30572 12 30628
rect 12 30572 68 30628
rect 68 30572 72 30628
rect 8 30568 72 30572
rect 8 30468 72 30472
rect 8 30412 12 30468
rect 12 30412 68 30468
rect 68 30412 72 30468
rect 8 30408 72 30412
rect 8 30308 72 30312
rect 8 30252 12 30308
rect 12 30252 68 30308
rect 68 30252 72 30308
rect 8 30248 72 30252
rect 8 30148 72 30152
rect 8 30092 12 30148
rect 12 30092 68 30148
rect 68 30092 72 30148
rect 8 30088 72 30092
rect 8 29988 72 29992
rect 8 29932 12 29988
rect 12 29932 68 29988
rect 68 29932 72 29988
rect 8 29928 72 29932
rect 8 29828 72 29832
rect 8 29772 12 29828
rect 12 29772 68 29828
rect 68 29772 72 29828
rect 8 29768 72 29772
rect 8 29668 72 29672
rect 8 29612 12 29668
rect 12 29612 68 29668
rect 68 29612 72 29668
rect 8 29608 72 29612
rect 8 29508 72 29512
rect 8 29452 12 29508
rect 12 29452 68 29508
rect 68 29452 72 29508
rect 8 29448 72 29452
rect 8 29348 72 29352
rect 8 29292 12 29348
rect 12 29292 68 29348
rect 68 29292 72 29348
rect 8 29288 72 29292
rect 8 29188 72 29192
rect 8 29132 12 29188
rect 12 29132 68 29188
rect 68 29132 72 29188
rect 8 29128 72 29132
rect 8 29028 72 29032
rect 8 28972 12 29028
rect 12 28972 68 29028
rect 68 28972 72 29028
rect 8 28968 72 28972
rect 8 28868 72 28872
rect 8 28812 12 28868
rect 12 28812 68 28868
rect 68 28812 72 28868
rect 8 28808 72 28812
rect 8 28708 72 28712
rect 8 28652 12 28708
rect 12 28652 68 28708
rect 68 28652 72 28708
rect 8 28648 72 28652
rect 8 28548 72 28552
rect 8 28492 12 28548
rect 12 28492 68 28548
rect 68 28492 72 28548
rect 8 28488 72 28492
rect 8 28388 72 28392
rect 8 28332 12 28388
rect 12 28332 68 28388
rect 68 28332 72 28388
rect 8 28328 72 28332
rect 8 28228 72 28232
rect 8 28172 12 28228
rect 12 28172 68 28228
rect 68 28172 72 28228
rect 8 28168 72 28172
rect 8 28068 72 28072
rect 8 28012 12 28068
rect 12 28012 68 28068
rect 68 28012 72 28068
rect 8 28008 72 28012
rect 8 27908 72 27912
rect 8 27852 12 27908
rect 12 27852 68 27908
rect 68 27852 72 27908
rect 8 27848 72 27852
rect 8 27748 72 27752
rect 8 27692 12 27748
rect 12 27692 68 27748
rect 68 27692 72 27748
rect 8 27688 72 27692
rect 8 27588 72 27592
rect 8 27532 12 27588
rect 12 27532 68 27588
rect 68 27532 72 27588
rect 8 27528 72 27532
rect 8 27428 72 27432
rect 8 27372 12 27428
rect 12 27372 68 27428
rect 68 27372 72 27428
rect 8 27368 72 27372
rect 8 27268 72 27272
rect 8 27212 12 27268
rect 12 27212 68 27268
rect 68 27212 72 27268
rect 8 27208 72 27212
rect 8 27108 72 27112
rect 8 27052 12 27108
rect 12 27052 68 27108
rect 68 27052 72 27108
rect 8 27048 72 27052
rect 8 26948 72 26952
rect 8 26892 12 26948
rect 12 26892 68 26948
rect 68 26892 72 26948
rect 8 26888 72 26892
rect 8 26788 72 26792
rect 8 26732 12 26788
rect 12 26732 68 26788
rect 68 26732 72 26788
rect 8 26728 72 26732
rect 8 26628 72 26632
rect 8 26572 12 26628
rect 12 26572 68 26628
rect 68 26572 72 26628
rect 8 26568 72 26572
rect 8 26468 72 26472
rect 8 26412 12 26468
rect 12 26412 68 26468
rect 68 26412 72 26468
rect 8 26408 72 26412
rect 8 26308 72 26312
rect 8 26252 12 26308
rect 12 26252 68 26308
rect 68 26252 72 26308
rect 8 26248 72 26252
rect 8 26148 72 26152
rect 8 26092 12 26148
rect 12 26092 68 26148
rect 68 26092 72 26148
rect 8 26088 72 26092
rect 8 25988 72 25992
rect 8 25932 12 25988
rect 12 25932 68 25988
rect 68 25932 72 25988
rect 8 25928 72 25932
rect 8 25828 72 25832
rect 8 25772 12 25828
rect 12 25772 68 25828
rect 68 25772 72 25828
rect 8 25768 72 25772
rect 8 25668 72 25672
rect 8 25612 12 25668
rect 12 25612 68 25668
rect 68 25612 72 25668
rect 8 25608 72 25612
rect 8 25508 72 25512
rect 8 25452 12 25508
rect 12 25452 68 25508
rect 68 25452 72 25508
rect 8 25448 72 25452
rect 8 25348 72 25352
rect 8 25292 12 25348
rect 12 25292 68 25348
rect 68 25292 72 25348
rect 8 25288 72 25292
rect 8 25188 72 25192
rect 8 25132 12 25188
rect 12 25132 68 25188
rect 68 25132 72 25188
rect 8 25128 72 25132
rect 8 25028 72 25032
rect 8 24972 12 25028
rect 12 24972 68 25028
rect 68 24972 72 25028
rect 8 24968 72 24972
rect 8 24868 72 24872
rect 8 24812 12 24868
rect 12 24812 68 24868
rect 68 24812 72 24868
rect 8 24808 72 24812
rect 8 24708 72 24712
rect 8 24652 12 24708
rect 12 24652 68 24708
rect 68 24652 72 24708
rect 8 24648 72 24652
rect 8 24548 72 24552
rect 8 24492 12 24548
rect 12 24492 68 24548
rect 68 24492 72 24548
rect 8 24488 72 24492
rect 8 24388 72 24392
rect 8 24332 12 24388
rect 12 24332 68 24388
rect 68 24332 72 24388
rect 8 24328 72 24332
rect 8 24228 72 24232
rect 8 24172 12 24228
rect 12 24172 68 24228
rect 68 24172 72 24228
rect 8 24168 72 24172
rect 8 24068 72 24072
rect 8 24012 12 24068
rect 12 24012 68 24068
rect 68 24012 72 24068
rect 8 24008 72 24012
rect 8 23908 72 23912
rect 8 23852 12 23908
rect 12 23852 68 23908
rect 68 23852 72 23908
rect 8 23848 72 23852
rect 8 23748 72 23752
rect 8 23692 12 23748
rect 12 23692 68 23748
rect 68 23692 72 23748
rect 8 23688 72 23692
rect 8 23588 72 23592
rect 8 23532 12 23588
rect 12 23532 68 23588
rect 68 23532 72 23588
rect 8 23528 72 23532
rect 8 23428 72 23432
rect 8 23372 12 23428
rect 12 23372 68 23428
rect 68 23372 72 23428
rect 8 23368 72 23372
rect 8 23268 72 23272
rect 8 23212 12 23268
rect 12 23212 68 23268
rect 68 23212 72 23268
rect 8 23208 72 23212
rect 8 23108 72 23112
rect 8 23052 12 23108
rect 12 23052 68 23108
rect 68 23052 72 23108
rect 8 23048 72 23052
rect 8 22948 72 22952
rect 8 22892 12 22948
rect 12 22892 68 22948
rect 68 22892 72 22948
rect 8 22888 72 22892
rect 8 22788 72 22792
rect 8 22732 12 22788
rect 12 22732 68 22788
rect 68 22732 72 22788
rect 8 22728 72 22732
rect 8 22468 72 22472
rect 8 22412 12 22468
rect 12 22412 68 22468
rect 68 22412 72 22468
rect 8 22408 72 22412
rect 8 22308 72 22312
rect 8 22252 12 22308
rect 12 22252 68 22308
rect 68 22252 72 22308
rect 8 22248 72 22252
rect 8 22148 72 22152
rect 8 22092 12 22148
rect 12 22092 68 22148
rect 68 22092 72 22148
rect 8 22088 72 22092
rect 8 21988 72 21992
rect 8 21932 12 21988
rect 12 21932 68 21988
rect 68 21932 72 21988
rect 8 21928 72 21932
rect 8 21828 72 21832
rect 8 21772 12 21828
rect 12 21772 68 21828
rect 68 21772 72 21828
rect 8 21768 72 21772
rect 8 21668 72 21672
rect 8 21612 12 21668
rect 12 21612 68 21668
rect 68 21612 72 21668
rect 8 21608 72 21612
rect 8 21508 72 21512
rect 8 21452 12 21508
rect 12 21452 68 21508
rect 68 21452 72 21508
rect 8 21448 72 21452
rect 8 21348 72 21352
rect 8 21292 12 21348
rect 12 21292 68 21348
rect 68 21292 72 21348
rect 8 21288 72 21292
rect 8 21188 72 21192
rect 8 21132 12 21188
rect 12 21132 68 21188
rect 68 21132 72 21188
rect 8 21128 72 21132
rect 8 21028 72 21032
rect 8 20972 12 21028
rect 12 20972 68 21028
rect 68 20972 72 21028
rect 8 20968 72 20972
rect 8 20868 72 20872
rect 8 20812 12 20868
rect 12 20812 68 20868
rect 68 20812 72 20868
rect 8 20808 72 20812
rect 8 20708 72 20712
rect 8 20652 12 20708
rect 12 20652 68 20708
rect 68 20652 72 20708
rect 8 20648 72 20652
rect 8 20548 72 20552
rect 8 20492 12 20548
rect 12 20492 68 20548
rect 68 20492 72 20548
rect 8 20488 72 20492
rect 8 20388 72 20392
rect 8 20332 12 20388
rect 12 20332 68 20388
rect 68 20332 72 20388
rect 8 20328 72 20332
rect 8 20228 72 20232
rect 8 20172 12 20228
rect 12 20172 68 20228
rect 68 20172 72 20228
rect 8 20168 72 20172
rect 8 20068 72 20072
rect 8 20012 12 20068
rect 12 20012 68 20068
rect 68 20012 72 20068
rect 8 20008 72 20012
rect 8 19908 72 19912
rect 8 19852 12 19908
rect 12 19852 68 19908
rect 68 19852 72 19908
rect 8 19848 72 19852
rect 8 19748 72 19752
rect 8 19692 12 19748
rect 12 19692 68 19748
rect 68 19692 72 19748
rect 8 19688 72 19692
rect 8 19588 72 19592
rect 8 19532 12 19588
rect 12 19532 68 19588
rect 68 19532 72 19588
rect 8 19528 72 19532
rect 8 19428 72 19432
rect 8 19372 12 19428
rect 12 19372 68 19428
rect 68 19372 72 19428
rect 8 19368 72 19372
rect 8 19268 72 19272
rect 8 19212 12 19268
rect 12 19212 68 19268
rect 68 19212 72 19268
rect 8 19208 72 19212
rect 8 19108 72 19112
rect 8 19052 12 19108
rect 12 19052 68 19108
rect 68 19052 72 19108
rect 8 19048 72 19052
rect 8 18948 72 18952
rect 8 18892 12 18948
rect 12 18892 68 18948
rect 68 18892 72 18948
rect 8 18888 72 18892
rect 8 18788 72 18792
rect 8 18732 12 18788
rect 12 18732 68 18788
rect 68 18732 72 18788
rect 8 18728 72 18732
rect 8 18628 72 18632
rect 8 18572 12 18628
rect 12 18572 68 18628
rect 68 18572 72 18628
rect 8 18568 72 18572
rect 8 18468 72 18472
rect 8 18412 12 18468
rect 12 18412 68 18468
rect 68 18412 72 18468
rect 8 18408 72 18412
rect 8 18308 72 18312
rect 8 18252 12 18308
rect 12 18252 68 18308
rect 68 18252 72 18308
rect 8 18248 72 18252
rect 8 18148 72 18152
rect 8 18092 12 18148
rect 12 18092 68 18148
rect 68 18092 72 18148
rect 8 18088 72 18092
rect 8 17988 72 17992
rect 8 17932 12 17988
rect 12 17932 68 17988
rect 68 17932 72 17988
rect 8 17928 72 17932
rect 8 17828 72 17832
rect 8 17772 12 17828
rect 12 17772 68 17828
rect 68 17772 72 17828
rect 8 17768 72 17772
rect 8 17668 72 17672
rect 8 17612 12 17668
rect 12 17612 68 17668
rect 68 17612 72 17668
rect 8 17608 72 17612
rect 8 17508 72 17512
rect 8 17452 12 17508
rect 12 17452 68 17508
rect 68 17452 72 17508
rect 8 17448 72 17452
rect 8 17348 72 17352
rect 8 17292 12 17348
rect 12 17292 68 17348
rect 68 17292 72 17348
rect 8 17288 72 17292
rect 8 17188 72 17192
rect 8 17132 12 17188
rect 12 17132 68 17188
rect 68 17132 72 17188
rect 8 17128 72 17132
rect 8 17028 72 17032
rect 8 16972 12 17028
rect 12 16972 68 17028
rect 68 16972 72 17028
rect 8 16968 72 16972
rect 8 16708 72 16712
rect 8 16652 12 16708
rect 12 16652 68 16708
rect 68 16652 72 16708
rect 8 16648 72 16652
rect 8 16548 72 16552
rect 8 16492 12 16548
rect 12 16492 68 16548
rect 68 16492 72 16548
rect 8 16488 72 16492
rect 8 16388 72 16392
rect 8 16332 12 16388
rect 12 16332 68 16388
rect 68 16332 72 16388
rect 8 16328 72 16332
rect 8 16228 72 16232
rect 8 16172 12 16228
rect 12 16172 68 16228
rect 68 16172 72 16228
rect 8 16168 72 16172
rect 8 15908 72 15912
rect 8 15852 12 15908
rect 12 15852 68 15908
rect 68 15852 72 15908
rect 8 15848 72 15852
rect 8 15748 72 15752
rect 8 15692 12 15748
rect 12 15692 68 15748
rect 68 15692 72 15748
rect 8 15688 72 15692
rect 8 15588 72 15592
rect 8 15532 12 15588
rect 12 15532 68 15588
rect 68 15532 72 15588
rect 8 15528 72 15532
rect 8 15428 72 15432
rect 8 15372 12 15428
rect 12 15372 68 15428
rect 68 15372 72 15428
rect 8 15368 72 15372
rect 8 15268 72 15272
rect 8 15212 12 15268
rect 12 15212 68 15268
rect 68 15212 72 15268
rect 8 15208 72 15212
rect 8 15108 72 15112
rect 8 15052 12 15108
rect 12 15052 68 15108
rect 68 15052 72 15108
rect 8 15048 72 15052
rect 8 14948 72 14952
rect 8 14892 12 14948
rect 12 14892 68 14948
rect 68 14892 72 14948
rect 8 14888 72 14892
rect 8 14788 72 14792
rect 8 14732 12 14788
rect 12 14732 68 14788
rect 68 14732 72 14788
rect 8 14728 72 14732
rect 8 14628 72 14632
rect 8 14572 12 14628
rect 12 14572 68 14628
rect 68 14572 72 14628
rect 8 14568 72 14572
rect 8 14468 72 14472
rect 8 14412 12 14468
rect 12 14412 68 14468
rect 68 14412 72 14468
rect 8 14408 72 14412
rect 8 14308 72 14312
rect 8 14252 12 14308
rect 12 14252 68 14308
rect 68 14252 72 14308
rect 8 14248 72 14252
rect 8 14148 72 14152
rect 8 14092 12 14148
rect 12 14092 68 14148
rect 68 14092 72 14148
rect 8 14088 72 14092
rect 8 13988 72 13992
rect 8 13932 12 13988
rect 12 13932 68 13988
rect 68 13932 72 13988
rect 8 13928 72 13932
rect 8 13828 72 13832
rect 8 13772 12 13828
rect 12 13772 68 13828
rect 68 13772 72 13828
rect 8 13768 72 13772
rect 8 13668 72 13672
rect 8 13612 12 13668
rect 12 13612 68 13668
rect 68 13612 72 13668
rect 8 13608 72 13612
rect 8 13508 72 13512
rect 8 13452 12 13508
rect 12 13452 68 13508
rect 68 13452 72 13508
rect 8 13448 72 13452
rect 8 13348 72 13352
rect 8 13292 12 13348
rect 12 13292 68 13348
rect 68 13292 72 13348
rect 8 13288 72 13292
rect 8 13188 72 13192
rect 8 13132 12 13188
rect 12 13132 68 13188
rect 68 13132 72 13188
rect 8 13128 72 13132
rect 8 13028 72 13032
rect 8 12972 12 13028
rect 12 12972 68 13028
rect 68 12972 72 13028
rect 8 12968 72 12972
rect 8 12868 72 12872
rect 8 12812 12 12868
rect 12 12812 68 12868
rect 68 12812 72 12868
rect 8 12808 72 12812
rect 8 12708 72 12712
rect 8 12652 12 12708
rect 12 12652 68 12708
rect 68 12652 72 12708
rect 8 12648 72 12652
rect 8 12548 72 12552
rect 8 12492 12 12548
rect 12 12492 68 12548
rect 68 12492 72 12548
rect 8 12488 72 12492
rect 8 12388 72 12392
rect 8 12332 12 12388
rect 12 12332 68 12388
rect 68 12332 72 12388
rect 8 12328 72 12332
rect 8 12228 72 12232
rect 8 12172 12 12228
rect 12 12172 68 12228
rect 68 12172 72 12228
rect 8 12168 72 12172
rect 8 12068 72 12072
rect 8 12012 12 12068
rect 12 12012 68 12068
rect 68 12012 72 12068
rect 8 12008 72 12012
rect 8 11908 72 11912
rect 8 11852 12 11908
rect 12 11852 68 11908
rect 68 11852 72 11908
rect 8 11848 72 11852
rect 8 11748 72 11752
rect 8 11692 12 11748
rect 12 11692 68 11748
rect 68 11692 72 11748
rect 8 11688 72 11692
rect 8 11588 72 11592
rect 8 11532 12 11588
rect 12 11532 68 11588
rect 68 11532 72 11588
rect 8 11528 72 11532
rect 8 11428 72 11432
rect 8 11372 12 11428
rect 12 11372 68 11428
rect 68 11372 72 11428
rect 8 11368 72 11372
rect 8 11268 72 11272
rect 8 11212 12 11268
rect 12 11212 68 11268
rect 68 11212 72 11268
rect 8 11208 72 11212
rect 8 11108 72 11112
rect 8 11052 12 11108
rect 12 11052 68 11108
rect 68 11052 72 11108
rect 8 11048 72 11052
rect 8 10948 72 10952
rect 8 10892 12 10948
rect 12 10892 68 10948
rect 68 10892 72 10948
rect 8 10888 72 10892
rect 8 10788 72 10792
rect 8 10732 12 10788
rect 12 10732 68 10788
rect 68 10732 72 10788
rect 8 10728 72 10732
rect 8 10628 72 10632
rect 8 10572 12 10628
rect 12 10572 68 10628
rect 68 10572 72 10628
rect 8 10568 72 10572
rect 8 10468 72 10472
rect 8 10412 12 10468
rect 12 10412 68 10468
rect 68 10412 72 10468
rect 8 10408 72 10412
rect 8 10148 72 10152
rect 8 10092 12 10148
rect 12 10092 68 10148
rect 68 10092 72 10148
rect 8 10088 72 10092
rect 8 9988 72 9992
rect 8 9932 12 9988
rect 12 9932 68 9988
rect 68 9932 72 9988
rect 8 9928 72 9932
rect 8 9828 72 9832
rect 8 9772 12 9828
rect 12 9772 68 9828
rect 68 9772 72 9828
rect 8 9768 72 9772
rect 8 9668 72 9672
rect 8 9612 12 9668
rect 12 9612 68 9668
rect 68 9612 72 9668
rect 8 9608 72 9612
rect 8 9508 72 9512
rect 8 9452 12 9508
rect 12 9452 68 9508
rect 68 9452 72 9508
rect 8 9448 72 9452
rect 8 9348 72 9352
rect 8 9292 12 9348
rect 12 9292 68 9348
rect 68 9292 72 9348
rect 8 9288 72 9292
rect 8 9188 72 9192
rect 8 9132 12 9188
rect 12 9132 68 9188
rect 68 9132 72 9188
rect 8 9128 72 9132
rect 8 9028 72 9032
rect 8 8972 12 9028
rect 12 8972 68 9028
rect 68 8972 72 9028
rect 8 8968 72 8972
rect 8 8868 72 8872
rect 8 8812 12 8868
rect 12 8812 68 8868
rect 68 8812 72 8868
rect 8 8808 72 8812
rect 8 8708 72 8712
rect 8 8652 12 8708
rect 12 8652 68 8708
rect 68 8652 72 8708
rect 8 8648 72 8652
rect 8 8548 72 8552
rect 8 8492 12 8548
rect 12 8492 68 8548
rect 68 8492 72 8548
rect 8 8488 72 8492
rect 8 8388 72 8392
rect 8 8332 12 8388
rect 12 8332 68 8388
rect 68 8332 72 8388
rect 8 8328 72 8332
rect 8 8228 72 8232
rect 8 8172 12 8228
rect 12 8172 68 8228
rect 68 8172 72 8228
rect 8 8168 72 8172
rect 8 8068 72 8072
rect 8 8012 12 8068
rect 12 8012 68 8068
rect 68 8012 72 8068
rect 8 8008 72 8012
rect 8 7908 72 7912
rect 8 7852 12 7908
rect 12 7852 68 7908
rect 68 7852 72 7908
rect 8 7848 72 7852
rect 8 7748 72 7752
rect 8 7692 12 7748
rect 12 7692 68 7748
rect 68 7692 72 7748
rect 8 7688 72 7692
rect 8 7588 72 7592
rect 8 7532 12 7588
rect 12 7532 68 7588
rect 68 7532 72 7588
rect 8 7528 72 7532
rect 8 7428 72 7432
rect 8 7372 12 7428
rect 12 7372 68 7428
rect 68 7372 72 7428
rect 8 7368 72 7372
rect 8 7268 72 7272
rect 8 7212 12 7268
rect 12 7212 68 7268
rect 68 7212 72 7268
rect 8 7208 72 7212
rect 8 7108 72 7112
rect 8 7052 12 7108
rect 12 7052 68 7108
rect 68 7052 72 7108
rect 8 7048 72 7052
rect 8 6948 72 6952
rect 8 6892 12 6948
rect 12 6892 68 6948
rect 68 6892 72 6948
rect 8 6888 72 6892
rect 8 6788 72 6792
rect 8 6732 12 6788
rect 12 6732 68 6788
rect 68 6732 72 6788
rect 8 6728 72 6732
rect 8 6628 72 6632
rect 8 6572 12 6628
rect 12 6572 68 6628
rect 68 6572 72 6628
rect 8 6568 72 6572
rect 8 6468 72 6472
rect 8 6412 12 6468
rect 12 6412 68 6468
rect 68 6412 72 6468
rect 8 6408 72 6412
rect 8 6308 72 6312
rect 8 6252 12 6308
rect 12 6252 68 6308
rect 68 6252 72 6308
rect 8 6248 72 6252
rect 8 6148 72 6152
rect 8 6092 12 6148
rect 12 6092 68 6148
rect 68 6092 72 6148
rect 8 6088 72 6092
rect 8 5988 72 5992
rect 8 5932 12 5988
rect 12 5932 68 5988
rect 68 5932 72 5988
rect 8 5928 72 5932
rect 8 5828 72 5832
rect 8 5772 12 5828
rect 12 5772 68 5828
rect 68 5772 72 5828
rect 8 5768 72 5772
rect 8 5668 72 5672
rect 8 5612 12 5668
rect 12 5612 68 5668
rect 68 5612 72 5668
rect 8 5608 72 5612
rect 8 5508 72 5512
rect 8 5452 12 5508
rect 12 5452 68 5508
rect 68 5452 72 5508
rect 8 5448 72 5452
rect 8 5348 72 5352
rect 8 5292 12 5348
rect 12 5292 68 5348
rect 68 5292 72 5348
rect 8 5288 72 5292
rect 8 5188 72 5192
rect 8 5132 12 5188
rect 12 5132 68 5188
rect 68 5132 72 5188
rect 8 5128 72 5132
rect 8 5028 72 5032
rect 8 4972 12 5028
rect 12 4972 68 5028
rect 68 4972 72 5028
rect 8 4968 72 4972
rect 8 4868 72 4872
rect 8 4812 12 4868
rect 12 4812 68 4868
rect 68 4812 72 4868
rect 8 4808 72 4812
rect 8 4708 72 4712
rect 8 4652 12 4708
rect 12 4652 68 4708
rect 68 4652 72 4708
rect 8 4648 72 4652
rect 8 4548 72 4552
rect 8 4492 12 4548
rect 12 4492 68 4548
rect 68 4492 72 4548
rect 8 4488 72 4492
rect 8 4388 72 4392
rect 8 4332 12 4388
rect 12 4332 68 4388
rect 68 4332 72 4388
rect 8 4328 72 4332
rect 8 4228 72 4232
rect 8 4172 12 4228
rect 12 4172 68 4228
rect 68 4172 72 4228
rect 8 4168 72 4172
rect 8 4068 72 4072
rect 8 4012 12 4068
rect 12 4012 68 4068
rect 68 4012 72 4068
rect 8 4008 72 4012
rect 8 3908 72 3912
rect 8 3852 12 3908
rect 12 3852 68 3908
rect 68 3852 72 3908
rect 8 3848 72 3852
rect 8 3748 72 3752
rect 8 3692 12 3748
rect 12 3692 68 3748
rect 68 3692 72 3748
rect 8 3688 72 3692
rect 8 3588 72 3592
rect 8 3532 12 3588
rect 12 3532 68 3588
rect 68 3532 72 3588
rect 8 3528 72 3532
rect 8 3428 72 3432
rect 8 3372 12 3428
rect 12 3372 68 3428
rect 68 3372 72 3428
rect 8 3368 72 3372
rect 8 3268 72 3272
rect 8 3212 12 3268
rect 12 3212 68 3268
rect 68 3212 72 3268
rect 8 3208 72 3212
rect 8 3108 72 3112
rect 8 3052 12 3108
rect 12 3052 68 3108
rect 68 3052 72 3108
rect 8 3048 72 3052
rect 8 2948 72 2952
rect 8 2892 12 2948
rect 12 2892 68 2948
rect 68 2892 72 2948
rect 8 2888 72 2892
rect 8 2788 72 2792
rect 8 2732 12 2788
rect 12 2732 68 2788
rect 68 2732 72 2788
rect 8 2728 72 2732
rect 8 2628 72 2632
rect 8 2572 12 2628
rect 12 2572 68 2628
rect 68 2572 72 2628
rect 8 2568 72 2572
rect 8 2468 72 2472
rect 8 2412 12 2468
rect 12 2412 68 2468
rect 68 2412 72 2468
rect 8 2408 72 2412
rect 8 2308 72 2312
rect 8 2252 12 2308
rect 12 2252 68 2308
rect 68 2252 72 2308
rect 8 2248 72 2252
rect 8 2148 72 2152
rect 8 2092 12 2148
rect 12 2092 68 2148
rect 68 2092 72 2148
rect 8 2088 72 2092
rect 8 1988 72 1992
rect 8 1932 12 1988
rect 12 1932 68 1988
rect 68 1932 72 1988
rect 8 1928 72 1932
rect 8 1828 72 1832
rect 8 1772 12 1828
rect 12 1772 68 1828
rect 68 1772 72 1828
rect 8 1768 72 1772
rect 8 1668 72 1672
rect 8 1612 12 1668
rect 12 1612 68 1668
rect 68 1612 72 1668
rect 8 1608 72 1612
rect 8 1508 72 1512
rect 8 1452 12 1508
rect 12 1452 68 1508
rect 68 1452 72 1508
rect 8 1448 72 1452
rect 8 1348 72 1352
rect 8 1292 12 1348
rect 12 1292 68 1348
rect 68 1292 72 1348
rect 8 1288 72 1292
rect 8 1188 72 1192
rect 8 1132 12 1188
rect 12 1132 68 1188
rect 68 1132 72 1188
rect 8 1128 72 1132
rect 8 1028 72 1032
rect 8 972 12 1028
rect 12 972 68 1028
rect 68 972 72 1028
rect 8 968 72 972
rect 168 22568 232 22632
rect 168 16808 232 16872
rect 168 16008 232 16072
rect 168 10248 232 10312
rect 328 31908 392 31912
rect 328 31852 332 31908
rect 332 31852 388 31908
rect 388 31852 392 31908
rect 328 31848 392 31852
rect 328 31748 392 31752
rect 328 31692 332 31748
rect 332 31692 388 31748
rect 388 31692 392 31748
rect 328 31688 392 31692
rect 328 31588 392 31592
rect 328 31532 332 31588
rect 332 31532 388 31588
rect 388 31532 392 31588
rect 328 31528 392 31532
rect 328 31428 392 31432
rect 328 31372 332 31428
rect 332 31372 388 31428
rect 388 31372 392 31428
rect 328 31368 392 31372
rect 328 31268 392 31272
rect 328 31212 332 31268
rect 332 31212 388 31268
rect 388 31212 392 31268
rect 328 31208 392 31212
rect 328 31108 392 31112
rect 328 31052 332 31108
rect 332 31052 388 31108
rect 388 31052 392 31108
rect 328 31048 392 31052
rect 328 30948 392 30952
rect 328 30892 332 30948
rect 332 30892 388 30948
rect 388 30892 392 30948
rect 328 30888 392 30892
rect 328 30788 392 30792
rect 328 30732 332 30788
rect 332 30732 388 30788
rect 388 30732 392 30788
rect 328 30728 392 30732
rect 328 30628 392 30632
rect 328 30572 332 30628
rect 332 30572 388 30628
rect 388 30572 392 30628
rect 328 30568 392 30572
rect 328 30468 392 30472
rect 328 30412 332 30468
rect 332 30412 388 30468
rect 388 30412 392 30468
rect 328 30408 392 30412
rect 328 30308 392 30312
rect 328 30252 332 30308
rect 332 30252 388 30308
rect 388 30252 392 30308
rect 328 30248 392 30252
rect 328 30148 392 30152
rect 328 30092 332 30148
rect 332 30092 388 30148
rect 388 30092 392 30148
rect 328 30088 392 30092
rect 328 29988 392 29992
rect 328 29932 332 29988
rect 332 29932 388 29988
rect 388 29932 392 29988
rect 328 29928 392 29932
rect 328 29828 392 29832
rect 328 29772 332 29828
rect 332 29772 388 29828
rect 388 29772 392 29828
rect 328 29768 392 29772
rect 328 29668 392 29672
rect 328 29612 332 29668
rect 332 29612 388 29668
rect 388 29612 392 29668
rect 328 29608 392 29612
rect 328 29508 392 29512
rect 328 29452 332 29508
rect 332 29452 388 29508
rect 388 29452 392 29508
rect 328 29448 392 29452
rect 328 29348 392 29352
rect 328 29292 332 29348
rect 332 29292 388 29348
rect 388 29292 392 29348
rect 328 29288 392 29292
rect 328 29188 392 29192
rect 328 29132 332 29188
rect 332 29132 388 29188
rect 388 29132 392 29188
rect 328 29128 392 29132
rect 328 29028 392 29032
rect 328 28972 332 29028
rect 332 28972 388 29028
rect 388 28972 392 29028
rect 328 28968 392 28972
rect 328 28868 392 28872
rect 328 28812 332 28868
rect 332 28812 388 28868
rect 388 28812 392 28868
rect 328 28808 392 28812
rect 328 28708 392 28712
rect 328 28652 332 28708
rect 332 28652 388 28708
rect 388 28652 392 28708
rect 328 28648 392 28652
rect 328 28548 392 28552
rect 328 28492 332 28548
rect 332 28492 388 28548
rect 388 28492 392 28548
rect 328 28488 392 28492
rect 328 28388 392 28392
rect 328 28332 332 28388
rect 332 28332 388 28388
rect 388 28332 392 28388
rect 328 28328 392 28332
rect 328 28228 392 28232
rect 328 28172 332 28228
rect 332 28172 388 28228
rect 388 28172 392 28228
rect 328 28168 392 28172
rect 328 28068 392 28072
rect 328 28012 332 28068
rect 332 28012 388 28068
rect 388 28012 392 28068
rect 328 28008 392 28012
rect 328 27908 392 27912
rect 328 27852 332 27908
rect 332 27852 388 27908
rect 388 27852 392 27908
rect 328 27848 392 27852
rect 328 27748 392 27752
rect 328 27692 332 27748
rect 332 27692 388 27748
rect 388 27692 392 27748
rect 328 27688 392 27692
rect 328 27588 392 27592
rect 328 27532 332 27588
rect 332 27532 388 27588
rect 388 27532 392 27588
rect 328 27528 392 27532
rect 328 27428 392 27432
rect 328 27372 332 27428
rect 332 27372 388 27428
rect 388 27372 392 27428
rect 328 27368 392 27372
rect 328 27268 392 27272
rect 328 27212 332 27268
rect 332 27212 388 27268
rect 388 27212 392 27268
rect 328 27208 392 27212
rect 328 27108 392 27112
rect 328 27052 332 27108
rect 332 27052 388 27108
rect 388 27052 392 27108
rect 328 27048 392 27052
rect 328 26948 392 26952
rect 328 26892 332 26948
rect 332 26892 388 26948
rect 388 26892 392 26948
rect 328 26888 392 26892
rect 328 26788 392 26792
rect 328 26732 332 26788
rect 332 26732 388 26788
rect 388 26732 392 26788
rect 328 26728 392 26732
rect 328 26628 392 26632
rect 328 26572 332 26628
rect 332 26572 388 26628
rect 388 26572 392 26628
rect 328 26568 392 26572
rect 328 26468 392 26472
rect 328 26412 332 26468
rect 332 26412 388 26468
rect 388 26412 392 26468
rect 328 26408 392 26412
rect 328 26308 392 26312
rect 328 26252 332 26308
rect 332 26252 388 26308
rect 388 26252 392 26308
rect 328 26248 392 26252
rect 328 26148 392 26152
rect 328 26092 332 26148
rect 332 26092 388 26148
rect 388 26092 392 26148
rect 328 26088 392 26092
rect 328 25988 392 25992
rect 328 25932 332 25988
rect 332 25932 388 25988
rect 388 25932 392 25988
rect 328 25928 392 25932
rect 328 25828 392 25832
rect 328 25772 332 25828
rect 332 25772 388 25828
rect 388 25772 392 25828
rect 328 25768 392 25772
rect 328 25668 392 25672
rect 328 25612 332 25668
rect 332 25612 388 25668
rect 388 25612 392 25668
rect 328 25608 392 25612
rect 328 25508 392 25512
rect 328 25452 332 25508
rect 332 25452 388 25508
rect 388 25452 392 25508
rect 328 25448 392 25452
rect 328 25348 392 25352
rect 328 25292 332 25348
rect 332 25292 388 25348
rect 388 25292 392 25348
rect 328 25288 392 25292
rect 328 25188 392 25192
rect 328 25132 332 25188
rect 332 25132 388 25188
rect 388 25132 392 25188
rect 328 25128 392 25132
rect 328 25028 392 25032
rect 328 24972 332 25028
rect 332 24972 388 25028
rect 388 24972 392 25028
rect 328 24968 392 24972
rect 328 24868 392 24872
rect 328 24812 332 24868
rect 332 24812 388 24868
rect 388 24812 392 24868
rect 328 24808 392 24812
rect 328 24708 392 24712
rect 328 24652 332 24708
rect 332 24652 388 24708
rect 388 24652 392 24708
rect 328 24648 392 24652
rect 328 24548 392 24552
rect 328 24492 332 24548
rect 332 24492 388 24548
rect 388 24492 392 24548
rect 328 24488 392 24492
rect 328 24388 392 24392
rect 328 24332 332 24388
rect 332 24332 388 24388
rect 388 24332 392 24388
rect 328 24328 392 24332
rect 328 24228 392 24232
rect 328 24172 332 24228
rect 332 24172 388 24228
rect 388 24172 392 24228
rect 328 24168 392 24172
rect 328 24068 392 24072
rect 328 24012 332 24068
rect 332 24012 388 24068
rect 388 24012 392 24068
rect 328 24008 392 24012
rect 328 23908 392 23912
rect 328 23852 332 23908
rect 332 23852 388 23908
rect 388 23852 392 23908
rect 328 23848 392 23852
rect 328 23748 392 23752
rect 328 23692 332 23748
rect 332 23692 388 23748
rect 388 23692 392 23748
rect 328 23688 392 23692
rect 328 23588 392 23592
rect 328 23532 332 23588
rect 332 23532 388 23588
rect 388 23532 392 23588
rect 328 23528 392 23532
rect 328 23428 392 23432
rect 328 23372 332 23428
rect 332 23372 388 23428
rect 388 23372 392 23428
rect 328 23368 392 23372
rect 328 23268 392 23272
rect 328 23212 332 23268
rect 332 23212 388 23268
rect 388 23212 392 23268
rect 328 23208 392 23212
rect 328 23108 392 23112
rect 328 23052 332 23108
rect 332 23052 388 23108
rect 388 23052 392 23108
rect 328 23048 392 23052
rect 328 22948 392 22952
rect 328 22892 332 22948
rect 332 22892 388 22948
rect 388 22892 392 22948
rect 328 22888 392 22892
rect 328 22788 392 22792
rect 328 22732 332 22788
rect 332 22732 388 22788
rect 388 22732 392 22788
rect 328 22728 392 22732
rect 328 22468 392 22472
rect 328 22412 332 22468
rect 332 22412 388 22468
rect 388 22412 392 22468
rect 328 22408 392 22412
rect 328 22308 392 22312
rect 328 22252 332 22308
rect 332 22252 388 22308
rect 388 22252 392 22308
rect 328 22248 392 22252
rect 328 22148 392 22152
rect 328 22092 332 22148
rect 332 22092 388 22148
rect 388 22092 392 22148
rect 328 22088 392 22092
rect 328 21988 392 21992
rect 328 21932 332 21988
rect 332 21932 388 21988
rect 388 21932 392 21988
rect 328 21928 392 21932
rect 328 21828 392 21832
rect 328 21772 332 21828
rect 332 21772 388 21828
rect 388 21772 392 21828
rect 328 21768 392 21772
rect 328 21668 392 21672
rect 328 21612 332 21668
rect 332 21612 388 21668
rect 388 21612 392 21668
rect 328 21608 392 21612
rect 328 21508 392 21512
rect 328 21452 332 21508
rect 332 21452 388 21508
rect 388 21452 392 21508
rect 328 21448 392 21452
rect 328 21348 392 21352
rect 328 21292 332 21348
rect 332 21292 388 21348
rect 388 21292 392 21348
rect 328 21288 392 21292
rect 328 21188 392 21192
rect 328 21132 332 21188
rect 332 21132 388 21188
rect 388 21132 392 21188
rect 328 21128 392 21132
rect 328 21028 392 21032
rect 328 20972 332 21028
rect 332 20972 388 21028
rect 388 20972 392 21028
rect 328 20968 392 20972
rect 328 20868 392 20872
rect 328 20812 332 20868
rect 332 20812 388 20868
rect 388 20812 392 20868
rect 328 20808 392 20812
rect 328 20708 392 20712
rect 328 20652 332 20708
rect 332 20652 388 20708
rect 388 20652 392 20708
rect 328 20648 392 20652
rect 328 20548 392 20552
rect 328 20492 332 20548
rect 332 20492 388 20548
rect 388 20492 392 20548
rect 328 20488 392 20492
rect 328 20388 392 20392
rect 328 20332 332 20388
rect 332 20332 388 20388
rect 388 20332 392 20388
rect 328 20328 392 20332
rect 328 20228 392 20232
rect 328 20172 332 20228
rect 332 20172 388 20228
rect 388 20172 392 20228
rect 328 20168 392 20172
rect 328 20068 392 20072
rect 328 20012 332 20068
rect 332 20012 388 20068
rect 388 20012 392 20068
rect 328 20008 392 20012
rect 328 19908 392 19912
rect 328 19852 332 19908
rect 332 19852 388 19908
rect 388 19852 392 19908
rect 328 19848 392 19852
rect 328 19748 392 19752
rect 328 19692 332 19748
rect 332 19692 388 19748
rect 388 19692 392 19748
rect 328 19688 392 19692
rect 328 19588 392 19592
rect 328 19532 332 19588
rect 332 19532 388 19588
rect 388 19532 392 19588
rect 328 19528 392 19532
rect 328 19428 392 19432
rect 328 19372 332 19428
rect 332 19372 388 19428
rect 388 19372 392 19428
rect 328 19368 392 19372
rect 328 19268 392 19272
rect 328 19212 332 19268
rect 332 19212 388 19268
rect 388 19212 392 19268
rect 328 19208 392 19212
rect 328 19108 392 19112
rect 328 19052 332 19108
rect 332 19052 388 19108
rect 388 19052 392 19108
rect 328 19048 392 19052
rect 328 18948 392 18952
rect 328 18892 332 18948
rect 332 18892 388 18948
rect 388 18892 392 18948
rect 328 18888 392 18892
rect 328 18788 392 18792
rect 328 18732 332 18788
rect 332 18732 388 18788
rect 388 18732 392 18788
rect 328 18728 392 18732
rect 328 18628 392 18632
rect 328 18572 332 18628
rect 332 18572 388 18628
rect 388 18572 392 18628
rect 328 18568 392 18572
rect 328 18468 392 18472
rect 328 18412 332 18468
rect 332 18412 388 18468
rect 388 18412 392 18468
rect 328 18408 392 18412
rect 328 18308 392 18312
rect 328 18252 332 18308
rect 332 18252 388 18308
rect 388 18252 392 18308
rect 328 18248 392 18252
rect 328 18148 392 18152
rect 328 18092 332 18148
rect 332 18092 388 18148
rect 388 18092 392 18148
rect 328 18088 392 18092
rect 328 17988 392 17992
rect 328 17932 332 17988
rect 332 17932 388 17988
rect 388 17932 392 17988
rect 328 17928 392 17932
rect 328 17828 392 17832
rect 328 17772 332 17828
rect 332 17772 388 17828
rect 388 17772 392 17828
rect 328 17768 392 17772
rect 328 17668 392 17672
rect 328 17612 332 17668
rect 332 17612 388 17668
rect 388 17612 392 17668
rect 328 17608 392 17612
rect 328 17508 392 17512
rect 328 17452 332 17508
rect 332 17452 388 17508
rect 388 17452 392 17508
rect 328 17448 392 17452
rect 328 17348 392 17352
rect 328 17292 332 17348
rect 332 17292 388 17348
rect 388 17292 392 17348
rect 328 17288 392 17292
rect 328 17188 392 17192
rect 328 17132 332 17188
rect 332 17132 388 17188
rect 388 17132 392 17188
rect 328 17128 392 17132
rect 328 17028 392 17032
rect 328 16972 332 17028
rect 332 16972 388 17028
rect 388 16972 392 17028
rect 328 16968 392 16972
rect 328 16708 392 16712
rect 328 16652 332 16708
rect 332 16652 388 16708
rect 388 16652 392 16708
rect 328 16648 392 16652
rect 328 16548 392 16552
rect 328 16492 332 16548
rect 332 16492 388 16548
rect 388 16492 392 16548
rect 328 16488 392 16492
rect 328 16388 392 16392
rect 328 16332 332 16388
rect 332 16332 388 16388
rect 388 16332 392 16388
rect 328 16328 392 16332
rect 328 16228 392 16232
rect 328 16172 332 16228
rect 332 16172 388 16228
rect 388 16172 392 16228
rect 328 16168 392 16172
rect 328 15908 392 15912
rect 328 15852 332 15908
rect 332 15852 388 15908
rect 388 15852 392 15908
rect 328 15848 392 15852
rect 328 15748 392 15752
rect 328 15692 332 15748
rect 332 15692 388 15748
rect 388 15692 392 15748
rect 328 15688 392 15692
rect 328 15588 392 15592
rect 328 15532 332 15588
rect 332 15532 388 15588
rect 388 15532 392 15588
rect 328 15528 392 15532
rect 328 15428 392 15432
rect 328 15372 332 15428
rect 332 15372 388 15428
rect 388 15372 392 15428
rect 328 15368 392 15372
rect 328 15268 392 15272
rect 328 15212 332 15268
rect 332 15212 388 15268
rect 388 15212 392 15268
rect 328 15208 392 15212
rect 328 15108 392 15112
rect 328 15052 332 15108
rect 332 15052 388 15108
rect 388 15052 392 15108
rect 328 15048 392 15052
rect 328 14948 392 14952
rect 328 14892 332 14948
rect 332 14892 388 14948
rect 388 14892 392 14948
rect 328 14888 392 14892
rect 328 14788 392 14792
rect 328 14732 332 14788
rect 332 14732 388 14788
rect 388 14732 392 14788
rect 328 14728 392 14732
rect 328 14628 392 14632
rect 328 14572 332 14628
rect 332 14572 388 14628
rect 388 14572 392 14628
rect 328 14568 392 14572
rect 328 14468 392 14472
rect 328 14412 332 14468
rect 332 14412 388 14468
rect 388 14412 392 14468
rect 328 14408 392 14412
rect 328 14308 392 14312
rect 328 14252 332 14308
rect 332 14252 388 14308
rect 388 14252 392 14308
rect 328 14248 392 14252
rect 328 14148 392 14152
rect 328 14092 332 14148
rect 332 14092 388 14148
rect 388 14092 392 14148
rect 328 14088 392 14092
rect 328 13988 392 13992
rect 328 13932 332 13988
rect 332 13932 388 13988
rect 388 13932 392 13988
rect 328 13928 392 13932
rect 328 13828 392 13832
rect 328 13772 332 13828
rect 332 13772 388 13828
rect 388 13772 392 13828
rect 328 13768 392 13772
rect 328 13668 392 13672
rect 328 13612 332 13668
rect 332 13612 388 13668
rect 388 13612 392 13668
rect 328 13608 392 13612
rect 328 13508 392 13512
rect 328 13452 332 13508
rect 332 13452 388 13508
rect 388 13452 392 13508
rect 328 13448 392 13452
rect 328 13348 392 13352
rect 328 13292 332 13348
rect 332 13292 388 13348
rect 388 13292 392 13348
rect 328 13288 392 13292
rect 328 13188 392 13192
rect 328 13132 332 13188
rect 332 13132 388 13188
rect 388 13132 392 13188
rect 328 13128 392 13132
rect 328 13028 392 13032
rect 328 12972 332 13028
rect 332 12972 388 13028
rect 388 12972 392 13028
rect 328 12968 392 12972
rect 328 12868 392 12872
rect 328 12812 332 12868
rect 332 12812 388 12868
rect 388 12812 392 12868
rect 328 12808 392 12812
rect 328 12708 392 12712
rect 328 12652 332 12708
rect 332 12652 388 12708
rect 388 12652 392 12708
rect 328 12648 392 12652
rect 328 12548 392 12552
rect 328 12492 332 12548
rect 332 12492 388 12548
rect 388 12492 392 12548
rect 328 12488 392 12492
rect 328 12388 392 12392
rect 328 12332 332 12388
rect 332 12332 388 12388
rect 388 12332 392 12388
rect 328 12328 392 12332
rect 328 12228 392 12232
rect 328 12172 332 12228
rect 332 12172 388 12228
rect 388 12172 392 12228
rect 328 12168 392 12172
rect 328 12068 392 12072
rect 328 12012 332 12068
rect 332 12012 388 12068
rect 388 12012 392 12068
rect 328 12008 392 12012
rect 328 11908 392 11912
rect 328 11852 332 11908
rect 332 11852 388 11908
rect 388 11852 392 11908
rect 328 11848 392 11852
rect 328 11748 392 11752
rect 328 11692 332 11748
rect 332 11692 388 11748
rect 388 11692 392 11748
rect 328 11688 392 11692
rect 328 11588 392 11592
rect 328 11532 332 11588
rect 332 11532 388 11588
rect 388 11532 392 11588
rect 328 11528 392 11532
rect 328 11428 392 11432
rect 328 11372 332 11428
rect 332 11372 388 11428
rect 388 11372 392 11428
rect 328 11368 392 11372
rect 328 11268 392 11272
rect 328 11212 332 11268
rect 332 11212 388 11268
rect 388 11212 392 11268
rect 328 11208 392 11212
rect 328 11108 392 11112
rect 328 11052 332 11108
rect 332 11052 388 11108
rect 388 11052 392 11108
rect 328 11048 392 11052
rect 328 10948 392 10952
rect 328 10892 332 10948
rect 332 10892 388 10948
rect 388 10892 392 10948
rect 328 10888 392 10892
rect 328 10788 392 10792
rect 328 10732 332 10788
rect 332 10732 388 10788
rect 388 10732 392 10788
rect 328 10728 392 10732
rect 328 10628 392 10632
rect 328 10572 332 10628
rect 332 10572 388 10628
rect 388 10572 392 10628
rect 328 10568 392 10572
rect 328 10468 392 10472
rect 328 10412 332 10468
rect 332 10412 388 10468
rect 388 10412 392 10468
rect 328 10408 392 10412
rect 328 10148 392 10152
rect 328 10092 332 10148
rect 332 10092 388 10148
rect 388 10092 392 10148
rect 328 10088 392 10092
rect 328 9988 392 9992
rect 328 9932 332 9988
rect 332 9932 388 9988
rect 388 9932 392 9988
rect 328 9928 392 9932
rect 328 9828 392 9832
rect 328 9772 332 9828
rect 332 9772 388 9828
rect 388 9772 392 9828
rect 328 9768 392 9772
rect 328 9668 392 9672
rect 328 9612 332 9668
rect 332 9612 388 9668
rect 388 9612 392 9668
rect 328 9608 392 9612
rect 328 9508 392 9512
rect 328 9452 332 9508
rect 332 9452 388 9508
rect 388 9452 392 9508
rect 328 9448 392 9452
rect 328 9348 392 9352
rect 328 9292 332 9348
rect 332 9292 388 9348
rect 388 9292 392 9348
rect 328 9288 392 9292
rect 328 9188 392 9192
rect 328 9132 332 9188
rect 332 9132 388 9188
rect 388 9132 392 9188
rect 328 9128 392 9132
rect 328 9028 392 9032
rect 328 8972 332 9028
rect 332 8972 388 9028
rect 388 8972 392 9028
rect 328 8968 392 8972
rect 328 8868 392 8872
rect 328 8812 332 8868
rect 332 8812 388 8868
rect 388 8812 392 8868
rect 328 8808 392 8812
rect 328 8708 392 8712
rect 328 8652 332 8708
rect 332 8652 388 8708
rect 388 8652 392 8708
rect 328 8648 392 8652
rect 328 8548 392 8552
rect 328 8492 332 8548
rect 332 8492 388 8548
rect 388 8492 392 8548
rect 328 8488 392 8492
rect 328 8388 392 8392
rect 328 8332 332 8388
rect 332 8332 388 8388
rect 388 8332 392 8388
rect 328 8328 392 8332
rect 328 8228 392 8232
rect 328 8172 332 8228
rect 332 8172 388 8228
rect 388 8172 392 8228
rect 328 8168 392 8172
rect 328 8068 392 8072
rect 328 8012 332 8068
rect 332 8012 388 8068
rect 388 8012 392 8068
rect 328 8008 392 8012
rect 328 7908 392 7912
rect 328 7852 332 7908
rect 332 7852 388 7908
rect 388 7852 392 7908
rect 328 7848 392 7852
rect 328 7748 392 7752
rect 328 7692 332 7748
rect 332 7692 388 7748
rect 388 7692 392 7748
rect 328 7688 392 7692
rect 328 7588 392 7592
rect 328 7532 332 7588
rect 332 7532 388 7588
rect 388 7532 392 7588
rect 328 7528 392 7532
rect 328 7428 392 7432
rect 328 7372 332 7428
rect 332 7372 388 7428
rect 388 7372 392 7428
rect 328 7368 392 7372
rect 328 7268 392 7272
rect 328 7212 332 7268
rect 332 7212 388 7268
rect 388 7212 392 7268
rect 328 7208 392 7212
rect 328 7108 392 7112
rect 328 7052 332 7108
rect 332 7052 388 7108
rect 388 7052 392 7108
rect 328 7048 392 7052
rect 328 6948 392 6952
rect 328 6892 332 6948
rect 332 6892 388 6948
rect 388 6892 392 6948
rect 328 6888 392 6892
rect 328 6788 392 6792
rect 328 6732 332 6788
rect 332 6732 388 6788
rect 388 6732 392 6788
rect 328 6728 392 6732
rect 328 6628 392 6632
rect 328 6572 332 6628
rect 332 6572 388 6628
rect 388 6572 392 6628
rect 328 6568 392 6572
rect 328 6468 392 6472
rect 328 6412 332 6468
rect 332 6412 388 6468
rect 388 6412 392 6468
rect 328 6408 392 6412
rect 328 6308 392 6312
rect 328 6252 332 6308
rect 332 6252 388 6308
rect 388 6252 392 6308
rect 328 6248 392 6252
rect 328 6148 392 6152
rect 328 6092 332 6148
rect 332 6092 388 6148
rect 388 6092 392 6148
rect 328 6088 392 6092
rect 328 5988 392 5992
rect 328 5932 332 5988
rect 332 5932 388 5988
rect 388 5932 392 5988
rect 328 5928 392 5932
rect 328 5828 392 5832
rect 328 5772 332 5828
rect 332 5772 388 5828
rect 388 5772 392 5828
rect 328 5768 392 5772
rect 328 5668 392 5672
rect 328 5612 332 5668
rect 332 5612 388 5668
rect 388 5612 392 5668
rect 328 5608 392 5612
rect 328 5508 392 5512
rect 328 5452 332 5508
rect 332 5452 388 5508
rect 388 5452 392 5508
rect 328 5448 392 5452
rect 328 5348 392 5352
rect 328 5292 332 5348
rect 332 5292 388 5348
rect 388 5292 392 5348
rect 328 5288 392 5292
rect 328 5188 392 5192
rect 328 5132 332 5188
rect 332 5132 388 5188
rect 388 5132 392 5188
rect 328 5128 392 5132
rect 328 5028 392 5032
rect 328 4972 332 5028
rect 332 4972 388 5028
rect 388 4972 392 5028
rect 328 4968 392 4972
rect 328 4868 392 4872
rect 328 4812 332 4868
rect 332 4812 388 4868
rect 388 4812 392 4868
rect 328 4808 392 4812
rect 328 4708 392 4712
rect 328 4652 332 4708
rect 332 4652 388 4708
rect 388 4652 392 4708
rect 328 4648 392 4652
rect 328 4548 392 4552
rect 328 4492 332 4548
rect 332 4492 388 4548
rect 388 4492 392 4548
rect 328 4488 392 4492
rect 328 4388 392 4392
rect 328 4332 332 4388
rect 332 4332 388 4388
rect 388 4332 392 4388
rect 328 4328 392 4332
rect 328 4228 392 4232
rect 328 4172 332 4228
rect 332 4172 388 4228
rect 388 4172 392 4228
rect 328 4168 392 4172
rect 328 4068 392 4072
rect 328 4012 332 4068
rect 332 4012 388 4068
rect 388 4012 392 4068
rect 328 4008 392 4012
rect 328 3908 392 3912
rect 328 3852 332 3908
rect 332 3852 388 3908
rect 388 3852 392 3908
rect 328 3848 392 3852
rect 328 3748 392 3752
rect 328 3692 332 3748
rect 332 3692 388 3748
rect 388 3692 392 3748
rect 328 3688 392 3692
rect 328 3588 392 3592
rect 328 3532 332 3588
rect 332 3532 388 3588
rect 388 3532 392 3588
rect 328 3528 392 3532
rect 328 3428 392 3432
rect 328 3372 332 3428
rect 332 3372 388 3428
rect 388 3372 392 3428
rect 328 3368 392 3372
rect 328 3268 392 3272
rect 328 3212 332 3268
rect 332 3212 388 3268
rect 388 3212 392 3268
rect 328 3208 392 3212
rect 328 3108 392 3112
rect 328 3052 332 3108
rect 332 3052 388 3108
rect 388 3052 392 3108
rect 328 3048 392 3052
rect 328 2948 392 2952
rect 328 2892 332 2948
rect 332 2892 388 2948
rect 388 2892 392 2948
rect 328 2888 392 2892
rect 328 2788 392 2792
rect 328 2732 332 2788
rect 332 2732 388 2788
rect 388 2732 392 2788
rect 328 2728 392 2732
rect 328 2628 392 2632
rect 328 2572 332 2628
rect 332 2572 388 2628
rect 388 2572 392 2628
rect 328 2568 392 2572
rect 328 2468 392 2472
rect 328 2412 332 2468
rect 332 2412 388 2468
rect 388 2412 392 2468
rect 328 2408 392 2412
rect 328 2308 392 2312
rect 328 2252 332 2308
rect 332 2252 388 2308
rect 388 2252 392 2308
rect 328 2248 392 2252
rect 328 2148 392 2152
rect 328 2092 332 2148
rect 332 2092 388 2148
rect 388 2092 392 2148
rect 328 2088 392 2092
rect 328 1988 392 1992
rect 328 1932 332 1988
rect 332 1932 388 1988
rect 388 1932 392 1988
rect 328 1928 392 1932
rect 328 1828 392 1832
rect 328 1772 332 1828
rect 332 1772 388 1828
rect 388 1772 392 1828
rect 328 1768 392 1772
rect 328 1668 392 1672
rect 328 1612 332 1668
rect 332 1612 388 1668
rect 388 1612 392 1668
rect 328 1608 392 1612
rect 328 1508 392 1512
rect 328 1452 332 1508
rect 332 1452 388 1508
rect 388 1452 392 1508
rect 328 1448 392 1452
rect 328 1348 392 1352
rect 328 1292 332 1348
rect 332 1292 388 1348
rect 388 1292 392 1348
rect 328 1288 392 1292
rect 328 1188 392 1192
rect 328 1132 332 1188
rect 332 1132 388 1188
rect 388 1132 392 1188
rect 328 1128 392 1132
rect 328 1028 392 1032
rect 328 972 332 1028
rect 332 972 388 1028
rect 388 972 392 1028
rect 328 968 392 972
rect 8 808 72 872
rect 8 728 72 792
rect 8 648 72 712
rect 8 568 72 632
rect 8 488 72 552
rect 488 22248 552 22312
rect 488 17128 552 17192
rect 488 15688 552 15752
rect 488 10568 552 10632
rect 648 31908 712 31912
rect 648 31852 652 31908
rect 652 31852 708 31908
rect 708 31852 712 31908
rect 648 31848 712 31852
rect 648 31748 712 31752
rect 648 31692 652 31748
rect 652 31692 708 31748
rect 708 31692 712 31748
rect 648 31688 712 31692
rect 648 31588 712 31592
rect 648 31532 652 31588
rect 652 31532 708 31588
rect 708 31532 712 31588
rect 648 31528 712 31532
rect 648 31428 712 31432
rect 648 31372 652 31428
rect 652 31372 708 31428
rect 708 31372 712 31428
rect 648 31368 712 31372
rect 648 31268 712 31272
rect 648 31212 652 31268
rect 652 31212 708 31268
rect 708 31212 712 31268
rect 648 31208 712 31212
rect 648 31108 712 31112
rect 648 31052 652 31108
rect 652 31052 708 31108
rect 708 31052 712 31108
rect 648 31048 712 31052
rect 648 30948 712 30952
rect 648 30892 652 30948
rect 652 30892 708 30948
rect 708 30892 712 30948
rect 648 30888 712 30892
rect 648 30788 712 30792
rect 648 30732 652 30788
rect 652 30732 708 30788
rect 708 30732 712 30788
rect 648 30728 712 30732
rect 648 30628 712 30632
rect 648 30572 652 30628
rect 652 30572 708 30628
rect 708 30572 712 30628
rect 648 30568 712 30572
rect 648 30468 712 30472
rect 648 30412 652 30468
rect 652 30412 708 30468
rect 708 30412 712 30468
rect 648 30408 712 30412
rect 648 30308 712 30312
rect 648 30252 652 30308
rect 652 30252 708 30308
rect 708 30252 712 30308
rect 648 30248 712 30252
rect 648 30148 712 30152
rect 648 30092 652 30148
rect 652 30092 708 30148
rect 708 30092 712 30148
rect 648 30088 712 30092
rect 648 29988 712 29992
rect 648 29932 652 29988
rect 652 29932 708 29988
rect 708 29932 712 29988
rect 648 29928 712 29932
rect 648 29828 712 29832
rect 648 29772 652 29828
rect 652 29772 708 29828
rect 708 29772 712 29828
rect 648 29768 712 29772
rect 648 29668 712 29672
rect 648 29612 652 29668
rect 652 29612 708 29668
rect 708 29612 712 29668
rect 648 29608 712 29612
rect 648 29508 712 29512
rect 648 29452 652 29508
rect 652 29452 708 29508
rect 708 29452 712 29508
rect 648 29448 712 29452
rect 648 29348 712 29352
rect 648 29292 652 29348
rect 652 29292 708 29348
rect 708 29292 712 29348
rect 648 29288 712 29292
rect 648 29188 712 29192
rect 648 29132 652 29188
rect 652 29132 708 29188
rect 708 29132 712 29188
rect 648 29128 712 29132
rect 648 29028 712 29032
rect 648 28972 652 29028
rect 652 28972 708 29028
rect 708 28972 712 29028
rect 648 28968 712 28972
rect 648 28868 712 28872
rect 648 28812 652 28868
rect 652 28812 708 28868
rect 708 28812 712 28868
rect 648 28808 712 28812
rect 648 28708 712 28712
rect 648 28652 652 28708
rect 652 28652 708 28708
rect 708 28652 712 28708
rect 648 28648 712 28652
rect 648 28548 712 28552
rect 648 28492 652 28548
rect 652 28492 708 28548
rect 708 28492 712 28548
rect 648 28488 712 28492
rect 648 28388 712 28392
rect 648 28332 652 28388
rect 652 28332 708 28388
rect 708 28332 712 28388
rect 648 28328 712 28332
rect 648 28228 712 28232
rect 648 28172 652 28228
rect 652 28172 708 28228
rect 708 28172 712 28228
rect 648 28168 712 28172
rect 648 28068 712 28072
rect 648 28012 652 28068
rect 652 28012 708 28068
rect 708 28012 712 28068
rect 648 28008 712 28012
rect 648 27908 712 27912
rect 648 27852 652 27908
rect 652 27852 708 27908
rect 708 27852 712 27908
rect 648 27848 712 27852
rect 648 27748 712 27752
rect 648 27692 652 27748
rect 652 27692 708 27748
rect 708 27692 712 27748
rect 648 27688 712 27692
rect 648 27588 712 27592
rect 648 27532 652 27588
rect 652 27532 708 27588
rect 708 27532 712 27588
rect 648 27528 712 27532
rect 648 27428 712 27432
rect 648 27372 652 27428
rect 652 27372 708 27428
rect 708 27372 712 27428
rect 648 27368 712 27372
rect 648 27268 712 27272
rect 648 27212 652 27268
rect 652 27212 708 27268
rect 708 27212 712 27268
rect 648 27208 712 27212
rect 648 27108 712 27112
rect 648 27052 652 27108
rect 652 27052 708 27108
rect 708 27052 712 27108
rect 648 27048 712 27052
rect 648 26948 712 26952
rect 648 26892 652 26948
rect 652 26892 708 26948
rect 708 26892 712 26948
rect 648 26888 712 26892
rect 648 26788 712 26792
rect 648 26732 652 26788
rect 652 26732 708 26788
rect 708 26732 712 26788
rect 648 26728 712 26732
rect 648 26628 712 26632
rect 648 26572 652 26628
rect 652 26572 708 26628
rect 708 26572 712 26628
rect 648 26568 712 26572
rect 648 26468 712 26472
rect 648 26412 652 26468
rect 652 26412 708 26468
rect 708 26412 712 26468
rect 648 26408 712 26412
rect 648 26308 712 26312
rect 648 26252 652 26308
rect 652 26252 708 26308
rect 708 26252 712 26308
rect 648 26248 712 26252
rect 648 26148 712 26152
rect 648 26092 652 26148
rect 652 26092 708 26148
rect 708 26092 712 26148
rect 648 26088 712 26092
rect 648 25988 712 25992
rect 648 25932 652 25988
rect 652 25932 708 25988
rect 708 25932 712 25988
rect 648 25928 712 25932
rect 648 25828 712 25832
rect 648 25772 652 25828
rect 652 25772 708 25828
rect 708 25772 712 25828
rect 648 25768 712 25772
rect 648 25668 712 25672
rect 648 25612 652 25668
rect 652 25612 708 25668
rect 708 25612 712 25668
rect 648 25608 712 25612
rect 648 25508 712 25512
rect 648 25452 652 25508
rect 652 25452 708 25508
rect 708 25452 712 25508
rect 648 25448 712 25452
rect 648 25348 712 25352
rect 648 25292 652 25348
rect 652 25292 708 25348
rect 708 25292 712 25348
rect 648 25288 712 25292
rect 648 25188 712 25192
rect 648 25132 652 25188
rect 652 25132 708 25188
rect 708 25132 712 25188
rect 648 25128 712 25132
rect 648 25028 712 25032
rect 648 24972 652 25028
rect 652 24972 708 25028
rect 708 24972 712 25028
rect 648 24968 712 24972
rect 648 24868 712 24872
rect 648 24812 652 24868
rect 652 24812 708 24868
rect 708 24812 712 24868
rect 648 24808 712 24812
rect 648 24708 712 24712
rect 648 24652 652 24708
rect 652 24652 708 24708
rect 708 24652 712 24708
rect 648 24648 712 24652
rect 648 24548 712 24552
rect 648 24492 652 24548
rect 652 24492 708 24548
rect 708 24492 712 24548
rect 648 24488 712 24492
rect 648 24388 712 24392
rect 648 24332 652 24388
rect 652 24332 708 24388
rect 708 24332 712 24388
rect 648 24328 712 24332
rect 648 24228 712 24232
rect 648 24172 652 24228
rect 652 24172 708 24228
rect 708 24172 712 24228
rect 648 24168 712 24172
rect 648 24068 712 24072
rect 648 24012 652 24068
rect 652 24012 708 24068
rect 708 24012 712 24068
rect 648 24008 712 24012
rect 648 23908 712 23912
rect 648 23852 652 23908
rect 652 23852 708 23908
rect 708 23852 712 23908
rect 648 23848 712 23852
rect 648 23748 712 23752
rect 648 23692 652 23748
rect 652 23692 708 23748
rect 708 23692 712 23748
rect 648 23688 712 23692
rect 648 23588 712 23592
rect 648 23532 652 23588
rect 652 23532 708 23588
rect 708 23532 712 23588
rect 648 23528 712 23532
rect 648 23428 712 23432
rect 648 23372 652 23428
rect 652 23372 708 23428
rect 708 23372 712 23428
rect 648 23368 712 23372
rect 648 23268 712 23272
rect 648 23212 652 23268
rect 652 23212 708 23268
rect 708 23212 712 23268
rect 648 23208 712 23212
rect 648 23108 712 23112
rect 648 23052 652 23108
rect 652 23052 708 23108
rect 708 23052 712 23108
rect 648 23048 712 23052
rect 648 22948 712 22952
rect 648 22892 652 22948
rect 652 22892 708 22948
rect 708 22892 712 22948
rect 648 22888 712 22892
rect 648 22788 712 22792
rect 648 22732 652 22788
rect 652 22732 708 22788
rect 708 22732 712 22788
rect 648 22728 712 22732
rect 648 22468 712 22472
rect 648 22412 652 22468
rect 652 22412 708 22468
rect 708 22412 712 22468
rect 648 22408 712 22412
rect 648 22148 712 22152
rect 648 22092 652 22148
rect 652 22092 708 22148
rect 708 22092 712 22148
rect 648 22088 712 22092
rect 648 21988 712 21992
rect 648 21932 652 21988
rect 652 21932 708 21988
rect 708 21932 712 21988
rect 648 21928 712 21932
rect 648 21828 712 21832
rect 648 21772 652 21828
rect 652 21772 708 21828
rect 708 21772 712 21828
rect 648 21768 712 21772
rect 648 21668 712 21672
rect 648 21612 652 21668
rect 652 21612 708 21668
rect 708 21612 712 21668
rect 648 21608 712 21612
rect 648 21508 712 21512
rect 648 21452 652 21508
rect 652 21452 708 21508
rect 708 21452 712 21508
rect 648 21448 712 21452
rect 648 21348 712 21352
rect 648 21292 652 21348
rect 652 21292 708 21348
rect 708 21292 712 21348
rect 648 21288 712 21292
rect 648 21188 712 21192
rect 648 21132 652 21188
rect 652 21132 708 21188
rect 708 21132 712 21188
rect 648 21128 712 21132
rect 648 21028 712 21032
rect 648 20972 652 21028
rect 652 20972 708 21028
rect 708 20972 712 21028
rect 648 20968 712 20972
rect 648 20868 712 20872
rect 648 20812 652 20868
rect 652 20812 708 20868
rect 708 20812 712 20868
rect 648 20808 712 20812
rect 648 20708 712 20712
rect 648 20652 652 20708
rect 652 20652 708 20708
rect 708 20652 712 20708
rect 648 20648 712 20652
rect 648 20548 712 20552
rect 648 20492 652 20548
rect 652 20492 708 20548
rect 708 20492 712 20548
rect 648 20488 712 20492
rect 648 20388 712 20392
rect 648 20332 652 20388
rect 652 20332 708 20388
rect 708 20332 712 20388
rect 648 20328 712 20332
rect 648 20228 712 20232
rect 648 20172 652 20228
rect 652 20172 708 20228
rect 708 20172 712 20228
rect 648 20168 712 20172
rect 648 20068 712 20072
rect 648 20012 652 20068
rect 652 20012 708 20068
rect 708 20012 712 20068
rect 648 20008 712 20012
rect 648 19908 712 19912
rect 648 19852 652 19908
rect 652 19852 708 19908
rect 708 19852 712 19908
rect 648 19848 712 19852
rect 648 19748 712 19752
rect 648 19692 652 19748
rect 652 19692 708 19748
rect 708 19692 712 19748
rect 648 19688 712 19692
rect 648 19588 712 19592
rect 648 19532 652 19588
rect 652 19532 708 19588
rect 708 19532 712 19588
rect 648 19528 712 19532
rect 648 19428 712 19432
rect 648 19372 652 19428
rect 652 19372 708 19428
rect 708 19372 712 19428
rect 648 19368 712 19372
rect 648 19268 712 19272
rect 648 19212 652 19268
rect 652 19212 708 19268
rect 708 19212 712 19268
rect 648 19208 712 19212
rect 648 19108 712 19112
rect 648 19052 652 19108
rect 652 19052 708 19108
rect 708 19052 712 19108
rect 648 19048 712 19052
rect 648 18948 712 18952
rect 648 18892 652 18948
rect 652 18892 708 18948
rect 708 18892 712 18948
rect 648 18888 712 18892
rect 648 18788 712 18792
rect 648 18732 652 18788
rect 652 18732 708 18788
rect 708 18732 712 18788
rect 648 18728 712 18732
rect 648 18628 712 18632
rect 648 18572 652 18628
rect 652 18572 708 18628
rect 708 18572 712 18628
rect 648 18568 712 18572
rect 648 18468 712 18472
rect 648 18412 652 18468
rect 652 18412 708 18468
rect 708 18412 712 18468
rect 648 18408 712 18412
rect 648 18308 712 18312
rect 648 18252 652 18308
rect 652 18252 708 18308
rect 708 18252 712 18308
rect 648 18248 712 18252
rect 648 18148 712 18152
rect 648 18092 652 18148
rect 652 18092 708 18148
rect 708 18092 712 18148
rect 648 18088 712 18092
rect 648 17988 712 17992
rect 648 17932 652 17988
rect 652 17932 708 17988
rect 708 17932 712 17988
rect 648 17928 712 17932
rect 648 17828 712 17832
rect 648 17772 652 17828
rect 652 17772 708 17828
rect 708 17772 712 17828
rect 648 17768 712 17772
rect 648 17668 712 17672
rect 648 17612 652 17668
rect 652 17612 708 17668
rect 708 17612 712 17668
rect 648 17608 712 17612
rect 648 17508 712 17512
rect 648 17452 652 17508
rect 652 17452 708 17508
rect 708 17452 712 17508
rect 648 17448 712 17452
rect 648 17348 712 17352
rect 648 17292 652 17348
rect 652 17292 708 17348
rect 708 17292 712 17348
rect 648 17288 712 17292
rect 648 17028 712 17032
rect 648 16972 652 17028
rect 652 16972 708 17028
rect 708 16972 712 17028
rect 648 16968 712 16972
rect 648 16708 712 16712
rect 648 16652 652 16708
rect 652 16652 708 16708
rect 708 16652 712 16708
rect 648 16648 712 16652
rect 648 16548 712 16552
rect 648 16492 652 16548
rect 652 16492 708 16548
rect 708 16492 712 16548
rect 648 16488 712 16492
rect 648 16388 712 16392
rect 648 16332 652 16388
rect 652 16332 708 16388
rect 708 16332 712 16388
rect 648 16328 712 16332
rect 648 16228 712 16232
rect 648 16172 652 16228
rect 652 16172 708 16228
rect 708 16172 712 16228
rect 648 16168 712 16172
rect 648 15908 712 15912
rect 648 15852 652 15908
rect 652 15852 708 15908
rect 708 15852 712 15908
rect 648 15848 712 15852
rect 648 15588 712 15592
rect 648 15532 652 15588
rect 652 15532 708 15588
rect 708 15532 712 15588
rect 648 15528 712 15532
rect 648 15428 712 15432
rect 648 15372 652 15428
rect 652 15372 708 15428
rect 708 15372 712 15428
rect 648 15368 712 15372
rect 648 15268 712 15272
rect 648 15212 652 15268
rect 652 15212 708 15268
rect 708 15212 712 15268
rect 648 15208 712 15212
rect 648 15108 712 15112
rect 648 15052 652 15108
rect 652 15052 708 15108
rect 708 15052 712 15108
rect 648 15048 712 15052
rect 648 14948 712 14952
rect 648 14892 652 14948
rect 652 14892 708 14948
rect 708 14892 712 14948
rect 648 14888 712 14892
rect 648 14788 712 14792
rect 648 14732 652 14788
rect 652 14732 708 14788
rect 708 14732 712 14788
rect 648 14728 712 14732
rect 648 14628 712 14632
rect 648 14572 652 14628
rect 652 14572 708 14628
rect 708 14572 712 14628
rect 648 14568 712 14572
rect 648 14468 712 14472
rect 648 14412 652 14468
rect 652 14412 708 14468
rect 708 14412 712 14468
rect 648 14408 712 14412
rect 648 14308 712 14312
rect 648 14252 652 14308
rect 652 14252 708 14308
rect 708 14252 712 14308
rect 648 14248 712 14252
rect 648 14148 712 14152
rect 648 14092 652 14148
rect 652 14092 708 14148
rect 708 14092 712 14148
rect 648 14088 712 14092
rect 648 13988 712 13992
rect 648 13932 652 13988
rect 652 13932 708 13988
rect 708 13932 712 13988
rect 648 13928 712 13932
rect 648 13828 712 13832
rect 648 13772 652 13828
rect 652 13772 708 13828
rect 708 13772 712 13828
rect 648 13768 712 13772
rect 648 13668 712 13672
rect 648 13612 652 13668
rect 652 13612 708 13668
rect 708 13612 712 13668
rect 648 13608 712 13612
rect 648 13508 712 13512
rect 648 13452 652 13508
rect 652 13452 708 13508
rect 708 13452 712 13508
rect 648 13448 712 13452
rect 648 13348 712 13352
rect 648 13292 652 13348
rect 652 13292 708 13348
rect 708 13292 712 13348
rect 648 13288 712 13292
rect 648 13188 712 13192
rect 648 13132 652 13188
rect 652 13132 708 13188
rect 708 13132 712 13188
rect 648 13128 712 13132
rect 648 13028 712 13032
rect 648 12972 652 13028
rect 652 12972 708 13028
rect 708 12972 712 13028
rect 648 12968 712 12972
rect 648 12868 712 12872
rect 648 12812 652 12868
rect 652 12812 708 12868
rect 708 12812 712 12868
rect 648 12808 712 12812
rect 648 12708 712 12712
rect 648 12652 652 12708
rect 652 12652 708 12708
rect 708 12652 712 12708
rect 648 12648 712 12652
rect 648 12548 712 12552
rect 648 12492 652 12548
rect 652 12492 708 12548
rect 708 12492 712 12548
rect 648 12488 712 12492
rect 648 12388 712 12392
rect 648 12332 652 12388
rect 652 12332 708 12388
rect 708 12332 712 12388
rect 648 12328 712 12332
rect 648 12228 712 12232
rect 648 12172 652 12228
rect 652 12172 708 12228
rect 708 12172 712 12228
rect 648 12168 712 12172
rect 648 12068 712 12072
rect 648 12012 652 12068
rect 652 12012 708 12068
rect 708 12012 712 12068
rect 648 12008 712 12012
rect 648 11908 712 11912
rect 648 11852 652 11908
rect 652 11852 708 11908
rect 708 11852 712 11908
rect 648 11848 712 11852
rect 648 11748 712 11752
rect 648 11692 652 11748
rect 652 11692 708 11748
rect 708 11692 712 11748
rect 648 11688 712 11692
rect 648 11588 712 11592
rect 648 11532 652 11588
rect 652 11532 708 11588
rect 708 11532 712 11588
rect 648 11528 712 11532
rect 648 11428 712 11432
rect 648 11372 652 11428
rect 652 11372 708 11428
rect 708 11372 712 11428
rect 648 11368 712 11372
rect 648 11268 712 11272
rect 648 11212 652 11268
rect 652 11212 708 11268
rect 708 11212 712 11268
rect 648 11208 712 11212
rect 648 11108 712 11112
rect 648 11052 652 11108
rect 652 11052 708 11108
rect 708 11052 712 11108
rect 648 11048 712 11052
rect 648 10948 712 10952
rect 648 10892 652 10948
rect 652 10892 708 10948
rect 708 10892 712 10948
rect 648 10888 712 10892
rect 648 10788 712 10792
rect 648 10732 652 10788
rect 652 10732 708 10788
rect 708 10732 712 10788
rect 648 10728 712 10732
rect 648 10468 712 10472
rect 648 10412 652 10468
rect 652 10412 708 10468
rect 708 10412 712 10468
rect 648 10408 712 10412
rect 648 10148 712 10152
rect 648 10092 652 10148
rect 652 10092 708 10148
rect 708 10092 712 10148
rect 648 10088 712 10092
rect 648 9988 712 9992
rect 648 9932 652 9988
rect 652 9932 708 9988
rect 708 9932 712 9988
rect 648 9928 712 9932
rect 648 9828 712 9832
rect 648 9772 652 9828
rect 652 9772 708 9828
rect 708 9772 712 9828
rect 648 9768 712 9772
rect 648 9668 712 9672
rect 648 9612 652 9668
rect 652 9612 708 9668
rect 708 9612 712 9668
rect 648 9608 712 9612
rect 648 9508 712 9512
rect 648 9452 652 9508
rect 652 9452 708 9508
rect 708 9452 712 9508
rect 648 9448 712 9452
rect 648 9348 712 9352
rect 648 9292 652 9348
rect 652 9292 708 9348
rect 708 9292 712 9348
rect 648 9288 712 9292
rect 648 9188 712 9192
rect 648 9132 652 9188
rect 652 9132 708 9188
rect 708 9132 712 9188
rect 648 9128 712 9132
rect 648 9028 712 9032
rect 648 8972 652 9028
rect 652 8972 708 9028
rect 708 8972 712 9028
rect 648 8968 712 8972
rect 648 8868 712 8872
rect 648 8812 652 8868
rect 652 8812 708 8868
rect 708 8812 712 8868
rect 648 8808 712 8812
rect 648 8708 712 8712
rect 648 8652 652 8708
rect 652 8652 708 8708
rect 708 8652 712 8708
rect 648 8648 712 8652
rect 648 8548 712 8552
rect 648 8492 652 8548
rect 652 8492 708 8548
rect 708 8492 712 8548
rect 648 8488 712 8492
rect 648 8388 712 8392
rect 648 8332 652 8388
rect 652 8332 708 8388
rect 708 8332 712 8388
rect 648 8328 712 8332
rect 648 8228 712 8232
rect 648 8172 652 8228
rect 652 8172 708 8228
rect 708 8172 712 8228
rect 648 8168 712 8172
rect 648 8068 712 8072
rect 648 8012 652 8068
rect 652 8012 708 8068
rect 708 8012 712 8068
rect 648 8008 712 8012
rect 648 7908 712 7912
rect 648 7852 652 7908
rect 652 7852 708 7908
rect 708 7852 712 7908
rect 648 7848 712 7852
rect 648 7748 712 7752
rect 648 7692 652 7748
rect 652 7692 708 7748
rect 708 7692 712 7748
rect 648 7688 712 7692
rect 648 7588 712 7592
rect 648 7532 652 7588
rect 652 7532 708 7588
rect 708 7532 712 7588
rect 648 7528 712 7532
rect 648 7428 712 7432
rect 648 7372 652 7428
rect 652 7372 708 7428
rect 708 7372 712 7428
rect 648 7368 712 7372
rect 648 7268 712 7272
rect 648 7212 652 7268
rect 652 7212 708 7268
rect 708 7212 712 7268
rect 648 7208 712 7212
rect 648 7108 712 7112
rect 648 7052 652 7108
rect 652 7052 708 7108
rect 708 7052 712 7108
rect 648 7048 712 7052
rect 648 6948 712 6952
rect 648 6892 652 6948
rect 652 6892 708 6948
rect 708 6892 712 6948
rect 648 6888 712 6892
rect 648 6788 712 6792
rect 648 6732 652 6788
rect 652 6732 708 6788
rect 708 6732 712 6788
rect 648 6728 712 6732
rect 648 6628 712 6632
rect 648 6572 652 6628
rect 652 6572 708 6628
rect 708 6572 712 6628
rect 648 6568 712 6572
rect 648 6468 712 6472
rect 648 6412 652 6468
rect 652 6412 708 6468
rect 708 6412 712 6468
rect 648 6408 712 6412
rect 648 6308 712 6312
rect 648 6252 652 6308
rect 652 6252 708 6308
rect 708 6252 712 6308
rect 648 6248 712 6252
rect 648 6148 712 6152
rect 648 6092 652 6148
rect 652 6092 708 6148
rect 708 6092 712 6148
rect 648 6088 712 6092
rect 648 5988 712 5992
rect 648 5932 652 5988
rect 652 5932 708 5988
rect 708 5932 712 5988
rect 648 5928 712 5932
rect 648 5828 712 5832
rect 648 5772 652 5828
rect 652 5772 708 5828
rect 708 5772 712 5828
rect 648 5768 712 5772
rect 648 5668 712 5672
rect 648 5612 652 5668
rect 652 5612 708 5668
rect 708 5612 712 5668
rect 648 5608 712 5612
rect 648 5508 712 5512
rect 648 5452 652 5508
rect 652 5452 708 5508
rect 708 5452 712 5508
rect 648 5448 712 5452
rect 648 5348 712 5352
rect 648 5292 652 5348
rect 652 5292 708 5348
rect 708 5292 712 5348
rect 648 5288 712 5292
rect 648 5188 712 5192
rect 648 5132 652 5188
rect 652 5132 708 5188
rect 708 5132 712 5188
rect 648 5128 712 5132
rect 648 5028 712 5032
rect 648 4972 652 5028
rect 652 4972 708 5028
rect 708 4972 712 5028
rect 648 4968 712 4972
rect 648 4868 712 4872
rect 648 4812 652 4868
rect 652 4812 708 4868
rect 708 4812 712 4868
rect 648 4808 712 4812
rect 648 4708 712 4712
rect 648 4652 652 4708
rect 652 4652 708 4708
rect 708 4652 712 4708
rect 648 4648 712 4652
rect 648 4548 712 4552
rect 648 4492 652 4548
rect 652 4492 708 4548
rect 708 4492 712 4548
rect 648 4488 712 4492
rect 648 4388 712 4392
rect 648 4332 652 4388
rect 652 4332 708 4388
rect 708 4332 712 4388
rect 648 4328 712 4332
rect 648 4228 712 4232
rect 648 4172 652 4228
rect 652 4172 708 4228
rect 708 4172 712 4228
rect 648 4168 712 4172
rect 648 4068 712 4072
rect 648 4012 652 4068
rect 652 4012 708 4068
rect 708 4012 712 4068
rect 648 4008 712 4012
rect 648 3908 712 3912
rect 648 3852 652 3908
rect 652 3852 708 3908
rect 708 3852 712 3908
rect 648 3848 712 3852
rect 648 3748 712 3752
rect 648 3692 652 3748
rect 652 3692 708 3748
rect 708 3692 712 3748
rect 648 3688 712 3692
rect 648 3588 712 3592
rect 648 3532 652 3588
rect 652 3532 708 3588
rect 708 3532 712 3588
rect 648 3528 712 3532
rect 648 3428 712 3432
rect 648 3372 652 3428
rect 652 3372 708 3428
rect 708 3372 712 3428
rect 648 3368 712 3372
rect 648 3268 712 3272
rect 648 3212 652 3268
rect 652 3212 708 3268
rect 708 3212 712 3268
rect 648 3208 712 3212
rect 648 3108 712 3112
rect 648 3052 652 3108
rect 652 3052 708 3108
rect 708 3052 712 3108
rect 648 3048 712 3052
rect 648 2948 712 2952
rect 648 2892 652 2948
rect 652 2892 708 2948
rect 708 2892 712 2948
rect 648 2888 712 2892
rect 648 2788 712 2792
rect 648 2732 652 2788
rect 652 2732 708 2788
rect 708 2732 712 2788
rect 648 2728 712 2732
rect 648 2628 712 2632
rect 648 2572 652 2628
rect 652 2572 708 2628
rect 708 2572 712 2628
rect 648 2568 712 2572
rect 648 2468 712 2472
rect 648 2412 652 2468
rect 652 2412 708 2468
rect 708 2412 712 2468
rect 648 2408 712 2412
rect 648 2308 712 2312
rect 648 2252 652 2308
rect 652 2252 708 2308
rect 708 2252 712 2308
rect 648 2248 712 2252
rect 648 2148 712 2152
rect 648 2092 652 2148
rect 652 2092 708 2148
rect 708 2092 712 2148
rect 648 2088 712 2092
rect 648 1988 712 1992
rect 648 1932 652 1988
rect 652 1932 708 1988
rect 708 1932 712 1988
rect 648 1928 712 1932
rect 648 1828 712 1832
rect 648 1772 652 1828
rect 652 1772 708 1828
rect 708 1772 712 1828
rect 648 1768 712 1772
rect 648 1668 712 1672
rect 648 1612 652 1668
rect 652 1612 708 1668
rect 708 1612 712 1668
rect 648 1608 712 1612
rect 648 1508 712 1512
rect 648 1452 652 1508
rect 652 1452 708 1508
rect 708 1452 712 1508
rect 648 1448 712 1452
rect 648 1348 712 1352
rect 648 1292 652 1348
rect 652 1292 708 1348
rect 708 1292 712 1348
rect 648 1288 712 1292
rect 648 1188 712 1192
rect 648 1132 652 1188
rect 652 1132 708 1188
rect 708 1132 712 1188
rect 648 1128 712 1132
rect 648 1028 712 1032
rect 648 972 652 1028
rect 652 972 708 1028
rect 708 972 712 1028
rect 648 968 712 972
rect 328 808 392 872
rect 328 728 392 792
rect 328 648 392 712
rect 328 568 392 632
rect 328 488 392 552
rect 808 19688 872 19752
rect 808 13128 872 13192
rect 968 31908 1032 31912
rect 968 31852 972 31908
rect 972 31852 1028 31908
rect 1028 31852 1032 31908
rect 968 31848 1032 31852
rect 968 31748 1032 31752
rect 968 31692 972 31748
rect 972 31692 1028 31748
rect 1028 31692 1032 31748
rect 968 31688 1032 31692
rect 968 31588 1032 31592
rect 968 31532 972 31588
rect 972 31532 1028 31588
rect 1028 31532 1032 31588
rect 968 31528 1032 31532
rect 968 31428 1032 31432
rect 968 31372 972 31428
rect 972 31372 1028 31428
rect 1028 31372 1032 31428
rect 968 31368 1032 31372
rect 968 31268 1032 31272
rect 968 31212 972 31268
rect 972 31212 1028 31268
rect 1028 31212 1032 31268
rect 968 31208 1032 31212
rect 968 31108 1032 31112
rect 968 31052 972 31108
rect 972 31052 1028 31108
rect 1028 31052 1032 31108
rect 968 31048 1032 31052
rect 968 30948 1032 30952
rect 968 30892 972 30948
rect 972 30892 1028 30948
rect 1028 30892 1032 30948
rect 968 30888 1032 30892
rect 968 30788 1032 30792
rect 968 30732 972 30788
rect 972 30732 1028 30788
rect 1028 30732 1032 30788
rect 968 30728 1032 30732
rect 968 30628 1032 30632
rect 968 30572 972 30628
rect 972 30572 1028 30628
rect 1028 30572 1032 30628
rect 968 30568 1032 30572
rect 968 30468 1032 30472
rect 968 30412 972 30468
rect 972 30412 1028 30468
rect 1028 30412 1032 30468
rect 968 30408 1032 30412
rect 968 30308 1032 30312
rect 968 30252 972 30308
rect 972 30252 1028 30308
rect 1028 30252 1032 30308
rect 968 30248 1032 30252
rect 968 30148 1032 30152
rect 968 30092 972 30148
rect 972 30092 1028 30148
rect 1028 30092 1032 30148
rect 968 30088 1032 30092
rect 968 29988 1032 29992
rect 968 29932 972 29988
rect 972 29932 1028 29988
rect 1028 29932 1032 29988
rect 968 29928 1032 29932
rect 968 29828 1032 29832
rect 968 29772 972 29828
rect 972 29772 1028 29828
rect 1028 29772 1032 29828
rect 968 29768 1032 29772
rect 968 29668 1032 29672
rect 968 29612 972 29668
rect 972 29612 1028 29668
rect 1028 29612 1032 29668
rect 968 29608 1032 29612
rect 968 29508 1032 29512
rect 968 29452 972 29508
rect 972 29452 1028 29508
rect 1028 29452 1032 29508
rect 968 29448 1032 29452
rect 968 29348 1032 29352
rect 968 29292 972 29348
rect 972 29292 1028 29348
rect 1028 29292 1032 29348
rect 968 29288 1032 29292
rect 968 29188 1032 29192
rect 968 29132 972 29188
rect 972 29132 1028 29188
rect 1028 29132 1032 29188
rect 968 29128 1032 29132
rect 968 29028 1032 29032
rect 968 28972 972 29028
rect 972 28972 1028 29028
rect 1028 28972 1032 29028
rect 968 28968 1032 28972
rect 968 28868 1032 28872
rect 968 28812 972 28868
rect 972 28812 1028 28868
rect 1028 28812 1032 28868
rect 968 28808 1032 28812
rect 968 28708 1032 28712
rect 968 28652 972 28708
rect 972 28652 1028 28708
rect 1028 28652 1032 28708
rect 968 28648 1032 28652
rect 968 28548 1032 28552
rect 968 28492 972 28548
rect 972 28492 1028 28548
rect 1028 28492 1032 28548
rect 968 28488 1032 28492
rect 968 28388 1032 28392
rect 968 28332 972 28388
rect 972 28332 1028 28388
rect 1028 28332 1032 28388
rect 968 28328 1032 28332
rect 968 28228 1032 28232
rect 968 28172 972 28228
rect 972 28172 1028 28228
rect 1028 28172 1032 28228
rect 968 28168 1032 28172
rect 968 28068 1032 28072
rect 968 28012 972 28068
rect 972 28012 1028 28068
rect 1028 28012 1032 28068
rect 968 28008 1032 28012
rect 968 27908 1032 27912
rect 968 27852 972 27908
rect 972 27852 1028 27908
rect 1028 27852 1032 27908
rect 968 27848 1032 27852
rect 968 27748 1032 27752
rect 968 27692 972 27748
rect 972 27692 1028 27748
rect 1028 27692 1032 27748
rect 968 27688 1032 27692
rect 968 27588 1032 27592
rect 968 27532 972 27588
rect 972 27532 1028 27588
rect 1028 27532 1032 27588
rect 968 27528 1032 27532
rect 968 27428 1032 27432
rect 968 27372 972 27428
rect 972 27372 1028 27428
rect 1028 27372 1032 27428
rect 968 27368 1032 27372
rect 968 27268 1032 27272
rect 968 27212 972 27268
rect 972 27212 1028 27268
rect 1028 27212 1032 27268
rect 968 27208 1032 27212
rect 968 27108 1032 27112
rect 968 27052 972 27108
rect 972 27052 1028 27108
rect 1028 27052 1032 27108
rect 968 27048 1032 27052
rect 968 26948 1032 26952
rect 968 26892 972 26948
rect 972 26892 1028 26948
rect 1028 26892 1032 26948
rect 968 26888 1032 26892
rect 968 26788 1032 26792
rect 968 26732 972 26788
rect 972 26732 1028 26788
rect 1028 26732 1032 26788
rect 968 26728 1032 26732
rect 968 26628 1032 26632
rect 968 26572 972 26628
rect 972 26572 1028 26628
rect 1028 26572 1032 26628
rect 968 26568 1032 26572
rect 968 26468 1032 26472
rect 968 26412 972 26468
rect 972 26412 1028 26468
rect 1028 26412 1032 26468
rect 968 26408 1032 26412
rect 968 26308 1032 26312
rect 968 26252 972 26308
rect 972 26252 1028 26308
rect 1028 26252 1032 26308
rect 968 26248 1032 26252
rect 968 26148 1032 26152
rect 968 26092 972 26148
rect 972 26092 1028 26148
rect 1028 26092 1032 26148
rect 968 26088 1032 26092
rect 968 25988 1032 25992
rect 968 25932 972 25988
rect 972 25932 1028 25988
rect 1028 25932 1032 25988
rect 968 25928 1032 25932
rect 968 25828 1032 25832
rect 968 25772 972 25828
rect 972 25772 1028 25828
rect 1028 25772 1032 25828
rect 968 25768 1032 25772
rect 968 25668 1032 25672
rect 968 25612 972 25668
rect 972 25612 1028 25668
rect 1028 25612 1032 25668
rect 968 25608 1032 25612
rect 968 25508 1032 25512
rect 968 25452 972 25508
rect 972 25452 1028 25508
rect 1028 25452 1032 25508
rect 968 25448 1032 25452
rect 968 25348 1032 25352
rect 968 25292 972 25348
rect 972 25292 1028 25348
rect 1028 25292 1032 25348
rect 968 25288 1032 25292
rect 968 25188 1032 25192
rect 968 25132 972 25188
rect 972 25132 1028 25188
rect 1028 25132 1032 25188
rect 968 25128 1032 25132
rect 968 25028 1032 25032
rect 968 24972 972 25028
rect 972 24972 1028 25028
rect 1028 24972 1032 25028
rect 968 24968 1032 24972
rect 968 24868 1032 24872
rect 968 24812 972 24868
rect 972 24812 1028 24868
rect 1028 24812 1032 24868
rect 968 24808 1032 24812
rect 968 24708 1032 24712
rect 968 24652 972 24708
rect 972 24652 1028 24708
rect 1028 24652 1032 24708
rect 968 24648 1032 24652
rect 968 24548 1032 24552
rect 968 24492 972 24548
rect 972 24492 1028 24548
rect 1028 24492 1032 24548
rect 968 24488 1032 24492
rect 968 24388 1032 24392
rect 968 24332 972 24388
rect 972 24332 1028 24388
rect 1028 24332 1032 24388
rect 968 24328 1032 24332
rect 968 24228 1032 24232
rect 968 24172 972 24228
rect 972 24172 1028 24228
rect 1028 24172 1032 24228
rect 968 24168 1032 24172
rect 968 24068 1032 24072
rect 968 24012 972 24068
rect 972 24012 1028 24068
rect 1028 24012 1032 24068
rect 968 24008 1032 24012
rect 968 23908 1032 23912
rect 968 23852 972 23908
rect 972 23852 1028 23908
rect 1028 23852 1032 23908
rect 968 23848 1032 23852
rect 968 23748 1032 23752
rect 968 23692 972 23748
rect 972 23692 1028 23748
rect 1028 23692 1032 23748
rect 968 23688 1032 23692
rect 968 23588 1032 23592
rect 968 23532 972 23588
rect 972 23532 1028 23588
rect 1028 23532 1032 23588
rect 968 23528 1032 23532
rect 968 23428 1032 23432
rect 968 23372 972 23428
rect 972 23372 1028 23428
rect 1028 23372 1032 23428
rect 968 23368 1032 23372
rect 968 23268 1032 23272
rect 968 23212 972 23268
rect 972 23212 1028 23268
rect 1028 23212 1032 23268
rect 968 23208 1032 23212
rect 968 23108 1032 23112
rect 968 23052 972 23108
rect 972 23052 1028 23108
rect 1028 23052 1032 23108
rect 968 23048 1032 23052
rect 968 22948 1032 22952
rect 968 22892 972 22948
rect 972 22892 1028 22948
rect 1028 22892 1032 22948
rect 968 22888 1032 22892
rect 968 22788 1032 22792
rect 968 22732 972 22788
rect 972 22732 1028 22788
rect 1028 22732 1032 22788
rect 968 22728 1032 22732
rect 968 22468 1032 22472
rect 968 22412 972 22468
rect 972 22412 1028 22468
rect 1028 22412 1032 22468
rect 968 22408 1032 22412
rect 968 22148 1032 22152
rect 968 22092 972 22148
rect 972 22092 1028 22148
rect 1028 22092 1032 22148
rect 968 22088 1032 22092
rect 968 21988 1032 21992
rect 968 21932 972 21988
rect 972 21932 1028 21988
rect 1028 21932 1032 21988
rect 968 21928 1032 21932
rect 968 21828 1032 21832
rect 968 21772 972 21828
rect 972 21772 1028 21828
rect 1028 21772 1032 21828
rect 968 21768 1032 21772
rect 968 21668 1032 21672
rect 968 21612 972 21668
rect 972 21612 1028 21668
rect 1028 21612 1032 21668
rect 968 21608 1032 21612
rect 968 21508 1032 21512
rect 968 21452 972 21508
rect 972 21452 1028 21508
rect 1028 21452 1032 21508
rect 968 21448 1032 21452
rect 968 21348 1032 21352
rect 968 21292 972 21348
rect 972 21292 1028 21348
rect 1028 21292 1032 21348
rect 968 21288 1032 21292
rect 968 21188 1032 21192
rect 968 21132 972 21188
rect 972 21132 1028 21188
rect 1028 21132 1032 21188
rect 968 21128 1032 21132
rect 968 21028 1032 21032
rect 968 20972 972 21028
rect 972 20972 1028 21028
rect 1028 20972 1032 21028
rect 968 20968 1032 20972
rect 968 20868 1032 20872
rect 968 20812 972 20868
rect 972 20812 1028 20868
rect 1028 20812 1032 20868
rect 968 20808 1032 20812
rect 968 20708 1032 20712
rect 968 20652 972 20708
rect 972 20652 1028 20708
rect 1028 20652 1032 20708
rect 968 20648 1032 20652
rect 968 20548 1032 20552
rect 968 20492 972 20548
rect 972 20492 1028 20548
rect 1028 20492 1032 20548
rect 968 20488 1032 20492
rect 968 20388 1032 20392
rect 968 20332 972 20388
rect 972 20332 1028 20388
rect 1028 20332 1032 20388
rect 968 20328 1032 20332
rect 968 20228 1032 20232
rect 968 20172 972 20228
rect 972 20172 1028 20228
rect 1028 20172 1032 20228
rect 968 20168 1032 20172
rect 968 20068 1032 20072
rect 968 20012 972 20068
rect 972 20012 1028 20068
rect 1028 20012 1032 20068
rect 968 20008 1032 20012
rect 968 19908 1032 19912
rect 968 19852 972 19908
rect 972 19852 1028 19908
rect 1028 19852 1032 19908
rect 968 19848 1032 19852
rect 968 19588 1032 19592
rect 968 19532 972 19588
rect 972 19532 1028 19588
rect 1028 19532 1032 19588
rect 968 19528 1032 19532
rect 968 19428 1032 19432
rect 968 19372 972 19428
rect 972 19372 1028 19428
rect 1028 19372 1032 19428
rect 968 19368 1032 19372
rect 968 19268 1032 19272
rect 968 19212 972 19268
rect 972 19212 1028 19268
rect 1028 19212 1032 19268
rect 968 19208 1032 19212
rect 968 19108 1032 19112
rect 968 19052 972 19108
rect 972 19052 1028 19108
rect 1028 19052 1032 19108
rect 968 19048 1032 19052
rect 968 18948 1032 18952
rect 968 18892 972 18948
rect 972 18892 1028 18948
rect 1028 18892 1032 18948
rect 968 18888 1032 18892
rect 968 18788 1032 18792
rect 968 18732 972 18788
rect 972 18732 1028 18788
rect 1028 18732 1032 18788
rect 968 18728 1032 18732
rect 968 18628 1032 18632
rect 968 18572 972 18628
rect 972 18572 1028 18628
rect 1028 18572 1032 18628
rect 968 18568 1032 18572
rect 968 18468 1032 18472
rect 968 18412 972 18468
rect 972 18412 1028 18468
rect 1028 18412 1032 18468
rect 968 18408 1032 18412
rect 968 18308 1032 18312
rect 968 18252 972 18308
rect 972 18252 1028 18308
rect 1028 18252 1032 18308
rect 968 18248 1032 18252
rect 968 18148 1032 18152
rect 968 18092 972 18148
rect 972 18092 1028 18148
rect 1028 18092 1032 18148
rect 968 18088 1032 18092
rect 968 17988 1032 17992
rect 968 17932 972 17988
rect 972 17932 1028 17988
rect 1028 17932 1032 17988
rect 968 17928 1032 17932
rect 968 17828 1032 17832
rect 968 17772 972 17828
rect 972 17772 1028 17828
rect 1028 17772 1032 17828
rect 968 17768 1032 17772
rect 968 17668 1032 17672
rect 968 17612 972 17668
rect 972 17612 1028 17668
rect 1028 17612 1032 17668
rect 968 17608 1032 17612
rect 968 17508 1032 17512
rect 968 17452 972 17508
rect 972 17452 1028 17508
rect 1028 17452 1032 17508
rect 968 17448 1032 17452
rect 968 17348 1032 17352
rect 968 17292 972 17348
rect 972 17292 1028 17348
rect 1028 17292 1032 17348
rect 968 17288 1032 17292
rect 968 17028 1032 17032
rect 968 16972 972 17028
rect 972 16972 1028 17028
rect 1028 16972 1032 17028
rect 968 16968 1032 16972
rect 968 16708 1032 16712
rect 968 16652 972 16708
rect 972 16652 1028 16708
rect 1028 16652 1032 16708
rect 968 16648 1032 16652
rect 968 16548 1032 16552
rect 968 16492 972 16548
rect 972 16492 1028 16548
rect 1028 16492 1032 16548
rect 968 16488 1032 16492
rect 968 16388 1032 16392
rect 968 16332 972 16388
rect 972 16332 1028 16388
rect 1028 16332 1032 16388
rect 968 16328 1032 16332
rect 968 16228 1032 16232
rect 968 16172 972 16228
rect 972 16172 1028 16228
rect 1028 16172 1032 16228
rect 968 16168 1032 16172
rect 968 15908 1032 15912
rect 968 15852 972 15908
rect 972 15852 1028 15908
rect 1028 15852 1032 15908
rect 968 15848 1032 15852
rect 968 15588 1032 15592
rect 968 15532 972 15588
rect 972 15532 1028 15588
rect 1028 15532 1032 15588
rect 968 15528 1032 15532
rect 968 15428 1032 15432
rect 968 15372 972 15428
rect 972 15372 1028 15428
rect 1028 15372 1032 15428
rect 968 15368 1032 15372
rect 968 15268 1032 15272
rect 968 15212 972 15268
rect 972 15212 1028 15268
rect 1028 15212 1032 15268
rect 968 15208 1032 15212
rect 968 15108 1032 15112
rect 968 15052 972 15108
rect 972 15052 1028 15108
rect 1028 15052 1032 15108
rect 968 15048 1032 15052
rect 968 14948 1032 14952
rect 968 14892 972 14948
rect 972 14892 1028 14948
rect 1028 14892 1032 14948
rect 968 14888 1032 14892
rect 968 14788 1032 14792
rect 968 14732 972 14788
rect 972 14732 1028 14788
rect 1028 14732 1032 14788
rect 968 14728 1032 14732
rect 968 14628 1032 14632
rect 968 14572 972 14628
rect 972 14572 1028 14628
rect 1028 14572 1032 14628
rect 968 14568 1032 14572
rect 968 14468 1032 14472
rect 968 14412 972 14468
rect 972 14412 1028 14468
rect 1028 14412 1032 14468
rect 968 14408 1032 14412
rect 968 14308 1032 14312
rect 968 14252 972 14308
rect 972 14252 1028 14308
rect 1028 14252 1032 14308
rect 968 14248 1032 14252
rect 968 14148 1032 14152
rect 968 14092 972 14148
rect 972 14092 1028 14148
rect 1028 14092 1032 14148
rect 968 14088 1032 14092
rect 968 13988 1032 13992
rect 968 13932 972 13988
rect 972 13932 1028 13988
rect 1028 13932 1032 13988
rect 968 13928 1032 13932
rect 968 13828 1032 13832
rect 968 13772 972 13828
rect 972 13772 1028 13828
rect 1028 13772 1032 13828
rect 968 13768 1032 13772
rect 968 13668 1032 13672
rect 968 13612 972 13668
rect 972 13612 1028 13668
rect 1028 13612 1032 13668
rect 968 13608 1032 13612
rect 968 13508 1032 13512
rect 968 13452 972 13508
rect 972 13452 1028 13508
rect 1028 13452 1032 13508
rect 968 13448 1032 13452
rect 968 13348 1032 13352
rect 968 13292 972 13348
rect 972 13292 1028 13348
rect 1028 13292 1032 13348
rect 968 13288 1032 13292
rect 968 13028 1032 13032
rect 968 12972 972 13028
rect 972 12972 1028 13028
rect 1028 12972 1032 13028
rect 968 12968 1032 12972
rect 968 12868 1032 12872
rect 968 12812 972 12868
rect 972 12812 1028 12868
rect 1028 12812 1032 12868
rect 968 12808 1032 12812
rect 968 12708 1032 12712
rect 968 12652 972 12708
rect 972 12652 1028 12708
rect 1028 12652 1032 12708
rect 968 12648 1032 12652
rect 968 12548 1032 12552
rect 968 12492 972 12548
rect 972 12492 1028 12548
rect 1028 12492 1032 12548
rect 968 12488 1032 12492
rect 968 12388 1032 12392
rect 968 12332 972 12388
rect 972 12332 1028 12388
rect 1028 12332 1032 12388
rect 968 12328 1032 12332
rect 968 12228 1032 12232
rect 968 12172 972 12228
rect 972 12172 1028 12228
rect 1028 12172 1032 12228
rect 968 12168 1032 12172
rect 968 12068 1032 12072
rect 968 12012 972 12068
rect 972 12012 1028 12068
rect 1028 12012 1032 12068
rect 968 12008 1032 12012
rect 968 11908 1032 11912
rect 968 11852 972 11908
rect 972 11852 1028 11908
rect 1028 11852 1032 11908
rect 968 11848 1032 11852
rect 968 11748 1032 11752
rect 968 11692 972 11748
rect 972 11692 1028 11748
rect 1028 11692 1032 11748
rect 968 11688 1032 11692
rect 968 11588 1032 11592
rect 968 11532 972 11588
rect 972 11532 1028 11588
rect 1028 11532 1032 11588
rect 968 11528 1032 11532
rect 968 11428 1032 11432
rect 968 11372 972 11428
rect 972 11372 1028 11428
rect 1028 11372 1032 11428
rect 968 11368 1032 11372
rect 968 11268 1032 11272
rect 968 11212 972 11268
rect 972 11212 1028 11268
rect 1028 11212 1032 11268
rect 968 11208 1032 11212
rect 968 11108 1032 11112
rect 968 11052 972 11108
rect 972 11052 1028 11108
rect 1028 11052 1032 11108
rect 968 11048 1032 11052
rect 968 10948 1032 10952
rect 968 10892 972 10948
rect 972 10892 1028 10948
rect 1028 10892 1032 10948
rect 968 10888 1032 10892
rect 968 10788 1032 10792
rect 968 10732 972 10788
rect 972 10732 1028 10788
rect 1028 10732 1032 10788
rect 968 10728 1032 10732
rect 968 10468 1032 10472
rect 968 10412 972 10468
rect 972 10412 1028 10468
rect 1028 10412 1032 10468
rect 968 10408 1032 10412
rect 968 10148 1032 10152
rect 968 10092 972 10148
rect 972 10092 1028 10148
rect 1028 10092 1032 10148
rect 968 10088 1032 10092
rect 968 9988 1032 9992
rect 968 9932 972 9988
rect 972 9932 1028 9988
rect 1028 9932 1032 9988
rect 968 9928 1032 9932
rect 968 9828 1032 9832
rect 968 9772 972 9828
rect 972 9772 1028 9828
rect 1028 9772 1032 9828
rect 968 9768 1032 9772
rect 968 9668 1032 9672
rect 968 9612 972 9668
rect 972 9612 1028 9668
rect 1028 9612 1032 9668
rect 968 9608 1032 9612
rect 968 9508 1032 9512
rect 968 9452 972 9508
rect 972 9452 1028 9508
rect 1028 9452 1032 9508
rect 968 9448 1032 9452
rect 968 9348 1032 9352
rect 968 9292 972 9348
rect 972 9292 1028 9348
rect 1028 9292 1032 9348
rect 968 9288 1032 9292
rect 968 9188 1032 9192
rect 968 9132 972 9188
rect 972 9132 1028 9188
rect 1028 9132 1032 9188
rect 968 9128 1032 9132
rect 968 9028 1032 9032
rect 968 8972 972 9028
rect 972 8972 1028 9028
rect 1028 8972 1032 9028
rect 968 8968 1032 8972
rect 968 8868 1032 8872
rect 968 8812 972 8868
rect 972 8812 1028 8868
rect 1028 8812 1032 8868
rect 968 8808 1032 8812
rect 968 8708 1032 8712
rect 968 8652 972 8708
rect 972 8652 1028 8708
rect 1028 8652 1032 8708
rect 968 8648 1032 8652
rect 968 8548 1032 8552
rect 968 8492 972 8548
rect 972 8492 1028 8548
rect 1028 8492 1032 8548
rect 968 8488 1032 8492
rect 968 8388 1032 8392
rect 968 8332 972 8388
rect 972 8332 1028 8388
rect 1028 8332 1032 8388
rect 968 8328 1032 8332
rect 968 8228 1032 8232
rect 968 8172 972 8228
rect 972 8172 1028 8228
rect 1028 8172 1032 8228
rect 968 8168 1032 8172
rect 968 8068 1032 8072
rect 968 8012 972 8068
rect 972 8012 1028 8068
rect 1028 8012 1032 8068
rect 968 8008 1032 8012
rect 968 7908 1032 7912
rect 968 7852 972 7908
rect 972 7852 1028 7908
rect 1028 7852 1032 7908
rect 968 7848 1032 7852
rect 968 7748 1032 7752
rect 968 7692 972 7748
rect 972 7692 1028 7748
rect 1028 7692 1032 7748
rect 968 7688 1032 7692
rect 968 7588 1032 7592
rect 968 7532 972 7588
rect 972 7532 1028 7588
rect 1028 7532 1032 7588
rect 968 7528 1032 7532
rect 968 7428 1032 7432
rect 968 7372 972 7428
rect 972 7372 1028 7428
rect 1028 7372 1032 7428
rect 968 7368 1032 7372
rect 968 7268 1032 7272
rect 968 7212 972 7268
rect 972 7212 1028 7268
rect 1028 7212 1032 7268
rect 968 7208 1032 7212
rect 968 7108 1032 7112
rect 968 7052 972 7108
rect 972 7052 1028 7108
rect 1028 7052 1032 7108
rect 968 7048 1032 7052
rect 968 6948 1032 6952
rect 968 6892 972 6948
rect 972 6892 1028 6948
rect 1028 6892 1032 6948
rect 968 6888 1032 6892
rect 968 6788 1032 6792
rect 968 6732 972 6788
rect 972 6732 1028 6788
rect 1028 6732 1032 6788
rect 968 6728 1032 6732
rect 968 6628 1032 6632
rect 968 6572 972 6628
rect 972 6572 1028 6628
rect 1028 6572 1032 6628
rect 968 6568 1032 6572
rect 968 6468 1032 6472
rect 968 6412 972 6468
rect 972 6412 1028 6468
rect 1028 6412 1032 6468
rect 968 6408 1032 6412
rect 968 6308 1032 6312
rect 968 6252 972 6308
rect 972 6252 1028 6308
rect 1028 6252 1032 6308
rect 968 6248 1032 6252
rect 968 6148 1032 6152
rect 968 6092 972 6148
rect 972 6092 1028 6148
rect 1028 6092 1032 6148
rect 968 6088 1032 6092
rect 968 5988 1032 5992
rect 968 5932 972 5988
rect 972 5932 1028 5988
rect 1028 5932 1032 5988
rect 968 5928 1032 5932
rect 968 5828 1032 5832
rect 968 5772 972 5828
rect 972 5772 1028 5828
rect 1028 5772 1032 5828
rect 968 5768 1032 5772
rect 968 5668 1032 5672
rect 968 5612 972 5668
rect 972 5612 1028 5668
rect 1028 5612 1032 5668
rect 968 5608 1032 5612
rect 968 5508 1032 5512
rect 968 5452 972 5508
rect 972 5452 1028 5508
rect 1028 5452 1032 5508
rect 968 5448 1032 5452
rect 968 5348 1032 5352
rect 968 5292 972 5348
rect 972 5292 1028 5348
rect 1028 5292 1032 5348
rect 968 5288 1032 5292
rect 968 5188 1032 5192
rect 968 5132 972 5188
rect 972 5132 1028 5188
rect 1028 5132 1032 5188
rect 968 5128 1032 5132
rect 968 5028 1032 5032
rect 968 4972 972 5028
rect 972 4972 1028 5028
rect 1028 4972 1032 5028
rect 968 4968 1032 4972
rect 968 4868 1032 4872
rect 968 4812 972 4868
rect 972 4812 1028 4868
rect 1028 4812 1032 4868
rect 968 4808 1032 4812
rect 968 4708 1032 4712
rect 968 4652 972 4708
rect 972 4652 1028 4708
rect 1028 4652 1032 4708
rect 968 4648 1032 4652
rect 968 4548 1032 4552
rect 968 4492 972 4548
rect 972 4492 1028 4548
rect 1028 4492 1032 4548
rect 968 4488 1032 4492
rect 968 4388 1032 4392
rect 968 4332 972 4388
rect 972 4332 1028 4388
rect 1028 4332 1032 4388
rect 968 4328 1032 4332
rect 968 4228 1032 4232
rect 968 4172 972 4228
rect 972 4172 1028 4228
rect 1028 4172 1032 4228
rect 968 4168 1032 4172
rect 968 4068 1032 4072
rect 968 4012 972 4068
rect 972 4012 1028 4068
rect 1028 4012 1032 4068
rect 968 4008 1032 4012
rect 968 3908 1032 3912
rect 968 3852 972 3908
rect 972 3852 1028 3908
rect 1028 3852 1032 3908
rect 968 3848 1032 3852
rect 968 3748 1032 3752
rect 968 3692 972 3748
rect 972 3692 1028 3748
rect 1028 3692 1032 3748
rect 968 3688 1032 3692
rect 968 3588 1032 3592
rect 968 3532 972 3588
rect 972 3532 1028 3588
rect 1028 3532 1032 3588
rect 968 3528 1032 3532
rect 968 3428 1032 3432
rect 968 3372 972 3428
rect 972 3372 1028 3428
rect 1028 3372 1032 3428
rect 968 3368 1032 3372
rect 968 3268 1032 3272
rect 968 3212 972 3268
rect 972 3212 1028 3268
rect 1028 3212 1032 3268
rect 968 3208 1032 3212
rect 968 3108 1032 3112
rect 968 3052 972 3108
rect 972 3052 1028 3108
rect 1028 3052 1032 3108
rect 968 3048 1032 3052
rect 968 2948 1032 2952
rect 968 2892 972 2948
rect 972 2892 1028 2948
rect 1028 2892 1032 2948
rect 968 2888 1032 2892
rect 968 2788 1032 2792
rect 968 2732 972 2788
rect 972 2732 1028 2788
rect 1028 2732 1032 2788
rect 968 2728 1032 2732
rect 968 2628 1032 2632
rect 968 2572 972 2628
rect 972 2572 1028 2628
rect 1028 2572 1032 2628
rect 968 2568 1032 2572
rect 968 2468 1032 2472
rect 968 2412 972 2468
rect 972 2412 1028 2468
rect 1028 2412 1032 2468
rect 968 2408 1032 2412
rect 968 2308 1032 2312
rect 968 2252 972 2308
rect 972 2252 1028 2308
rect 1028 2252 1032 2308
rect 968 2248 1032 2252
rect 968 2148 1032 2152
rect 968 2092 972 2148
rect 972 2092 1028 2148
rect 1028 2092 1032 2148
rect 968 2088 1032 2092
rect 968 1988 1032 1992
rect 968 1932 972 1988
rect 972 1932 1028 1988
rect 1028 1932 1032 1988
rect 968 1928 1032 1932
rect 968 1828 1032 1832
rect 968 1772 972 1828
rect 972 1772 1028 1828
rect 1028 1772 1032 1828
rect 968 1768 1032 1772
rect 968 1668 1032 1672
rect 968 1612 972 1668
rect 972 1612 1028 1668
rect 1028 1612 1032 1668
rect 968 1608 1032 1612
rect 968 1508 1032 1512
rect 968 1452 972 1508
rect 972 1452 1028 1508
rect 1028 1452 1032 1508
rect 968 1448 1032 1452
rect 968 1348 1032 1352
rect 968 1292 972 1348
rect 972 1292 1028 1348
rect 1028 1292 1032 1348
rect 968 1288 1032 1292
rect 968 1188 1032 1192
rect 968 1132 972 1188
rect 972 1132 1028 1188
rect 1028 1132 1032 1188
rect 968 1128 1032 1132
rect 28968 31908 29032 31912
rect 28968 31852 28972 31908
rect 28972 31852 29028 31908
rect 29028 31852 29032 31908
rect 28968 31848 29032 31852
rect 28968 31748 29032 31752
rect 28968 31692 28972 31748
rect 28972 31692 29028 31748
rect 29028 31692 29032 31748
rect 28968 31688 29032 31692
rect 28968 31588 29032 31592
rect 28968 31532 28972 31588
rect 28972 31532 29028 31588
rect 29028 31532 29032 31588
rect 28968 31528 29032 31532
rect 28968 31428 29032 31432
rect 28968 31372 28972 31428
rect 28972 31372 29028 31428
rect 29028 31372 29032 31428
rect 28968 31368 29032 31372
rect 28968 31268 29032 31272
rect 28968 31212 28972 31268
rect 28972 31212 29028 31268
rect 29028 31212 29032 31268
rect 28968 31208 29032 31212
rect 28968 31108 29032 31112
rect 28968 31052 28972 31108
rect 28972 31052 29028 31108
rect 29028 31052 29032 31108
rect 28968 31048 29032 31052
rect 28968 30948 29032 30952
rect 28968 30892 28972 30948
rect 28972 30892 29028 30948
rect 29028 30892 29032 30948
rect 28968 30888 29032 30892
rect 28968 30788 29032 30792
rect 28968 30732 28972 30788
rect 28972 30732 29028 30788
rect 29028 30732 29032 30788
rect 28968 30728 29032 30732
rect 28968 30628 29032 30632
rect 28968 30572 28972 30628
rect 28972 30572 29028 30628
rect 29028 30572 29032 30628
rect 28968 30568 29032 30572
rect 28968 30468 29032 30472
rect 28968 30412 28972 30468
rect 28972 30412 29028 30468
rect 29028 30412 29032 30468
rect 28968 30408 29032 30412
rect 28968 30308 29032 30312
rect 28968 30252 28972 30308
rect 28972 30252 29028 30308
rect 29028 30252 29032 30308
rect 28968 30248 29032 30252
rect 28968 30148 29032 30152
rect 28968 30092 28972 30148
rect 28972 30092 29028 30148
rect 29028 30092 29032 30148
rect 28968 30088 29032 30092
rect 28968 29988 29032 29992
rect 28968 29932 28972 29988
rect 28972 29932 29028 29988
rect 29028 29932 29032 29988
rect 28968 29928 29032 29932
rect 28968 29828 29032 29832
rect 28968 29772 28972 29828
rect 28972 29772 29028 29828
rect 29028 29772 29032 29828
rect 28968 29768 29032 29772
rect 28968 29668 29032 29672
rect 28968 29612 28972 29668
rect 28972 29612 29028 29668
rect 29028 29612 29032 29668
rect 28968 29608 29032 29612
rect 28968 29508 29032 29512
rect 28968 29452 28972 29508
rect 28972 29452 29028 29508
rect 29028 29452 29032 29508
rect 28968 29448 29032 29452
rect 28968 29348 29032 29352
rect 28968 29292 28972 29348
rect 28972 29292 29028 29348
rect 29028 29292 29032 29348
rect 28968 29288 29032 29292
rect 28968 29028 29032 29032
rect 28968 28972 28972 29028
rect 28972 28972 29028 29028
rect 29028 28972 29032 29028
rect 28968 28968 29032 28972
rect 28968 28708 29032 28712
rect 28968 28652 28972 28708
rect 28972 28652 29028 28708
rect 29028 28652 29032 28708
rect 28968 28648 29032 28652
rect 28968 28548 29032 28552
rect 28968 28492 28972 28548
rect 28972 28492 29028 28548
rect 29028 28492 29032 28548
rect 28968 28488 29032 28492
rect 28968 28388 29032 28392
rect 28968 28332 28972 28388
rect 28972 28332 29028 28388
rect 29028 28332 29032 28388
rect 28968 28328 29032 28332
rect 28968 28228 29032 28232
rect 28968 28172 28972 28228
rect 28972 28172 29028 28228
rect 29028 28172 29032 28228
rect 28968 28168 29032 28172
rect 28968 28068 29032 28072
rect 28968 28012 28972 28068
rect 28972 28012 29028 28068
rect 29028 28012 29032 28068
rect 28968 28008 29032 28012
rect 28968 27908 29032 27912
rect 28968 27852 28972 27908
rect 28972 27852 29028 27908
rect 29028 27852 29032 27908
rect 28968 27848 29032 27852
rect 28968 27748 29032 27752
rect 28968 27692 28972 27748
rect 28972 27692 29028 27748
rect 29028 27692 29032 27748
rect 28968 27688 29032 27692
rect 28968 27588 29032 27592
rect 28968 27532 28972 27588
rect 28972 27532 29028 27588
rect 29028 27532 29032 27588
rect 28968 27528 29032 27532
rect 28968 27428 29032 27432
rect 28968 27372 28972 27428
rect 28972 27372 29028 27428
rect 29028 27372 29032 27428
rect 28968 27368 29032 27372
rect 28968 27268 29032 27272
rect 28968 27212 28972 27268
rect 28972 27212 29028 27268
rect 29028 27212 29032 27268
rect 28968 27208 29032 27212
rect 28968 27108 29032 27112
rect 28968 27052 28972 27108
rect 28972 27052 29028 27108
rect 29028 27052 29032 27108
rect 28968 27048 29032 27052
rect 28968 26948 29032 26952
rect 28968 26892 28972 26948
rect 28972 26892 29028 26948
rect 29028 26892 29032 26948
rect 28968 26888 29032 26892
rect 28968 26788 29032 26792
rect 28968 26732 28972 26788
rect 28972 26732 29028 26788
rect 29028 26732 29032 26788
rect 28968 26728 29032 26732
rect 28968 26628 29032 26632
rect 28968 26572 28972 26628
rect 28972 26572 29028 26628
rect 29028 26572 29032 26628
rect 28968 26568 29032 26572
rect 28968 26468 29032 26472
rect 28968 26412 28972 26468
rect 28972 26412 29028 26468
rect 29028 26412 29032 26468
rect 28968 26408 29032 26412
rect 28968 26148 29032 26152
rect 28968 26092 28972 26148
rect 28972 26092 29028 26148
rect 29028 26092 29032 26148
rect 28968 26088 29032 26092
rect 28968 25988 29032 25992
rect 28968 25932 28972 25988
rect 28972 25932 29028 25988
rect 29028 25932 29032 25988
rect 28968 25928 29032 25932
rect 28968 25828 29032 25832
rect 28968 25772 28972 25828
rect 28972 25772 29028 25828
rect 29028 25772 29032 25828
rect 28968 25768 29032 25772
rect 28968 25668 29032 25672
rect 28968 25612 28972 25668
rect 28972 25612 29028 25668
rect 29028 25612 29032 25668
rect 28968 25608 29032 25612
rect 28968 25508 29032 25512
rect 28968 25452 28972 25508
rect 28972 25452 29028 25508
rect 29028 25452 29032 25508
rect 28968 25448 29032 25452
rect 28968 25348 29032 25352
rect 28968 25292 28972 25348
rect 28972 25292 29028 25348
rect 29028 25292 29032 25348
rect 28968 25288 29032 25292
rect 28968 25188 29032 25192
rect 28968 25132 28972 25188
rect 28972 25132 29028 25188
rect 29028 25132 29032 25188
rect 28968 25128 29032 25132
rect 28968 25028 29032 25032
rect 28968 24972 28972 25028
rect 28972 24972 29028 25028
rect 29028 24972 29032 25028
rect 28968 24968 29032 24972
rect 28968 24868 29032 24872
rect 28968 24812 28972 24868
rect 28972 24812 29028 24868
rect 29028 24812 29032 24868
rect 28968 24808 29032 24812
rect 28968 24708 29032 24712
rect 28968 24652 28972 24708
rect 28972 24652 29028 24708
rect 29028 24652 29032 24708
rect 28968 24648 29032 24652
rect 28968 24548 29032 24552
rect 28968 24492 28972 24548
rect 28972 24492 29028 24548
rect 29028 24492 29032 24548
rect 28968 24488 29032 24492
rect 28968 24388 29032 24392
rect 28968 24332 28972 24388
rect 28972 24332 29028 24388
rect 29028 24332 29032 24388
rect 28968 24328 29032 24332
rect 28968 24228 29032 24232
rect 28968 24172 28972 24228
rect 28972 24172 29028 24228
rect 29028 24172 29032 24228
rect 28968 24168 29032 24172
rect 28968 24068 29032 24072
rect 28968 24012 28972 24068
rect 28972 24012 29028 24068
rect 29028 24012 29032 24068
rect 28968 24008 29032 24012
rect 28968 23908 29032 23912
rect 28968 23852 28972 23908
rect 28972 23852 29028 23908
rect 29028 23852 29032 23908
rect 28968 23848 29032 23852
rect 28968 23588 29032 23592
rect 28968 23532 28972 23588
rect 28972 23532 29028 23588
rect 29028 23532 29032 23588
rect 28968 23528 29032 23532
rect 28968 23268 29032 23272
rect 28968 23212 28972 23268
rect 28972 23212 29028 23268
rect 29028 23212 29032 23268
rect 28968 23208 29032 23212
rect 28968 23108 29032 23112
rect 28968 23052 28972 23108
rect 28972 23052 29028 23108
rect 29028 23052 29032 23108
rect 28968 23048 29032 23052
rect 28968 22948 29032 22952
rect 28968 22892 28972 22948
rect 28972 22892 29028 22948
rect 29028 22892 29032 22948
rect 28968 22888 29032 22892
rect 28968 22788 29032 22792
rect 28968 22732 28972 22788
rect 28972 22732 29028 22788
rect 29028 22732 29032 22788
rect 28968 22728 29032 22732
rect 28968 22628 29032 22632
rect 28968 22572 28972 22628
rect 28972 22572 29028 22628
rect 29028 22572 29032 22628
rect 28968 22568 29032 22572
rect 28968 22468 29032 22472
rect 28968 22412 28972 22468
rect 28972 22412 29028 22468
rect 29028 22412 29032 22468
rect 28968 22408 29032 22412
rect 28968 22308 29032 22312
rect 28968 22252 28972 22308
rect 28972 22252 29028 22308
rect 29028 22252 29032 22308
rect 28968 22248 29032 22252
rect 28968 22148 29032 22152
rect 28968 22092 28972 22148
rect 28972 22092 29028 22148
rect 29028 22092 29032 22148
rect 28968 22088 29032 22092
rect 28968 21988 29032 21992
rect 28968 21932 28972 21988
rect 28972 21932 29028 21988
rect 29028 21932 29032 21988
rect 28968 21928 29032 21932
rect 28968 21828 29032 21832
rect 28968 21772 28972 21828
rect 28972 21772 29028 21828
rect 29028 21772 29032 21828
rect 28968 21768 29032 21772
rect 28968 21668 29032 21672
rect 28968 21612 28972 21668
rect 28972 21612 29028 21668
rect 29028 21612 29032 21668
rect 28968 21608 29032 21612
rect 28968 21508 29032 21512
rect 28968 21452 28972 21508
rect 28972 21452 29028 21508
rect 29028 21452 29032 21508
rect 28968 21448 29032 21452
rect 28968 21348 29032 21352
rect 28968 21292 28972 21348
rect 28972 21292 29028 21348
rect 29028 21292 29032 21348
rect 28968 21288 29032 21292
rect 28968 21188 29032 21192
rect 28968 21132 28972 21188
rect 28972 21132 29028 21188
rect 29028 21132 29032 21188
rect 28968 21128 29032 21132
rect 28968 21028 29032 21032
rect 28968 20972 28972 21028
rect 28972 20972 29028 21028
rect 29028 20972 29032 21028
rect 28968 20968 29032 20972
rect 28968 20868 29032 20872
rect 28968 20812 28972 20868
rect 28972 20812 29028 20868
rect 29028 20812 29032 20868
rect 28968 20808 29032 20812
rect 28968 20708 29032 20712
rect 28968 20652 28972 20708
rect 28972 20652 29028 20708
rect 29028 20652 29032 20708
rect 28968 20648 29032 20652
rect 28968 20548 29032 20552
rect 28968 20492 28972 20548
rect 28972 20492 29028 20548
rect 29028 20492 29032 20548
rect 28968 20488 29032 20492
rect 28968 20388 29032 20392
rect 28968 20332 28972 20388
rect 28972 20332 29028 20388
rect 29028 20332 29032 20388
rect 28968 20328 29032 20332
rect 28968 20228 29032 20232
rect 28968 20172 28972 20228
rect 28972 20172 29028 20228
rect 29028 20172 29032 20228
rect 28968 20168 29032 20172
rect 28968 20068 29032 20072
rect 28968 20012 28972 20068
rect 28972 20012 29028 20068
rect 29028 20012 29032 20068
rect 28968 20008 29032 20012
rect 28968 19908 29032 19912
rect 28968 19852 28972 19908
rect 28972 19852 29028 19908
rect 29028 19852 29032 19908
rect 28968 19848 29032 19852
rect 28968 19748 29032 19752
rect 28968 19692 28972 19748
rect 28972 19692 29028 19748
rect 29028 19692 29032 19748
rect 28968 19688 29032 19692
rect 28968 19588 29032 19592
rect 28968 19532 28972 19588
rect 28972 19532 29028 19588
rect 29028 19532 29032 19588
rect 28968 19528 29032 19532
rect 28968 19428 29032 19432
rect 28968 19372 28972 19428
rect 28972 19372 29028 19428
rect 29028 19372 29032 19428
rect 28968 19368 29032 19372
rect 28968 19268 29032 19272
rect 28968 19212 28972 19268
rect 28972 19212 29028 19268
rect 29028 19212 29032 19268
rect 28968 19208 29032 19212
rect 28968 19108 29032 19112
rect 28968 19052 28972 19108
rect 28972 19052 29028 19108
rect 29028 19052 29032 19108
rect 28968 19048 29032 19052
rect 28968 18948 29032 18952
rect 28968 18892 28972 18948
rect 28972 18892 29028 18948
rect 29028 18892 29032 18948
rect 28968 18888 29032 18892
rect 28968 18788 29032 18792
rect 28968 18732 28972 18788
rect 28972 18732 29028 18788
rect 29028 18732 29032 18788
rect 28968 18728 29032 18732
rect 28968 18628 29032 18632
rect 28968 18572 28972 18628
rect 28972 18572 29028 18628
rect 29028 18572 29032 18628
rect 28968 18568 29032 18572
rect 28968 18468 29032 18472
rect 28968 18412 28972 18468
rect 28972 18412 29028 18468
rect 29028 18412 29032 18468
rect 28968 18408 29032 18412
rect 28968 18308 29032 18312
rect 28968 18252 28972 18308
rect 28972 18252 29028 18308
rect 29028 18252 29032 18308
rect 28968 18248 29032 18252
rect 28968 18148 29032 18152
rect 28968 18092 28972 18148
rect 28972 18092 29028 18148
rect 29028 18092 29032 18148
rect 28968 18088 29032 18092
rect 28968 17988 29032 17992
rect 28968 17932 28972 17988
rect 28972 17932 29028 17988
rect 29028 17932 29032 17988
rect 28968 17928 29032 17932
rect 28968 17828 29032 17832
rect 28968 17772 28972 17828
rect 28972 17772 29028 17828
rect 29028 17772 29032 17828
rect 28968 17768 29032 17772
rect 28968 17668 29032 17672
rect 28968 17612 28972 17668
rect 28972 17612 29028 17668
rect 29028 17612 29032 17668
rect 28968 17608 29032 17612
rect 28968 17508 29032 17512
rect 28968 17452 28972 17508
rect 28972 17452 29028 17508
rect 29028 17452 29032 17508
rect 28968 17448 29032 17452
rect 28968 17348 29032 17352
rect 28968 17292 28972 17348
rect 28972 17292 29028 17348
rect 29028 17292 29032 17348
rect 28968 17288 29032 17292
rect 28968 17188 29032 17192
rect 28968 17132 28972 17188
rect 28972 17132 29028 17188
rect 29028 17132 29032 17188
rect 28968 17128 29032 17132
rect 28968 17028 29032 17032
rect 28968 16972 28972 17028
rect 28972 16972 29028 17028
rect 29028 16972 29032 17028
rect 28968 16968 29032 16972
rect 28968 16868 29032 16872
rect 28968 16812 28972 16868
rect 28972 16812 29028 16868
rect 29028 16812 29032 16868
rect 28968 16808 29032 16812
rect 28968 16708 29032 16712
rect 28968 16652 28972 16708
rect 28972 16652 29028 16708
rect 29028 16652 29032 16708
rect 28968 16648 29032 16652
rect 28968 16548 29032 16552
rect 28968 16492 28972 16548
rect 28972 16492 29028 16548
rect 29028 16492 29032 16548
rect 28968 16488 29032 16492
rect 28968 16388 29032 16392
rect 28968 16332 28972 16388
rect 28972 16332 29028 16388
rect 29028 16332 29032 16388
rect 28968 16328 29032 16332
rect 28968 16228 29032 16232
rect 28968 16172 28972 16228
rect 28972 16172 29028 16228
rect 29028 16172 29032 16228
rect 28968 16168 29032 16172
rect 28968 16068 29032 16072
rect 28968 16012 28972 16068
rect 28972 16012 29028 16068
rect 29028 16012 29032 16068
rect 28968 16008 29032 16012
rect 28968 15908 29032 15912
rect 28968 15852 28972 15908
rect 28972 15852 29028 15908
rect 29028 15852 29032 15908
rect 28968 15848 29032 15852
rect 28968 15748 29032 15752
rect 28968 15692 28972 15748
rect 28972 15692 29028 15748
rect 29028 15692 29032 15748
rect 28968 15688 29032 15692
rect 28968 15588 29032 15592
rect 28968 15532 28972 15588
rect 28972 15532 29028 15588
rect 29028 15532 29032 15588
rect 28968 15528 29032 15532
rect 28968 15428 29032 15432
rect 28968 15372 28972 15428
rect 28972 15372 29028 15428
rect 29028 15372 29032 15428
rect 28968 15368 29032 15372
rect 28968 15268 29032 15272
rect 28968 15212 28972 15268
rect 28972 15212 29028 15268
rect 29028 15212 29032 15268
rect 28968 15208 29032 15212
rect 28968 15108 29032 15112
rect 28968 15052 28972 15108
rect 28972 15052 29028 15108
rect 29028 15052 29032 15108
rect 28968 15048 29032 15052
rect 28968 14948 29032 14952
rect 28968 14892 28972 14948
rect 28972 14892 29028 14948
rect 29028 14892 29032 14948
rect 28968 14888 29032 14892
rect 28968 14788 29032 14792
rect 28968 14732 28972 14788
rect 28972 14732 29028 14788
rect 29028 14732 29032 14788
rect 28968 14728 29032 14732
rect 28968 14628 29032 14632
rect 28968 14572 28972 14628
rect 28972 14572 29028 14628
rect 29028 14572 29032 14628
rect 28968 14568 29032 14572
rect 28968 14468 29032 14472
rect 28968 14412 28972 14468
rect 28972 14412 29028 14468
rect 29028 14412 29032 14468
rect 28968 14408 29032 14412
rect 28968 14308 29032 14312
rect 28968 14252 28972 14308
rect 28972 14252 29028 14308
rect 29028 14252 29032 14308
rect 28968 14248 29032 14252
rect 28968 14148 29032 14152
rect 28968 14092 28972 14148
rect 28972 14092 29028 14148
rect 29028 14092 29032 14148
rect 28968 14088 29032 14092
rect 28968 13988 29032 13992
rect 28968 13932 28972 13988
rect 28972 13932 29028 13988
rect 29028 13932 29032 13988
rect 28968 13928 29032 13932
rect 28968 13828 29032 13832
rect 28968 13772 28972 13828
rect 28972 13772 29028 13828
rect 29028 13772 29032 13828
rect 28968 13768 29032 13772
rect 28968 13668 29032 13672
rect 28968 13612 28972 13668
rect 28972 13612 29028 13668
rect 29028 13612 29032 13668
rect 28968 13608 29032 13612
rect 28968 13508 29032 13512
rect 28968 13452 28972 13508
rect 28972 13452 29028 13508
rect 29028 13452 29032 13508
rect 28968 13448 29032 13452
rect 28968 13348 29032 13352
rect 28968 13292 28972 13348
rect 28972 13292 29028 13348
rect 29028 13292 29032 13348
rect 28968 13288 29032 13292
rect 28968 13188 29032 13192
rect 28968 13132 28972 13188
rect 28972 13132 29028 13188
rect 29028 13132 29032 13188
rect 28968 13128 29032 13132
rect 28968 13028 29032 13032
rect 28968 12972 28972 13028
rect 28972 12972 29028 13028
rect 29028 12972 29032 13028
rect 28968 12968 29032 12972
rect 28968 12868 29032 12872
rect 28968 12812 28972 12868
rect 28972 12812 29028 12868
rect 29028 12812 29032 12868
rect 28968 12808 29032 12812
rect 28968 12708 29032 12712
rect 28968 12652 28972 12708
rect 28972 12652 29028 12708
rect 29028 12652 29032 12708
rect 28968 12648 29032 12652
rect 28968 12548 29032 12552
rect 28968 12492 28972 12548
rect 28972 12492 29028 12548
rect 29028 12492 29032 12548
rect 28968 12488 29032 12492
rect 28968 12388 29032 12392
rect 28968 12332 28972 12388
rect 28972 12332 29028 12388
rect 29028 12332 29032 12388
rect 28968 12328 29032 12332
rect 28968 12228 29032 12232
rect 28968 12172 28972 12228
rect 28972 12172 29028 12228
rect 29028 12172 29032 12228
rect 28968 12168 29032 12172
rect 28968 12068 29032 12072
rect 28968 12012 28972 12068
rect 28972 12012 29028 12068
rect 29028 12012 29032 12068
rect 28968 12008 29032 12012
rect 28968 11908 29032 11912
rect 28968 11852 28972 11908
rect 28972 11852 29028 11908
rect 29028 11852 29032 11908
rect 28968 11848 29032 11852
rect 28968 11748 29032 11752
rect 28968 11692 28972 11748
rect 28972 11692 29028 11748
rect 29028 11692 29032 11748
rect 28968 11688 29032 11692
rect 28968 11588 29032 11592
rect 28968 11532 28972 11588
rect 28972 11532 29028 11588
rect 29028 11532 29032 11588
rect 28968 11528 29032 11532
rect 28968 11428 29032 11432
rect 28968 11372 28972 11428
rect 28972 11372 29028 11428
rect 29028 11372 29032 11428
rect 28968 11368 29032 11372
rect 28968 11268 29032 11272
rect 28968 11212 28972 11268
rect 28972 11212 29028 11268
rect 29028 11212 29032 11268
rect 28968 11208 29032 11212
rect 28968 11108 29032 11112
rect 28968 11052 28972 11108
rect 28972 11052 29028 11108
rect 29028 11052 29032 11108
rect 28968 11048 29032 11052
rect 28968 10948 29032 10952
rect 28968 10892 28972 10948
rect 28972 10892 29028 10948
rect 29028 10892 29032 10948
rect 28968 10888 29032 10892
rect 28968 10788 29032 10792
rect 28968 10732 28972 10788
rect 28972 10732 29028 10788
rect 29028 10732 29032 10788
rect 28968 10728 29032 10732
rect 28968 10628 29032 10632
rect 28968 10572 28972 10628
rect 28972 10572 29028 10628
rect 29028 10572 29032 10628
rect 28968 10568 29032 10572
rect 28968 10468 29032 10472
rect 28968 10412 28972 10468
rect 28972 10412 29028 10468
rect 29028 10412 29032 10468
rect 28968 10408 29032 10412
rect 28968 10308 29032 10312
rect 28968 10252 28972 10308
rect 28972 10252 29028 10308
rect 29028 10252 29032 10308
rect 28968 10248 29032 10252
rect 28968 10148 29032 10152
rect 28968 10092 28972 10148
rect 28972 10092 29028 10148
rect 29028 10092 29032 10148
rect 28968 10088 29032 10092
rect 28968 9988 29032 9992
rect 28968 9932 28972 9988
rect 28972 9932 29028 9988
rect 29028 9932 29032 9988
rect 28968 9928 29032 9932
rect 28968 9828 29032 9832
rect 28968 9772 28972 9828
rect 28972 9772 29028 9828
rect 29028 9772 29032 9828
rect 28968 9768 29032 9772
rect 28968 9668 29032 9672
rect 28968 9612 28972 9668
rect 28972 9612 29028 9668
rect 29028 9612 29032 9668
rect 28968 9608 29032 9612
rect 28968 9348 29032 9352
rect 28968 9292 28972 9348
rect 28972 9292 29028 9348
rect 29028 9292 29032 9348
rect 28968 9288 29032 9292
rect 28968 9028 29032 9032
rect 28968 8972 28972 9028
rect 28972 8972 29028 9028
rect 29028 8972 29032 9028
rect 28968 8968 29032 8972
rect 28968 8868 29032 8872
rect 28968 8812 28972 8868
rect 28972 8812 29028 8868
rect 29028 8812 29032 8868
rect 28968 8808 29032 8812
rect 28968 8708 29032 8712
rect 28968 8652 28972 8708
rect 28972 8652 29028 8708
rect 29028 8652 29032 8708
rect 28968 8648 29032 8652
rect 28968 8548 29032 8552
rect 28968 8492 28972 8548
rect 28972 8492 29028 8548
rect 29028 8492 29032 8548
rect 28968 8488 29032 8492
rect 28968 8388 29032 8392
rect 28968 8332 28972 8388
rect 28972 8332 29028 8388
rect 29028 8332 29032 8388
rect 28968 8328 29032 8332
rect 28968 8228 29032 8232
rect 28968 8172 28972 8228
rect 28972 8172 29028 8228
rect 29028 8172 29032 8228
rect 28968 8168 29032 8172
rect 28968 8068 29032 8072
rect 28968 8012 28972 8068
rect 28972 8012 29028 8068
rect 29028 8012 29032 8068
rect 28968 8008 29032 8012
rect 28968 7908 29032 7912
rect 28968 7852 28972 7908
rect 28972 7852 29028 7908
rect 29028 7852 29032 7908
rect 28968 7848 29032 7852
rect 28968 7748 29032 7752
rect 28968 7692 28972 7748
rect 28972 7692 29028 7748
rect 29028 7692 29032 7748
rect 28968 7688 29032 7692
rect 28968 7588 29032 7592
rect 28968 7532 28972 7588
rect 28972 7532 29028 7588
rect 29028 7532 29032 7588
rect 28968 7528 29032 7532
rect 28968 7428 29032 7432
rect 28968 7372 28972 7428
rect 28972 7372 29028 7428
rect 29028 7372 29032 7428
rect 28968 7368 29032 7372
rect 28968 7268 29032 7272
rect 28968 7212 28972 7268
rect 28972 7212 29028 7268
rect 29028 7212 29032 7268
rect 28968 7208 29032 7212
rect 28968 7108 29032 7112
rect 28968 7052 28972 7108
rect 28972 7052 29028 7108
rect 29028 7052 29032 7108
rect 28968 7048 29032 7052
rect 28968 6948 29032 6952
rect 28968 6892 28972 6948
rect 28972 6892 29028 6948
rect 29028 6892 29032 6948
rect 28968 6888 29032 6892
rect 28968 6788 29032 6792
rect 28968 6732 28972 6788
rect 28972 6732 29028 6788
rect 29028 6732 29032 6788
rect 28968 6728 29032 6732
rect 28968 6468 29032 6472
rect 28968 6412 28972 6468
rect 28972 6412 29028 6468
rect 29028 6412 29032 6468
rect 28968 6408 29032 6412
rect 28968 6308 29032 6312
rect 28968 6252 28972 6308
rect 28972 6252 29028 6308
rect 29028 6252 29032 6308
rect 28968 6248 29032 6252
rect 28968 6148 29032 6152
rect 28968 6092 28972 6148
rect 28972 6092 29028 6148
rect 29028 6092 29032 6148
rect 28968 6088 29032 6092
rect 28968 5988 29032 5992
rect 28968 5932 28972 5988
rect 28972 5932 29028 5988
rect 29028 5932 29032 5988
rect 28968 5928 29032 5932
rect 28968 5828 29032 5832
rect 28968 5772 28972 5828
rect 28972 5772 29028 5828
rect 29028 5772 29032 5828
rect 28968 5768 29032 5772
rect 28968 5668 29032 5672
rect 28968 5612 28972 5668
rect 28972 5612 29028 5668
rect 29028 5612 29032 5668
rect 28968 5608 29032 5612
rect 28968 5508 29032 5512
rect 28968 5452 28972 5508
rect 28972 5452 29028 5508
rect 29028 5452 29032 5508
rect 28968 5448 29032 5452
rect 28968 5348 29032 5352
rect 28968 5292 28972 5348
rect 28972 5292 29028 5348
rect 29028 5292 29032 5348
rect 28968 5288 29032 5292
rect 28968 5188 29032 5192
rect 28968 5132 28972 5188
rect 28972 5132 29028 5188
rect 29028 5132 29032 5188
rect 28968 5128 29032 5132
rect 28968 5028 29032 5032
rect 28968 4972 28972 5028
rect 28972 4972 29028 5028
rect 29028 4972 29032 5028
rect 28968 4968 29032 4972
rect 28968 4868 29032 4872
rect 28968 4812 28972 4868
rect 28972 4812 29028 4868
rect 29028 4812 29032 4868
rect 28968 4808 29032 4812
rect 28968 4708 29032 4712
rect 28968 4652 28972 4708
rect 28972 4652 29028 4708
rect 29028 4652 29032 4708
rect 28968 4648 29032 4652
rect 28968 4548 29032 4552
rect 28968 4492 28972 4548
rect 28972 4492 29028 4548
rect 29028 4492 29032 4548
rect 28968 4488 29032 4492
rect 28968 4388 29032 4392
rect 28968 4332 28972 4388
rect 28972 4332 29028 4388
rect 29028 4332 29032 4388
rect 28968 4328 29032 4332
rect 28968 4228 29032 4232
rect 28968 4172 28972 4228
rect 28972 4172 29028 4228
rect 29028 4172 29032 4228
rect 28968 4168 29032 4172
rect 28968 3908 29032 3912
rect 28968 3852 28972 3908
rect 28972 3852 29028 3908
rect 29028 3852 29032 3908
rect 28968 3848 29032 3852
rect 28968 3588 29032 3592
rect 28968 3532 28972 3588
rect 28972 3532 29028 3588
rect 29028 3532 29032 3588
rect 28968 3528 29032 3532
rect 28968 3428 29032 3432
rect 28968 3372 28972 3428
rect 28972 3372 29028 3428
rect 29028 3372 29032 3428
rect 28968 3368 29032 3372
rect 28968 3268 29032 3272
rect 28968 3212 28972 3268
rect 28972 3212 29028 3268
rect 29028 3212 29032 3268
rect 28968 3208 29032 3212
rect 28968 3108 29032 3112
rect 28968 3052 28972 3108
rect 28972 3052 29028 3108
rect 29028 3052 29032 3108
rect 28968 3048 29032 3052
rect 28968 2948 29032 2952
rect 28968 2892 28972 2948
rect 28972 2892 29028 2948
rect 29028 2892 29032 2948
rect 28968 2888 29032 2892
rect 28968 2788 29032 2792
rect 28968 2732 28972 2788
rect 28972 2732 29028 2788
rect 29028 2732 29032 2788
rect 28968 2728 29032 2732
rect 28968 2628 29032 2632
rect 28968 2572 28972 2628
rect 28972 2572 29028 2628
rect 29028 2572 29032 2628
rect 28968 2568 29032 2572
rect 28968 2468 29032 2472
rect 28968 2412 28972 2468
rect 28972 2412 29028 2468
rect 29028 2412 29032 2468
rect 28968 2408 29032 2412
rect 28968 2308 29032 2312
rect 28968 2252 28972 2308
rect 28972 2252 29028 2308
rect 29028 2252 29032 2308
rect 28968 2248 29032 2252
rect 28968 2148 29032 2152
rect 28968 2092 28972 2148
rect 28972 2092 29028 2148
rect 29028 2092 29032 2148
rect 28968 2088 29032 2092
rect 28968 1988 29032 1992
rect 28968 1932 28972 1988
rect 28972 1932 29028 1988
rect 29028 1932 29032 1988
rect 28968 1928 29032 1932
rect 28968 1828 29032 1832
rect 28968 1772 28972 1828
rect 28972 1772 29028 1828
rect 29028 1772 29032 1828
rect 28968 1768 29032 1772
rect 28968 1668 29032 1672
rect 28968 1612 28972 1668
rect 28972 1612 29028 1668
rect 29028 1612 29032 1668
rect 28968 1608 29032 1612
rect 28968 1508 29032 1512
rect 28968 1452 28972 1508
rect 28972 1452 29028 1508
rect 29028 1452 29032 1508
rect 28968 1448 29032 1452
rect 28968 1348 29032 1352
rect 28968 1292 28972 1348
rect 28972 1292 29028 1348
rect 29028 1292 29032 1348
rect 28968 1288 29032 1292
rect 28968 1188 29032 1192
rect 28968 1132 28972 1188
rect 28972 1132 29028 1188
rect 29028 1132 29032 1188
rect 28968 1128 29032 1132
rect 968 1028 1032 1032
rect 968 972 972 1028
rect 972 972 1028 1028
rect 1028 972 1032 1028
rect 968 968 1032 972
rect 648 808 712 872
rect 648 728 712 792
rect 648 648 712 712
rect 648 568 712 632
rect 648 488 712 552
rect 968 808 1032 872
rect 968 728 1032 792
rect 968 648 1032 712
rect 968 568 1032 632
rect 968 488 1032 552
rect 1128 328 1192 392
rect 1128 248 1192 312
rect 1128 168 1192 232
rect 1128 88 1192 152
rect 1128 8 1192 72
rect 28968 1028 29032 1032
rect 28968 972 28972 1028
rect 28972 972 29028 1028
rect 29028 972 29032 1028
rect 28968 968 29032 972
rect 29128 26248 29192 26312
rect 29128 6568 29192 6632
rect 29288 31908 29352 31912
rect 29288 31852 29292 31908
rect 29292 31852 29348 31908
rect 29348 31852 29352 31908
rect 29288 31848 29352 31852
rect 29288 31748 29352 31752
rect 29288 31692 29292 31748
rect 29292 31692 29348 31748
rect 29348 31692 29352 31748
rect 29288 31688 29352 31692
rect 29288 31588 29352 31592
rect 29288 31532 29292 31588
rect 29292 31532 29348 31588
rect 29348 31532 29352 31588
rect 29288 31528 29352 31532
rect 29288 31428 29352 31432
rect 29288 31372 29292 31428
rect 29292 31372 29348 31428
rect 29348 31372 29352 31428
rect 29288 31368 29352 31372
rect 29288 31268 29352 31272
rect 29288 31212 29292 31268
rect 29292 31212 29348 31268
rect 29348 31212 29352 31268
rect 29288 31208 29352 31212
rect 29288 31108 29352 31112
rect 29288 31052 29292 31108
rect 29292 31052 29348 31108
rect 29348 31052 29352 31108
rect 29288 31048 29352 31052
rect 29288 30948 29352 30952
rect 29288 30892 29292 30948
rect 29292 30892 29348 30948
rect 29348 30892 29352 30948
rect 29288 30888 29352 30892
rect 29288 30788 29352 30792
rect 29288 30732 29292 30788
rect 29292 30732 29348 30788
rect 29348 30732 29352 30788
rect 29288 30728 29352 30732
rect 29288 30628 29352 30632
rect 29288 30572 29292 30628
rect 29292 30572 29348 30628
rect 29348 30572 29352 30628
rect 29288 30568 29352 30572
rect 29288 30468 29352 30472
rect 29288 30412 29292 30468
rect 29292 30412 29348 30468
rect 29348 30412 29352 30468
rect 29288 30408 29352 30412
rect 29288 30308 29352 30312
rect 29288 30252 29292 30308
rect 29292 30252 29348 30308
rect 29348 30252 29352 30308
rect 29288 30248 29352 30252
rect 29288 30148 29352 30152
rect 29288 30092 29292 30148
rect 29292 30092 29348 30148
rect 29348 30092 29352 30148
rect 29288 30088 29352 30092
rect 29288 29988 29352 29992
rect 29288 29932 29292 29988
rect 29292 29932 29348 29988
rect 29348 29932 29352 29988
rect 29288 29928 29352 29932
rect 29288 29828 29352 29832
rect 29288 29772 29292 29828
rect 29292 29772 29348 29828
rect 29348 29772 29352 29828
rect 29288 29768 29352 29772
rect 29288 29668 29352 29672
rect 29288 29612 29292 29668
rect 29292 29612 29348 29668
rect 29348 29612 29352 29668
rect 29288 29608 29352 29612
rect 29288 29508 29352 29512
rect 29288 29452 29292 29508
rect 29292 29452 29348 29508
rect 29348 29452 29352 29508
rect 29288 29448 29352 29452
rect 29288 29348 29352 29352
rect 29288 29292 29292 29348
rect 29292 29292 29348 29348
rect 29348 29292 29352 29348
rect 29288 29288 29352 29292
rect 29288 29028 29352 29032
rect 29288 28972 29292 29028
rect 29292 28972 29348 29028
rect 29348 28972 29352 29028
rect 29288 28968 29352 28972
rect 29288 28708 29352 28712
rect 29288 28652 29292 28708
rect 29292 28652 29348 28708
rect 29348 28652 29352 28708
rect 29288 28648 29352 28652
rect 29288 28548 29352 28552
rect 29288 28492 29292 28548
rect 29292 28492 29348 28548
rect 29348 28492 29352 28548
rect 29288 28488 29352 28492
rect 29288 28388 29352 28392
rect 29288 28332 29292 28388
rect 29292 28332 29348 28388
rect 29348 28332 29352 28388
rect 29288 28328 29352 28332
rect 29288 28228 29352 28232
rect 29288 28172 29292 28228
rect 29292 28172 29348 28228
rect 29348 28172 29352 28228
rect 29288 28168 29352 28172
rect 29288 28068 29352 28072
rect 29288 28012 29292 28068
rect 29292 28012 29348 28068
rect 29348 28012 29352 28068
rect 29288 28008 29352 28012
rect 29288 27908 29352 27912
rect 29288 27852 29292 27908
rect 29292 27852 29348 27908
rect 29348 27852 29352 27908
rect 29288 27848 29352 27852
rect 29288 27748 29352 27752
rect 29288 27692 29292 27748
rect 29292 27692 29348 27748
rect 29348 27692 29352 27748
rect 29288 27688 29352 27692
rect 29288 27588 29352 27592
rect 29288 27532 29292 27588
rect 29292 27532 29348 27588
rect 29348 27532 29352 27588
rect 29288 27528 29352 27532
rect 29288 27428 29352 27432
rect 29288 27372 29292 27428
rect 29292 27372 29348 27428
rect 29348 27372 29352 27428
rect 29288 27368 29352 27372
rect 29288 27268 29352 27272
rect 29288 27212 29292 27268
rect 29292 27212 29348 27268
rect 29348 27212 29352 27268
rect 29288 27208 29352 27212
rect 29288 27108 29352 27112
rect 29288 27052 29292 27108
rect 29292 27052 29348 27108
rect 29348 27052 29352 27108
rect 29288 27048 29352 27052
rect 29288 26948 29352 26952
rect 29288 26892 29292 26948
rect 29292 26892 29348 26948
rect 29348 26892 29352 26948
rect 29288 26888 29352 26892
rect 29288 26788 29352 26792
rect 29288 26732 29292 26788
rect 29292 26732 29348 26788
rect 29348 26732 29352 26788
rect 29288 26728 29352 26732
rect 29288 26628 29352 26632
rect 29288 26572 29292 26628
rect 29292 26572 29348 26628
rect 29348 26572 29352 26628
rect 29288 26568 29352 26572
rect 29288 26468 29352 26472
rect 29288 26412 29292 26468
rect 29292 26412 29348 26468
rect 29348 26412 29352 26468
rect 29288 26408 29352 26412
rect 29288 26308 29352 26312
rect 29288 26252 29292 26308
rect 29292 26252 29348 26308
rect 29348 26252 29352 26308
rect 29288 26248 29352 26252
rect 29288 26148 29352 26152
rect 29288 26092 29292 26148
rect 29292 26092 29348 26148
rect 29348 26092 29352 26148
rect 29288 26088 29352 26092
rect 29288 25988 29352 25992
rect 29288 25932 29292 25988
rect 29292 25932 29348 25988
rect 29348 25932 29352 25988
rect 29288 25928 29352 25932
rect 29288 25828 29352 25832
rect 29288 25772 29292 25828
rect 29292 25772 29348 25828
rect 29348 25772 29352 25828
rect 29288 25768 29352 25772
rect 29288 25668 29352 25672
rect 29288 25612 29292 25668
rect 29292 25612 29348 25668
rect 29348 25612 29352 25668
rect 29288 25608 29352 25612
rect 29288 25508 29352 25512
rect 29288 25452 29292 25508
rect 29292 25452 29348 25508
rect 29348 25452 29352 25508
rect 29288 25448 29352 25452
rect 29288 25348 29352 25352
rect 29288 25292 29292 25348
rect 29292 25292 29348 25348
rect 29348 25292 29352 25348
rect 29288 25288 29352 25292
rect 29288 25188 29352 25192
rect 29288 25132 29292 25188
rect 29292 25132 29348 25188
rect 29348 25132 29352 25188
rect 29288 25128 29352 25132
rect 29288 25028 29352 25032
rect 29288 24972 29292 25028
rect 29292 24972 29348 25028
rect 29348 24972 29352 25028
rect 29288 24968 29352 24972
rect 29288 24868 29352 24872
rect 29288 24812 29292 24868
rect 29292 24812 29348 24868
rect 29348 24812 29352 24868
rect 29288 24808 29352 24812
rect 29288 24708 29352 24712
rect 29288 24652 29292 24708
rect 29292 24652 29348 24708
rect 29348 24652 29352 24708
rect 29288 24648 29352 24652
rect 29288 24548 29352 24552
rect 29288 24492 29292 24548
rect 29292 24492 29348 24548
rect 29348 24492 29352 24548
rect 29288 24488 29352 24492
rect 29288 24388 29352 24392
rect 29288 24332 29292 24388
rect 29292 24332 29348 24388
rect 29348 24332 29352 24388
rect 29288 24328 29352 24332
rect 29288 24228 29352 24232
rect 29288 24172 29292 24228
rect 29292 24172 29348 24228
rect 29348 24172 29352 24228
rect 29288 24168 29352 24172
rect 29288 24068 29352 24072
rect 29288 24012 29292 24068
rect 29292 24012 29348 24068
rect 29348 24012 29352 24068
rect 29288 24008 29352 24012
rect 29288 23908 29352 23912
rect 29288 23852 29292 23908
rect 29292 23852 29348 23908
rect 29348 23852 29352 23908
rect 29288 23848 29352 23852
rect 29288 23588 29352 23592
rect 29288 23532 29292 23588
rect 29292 23532 29348 23588
rect 29348 23532 29352 23588
rect 29288 23528 29352 23532
rect 29288 23268 29352 23272
rect 29288 23212 29292 23268
rect 29292 23212 29348 23268
rect 29348 23212 29352 23268
rect 29288 23208 29352 23212
rect 29288 23108 29352 23112
rect 29288 23052 29292 23108
rect 29292 23052 29348 23108
rect 29348 23052 29352 23108
rect 29288 23048 29352 23052
rect 29288 22948 29352 22952
rect 29288 22892 29292 22948
rect 29292 22892 29348 22948
rect 29348 22892 29352 22948
rect 29288 22888 29352 22892
rect 29288 22788 29352 22792
rect 29288 22732 29292 22788
rect 29292 22732 29348 22788
rect 29348 22732 29352 22788
rect 29288 22728 29352 22732
rect 29288 22628 29352 22632
rect 29288 22572 29292 22628
rect 29292 22572 29348 22628
rect 29348 22572 29352 22628
rect 29288 22568 29352 22572
rect 29288 22468 29352 22472
rect 29288 22412 29292 22468
rect 29292 22412 29348 22468
rect 29348 22412 29352 22468
rect 29288 22408 29352 22412
rect 29288 22308 29352 22312
rect 29288 22252 29292 22308
rect 29292 22252 29348 22308
rect 29348 22252 29352 22308
rect 29288 22248 29352 22252
rect 29288 22148 29352 22152
rect 29288 22092 29292 22148
rect 29292 22092 29348 22148
rect 29348 22092 29352 22148
rect 29288 22088 29352 22092
rect 29288 21988 29352 21992
rect 29288 21932 29292 21988
rect 29292 21932 29348 21988
rect 29348 21932 29352 21988
rect 29288 21928 29352 21932
rect 29288 21828 29352 21832
rect 29288 21772 29292 21828
rect 29292 21772 29348 21828
rect 29348 21772 29352 21828
rect 29288 21768 29352 21772
rect 29288 21668 29352 21672
rect 29288 21612 29292 21668
rect 29292 21612 29348 21668
rect 29348 21612 29352 21668
rect 29288 21608 29352 21612
rect 29288 21508 29352 21512
rect 29288 21452 29292 21508
rect 29292 21452 29348 21508
rect 29348 21452 29352 21508
rect 29288 21448 29352 21452
rect 29288 21348 29352 21352
rect 29288 21292 29292 21348
rect 29292 21292 29348 21348
rect 29348 21292 29352 21348
rect 29288 21288 29352 21292
rect 29288 21188 29352 21192
rect 29288 21132 29292 21188
rect 29292 21132 29348 21188
rect 29348 21132 29352 21188
rect 29288 21128 29352 21132
rect 29288 21028 29352 21032
rect 29288 20972 29292 21028
rect 29292 20972 29348 21028
rect 29348 20972 29352 21028
rect 29288 20968 29352 20972
rect 29288 20868 29352 20872
rect 29288 20812 29292 20868
rect 29292 20812 29348 20868
rect 29348 20812 29352 20868
rect 29288 20808 29352 20812
rect 29288 20708 29352 20712
rect 29288 20652 29292 20708
rect 29292 20652 29348 20708
rect 29348 20652 29352 20708
rect 29288 20648 29352 20652
rect 29288 20548 29352 20552
rect 29288 20492 29292 20548
rect 29292 20492 29348 20548
rect 29348 20492 29352 20548
rect 29288 20488 29352 20492
rect 29288 20388 29352 20392
rect 29288 20332 29292 20388
rect 29292 20332 29348 20388
rect 29348 20332 29352 20388
rect 29288 20328 29352 20332
rect 29288 20228 29352 20232
rect 29288 20172 29292 20228
rect 29292 20172 29348 20228
rect 29348 20172 29352 20228
rect 29288 20168 29352 20172
rect 29288 20068 29352 20072
rect 29288 20012 29292 20068
rect 29292 20012 29348 20068
rect 29348 20012 29352 20068
rect 29288 20008 29352 20012
rect 29288 19908 29352 19912
rect 29288 19852 29292 19908
rect 29292 19852 29348 19908
rect 29348 19852 29352 19908
rect 29288 19848 29352 19852
rect 29288 19748 29352 19752
rect 29288 19692 29292 19748
rect 29292 19692 29348 19748
rect 29348 19692 29352 19748
rect 29288 19688 29352 19692
rect 29288 19588 29352 19592
rect 29288 19532 29292 19588
rect 29292 19532 29348 19588
rect 29348 19532 29352 19588
rect 29288 19528 29352 19532
rect 29288 19428 29352 19432
rect 29288 19372 29292 19428
rect 29292 19372 29348 19428
rect 29348 19372 29352 19428
rect 29288 19368 29352 19372
rect 29288 19268 29352 19272
rect 29288 19212 29292 19268
rect 29292 19212 29348 19268
rect 29348 19212 29352 19268
rect 29288 19208 29352 19212
rect 29288 19108 29352 19112
rect 29288 19052 29292 19108
rect 29292 19052 29348 19108
rect 29348 19052 29352 19108
rect 29288 19048 29352 19052
rect 29288 18948 29352 18952
rect 29288 18892 29292 18948
rect 29292 18892 29348 18948
rect 29348 18892 29352 18948
rect 29288 18888 29352 18892
rect 29288 18788 29352 18792
rect 29288 18732 29292 18788
rect 29292 18732 29348 18788
rect 29348 18732 29352 18788
rect 29288 18728 29352 18732
rect 29288 18628 29352 18632
rect 29288 18572 29292 18628
rect 29292 18572 29348 18628
rect 29348 18572 29352 18628
rect 29288 18568 29352 18572
rect 29288 18468 29352 18472
rect 29288 18412 29292 18468
rect 29292 18412 29348 18468
rect 29348 18412 29352 18468
rect 29288 18408 29352 18412
rect 29288 18308 29352 18312
rect 29288 18252 29292 18308
rect 29292 18252 29348 18308
rect 29348 18252 29352 18308
rect 29288 18248 29352 18252
rect 29288 18148 29352 18152
rect 29288 18092 29292 18148
rect 29292 18092 29348 18148
rect 29348 18092 29352 18148
rect 29288 18088 29352 18092
rect 29288 17988 29352 17992
rect 29288 17932 29292 17988
rect 29292 17932 29348 17988
rect 29348 17932 29352 17988
rect 29288 17928 29352 17932
rect 29288 17828 29352 17832
rect 29288 17772 29292 17828
rect 29292 17772 29348 17828
rect 29348 17772 29352 17828
rect 29288 17768 29352 17772
rect 29288 17668 29352 17672
rect 29288 17612 29292 17668
rect 29292 17612 29348 17668
rect 29348 17612 29352 17668
rect 29288 17608 29352 17612
rect 29288 17508 29352 17512
rect 29288 17452 29292 17508
rect 29292 17452 29348 17508
rect 29348 17452 29352 17508
rect 29288 17448 29352 17452
rect 29288 17348 29352 17352
rect 29288 17292 29292 17348
rect 29292 17292 29348 17348
rect 29348 17292 29352 17348
rect 29288 17288 29352 17292
rect 29288 17188 29352 17192
rect 29288 17132 29292 17188
rect 29292 17132 29348 17188
rect 29348 17132 29352 17188
rect 29288 17128 29352 17132
rect 29288 17028 29352 17032
rect 29288 16972 29292 17028
rect 29292 16972 29348 17028
rect 29348 16972 29352 17028
rect 29288 16968 29352 16972
rect 29288 16868 29352 16872
rect 29288 16812 29292 16868
rect 29292 16812 29348 16868
rect 29348 16812 29352 16868
rect 29288 16808 29352 16812
rect 29288 16708 29352 16712
rect 29288 16652 29292 16708
rect 29292 16652 29348 16708
rect 29348 16652 29352 16708
rect 29288 16648 29352 16652
rect 29288 16548 29352 16552
rect 29288 16492 29292 16548
rect 29292 16492 29348 16548
rect 29348 16492 29352 16548
rect 29288 16488 29352 16492
rect 29288 16388 29352 16392
rect 29288 16332 29292 16388
rect 29292 16332 29348 16388
rect 29348 16332 29352 16388
rect 29288 16328 29352 16332
rect 29288 16228 29352 16232
rect 29288 16172 29292 16228
rect 29292 16172 29348 16228
rect 29348 16172 29352 16228
rect 29288 16168 29352 16172
rect 29288 16068 29352 16072
rect 29288 16012 29292 16068
rect 29292 16012 29348 16068
rect 29348 16012 29352 16068
rect 29288 16008 29352 16012
rect 29288 15908 29352 15912
rect 29288 15852 29292 15908
rect 29292 15852 29348 15908
rect 29348 15852 29352 15908
rect 29288 15848 29352 15852
rect 29288 15748 29352 15752
rect 29288 15692 29292 15748
rect 29292 15692 29348 15748
rect 29348 15692 29352 15748
rect 29288 15688 29352 15692
rect 29288 15588 29352 15592
rect 29288 15532 29292 15588
rect 29292 15532 29348 15588
rect 29348 15532 29352 15588
rect 29288 15528 29352 15532
rect 29288 15428 29352 15432
rect 29288 15372 29292 15428
rect 29292 15372 29348 15428
rect 29348 15372 29352 15428
rect 29288 15368 29352 15372
rect 29288 15268 29352 15272
rect 29288 15212 29292 15268
rect 29292 15212 29348 15268
rect 29348 15212 29352 15268
rect 29288 15208 29352 15212
rect 29288 15108 29352 15112
rect 29288 15052 29292 15108
rect 29292 15052 29348 15108
rect 29348 15052 29352 15108
rect 29288 15048 29352 15052
rect 29288 14948 29352 14952
rect 29288 14892 29292 14948
rect 29292 14892 29348 14948
rect 29348 14892 29352 14948
rect 29288 14888 29352 14892
rect 29288 14788 29352 14792
rect 29288 14732 29292 14788
rect 29292 14732 29348 14788
rect 29348 14732 29352 14788
rect 29288 14728 29352 14732
rect 29288 14628 29352 14632
rect 29288 14572 29292 14628
rect 29292 14572 29348 14628
rect 29348 14572 29352 14628
rect 29288 14568 29352 14572
rect 29288 14468 29352 14472
rect 29288 14412 29292 14468
rect 29292 14412 29348 14468
rect 29348 14412 29352 14468
rect 29288 14408 29352 14412
rect 29288 14308 29352 14312
rect 29288 14252 29292 14308
rect 29292 14252 29348 14308
rect 29348 14252 29352 14308
rect 29288 14248 29352 14252
rect 29288 14148 29352 14152
rect 29288 14092 29292 14148
rect 29292 14092 29348 14148
rect 29348 14092 29352 14148
rect 29288 14088 29352 14092
rect 29288 13988 29352 13992
rect 29288 13932 29292 13988
rect 29292 13932 29348 13988
rect 29348 13932 29352 13988
rect 29288 13928 29352 13932
rect 29288 13828 29352 13832
rect 29288 13772 29292 13828
rect 29292 13772 29348 13828
rect 29348 13772 29352 13828
rect 29288 13768 29352 13772
rect 29288 13668 29352 13672
rect 29288 13612 29292 13668
rect 29292 13612 29348 13668
rect 29348 13612 29352 13668
rect 29288 13608 29352 13612
rect 29288 13508 29352 13512
rect 29288 13452 29292 13508
rect 29292 13452 29348 13508
rect 29348 13452 29352 13508
rect 29288 13448 29352 13452
rect 29288 13348 29352 13352
rect 29288 13292 29292 13348
rect 29292 13292 29348 13348
rect 29348 13292 29352 13348
rect 29288 13288 29352 13292
rect 29288 13188 29352 13192
rect 29288 13132 29292 13188
rect 29292 13132 29348 13188
rect 29348 13132 29352 13188
rect 29288 13128 29352 13132
rect 29288 13028 29352 13032
rect 29288 12972 29292 13028
rect 29292 12972 29348 13028
rect 29348 12972 29352 13028
rect 29288 12968 29352 12972
rect 29288 12868 29352 12872
rect 29288 12812 29292 12868
rect 29292 12812 29348 12868
rect 29348 12812 29352 12868
rect 29288 12808 29352 12812
rect 29288 12708 29352 12712
rect 29288 12652 29292 12708
rect 29292 12652 29348 12708
rect 29348 12652 29352 12708
rect 29288 12648 29352 12652
rect 29288 12548 29352 12552
rect 29288 12492 29292 12548
rect 29292 12492 29348 12548
rect 29348 12492 29352 12548
rect 29288 12488 29352 12492
rect 29288 12388 29352 12392
rect 29288 12332 29292 12388
rect 29292 12332 29348 12388
rect 29348 12332 29352 12388
rect 29288 12328 29352 12332
rect 29288 12228 29352 12232
rect 29288 12172 29292 12228
rect 29292 12172 29348 12228
rect 29348 12172 29352 12228
rect 29288 12168 29352 12172
rect 29288 12068 29352 12072
rect 29288 12012 29292 12068
rect 29292 12012 29348 12068
rect 29348 12012 29352 12068
rect 29288 12008 29352 12012
rect 29288 11908 29352 11912
rect 29288 11852 29292 11908
rect 29292 11852 29348 11908
rect 29348 11852 29352 11908
rect 29288 11848 29352 11852
rect 29288 11748 29352 11752
rect 29288 11692 29292 11748
rect 29292 11692 29348 11748
rect 29348 11692 29352 11748
rect 29288 11688 29352 11692
rect 29288 11588 29352 11592
rect 29288 11532 29292 11588
rect 29292 11532 29348 11588
rect 29348 11532 29352 11588
rect 29288 11528 29352 11532
rect 29288 11428 29352 11432
rect 29288 11372 29292 11428
rect 29292 11372 29348 11428
rect 29348 11372 29352 11428
rect 29288 11368 29352 11372
rect 29288 11268 29352 11272
rect 29288 11212 29292 11268
rect 29292 11212 29348 11268
rect 29348 11212 29352 11268
rect 29288 11208 29352 11212
rect 29288 11108 29352 11112
rect 29288 11052 29292 11108
rect 29292 11052 29348 11108
rect 29348 11052 29352 11108
rect 29288 11048 29352 11052
rect 29288 10948 29352 10952
rect 29288 10892 29292 10948
rect 29292 10892 29348 10948
rect 29348 10892 29352 10948
rect 29288 10888 29352 10892
rect 29288 10788 29352 10792
rect 29288 10732 29292 10788
rect 29292 10732 29348 10788
rect 29348 10732 29352 10788
rect 29288 10728 29352 10732
rect 29288 10628 29352 10632
rect 29288 10572 29292 10628
rect 29292 10572 29348 10628
rect 29348 10572 29352 10628
rect 29288 10568 29352 10572
rect 29288 10468 29352 10472
rect 29288 10412 29292 10468
rect 29292 10412 29348 10468
rect 29348 10412 29352 10468
rect 29288 10408 29352 10412
rect 29288 10308 29352 10312
rect 29288 10252 29292 10308
rect 29292 10252 29348 10308
rect 29348 10252 29352 10308
rect 29288 10248 29352 10252
rect 29288 10148 29352 10152
rect 29288 10092 29292 10148
rect 29292 10092 29348 10148
rect 29348 10092 29352 10148
rect 29288 10088 29352 10092
rect 29288 9988 29352 9992
rect 29288 9932 29292 9988
rect 29292 9932 29348 9988
rect 29348 9932 29352 9988
rect 29288 9928 29352 9932
rect 29288 9828 29352 9832
rect 29288 9772 29292 9828
rect 29292 9772 29348 9828
rect 29348 9772 29352 9828
rect 29288 9768 29352 9772
rect 29288 9668 29352 9672
rect 29288 9612 29292 9668
rect 29292 9612 29348 9668
rect 29348 9612 29352 9668
rect 29288 9608 29352 9612
rect 29288 9348 29352 9352
rect 29288 9292 29292 9348
rect 29292 9292 29348 9348
rect 29348 9292 29352 9348
rect 29288 9288 29352 9292
rect 29288 9028 29352 9032
rect 29288 8972 29292 9028
rect 29292 8972 29348 9028
rect 29348 8972 29352 9028
rect 29288 8968 29352 8972
rect 29288 8868 29352 8872
rect 29288 8812 29292 8868
rect 29292 8812 29348 8868
rect 29348 8812 29352 8868
rect 29288 8808 29352 8812
rect 29288 8708 29352 8712
rect 29288 8652 29292 8708
rect 29292 8652 29348 8708
rect 29348 8652 29352 8708
rect 29288 8648 29352 8652
rect 29288 8548 29352 8552
rect 29288 8492 29292 8548
rect 29292 8492 29348 8548
rect 29348 8492 29352 8548
rect 29288 8488 29352 8492
rect 29288 8388 29352 8392
rect 29288 8332 29292 8388
rect 29292 8332 29348 8388
rect 29348 8332 29352 8388
rect 29288 8328 29352 8332
rect 29288 8228 29352 8232
rect 29288 8172 29292 8228
rect 29292 8172 29348 8228
rect 29348 8172 29352 8228
rect 29288 8168 29352 8172
rect 29288 8068 29352 8072
rect 29288 8012 29292 8068
rect 29292 8012 29348 8068
rect 29348 8012 29352 8068
rect 29288 8008 29352 8012
rect 29288 7908 29352 7912
rect 29288 7852 29292 7908
rect 29292 7852 29348 7908
rect 29348 7852 29352 7908
rect 29288 7848 29352 7852
rect 29288 7748 29352 7752
rect 29288 7692 29292 7748
rect 29292 7692 29348 7748
rect 29348 7692 29352 7748
rect 29288 7688 29352 7692
rect 29288 7588 29352 7592
rect 29288 7532 29292 7588
rect 29292 7532 29348 7588
rect 29348 7532 29352 7588
rect 29288 7528 29352 7532
rect 29288 7428 29352 7432
rect 29288 7372 29292 7428
rect 29292 7372 29348 7428
rect 29348 7372 29352 7428
rect 29288 7368 29352 7372
rect 29288 7268 29352 7272
rect 29288 7212 29292 7268
rect 29292 7212 29348 7268
rect 29348 7212 29352 7268
rect 29288 7208 29352 7212
rect 29288 7108 29352 7112
rect 29288 7052 29292 7108
rect 29292 7052 29348 7108
rect 29348 7052 29352 7108
rect 29288 7048 29352 7052
rect 29288 6948 29352 6952
rect 29288 6892 29292 6948
rect 29292 6892 29348 6948
rect 29348 6892 29352 6948
rect 29288 6888 29352 6892
rect 29288 6788 29352 6792
rect 29288 6732 29292 6788
rect 29292 6732 29348 6788
rect 29348 6732 29352 6788
rect 29288 6728 29352 6732
rect 29288 6628 29352 6632
rect 29288 6572 29292 6628
rect 29292 6572 29348 6628
rect 29348 6572 29352 6628
rect 29288 6568 29352 6572
rect 29288 6468 29352 6472
rect 29288 6412 29292 6468
rect 29292 6412 29348 6468
rect 29348 6412 29352 6468
rect 29288 6408 29352 6412
rect 29288 6308 29352 6312
rect 29288 6252 29292 6308
rect 29292 6252 29348 6308
rect 29348 6252 29352 6308
rect 29288 6248 29352 6252
rect 29288 6148 29352 6152
rect 29288 6092 29292 6148
rect 29292 6092 29348 6148
rect 29348 6092 29352 6148
rect 29288 6088 29352 6092
rect 29288 5988 29352 5992
rect 29288 5932 29292 5988
rect 29292 5932 29348 5988
rect 29348 5932 29352 5988
rect 29288 5928 29352 5932
rect 29288 5828 29352 5832
rect 29288 5772 29292 5828
rect 29292 5772 29348 5828
rect 29348 5772 29352 5828
rect 29288 5768 29352 5772
rect 29288 5668 29352 5672
rect 29288 5612 29292 5668
rect 29292 5612 29348 5668
rect 29348 5612 29352 5668
rect 29288 5608 29352 5612
rect 29288 5508 29352 5512
rect 29288 5452 29292 5508
rect 29292 5452 29348 5508
rect 29348 5452 29352 5508
rect 29288 5448 29352 5452
rect 29288 5348 29352 5352
rect 29288 5292 29292 5348
rect 29292 5292 29348 5348
rect 29348 5292 29352 5348
rect 29288 5288 29352 5292
rect 29288 5188 29352 5192
rect 29288 5132 29292 5188
rect 29292 5132 29348 5188
rect 29348 5132 29352 5188
rect 29288 5128 29352 5132
rect 29288 5028 29352 5032
rect 29288 4972 29292 5028
rect 29292 4972 29348 5028
rect 29348 4972 29352 5028
rect 29288 4968 29352 4972
rect 29288 4868 29352 4872
rect 29288 4812 29292 4868
rect 29292 4812 29348 4868
rect 29348 4812 29352 4868
rect 29288 4808 29352 4812
rect 29288 4708 29352 4712
rect 29288 4652 29292 4708
rect 29292 4652 29348 4708
rect 29348 4652 29352 4708
rect 29288 4648 29352 4652
rect 29288 4548 29352 4552
rect 29288 4492 29292 4548
rect 29292 4492 29348 4548
rect 29348 4492 29352 4548
rect 29288 4488 29352 4492
rect 29288 4388 29352 4392
rect 29288 4332 29292 4388
rect 29292 4332 29348 4388
rect 29348 4332 29352 4388
rect 29288 4328 29352 4332
rect 29288 4228 29352 4232
rect 29288 4172 29292 4228
rect 29292 4172 29348 4228
rect 29348 4172 29352 4228
rect 29288 4168 29352 4172
rect 29288 3908 29352 3912
rect 29288 3852 29292 3908
rect 29292 3852 29348 3908
rect 29348 3852 29352 3908
rect 29288 3848 29352 3852
rect 29288 3588 29352 3592
rect 29288 3532 29292 3588
rect 29292 3532 29348 3588
rect 29348 3532 29352 3588
rect 29288 3528 29352 3532
rect 29288 3428 29352 3432
rect 29288 3372 29292 3428
rect 29292 3372 29348 3428
rect 29348 3372 29352 3428
rect 29288 3368 29352 3372
rect 29288 3268 29352 3272
rect 29288 3212 29292 3268
rect 29292 3212 29348 3268
rect 29348 3212 29352 3268
rect 29288 3208 29352 3212
rect 29288 3108 29352 3112
rect 29288 3052 29292 3108
rect 29292 3052 29348 3108
rect 29348 3052 29352 3108
rect 29288 3048 29352 3052
rect 29288 2948 29352 2952
rect 29288 2892 29292 2948
rect 29292 2892 29348 2948
rect 29348 2892 29352 2948
rect 29288 2888 29352 2892
rect 29288 2788 29352 2792
rect 29288 2732 29292 2788
rect 29292 2732 29348 2788
rect 29348 2732 29352 2788
rect 29288 2728 29352 2732
rect 29288 2628 29352 2632
rect 29288 2572 29292 2628
rect 29292 2572 29348 2628
rect 29348 2572 29352 2628
rect 29288 2568 29352 2572
rect 29288 2468 29352 2472
rect 29288 2412 29292 2468
rect 29292 2412 29348 2468
rect 29348 2412 29352 2468
rect 29288 2408 29352 2412
rect 29288 2308 29352 2312
rect 29288 2252 29292 2308
rect 29292 2252 29348 2308
rect 29348 2252 29352 2308
rect 29288 2248 29352 2252
rect 29288 2148 29352 2152
rect 29288 2092 29292 2148
rect 29292 2092 29348 2148
rect 29348 2092 29352 2148
rect 29288 2088 29352 2092
rect 29288 1988 29352 1992
rect 29288 1932 29292 1988
rect 29292 1932 29348 1988
rect 29348 1932 29352 1988
rect 29288 1928 29352 1932
rect 29288 1828 29352 1832
rect 29288 1772 29292 1828
rect 29292 1772 29348 1828
rect 29348 1772 29352 1828
rect 29288 1768 29352 1772
rect 29288 1668 29352 1672
rect 29288 1612 29292 1668
rect 29292 1612 29348 1668
rect 29348 1612 29352 1668
rect 29288 1608 29352 1612
rect 29288 1508 29352 1512
rect 29288 1452 29292 1508
rect 29292 1452 29348 1508
rect 29348 1452 29352 1508
rect 29288 1448 29352 1452
rect 29288 1348 29352 1352
rect 29288 1292 29292 1348
rect 29292 1292 29348 1348
rect 29348 1292 29352 1348
rect 29288 1288 29352 1292
rect 29288 1188 29352 1192
rect 29288 1132 29292 1188
rect 29292 1132 29348 1188
rect 29348 1132 29352 1188
rect 29288 1128 29352 1132
rect 29288 1028 29352 1032
rect 29288 972 29292 1028
rect 29292 972 29348 1028
rect 29348 972 29352 1028
rect 29288 968 29352 972
rect 28968 808 29032 872
rect 28968 728 29032 792
rect 28968 648 29032 712
rect 28968 568 29032 632
rect 28968 488 29032 552
rect 29448 28808 29512 28872
rect 29448 23688 29512 23752
rect 29448 9128 29512 9192
rect 29448 4008 29512 4072
rect 29608 31908 29672 31912
rect 29608 31852 29612 31908
rect 29612 31852 29668 31908
rect 29668 31852 29672 31908
rect 29608 31848 29672 31852
rect 29608 31748 29672 31752
rect 29608 31692 29612 31748
rect 29612 31692 29668 31748
rect 29668 31692 29672 31748
rect 29608 31688 29672 31692
rect 29608 31588 29672 31592
rect 29608 31532 29612 31588
rect 29612 31532 29668 31588
rect 29668 31532 29672 31588
rect 29608 31528 29672 31532
rect 29608 31428 29672 31432
rect 29608 31372 29612 31428
rect 29612 31372 29668 31428
rect 29668 31372 29672 31428
rect 29608 31368 29672 31372
rect 29608 31268 29672 31272
rect 29608 31212 29612 31268
rect 29612 31212 29668 31268
rect 29668 31212 29672 31268
rect 29608 31208 29672 31212
rect 29608 31108 29672 31112
rect 29608 31052 29612 31108
rect 29612 31052 29668 31108
rect 29668 31052 29672 31108
rect 29608 31048 29672 31052
rect 29608 30948 29672 30952
rect 29608 30892 29612 30948
rect 29612 30892 29668 30948
rect 29668 30892 29672 30948
rect 29608 30888 29672 30892
rect 29608 30788 29672 30792
rect 29608 30732 29612 30788
rect 29612 30732 29668 30788
rect 29668 30732 29672 30788
rect 29608 30728 29672 30732
rect 29608 30628 29672 30632
rect 29608 30572 29612 30628
rect 29612 30572 29668 30628
rect 29668 30572 29672 30628
rect 29608 30568 29672 30572
rect 29608 30468 29672 30472
rect 29608 30412 29612 30468
rect 29612 30412 29668 30468
rect 29668 30412 29672 30468
rect 29608 30408 29672 30412
rect 29608 30308 29672 30312
rect 29608 30252 29612 30308
rect 29612 30252 29668 30308
rect 29668 30252 29672 30308
rect 29608 30248 29672 30252
rect 29608 30148 29672 30152
rect 29608 30092 29612 30148
rect 29612 30092 29668 30148
rect 29668 30092 29672 30148
rect 29608 30088 29672 30092
rect 29608 29988 29672 29992
rect 29608 29932 29612 29988
rect 29612 29932 29668 29988
rect 29668 29932 29672 29988
rect 29608 29928 29672 29932
rect 29608 29828 29672 29832
rect 29608 29772 29612 29828
rect 29612 29772 29668 29828
rect 29668 29772 29672 29828
rect 29608 29768 29672 29772
rect 29608 29668 29672 29672
rect 29608 29612 29612 29668
rect 29612 29612 29668 29668
rect 29668 29612 29672 29668
rect 29608 29608 29672 29612
rect 29608 29508 29672 29512
rect 29608 29452 29612 29508
rect 29612 29452 29668 29508
rect 29668 29452 29672 29508
rect 29608 29448 29672 29452
rect 29608 29348 29672 29352
rect 29608 29292 29612 29348
rect 29612 29292 29668 29348
rect 29668 29292 29672 29348
rect 29608 29288 29672 29292
rect 29608 29028 29672 29032
rect 29608 28972 29612 29028
rect 29612 28972 29668 29028
rect 29668 28972 29672 29028
rect 29608 28968 29672 28972
rect 29608 28868 29672 28872
rect 29608 28812 29612 28868
rect 29612 28812 29668 28868
rect 29668 28812 29672 28868
rect 29608 28808 29672 28812
rect 29608 28708 29672 28712
rect 29608 28652 29612 28708
rect 29612 28652 29668 28708
rect 29668 28652 29672 28708
rect 29608 28648 29672 28652
rect 29608 28548 29672 28552
rect 29608 28492 29612 28548
rect 29612 28492 29668 28548
rect 29668 28492 29672 28548
rect 29608 28488 29672 28492
rect 29608 28388 29672 28392
rect 29608 28332 29612 28388
rect 29612 28332 29668 28388
rect 29668 28332 29672 28388
rect 29608 28328 29672 28332
rect 29608 28228 29672 28232
rect 29608 28172 29612 28228
rect 29612 28172 29668 28228
rect 29668 28172 29672 28228
rect 29608 28168 29672 28172
rect 29608 28068 29672 28072
rect 29608 28012 29612 28068
rect 29612 28012 29668 28068
rect 29668 28012 29672 28068
rect 29608 28008 29672 28012
rect 29608 27908 29672 27912
rect 29608 27852 29612 27908
rect 29612 27852 29668 27908
rect 29668 27852 29672 27908
rect 29608 27848 29672 27852
rect 29608 27748 29672 27752
rect 29608 27692 29612 27748
rect 29612 27692 29668 27748
rect 29668 27692 29672 27748
rect 29608 27688 29672 27692
rect 29608 27588 29672 27592
rect 29608 27532 29612 27588
rect 29612 27532 29668 27588
rect 29668 27532 29672 27588
rect 29608 27528 29672 27532
rect 29608 27428 29672 27432
rect 29608 27372 29612 27428
rect 29612 27372 29668 27428
rect 29668 27372 29672 27428
rect 29608 27368 29672 27372
rect 29608 27268 29672 27272
rect 29608 27212 29612 27268
rect 29612 27212 29668 27268
rect 29668 27212 29672 27268
rect 29608 27208 29672 27212
rect 29608 27108 29672 27112
rect 29608 27052 29612 27108
rect 29612 27052 29668 27108
rect 29668 27052 29672 27108
rect 29608 27048 29672 27052
rect 29608 26948 29672 26952
rect 29608 26892 29612 26948
rect 29612 26892 29668 26948
rect 29668 26892 29672 26948
rect 29608 26888 29672 26892
rect 29608 26788 29672 26792
rect 29608 26732 29612 26788
rect 29612 26732 29668 26788
rect 29668 26732 29672 26788
rect 29608 26728 29672 26732
rect 29608 26628 29672 26632
rect 29608 26572 29612 26628
rect 29612 26572 29668 26628
rect 29668 26572 29672 26628
rect 29608 26568 29672 26572
rect 29608 26468 29672 26472
rect 29608 26412 29612 26468
rect 29612 26412 29668 26468
rect 29668 26412 29672 26468
rect 29608 26408 29672 26412
rect 29608 26308 29672 26312
rect 29608 26252 29612 26308
rect 29612 26252 29668 26308
rect 29668 26252 29672 26308
rect 29608 26248 29672 26252
rect 29608 26148 29672 26152
rect 29608 26092 29612 26148
rect 29612 26092 29668 26148
rect 29668 26092 29672 26148
rect 29608 26088 29672 26092
rect 29608 25988 29672 25992
rect 29608 25932 29612 25988
rect 29612 25932 29668 25988
rect 29668 25932 29672 25988
rect 29608 25928 29672 25932
rect 29608 25828 29672 25832
rect 29608 25772 29612 25828
rect 29612 25772 29668 25828
rect 29668 25772 29672 25828
rect 29608 25768 29672 25772
rect 29608 25668 29672 25672
rect 29608 25612 29612 25668
rect 29612 25612 29668 25668
rect 29668 25612 29672 25668
rect 29608 25608 29672 25612
rect 29608 25508 29672 25512
rect 29608 25452 29612 25508
rect 29612 25452 29668 25508
rect 29668 25452 29672 25508
rect 29608 25448 29672 25452
rect 29608 25348 29672 25352
rect 29608 25292 29612 25348
rect 29612 25292 29668 25348
rect 29668 25292 29672 25348
rect 29608 25288 29672 25292
rect 29608 25188 29672 25192
rect 29608 25132 29612 25188
rect 29612 25132 29668 25188
rect 29668 25132 29672 25188
rect 29608 25128 29672 25132
rect 29608 25028 29672 25032
rect 29608 24972 29612 25028
rect 29612 24972 29668 25028
rect 29668 24972 29672 25028
rect 29608 24968 29672 24972
rect 29608 24868 29672 24872
rect 29608 24812 29612 24868
rect 29612 24812 29668 24868
rect 29668 24812 29672 24868
rect 29608 24808 29672 24812
rect 29608 24708 29672 24712
rect 29608 24652 29612 24708
rect 29612 24652 29668 24708
rect 29668 24652 29672 24708
rect 29608 24648 29672 24652
rect 29608 24548 29672 24552
rect 29608 24492 29612 24548
rect 29612 24492 29668 24548
rect 29668 24492 29672 24548
rect 29608 24488 29672 24492
rect 29608 24388 29672 24392
rect 29608 24332 29612 24388
rect 29612 24332 29668 24388
rect 29668 24332 29672 24388
rect 29608 24328 29672 24332
rect 29608 24228 29672 24232
rect 29608 24172 29612 24228
rect 29612 24172 29668 24228
rect 29668 24172 29672 24228
rect 29608 24168 29672 24172
rect 29608 24068 29672 24072
rect 29608 24012 29612 24068
rect 29612 24012 29668 24068
rect 29668 24012 29672 24068
rect 29608 24008 29672 24012
rect 29608 23908 29672 23912
rect 29608 23852 29612 23908
rect 29612 23852 29668 23908
rect 29668 23852 29672 23908
rect 29608 23848 29672 23852
rect 29608 23748 29672 23752
rect 29608 23692 29612 23748
rect 29612 23692 29668 23748
rect 29668 23692 29672 23748
rect 29608 23688 29672 23692
rect 29608 23588 29672 23592
rect 29608 23532 29612 23588
rect 29612 23532 29668 23588
rect 29668 23532 29672 23588
rect 29608 23528 29672 23532
rect 29608 23268 29672 23272
rect 29608 23212 29612 23268
rect 29612 23212 29668 23268
rect 29668 23212 29672 23268
rect 29608 23208 29672 23212
rect 29608 23108 29672 23112
rect 29608 23052 29612 23108
rect 29612 23052 29668 23108
rect 29668 23052 29672 23108
rect 29608 23048 29672 23052
rect 29608 22948 29672 22952
rect 29608 22892 29612 22948
rect 29612 22892 29668 22948
rect 29668 22892 29672 22948
rect 29608 22888 29672 22892
rect 29608 22788 29672 22792
rect 29608 22732 29612 22788
rect 29612 22732 29668 22788
rect 29668 22732 29672 22788
rect 29608 22728 29672 22732
rect 29608 22628 29672 22632
rect 29608 22572 29612 22628
rect 29612 22572 29668 22628
rect 29668 22572 29672 22628
rect 29608 22568 29672 22572
rect 29608 22468 29672 22472
rect 29608 22412 29612 22468
rect 29612 22412 29668 22468
rect 29668 22412 29672 22468
rect 29608 22408 29672 22412
rect 29608 22308 29672 22312
rect 29608 22252 29612 22308
rect 29612 22252 29668 22308
rect 29668 22252 29672 22308
rect 29608 22248 29672 22252
rect 29608 22148 29672 22152
rect 29608 22092 29612 22148
rect 29612 22092 29668 22148
rect 29668 22092 29672 22148
rect 29608 22088 29672 22092
rect 29608 21988 29672 21992
rect 29608 21932 29612 21988
rect 29612 21932 29668 21988
rect 29668 21932 29672 21988
rect 29608 21928 29672 21932
rect 29608 21828 29672 21832
rect 29608 21772 29612 21828
rect 29612 21772 29668 21828
rect 29668 21772 29672 21828
rect 29608 21768 29672 21772
rect 29608 21668 29672 21672
rect 29608 21612 29612 21668
rect 29612 21612 29668 21668
rect 29668 21612 29672 21668
rect 29608 21608 29672 21612
rect 29608 21508 29672 21512
rect 29608 21452 29612 21508
rect 29612 21452 29668 21508
rect 29668 21452 29672 21508
rect 29608 21448 29672 21452
rect 29608 21348 29672 21352
rect 29608 21292 29612 21348
rect 29612 21292 29668 21348
rect 29668 21292 29672 21348
rect 29608 21288 29672 21292
rect 29608 21188 29672 21192
rect 29608 21132 29612 21188
rect 29612 21132 29668 21188
rect 29668 21132 29672 21188
rect 29608 21128 29672 21132
rect 29608 21028 29672 21032
rect 29608 20972 29612 21028
rect 29612 20972 29668 21028
rect 29668 20972 29672 21028
rect 29608 20968 29672 20972
rect 29608 20868 29672 20872
rect 29608 20812 29612 20868
rect 29612 20812 29668 20868
rect 29668 20812 29672 20868
rect 29608 20808 29672 20812
rect 29608 20708 29672 20712
rect 29608 20652 29612 20708
rect 29612 20652 29668 20708
rect 29668 20652 29672 20708
rect 29608 20648 29672 20652
rect 29608 20548 29672 20552
rect 29608 20492 29612 20548
rect 29612 20492 29668 20548
rect 29668 20492 29672 20548
rect 29608 20488 29672 20492
rect 29608 20388 29672 20392
rect 29608 20332 29612 20388
rect 29612 20332 29668 20388
rect 29668 20332 29672 20388
rect 29608 20328 29672 20332
rect 29608 20228 29672 20232
rect 29608 20172 29612 20228
rect 29612 20172 29668 20228
rect 29668 20172 29672 20228
rect 29608 20168 29672 20172
rect 29608 20068 29672 20072
rect 29608 20012 29612 20068
rect 29612 20012 29668 20068
rect 29668 20012 29672 20068
rect 29608 20008 29672 20012
rect 29608 19908 29672 19912
rect 29608 19852 29612 19908
rect 29612 19852 29668 19908
rect 29668 19852 29672 19908
rect 29608 19848 29672 19852
rect 29608 19748 29672 19752
rect 29608 19692 29612 19748
rect 29612 19692 29668 19748
rect 29668 19692 29672 19748
rect 29608 19688 29672 19692
rect 29608 19588 29672 19592
rect 29608 19532 29612 19588
rect 29612 19532 29668 19588
rect 29668 19532 29672 19588
rect 29608 19528 29672 19532
rect 29608 19428 29672 19432
rect 29608 19372 29612 19428
rect 29612 19372 29668 19428
rect 29668 19372 29672 19428
rect 29608 19368 29672 19372
rect 29608 19268 29672 19272
rect 29608 19212 29612 19268
rect 29612 19212 29668 19268
rect 29668 19212 29672 19268
rect 29608 19208 29672 19212
rect 29608 19108 29672 19112
rect 29608 19052 29612 19108
rect 29612 19052 29668 19108
rect 29668 19052 29672 19108
rect 29608 19048 29672 19052
rect 29608 18948 29672 18952
rect 29608 18892 29612 18948
rect 29612 18892 29668 18948
rect 29668 18892 29672 18948
rect 29608 18888 29672 18892
rect 29608 18788 29672 18792
rect 29608 18732 29612 18788
rect 29612 18732 29668 18788
rect 29668 18732 29672 18788
rect 29608 18728 29672 18732
rect 29608 18628 29672 18632
rect 29608 18572 29612 18628
rect 29612 18572 29668 18628
rect 29668 18572 29672 18628
rect 29608 18568 29672 18572
rect 29608 18468 29672 18472
rect 29608 18412 29612 18468
rect 29612 18412 29668 18468
rect 29668 18412 29672 18468
rect 29608 18408 29672 18412
rect 29608 18308 29672 18312
rect 29608 18252 29612 18308
rect 29612 18252 29668 18308
rect 29668 18252 29672 18308
rect 29608 18248 29672 18252
rect 29608 18148 29672 18152
rect 29608 18092 29612 18148
rect 29612 18092 29668 18148
rect 29668 18092 29672 18148
rect 29608 18088 29672 18092
rect 29608 17988 29672 17992
rect 29608 17932 29612 17988
rect 29612 17932 29668 17988
rect 29668 17932 29672 17988
rect 29608 17928 29672 17932
rect 29608 17828 29672 17832
rect 29608 17772 29612 17828
rect 29612 17772 29668 17828
rect 29668 17772 29672 17828
rect 29608 17768 29672 17772
rect 29608 17668 29672 17672
rect 29608 17612 29612 17668
rect 29612 17612 29668 17668
rect 29668 17612 29672 17668
rect 29608 17608 29672 17612
rect 29608 17508 29672 17512
rect 29608 17452 29612 17508
rect 29612 17452 29668 17508
rect 29668 17452 29672 17508
rect 29608 17448 29672 17452
rect 29608 17348 29672 17352
rect 29608 17292 29612 17348
rect 29612 17292 29668 17348
rect 29668 17292 29672 17348
rect 29608 17288 29672 17292
rect 29608 17188 29672 17192
rect 29608 17132 29612 17188
rect 29612 17132 29668 17188
rect 29668 17132 29672 17188
rect 29608 17128 29672 17132
rect 29608 17028 29672 17032
rect 29608 16972 29612 17028
rect 29612 16972 29668 17028
rect 29668 16972 29672 17028
rect 29608 16968 29672 16972
rect 29608 16868 29672 16872
rect 29608 16812 29612 16868
rect 29612 16812 29668 16868
rect 29668 16812 29672 16868
rect 29608 16808 29672 16812
rect 29608 16708 29672 16712
rect 29608 16652 29612 16708
rect 29612 16652 29668 16708
rect 29668 16652 29672 16708
rect 29608 16648 29672 16652
rect 29608 16548 29672 16552
rect 29608 16492 29612 16548
rect 29612 16492 29668 16548
rect 29668 16492 29672 16548
rect 29608 16488 29672 16492
rect 29608 16388 29672 16392
rect 29608 16332 29612 16388
rect 29612 16332 29668 16388
rect 29668 16332 29672 16388
rect 29608 16328 29672 16332
rect 29608 16228 29672 16232
rect 29608 16172 29612 16228
rect 29612 16172 29668 16228
rect 29668 16172 29672 16228
rect 29608 16168 29672 16172
rect 29608 16068 29672 16072
rect 29608 16012 29612 16068
rect 29612 16012 29668 16068
rect 29668 16012 29672 16068
rect 29608 16008 29672 16012
rect 29608 15908 29672 15912
rect 29608 15852 29612 15908
rect 29612 15852 29668 15908
rect 29668 15852 29672 15908
rect 29608 15848 29672 15852
rect 29608 15748 29672 15752
rect 29608 15692 29612 15748
rect 29612 15692 29668 15748
rect 29668 15692 29672 15748
rect 29608 15688 29672 15692
rect 29608 15588 29672 15592
rect 29608 15532 29612 15588
rect 29612 15532 29668 15588
rect 29668 15532 29672 15588
rect 29608 15528 29672 15532
rect 29608 15428 29672 15432
rect 29608 15372 29612 15428
rect 29612 15372 29668 15428
rect 29668 15372 29672 15428
rect 29608 15368 29672 15372
rect 29608 15268 29672 15272
rect 29608 15212 29612 15268
rect 29612 15212 29668 15268
rect 29668 15212 29672 15268
rect 29608 15208 29672 15212
rect 29608 15108 29672 15112
rect 29608 15052 29612 15108
rect 29612 15052 29668 15108
rect 29668 15052 29672 15108
rect 29608 15048 29672 15052
rect 29608 14948 29672 14952
rect 29608 14892 29612 14948
rect 29612 14892 29668 14948
rect 29668 14892 29672 14948
rect 29608 14888 29672 14892
rect 29608 14788 29672 14792
rect 29608 14732 29612 14788
rect 29612 14732 29668 14788
rect 29668 14732 29672 14788
rect 29608 14728 29672 14732
rect 29608 14628 29672 14632
rect 29608 14572 29612 14628
rect 29612 14572 29668 14628
rect 29668 14572 29672 14628
rect 29608 14568 29672 14572
rect 29608 14468 29672 14472
rect 29608 14412 29612 14468
rect 29612 14412 29668 14468
rect 29668 14412 29672 14468
rect 29608 14408 29672 14412
rect 29608 14308 29672 14312
rect 29608 14252 29612 14308
rect 29612 14252 29668 14308
rect 29668 14252 29672 14308
rect 29608 14248 29672 14252
rect 29608 14148 29672 14152
rect 29608 14092 29612 14148
rect 29612 14092 29668 14148
rect 29668 14092 29672 14148
rect 29608 14088 29672 14092
rect 29608 13988 29672 13992
rect 29608 13932 29612 13988
rect 29612 13932 29668 13988
rect 29668 13932 29672 13988
rect 29608 13928 29672 13932
rect 29608 13828 29672 13832
rect 29608 13772 29612 13828
rect 29612 13772 29668 13828
rect 29668 13772 29672 13828
rect 29608 13768 29672 13772
rect 29608 13668 29672 13672
rect 29608 13612 29612 13668
rect 29612 13612 29668 13668
rect 29668 13612 29672 13668
rect 29608 13608 29672 13612
rect 29608 13508 29672 13512
rect 29608 13452 29612 13508
rect 29612 13452 29668 13508
rect 29668 13452 29672 13508
rect 29608 13448 29672 13452
rect 29608 13348 29672 13352
rect 29608 13292 29612 13348
rect 29612 13292 29668 13348
rect 29668 13292 29672 13348
rect 29608 13288 29672 13292
rect 29608 13188 29672 13192
rect 29608 13132 29612 13188
rect 29612 13132 29668 13188
rect 29668 13132 29672 13188
rect 29608 13128 29672 13132
rect 29608 13028 29672 13032
rect 29608 12972 29612 13028
rect 29612 12972 29668 13028
rect 29668 12972 29672 13028
rect 29608 12968 29672 12972
rect 29608 12868 29672 12872
rect 29608 12812 29612 12868
rect 29612 12812 29668 12868
rect 29668 12812 29672 12868
rect 29608 12808 29672 12812
rect 29608 12708 29672 12712
rect 29608 12652 29612 12708
rect 29612 12652 29668 12708
rect 29668 12652 29672 12708
rect 29608 12648 29672 12652
rect 29608 12548 29672 12552
rect 29608 12492 29612 12548
rect 29612 12492 29668 12548
rect 29668 12492 29672 12548
rect 29608 12488 29672 12492
rect 29608 12388 29672 12392
rect 29608 12332 29612 12388
rect 29612 12332 29668 12388
rect 29668 12332 29672 12388
rect 29608 12328 29672 12332
rect 29608 12228 29672 12232
rect 29608 12172 29612 12228
rect 29612 12172 29668 12228
rect 29668 12172 29672 12228
rect 29608 12168 29672 12172
rect 29608 12068 29672 12072
rect 29608 12012 29612 12068
rect 29612 12012 29668 12068
rect 29668 12012 29672 12068
rect 29608 12008 29672 12012
rect 29608 11908 29672 11912
rect 29608 11852 29612 11908
rect 29612 11852 29668 11908
rect 29668 11852 29672 11908
rect 29608 11848 29672 11852
rect 29608 11748 29672 11752
rect 29608 11692 29612 11748
rect 29612 11692 29668 11748
rect 29668 11692 29672 11748
rect 29608 11688 29672 11692
rect 29608 11588 29672 11592
rect 29608 11532 29612 11588
rect 29612 11532 29668 11588
rect 29668 11532 29672 11588
rect 29608 11528 29672 11532
rect 29608 11428 29672 11432
rect 29608 11372 29612 11428
rect 29612 11372 29668 11428
rect 29668 11372 29672 11428
rect 29608 11368 29672 11372
rect 29608 11268 29672 11272
rect 29608 11212 29612 11268
rect 29612 11212 29668 11268
rect 29668 11212 29672 11268
rect 29608 11208 29672 11212
rect 29608 11108 29672 11112
rect 29608 11052 29612 11108
rect 29612 11052 29668 11108
rect 29668 11052 29672 11108
rect 29608 11048 29672 11052
rect 29608 10948 29672 10952
rect 29608 10892 29612 10948
rect 29612 10892 29668 10948
rect 29668 10892 29672 10948
rect 29608 10888 29672 10892
rect 29608 10788 29672 10792
rect 29608 10732 29612 10788
rect 29612 10732 29668 10788
rect 29668 10732 29672 10788
rect 29608 10728 29672 10732
rect 29608 10628 29672 10632
rect 29608 10572 29612 10628
rect 29612 10572 29668 10628
rect 29668 10572 29672 10628
rect 29608 10568 29672 10572
rect 29608 10468 29672 10472
rect 29608 10412 29612 10468
rect 29612 10412 29668 10468
rect 29668 10412 29672 10468
rect 29608 10408 29672 10412
rect 29608 10308 29672 10312
rect 29608 10252 29612 10308
rect 29612 10252 29668 10308
rect 29668 10252 29672 10308
rect 29608 10248 29672 10252
rect 29608 10148 29672 10152
rect 29608 10092 29612 10148
rect 29612 10092 29668 10148
rect 29668 10092 29672 10148
rect 29608 10088 29672 10092
rect 29608 9988 29672 9992
rect 29608 9932 29612 9988
rect 29612 9932 29668 9988
rect 29668 9932 29672 9988
rect 29608 9928 29672 9932
rect 29608 9828 29672 9832
rect 29608 9772 29612 9828
rect 29612 9772 29668 9828
rect 29668 9772 29672 9828
rect 29608 9768 29672 9772
rect 29608 9668 29672 9672
rect 29608 9612 29612 9668
rect 29612 9612 29668 9668
rect 29668 9612 29672 9668
rect 29608 9608 29672 9612
rect 29608 9348 29672 9352
rect 29608 9292 29612 9348
rect 29612 9292 29668 9348
rect 29668 9292 29672 9348
rect 29608 9288 29672 9292
rect 29608 9188 29672 9192
rect 29608 9132 29612 9188
rect 29612 9132 29668 9188
rect 29668 9132 29672 9188
rect 29608 9128 29672 9132
rect 29608 9028 29672 9032
rect 29608 8972 29612 9028
rect 29612 8972 29668 9028
rect 29668 8972 29672 9028
rect 29608 8968 29672 8972
rect 29608 8868 29672 8872
rect 29608 8812 29612 8868
rect 29612 8812 29668 8868
rect 29668 8812 29672 8868
rect 29608 8808 29672 8812
rect 29608 8708 29672 8712
rect 29608 8652 29612 8708
rect 29612 8652 29668 8708
rect 29668 8652 29672 8708
rect 29608 8648 29672 8652
rect 29608 8548 29672 8552
rect 29608 8492 29612 8548
rect 29612 8492 29668 8548
rect 29668 8492 29672 8548
rect 29608 8488 29672 8492
rect 29608 8388 29672 8392
rect 29608 8332 29612 8388
rect 29612 8332 29668 8388
rect 29668 8332 29672 8388
rect 29608 8328 29672 8332
rect 29608 8228 29672 8232
rect 29608 8172 29612 8228
rect 29612 8172 29668 8228
rect 29668 8172 29672 8228
rect 29608 8168 29672 8172
rect 29608 8068 29672 8072
rect 29608 8012 29612 8068
rect 29612 8012 29668 8068
rect 29668 8012 29672 8068
rect 29608 8008 29672 8012
rect 29608 7908 29672 7912
rect 29608 7852 29612 7908
rect 29612 7852 29668 7908
rect 29668 7852 29672 7908
rect 29608 7848 29672 7852
rect 29608 7748 29672 7752
rect 29608 7692 29612 7748
rect 29612 7692 29668 7748
rect 29668 7692 29672 7748
rect 29608 7688 29672 7692
rect 29608 7588 29672 7592
rect 29608 7532 29612 7588
rect 29612 7532 29668 7588
rect 29668 7532 29672 7588
rect 29608 7528 29672 7532
rect 29608 7428 29672 7432
rect 29608 7372 29612 7428
rect 29612 7372 29668 7428
rect 29668 7372 29672 7428
rect 29608 7368 29672 7372
rect 29608 7268 29672 7272
rect 29608 7212 29612 7268
rect 29612 7212 29668 7268
rect 29668 7212 29672 7268
rect 29608 7208 29672 7212
rect 29608 7108 29672 7112
rect 29608 7052 29612 7108
rect 29612 7052 29668 7108
rect 29668 7052 29672 7108
rect 29608 7048 29672 7052
rect 29608 6948 29672 6952
rect 29608 6892 29612 6948
rect 29612 6892 29668 6948
rect 29668 6892 29672 6948
rect 29608 6888 29672 6892
rect 29608 6788 29672 6792
rect 29608 6732 29612 6788
rect 29612 6732 29668 6788
rect 29668 6732 29672 6788
rect 29608 6728 29672 6732
rect 29608 6628 29672 6632
rect 29608 6572 29612 6628
rect 29612 6572 29668 6628
rect 29668 6572 29672 6628
rect 29608 6568 29672 6572
rect 29608 6468 29672 6472
rect 29608 6412 29612 6468
rect 29612 6412 29668 6468
rect 29668 6412 29672 6468
rect 29608 6408 29672 6412
rect 29608 6308 29672 6312
rect 29608 6252 29612 6308
rect 29612 6252 29668 6308
rect 29668 6252 29672 6308
rect 29608 6248 29672 6252
rect 29608 6148 29672 6152
rect 29608 6092 29612 6148
rect 29612 6092 29668 6148
rect 29668 6092 29672 6148
rect 29608 6088 29672 6092
rect 29608 5988 29672 5992
rect 29608 5932 29612 5988
rect 29612 5932 29668 5988
rect 29668 5932 29672 5988
rect 29608 5928 29672 5932
rect 29608 5828 29672 5832
rect 29608 5772 29612 5828
rect 29612 5772 29668 5828
rect 29668 5772 29672 5828
rect 29608 5768 29672 5772
rect 29608 5668 29672 5672
rect 29608 5612 29612 5668
rect 29612 5612 29668 5668
rect 29668 5612 29672 5668
rect 29608 5608 29672 5612
rect 29608 5508 29672 5512
rect 29608 5452 29612 5508
rect 29612 5452 29668 5508
rect 29668 5452 29672 5508
rect 29608 5448 29672 5452
rect 29608 5348 29672 5352
rect 29608 5292 29612 5348
rect 29612 5292 29668 5348
rect 29668 5292 29672 5348
rect 29608 5288 29672 5292
rect 29608 5188 29672 5192
rect 29608 5132 29612 5188
rect 29612 5132 29668 5188
rect 29668 5132 29672 5188
rect 29608 5128 29672 5132
rect 29608 5028 29672 5032
rect 29608 4972 29612 5028
rect 29612 4972 29668 5028
rect 29668 4972 29672 5028
rect 29608 4968 29672 4972
rect 29608 4868 29672 4872
rect 29608 4812 29612 4868
rect 29612 4812 29668 4868
rect 29668 4812 29672 4868
rect 29608 4808 29672 4812
rect 29608 4708 29672 4712
rect 29608 4652 29612 4708
rect 29612 4652 29668 4708
rect 29668 4652 29672 4708
rect 29608 4648 29672 4652
rect 29608 4548 29672 4552
rect 29608 4492 29612 4548
rect 29612 4492 29668 4548
rect 29668 4492 29672 4548
rect 29608 4488 29672 4492
rect 29608 4388 29672 4392
rect 29608 4332 29612 4388
rect 29612 4332 29668 4388
rect 29668 4332 29672 4388
rect 29608 4328 29672 4332
rect 29608 4228 29672 4232
rect 29608 4172 29612 4228
rect 29612 4172 29668 4228
rect 29668 4172 29672 4228
rect 29608 4168 29672 4172
rect 29608 4068 29672 4072
rect 29608 4012 29612 4068
rect 29612 4012 29668 4068
rect 29668 4012 29672 4068
rect 29608 4008 29672 4012
rect 29608 3908 29672 3912
rect 29608 3852 29612 3908
rect 29612 3852 29668 3908
rect 29668 3852 29672 3908
rect 29608 3848 29672 3852
rect 29608 3588 29672 3592
rect 29608 3532 29612 3588
rect 29612 3532 29668 3588
rect 29668 3532 29672 3588
rect 29608 3528 29672 3532
rect 29608 3428 29672 3432
rect 29608 3372 29612 3428
rect 29612 3372 29668 3428
rect 29668 3372 29672 3428
rect 29608 3368 29672 3372
rect 29608 3268 29672 3272
rect 29608 3212 29612 3268
rect 29612 3212 29668 3268
rect 29668 3212 29672 3268
rect 29608 3208 29672 3212
rect 29608 3108 29672 3112
rect 29608 3052 29612 3108
rect 29612 3052 29668 3108
rect 29668 3052 29672 3108
rect 29608 3048 29672 3052
rect 29608 2948 29672 2952
rect 29608 2892 29612 2948
rect 29612 2892 29668 2948
rect 29668 2892 29672 2948
rect 29608 2888 29672 2892
rect 29608 2788 29672 2792
rect 29608 2732 29612 2788
rect 29612 2732 29668 2788
rect 29668 2732 29672 2788
rect 29608 2728 29672 2732
rect 29608 2628 29672 2632
rect 29608 2572 29612 2628
rect 29612 2572 29668 2628
rect 29668 2572 29672 2628
rect 29608 2568 29672 2572
rect 29608 2468 29672 2472
rect 29608 2412 29612 2468
rect 29612 2412 29668 2468
rect 29668 2412 29672 2468
rect 29608 2408 29672 2412
rect 29608 2308 29672 2312
rect 29608 2252 29612 2308
rect 29612 2252 29668 2308
rect 29668 2252 29672 2308
rect 29608 2248 29672 2252
rect 29608 2148 29672 2152
rect 29608 2092 29612 2148
rect 29612 2092 29668 2148
rect 29668 2092 29672 2148
rect 29608 2088 29672 2092
rect 29608 1988 29672 1992
rect 29608 1932 29612 1988
rect 29612 1932 29668 1988
rect 29668 1932 29672 1988
rect 29608 1928 29672 1932
rect 29608 1828 29672 1832
rect 29608 1772 29612 1828
rect 29612 1772 29668 1828
rect 29668 1772 29672 1828
rect 29608 1768 29672 1772
rect 29608 1668 29672 1672
rect 29608 1612 29612 1668
rect 29612 1612 29668 1668
rect 29668 1612 29672 1668
rect 29608 1608 29672 1612
rect 29608 1508 29672 1512
rect 29608 1452 29612 1508
rect 29612 1452 29668 1508
rect 29668 1452 29672 1508
rect 29608 1448 29672 1452
rect 29608 1348 29672 1352
rect 29608 1292 29612 1348
rect 29612 1292 29668 1348
rect 29668 1292 29672 1348
rect 29608 1288 29672 1292
rect 29608 1188 29672 1192
rect 29608 1132 29612 1188
rect 29612 1132 29668 1188
rect 29668 1132 29672 1188
rect 29608 1128 29672 1132
rect 29608 1028 29672 1032
rect 29608 972 29612 1028
rect 29612 972 29668 1028
rect 29668 972 29672 1028
rect 29608 968 29672 972
rect 29288 808 29352 872
rect 29288 728 29352 792
rect 29288 648 29352 712
rect 29288 568 29352 632
rect 29288 488 29352 552
rect 29768 29128 29832 29192
rect 29768 23368 29832 23432
rect 29768 9448 29832 9512
rect 29768 3688 29832 3752
rect 29928 31908 29992 31912
rect 29928 31852 29932 31908
rect 29932 31852 29988 31908
rect 29988 31852 29992 31908
rect 29928 31848 29992 31852
rect 29928 31748 29992 31752
rect 29928 31692 29932 31748
rect 29932 31692 29988 31748
rect 29988 31692 29992 31748
rect 29928 31688 29992 31692
rect 29928 31588 29992 31592
rect 29928 31532 29932 31588
rect 29932 31532 29988 31588
rect 29988 31532 29992 31588
rect 29928 31528 29992 31532
rect 29928 31428 29992 31432
rect 29928 31372 29932 31428
rect 29932 31372 29988 31428
rect 29988 31372 29992 31428
rect 29928 31368 29992 31372
rect 29928 31268 29992 31272
rect 29928 31212 29932 31268
rect 29932 31212 29988 31268
rect 29988 31212 29992 31268
rect 29928 31208 29992 31212
rect 29928 31108 29992 31112
rect 29928 31052 29932 31108
rect 29932 31052 29988 31108
rect 29988 31052 29992 31108
rect 29928 31048 29992 31052
rect 29928 30948 29992 30952
rect 29928 30892 29932 30948
rect 29932 30892 29988 30948
rect 29988 30892 29992 30948
rect 29928 30888 29992 30892
rect 29928 30788 29992 30792
rect 29928 30732 29932 30788
rect 29932 30732 29988 30788
rect 29988 30732 29992 30788
rect 29928 30728 29992 30732
rect 29928 30628 29992 30632
rect 29928 30572 29932 30628
rect 29932 30572 29988 30628
rect 29988 30572 29992 30628
rect 29928 30568 29992 30572
rect 29928 30468 29992 30472
rect 29928 30412 29932 30468
rect 29932 30412 29988 30468
rect 29988 30412 29992 30468
rect 29928 30408 29992 30412
rect 29928 30308 29992 30312
rect 29928 30252 29932 30308
rect 29932 30252 29988 30308
rect 29988 30252 29992 30308
rect 29928 30248 29992 30252
rect 29928 30148 29992 30152
rect 29928 30092 29932 30148
rect 29932 30092 29988 30148
rect 29988 30092 29992 30148
rect 29928 30088 29992 30092
rect 29928 29988 29992 29992
rect 29928 29932 29932 29988
rect 29932 29932 29988 29988
rect 29988 29932 29992 29988
rect 29928 29928 29992 29932
rect 29928 29828 29992 29832
rect 29928 29772 29932 29828
rect 29932 29772 29988 29828
rect 29988 29772 29992 29828
rect 29928 29768 29992 29772
rect 29928 29668 29992 29672
rect 29928 29612 29932 29668
rect 29932 29612 29988 29668
rect 29988 29612 29992 29668
rect 29928 29608 29992 29612
rect 29928 29508 29992 29512
rect 29928 29452 29932 29508
rect 29932 29452 29988 29508
rect 29988 29452 29992 29508
rect 29928 29448 29992 29452
rect 29928 29348 29992 29352
rect 29928 29292 29932 29348
rect 29932 29292 29988 29348
rect 29988 29292 29992 29348
rect 29928 29288 29992 29292
rect 29928 29028 29992 29032
rect 29928 28972 29932 29028
rect 29932 28972 29988 29028
rect 29988 28972 29992 29028
rect 29928 28968 29992 28972
rect 29928 28868 29992 28872
rect 29928 28812 29932 28868
rect 29932 28812 29988 28868
rect 29988 28812 29992 28868
rect 29928 28808 29992 28812
rect 29928 28708 29992 28712
rect 29928 28652 29932 28708
rect 29932 28652 29988 28708
rect 29988 28652 29992 28708
rect 29928 28648 29992 28652
rect 29928 28548 29992 28552
rect 29928 28492 29932 28548
rect 29932 28492 29988 28548
rect 29988 28492 29992 28548
rect 29928 28488 29992 28492
rect 29928 28388 29992 28392
rect 29928 28332 29932 28388
rect 29932 28332 29988 28388
rect 29988 28332 29992 28388
rect 29928 28328 29992 28332
rect 29928 28228 29992 28232
rect 29928 28172 29932 28228
rect 29932 28172 29988 28228
rect 29988 28172 29992 28228
rect 29928 28168 29992 28172
rect 29928 28068 29992 28072
rect 29928 28012 29932 28068
rect 29932 28012 29988 28068
rect 29988 28012 29992 28068
rect 29928 28008 29992 28012
rect 29928 27908 29992 27912
rect 29928 27852 29932 27908
rect 29932 27852 29988 27908
rect 29988 27852 29992 27908
rect 29928 27848 29992 27852
rect 29928 27748 29992 27752
rect 29928 27692 29932 27748
rect 29932 27692 29988 27748
rect 29988 27692 29992 27748
rect 29928 27688 29992 27692
rect 29928 27588 29992 27592
rect 29928 27532 29932 27588
rect 29932 27532 29988 27588
rect 29988 27532 29992 27588
rect 29928 27528 29992 27532
rect 29928 27428 29992 27432
rect 29928 27372 29932 27428
rect 29932 27372 29988 27428
rect 29988 27372 29992 27428
rect 29928 27368 29992 27372
rect 29928 27268 29992 27272
rect 29928 27212 29932 27268
rect 29932 27212 29988 27268
rect 29988 27212 29992 27268
rect 29928 27208 29992 27212
rect 29928 27108 29992 27112
rect 29928 27052 29932 27108
rect 29932 27052 29988 27108
rect 29988 27052 29992 27108
rect 29928 27048 29992 27052
rect 29928 26948 29992 26952
rect 29928 26892 29932 26948
rect 29932 26892 29988 26948
rect 29988 26892 29992 26948
rect 29928 26888 29992 26892
rect 29928 26788 29992 26792
rect 29928 26732 29932 26788
rect 29932 26732 29988 26788
rect 29988 26732 29992 26788
rect 29928 26728 29992 26732
rect 29928 26628 29992 26632
rect 29928 26572 29932 26628
rect 29932 26572 29988 26628
rect 29988 26572 29992 26628
rect 29928 26568 29992 26572
rect 29928 26468 29992 26472
rect 29928 26412 29932 26468
rect 29932 26412 29988 26468
rect 29988 26412 29992 26468
rect 29928 26408 29992 26412
rect 29928 26308 29992 26312
rect 29928 26252 29932 26308
rect 29932 26252 29988 26308
rect 29988 26252 29992 26308
rect 29928 26248 29992 26252
rect 29928 26148 29992 26152
rect 29928 26092 29932 26148
rect 29932 26092 29988 26148
rect 29988 26092 29992 26148
rect 29928 26088 29992 26092
rect 29928 25988 29992 25992
rect 29928 25932 29932 25988
rect 29932 25932 29988 25988
rect 29988 25932 29992 25988
rect 29928 25928 29992 25932
rect 29928 25828 29992 25832
rect 29928 25772 29932 25828
rect 29932 25772 29988 25828
rect 29988 25772 29992 25828
rect 29928 25768 29992 25772
rect 29928 25668 29992 25672
rect 29928 25612 29932 25668
rect 29932 25612 29988 25668
rect 29988 25612 29992 25668
rect 29928 25608 29992 25612
rect 29928 25508 29992 25512
rect 29928 25452 29932 25508
rect 29932 25452 29988 25508
rect 29988 25452 29992 25508
rect 29928 25448 29992 25452
rect 29928 25348 29992 25352
rect 29928 25292 29932 25348
rect 29932 25292 29988 25348
rect 29988 25292 29992 25348
rect 29928 25288 29992 25292
rect 29928 25188 29992 25192
rect 29928 25132 29932 25188
rect 29932 25132 29988 25188
rect 29988 25132 29992 25188
rect 29928 25128 29992 25132
rect 29928 25028 29992 25032
rect 29928 24972 29932 25028
rect 29932 24972 29988 25028
rect 29988 24972 29992 25028
rect 29928 24968 29992 24972
rect 29928 24868 29992 24872
rect 29928 24812 29932 24868
rect 29932 24812 29988 24868
rect 29988 24812 29992 24868
rect 29928 24808 29992 24812
rect 29928 24708 29992 24712
rect 29928 24652 29932 24708
rect 29932 24652 29988 24708
rect 29988 24652 29992 24708
rect 29928 24648 29992 24652
rect 29928 24548 29992 24552
rect 29928 24492 29932 24548
rect 29932 24492 29988 24548
rect 29988 24492 29992 24548
rect 29928 24488 29992 24492
rect 29928 24388 29992 24392
rect 29928 24332 29932 24388
rect 29932 24332 29988 24388
rect 29988 24332 29992 24388
rect 29928 24328 29992 24332
rect 29928 24228 29992 24232
rect 29928 24172 29932 24228
rect 29932 24172 29988 24228
rect 29988 24172 29992 24228
rect 29928 24168 29992 24172
rect 29928 24068 29992 24072
rect 29928 24012 29932 24068
rect 29932 24012 29988 24068
rect 29988 24012 29992 24068
rect 29928 24008 29992 24012
rect 29928 23908 29992 23912
rect 29928 23852 29932 23908
rect 29932 23852 29988 23908
rect 29988 23852 29992 23908
rect 29928 23848 29992 23852
rect 29928 23748 29992 23752
rect 29928 23692 29932 23748
rect 29932 23692 29988 23748
rect 29988 23692 29992 23748
rect 29928 23688 29992 23692
rect 29928 23588 29992 23592
rect 29928 23532 29932 23588
rect 29932 23532 29988 23588
rect 29988 23532 29992 23588
rect 29928 23528 29992 23532
rect 29928 23268 29992 23272
rect 29928 23212 29932 23268
rect 29932 23212 29988 23268
rect 29988 23212 29992 23268
rect 29928 23208 29992 23212
rect 29928 23108 29992 23112
rect 29928 23052 29932 23108
rect 29932 23052 29988 23108
rect 29988 23052 29992 23108
rect 29928 23048 29992 23052
rect 29928 22948 29992 22952
rect 29928 22892 29932 22948
rect 29932 22892 29988 22948
rect 29988 22892 29992 22948
rect 29928 22888 29992 22892
rect 29928 22788 29992 22792
rect 29928 22732 29932 22788
rect 29932 22732 29988 22788
rect 29988 22732 29992 22788
rect 29928 22728 29992 22732
rect 29928 22628 29992 22632
rect 29928 22572 29932 22628
rect 29932 22572 29988 22628
rect 29988 22572 29992 22628
rect 29928 22568 29992 22572
rect 29928 22468 29992 22472
rect 29928 22412 29932 22468
rect 29932 22412 29988 22468
rect 29988 22412 29992 22468
rect 29928 22408 29992 22412
rect 29928 22308 29992 22312
rect 29928 22252 29932 22308
rect 29932 22252 29988 22308
rect 29988 22252 29992 22308
rect 29928 22248 29992 22252
rect 29928 22148 29992 22152
rect 29928 22092 29932 22148
rect 29932 22092 29988 22148
rect 29988 22092 29992 22148
rect 29928 22088 29992 22092
rect 29928 21988 29992 21992
rect 29928 21932 29932 21988
rect 29932 21932 29988 21988
rect 29988 21932 29992 21988
rect 29928 21928 29992 21932
rect 29928 21828 29992 21832
rect 29928 21772 29932 21828
rect 29932 21772 29988 21828
rect 29988 21772 29992 21828
rect 29928 21768 29992 21772
rect 29928 21668 29992 21672
rect 29928 21612 29932 21668
rect 29932 21612 29988 21668
rect 29988 21612 29992 21668
rect 29928 21608 29992 21612
rect 29928 21508 29992 21512
rect 29928 21452 29932 21508
rect 29932 21452 29988 21508
rect 29988 21452 29992 21508
rect 29928 21448 29992 21452
rect 29928 21348 29992 21352
rect 29928 21292 29932 21348
rect 29932 21292 29988 21348
rect 29988 21292 29992 21348
rect 29928 21288 29992 21292
rect 29928 21188 29992 21192
rect 29928 21132 29932 21188
rect 29932 21132 29988 21188
rect 29988 21132 29992 21188
rect 29928 21128 29992 21132
rect 29928 21028 29992 21032
rect 29928 20972 29932 21028
rect 29932 20972 29988 21028
rect 29988 20972 29992 21028
rect 29928 20968 29992 20972
rect 29928 20868 29992 20872
rect 29928 20812 29932 20868
rect 29932 20812 29988 20868
rect 29988 20812 29992 20868
rect 29928 20808 29992 20812
rect 29928 20708 29992 20712
rect 29928 20652 29932 20708
rect 29932 20652 29988 20708
rect 29988 20652 29992 20708
rect 29928 20648 29992 20652
rect 29928 20548 29992 20552
rect 29928 20492 29932 20548
rect 29932 20492 29988 20548
rect 29988 20492 29992 20548
rect 29928 20488 29992 20492
rect 29928 20388 29992 20392
rect 29928 20332 29932 20388
rect 29932 20332 29988 20388
rect 29988 20332 29992 20388
rect 29928 20328 29992 20332
rect 29928 20228 29992 20232
rect 29928 20172 29932 20228
rect 29932 20172 29988 20228
rect 29988 20172 29992 20228
rect 29928 20168 29992 20172
rect 29928 20068 29992 20072
rect 29928 20012 29932 20068
rect 29932 20012 29988 20068
rect 29988 20012 29992 20068
rect 29928 20008 29992 20012
rect 29928 19908 29992 19912
rect 29928 19852 29932 19908
rect 29932 19852 29988 19908
rect 29988 19852 29992 19908
rect 29928 19848 29992 19852
rect 29928 19748 29992 19752
rect 29928 19692 29932 19748
rect 29932 19692 29988 19748
rect 29988 19692 29992 19748
rect 29928 19688 29992 19692
rect 29928 19588 29992 19592
rect 29928 19532 29932 19588
rect 29932 19532 29988 19588
rect 29988 19532 29992 19588
rect 29928 19528 29992 19532
rect 29928 19428 29992 19432
rect 29928 19372 29932 19428
rect 29932 19372 29988 19428
rect 29988 19372 29992 19428
rect 29928 19368 29992 19372
rect 29928 19268 29992 19272
rect 29928 19212 29932 19268
rect 29932 19212 29988 19268
rect 29988 19212 29992 19268
rect 29928 19208 29992 19212
rect 29928 19108 29992 19112
rect 29928 19052 29932 19108
rect 29932 19052 29988 19108
rect 29988 19052 29992 19108
rect 29928 19048 29992 19052
rect 29928 18948 29992 18952
rect 29928 18892 29932 18948
rect 29932 18892 29988 18948
rect 29988 18892 29992 18948
rect 29928 18888 29992 18892
rect 29928 18788 29992 18792
rect 29928 18732 29932 18788
rect 29932 18732 29988 18788
rect 29988 18732 29992 18788
rect 29928 18728 29992 18732
rect 29928 18628 29992 18632
rect 29928 18572 29932 18628
rect 29932 18572 29988 18628
rect 29988 18572 29992 18628
rect 29928 18568 29992 18572
rect 29928 18468 29992 18472
rect 29928 18412 29932 18468
rect 29932 18412 29988 18468
rect 29988 18412 29992 18468
rect 29928 18408 29992 18412
rect 29928 18308 29992 18312
rect 29928 18252 29932 18308
rect 29932 18252 29988 18308
rect 29988 18252 29992 18308
rect 29928 18248 29992 18252
rect 29928 18148 29992 18152
rect 29928 18092 29932 18148
rect 29932 18092 29988 18148
rect 29988 18092 29992 18148
rect 29928 18088 29992 18092
rect 29928 17988 29992 17992
rect 29928 17932 29932 17988
rect 29932 17932 29988 17988
rect 29988 17932 29992 17988
rect 29928 17928 29992 17932
rect 29928 17828 29992 17832
rect 29928 17772 29932 17828
rect 29932 17772 29988 17828
rect 29988 17772 29992 17828
rect 29928 17768 29992 17772
rect 29928 17668 29992 17672
rect 29928 17612 29932 17668
rect 29932 17612 29988 17668
rect 29988 17612 29992 17668
rect 29928 17608 29992 17612
rect 29928 17508 29992 17512
rect 29928 17452 29932 17508
rect 29932 17452 29988 17508
rect 29988 17452 29992 17508
rect 29928 17448 29992 17452
rect 29928 17348 29992 17352
rect 29928 17292 29932 17348
rect 29932 17292 29988 17348
rect 29988 17292 29992 17348
rect 29928 17288 29992 17292
rect 29928 17188 29992 17192
rect 29928 17132 29932 17188
rect 29932 17132 29988 17188
rect 29988 17132 29992 17188
rect 29928 17128 29992 17132
rect 29928 17028 29992 17032
rect 29928 16972 29932 17028
rect 29932 16972 29988 17028
rect 29988 16972 29992 17028
rect 29928 16968 29992 16972
rect 29928 16868 29992 16872
rect 29928 16812 29932 16868
rect 29932 16812 29988 16868
rect 29988 16812 29992 16868
rect 29928 16808 29992 16812
rect 29928 16708 29992 16712
rect 29928 16652 29932 16708
rect 29932 16652 29988 16708
rect 29988 16652 29992 16708
rect 29928 16648 29992 16652
rect 29928 16548 29992 16552
rect 29928 16492 29932 16548
rect 29932 16492 29988 16548
rect 29988 16492 29992 16548
rect 29928 16488 29992 16492
rect 29928 16388 29992 16392
rect 29928 16332 29932 16388
rect 29932 16332 29988 16388
rect 29988 16332 29992 16388
rect 29928 16328 29992 16332
rect 29928 16228 29992 16232
rect 29928 16172 29932 16228
rect 29932 16172 29988 16228
rect 29988 16172 29992 16228
rect 29928 16168 29992 16172
rect 29928 16068 29992 16072
rect 29928 16012 29932 16068
rect 29932 16012 29988 16068
rect 29988 16012 29992 16068
rect 29928 16008 29992 16012
rect 29928 15908 29992 15912
rect 29928 15852 29932 15908
rect 29932 15852 29988 15908
rect 29988 15852 29992 15908
rect 29928 15848 29992 15852
rect 29928 15748 29992 15752
rect 29928 15692 29932 15748
rect 29932 15692 29988 15748
rect 29988 15692 29992 15748
rect 29928 15688 29992 15692
rect 29928 15588 29992 15592
rect 29928 15532 29932 15588
rect 29932 15532 29988 15588
rect 29988 15532 29992 15588
rect 29928 15528 29992 15532
rect 29928 15428 29992 15432
rect 29928 15372 29932 15428
rect 29932 15372 29988 15428
rect 29988 15372 29992 15428
rect 29928 15368 29992 15372
rect 29928 15268 29992 15272
rect 29928 15212 29932 15268
rect 29932 15212 29988 15268
rect 29988 15212 29992 15268
rect 29928 15208 29992 15212
rect 29928 15108 29992 15112
rect 29928 15052 29932 15108
rect 29932 15052 29988 15108
rect 29988 15052 29992 15108
rect 29928 15048 29992 15052
rect 29928 14948 29992 14952
rect 29928 14892 29932 14948
rect 29932 14892 29988 14948
rect 29988 14892 29992 14948
rect 29928 14888 29992 14892
rect 29928 14788 29992 14792
rect 29928 14732 29932 14788
rect 29932 14732 29988 14788
rect 29988 14732 29992 14788
rect 29928 14728 29992 14732
rect 29928 14628 29992 14632
rect 29928 14572 29932 14628
rect 29932 14572 29988 14628
rect 29988 14572 29992 14628
rect 29928 14568 29992 14572
rect 29928 14468 29992 14472
rect 29928 14412 29932 14468
rect 29932 14412 29988 14468
rect 29988 14412 29992 14468
rect 29928 14408 29992 14412
rect 29928 14308 29992 14312
rect 29928 14252 29932 14308
rect 29932 14252 29988 14308
rect 29988 14252 29992 14308
rect 29928 14248 29992 14252
rect 29928 14148 29992 14152
rect 29928 14092 29932 14148
rect 29932 14092 29988 14148
rect 29988 14092 29992 14148
rect 29928 14088 29992 14092
rect 29928 13988 29992 13992
rect 29928 13932 29932 13988
rect 29932 13932 29988 13988
rect 29988 13932 29992 13988
rect 29928 13928 29992 13932
rect 29928 13828 29992 13832
rect 29928 13772 29932 13828
rect 29932 13772 29988 13828
rect 29988 13772 29992 13828
rect 29928 13768 29992 13772
rect 29928 13668 29992 13672
rect 29928 13612 29932 13668
rect 29932 13612 29988 13668
rect 29988 13612 29992 13668
rect 29928 13608 29992 13612
rect 29928 13508 29992 13512
rect 29928 13452 29932 13508
rect 29932 13452 29988 13508
rect 29988 13452 29992 13508
rect 29928 13448 29992 13452
rect 29928 13348 29992 13352
rect 29928 13292 29932 13348
rect 29932 13292 29988 13348
rect 29988 13292 29992 13348
rect 29928 13288 29992 13292
rect 29928 13188 29992 13192
rect 29928 13132 29932 13188
rect 29932 13132 29988 13188
rect 29988 13132 29992 13188
rect 29928 13128 29992 13132
rect 29928 13028 29992 13032
rect 29928 12972 29932 13028
rect 29932 12972 29988 13028
rect 29988 12972 29992 13028
rect 29928 12968 29992 12972
rect 29928 12868 29992 12872
rect 29928 12812 29932 12868
rect 29932 12812 29988 12868
rect 29988 12812 29992 12868
rect 29928 12808 29992 12812
rect 29928 12708 29992 12712
rect 29928 12652 29932 12708
rect 29932 12652 29988 12708
rect 29988 12652 29992 12708
rect 29928 12648 29992 12652
rect 29928 12548 29992 12552
rect 29928 12492 29932 12548
rect 29932 12492 29988 12548
rect 29988 12492 29992 12548
rect 29928 12488 29992 12492
rect 29928 12388 29992 12392
rect 29928 12332 29932 12388
rect 29932 12332 29988 12388
rect 29988 12332 29992 12388
rect 29928 12328 29992 12332
rect 29928 12228 29992 12232
rect 29928 12172 29932 12228
rect 29932 12172 29988 12228
rect 29988 12172 29992 12228
rect 29928 12168 29992 12172
rect 29928 12068 29992 12072
rect 29928 12012 29932 12068
rect 29932 12012 29988 12068
rect 29988 12012 29992 12068
rect 29928 12008 29992 12012
rect 29928 11908 29992 11912
rect 29928 11852 29932 11908
rect 29932 11852 29988 11908
rect 29988 11852 29992 11908
rect 29928 11848 29992 11852
rect 29928 11748 29992 11752
rect 29928 11692 29932 11748
rect 29932 11692 29988 11748
rect 29988 11692 29992 11748
rect 29928 11688 29992 11692
rect 29928 11588 29992 11592
rect 29928 11532 29932 11588
rect 29932 11532 29988 11588
rect 29988 11532 29992 11588
rect 29928 11528 29992 11532
rect 29928 11428 29992 11432
rect 29928 11372 29932 11428
rect 29932 11372 29988 11428
rect 29988 11372 29992 11428
rect 29928 11368 29992 11372
rect 29928 11268 29992 11272
rect 29928 11212 29932 11268
rect 29932 11212 29988 11268
rect 29988 11212 29992 11268
rect 29928 11208 29992 11212
rect 29928 11108 29992 11112
rect 29928 11052 29932 11108
rect 29932 11052 29988 11108
rect 29988 11052 29992 11108
rect 29928 11048 29992 11052
rect 29928 10948 29992 10952
rect 29928 10892 29932 10948
rect 29932 10892 29988 10948
rect 29988 10892 29992 10948
rect 29928 10888 29992 10892
rect 29928 10788 29992 10792
rect 29928 10732 29932 10788
rect 29932 10732 29988 10788
rect 29988 10732 29992 10788
rect 29928 10728 29992 10732
rect 29928 10628 29992 10632
rect 29928 10572 29932 10628
rect 29932 10572 29988 10628
rect 29988 10572 29992 10628
rect 29928 10568 29992 10572
rect 29928 10468 29992 10472
rect 29928 10412 29932 10468
rect 29932 10412 29988 10468
rect 29988 10412 29992 10468
rect 29928 10408 29992 10412
rect 29928 10308 29992 10312
rect 29928 10252 29932 10308
rect 29932 10252 29988 10308
rect 29988 10252 29992 10308
rect 29928 10248 29992 10252
rect 29928 10148 29992 10152
rect 29928 10092 29932 10148
rect 29932 10092 29988 10148
rect 29988 10092 29992 10148
rect 29928 10088 29992 10092
rect 29928 9988 29992 9992
rect 29928 9932 29932 9988
rect 29932 9932 29988 9988
rect 29988 9932 29992 9988
rect 29928 9928 29992 9932
rect 29928 9828 29992 9832
rect 29928 9772 29932 9828
rect 29932 9772 29988 9828
rect 29988 9772 29992 9828
rect 29928 9768 29992 9772
rect 29928 9668 29992 9672
rect 29928 9612 29932 9668
rect 29932 9612 29988 9668
rect 29988 9612 29992 9668
rect 29928 9608 29992 9612
rect 29928 9348 29992 9352
rect 29928 9292 29932 9348
rect 29932 9292 29988 9348
rect 29988 9292 29992 9348
rect 29928 9288 29992 9292
rect 29928 9188 29992 9192
rect 29928 9132 29932 9188
rect 29932 9132 29988 9188
rect 29988 9132 29992 9188
rect 29928 9128 29992 9132
rect 29928 9028 29992 9032
rect 29928 8972 29932 9028
rect 29932 8972 29988 9028
rect 29988 8972 29992 9028
rect 29928 8968 29992 8972
rect 29928 8868 29992 8872
rect 29928 8812 29932 8868
rect 29932 8812 29988 8868
rect 29988 8812 29992 8868
rect 29928 8808 29992 8812
rect 29928 8708 29992 8712
rect 29928 8652 29932 8708
rect 29932 8652 29988 8708
rect 29988 8652 29992 8708
rect 29928 8648 29992 8652
rect 29928 8548 29992 8552
rect 29928 8492 29932 8548
rect 29932 8492 29988 8548
rect 29988 8492 29992 8548
rect 29928 8488 29992 8492
rect 29928 8388 29992 8392
rect 29928 8332 29932 8388
rect 29932 8332 29988 8388
rect 29988 8332 29992 8388
rect 29928 8328 29992 8332
rect 29928 8228 29992 8232
rect 29928 8172 29932 8228
rect 29932 8172 29988 8228
rect 29988 8172 29992 8228
rect 29928 8168 29992 8172
rect 29928 8068 29992 8072
rect 29928 8012 29932 8068
rect 29932 8012 29988 8068
rect 29988 8012 29992 8068
rect 29928 8008 29992 8012
rect 29928 7908 29992 7912
rect 29928 7852 29932 7908
rect 29932 7852 29988 7908
rect 29988 7852 29992 7908
rect 29928 7848 29992 7852
rect 29928 7748 29992 7752
rect 29928 7692 29932 7748
rect 29932 7692 29988 7748
rect 29988 7692 29992 7748
rect 29928 7688 29992 7692
rect 29928 7588 29992 7592
rect 29928 7532 29932 7588
rect 29932 7532 29988 7588
rect 29988 7532 29992 7588
rect 29928 7528 29992 7532
rect 29928 7428 29992 7432
rect 29928 7372 29932 7428
rect 29932 7372 29988 7428
rect 29988 7372 29992 7428
rect 29928 7368 29992 7372
rect 29928 7268 29992 7272
rect 29928 7212 29932 7268
rect 29932 7212 29988 7268
rect 29988 7212 29992 7268
rect 29928 7208 29992 7212
rect 29928 7108 29992 7112
rect 29928 7052 29932 7108
rect 29932 7052 29988 7108
rect 29988 7052 29992 7108
rect 29928 7048 29992 7052
rect 29928 6948 29992 6952
rect 29928 6892 29932 6948
rect 29932 6892 29988 6948
rect 29988 6892 29992 6948
rect 29928 6888 29992 6892
rect 29928 6788 29992 6792
rect 29928 6732 29932 6788
rect 29932 6732 29988 6788
rect 29988 6732 29992 6788
rect 29928 6728 29992 6732
rect 29928 6628 29992 6632
rect 29928 6572 29932 6628
rect 29932 6572 29988 6628
rect 29988 6572 29992 6628
rect 29928 6568 29992 6572
rect 29928 6468 29992 6472
rect 29928 6412 29932 6468
rect 29932 6412 29988 6468
rect 29988 6412 29992 6468
rect 29928 6408 29992 6412
rect 29928 6308 29992 6312
rect 29928 6252 29932 6308
rect 29932 6252 29988 6308
rect 29988 6252 29992 6308
rect 29928 6248 29992 6252
rect 29928 6148 29992 6152
rect 29928 6092 29932 6148
rect 29932 6092 29988 6148
rect 29988 6092 29992 6148
rect 29928 6088 29992 6092
rect 29928 5988 29992 5992
rect 29928 5932 29932 5988
rect 29932 5932 29988 5988
rect 29988 5932 29992 5988
rect 29928 5928 29992 5932
rect 29928 5828 29992 5832
rect 29928 5772 29932 5828
rect 29932 5772 29988 5828
rect 29988 5772 29992 5828
rect 29928 5768 29992 5772
rect 29928 5668 29992 5672
rect 29928 5612 29932 5668
rect 29932 5612 29988 5668
rect 29988 5612 29992 5668
rect 29928 5608 29992 5612
rect 29928 5508 29992 5512
rect 29928 5452 29932 5508
rect 29932 5452 29988 5508
rect 29988 5452 29992 5508
rect 29928 5448 29992 5452
rect 29928 5348 29992 5352
rect 29928 5292 29932 5348
rect 29932 5292 29988 5348
rect 29988 5292 29992 5348
rect 29928 5288 29992 5292
rect 29928 5188 29992 5192
rect 29928 5132 29932 5188
rect 29932 5132 29988 5188
rect 29988 5132 29992 5188
rect 29928 5128 29992 5132
rect 29928 5028 29992 5032
rect 29928 4972 29932 5028
rect 29932 4972 29988 5028
rect 29988 4972 29992 5028
rect 29928 4968 29992 4972
rect 29928 4868 29992 4872
rect 29928 4812 29932 4868
rect 29932 4812 29988 4868
rect 29988 4812 29992 4868
rect 29928 4808 29992 4812
rect 29928 4708 29992 4712
rect 29928 4652 29932 4708
rect 29932 4652 29988 4708
rect 29988 4652 29992 4708
rect 29928 4648 29992 4652
rect 29928 4548 29992 4552
rect 29928 4492 29932 4548
rect 29932 4492 29988 4548
rect 29988 4492 29992 4548
rect 29928 4488 29992 4492
rect 29928 4388 29992 4392
rect 29928 4332 29932 4388
rect 29932 4332 29988 4388
rect 29988 4332 29992 4388
rect 29928 4328 29992 4332
rect 29928 4228 29992 4232
rect 29928 4172 29932 4228
rect 29932 4172 29988 4228
rect 29988 4172 29992 4228
rect 29928 4168 29992 4172
rect 29928 4068 29992 4072
rect 29928 4012 29932 4068
rect 29932 4012 29988 4068
rect 29988 4012 29992 4068
rect 29928 4008 29992 4012
rect 29928 3908 29992 3912
rect 29928 3852 29932 3908
rect 29932 3852 29988 3908
rect 29988 3852 29992 3908
rect 29928 3848 29992 3852
rect 29928 3588 29992 3592
rect 29928 3532 29932 3588
rect 29932 3532 29988 3588
rect 29988 3532 29992 3588
rect 29928 3528 29992 3532
rect 29928 3428 29992 3432
rect 29928 3372 29932 3428
rect 29932 3372 29988 3428
rect 29988 3372 29992 3428
rect 29928 3368 29992 3372
rect 29928 3268 29992 3272
rect 29928 3212 29932 3268
rect 29932 3212 29988 3268
rect 29988 3212 29992 3268
rect 29928 3208 29992 3212
rect 29928 3108 29992 3112
rect 29928 3052 29932 3108
rect 29932 3052 29988 3108
rect 29988 3052 29992 3108
rect 29928 3048 29992 3052
rect 29928 2948 29992 2952
rect 29928 2892 29932 2948
rect 29932 2892 29988 2948
rect 29988 2892 29992 2948
rect 29928 2888 29992 2892
rect 29928 2788 29992 2792
rect 29928 2732 29932 2788
rect 29932 2732 29988 2788
rect 29988 2732 29992 2788
rect 29928 2728 29992 2732
rect 29928 2628 29992 2632
rect 29928 2572 29932 2628
rect 29932 2572 29988 2628
rect 29988 2572 29992 2628
rect 29928 2568 29992 2572
rect 29928 2468 29992 2472
rect 29928 2412 29932 2468
rect 29932 2412 29988 2468
rect 29988 2412 29992 2468
rect 29928 2408 29992 2412
rect 29928 2308 29992 2312
rect 29928 2252 29932 2308
rect 29932 2252 29988 2308
rect 29988 2252 29992 2308
rect 29928 2248 29992 2252
rect 29928 2148 29992 2152
rect 29928 2092 29932 2148
rect 29932 2092 29988 2148
rect 29988 2092 29992 2148
rect 29928 2088 29992 2092
rect 29928 1988 29992 1992
rect 29928 1932 29932 1988
rect 29932 1932 29988 1988
rect 29988 1932 29992 1988
rect 29928 1928 29992 1932
rect 29928 1828 29992 1832
rect 29928 1772 29932 1828
rect 29932 1772 29988 1828
rect 29988 1772 29992 1828
rect 29928 1768 29992 1772
rect 29928 1668 29992 1672
rect 29928 1612 29932 1668
rect 29932 1612 29988 1668
rect 29988 1612 29992 1668
rect 29928 1608 29992 1612
rect 29928 1508 29992 1512
rect 29928 1452 29932 1508
rect 29932 1452 29988 1508
rect 29988 1452 29992 1508
rect 29928 1448 29992 1452
rect 29928 1348 29992 1352
rect 29928 1292 29932 1348
rect 29932 1292 29988 1348
rect 29988 1292 29992 1348
rect 29928 1288 29992 1292
rect 29928 1188 29992 1192
rect 29928 1132 29932 1188
rect 29932 1132 29988 1188
rect 29988 1132 29992 1188
rect 29928 1128 29992 1132
rect 29928 1028 29992 1032
rect 29928 972 29932 1028
rect 29932 972 29988 1028
rect 29988 972 29992 1028
rect 29928 968 29992 972
rect 29608 808 29672 872
rect 29608 728 29672 792
rect 29608 648 29672 712
rect 29608 568 29672 632
rect 29608 488 29672 552
rect 29928 808 29992 872
rect 29928 728 29992 792
rect 29928 648 29992 712
rect 29928 568 29992 632
rect 29928 488 29992 552
rect 28808 328 28872 392
rect 28808 248 28872 312
rect 28808 168 28872 232
rect 28808 88 28872 152
rect 28808 8 28872 72
<< metal4 >>
rect 0 31912 1040 31920
rect 0 31848 8 31912
rect 72 31848 328 31912
rect 392 31848 648 31912
rect 712 31848 968 31912
rect 1032 31848 1040 31912
rect 0 31840 1040 31848
rect 28960 31912 30000 31920
rect 28960 31848 28968 31912
rect 29032 31848 29288 31912
rect 29352 31848 29608 31912
rect 29672 31848 29928 31912
rect 29992 31848 30000 31912
rect 28960 31840 30000 31848
rect 0 31752 1360 31760
rect 0 31688 8 31752
rect 72 31688 328 31752
rect 392 31688 648 31752
rect 712 31688 968 31752
rect 1032 31688 1360 31752
rect 0 31680 1360 31688
rect 28640 31752 30000 31760
rect 28640 31688 28968 31752
rect 29032 31688 29288 31752
rect 29352 31688 29608 31752
rect 29672 31688 29928 31752
rect 29992 31688 30000 31752
rect 28640 31680 30000 31688
rect 0 31592 1360 31600
rect 0 31528 8 31592
rect 72 31528 328 31592
rect 392 31528 648 31592
rect 712 31528 968 31592
rect 1032 31528 1360 31592
rect 0 31520 1360 31528
rect 28640 31592 30000 31600
rect 28640 31528 28968 31592
rect 29032 31528 29288 31592
rect 29352 31528 29608 31592
rect 29672 31528 29928 31592
rect 29992 31528 30000 31592
rect 28640 31520 30000 31528
rect 0 31432 1360 31440
rect 0 31368 8 31432
rect 72 31368 328 31432
rect 392 31368 648 31432
rect 712 31368 968 31432
rect 1032 31368 1360 31432
rect 0 31360 1360 31368
rect 28640 31432 30000 31440
rect 28640 31368 28968 31432
rect 29032 31368 29288 31432
rect 29352 31368 29608 31432
rect 29672 31368 29928 31432
rect 29992 31368 30000 31432
rect 28640 31360 30000 31368
rect 0 31272 1360 31280
rect 0 31208 8 31272
rect 72 31208 328 31272
rect 392 31208 648 31272
rect 712 31208 968 31272
rect 1032 31208 1360 31272
rect 0 31200 1360 31208
rect 28640 31272 30000 31280
rect 28640 31208 28968 31272
rect 29032 31208 29288 31272
rect 29352 31208 29608 31272
rect 29672 31208 29928 31272
rect 29992 31208 30000 31272
rect 28640 31200 30000 31208
rect 0 31112 1360 31120
rect 0 31048 8 31112
rect 72 31048 328 31112
rect 392 31048 648 31112
rect 712 31048 968 31112
rect 1032 31048 1360 31112
rect 0 31040 1360 31048
rect 28640 31112 30000 31120
rect 28640 31048 28968 31112
rect 29032 31048 29288 31112
rect 29352 31048 29608 31112
rect 29672 31048 29928 31112
rect 29992 31048 30000 31112
rect 28640 31040 30000 31048
rect 0 30952 1040 30960
rect 0 30888 8 30952
rect 72 30888 328 30952
rect 392 30888 648 30952
rect 712 30888 968 30952
rect 1032 30888 1040 30952
rect 0 30880 1040 30888
rect 28960 30952 30000 30960
rect 28960 30888 28968 30952
rect 29032 30888 29288 30952
rect 29352 30888 29608 30952
rect 29672 30888 29928 30952
rect 29992 30888 30000 30952
rect 28960 30880 30000 30888
rect 0 30792 1040 30800
rect 0 30728 8 30792
rect 72 30728 328 30792
rect 392 30728 648 30792
rect 712 30728 968 30792
rect 1032 30728 1040 30792
rect 0 30720 1040 30728
rect 28960 30792 30000 30800
rect 28960 30728 28968 30792
rect 29032 30728 29288 30792
rect 29352 30728 29608 30792
rect 29672 30728 29928 30792
rect 29992 30728 30000 30792
rect 28960 30720 30000 30728
rect 0 30632 1040 30640
rect 0 30568 8 30632
rect 72 30568 328 30632
rect 392 30568 648 30632
rect 712 30568 968 30632
rect 1032 30568 1040 30632
rect 0 30560 1040 30568
rect 28960 30632 30000 30640
rect 28960 30568 28968 30632
rect 29032 30568 29288 30632
rect 29352 30568 29608 30632
rect 29672 30568 29928 30632
rect 29992 30568 30000 30632
rect 28960 30560 30000 30568
rect 0 30472 1360 30480
rect 0 30408 8 30472
rect 72 30408 328 30472
rect 392 30408 648 30472
rect 712 30408 968 30472
rect 1032 30408 1360 30472
rect 0 30400 1360 30408
rect 28640 30472 30000 30480
rect 28640 30408 28968 30472
rect 29032 30408 29288 30472
rect 29352 30408 29608 30472
rect 29672 30408 29928 30472
rect 29992 30408 30000 30472
rect 28640 30400 30000 30408
rect 0 30312 1360 30320
rect 0 30248 8 30312
rect 72 30248 328 30312
rect 392 30248 648 30312
rect 712 30248 968 30312
rect 1032 30248 1360 30312
rect 0 30240 1360 30248
rect 28640 30312 30000 30320
rect 28640 30248 28968 30312
rect 29032 30248 29288 30312
rect 29352 30248 29608 30312
rect 29672 30248 29928 30312
rect 29992 30248 30000 30312
rect 28640 30240 30000 30248
rect 0 30152 1360 30160
rect 0 30088 8 30152
rect 72 30088 328 30152
rect 392 30088 648 30152
rect 712 30088 968 30152
rect 1032 30088 1360 30152
rect 0 30080 1360 30088
rect 28640 30152 30000 30160
rect 28640 30088 28968 30152
rect 29032 30088 29288 30152
rect 29352 30088 29608 30152
rect 29672 30088 29928 30152
rect 29992 30088 30000 30152
rect 28640 30080 30000 30088
rect 0 29992 1360 30000
rect 0 29928 8 29992
rect 72 29928 328 29992
rect 392 29928 648 29992
rect 712 29928 968 29992
rect 1032 29928 1360 29992
rect 0 29920 1360 29928
rect 28640 29992 30000 30000
rect 28640 29928 28968 29992
rect 29032 29928 29288 29992
rect 29352 29928 29608 29992
rect 29672 29928 29928 29992
rect 29992 29928 30000 29992
rect 28640 29920 30000 29928
rect 0 29832 1360 29840
rect 0 29768 8 29832
rect 72 29768 328 29832
rect 392 29768 648 29832
rect 712 29768 968 29832
rect 1032 29768 1360 29832
rect 0 29760 1360 29768
rect 28640 29832 30000 29840
rect 28640 29768 28968 29832
rect 29032 29768 29288 29832
rect 29352 29768 29608 29832
rect 29672 29768 29928 29832
rect 29992 29768 30000 29832
rect 28640 29760 30000 29768
rect 0 29672 1040 29680
rect 0 29608 8 29672
rect 72 29608 328 29672
rect 392 29608 648 29672
rect 712 29608 968 29672
rect 1032 29608 1040 29672
rect 0 29600 1040 29608
rect 28960 29672 30000 29680
rect 28960 29608 28968 29672
rect 29032 29608 29288 29672
rect 29352 29608 29608 29672
rect 29672 29608 29928 29672
rect 29992 29608 30000 29672
rect 28960 29600 30000 29608
rect 0 29512 1040 29520
rect 0 29448 8 29512
rect 72 29448 328 29512
rect 392 29448 648 29512
rect 712 29448 968 29512
rect 1032 29448 1040 29512
rect 0 29440 1040 29448
rect 28960 29512 30000 29520
rect 28960 29448 28968 29512
rect 29032 29448 29288 29512
rect 29352 29448 29608 29512
rect 29672 29448 29928 29512
rect 29992 29448 30000 29512
rect 28960 29440 30000 29448
rect 0 29352 1360 29360
rect 0 29288 8 29352
rect 72 29288 328 29352
rect 392 29288 648 29352
rect 712 29288 968 29352
rect 1032 29288 1360 29352
rect 0 29280 1360 29288
rect 28720 29352 30000 29360
rect 28720 29288 28968 29352
rect 29032 29288 29288 29352
rect 29352 29288 29608 29352
rect 29672 29288 29928 29352
rect 29992 29288 30000 29352
rect 28720 29280 30000 29288
rect 0 29192 1040 29200
rect 0 29128 8 29192
rect 72 29128 328 29192
rect 392 29128 648 29192
rect 712 29128 968 29192
rect 1032 29128 1040 29192
rect 0 29120 1040 29128
rect 28640 29192 29840 29200
rect 28640 29128 29768 29192
rect 29832 29128 29840 29192
rect 28640 29120 29840 29128
rect 0 29032 1360 29040
rect 0 28968 8 29032
rect 72 28968 328 29032
rect 392 28968 648 29032
rect 712 28968 968 29032
rect 1032 28968 1360 29032
rect 0 28960 1360 28968
rect 28640 29032 30000 29040
rect 28640 28968 28968 29032
rect 29032 28968 29288 29032
rect 29352 28968 29608 29032
rect 29672 28968 29928 29032
rect 29992 28968 30000 29032
rect 28640 28960 30000 28968
rect 0 28872 1040 28880
rect 0 28808 8 28872
rect 72 28808 328 28872
rect 392 28808 648 28872
rect 712 28808 968 28872
rect 1032 28808 1040 28872
rect 0 28800 1040 28808
rect 28640 28872 29520 28880
rect 28640 28808 29448 28872
rect 29512 28808 29520 28872
rect 28640 28800 29520 28808
rect 29600 28872 30000 28880
rect 29600 28808 29608 28872
rect 29672 28808 29928 28872
rect 29992 28808 30000 28872
rect 29600 28800 30000 28808
rect 0 28712 1360 28720
rect 0 28648 8 28712
rect 72 28648 328 28712
rect 392 28648 648 28712
rect 712 28648 968 28712
rect 1032 28648 1360 28712
rect 0 28640 1360 28648
rect 28640 28712 30000 28720
rect 28640 28648 28968 28712
rect 29032 28648 29288 28712
rect 29352 28648 29608 28712
rect 29672 28648 29928 28712
rect 29992 28648 30000 28712
rect 28640 28640 30000 28648
rect 0 28552 1040 28560
rect 0 28488 8 28552
rect 72 28488 328 28552
rect 392 28488 648 28552
rect 712 28488 968 28552
rect 1032 28488 1040 28552
rect 0 28480 1040 28488
rect 28960 28552 30000 28560
rect 28960 28488 28968 28552
rect 29032 28488 29288 28552
rect 29352 28488 29608 28552
rect 29672 28488 29928 28552
rect 29992 28488 30000 28552
rect 28960 28480 30000 28488
rect 0 28392 1040 28400
rect 0 28328 8 28392
rect 72 28328 328 28392
rect 392 28328 648 28392
rect 712 28328 968 28392
rect 1032 28328 1040 28392
rect 0 28320 1040 28328
rect 28960 28392 30000 28400
rect 28960 28328 28968 28392
rect 29032 28328 29288 28392
rect 29352 28328 29608 28392
rect 29672 28328 29928 28392
rect 29992 28328 30000 28392
rect 28960 28320 30000 28328
rect 0 28232 1040 28240
rect 0 28168 8 28232
rect 72 28168 328 28232
rect 392 28168 648 28232
rect 712 28168 968 28232
rect 1032 28168 1040 28232
rect 0 28160 1040 28168
rect 28960 28232 30000 28240
rect 28960 28168 28968 28232
rect 29032 28168 29288 28232
rect 29352 28168 29608 28232
rect 29672 28168 29928 28232
rect 29992 28168 30000 28232
rect 28960 28160 30000 28168
rect 0 28072 1040 28080
rect 0 28008 8 28072
rect 72 28008 328 28072
rect 392 28008 648 28072
rect 712 28008 968 28072
rect 1032 28008 1040 28072
rect 0 28000 1040 28008
rect 28960 28072 30000 28080
rect 28960 28008 28968 28072
rect 29032 28008 29288 28072
rect 29352 28008 29608 28072
rect 29672 28008 29928 28072
rect 29992 28008 30000 28072
rect 28960 28000 30000 28008
rect 0 27912 1040 27920
rect 0 27848 8 27912
rect 72 27848 328 27912
rect 392 27848 648 27912
rect 712 27848 968 27912
rect 1032 27848 1040 27912
rect 0 27840 1040 27848
rect 28960 27912 30000 27920
rect 28960 27848 28968 27912
rect 29032 27848 29288 27912
rect 29352 27848 29608 27912
rect 29672 27848 29928 27912
rect 29992 27848 30000 27912
rect 28960 27840 30000 27848
rect 0 27752 1040 27760
rect 0 27688 8 27752
rect 72 27688 328 27752
rect 392 27688 648 27752
rect 712 27688 968 27752
rect 1032 27688 1040 27752
rect 0 27680 1040 27688
rect 28960 27752 30000 27760
rect 28960 27688 28968 27752
rect 29032 27688 29288 27752
rect 29352 27688 29608 27752
rect 29672 27688 29928 27752
rect 29992 27688 30000 27752
rect 28960 27680 30000 27688
rect 0 27592 1040 27600
rect 0 27528 8 27592
rect 72 27528 328 27592
rect 392 27528 648 27592
rect 712 27528 968 27592
rect 1032 27528 1040 27592
rect 0 27520 1040 27528
rect 28960 27592 30000 27600
rect 28960 27528 28968 27592
rect 29032 27528 29288 27592
rect 29352 27528 29608 27592
rect 29672 27528 29928 27592
rect 29992 27528 30000 27592
rect 28960 27520 30000 27528
rect 0 27432 1040 27440
rect 0 27368 8 27432
rect 72 27368 328 27432
rect 392 27368 648 27432
rect 712 27368 968 27432
rect 1032 27368 1040 27432
rect 0 27360 1040 27368
rect 28960 27432 30000 27440
rect 28960 27368 28968 27432
rect 29032 27368 29288 27432
rect 29352 27368 29608 27432
rect 29672 27368 29928 27432
rect 29992 27368 30000 27432
rect 28960 27360 30000 27368
rect 0 27272 1040 27280
rect 0 27208 8 27272
rect 72 27208 328 27272
rect 392 27208 648 27272
rect 712 27208 968 27272
rect 1032 27208 1040 27272
rect 0 27200 1040 27208
rect 28960 27272 30000 27280
rect 28960 27208 28968 27272
rect 29032 27208 29288 27272
rect 29352 27208 29608 27272
rect 29672 27208 29928 27272
rect 29992 27208 30000 27272
rect 28960 27200 30000 27208
rect 0 27112 1040 27120
rect 0 27048 8 27112
rect 72 27048 328 27112
rect 392 27048 648 27112
rect 712 27048 968 27112
rect 1032 27048 1040 27112
rect 0 27040 1040 27048
rect 28960 27112 30000 27120
rect 28960 27048 28968 27112
rect 29032 27048 29288 27112
rect 29352 27048 29608 27112
rect 29672 27048 29928 27112
rect 29992 27048 30000 27112
rect 28960 27040 30000 27048
rect 0 26952 1040 26960
rect 0 26888 8 26952
rect 72 26888 328 26952
rect 392 26888 648 26952
rect 712 26888 968 26952
rect 1032 26888 1040 26952
rect 0 26880 1040 26888
rect 28960 26952 30000 26960
rect 28960 26888 28968 26952
rect 29032 26888 29288 26952
rect 29352 26888 29608 26952
rect 29672 26888 29928 26952
rect 29992 26888 30000 26952
rect 28960 26880 30000 26888
rect 0 26792 1040 26800
rect 0 26728 8 26792
rect 72 26728 328 26792
rect 392 26728 648 26792
rect 712 26728 968 26792
rect 1032 26728 1040 26792
rect 0 26720 1040 26728
rect 28960 26792 30000 26800
rect 28960 26728 28968 26792
rect 29032 26728 29288 26792
rect 29352 26728 29608 26792
rect 29672 26728 29928 26792
rect 29992 26728 30000 26792
rect 28960 26720 30000 26728
rect 0 26632 1040 26640
rect 0 26568 8 26632
rect 72 26568 328 26632
rect 392 26568 648 26632
rect 712 26568 968 26632
rect 1032 26568 1040 26632
rect 0 26560 1040 26568
rect 28960 26632 30000 26640
rect 28960 26568 28968 26632
rect 29032 26568 29288 26632
rect 29352 26568 29608 26632
rect 29672 26568 29928 26632
rect 29992 26568 30000 26632
rect 28960 26560 30000 26568
rect 0 26472 1040 26480
rect 0 26408 8 26472
rect 72 26408 328 26472
rect 392 26408 648 26472
rect 712 26408 968 26472
rect 1032 26408 1040 26472
rect 0 26400 1040 26408
rect 28960 26472 30000 26480
rect 28960 26408 28968 26472
rect 29032 26408 29288 26472
rect 29352 26408 29608 26472
rect 29672 26408 29928 26472
rect 29992 26408 30000 26472
rect 28960 26400 30000 26408
rect 0 26312 1040 26320
rect 0 26248 8 26312
rect 72 26248 328 26312
rect 392 26248 648 26312
rect 712 26248 968 26312
rect 1032 26248 1040 26312
rect 0 26240 1040 26248
rect 28720 26312 29200 26320
rect 28720 26248 29128 26312
rect 29192 26248 29200 26312
rect 28720 26240 29200 26248
rect 29280 26312 30000 26320
rect 29280 26248 29288 26312
rect 29352 26248 29608 26312
rect 29672 26248 29928 26312
rect 29992 26248 30000 26312
rect 29280 26240 30000 26248
rect 0 26152 1040 26160
rect 0 26088 8 26152
rect 72 26088 328 26152
rect 392 26088 648 26152
rect 712 26088 968 26152
rect 1032 26088 1040 26152
rect 0 26080 1040 26088
rect 28960 26152 30000 26160
rect 28960 26088 28968 26152
rect 29032 26088 29288 26152
rect 29352 26088 29608 26152
rect 29672 26088 29928 26152
rect 29992 26088 30000 26152
rect 28960 26080 30000 26088
rect 0 25992 1040 26000
rect 0 25928 8 25992
rect 72 25928 328 25992
rect 392 25928 648 25992
rect 712 25928 968 25992
rect 1032 25928 1040 25992
rect 0 25920 1040 25928
rect 28960 25992 30000 26000
rect 28960 25928 28968 25992
rect 29032 25928 29288 25992
rect 29352 25928 29608 25992
rect 29672 25928 29928 25992
rect 29992 25928 30000 25992
rect 28960 25920 30000 25928
rect 0 25832 1040 25840
rect 0 25768 8 25832
rect 72 25768 328 25832
rect 392 25768 648 25832
rect 712 25768 968 25832
rect 1032 25768 1040 25832
rect 0 25760 1040 25768
rect 28960 25832 30000 25840
rect 28960 25768 28968 25832
rect 29032 25768 29288 25832
rect 29352 25768 29608 25832
rect 29672 25768 29928 25832
rect 29992 25768 30000 25832
rect 28960 25760 30000 25768
rect 0 25672 1040 25680
rect 0 25608 8 25672
rect 72 25608 328 25672
rect 392 25608 648 25672
rect 712 25608 968 25672
rect 1032 25608 1040 25672
rect 0 25600 1040 25608
rect 28960 25672 30000 25680
rect 28960 25608 28968 25672
rect 29032 25608 29288 25672
rect 29352 25608 29608 25672
rect 29672 25608 29928 25672
rect 29992 25608 30000 25672
rect 28960 25600 30000 25608
rect 0 25512 1040 25520
rect 0 25448 8 25512
rect 72 25448 328 25512
rect 392 25448 648 25512
rect 712 25448 968 25512
rect 1032 25448 1040 25512
rect 0 25440 1040 25448
rect 28960 25512 30000 25520
rect 28960 25448 28968 25512
rect 29032 25448 29288 25512
rect 29352 25448 29608 25512
rect 29672 25448 29928 25512
rect 29992 25448 30000 25512
rect 28960 25440 30000 25448
rect 0 25352 1040 25360
rect 0 25288 8 25352
rect 72 25288 328 25352
rect 392 25288 648 25352
rect 712 25288 968 25352
rect 1032 25288 1040 25352
rect 0 25280 1040 25288
rect 28960 25352 30000 25360
rect 28960 25288 28968 25352
rect 29032 25288 29288 25352
rect 29352 25288 29608 25352
rect 29672 25288 29928 25352
rect 29992 25288 30000 25352
rect 28960 25280 30000 25288
rect 0 25192 1040 25200
rect 0 25128 8 25192
rect 72 25128 328 25192
rect 392 25128 648 25192
rect 712 25128 968 25192
rect 1032 25128 1040 25192
rect 0 25120 1040 25128
rect 28960 25192 30000 25200
rect 28960 25128 28968 25192
rect 29032 25128 29288 25192
rect 29352 25128 29608 25192
rect 29672 25128 29928 25192
rect 29992 25128 30000 25192
rect 28960 25120 30000 25128
rect 0 25032 1040 25040
rect 0 24968 8 25032
rect 72 24968 328 25032
rect 392 24968 648 25032
rect 712 24968 968 25032
rect 1032 24968 1040 25032
rect 0 24960 1040 24968
rect 28960 25032 30000 25040
rect 28960 24968 28968 25032
rect 29032 24968 29288 25032
rect 29352 24968 29608 25032
rect 29672 24968 29928 25032
rect 29992 24968 30000 25032
rect 28960 24960 30000 24968
rect 0 24872 1040 24880
rect 0 24808 8 24872
rect 72 24808 328 24872
rect 392 24808 648 24872
rect 712 24808 968 24872
rect 1032 24808 1040 24872
rect 0 24800 1040 24808
rect 28960 24872 30000 24880
rect 28960 24808 28968 24872
rect 29032 24808 29288 24872
rect 29352 24808 29608 24872
rect 29672 24808 29928 24872
rect 29992 24808 30000 24872
rect 28960 24800 30000 24808
rect 0 24712 1040 24720
rect 0 24648 8 24712
rect 72 24648 328 24712
rect 392 24648 648 24712
rect 712 24648 968 24712
rect 1032 24648 1040 24712
rect 0 24640 1040 24648
rect 28960 24712 30000 24720
rect 28960 24648 28968 24712
rect 29032 24648 29288 24712
rect 29352 24648 29608 24712
rect 29672 24648 29928 24712
rect 29992 24648 30000 24712
rect 28960 24640 30000 24648
rect 0 24552 1040 24560
rect 0 24488 8 24552
rect 72 24488 328 24552
rect 392 24488 648 24552
rect 712 24488 968 24552
rect 1032 24488 1040 24552
rect 0 24480 1040 24488
rect 28960 24552 30000 24560
rect 28960 24488 28968 24552
rect 29032 24488 29288 24552
rect 29352 24488 29608 24552
rect 29672 24488 29928 24552
rect 29992 24488 30000 24552
rect 28960 24480 30000 24488
rect 0 24392 1040 24400
rect 0 24328 8 24392
rect 72 24328 328 24392
rect 392 24328 648 24392
rect 712 24328 968 24392
rect 1032 24328 1040 24392
rect 0 24320 1040 24328
rect 28960 24392 30000 24400
rect 28960 24328 28968 24392
rect 29032 24328 29288 24392
rect 29352 24328 29608 24392
rect 29672 24328 29928 24392
rect 29992 24328 30000 24392
rect 28960 24320 30000 24328
rect 0 24232 1040 24240
rect 0 24168 8 24232
rect 72 24168 328 24232
rect 392 24168 648 24232
rect 712 24168 968 24232
rect 1032 24168 1040 24232
rect 0 24160 1040 24168
rect 28960 24232 30000 24240
rect 28960 24168 28968 24232
rect 29032 24168 29288 24232
rect 29352 24168 29608 24232
rect 29672 24168 29928 24232
rect 29992 24168 30000 24232
rect 28960 24160 30000 24168
rect 0 24072 1040 24080
rect 0 24008 8 24072
rect 72 24008 328 24072
rect 392 24008 648 24072
rect 712 24008 968 24072
rect 1032 24008 1040 24072
rect 0 24000 1040 24008
rect 28960 24072 30000 24080
rect 28960 24008 28968 24072
rect 29032 24008 29288 24072
rect 29352 24008 29608 24072
rect 29672 24008 29928 24072
rect 29992 24008 30000 24072
rect 28960 24000 30000 24008
rect 0 23912 1360 23920
rect 0 23848 8 23912
rect 72 23848 328 23912
rect 392 23848 648 23912
rect 712 23848 968 23912
rect 1032 23848 1360 23912
rect 0 23840 1360 23848
rect 28720 23912 30000 23920
rect 28720 23848 28968 23912
rect 29032 23848 29288 23912
rect 29352 23848 29608 23912
rect 29672 23848 29928 23912
rect 29992 23848 30000 23912
rect 28720 23840 30000 23848
rect 0 23752 1040 23760
rect 0 23688 8 23752
rect 72 23688 328 23752
rect 392 23688 648 23752
rect 712 23688 968 23752
rect 1032 23688 1040 23752
rect 0 23680 1040 23688
rect 28640 23752 29520 23760
rect 28640 23688 29448 23752
rect 29512 23688 29520 23752
rect 28640 23680 29520 23688
rect 29600 23752 30000 23760
rect 29600 23688 29608 23752
rect 29672 23688 29928 23752
rect 29992 23688 30000 23752
rect 29600 23680 30000 23688
rect 0 23592 1360 23600
rect 0 23528 8 23592
rect 72 23528 328 23592
rect 392 23528 648 23592
rect 712 23528 968 23592
rect 1032 23528 1360 23592
rect 0 23520 1360 23528
rect 28720 23592 30000 23600
rect 28720 23528 28968 23592
rect 29032 23528 29288 23592
rect 29352 23528 29608 23592
rect 29672 23528 29928 23592
rect 29992 23528 30000 23592
rect 28720 23520 30000 23528
rect 0 23432 1040 23440
rect 0 23368 8 23432
rect 72 23368 328 23432
rect 392 23368 648 23432
rect 712 23368 968 23432
rect 1032 23368 1040 23432
rect 0 23360 1040 23368
rect 28640 23432 29840 23440
rect 28640 23368 29768 23432
rect 29832 23368 29840 23432
rect 28640 23360 29840 23368
rect 0 23272 1360 23280
rect 0 23208 8 23272
rect 72 23208 328 23272
rect 392 23208 648 23272
rect 712 23208 968 23272
rect 1032 23208 1360 23272
rect 0 23200 1360 23208
rect 28720 23272 30000 23280
rect 28720 23208 28968 23272
rect 29032 23208 29288 23272
rect 29352 23208 29608 23272
rect 29672 23208 29928 23272
rect 29992 23208 30000 23272
rect 28720 23200 30000 23208
rect 0 23112 1040 23120
rect 0 23048 8 23112
rect 72 23048 328 23112
rect 392 23048 648 23112
rect 712 23048 968 23112
rect 1032 23048 1040 23112
rect 0 23040 1040 23048
rect 28960 23112 30000 23120
rect 28960 23048 28968 23112
rect 29032 23048 29288 23112
rect 29352 23048 29608 23112
rect 29672 23048 29928 23112
rect 29992 23048 30000 23112
rect 28960 23040 30000 23048
rect 0 22952 1040 22960
rect 0 22888 8 22952
rect 72 22888 328 22952
rect 392 22888 648 22952
rect 712 22888 968 22952
rect 1032 22888 1040 22952
rect 0 22880 1040 22888
rect 28960 22952 30000 22960
rect 28960 22888 28968 22952
rect 29032 22888 29288 22952
rect 29352 22888 29608 22952
rect 29672 22888 29928 22952
rect 29992 22888 30000 22952
rect 28960 22880 30000 22888
rect 0 22792 1360 22800
rect 0 22728 8 22792
rect 72 22728 328 22792
rect 392 22728 648 22792
rect 712 22728 968 22792
rect 1032 22728 1360 22792
rect 0 22720 1360 22728
rect 28640 22792 30000 22800
rect 28640 22728 28968 22792
rect 29032 22728 29288 22792
rect 29352 22728 29608 22792
rect 29672 22728 29928 22792
rect 29992 22728 30000 22792
rect 28640 22720 30000 22728
rect 160 22632 1360 22640
rect 160 22568 168 22632
rect 232 22568 1360 22632
rect 160 22560 1360 22568
rect 28960 22632 30000 22640
rect 28960 22568 28968 22632
rect 29032 22568 29288 22632
rect 29352 22568 29608 22632
rect 29672 22568 29928 22632
rect 29992 22568 30000 22632
rect 28960 22560 30000 22568
rect 0 22472 1360 22480
rect 0 22408 8 22472
rect 72 22408 328 22472
rect 392 22408 648 22472
rect 712 22408 968 22472
rect 1032 22408 1360 22472
rect 0 22400 1360 22408
rect 28640 22472 30000 22480
rect 28640 22408 28968 22472
rect 29032 22408 29288 22472
rect 29352 22408 29608 22472
rect 29672 22408 29928 22472
rect 29992 22408 30000 22472
rect 28640 22400 30000 22408
rect 0 22312 400 22320
rect 0 22248 8 22312
rect 72 22248 328 22312
rect 392 22248 400 22312
rect 0 22240 400 22248
rect 480 22312 1360 22320
rect 480 22248 488 22312
rect 552 22248 1360 22312
rect 480 22240 1360 22248
rect 28960 22312 30000 22320
rect 28960 22248 28968 22312
rect 29032 22248 29288 22312
rect 29352 22248 29608 22312
rect 29672 22248 29928 22312
rect 29992 22248 30000 22312
rect 28960 22240 30000 22248
rect 0 22152 1040 22160
rect 0 22088 8 22152
rect 72 22088 328 22152
rect 392 22088 648 22152
rect 712 22088 968 22152
rect 1032 22088 1040 22152
rect 0 22080 1040 22088
rect 28640 22152 30000 22160
rect 28640 22088 28968 22152
rect 29032 22088 29288 22152
rect 29352 22088 29608 22152
rect 29672 22088 29928 22152
rect 29992 22088 30000 22152
rect 28640 22080 30000 22088
rect 0 21992 1040 22000
rect 0 21928 8 21992
rect 72 21928 328 21992
rect 392 21928 648 21992
rect 712 21928 968 21992
rect 1032 21928 1040 21992
rect 0 21920 1040 21928
rect 28960 21992 30000 22000
rect 28960 21928 28968 21992
rect 29032 21928 29288 21992
rect 29352 21928 29608 21992
rect 29672 21928 29928 21992
rect 29992 21928 30000 21992
rect 28960 21920 30000 21928
rect 0 21832 1040 21840
rect 0 21768 8 21832
rect 72 21768 328 21832
rect 392 21768 648 21832
rect 712 21768 968 21832
rect 1032 21768 1040 21832
rect 0 21760 1040 21768
rect 28960 21832 30000 21840
rect 28960 21768 28968 21832
rect 29032 21768 29288 21832
rect 29352 21768 29608 21832
rect 29672 21768 29928 21832
rect 29992 21768 30000 21832
rect 28960 21760 30000 21768
rect 0 21672 1040 21680
rect 0 21608 8 21672
rect 72 21608 328 21672
rect 392 21608 648 21672
rect 712 21608 968 21672
rect 1032 21608 1040 21672
rect 0 21600 1040 21608
rect 28960 21672 30000 21680
rect 28960 21608 28968 21672
rect 29032 21608 29288 21672
rect 29352 21608 29608 21672
rect 29672 21608 29928 21672
rect 29992 21608 30000 21672
rect 28960 21600 30000 21608
rect 0 21512 1040 21520
rect 0 21448 8 21512
rect 72 21448 328 21512
rect 392 21448 648 21512
rect 712 21448 968 21512
rect 1032 21448 1040 21512
rect 0 21440 1040 21448
rect 28960 21512 30000 21520
rect 28960 21448 28968 21512
rect 29032 21448 29288 21512
rect 29352 21448 29608 21512
rect 29672 21448 29928 21512
rect 29992 21448 30000 21512
rect 28960 21440 30000 21448
rect 0 21352 1040 21360
rect 0 21288 8 21352
rect 72 21288 328 21352
rect 392 21288 648 21352
rect 712 21288 968 21352
rect 1032 21288 1040 21352
rect 0 21280 1040 21288
rect 28960 21352 30000 21360
rect 28960 21288 28968 21352
rect 29032 21288 29288 21352
rect 29352 21288 29608 21352
rect 29672 21288 29928 21352
rect 29992 21288 30000 21352
rect 28960 21280 30000 21288
rect 0 21192 1040 21200
rect 0 21128 8 21192
rect 72 21128 328 21192
rect 392 21128 648 21192
rect 712 21128 968 21192
rect 1032 21128 1040 21192
rect 0 21120 1040 21128
rect 28960 21192 30000 21200
rect 28960 21128 28968 21192
rect 29032 21128 29288 21192
rect 29352 21128 29608 21192
rect 29672 21128 29928 21192
rect 29992 21128 30000 21192
rect 28960 21120 30000 21128
rect 0 21032 1040 21040
rect 0 20968 8 21032
rect 72 20968 328 21032
rect 392 20968 648 21032
rect 712 20968 968 21032
rect 1032 20968 1040 21032
rect 0 20960 1040 20968
rect 28960 21032 30000 21040
rect 28960 20968 28968 21032
rect 29032 20968 29288 21032
rect 29352 20968 29608 21032
rect 29672 20968 29928 21032
rect 29992 20968 30000 21032
rect 28960 20960 30000 20968
rect 0 20872 1040 20880
rect 0 20808 8 20872
rect 72 20808 328 20872
rect 392 20808 648 20872
rect 712 20808 968 20872
rect 1032 20808 1040 20872
rect 0 20800 1040 20808
rect 28960 20872 30000 20880
rect 28960 20808 28968 20872
rect 29032 20808 29288 20872
rect 29352 20808 29608 20872
rect 29672 20808 29928 20872
rect 29992 20808 30000 20872
rect 28960 20800 30000 20808
rect 0 20712 1040 20720
rect 0 20648 8 20712
rect 72 20648 328 20712
rect 392 20648 648 20712
rect 712 20648 968 20712
rect 1032 20648 1040 20712
rect 0 20640 1040 20648
rect 28960 20712 30000 20720
rect 28960 20648 28968 20712
rect 29032 20648 29288 20712
rect 29352 20648 29608 20712
rect 29672 20648 29928 20712
rect 29992 20648 30000 20712
rect 28960 20640 30000 20648
rect 0 20552 1040 20560
rect 0 20488 8 20552
rect 72 20488 328 20552
rect 392 20488 648 20552
rect 712 20488 968 20552
rect 1032 20488 1040 20552
rect 0 20480 1040 20488
rect 28960 20552 30000 20560
rect 28960 20488 28968 20552
rect 29032 20488 29288 20552
rect 29352 20488 29608 20552
rect 29672 20488 29928 20552
rect 29992 20488 30000 20552
rect 28960 20480 30000 20488
rect 0 20392 1040 20400
rect 0 20328 8 20392
rect 72 20328 328 20392
rect 392 20328 648 20392
rect 712 20328 968 20392
rect 1032 20328 1040 20392
rect 0 20320 1040 20328
rect 28960 20392 30000 20400
rect 28960 20328 28968 20392
rect 29032 20328 29288 20392
rect 29352 20328 29608 20392
rect 29672 20328 29928 20392
rect 29992 20328 30000 20392
rect 28960 20320 30000 20328
rect 0 20232 1040 20240
rect 0 20168 8 20232
rect 72 20168 328 20232
rect 392 20168 648 20232
rect 712 20168 968 20232
rect 1032 20168 1040 20232
rect 0 20160 1040 20168
rect 28960 20232 30000 20240
rect 28960 20168 28968 20232
rect 29032 20168 29288 20232
rect 29352 20168 29608 20232
rect 29672 20168 29928 20232
rect 29992 20168 30000 20232
rect 28960 20160 30000 20168
rect 0 20072 1040 20080
rect 0 20008 8 20072
rect 72 20008 328 20072
rect 392 20008 648 20072
rect 712 20008 968 20072
rect 1032 20008 1040 20072
rect 0 20000 1040 20008
rect 28960 20072 30000 20080
rect 28960 20008 28968 20072
rect 29032 20008 29288 20072
rect 29352 20008 29608 20072
rect 29672 20008 29928 20072
rect 29992 20008 30000 20072
rect 28960 20000 30000 20008
rect 0 19912 1040 19920
rect 0 19848 8 19912
rect 72 19848 328 19912
rect 392 19848 648 19912
rect 712 19848 968 19912
rect 1032 19848 1040 19912
rect 0 19840 1040 19848
rect 28960 19912 30000 19920
rect 28960 19848 28968 19912
rect 29032 19848 29288 19912
rect 29352 19848 29608 19912
rect 29672 19848 29928 19912
rect 29992 19848 30000 19912
rect 28960 19840 30000 19848
rect 0 19752 720 19760
rect 0 19688 8 19752
rect 72 19688 328 19752
rect 392 19688 648 19752
rect 712 19688 720 19752
rect 0 19680 720 19688
rect 800 19752 1360 19760
rect 800 19688 808 19752
rect 872 19688 1360 19752
rect 800 19680 1360 19688
rect 28960 19752 30000 19760
rect 28960 19688 28968 19752
rect 29032 19688 29288 19752
rect 29352 19688 29608 19752
rect 29672 19688 29928 19752
rect 29992 19688 30000 19752
rect 28960 19680 30000 19688
rect 0 19592 1040 19600
rect 0 19528 8 19592
rect 72 19528 328 19592
rect 392 19528 648 19592
rect 712 19528 968 19592
rect 1032 19528 1040 19592
rect 0 19520 1040 19528
rect 28960 19592 30000 19600
rect 28960 19528 28968 19592
rect 29032 19528 29288 19592
rect 29352 19528 29608 19592
rect 29672 19528 29928 19592
rect 29992 19528 30000 19592
rect 28960 19520 30000 19528
rect 0 19432 1040 19440
rect 0 19368 8 19432
rect 72 19368 328 19432
rect 392 19368 648 19432
rect 712 19368 968 19432
rect 1032 19368 1040 19432
rect 0 19360 1040 19368
rect 28960 19432 30000 19440
rect 28960 19368 28968 19432
rect 29032 19368 29288 19432
rect 29352 19368 29608 19432
rect 29672 19368 29928 19432
rect 29992 19368 30000 19432
rect 28960 19360 30000 19368
rect 0 19272 1040 19280
rect 0 19208 8 19272
rect 72 19208 328 19272
rect 392 19208 648 19272
rect 712 19208 968 19272
rect 1032 19208 1040 19272
rect 0 19200 1040 19208
rect 28960 19272 30000 19280
rect 28960 19208 28968 19272
rect 29032 19208 29288 19272
rect 29352 19208 29608 19272
rect 29672 19208 29928 19272
rect 29992 19208 30000 19272
rect 28960 19200 30000 19208
rect 0 19112 1040 19120
rect 0 19048 8 19112
rect 72 19048 328 19112
rect 392 19048 648 19112
rect 712 19048 968 19112
rect 1032 19048 1040 19112
rect 0 19040 1040 19048
rect 28960 19112 30000 19120
rect 28960 19048 28968 19112
rect 29032 19048 29288 19112
rect 29352 19048 29608 19112
rect 29672 19048 29928 19112
rect 29992 19048 30000 19112
rect 28960 19040 30000 19048
rect 0 18952 1040 18960
rect 0 18888 8 18952
rect 72 18888 328 18952
rect 392 18888 648 18952
rect 712 18888 968 18952
rect 1032 18888 1040 18952
rect 0 18880 1040 18888
rect 28960 18952 30000 18960
rect 28960 18888 28968 18952
rect 29032 18888 29288 18952
rect 29352 18888 29608 18952
rect 29672 18888 29928 18952
rect 29992 18888 30000 18952
rect 28960 18880 30000 18888
rect 0 18792 1040 18800
rect 0 18728 8 18792
rect 72 18728 328 18792
rect 392 18728 648 18792
rect 712 18728 968 18792
rect 1032 18728 1040 18792
rect 0 18720 1040 18728
rect 28960 18792 30000 18800
rect 28960 18728 28968 18792
rect 29032 18728 29288 18792
rect 29352 18728 29608 18792
rect 29672 18728 29928 18792
rect 29992 18728 30000 18792
rect 28960 18720 30000 18728
rect 0 18632 1040 18640
rect 0 18568 8 18632
rect 72 18568 328 18632
rect 392 18568 648 18632
rect 712 18568 968 18632
rect 1032 18568 1040 18632
rect 0 18560 1040 18568
rect 28960 18632 30000 18640
rect 28960 18568 28968 18632
rect 29032 18568 29288 18632
rect 29352 18568 29608 18632
rect 29672 18568 29928 18632
rect 29992 18568 30000 18632
rect 28960 18560 30000 18568
rect 0 18472 1040 18480
rect 0 18408 8 18472
rect 72 18408 328 18472
rect 392 18408 648 18472
rect 712 18408 968 18472
rect 1032 18408 1040 18472
rect 0 18400 1040 18408
rect 28960 18472 30000 18480
rect 28960 18408 28968 18472
rect 29032 18408 29288 18472
rect 29352 18408 29608 18472
rect 29672 18408 29928 18472
rect 29992 18408 30000 18472
rect 28960 18400 30000 18408
rect 0 18312 1040 18320
rect 0 18248 8 18312
rect 72 18248 328 18312
rect 392 18248 648 18312
rect 712 18248 968 18312
rect 1032 18248 1040 18312
rect 0 18240 1040 18248
rect 28960 18312 30000 18320
rect 28960 18248 28968 18312
rect 29032 18248 29288 18312
rect 29352 18248 29608 18312
rect 29672 18248 29928 18312
rect 29992 18248 30000 18312
rect 28960 18240 30000 18248
rect 0 18152 1040 18160
rect 0 18088 8 18152
rect 72 18088 328 18152
rect 392 18088 648 18152
rect 712 18088 968 18152
rect 1032 18088 1040 18152
rect 0 18080 1040 18088
rect 28960 18152 30000 18160
rect 28960 18088 28968 18152
rect 29032 18088 29288 18152
rect 29352 18088 29608 18152
rect 29672 18088 29928 18152
rect 29992 18088 30000 18152
rect 28960 18080 30000 18088
rect 0 17992 1040 18000
rect 0 17928 8 17992
rect 72 17928 328 17992
rect 392 17928 648 17992
rect 712 17928 968 17992
rect 1032 17928 1040 17992
rect 0 17920 1040 17928
rect 28960 17992 30000 18000
rect 28960 17928 28968 17992
rect 29032 17928 29288 17992
rect 29352 17928 29608 17992
rect 29672 17928 29928 17992
rect 29992 17928 30000 17992
rect 28960 17920 30000 17928
rect 0 17832 1040 17840
rect 0 17768 8 17832
rect 72 17768 328 17832
rect 392 17768 648 17832
rect 712 17768 968 17832
rect 1032 17768 1040 17832
rect 0 17760 1040 17768
rect 28960 17832 30000 17840
rect 28960 17768 28968 17832
rect 29032 17768 29288 17832
rect 29352 17768 29608 17832
rect 29672 17768 29928 17832
rect 29992 17768 30000 17832
rect 28960 17760 30000 17768
rect 0 17672 1040 17680
rect 0 17608 8 17672
rect 72 17608 328 17672
rect 392 17608 648 17672
rect 712 17608 968 17672
rect 1032 17608 1040 17672
rect 0 17600 1040 17608
rect 28960 17672 30000 17680
rect 28960 17608 28968 17672
rect 29032 17608 29288 17672
rect 29352 17608 29608 17672
rect 29672 17608 29928 17672
rect 29992 17608 30000 17672
rect 28960 17600 30000 17608
rect 0 17512 1040 17520
rect 0 17448 8 17512
rect 72 17448 328 17512
rect 392 17448 648 17512
rect 712 17448 968 17512
rect 1032 17448 1040 17512
rect 0 17440 1040 17448
rect 28960 17512 30000 17520
rect 28960 17448 28968 17512
rect 29032 17448 29288 17512
rect 29352 17448 29608 17512
rect 29672 17448 29928 17512
rect 29992 17448 30000 17512
rect 28960 17440 30000 17448
rect 0 17352 1360 17360
rect 0 17288 8 17352
rect 72 17288 328 17352
rect 392 17288 648 17352
rect 712 17288 968 17352
rect 1032 17288 1360 17352
rect 0 17280 1360 17288
rect 28640 17352 30000 17360
rect 28640 17288 28968 17352
rect 29032 17288 29288 17352
rect 29352 17288 29608 17352
rect 29672 17288 29928 17352
rect 29992 17288 30000 17352
rect 28640 17280 30000 17288
rect 0 17192 400 17200
rect 0 17128 8 17192
rect 72 17128 328 17192
rect 392 17128 400 17192
rect 0 17120 400 17128
rect 480 17192 1360 17200
rect 480 17128 488 17192
rect 552 17128 1360 17192
rect 480 17120 1360 17128
rect 28960 17192 30000 17200
rect 28960 17128 28968 17192
rect 29032 17128 29288 17192
rect 29352 17128 29608 17192
rect 29672 17128 29928 17192
rect 29992 17128 30000 17192
rect 28960 17120 30000 17128
rect 0 17032 1360 17040
rect 0 16968 8 17032
rect 72 16968 328 17032
rect 392 16968 648 17032
rect 712 16968 968 17032
rect 1032 16968 1360 17032
rect 0 16960 1360 16968
rect 28640 17032 30000 17040
rect 28640 16968 28968 17032
rect 29032 16968 29288 17032
rect 29352 16968 29608 17032
rect 29672 16968 29928 17032
rect 29992 16968 30000 17032
rect 28640 16960 30000 16968
rect 160 16872 1360 16880
rect 160 16808 168 16872
rect 232 16808 1360 16872
rect 160 16800 1360 16808
rect 28960 16872 30000 16880
rect 28960 16808 28968 16872
rect 29032 16808 29288 16872
rect 29352 16808 29608 16872
rect 29672 16808 29928 16872
rect 29992 16808 30000 16872
rect 28960 16800 30000 16808
rect 0 16712 1360 16720
rect 0 16648 8 16712
rect 72 16648 328 16712
rect 392 16648 648 16712
rect 712 16648 968 16712
rect 1032 16648 1360 16712
rect 0 16640 1360 16648
rect 28640 16712 30000 16720
rect 28640 16648 28968 16712
rect 29032 16648 29288 16712
rect 29352 16648 29608 16712
rect 29672 16648 29928 16712
rect 29992 16648 30000 16712
rect 28640 16640 30000 16648
rect 0 16552 1040 16560
rect 0 16488 8 16552
rect 72 16488 328 16552
rect 392 16488 648 16552
rect 712 16488 968 16552
rect 1032 16488 1040 16552
rect 0 16480 1040 16488
rect 28960 16552 30000 16560
rect 28960 16488 28968 16552
rect 29032 16488 29288 16552
rect 29352 16488 29608 16552
rect 29672 16488 29928 16552
rect 29992 16488 30000 16552
rect 28960 16480 30000 16488
rect 0 16392 1040 16400
rect 0 16328 8 16392
rect 72 16328 328 16392
rect 392 16328 648 16392
rect 712 16328 968 16392
rect 1032 16328 1040 16392
rect 0 16320 1040 16328
rect 28960 16392 30000 16400
rect 28960 16328 28968 16392
rect 29032 16328 29288 16392
rect 29352 16328 29608 16392
rect 29672 16328 29928 16392
rect 29992 16328 30000 16392
rect 28960 16320 30000 16328
rect 0 16232 1360 16240
rect 0 16168 8 16232
rect 72 16168 328 16232
rect 392 16168 648 16232
rect 712 16168 968 16232
rect 1032 16168 1360 16232
rect 0 16160 1360 16168
rect 28640 16232 30000 16240
rect 28640 16168 28968 16232
rect 29032 16168 29288 16232
rect 29352 16168 29608 16232
rect 29672 16168 29928 16232
rect 29992 16168 30000 16232
rect 28640 16160 30000 16168
rect 160 16072 1360 16080
rect 160 16008 168 16072
rect 232 16008 1360 16072
rect 160 16000 1360 16008
rect 28960 16072 30000 16080
rect 28960 16008 28968 16072
rect 29032 16008 29288 16072
rect 29352 16008 29608 16072
rect 29672 16008 29928 16072
rect 29992 16008 30000 16072
rect 28960 16000 30000 16008
rect 0 15912 1360 15920
rect 0 15848 8 15912
rect 72 15848 328 15912
rect 392 15848 648 15912
rect 712 15848 968 15912
rect 1032 15848 1360 15912
rect 0 15840 1360 15848
rect 28640 15912 30000 15920
rect 28640 15848 28968 15912
rect 29032 15848 29288 15912
rect 29352 15848 29608 15912
rect 29672 15848 29928 15912
rect 29992 15848 30000 15912
rect 28640 15840 30000 15848
rect 0 15752 400 15760
rect 0 15688 8 15752
rect 72 15688 328 15752
rect 392 15688 400 15752
rect 0 15680 400 15688
rect 480 15752 1360 15760
rect 480 15688 488 15752
rect 552 15688 1360 15752
rect 480 15680 1360 15688
rect 28960 15752 30000 15760
rect 28960 15688 28968 15752
rect 29032 15688 29288 15752
rect 29352 15688 29608 15752
rect 29672 15688 29928 15752
rect 29992 15688 30000 15752
rect 28960 15680 30000 15688
rect 0 15592 1360 15600
rect 0 15528 8 15592
rect 72 15528 328 15592
rect 392 15528 648 15592
rect 712 15528 968 15592
rect 1032 15528 1360 15592
rect 0 15520 1360 15528
rect 28640 15592 30000 15600
rect 28640 15528 28968 15592
rect 29032 15528 29288 15592
rect 29352 15528 29608 15592
rect 29672 15528 29928 15592
rect 29992 15528 30000 15592
rect 28640 15520 30000 15528
rect 0 15432 1040 15440
rect 0 15368 8 15432
rect 72 15368 328 15432
rect 392 15368 648 15432
rect 712 15368 968 15432
rect 1032 15368 1040 15432
rect 0 15360 1040 15368
rect 28960 15432 30000 15440
rect 28960 15368 28968 15432
rect 29032 15368 29288 15432
rect 29352 15368 29608 15432
rect 29672 15368 29928 15432
rect 29992 15368 30000 15432
rect 28960 15360 30000 15368
rect 0 15272 1040 15280
rect 0 15208 8 15272
rect 72 15208 328 15272
rect 392 15208 648 15272
rect 712 15208 968 15272
rect 1032 15208 1040 15272
rect 0 15200 1040 15208
rect 28960 15272 30000 15280
rect 28960 15208 28968 15272
rect 29032 15208 29288 15272
rect 29352 15208 29608 15272
rect 29672 15208 29928 15272
rect 29992 15208 30000 15272
rect 28960 15200 30000 15208
rect 0 15112 1040 15120
rect 0 15048 8 15112
rect 72 15048 328 15112
rect 392 15048 648 15112
rect 712 15048 968 15112
rect 1032 15048 1040 15112
rect 0 15040 1040 15048
rect 28960 15112 30000 15120
rect 28960 15048 28968 15112
rect 29032 15048 29288 15112
rect 29352 15048 29608 15112
rect 29672 15048 29928 15112
rect 29992 15048 30000 15112
rect 28960 15040 30000 15048
rect 0 14952 1040 14960
rect 0 14888 8 14952
rect 72 14888 328 14952
rect 392 14888 648 14952
rect 712 14888 968 14952
rect 1032 14888 1040 14952
rect 0 14880 1040 14888
rect 28960 14952 30000 14960
rect 28960 14888 28968 14952
rect 29032 14888 29288 14952
rect 29352 14888 29608 14952
rect 29672 14888 29928 14952
rect 29992 14888 30000 14952
rect 28960 14880 30000 14888
rect 0 14792 1040 14800
rect 0 14728 8 14792
rect 72 14728 328 14792
rect 392 14728 648 14792
rect 712 14728 968 14792
rect 1032 14728 1040 14792
rect 0 14720 1040 14728
rect 28960 14792 30000 14800
rect 28960 14728 28968 14792
rect 29032 14728 29288 14792
rect 29352 14728 29608 14792
rect 29672 14728 29928 14792
rect 29992 14728 30000 14792
rect 28960 14720 30000 14728
rect 0 14632 1040 14640
rect 0 14568 8 14632
rect 72 14568 328 14632
rect 392 14568 648 14632
rect 712 14568 968 14632
rect 1032 14568 1040 14632
rect 0 14560 1040 14568
rect 28960 14632 30000 14640
rect 28960 14568 28968 14632
rect 29032 14568 29288 14632
rect 29352 14568 29608 14632
rect 29672 14568 29928 14632
rect 29992 14568 30000 14632
rect 28960 14560 30000 14568
rect 0 14472 1040 14480
rect 0 14408 8 14472
rect 72 14408 328 14472
rect 392 14408 648 14472
rect 712 14408 968 14472
rect 1032 14408 1040 14472
rect 0 14400 1040 14408
rect 28960 14472 30000 14480
rect 28960 14408 28968 14472
rect 29032 14408 29288 14472
rect 29352 14408 29608 14472
rect 29672 14408 29928 14472
rect 29992 14408 30000 14472
rect 28960 14400 30000 14408
rect 0 14312 1040 14320
rect 0 14248 8 14312
rect 72 14248 328 14312
rect 392 14248 648 14312
rect 712 14248 968 14312
rect 1032 14248 1040 14312
rect 0 14240 1040 14248
rect 28960 14312 30000 14320
rect 28960 14248 28968 14312
rect 29032 14248 29288 14312
rect 29352 14248 29608 14312
rect 29672 14248 29928 14312
rect 29992 14248 30000 14312
rect 28960 14240 30000 14248
rect 0 14152 1040 14160
rect 0 14088 8 14152
rect 72 14088 328 14152
rect 392 14088 648 14152
rect 712 14088 968 14152
rect 1032 14088 1040 14152
rect 0 14080 1040 14088
rect 28960 14152 30000 14160
rect 28960 14088 28968 14152
rect 29032 14088 29288 14152
rect 29352 14088 29608 14152
rect 29672 14088 29928 14152
rect 29992 14088 30000 14152
rect 28960 14080 30000 14088
rect 0 13992 1040 14000
rect 0 13928 8 13992
rect 72 13928 328 13992
rect 392 13928 648 13992
rect 712 13928 968 13992
rect 1032 13928 1040 13992
rect 0 13920 1040 13928
rect 28960 13992 30000 14000
rect 28960 13928 28968 13992
rect 29032 13928 29288 13992
rect 29352 13928 29608 13992
rect 29672 13928 29928 13992
rect 29992 13928 30000 13992
rect 28960 13920 30000 13928
rect 0 13832 1040 13840
rect 0 13768 8 13832
rect 72 13768 328 13832
rect 392 13768 648 13832
rect 712 13768 968 13832
rect 1032 13768 1040 13832
rect 0 13760 1040 13768
rect 28960 13832 30000 13840
rect 28960 13768 28968 13832
rect 29032 13768 29288 13832
rect 29352 13768 29608 13832
rect 29672 13768 29928 13832
rect 29992 13768 30000 13832
rect 28960 13760 30000 13768
rect 0 13672 1040 13680
rect 0 13608 8 13672
rect 72 13608 328 13672
rect 392 13608 648 13672
rect 712 13608 968 13672
rect 1032 13608 1040 13672
rect 0 13600 1040 13608
rect 28960 13672 30000 13680
rect 28960 13608 28968 13672
rect 29032 13608 29288 13672
rect 29352 13608 29608 13672
rect 29672 13608 29928 13672
rect 29992 13608 30000 13672
rect 28960 13600 30000 13608
rect 0 13512 1040 13520
rect 0 13448 8 13512
rect 72 13448 328 13512
rect 392 13448 648 13512
rect 712 13448 968 13512
rect 1032 13448 1040 13512
rect 0 13440 1040 13448
rect 28960 13512 30000 13520
rect 28960 13448 28968 13512
rect 29032 13448 29288 13512
rect 29352 13448 29608 13512
rect 29672 13448 29928 13512
rect 29992 13448 30000 13512
rect 28960 13440 30000 13448
rect 0 13352 1040 13360
rect 0 13288 8 13352
rect 72 13288 328 13352
rect 392 13288 648 13352
rect 712 13288 968 13352
rect 1032 13288 1040 13352
rect 0 13280 1040 13288
rect 28960 13352 30000 13360
rect 28960 13288 28968 13352
rect 29032 13288 29288 13352
rect 29352 13288 29608 13352
rect 29672 13288 29928 13352
rect 29992 13288 30000 13352
rect 28960 13280 30000 13288
rect 0 13192 720 13200
rect 0 13128 8 13192
rect 72 13128 328 13192
rect 392 13128 648 13192
rect 712 13128 720 13192
rect 0 13120 720 13128
rect 800 13192 1360 13200
rect 800 13128 808 13192
rect 872 13128 1360 13192
rect 800 13120 1360 13128
rect 28960 13192 30000 13200
rect 28960 13128 28968 13192
rect 29032 13128 29288 13192
rect 29352 13128 29608 13192
rect 29672 13128 29928 13192
rect 29992 13128 30000 13192
rect 28960 13120 30000 13128
rect 0 13032 1040 13040
rect 0 12968 8 13032
rect 72 12968 328 13032
rect 392 12968 648 13032
rect 712 12968 968 13032
rect 1032 12968 1040 13032
rect 0 12960 1040 12968
rect 28960 13032 30000 13040
rect 28960 12968 28968 13032
rect 29032 12968 29288 13032
rect 29352 12968 29608 13032
rect 29672 12968 29928 13032
rect 29992 12968 30000 13032
rect 28960 12960 30000 12968
rect 0 12872 1040 12880
rect 0 12808 8 12872
rect 72 12808 328 12872
rect 392 12808 648 12872
rect 712 12808 968 12872
rect 1032 12808 1040 12872
rect 0 12800 1040 12808
rect 28960 12872 30000 12880
rect 28960 12808 28968 12872
rect 29032 12808 29288 12872
rect 29352 12808 29608 12872
rect 29672 12808 29928 12872
rect 29992 12808 30000 12872
rect 28960 12800 30000 12808
rect 0 12712 1040 12720
rect 0 12648 8 12712
rect 72 12648 328 12712
rect 392 12648 648 12712
rect 712 12648 968 12712
rect 1032 12648 1040 12712
rect 0 12640 1040 12648
rect 28960 12712 30000 12720
rect 28960 12648 28968 12712
rect 29032 12648 29288 12712
rect 29352 12648 29608 12712
rect 29672 12648 29928 12712
rect 29992 12648 30000 12712
rect 28960 12640 30000 12648
rect 0 12552 1040 12560
rect 0 12488 8 12552
rect 72 12488 328 12552
rect 392 12488 648 12552
rect 712 12488 968 12552
rect 1032 12488 1040 12552
rect 0 12480 1040 12488
rect 28960 12552 30000 12560
rect 28960 12488 28968 12552
rect 29032 12488 29288 12552
rect 29352 12488 29608 12552
rect 29672 12488 29928 12552
rect 29992 12488 30000 12552
rect 28960 12480 30000 12488
rect 0 12392 1040 12400
rect 0 12328 8 12392
rect 72 12328 328 12392
rect 392 12328 648 12392
rect 712 12328 968 12392
rect 1032 12328 1040 12392
rect 0 12320 1040 12328
rect 28960 12392 30000 12400
rect 28960 12328 28968 12392
rect 29032 12328 29288 12392
rect 29352 12328 29608 12392
rect 29672 12328 29928 12392
rect 29992 12328 30000 12392
rect 28960 12320 30000 12328
rect 0 12232 1040 12240
rect 0 12168 8 12232
rect 72 12168 328 12232
rect 392 12168 648 12232
rect 712 12168 968 12232
rect 1032 12168 1040 12232
rect 0 12160 1040 12168
rect 28960 12232 30000 12240
rect 28960 12168 28968 12232
rect 29032 12168 29288 12232
rect 29352 12168 29608 12232
rect 29672 12168 29928 12232
rect 29992 12168 30000 12232
rect 28960 12160 30000 12168
rect 0 12072 1040 12080
rect 0 12008 8 12072
rect 72 12008 328 12072
rect 392 12008 648 12072
rect 712 12008 968 12072
rect 1032 12008 1040 12072
rect 0 12000 1040 12008
rect 28960 12072 30000 12080
rect 28960 12008 28968 12072
rect 29032 12008 29288 12072
rect 29352 12008 29608 12072
rect 29672 12008 29928 12072
rect 29992 12008 30000 12072
rect 28960 12000 30000 12008
rect 0 11912 1040 11920
rect 0 11848 8 11912
rect 72 11848 328 11912
rect 392 11848 648 11912
rect 712 11848 968 11912
rect 1032 11848 1040 11912
rect 0 11840 1040 11848
rect 28960 11912 30000 11920
rect 28960 11848 28968 11912
rect 29032 11848 29288 11912
rect 29352 11848 29608 11912
rect 29672 11848 29928 11912
rect 29992 11848 30000 11912
rect 28960 11840 30000 11848
rect 0 11752 1040 11760
rect 0 11688 8 11752
rect 72 11688 328 11752
rect 392 11688 648 11752
rect 712 11688 968 11752
rect 1032 11688 1040 11752
rect 0 11680 1040 11688
rect 28960 11752 30000 11760
rect 28960 11688 28968 11752
rect 29032 11688 29288 11752
rect 29352 11688 29608 11752
rect 29672 11688 29928 11752
rect 29992 11688 30000 11752
rect 28960 11680 30000 11688
rect 0 11592 1040 11600
rect 0 11528 8 11592
rect 72 11528 328 11592
rect 392 11528 648 11592
rect 712 11528 968 11592
rect 1032 11528 1040 11592
rect 0 11520 1040 11528
rect 28960 11592 30000 11600
rect 28960 11528 28968 11592
rect 29032 11528 29288 11592
rect 29352 11528 29608 11592
rect 29672 11528 29928 11592
rect 29992 11528 30000 11592
rect 28960 11520 30000 11528
rect 0 11432 1040 11440
rect 0 11368 8 11432
rect 72 11368 328 11432
rect 392 11368 648 11432
rect 712 11368 968 11432
rect 1032 11368 1040 11432
rect 0 11360 1040 11368
rect 28960 11432 30000 11440
rect 28960 11368 28968 11432
rect 29032 11368 29288 11432
rect 29352 11368 29608 11432
rect 29672 11368 29928 11432
rect 29992 11368 30000 11432
rect 28960 11360 30000 11368
rect 0 11272 1040 11280
rect 0 11208 8 11272
rect 72 11208 328 11272
rect 392 11208 648 11272
rect 712 11208 968 11272
rect 1032 11208 1040 11272
rect 0 11200 1040 11208
rect 28960 11272 30000 11280
rect 28960 11208 28968 11272
rect 29032 11208 29288 11272
rect 29352 11208 29608 11272
rect 29672 11208 29928 11272
rect 29992 11208 30000 11272
rect 28960 11200 30000 11208
rect 0 11112 1040 11120
rect 0 11048 8 11112
rect 72 11048 328 11112
rect 392 11048 648 11112
rect 712 11048 968 11112
rect 1032 11048 1040 11112
rect 0 11040 1040 11048
rect 28960 11112 30000 11120
rect 28960 11048 28968 11112
rect 29032 11048 29288 11112
rect 29352 11048 29608 11112
rect 29672 11048 29928 11112
rect 29992 11048 30000 11112
rect 28960 11040 30000 11048
rect 0 10952 1040 10960
rect 0 10888 8 10952
rect 72 10888 328 10952
rect 392 10888 648 10952
rect 712 10888 968 10952
rect 1032 10888 1040 10952
rect 0 10880 1040 10888
rect 28960 10952 30000 10960
rect 28960 10888 28968 10952
rect 29032 10888 29288 10952
rect 29352 10888 29608 10952
rect 29672 10888 29928 10952
rect 29992 10888 30000 10952
rect 28960 10880 30000 10888
rect 0 10792 1360 10800
rect 0 10728 8 10792
rect 72 10728 328 10792
rect 392 10728 648 10792
rect 712 10728 968 10792
rect 1032 10728 1360 10792
rect 0 10720 1360 10728
rect 28640 10792 30000 10800
rect 28640 10728 28968 10792
rect 29032 10728 29288 10792
rect 29352 10728 29608 10792
rect 29672 10728 29928 10792
rect 29992 10728 30000 10792
rect 28640 10720 30000 10728
rect 0 10632 400 10640
rect 0 10568 8 10632
rect 72 10568 328 10632
rect 392 10568 400 10632
rect 0 10560 400 10568
rect 480 10632 1360 10640
rect 480 10568 488 10632
rect 552 10568 1360 10632
rect 480 10560 1360 10568
rect 28960 10632 30000 10640
rect 28960 10568 28968 10632
rect 29032 10568 29288 10632
rect 29352 10568 29608 10632
rect 29672 10568 29928 10632
rect 29992 10568 30000 10632
rect 28960 10560 30000 10568
rect 0 10472 1360 10480
rect 0 10408 8 10472
rect 72 10408 328 10472
rect 392 10408 648 10472
rect 712 10408 968 10472
rect 1032 10408 1360 10472
rect 0 10400 1360 10408
rect 28640 10472 30000 10480
rect 28640 10408 28968 10472
rect 29032 10408 29288 10472
rect 29352 10408 29608 10472
rect 29672 10408 29928 10472
rect 29992 10408 30000 10472
rect 28640 10400 30000 10408
rect 160 10312 1360 10320
rect 160 10248 168 10312
rect 232 10248 1360 10312
rect 160 10240 1360 10248
rect 28960 10312 30000 10320
rect 28960 10248 28968 10312
rect 29032 10248 29288 10312
rect 29352 10248 29608 10312
rect 29672 10248 29928 10312
rect 29992 10248 30000 10312
rect 28960 10240 30000 10248
rect 0 10152 1360 10160
rect 0 10088 8 10152
rect 72 10088 328 10152
rect 392 10088 648 10152
rect 712 10088 968 10152
rect 1032 10088 1360 10152
rect 0 10080 1360 10088
rect 28640 10152 30000 10160
rect 28640 10088 28968 10152
rect 29032 10088 29288 10152
rect 29352 10088 29608 10152
rect 29672 10088 29928 10152
rect 29992 10088 30000 10152
rect 28640 10080 30000 10088
rect 0 9992 1040 10000
rect 0 9928 8 9992
rect 72 9928 328 9992
rect 392 9928 648 9992
rect 712 9928 968 9992
rect 1032 9928 1040 9992
rect 0 9920 1040 9928
rect 28960 9992 30000 10000
rect 28960 9928 28968 9992
rect 29032 9928 29288 9992
rect 29352 9928 29608 9992
rect 29672 9928 29928 9992
rect 29992 9928 30000 9992
rect 28960 9920 30000 9928
rect 0 9832 1040 9840
rect 0 9768 8 9832
rect 72 9768 328 9832
rect 392 9768 648 9832
rect 712 9768 968 9832
rect 1032 9768 1040 9832
rect 0 9760 1040 9768
rect 28960 9832 30000 9840
rect 28960 9768 28968 9832
rect 29032 9768 29288 9832
rect 29352 9768 29608 9832
rect 29672 9768 29928 9832
rect 29992 9768 30000 9832
rect 28960 9760 30000 9768
rect 0 9672 1360 9680
rect 0 9608 8 9672
rect 72 9608 328 9672
rect 392 9608 648 9672
rect 712 9608 968 9672
rect 1032 9608 1360 9672
rect 0 9600 1360 9608
rect 28640 9672 30000 9680
rect 28640 9608 28968 9672
rect 29032 9608 29288 9672
rect 29352 9608 29608 9672
rect 29672 9608 29928 9672
rect 29992 9608 30000 9672
rect 28640 9600 30000 9608
rect 0 9512 1040 9520
rect 0 9448 8 9512
rect 72 9448 328 9512
rect 392 9448 648 9512
rect 712 9448 968 9512
rect 1032 9448 1040 9512
rect 0 9440 1040 9448
rect 28640 9512 30000 9520
rect 28640 9448 29768 9512
rect 29832 9448 30000 9512
rect 28640 9440 30000 9448
rect 0 9352 1360 9360
rect 0 9288 8 9352
rect 72 9288 328 9352
rect 392 9288 648 9352
rect 712 9288 968 9352
rect 1032 9288 1360 9352
rect 0 9280 1360 9288
rect 28640 9352 30000 9360
rect 28640 9288 28968 9352
rect 29032 9288 29288 9352
rect 29352 9288 29608 9352
rect 29672 9288 29928 9352
rect 29992 9288 30000 9352
rect 28640 9280 30000 9288
rect 0 9192 1040 9200
rect 0 9128 8 9192
rect 72 9128 328 9192
rect 392 9128 648 9192
rect 712 9128 968 9192
rect 1032 9128 1040 9192
rect 0 9120 1040 9128
rect 28640 9192 29520 9200
rect 28640 9128 29448 9192
rect 29512 9128 29520 9192
rect 28640 9120 29520 9128
rect 29600 9192 30000 9200
rect 29600 9128 29608 9192
rect 29672 9128 29928 9192
rect 29992 9128 30000 9192
rect 29600 9120 30000 9128
rect 0 9032 1360 9040
rect 0 8968 8 9032
rect 72 8968 328 9032
rect 392 8968 648 9032
rect 712 8968 968 9032
rect 1032 8968 1360 9032
rect 0 8960 1360 8968
rect 28640 9032 30000 9040
rect 28640 8968 28968 9032
rect 29032 8968 29288 9032
rect 29352 8968 29608 9032
rect 29672 8968 29928 9032
rect 29992 8968 30000 9032
rect 28640 8960 30000 8968
rect 0 8872 1040 8880
rect 0 8808 8 8872
rect 72 8808 328 8872
rect 392 8808 648 8872
rect 712 8808 968 8872
rect 1032 8808 1040 8872
rect 0 8800 1040 8808
rect 28960 8872 30000 8880
rect 28960 8808 28968 8872
rect 29032 8808 29288 8872
rect 29352 8808 29608 8872
rect 29672 8808 29928 8872
rect 29992 8808 30000 8872
rect 28960 8800 30000 8808
rect 0 8712 1040 8720
rect 0 8648 8 8712
rect 72 8648 328 8712
rect 392 8648 648 8712
rect 712 8648 968 8712
rect 1032 8648 1040 8712
rect 0 8640 1040 8648
rect 28960 8712 30000 8720
rect 28960 8648 28968 8712
rect 29032 8648 29288 8712
rect 29352 8648 29608 8712
rect 29672 8648 29928 8712
rect 29992 8648 30000 8712
rect 28960 8640 30000 8648
rect 0 8552 1040 8560
rect 0 8488 8 8552
rect 72 8488 328 8552
rect 392 8488 648 8552
rect 712 8488 968 8552
rect 1032 8488 1040 8552
rect 0 8480 1040 8488
rect 28960 8552 30000 8560
rect 28960 8488 28968 8552
rect 29032 8488 29288 8552
rect 29352 8488 29608 8552
rect 29672 8488 29928 8552
rect 29992 8488 30000 8552
rect 28960 8480 30000 8488
rect 0 8392 1040 8400
rect 0 8328 8 8392
rect 72 8328 328 8392
rect 392 8328 648 8392
rect 712 8328 968 8392
rect 1032 8328 1040 8392
rect 0 8320 1040 8328
rect 28960 8392 30000 8400
rect 28960 8328 28968 8392
rect 29032 8328 29288 8392
rect 29352 8328 29608 8392
rect 29672 8328 29928 8392
rect 29992 8328 30000 8392
rect 28960 8320 30000 8328
rect 0 8232 1040 8240
rect 0 8168 8 8232
rect 72 8168 328 8232
rect 392 8168 648 8232
rect 712 8168 968 8232
rect 1032 8168 1040 8232
rect 0 8160 1040 8168
rect 28960 8232 30000 8240
rect 28960 8168 28968 8232
rect 29032 8168 29288 8232
rect 29352 8168 29608 8232
rect 29672 8168 29928 8232
rect 29992 8168 30000 8232
rect 28960 8160 30000 8168
rect 0 8072 1040 8080
rect 0 8008 8 8072
rect 72 8008 328 8072
rect 392 8008 648 8072
rect 712 8008 968 8072
rect 1032 8008 1040 8072
rect 0 8000 1040 8008
rect 28960 8072 30000 8080
rect 28960 8008 28968 8072
rect 29032 8008 29288 8072
rect 29352 8008 29608 8072
rect 29672 8008 29928 8072
rect 29992 8008 30000 8072
rect 28960 8000 30000 8008
rect 0 7912 1040 7920
rect 0 7848 8 7912
rect 72 7848 328 7912
rect 392 7848 648 7912
rect 712 7848 968 7912
rect 1032 7848 1040 7912
rect 0 7840 1040 7848
rect 28960 7912 30000 7920
rect 28960 7848 28968 7912
rect 29032 7848 29288 7912
rect 29352 7848 29608 7912
rect 29672 7848 29928 7912
rect 29992 7848 30000 7912
rect 28960 7840 30000 7848
rect 0 7752 1040 7760
rect 0 7688 8 7752
rect 72 7688 328 7752
rect 392 7688 648 7752
rect 712 7688 968 7752
rect 1032 7688 1040 7752
rect 0 7680 1040 7688
rect 28960 7752 30000 7760
rect 28960 7688 28968 7752
rect 29032 7688 29288 7752
rect 29352 7688 29608 7752
rect 29672 7688 29928 7752
rect 29992 7688 30000 7752
rect 28960 7680 30000 7688
rect 0 7592 1040 7600
rect 0 7528 8 7592
rect 72 7528 328 7592
rect 392 7528 648 7592
rect 712 7528 968 7592
rect 1032 7528 1040 7592
rect 0 7520 1040 7528
rect 28960 7592 30000 7600
rect 28960 7528 28968 7592
rect 29032 7528 29288 7592
rect 29352 7528 29608 7592
rect 29672 7528 29928 7592
rect 29992 7528 30000 7592
rect 28960 7520 30000 7528
rect 0 7432 1040 7440
rect 0 7368 8 7432
rect 72 7368 328 7432
rect 392 7368 648 7432
rect 712 7368 968 7432
rect 1032 7368 1040 7432
rect 0 7360 1040 7368
rect 28960 7432 30000 7440
rect 28960 7368 28968 7432
rect 29032 7368 29288 7432
rect 29352 7368 29608 7432
rect 29672 7368 29928 7432
rect 29992 7368 30000 7432
rect 28960 7360 30000 7368
rect 0 7272 1040 7280
rect 0 7208 8 7272
rect 72 7208 328 7272
rect 392 7208 648 7272
rect 712 7208 968 7272
rect 1032 7208 1040 7272
rect 0 7200 1040 7208
rect 28960 7272 30000 7280
rect 28960 7208 28968 7272
rect 29032 7208 29288 7272
rect 29352 7208 29608 7272
rect 29672 7208 29928 7272
rect 29992 7208 30000 7272
rect 28960 7200 30000 7208
rect 0 7112 1040 7120
rect 0 7048 8 7112
rect 72 7048 328 7112
rect 392 7048 648 7112
rect 712 7048 968 7112
rect 1032 7048 1040 7112
rect 0 7040 1040 7048
rect 28960 7112 30000 7120
rect 28960 7048 28968 7112
rect 29032 7048 29288 7112
rect 29352 7048 29608 7112
rect 29672 7048 29928 7112
rect 29992 7048 30000 7112
rect 28960 7040 30000 7048
rect 0 6952 1040 6960
rect 0 6888 8 6952
rect 72 6888 328 6952
rect 392 6888 648 6952
rect 712 6888 968 6952
rect 1032 6888 1040 6952
rect 0 6880 1040 6888
rect 28960 6952 30000 6960
rect 28960 6888 28968 6952
rect 29032 6888 29288 6952
rect 29352 6888 29608 6952
rect 29672 6888 29928 6952
rect 29992 6888 30000 6952
rect 28960 6880 30000 6888
rect 0 6792 1040 6800
rect 0 6728 8 6792
rect 72 6728 328 6792
rect 392 6728 648 6792
rect 712 6728 968 6792
rect 1032 6728 1040 6792
rect 0 6720 1040 6728
rect 28960 6792 30000 6800
rect 28960 6728 28968 6792
rect 29032 6728 29288 6792
rect 29352 6728 29608 6792
rect 29672 6728 29928 6792
rect 29992 6728 30000 6792
rect 28960 6720 30000 6728
rect 0 6632 1040 6640
rect 0 6568 8 6632
rect 72 6568 328 6632
rect 392 6568 648 6632
rect 712 6568 968 6632
rect 1032 6568 1040 6632
rect 0 6560 1040 6568
rect 28640 6632 29200 6640
rect 28640 6568 29128 6632
rect 29192 6568 29200 6632
rect 28640 6560 29200 6568
rect 29280 6632 30000 6640
rect 29280 6568 29288 6632
rect 29352 6568 29608 6632
rect 29672 6568 29928 6632
rect 29992 6568 30000 6632
rect 29280 6560 30000 6568
rect 0 6472 1040 6480
rect 0 6408 8 6472
rect 72 6408 328 6472
rect 392 6408 648 6472
rect 712 6408 968 6472
rect 1032 6408 1040 6472
rect 0 6400 1040 6408
rect 28960 6472 30000 6480
rect 28960 6408 28968 6472
rect 29032 6408 29288 6472
rect 29352 6408 29608 6472
rect 29672 6408 29928 6472
rect 29992 6408 30000 6472
rect 28960 6400 30000 6408
rect 0 6312 1040 6320
rect 0 6248 8 6312
rect 72 6248 328 6312
rect 392 6248 648 6312
rect 712 6248 968 6312
rect 1032 6248 1040 6312
rect 0 6240 1040 6248
rect 28960 6312 30000 6320
rect 28960 6248 28968 6312
rect 29032 6248 29288 6312
rect 29352 6248 29608 6312
rect 29672 6248 29928 6312
rect 29992 6248 30000 6312
rect 28960 6240 30000 6248
rect 0 6152 1040 6160
rect 0 6088 8 6152
rect 72 6088 328 6152
rect 392 6088 648 6152
rect 712 6088 968 6152
rect 1032 6088 1040 6152
rect 0 6080 1040 6088
rect 28960 6152 30000 6160
rect 28960 6088 28968 6152
rect 29032 6088 29288 6152
rect 29352 6088 29608 6152
rect 29672 6088 29928 6152
rect 29992 6088 30000 6152
rect 28960 6080 30000 6088
rect 0 5992 1040 6000
rect 0 5928 8 5992
rect 72 5928 328 5992
rect 392 5928 648 5992
rect 712 5928 968 5992
rect 1032 5928 1040 5992
rect 0 5920 1040 5928
rect 28960 5992 30000 6000
rect 28960 5928 28968 5992
rect 29032 5928 29288 5992
rect 29352 5928 29608 5992
rect 29672 5928 29928 5992
rect 29992 5928 30000 5992
rect 28960 5920 30000 5928
rect 0 5832 1040 5840
rect 0 5768 8 5832
rect 72 5768 328 5832
rect 392 5768 648 5832
rect 712 5768 968 5832
rect 1032 5768 1040 5832
rect 0 5760 1040 5768
rect 28960 5832 30000 5840
rect 28960 5768 28968 5832
rect 29032 5768 29288 5832
rect 29352 5768 29608 5832
rect 29672 5768 29928 5832
rect 29992 5768 30000 5832
rect 28960 5760 30000 5768
rect 0 5672 1040 5680
rect 0 5608 8 5672
rect 72 5608 328 5672
rect 392 5608 648 5672
rect 712 5608 968 5672
rect 1032 5608 1040 5672
rect 0 5600 1040 5608
rect 28960 5672 30000 5680
rect 28960 5608 28968 5672
rect 29032 5608 29288 5672
rect 29352 5608 29608 5672
rect 29672 5608 29928 5672
rect 29992 5608 30000 5672
rect 28960 5600 30000 5608
rect 0 5512 1040 5520
rect 0 5448 8 5512
rect 72 5448 328 5512
rect 392 5448 648 5512
rect 712 5448 968 5512
rect 1032 5448 1040 5512
rect 0 5440 1040 5448
rect 28960 5512 30000 5520
rect 28960 5448 28968 5512
rect 29032 5448 29288 5512
rect 29352 5448 29608 5512
rect 29672 5448 29928 5512
rect 29992 5448 30000 5512
rect 28960 5440 30000 5448
rect 0 5352 1040 5360
rect 0 5288 8 5352
rect 72 5288 328 5352
rect 392 5288 648 5352
rect 712 5288 968 5352
rect 1032 5288 1040 5352
rect 0 5280 1040 5288
rect 28960 5352 30000 5360
rect 28960 5288 28968 5352
rect 29032 5288 29288 5352
rect 29352 5288 29608 5352
rect 29672 5288 29928 5352
rect 29992 5288 30000 5352
rect 28960 5280 30000 5288
rect 0 5192 1040 5200
rect 0 5128 8 5192
rect 72 5128 328 5192
rect 392 5128 648 5192
rect 712 5128 968 5192
rect 1032 5128 1040 5192
rect 0 5120 1040 5128
rect 28960 5192 30000 5200
rect 28960 5128 28968 5192
rect 29032 5128 29288 5192
rect 29352 5128 29608 5192
rect 29672 5128 29928 5192
rect 29992 5128 30000 5192
rect 28960 5120 30000 5128
rect 0 5032 1040 5040
rect 0 4968 8 5032
rect 72 4968 328 5032
rect 392 4968 648 5032
rect 712 4968 968 5032
rect 1032 4968 1040 5032
rect 0 4960 1040 4968
rect 28960 5032 30000 5040
rect 28960 4968 28968 5032
rect 29032 4968 29288 5032
rect 29352 4968 29608 5032
rect 29672 4968 29928 5032
rect 29992 4968 30000 5032
rect 28960 4960 30000 4968
rect 0 4872 1040 4880
rect 0 4808 8 4872
rect 72 4808 328 4872
rect 392 4808 648 4872
rect 712 4808 968 4872
rect 1032 4808 1040 4872
rect 0 4800 1040 4808
rect 28960 4872 30000 4880
rect 28960 4808 28968 4872
rect 29032 4808 29288 4872
rect 29352 4808 29608 4872
rect 29672 4808 29928 4872
rect 29992 4808 30000 4872
rect 28960 4800 30000 4808
rect 0 4712 1040 4720
rect 0 4648 8 4712
rect 72 4648 328 4712
rect 392 4648 648 4712
rect 712 4648 968 4712
rect 1032 4648 1040 4712
rect 0 4640 1040 4648
rect 28960 4712 30000 4720
rect 28960 4648 28968 4712
rect 29032 4648 29288 4712
rect 29352 4648 29608 4712
rect 29672 4648 29928 4712
rect 29992 4648 30000 4712
rect 28960 4640 30000 4648
rect 0 4552 1040 4560
rect 0 4488 8 4552
rect 72 4488 328 4552
rect 392 4488 648 4552
rect 712 4488 968 4552
rect 1032 4488 1040 4552
rect 0 4480 1040 4488
rect 28960 4552 30000 4560
rect 28960 4488 28968 4552
rect 29032 4488 29288 4552
rect 29352 4488 29608 4552
rect 29672 4488 29928 4552
rect 29992 4488 30000 4552
rect 28960 4480 30000 4488
rect 0 4392 1040 4400
rect 0 4328 8 4392
rect 72 4328 328 4392
rect 392 4328 648 4392
rect 712 4328 968 4392
rect 1032 4328 1040 4392
rect 0 4320 1040 4328
rect 28960 4392 30000 4400
rect 28960 4328 28968 4392
rect 29032 4328 29288 4392
rect 29352 4328 29608 4392
rect 29672 4328 29928 4392
rect 29992 4328 30000 4392
rect 28960 4320 30000 4328
rect 0 4232 1360 4240
rect 0 4168 8 4232
rect 72 4168 328 4232
rect 392 4168 648 4232
rect 712 4168 968 4232
rect 1032 4168 1360 4232
rect 0 4160 1360 4168
rect 28720 4232 30000 4240
rect 28720 4168 28968 4232
rect 29032 4168 29288 4232
rect 29352 4168 29608 4232
rect 29672 4168 29928 4232
rect 29992 4168 30000 4232
rect 28720 4160 30000 4168
rect 0 4072 1040 4080
rect 0 4008 8 4072
rect 72 4008 328 4072
rect 392 4008 648 4072
rect 712 4008 968 4072
rect 1032 4008 1040 4072
rect 0 4000 1040 4008
rect 28640 4072 29520 4080
rect 28640 4008 29448 4072
rect 29512 4008 29520 4072
rect 28640 4000 29520 4008
rect 29600 4072 30000 4080
rect 29600 4008 29608 4072
rect 29672 4008 29928 4072
rect 29992 4008 30000 4072
rect 29600 4000 30000 4008
rect 0 3912 1360 3920
rect 0 3848 8 3912
rect 72 3848 328 3912
rect 392 3848 648 3912
rect 712 3848 968 3912
rect 1032 3848 1360 3912
rect 0 3840 1360 3848
rect 28640 3912 30000 3920
rect 28640 3848 28968 3912
rect 29032 3848 29288 3912
rect 29352 3848 29608 3912
rect 29672 3848 29928 3912
rect 29992 3848 30000 3912
rect 28640 3840 30000 3848
rect 0 3752 1040 3760
rect 0 3688 8 3752
rect 72 3688 328 3752
rect 392 3688 648 3752
rect 712 3688 968 3752
rect 1032 3688 1040 3752
rect 0 3680 1040 3688
rect 28640 3752 30000 3760
rect 28640 3688 29768 3752
rect 29832 3688 30000 3752
rect 28640 3680 30000 3688
rect 0 3592 1360 3600
rect 0 3528 8 3592
rect 72 3528 328 3592
rect 392 3528 648 3592
rect 712 3528 968 3592
rect 1032 3528 1360 3592
rect 0 3520 1360 3528
rect 28640 3592 30000 3600
rect 28640 3528 28968 3592
rect 29032 3528 29288 3592
rect 29352 3528 29608 3592
rect 29672 3528 29928 3592
rect 29992 3528 30000 3592
rect 28640 3520 30000 3528
rect 0 3432 1040 3440
rect 0 3368 8 3432
rect 72 3368 328 3432
rect 392 3368 648 3432
rect 712 3368 968 3432
rect 1032 3368 1040 3432
rect 0 3360 1040 3368
rect 28960 3432 30000 3440
rect 28960 3368 28968 3432
rect 29032 3368 29288 3432
rect 29352 3368 29608 3432
rect 29672 3368 29928 3432
rect 29992 3368 30000 3432
rect 28960 3360 30000 3368
rect 0 3272 1040 3280
rect 0 3208 8 3272
rect 72 3208 328 3272
rect 392 3208 648 3272
rect 712 3208 968 3272
rect 1032 3208 1040 3272
rect 0 3200 1040 3208
rect 28960 3272 30000 3280
rect 28960 3208 28968 3272
rect 29032 3208 29288 3272
rect 29352 3208 29608 3272
rect 29672 3208 29928 3272
rect 29992 3208 30000 3272
rect 28960 3200 30000 3208
rect 0 3112 1360 3120
rect 0 3048 8 3112
rect 72 3048 328 3112
rect 392 3048 648 3112
rect 712 3048 968 3112
rect 1032 3048 1360 3112
rect 0 3040 1360 3048
rect 28640 3112 30000 3120
rect 28640 3048 28968 3112
rect 29032 3048 29288 3112
rect 29352 3048 29608 3112
rect 29672 3048 29928 3112
rect 29992 3048 30000 3112
rect 28640 3040 30000 3048
rect 0 2952 1360 2960
rect 0 2888 8 2952
rect 72 2888 328 2952
rect 392 2888 648 2952
rect 712 2888 968 2952
rect 1032 2888 1360 2952
rect 0 2880 1360 2888
rect 28640 2952 30000 2960
rect 28640 2888 28968 2952
rect 29032 2888 29288 2952
rect 29352 2888 29608 2952
rect 29672 2888 29928 2952
rect 29992 2888 30000 2952
rect 28640 2880 30000 2888
rect 0 2792 1360 2800
rect 0 2728 8 2792
rect 72 2728 328 2792
rect 392 2728 648 2792
rect 712 2728 968 2792
rect 1032 2728 1360 2792
rect 0 2720 1360 2728
rect 28640 2792 30000 2800
rect 28640 2728 28968 2792
rect 29032 2728 29288 2792
rect 29352 2728 29608 2792
rect 29672 2728 29928 2792
rect 29992 2728 30000 2792
rect 28640 2720 30000 2728
rect 0 2632 1360 2640
rect 0 2568 8 2632
rect 72 2568 328 2632
rect 392 2568 648 2632
rect 712 2568 968 2632
rect 1032 2568 1360 2632
rect 0 2560 1360 2568
rect 28640 2632 30000 2640
rect 28640 2568 28968 2632
rect 29032 2568 29288 2632
rect 29352 2568 29608 2632
rect 29672 2568 29928 2632
rect 29992 2568 30000 2632
rect 28640 2560 30000 2568
rect 0 2472 1360 2480
rect 0 2408 8 2472
rect 72 2408 328 2472
rect 392 2408 648 2472
rect 712 2408 968 2472
rect 1032 2408 1360 2472
rect 0 2400 1360 2408
rect 28640 2472 30000 2480
rect 28640 2408 28968 2472
rect 29032 2408 29288 2472
rect 29352 2408 29608 2472
rect 29672 2408 29928 2472
rect 29992 2408 30000 2472
rect 28640 2400 30000 2408
rect 0 2312 1040 2320
rect 0 2248 8 2312
rect 72 2248 328 2312
rect 392 2248 648 2312
rect 712 2248 968 2312
rect 1032 2248 1040 2312
rect 0 2240 1040 2248
rect 28960 2312 30000 2320
rect 28960 2248 28968 2312
rect 29032 2248 29288 2312
rect 29352 2248 29608 2312
rect 29672 2248 29928 2312
rect 29992 2248 30000 2312
rect 28960 2240 30000 2248
rect 0 2152 1040 2160
rect 0 2088 8 2152
rect 72 2088 328 2152
rect 392 2088 648 2152
rect 712 2088 968 2152
rect 1032 2088 1040 2152
rect 0 2080 1040 2088
rect 28960 2152 30000 2160
rect 28960 2088 28968 2152
rect 29032 2088 29288 2152
rect 29352 2088 29608 2152
rect 29672 2088 29928 2152
rect 29992 2088 30000 2152
rect 28960 2080 30000 2088
rect 0 1992 1040 2000
rect 0 1928 8 1992
rect 72 1928 328 1992
rect 392 1928 648 1992
rect 712 1928 968 1992
rect 1032 1928 1040 1992
rect 0 1920 1040 1928
rect 28960 1992 30000 2000
rect 28960 1928 28968 1992
rect 29032 1928 29288 1992
rect 29352 1928 29608 1992
rect 29672 1928 29928 1992
rect 29992 1928 30000 1992
rect 28960 1920 30000 1928
rect 0 1832 1360 1840
rect 0 1768 8 1832
rect 72 1768 328 1832
rect 392 1768 648 1832
rect 712 1768 968 1832
rect 1032 1768 1360 1832
rect 0 1760 1360 1768
rect 28640 1832 30000 1840
rect 28640 1768 28968 1832
rect 29032 1768 29288 1832
rect 29352 1768 29608 1832
rect 29672 1768 29928 1832
rect 29992 1768 30000 1832
rect 28640 1760 30000 1768
rect 0 1672 1360 1680
rect 0 1608 8 1672
rect 72 1608 328 1672
rect 392 1608 648 1672
rect 712 1608 968 1672
rect 1032 1608 1360 1672
rect 0 1600 1360 1608
rect 28640 1672 30000 1680
rect 28640 1608 28968 1672
rect 29032 1608 29288 1672
rect 29352 1608 29608 1672
rect 29672 1608 29928 1672
rect 29992 1608 30000 1672
rect 28640 1600 30000 1608
rect 0 1512 1360 1520
rect 0 1448 8 1512
rect 72 1448 328 1512
rect 392 1448 648 1512
rect 712 1448 968 1512
rect 1032 1448 1360 1512
rect 0 1440 1360 1448
rect 28640 1512 30000 1520
rect 28640 1448 28968 1512
rect 29032 1448 29288 1512
rect 29352 1448 29608 1512
rect 29672 1448 29928 1512
rect 29992 1448 30000 1512
rect 28640 1440 30000 1448
rect 0 1352 1360 1360
rect 0 1288 8 1352
rect 72 1288 328 1352
rect 392 1288 648 1352
rect 712 1288 968 1352
rect 1032 1288 1360 1352
rect 0 1280 1360 1288
rect 28640 1352 30000 1360
rect 28640 1288 28968 1352
rect 29032 1288 29288 1352
rect 29352 1288 29608 1352
rect 29672 1288 29928 1352
rect 29992 1288 30000 1352
rect 28640 1280 30000 1288
rect 0 1192 1360 1200
rect 0 1128 8 1192
rect 72 1128 328 1192
rect 392 1128 648 1192
rect 712 1128 968 1192
rect 1032 1128 1360 1192
rect 0 1120 1360 1128
rect 28640 1192 30000 1200
rect 28640 1128 28968 1192
rect 29032 1128 29288 1192
rect 29352 1128 29608 1192
rect 29672 1128 29928 1192
rect 29992 1128 30000 1192
rect 28640 1120 30000 1128
rect 0 1032 1040 1040
rect 0 968 8 1032
rect 72 968 328 1032
rect 392 968 648 1032
rect 712 968 968 1032
rect 1032 968 1040 1032
rect 0 960 1040 968
rect 28960 1032 30000 1040
rect 28960 968 28968 1032
rect 29032 968 29288 1032
rect 29352 968 29608 1032
rect 29672 968 29928 1032
rect 29992 968 30000 1032
rect 28960 960 30000 968
rect 0 872 30000 880
rect 0 808 8 872
rect 72 808 328 872
rect 392 808 648 872
rect 712 808 968 872
rect 1032 808 28968 872
rect 29032 808 29288 872
rect 29352 808 29608 872
rect 29672 808 29928 872
rect 29992 808 30000 872
rect 0 792 30000 808
rect 0 728 8 792
rect 72 728 328 792
rect 392 728 648 792
rect 712 728 968 792
rect 1032 728 28968 792
rect 29032 728 29288 792
rect 29352 728 29608 792
rect 29672 728 29928 792
rect 29992 728 30000 792
rect 0 712 30000 728
rect 0 648 8 712
rect 72 648 328 712
rect 392 648 648 712
rect 712 648 968 712
rect 1032 648 28968 712
rect 29032 648 29288 712
rect 29352 648 29608 712
rect 29672 648 29928 712
rect 29992 648 30000 712
rect 0 632 30000 648
rect 0 568 8 632
rect 72 568 328 632
rect 392 568 648 632
rect 712 568 968 632
rect 1032 568 28968 632
rect 29032 568 29288 632
rect 29352 568 29608 632
rect 29672 568 29928 632
rect 29992 568 30000 632
rect 0 552 30000 568
rect 0 488 8 552
rect 72 488 328 552
rect 392 488 648 552
rect 712 488 968 552
rect 1032 488 28968 552
rect 29032 488 29288 552
rect 29352 488 29608 552
rect 29672 488 29928 552
rect 29992 488 30000 552
rect 0 480 30000 488
rect 0 392 30000 400
rect 0 328 1128 392
rect 1192 328 28808 392
rect 28872 328 30000 392
rect 0 312 30000 328
rect 0 248 1128 312
rect 1192 248 28808 312
rect 28872 248 30000 312
rect 0 232 30000 248
rect 0 168 1128 232
rect 1192 168 28808 232
rect 28872 168 30000 232
rect 0 152 30000 168
rect 0 88 1128 152
rect 1192 88 28808 152
rect 28872 88 30000 152
rect 0 72 30000 88
rect 0 8 1128 72
rect 1192 8 28808 72
rect 28872 8 30000 72
rect 0 0 30000 8
use cap1_10_core  p2
timestamp 1638148091
transform 1 0 14000 0 1 2000
box -12906 1334 14906 7866
use cap1_10_core  m2
timestamp 1638148091
transform 1 0 14000 0 1 8560
box -12906 1334 14906 7866
use cap1_10_core  m1
timestamp 1638148091
transform 1 0 14000 0 1 15120
box -12906 1334 14906 7866
use cap1_10_core  p1
timestamp 1638148091
transform 1 0 14000 0 1 21680
box -12906 1334 14906 7866
use cap1_10_dummy  dummy1
timestamp 1638148091
transform 1 0 14000 0 1 28240
box -12906 1334 14906 3706
use cap1_10_dummy  dummy2
timestamp 1638148091
transform 1 0 14000 0 1 -400
box -12906 1334 14906 3706
<< labels >>
rlabel metal3 s 29760 31840 29840 31920 4 ip
port 1 nsew
rlabel metal3 s 29120 31840 29200 31920 4 xp
port 2 nsew
rlabel metal3 s 29440 31840 29520 31920 4 om
port 3 nsew
rlabel metal3 s 160 31840 240 31920 4 im
port 4 nsew
rlabel metal3 s 800 31840 880 31920 4 xm
port 5 nsew
rlabel metal3 s 480 31840 560 31920 4 op
port 6 nsew
rlabel metal4 s 0 480 80 880 4 gnda
port 7 nsew
rlabel metal4 s 0 0 80 400 4 vssa
port 8 nsew
<< end >>
