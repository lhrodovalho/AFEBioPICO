* lna-ota buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "./afe_no_pseudo.spice"


* supply voltages
vdda	vdda 0 1.8
vgnda	gnda 0 0.9
vssa	vssa 0 0.0

* input signals
vin	in gnda dc 0 ac 1 SINE(0 50m 1 0 0 0)
einp	ip gnda in gnda  0.5
einm	im gnda in gnda -0.5

* DUT
x0 ip im om op fsb ib vdda gnda vssa lna
IB   vdda ib 10n
CLP  op gnda 10p
CLM  om gnda 10p

.option gmin=1e-12
*.option NOOPITER
.option NOINIT
.option METHOD=Gear
.control
	noise v(op,om) vin dec 10 1 100
	print inoise_total onoise_total
	setplot noise1
	plot inoise_spectrum loglog
    
.endc

.end
