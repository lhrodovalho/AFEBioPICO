* lna-ota buffer testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "lna_ota.spice"
.include "vga_ota.spice"

.subckt buffer in out ib vdda vssa

xpa0 ib  ib  vdda vdda vssa p1_8 m=8
xpb0 n   ib  vdda vdda vssa p1_8 m=8
xnb0 n   n   vssa vssa      n1_8 m=8

xpc0 yn  ib  vdda vdda vssa p1_8 m=8
xnc2 out out xn   vssa 	    n1_8 m=8
xnc1 yn  in  xn   vssa 	    n1_8 m=8
xnc0 xn  yn  vssa vssa 	    n1_8 m=16

xpd0 xp  yp  vdda vdda vssa p1_8 m=16
xpd1 yp  in  xp   vdda vssa p1_8 m=8
xpd2 out out xp   vdda vssa p1_8 m=8
xnd0 yp  n   vssa vssa      n1_8 m=8

.ends

.subckt vga_buf in out ib vdda gnda vssa

	Xamp x in outx ib vdda vssa vga_ota
	Xbuf outx out  ib vdda vssa buffer
	ri gnda x   1Meg
	rf x    out 10Meg

.ends


vdd vdd 0 1.8
vss vss 0 0.0
ecm cm vss vdd vss 0.5

vin in cm dc 0 ac 1 SINE(0 0.4 0.5k 0 0 0)

* DUT
IB ib vss 10n
X0 out0 in out0 ib vdd vss lna_ota
X1 out1 in out1 ib vdd vss vga_ota
CL0 out0 cm 1p
CL1 out1 cm 1p

*.save v(in) v(out0) v(out1) v(ib) v(x0.x) v(x0.y) i(vdd)
.nodeset v(ib) 1.4
*.option gmin=1e-12
.option scale=1e-6
.control

	op
	print in out ib x0.x x0.y i(vdd)

	dc vin -10m 10m 100u
	let dc_vi = v(in)
	let dc_vo = v(out)
	wrdata lna_ota_dc_vo.txt dc_vo
	plot in out0 out1

    
.endc

.end
