magic
tech sky130A
timestamp 1638020595
<< locali >>
rect 0 18670 40 18680
rect 0 18650 10 18670
rect 30 18650 40 18670
rect 0 18510 40 18650
rect 0 18490 10 18510
rect 30 18490 40 18510
rect 0 18480 40 18490
rect 80 18670 120 18680
rect 80 18650 90 18670
rect 110 18650 120 18670
rect 80 18510 120 18650
rect 80 18490 90 18510
rect 110 18490 120 18510
rect 80 18480 120 18490
rect 160 18670 200 18680
rect 160 18650 170 18670
rect 190 18650 200 18670
rect 160 18510 200 18650
rect 160 18490 170 18510
rect 190 18490 200 18510
rect 160 18480 200 18490
rect 240 18670 280 18680
rect 240 18650 250 18670
rect 270 18650 280 18670
rect 240 18510 280 18650
rect 240 18490 250 18510
rect 270 18490 280 18510
rect 240 18480 280 18490
rect 320 18670 360 18680
rect 320 18650 330 18670
rect 350 18650 360 18670
rect 320 18510 360 18650
rect 320 18490 330 18510
rect 350 18490 360 18510
rect 320 18480 360 18490
rect 400 18670 440 18680
rect 400 18650 410 18670
rect 430 18650 440 18670
rect 400 18510 440 18650
rect 400 18490 410 18510
rect 430 18490 440 18510
rect 400 18480 440 18490
rect 480 18670 520 18680
rect 480 18650 490 18670
rect 510 18650 520 18670
rect 480 18510 520 18650
rect 480 18490 490 18510
rect 510 18490 520 18510
rect 480 18480 520 18490
rect 560 18670 600 18680
rect 560 18650 570 18670
rect 590 18650 600 18670
rect 560 18510 600 18650
rect 560 18490 570 18510
rect 590 18490 600 18510
rect 560 18480 600 18490
rect 640 18670 680 18680
rect 640 18650 650 18670
rect 670 18650 680 18670
rect 640 18510 680 18650
rect 640 18490 650 18510
rect 670 18490 680 18510
rect 640 18480 680 18490
rect 720 18670 760 18680
rect 720 18650 730 18670
rect 750 18650 760 18670
rect 720 18510 760 18650
rect 720 18490 730 18510
rect 750 18490 760 18510
rect 720 18480 760 18490
rect 800 18670 840 18680
rect 800 18650 810 18670
rect 830 18650 840 18670
rect 800 18510 840 18650
rect 800 18490 810 18510
rect 830 18490 840 18510
rect 800 18480 840 18490
rect 880 18670 920 18680
rect 880 18650 890 18670
rect 910 18650 920 18670
rect 880 18510 920 18650
rect 880 18490 890 18510
rect 910 18490 920 18510
rect 880 18480 920 18490
rect 960 18670 1000 18680
rect 960 18650 970 18670
rect 990 18650 1000 18670
rect 960 18510 1000 18650
rect 960 18490 970 18510
rect 990 18490 1000 18510
rect 960 18480 1000 18490
rect 1040 18670 1080 18680
rect 1040 18650 1050 18670
rect 1070 18650 1080 18670
rect 1040 18510 1080 18650
rect 1040 18490 1050 18510
rect 1070 18490 1080 18510
rect 1040 18480 1080 18490
rect 1120 18670 1160 18680
rect 1120 18650 1130 18670
rect 1150 18650 1160 18670
rect 1120 18510 1160 18650
rect 1120 18490 1130 18510
rect 1150 18490 1160 18510
rect 1120 18480 1160 18490
rect 1200 18670 1240 18680
rect 1200 18650 1210 18670
rect 1230 18650 1240 18670
rect 1200 18510 1240 18650
rect 1200 18490 1210 18510
rect 1230 18490 1240 18510
rect 1200 18480 1240 18490
rect 1280 18670 1320 18680
rect 1280 18650 1290 18670
rect 1310 18650 1320 18670
rect 1280 18510 1320 18650
rect 1280 18490 1290 18510
rect 1310 18490 1320 18510
rect 1280 18480 1320 18490
rect 1360 18670 1400 18680
rect 1360 18650 1370 18670
rect 1390 18650 1400 18670
rect 1360 18510 1400 18650
rect 1360 18490 1370 18510
rect 1390 18490 1400 18510
rect 1360 18480 1400 18490
rect 1440 18670 1480 18680
rect 1440 18650 1450 18670
rect 1470 18650 1480 18670
rect 1440 18510 1480 18650
rect 1440 18490 1450 18510
rect 1470 18490 1480 18510
rect 1440 18480 1480 18490
rect 1520 18670 1560 18680
rect 1520 18650 1530 18670
rect 1550 18650 1560 18670
rect 1520 18510 1560 18650
rect 1520 18490 1530 18510
rect 1550 18490 1560 18510
rect 1520 18480 1560 18490
rect 1600 18670 1640 18680
rect 1600 18650 1610 18670
rect 1630 18650 1640 18670
rect 1600 18510 1640 18650
rect 1600 18490 1610 18510
rect 1630 18490 1640 18510
rect 1600 18480 1640 18490
rect 1680 18670 1720 18680
rect 1680 18650 1690 18670
rect 1710 18650 1720 18670
rect 1680 18510 1720 18650
rect 1680 18490 1690 18510
rect 1710 18490 1720 18510
rect 1680 18480 1720 18490
rect 1760 18670 1800 18680
rect 1760 18650 1770 18670
rect 1790 18650 1800 18670
rect 1760 18510 1800 18650
rect 1760 18490 1770 18510
rect 1790 18490 1800 18510
rect 1760 18480 1800 18490
rect 1840 18670 1880 18680
rect 1840 18650 1850 18670
rect 1870 18650 1880 18670
rect 1840 18510 1880 18650
rect 1840 18490 1850 18510
rect 1870 18490 1880 18510
rect 1840 18480 1880 18490
rect 1920 18670 1960 18680
rect 1920 18650 1930 18670
rect 1950 18650 1960 18670
rect 1920 18510 1960 18650
rect 1920 18490 1930 18510
rect 1950 18490 1960 18510
rect 1920 18480 1960 18490
rect 2000 18670 2040 18680
rect 2000 18650 2010 18670
rect 2030 18650 2040 18670
rect 2000 18510 2040 18650
rect 2000 18490 2010 18510
rect 2030 18490 2040 18510
rect 2000 18480 2040 18490
rect 2080 18670 2120 18680
rect 2080 18650 2090 18670
rect 2110 18650 2120 18670
rect 2080 18510 2120 18650
rect 2080 18490 2090 18510
rect 2110 18490 2120 18510
rect 2080 18480 2120 18490
rect 2160 18670 2200 18680
rect 2160 18650 2170 18670
rect 2190 18650 2200 18670
rect 2160 18510 2200 18650
rect 2160 18490 2170 18510
rect 2190 18490 2200 18510
rect 2160 18480 2200 18490
rect 2240 18670 2280 18680
rect 2240 18650 2250 18670
rect 2270 18650 2280 18670
rect 2240 18510 2280 18650
rect 2240 18490 2250 18510
rect 2270 18490 2280 18510
rect 2240 18480 2280 18490
rect 2320 18670 2360 18680
rect 2320 18650 2330 18670
rect 2350 18650 2360 18670
rect 2320 18510 2360 18650
rect 2320 18490 2330 18510
rect 2350 18490 2360 18510
rect 2320 18480 2360 18490
rect 2400 18670 2440 18680
rect 2400 18650 2410 18670
rect 2430 18650 2440 18670
rect 2400 18510 2440 18650
rect 2400 18490 2410 18510
rect 2430 18490 2440 18510
rect 2400 18480 2440 18490
rect 2480 18670 2520 18680
rect 2480 18650 2490 18670
rect 2510 18650 2520 18670
rect 2480 18510 2520 18650
rect 2480 18490 2490 18510
rect 2510 18490 2520 18510
rect 2480 18480 2520 18490
rect 2560 18670 2600 18680
rect 2560 18650 2570 18670
rect 2590 18650 2600 18670
rect 2560 18510 2600 18650
rect 2560 18490 2570 18510
rect 2590 18490 2600 18510
rect 2560 18480 2600 18490
rect 2640 18670 2680 18680
rect 2640 18650 2650 18670
rect 2670 18650 2680 18670
rect 2640 18510 2680 18650
rect 2640 18490 2650 18510
rect 2670 18490 2680 18510
rect 2640 18480 2680 18490
rect 2720 18670 2760 18680
rect 2720 18650 2730 18670
rect 2750 18650 2760 18670
rect 2720 18510 2760 18650
rect 2720 18490 2730 18510
rect 2750 18490 2760 18510
rect 2720 18480 2760 18490
rect 2800 18670 2840 18680
rect 2800 18650 2810 18670
rect 2830 18650 2840 18670
rect 2800 18510 2840 18650
rect 2800 18490 2810 18510
rect 2830 18490 2840 18510
rect 2800 18480 2840 18490
rect 2880 18670 2920 18680
rect 2880 18650 2890 18670
rect 2910 18650 2920 18670
rect 2880 18510 2920 18650
rect 2880 18490 2890 18510
rect 2910 18490 2920 18510
rect 2880 18480 2920 18490
rect 2960 18670 3000 18680
rect 2960 18650 2970 18670
rect 2990 18650 3000 18670
rect 2960 18510 3000 18650
rect 2960 18490 2970 18510
rect 2990 18490 3000 18510
rect 2960 18480 3000 18490
rect 3040 18670 3080 18680
rect 3040 18650 3050 18670
rect 3070 18650 3080 18670
rect 3040 18510 3080 18650
rect 3040 18490 3050 18510
rect 3070 18490 3080 18510
rect 3040 18480 3080 18490
rect 3120 18670 3160 18680
rect 3120 18650 3130 18670
rect 3150 18650 3160 18670
rect 3120 18510 3160 18650
rect 3120 18490 3130 18510
rect 3150 18490 3160 18510
rect 3120 18480 3160 18490
rect 3200 18670 3240 18680
rect 3200 18650 3210 18670
rect 3230 18650 3240 18670
rect 3200 18510 3240 18650
rect 3200 18490 3210 18510
rect 3230 18490 3240 18510
rect 3200 18480 3240 18490
rect 3280 18670 3320 18680
rect 3280 18650 3290 18670
rect 3310 18650 3320 18670
rect 3280 18510 3320 18650
rect 3280 18490 3290 18510
rect 3310 18490 3320 18510
rect 3280 18480 3320 18490
rect 3360 18670 3400 18680
rect 3360 18650 3370 18670
rect 3390 18650 3400 18670
rect 3360 18510 3400 18650
rect 3360 18490 3370 18510
rect 3390 18490 3400 18510
rect 3360 18480 3400 18490
rect 3440 18670 3480 18680
rect 3440 18650 3450 18670
rect 3470 18650 3480 18670
rect 3440 18510 3480 18650
rect 3440 18490 3450 18510
rect 3470 18490 3480 18510
rect 3440 18480 3480 18490
rect 3520 18670 3560 18680
rect 3520 18650 3530 18670
rect 3550 18650 3560 18670
rect 3520 18510 3560 18650
rect 3520 18490 3530 18510
rect 3550 18490 3560 18510
rect 3520 18480 3560 18490
rect 3600 18670 3640 18680
rect 3600 18650 3610 18670
rect 3630 18650 3640 18670
rect 3600 18510 3640 18650
rect 3600 18490 3610 18510
rect 3630 18490 3640 18510
rect 3600 18480 3640 18490
rect 3680 18670 3720 18680
rect 3680 18650 3690 18670
rect 3710 18650 3720 18670
rect 3680 18510 3720 18650
rect 3680 18490 3690 18510
rect 3710 18490 3720 18510
rect 3680 18480 3720 18490
rect 3760 18670 3800 18680
rect 3760 18650 3770 18670
rect 3790 18650 3800 18670
rect 3760 18510 3800 18650
rect 3760 18490 3770 18510
rect 3790 18490 3800 18510
rect 3760 18480 3800 18490
rect 3840 18670 3880 18680
rect 3840 18650 3850 18670
rect 3870 18650 3880 18670
rect 3840 18510 3880 18650
rect 3840 18490 3850 18510
rect 3870 18490 3880 18510
rect 3840 18480 3880 18490
rect 3920 18670 3960 18680
rect 3920 18650 3930 18670
rect 3950 18650 3960 18670
rect 3920 18510 3960 18650
rect 3920 18490 3930 18510
rect 3950 18490 3960 18510
rect 3920 18480 3960 18490
rect 4000 18670 4040 18680
rect 4000 18650 4010 18670
rect 4030 18650 4040 18670
rect 4000 18510 4040 18650
rect 4000 18490 4010 18510
rect 4030 18490 4040 18510
rect 4000 18480 4040 18490
rect 4080 18670 4120 18680
rect 4080 18650 4090 18670
rect 4110 18650 4120 18670
rect 4080 18510 4120 18650
rect 4080 18490 4090 18510
rect 4110 18490 4120 18510
rect 4080 18480 4120 18490
rect 4160 18670 4200 18680
rect 4160 18650 4170 18670
rect 4190 18650 4200 18670
rect 4160 18510 4200 18650
rect 4160 18490 4170 18510
rect 4190 18490 4200 18510
rect 4160 18480 4200 18490
rect 4240 18480 4280 18680
rect 4320 18480 4360 18680
rect 4400 18480 4440 18680
rect 4480 18480 4520 18680
rect 4560 18480 4600 18680
rect 4640 18480 4680 18680
rect 4720 18480 4760 18680
rect 4800 18480 4840 18680
rect 4880 18480 4920 18680
rect 4960 18480 5000 18680
rect 5040 18480 5080 18680
rect 5120 18480 5160 18680
rect 5200 18480 5240 18680
rect 5280 18480 5320 18680
rect 5360 18480 5400 18680
rect 5440 18480 5480 18680
rect 5520 18480 5560 18680
rect 5600 18480 5640 18680
rect 5680 18480 5720 18680
rect 5760 18480 5800 18680
rect 5840 18480 5880 18680
rect 5920 18480 5960 18680
rect 6000 18480 6040 18680
rect 6080 18480 6120 18680
rect 6160 18480 6200 18680
rect 6240 18670 6280 18680
rect 6240 18650 6250 18670
rect 6270 18650 6280 18670
rect 6240 18510 6280 18650
rect 6240 18490 6250 18510
rect 6270 18490 6280 18510
rect 6240 18480 6280 18490
rect 6320 18670 6360 18680
rect 6320 18650 6330 18670
rect 6350 18650 6360 18670
rect 6320 18510 6360 18650
rect 6320 18490 6330 18510
rect 6350 18490 6360 18510
rect 6320 18480 6360 18490
rect 6400 18670 6440 18680
rect 6400 18650 6410 18670
rect 6430 18650 6440 18670
rect 6400 18510 6440 18650
rect 6400 18490 6410 18510
rect 6430 18490 6440 18510
rect 6400 18480 6440 18490
rect 6480 18670 6520 18680
rect 6480 18650 6490 18670
rect 6510 18650 6520 18670
rect 6480 18510 6520 18650
rect 6480 18490 6490 18510
rect 6510 18490 6520 18510
rect 6480 18480 6520 18490
rect 6560 18670 6600 18680
rect 6560 18650 6570 18670
rect 6590 18650 6600 18670
rect 6560 18510 6600 18650
rect 6560 18490 6570 18510
rect 6590 18490 6600 18510
rect 6560 18480 6600 18490
rect 6640 18670 6680 18680
rect 6640 18650 6650 18670
rect 6670 18650 6680 18670
rect 6640 18510 6680 18650
rect 6640 18490 6650 18510
rect 6670 18490 6680 18510
rect 6640 18480 6680 18490
rect 6720 18670 6760 18680
rect 6720 18650 6730 18670
rect 6750 18650 6760 18670
rect 6720 18510 6760 18650
rect 6720 18490 6730 18510
rect 6750 18490 6760 18510
rect 6720 18480 6760 18490
rect 6800 18670 6840 18680
rect 6800 18650 6810 18670
rect 6830 18650 6840 18670
rect 6800 18510 6840 18650
rect 6800 18490 6810 18510
rect 6830 18490 6840 18510
rect 6800 18480 6840 18490
rect 6880 18670 6920 18680
rect 6880 18650 6890 18670
rect 6910 18650 6920 18670
rect 6880 18510 6920 18650
rect 6880 18490 6890 18510
rect 6910 18490 6920 18510
rect 6880 18480 6920 18490
rect 6960 18670 7000 18680
rect 6960 18650 6970 18670
rect 6990 18650 7000 18670
rect 6960 18510 7000 18650
rect 6960 18490 6970 18510
rect 6990 18490 7000 18510
rect 6960 18480 7000 18490
rect 7040 18670 7080 18680
rect 7040 18650 7050 18670
rect 7070 18650 7080 18670
rect 7040 18510 7080 18650
rect 7040 18490 7050 18510
rect 7070 18490 7080 18510
rect 7040 18480 7080 18490
rect 7120 18670 7160 18680
rect 7120 18650 7130 18670
rect 7150 18650 7160 18670
rect 7120 18510 7160 18650
rect 7120 18490 7130 18510
rect 7150 18490 7160 18510
rect 7120 18480 7160 18490
rect 7200 18670 7240 18680
rect 7200 18650 7210 18670
rect 7230 18650 7240 18670
rect 7200 18510 7240 18650
rect 7200 18490 7210 18510
rect 7230 18490 7240 18510
rect 7200 18480 7240 18490
rect 7280 18670 7320 18680
rect 7280 18650 7290 18670
rect 7310 18650 7320 18670
rect 7280 18510 7320 18650
rect 7280 18490 7290 18510
rect 7310 18490 7320 18510
rect 7280 18480 7320 18490
rect 7360 18670 7400 18680
rect 7360 18650 7370 18670
rect 7390 18650 7400 18670
rect 7360 18510 7400 18650
rect 7360 18490 7370 18510
rect 7390 18490 7400 18510
rect 7360 18480 7400 18490
rect 7440 18670 7480 18680
rect 7440 18650 7450 18670
rect 7470 18650 7480 18670
rect 7440 18510 7480 18650
rect 7440 18490 7450 18510
rect 7470 18490 7480 18510
rect 7440 18480 7480 18490
rect 7520 18670 7560 18680
rect 7520 18650 7530 18670
rect 7550 18650 7560 18670
rect 7520 18510 7560 18650
rect 7520 18490 7530 18510
rect 7550 18490 7560 18510
rect 7520 18480 7560 18490
rect 7600 18670 7640 18680
rect 7600 18650 7610 18670
rect 7630 18650 7640 18670
rect 7600 18510 7640 18650
rect 7600 18490 7610 18510
rect 7630 18490 7640 18510
rect 7600 18480 7640 18490
rect 7680 18670 7720 18680
rect 7680 18650 7690 18670
rect 7710 18650 7720 18670
rect 7680 18510 7720 18650
rect 7680 18490 7690 18510
rect 7710 18490 7720 18510
rect 7680 18480 7720 18490
rect 7760 18670 7800 18680
rect 7760 18650 7770 18670
rect 7790 18650 7800 18670
rect 7760 18510 7800 18650
rect 7760 18490 7770 18510
rect 7790 18490 7800 18510
rect 7760 18480 7800 18490
rect 7840 18670 7880 18680
rect 7840 18650 7850 18670
rect 7870 18650 7880 18670
rect 7840 18510 7880 18650
rect 7840 18490 7850 18510
rect 7870 18490 7880 18510
rect 7840 18480 7880 18490
rect 7920 18670 7960 18680
rect 7920 18650 7930 18670
rect 7950 18650 7960 18670
rect 7920 18510 7960 18650
rect 7920 18490 7930 18510
rect 7950 18490 7960 18510
rect 7920 18480 7960 18490
rect 8000 18670 8040 18680
rect 8000 18650 8010 18670
rect 8030 18650 8040 18670
rect 8000 18510 8040 18650
rect 8000 18490 8010 18510
rect 8030 18490 8040 18510
rect 8000 18480 8040 18490
rect 8080 18670 8120 18680
rect 8080 18650 8090 18670
rect 8110 18650 8120 18670
rect 8080 18510 8120 18650
rect 8080 18490 8090 18510
rect 8110 18490 8120 18510
rect 8080 18480 8120 18490
rect 8160 18670 8200 18680
rect 8160 18650 8170 18670
rect 8190 18650 8200 18670
rect 8160 18510 8200 18650
rect 8160 18490 8170 18510
rect 8190 18490 8200 18510
rect 8160 18480 8200 18490
rect 8240 18670 8280 18680
rect 8240 18650 8250 18670
rect 8270 18650 8280 18670
rect 8240 18510 8280 18650
rect 8240 18490 8250 18510
rect 8270 18490 8280 18510
rect 8240 18480 8280 18490
rect 8320 18670 8360 18680
rect 8320 18650 8330 18670
rect 8350 18650 8360 18670
rect 8320 18510 8360 18650
rect 8320 18490 8330 18510
rect 8350 18490 8360 18510
rect 8320 18480 8360 18490
rect 8400 18670 8440 18680
rect 8400 18650 8410 18670
rect 8430 18650 8440 18670
rect 8400 18510 8440 18650
rect 8400 18490 8410 18510
rect 8430 18490 8440 18510
rect 8400 18480 8440 18490
rect 8480 18670 8520 18680
rect 8480 18650 8490 18670
rect 8510 18650 8520 18670
rect 8480 18510 8520 18650
rect 8480 18490 8490 18510
rect 8510 18490 8520 18510
rect 8480 18480 8520 18490
rect 8560 18670 8600 18680
rect 8560 18650 8570 18670
rect 8590 18650 8600 18670
rect 8560 18510 8600 18650
rect 8560 18490 8570 18510
rect 8590 18490 8600 18510
rect 8560 18480 8600 18490
rect 8640 18670 8680 18680
rect 8640 18650 8650 18670
rect 8670 18650 8680 18670
rect 8640 18510 8680 18650
rect 8640 18490 8650 18510
rect 8670 18490 8680 18510
rect 8640 18480 8680 18490
rect 8720 18670 8760 18680
rect 8720 18650 8730 18670
rect 8750 18650 8760 18670
rect 8720 18510 8760 18650
rect 8720 18490 8730 18510
rect 8750 18490 8760 18510
rect 8720 18480 8760 18490
rect 8800 18670 8840 18680
rect 8800 18650 8810 18670
rect 8830 18650 8840 18670
rect 8800 18510 8840 18650
rect 8800 18490 8810 18510
rect 8830 18490 8840 18510
rect 8800 18480 8840 18490
rect 8880 18670 8920 18680
rect 8880 18650 8890 18670
rect 8910 18650 8920 18670
rect 8880 18510 8920 18650
rect 8880 18490 8890 18510
rect 8910 18490 8920 18510
rect 8880 18480 8920 18490
rect 8960 18670 9000 18680
rect 8960 18650 8970 18670
rect 8990 18650 9000 18670
rect 8960 18510 9000 18650
rect 8960 18490 8970 18510
rect 8990 18490 9000 18510
rect 8960 18480 9000 18490
rect 9040 18670 9080 18680
rect 9040 18650 9050 18670
rect 9070 18650 9080 18670
rect 9040 18510 9080 18650
rect 9040 18490 9050 18510
rect 9070 18490 9080 18510
rect 9040 18480 9080 18490
rect 9120 18670 9160 18680
rect 9120 18650 9130 18670
rect 9150 18650 9160 18670
rect 9120 18510 9160 18650
rect 9120 18490 9130 18510
rect 9150 18490 9160 18510
rect 9120 18480 9160 18490
rect 9200 18670 9240 18680
rect 9200 18650 9210 18670
rect 9230 18650 9240 18670
rect 9200 18510 9240 18650
rect 9200 18490 9210 18510
rect 9230 18490 9240 18510
rect 9200 18480 9240 18490
rect 9280 18670 9320 18680
rect 9280 18650 9290 18670
rect 9310 18650 9320 18670
rect 9280 18510 9320 18650
rect 9280 18490 9290 18510
rect 9310 18490 9320 18510
rect 9280 18480 9320 18490
rect 9360 18670 9400 18680
rect 9360 18650 9370 18670
rect 9390 18650 9400 18670
rect 9360 18510 9400 18650
rect 9360 18490 9370 18510
rect 9390 18490 9400 18510
rect 9360 18480 9400 18490
rect 9440 18670 9480 18680
rect 9440 18650 9450 18670
rect 9470 18650 9480 18670
rect 9440 18510 9480 18650
rect 9440 18490 9450 18510
rect 9470 18490 9480 18510
rect 9440 18480 9480 18490
rect 9520 18480 9560 18680
rect 9600 18480 9640 18680
rect 9680 18480 9720 18680
rect 9760 18480 9800 18680
rect 9840 18480 9880 18680
rect 9920 18480 9960 18680
rect 10000 18480 10040 18680
rect 10080 18480 10120 18680
rect 10160 18480 10200 18680
rect 10240 18480 10280 18680
rect 10320 18480 10360 18680
rect 10400 18480 10440 18680
rect 10480 18480 10520 18680
rect 10560 18480 10600 18680
rect 10640 18480 10680 18680
rect 10720 18480 10760 18680
rect 10800 18480 10840 18680
rect 10880 18480 10920 18680
rect 10960 18480 11000 18680
rect 11040 18480 11080 18680
rect 11120 18480 11160 18680
rect 11200 18480 11240 18680
rect 11280 18480 11320 18680
rect 11360 18480 11400 18680
rect 11440 18480 11480 18680
rect 11560 18670 11600 18680
rect 11560 18650 11570 18670
rect 11590 18650 11600 18670
rect 11560 18510 11600 18650
rect 11560 18490 11570 18510
rect 11590 18490 11600 18510
rect 11560 18480 11600 18490
rect 11640 18670 11680 18680
rect 11640 18650 11650 18670
rect 11670 18650 11680 18670
rect 11640 18510 11680 18650
rect 11640 18490 11650 18510
rect 11670 18490 11680 18510
rect 11640 18480 11680 18490
rect 11720 18670 11760 18680
rect 11720 18650 11730 18670
rect 11750 18650 11760 18670
rect 11720 18510 11760 18650
rect 11720 18490 11730 18510
rect 11750 18490 11760 18510
rect 11720 18480 11760 18490
rect 11800 18670 11840 18680
rect 11800 18650 11810 18670
rect 11830 18650 11840 18670
rect 11800 18510 11840 18650
rect 11800 18490 11810 18510
rect 11830 18490 11840 18510
rect 11800 18480 11840 18490
rect 11880 18670 11920 18680
rect 11880 18650 11890 18670
rect 11910 18650 11920 18670
rect 11880 18510 11920 18650
rect 11880 18490 11890 18510
rect 11910 18490 11920 18510
rect 11880 18480 11920 18490
rect 11960 18670 12000 18680
rect 11960 18650 11970 18670
rect 11990 18650 12000 18670
rect 11960 18510 12000 18650
rect 11960 18490 11970 18510
rect 11990 18490 12000 18510
rect 11960 18480 12000 18490
rect 12040 18670 12080 18680
rect 12040 18650 12050 18670
rect 12070 18650 12080 18670
rect 12040 18510 12080 18650
rect 12040 18490 12050 18510
rect 12070 18490 12080 18510
rect 12040 18480 12080 18490
rect 12120 18670 12160 18680
rect 12120 18650 12130 18670
rect 12150 18650 12160 18670
rect 12120 18510 12160 18650
rect 12120 18490 12130 18510
rect 12150 18490 12160 18510
rect 12120 18480 12160 18490
rect 12200 18670 12240 18680
rect 12200 18650 12210 18670
rect 12230 18650 12240 18670
rect 12200 18510 12240 18650
rect 12200 18490 12210 18510
rect 12230 18490 12240 18510
rect 12200 18480 12240 18490
rect 12280 18670 12320 18680
rect 12280 18650 12290 18670
rect 12310 18650 12320 18670
rect 12280 18510 12320 18650
rect 12280 18490 12290 18510
rect 12310 18490 12320 18510
rect 12280 18480 12320 18490
rect 12360 18670 12400 18680
rect 12360 18650 12370 18670
rect 12390 18650 12400 18670
rect 12360 18510 12400 18650
rect 12360 18490 12370 18510
rect 12390 18490 12400 18510
rect 12360 18480 12400 18490
rect 12440 18670 12480 18680
rect 12440 18650 12450 18670
rect 12470 18650 12480 18670
rect 12440 18510 12480 18650
rect 12440 18490 12450 18510
rect 12470 18490 12480 18510
rect 12440 18480 12480 18490
rect 12520 18670 12560 18680
rect 12520 18650 12530 18670
rect 12550 18650 12560 18670
rect 12520 18510 12560 18650
rect 12520 18490 12530 18510
rect 12550 18490 12560 18510
rect 12520 18480 12560 18490
rect 12600 18670 12640 18680
rect 12600 18650 12610 18670
rect 12630 18650 12640 18670
rect 12600 18510 12640 18650
rect 12600 18490 12610 18510
rect 12630 18490 12640 18510
rect 12600 18480 12640 18490
rect 12680 18670 12720 18680
rect 12680 18650 12690 18670
rect 12710 18650 12720 18670
rect 12680 18510 12720 18650
rect 12680 18490 12690 18510
rect 12710 18490 12720 18510
rect 12680 18480 12720 18490
rect 12760 18670 12800 18680
rect 12760 18650 12770 18670
rect 12790 18650 12800 18670
rect 12760 18510 12800 18650
rect 12760 18490 12770 18510
rect 12790 18490 12800 18510
rect 12760 18480 12800 18490
rect 12840 18670 12880 18680
rect 12840 18650 12850 18670
rect 12870 18650 12880 18670
rect 12840 18510 12880 18650
rect 12840 18490 12850 18510
rect 12870 18490 12880 18510
rect 12840 18480 12880 18490
rect 12920 18670 12960 18680
rect 12920 18650 12930 18670
rect 12950 18650 12960 18670
rect 12920 18510 12960 18650
rect 12920 18490 12930 18510
rect 12950 18490 12960 18510
rect 12920 18480 12960 18490
rect 13000 18670 13040 18680
rect 13000 18650 13010 18670
rect 13030 18650 13040 18670
rect 13000 18510 13040 18650
rect 13000 18490 13010 18510
rect 13030 18490 13040 18510
rect 13000 18480 13040 18490
rect 13080 18670 13120 18680
rect 13080 18650 13090 18670
rect 13110 18650 13120 18670
rect 13080 18510 13120 18650
rect 13080 18490 13090 18510
rect 13110 18490 13120 18510
rect 13080 18480 13120 18490
rect 13160 18670 13200 18680
rect 13160 18650 13170 18670
rect 13190 18650 13200 18670
rect 13160 18510 13200 18650
rect 13160 18490 13170 18510
rect 13190 18490 13200 18510
rect 13160 18480 13200 18490
rect 13240 18670 13280 18680
rect 13240 18650 13250 18670
rect 13270 18650 13280 18670
rect 13240 18510 13280 18650
rect 13240 18490 13250 18510
rect 13270 18490 13280 18510
rect 13240 18480 13280 18490
rect 13320 18670 13360 18680
rect 13320 18650 13330 18670
rect 13350 18650 13360 18670
rect 13320 18510 13360 18650
rect 13320 18490 13330 18510
rect 13350 18490 13360 18510
rect 13320 18480 13360 18490
rect 13400 18670 13440 18680
rect 13400 18650 13410 18670
rect 13430 18650 13440 18670
rect 13400 18510 13440 18650
rect 13400 18490 13410 18510
rect 13430 18490 13440 18510
rect 13400 18480 13440 18490
rect 13480 18670 13520 18680
rect 13480 18650 13490 18670
rect 13510 18650 13520 18670
rect 13480 18510 13520 18650
rect 13480 18490 13490 18510
rect 13510 18490 13520 18510
rect 13480 18480 13520 18490
rect 13560 18670 13600 18680
rect 13560 18650 13570 18670
rect 13590 18650 13600 18670
rect 13560 18510 13600 18650
rect 13560 18490 13570 18510
rect 13590 18490 13600 18510
rect 13560 18480 13600 18490
rect 13640 18670 13680 18680
rect 13640 18650 13650 18670
rect 13670 18650 13680 18670
rect 13640 18510 13680 18650
rect 13640 18490 13650 18510
rect 13670 18490 13680 18510
rect 13640 18480 13680 18490
rect 13720 18670 13760 18680
rect 13720 18650 13730 18670
rect 13750 18650 13760 18670
rect 13720 18510 13760 18650
rect 13720 18490 13730 18510
rect 13750 18490 13760 18510
rect 13720 18480 13760 18490
rect 13800 18670 13840 18680
rect 13800 18650 13810 18670
rect 13830 18650 13840 18670
rect 13800 18510 13840 18650
rect 13800 18490 13810 18510
rect 13830 18490 13840 18510
rect 13800 18480 13840 18490
rect 13880 18670 13920 18680
rect 13880 18650 13890 18670
rect 13910 18650 13920 18670
rect 13880 18510 13920 18650
rect 13880 18490 13890 18510
rect 13910 18490 13920 18510
rect 13880 18480 13920 18490
rect 13960 18670 14000 18680
rect 13960 18650 13970 18670
rect 13990 18650 14000 18670
rect 13960 18510 14000 18650
rect 13960 18490 13970 18510
rect 13990 18490 14000 18510
rect 13960 18480 14000 18490
rect 14040 18670 14080 18680
rect 14040 18650 14050 18670
rect 14070 18650 14080 18670
rect 14040 18510 14080 18650
rect 14040 18490 14050 18510
rect 14070 18490 14080 18510
rect 14040 18480 14080 18490
rect 14120 18670 14160 18680
rect 14120 18650 14130 18670
rect 14150 18650 14160 18670
rect 14120 18510 14160 18650
rect 14120 18490 14130 18510
rect 14150 18490 14160 18510
rect 14120 18480 14160 18490
rect 14200 18670 14240 18680
rect 14200 18650 14210 18670
rect 14230 18650 14240 18670
rect 14200 18510 14240 18650
rect 14200 18490 14210 18510
rect 14230 18490 14240 18510
rect 14200 18480 14240 18490
rect 14280 18670 14320 18680
rect 14280 18650 14290 18670
rect 14310 18650 14320 18670
rect 14280 18510 14320 18650
rect 14280 18490 14290 18510
rect 14310 18490 14320 18510
rect 14280 18480 14320 18490
rect 14360 18670 14400 18680
rect 14360 18650 14370 18670
rect 14390 18650 14400 18670
rect 14360 18510 14400 18650
rect 14360 18490 14370 18510
rect 14390 18490 14400 18510
rect 14360 18480 14400 18490
rect 14440 18670 14480 18680
rect 14440 18650 14450 18670
rect 14470 18650 14480 18670
rect 14440 18510 14480 18650
rect 14440 18490 14450 18510
rect 14470 18490 14480 18510
rect 14440 18480 14480 18490
rect 14520 18670 14560 18680
rect 14520 18650 14530 18670
rect 14550 18650 14560 18670
rect 14520 18510 14560 18650
rect 14520 18490 14530 18510
rect 14550 18490 14560 18510
rect 14520 18480 14560 18490
rect 14600 18670 14640 18680
rect 14600 18650 14610 18670
rect 14630 18650 14640 18670
rect 14600 18510 14640 18650
rect 14600 18490 14610 18510
rect 14630 18490 14640 18510
rect 14600 18480 14640 18490
rect 14680 18670 14720 18680
rect 14680 18650 14690 18670
rect 14710 18650 14720 18670
rect 14680 18510 14720 18650
rect 14680 18490 14690 18510
rect 14710 18490 14720 18510
rect 14680 18480 14720 18490
rect 14760 18480 14800 18680
rect 14840 18480 14880 18680
rect 14920 18480 14960 18680
rect 15000 18480 15040 18680
rect 15080 18480 15120 18680
rect 15160 18480 15200 18680
rect 15240 18480 15280 18680
rect 15320 18480 15360 18680
rect 15400 18480 15440 18680
rect 15480 18480 15520 18680
rect 15560 18480 15600 18680
rect 15640 18480 15680 18680
rect 15720 18480 15760 18680
rect 15800 18480 15840 18680
rect 15880 18480 15920 18680
rect 15960 18480 16000 18680
rect 16040 18480 16080 18680
rect 16120 18480 16160 18680
rect 16200 18480 16240 18680
rect 16280 18480 16320 18680
rect 16360 18480 16400 18680
rect 16440 18480 16480 18680
rect 16520 18480 16560 18680
rect 16600 18480 16640 18680
rect 16680 18480 16720 18680
rect 16760 18670 16800 18680
rect 16760 18650 16770 18670
rect 16790 18650 16800 18670
rect 16760 18510 16800 18650
rect 16760 18490 16770 18510
rect 16790 18490 16800 18510
rect 16760 18480 16800 18490
rect 16840 18670 16880 18680
rect 16840 18650 16850 18670
rect 16870 18650 16880 18670
rect 16840 18510 16880 18650
rect 16840 18490 16850 18510
rect 16870 18490 16880 18510
rect 16840 18480 16880 18490
rect 16920 18670 16960 18680
rect 16920 18650 16930 18670
rect 16950 18650 16960 18670
rect 16920 18510 16960 18650
rect 16920 18490 16930 18510
rect 16950 18490 16960 18510
rect 16920 18480 16960 18490
rect 17000 18670 17040 18680
rect 17000 18650 17010 18670
rect 17030 18650 17040 18670
rect 17000 18510 17040 18650
rect 17000 18490 17010 18510
rect 17030 18490 17040 18510
rect 17000 18480 17040 18490
rect 17080 18670 17120 18680
rect 17080 18650 17090 18670
rect 17110 18650 17120 18670
rect 17080 18510 17120 18650
rect 17080 18490 17090 18510
rect 17110 18490 17120 18510
rect 17080 18480 17120 18490
rect 17160 18670 17200 18680
rect 17160 18650 17170 18670
rect 17190 18650 17200 18670
rect 17160 18510 17200 18650
rect 17160 18490 17170 18510
rect 17190 18490 17200 18510
rect 17160 18480 17200 18490
rect 17240 18670 17280 18680
rect 17240 18650 17250 18670
rect 17270 18650 17280 18670
rect 17240 18510 17280 18650
rect 17240 18490 17250 18510
rect 17270 18490 17280 18510
rect 17240 18480 17280 18490
rect 17320 18670 17360 18680
rect 17320 18650 17330 18670
rect 17350 18650 17360 18670
rect 17320 18510 17360 18650
rect 17320 18490 17330 18510
rect 17350 18490 17360 18510
rect 17320 18480 17360 18490
rect 17400 18670 17440 18680
rect 17400 18650 17410 18670
rect 17430 18650 17440 18670
rect 17400 18510 17440 18650
rect 17400 18490 17410 18510
rect 17430 18490 17440 18510
rect 17400 18480 17440 18490
rect 17480 18670 17520 18680
rect 17480 18650 17490 18670
rect 17510 18650 17520 18670
rect 17480 18510 17520 18650
rect 17480 18490 17490 18510
rect 17510 18490 17520 18510
rect 17480 18480 17520 18490
rect 17560 18670 17600 18680
rect 17560 18650 17570 18670
rect 17590 18650 17600 18670
rect 17560 18510 17600 18650
rect 17560 18490 17570 18510
rect 17590 18490 17600 18510
rect 17560 18480 17600 18490
rect 17640 18670 17680 18680
rect 17640 18650 17650 18670
rect 17670 18650 17680 18670
rect 17640 18510 17680 18650
rect 17640 18490 17650 18510
rect 17670 18490 17680 18510
rect 17640 18480 17680 18490
rect 17720 18670 17760 18680
rect 17720 18650 17730 18670
rect 17750 18650 17760 18670
rect 17720 18510 17760 18650
rect 17720 18490 17730 18510
rect 17750 18490 17760 18510
rect 17720 18480 17760 18490
rect 17800 18670 17840 18680
rect 17800 18650 17810 18670
rect 17830 18650 17840 18670
rect 17800 18510 17840 18650
rect 17800 18490 17810 18510
rect 17830 18490 17840 18510
rect 17800 18480 17840 18490
rect 17880 18670 17920 18680
rect 17880 18650 17890 18670
rect 17910 18650 17920 18670
rect 17880 18510 17920 18650
rect 17880 18490 17890 18510
rect 17910 18490 17920 18510
rect 17880 18480 17920 18490
rect 17960 18670 18000 18680
rect 17960 18650 17970 18670
rect 17990 18650 18000 18670
rect 17960 18510 18000 18650
rect 17960 18490 17970 18510
rect 17990 18490 18000 18510
rect 17960 18480 18000 18490
rect 18040 18670 18080 18680
rect 18040 18650 18050 18670
rect 18070 18650 18080 18670
rect 18040 18510 18080 18650
rect 18040 18490 18050 18510
rect 18070 18490 18080 18510
rect 18040 18480 18080 18490
rect 18120 18670 18160 18680
rect 18120 18650 18130 18670
rect 18150 18650 18160 18670
rect 18120 18510 18160 18650
rect 18120 18490 18130 18510
rect 18150 18490 18160 18510
rect 18120 18480 18160 18490
rect 18200 18670 18240 18680
rect 18200 18650 18210 18670
rect 18230 18650 18240 18670
rect 18200 18510 18240 18650
rect 18200 18490 18210 18510
rect 18230 18490 18240 18510
rect 18200 18480 18240 18490
rect 18280 18670 18320 18680
rect 18280 18650 18290 18670
rect 18310 18650 18320 18670
rect 18280 18510 18320 18650
rect 18280 18490 18290 18510
rect 18310 18490 18320 18510
rect 18280 18480 18320 18490
rect 18360 18670 18400 18680
rect 18360 18650 18370 18670
rect 18390 18650 18400 18670
rect 18360 18510 18400 18650
rect 18360 18490 18370 18510
rect 18390 18490 18400 18510
rect 18360 18480 18400 18490
rect 18440 18670 18480 18680
rect 18440 18650 18450 18670
rect 18470 18650 18480 18670
rect 18440 18510 18480 18650
rect 18440 18490 18450 18510
rect 18470 18490 18480 18510
rect 18440 18480 18480 18490
rect 18520 18670 18560 18680
rect 18520 18650 18530 18670
rect 18550 18650 18560 18670
rect 18520 18510 18560 18650
rect 18520 18490 18530 18510
rect 18550 18490 18560 18510
rect 18520 18480 18560 18490
rect 18600 18670 18640 18680
rect 18600 18650 18610 18670
rect 18630 18650 18640 18670
rect 18600 18510 18640 18650
rect 18600 18490 18610 18510
rect 18630 18490 18640 18510
rect 18600 18480 18640 18490
rect 18680 18670 18720 18680
rect 18680 18650 18690 18670
rect 18710 18650 18720 18670
rect 18680 18510 18720 18650
rect 18680 18490 18690 18510
rect 18710 18490 18720 18510
rect 18680 18480 18720 18490
rect 18760 18670 18800 18680
rect 18760 18650 18770 18670
rect 18790 18650 18800 18670
rect 18760 18510 18800 18650
rect 18760 18490 18770 18510
rect 18790 18490 18800 18510
rect 18760 18480 18800 18490
rect 18840 18670 18880 18680
rect 18840 18650 18850 18670
rect 18870 18650 18880 18670
rect 18840 18510 18880 18650
rect 18840 18490 18850 18510
rect 18870 18490 18880 18510
rect 18840 18480 18880 18490
rect 18920 18670 18960 18680
rect 18920 18650 18930 18670
rect 18950 18650 18960 18670
rect 18920 18510 18960 18650
rect 18920 18490 18930 18510
rect 18950 18490 18960 18510
rect 18920 18480 18960 18490
rect 19000 18670 19040 18680
rect 19000 18650 19010 18670
rect 19030 18650 19040 18670
rect 19000 18510 19040 18650
rect 19000 18490 19010 18510
rect 19030 18490 19040 18510
rect 19000 18480 19040 18490
rect 19080 18670 19120 18680
rect 19080 18650 19090 18670
rect 19110 18650 19120 18670
rect 19080 18510 19120 18650
rect 19080 18490 19090 18510
rect 19110 18490 19120 18510
rect 19080 18480 19120 18490
rect 19160 18670 19200 18680
rect 19160 18650 19170 18670
rect 19190 18650 19200 18670
rect 19160 18510 19200 18650
rect 19160 18490 19170 18510
rect 19190 18490 19200 18510
rect 19160 18480 19200 18490
rect 19240 18670 19280 18680
rect 19240 18650 19250 18670
rect 19270 18650 19280 18670
rect 19240 18510 19280 18650
rect 19240 18490 19250 18510
rect 19270 18490 19280 18510
rect 19240 18480 19280 18490
rect 19320 18670 19360 18680
rect 19320 18650 19330 18670
rect 19350 18650 19360 18670
rect 19320 18510 19360 18650
rect 19320 18490 19330 18510
rect 19350 18490 19360 18510
rect 19320 18480 19360 18490
rect 19400 18670 19440 18680
rect 19400 18650 19410 18670
rect 19430 18650 19440 18670
rect 19400 18510 19440 18650
rect 19400 18490 19410 18510
rect 19430 18490 19440 18510
rect 19400 18480 19440 18490
rect 19480 18670 19520 18680
rect 19480 18650 19490 18670
rect 19510 18650 19520 18670
rect 19480 18510 19520 18650
rect 19480 18490 19490 18510
rect 19510 18490 19520 18510
rect 19480 18480 19520 18490
rect 19560 18670 19600 18680
rect 19560 18650 19570 18670
rect 19590 18650 19600 18670
rect 19560 18510 19600 18650
rect 19560 18490 19570 18510
rect 19590 18490 19600 18510
rect 19560 18480 19600 18490
rect 19640 18670 19680 18680
rect 19640 18650 19650 18670
rect 19670 18650 19680 18670
rect 19640 18510 19680 18650
rect 19640 18490 19650 18510
rect 19670 18490 19680 18510
rect 19640 18480 19680 18490
rect 19720 18670 19760 18680
rect 19720 18650 19730 18670
rect 19750 18650 19760 18670
rect 19720 18510 19760 18650
rect 19720 18490 19730 18510
rect 19750 18490 19760 18510
rect 19720 18480 19760 18490
rect 19800 18670 19840 18680
rect 19800 18650 19810 18670
rect 19830 18650 19840 18670
rect 19800 18510 19840 18650
rect 19800 18490 19810 18510
rect 19830 18490 19840 18510
rect 19800 18480 19840 18490
rect 19880 18670 19920 18680
rect 19880 18650 19890 18670
rect 19910 18650 19920 18670
rect 19880 18510 19920 18650
rect 19880 18490 19890 18510
rect 19910 18490 19920 18510
rect 19880 18480 19920 18490
rect 19960 18670 20000 18680
rect 19960 18650 19970 18670
rect 19990 18650 20000 18670
rect 19960 18510 20000 18650
rect 19960 18490 19970 18510
rect 19990 18490 20000 18510
rect 19960 18480 20000 18490
rect 20040 18670 20080 18680
rect 20040 18650 20050 18670
rect 20070 18650 20080 18670
rect 20040 18510 20080 18650
rect 20040 18490 20050 18510
rect 20070 18490 20080 18510
rect 20040 18480 20080 18490
rect 20120 18670 20160 18680
rect 20120 18650 20130 18670
rect 20150 18650 20160 18670
rect 20120 18510 20160 18650
rect 20120 18490 20130 18510
rect 20150 18490 20160 18510
rect 20120 18480 20160 18490
rect 20200 18670 20240 18680
rect 20200 18650 20210 18670
rect 20230 18650 20240 18670
rect 20200 18510 20240 18650
rect 20200 18490 20210 18510
rect 20230 18490 20240 18510
rect 20200 18480 20240 18490
rect 20280 18670 20320 18680
rect 20280 18650 20290 18670
rect 20310 18650 20320 18670
rect 20280 18510 20320 18650
rect 20280 18490 20290 18510
rect 20310 18490 20320 18510
rect 20280 18480 20320 18490
rect 20360 18670 20400 18680
rect 20360 18650 20370 18670
rect 20390 18650 20400 18670
rect 20360 18510 20400 18650
rect 20360 18490 20370 18510
rect 20390 18490 20400 18510
rect 20360 18480 20400 18490
rect 20440 18670 20480 18680
rect 20440 18650 20450 18670
rect 20470 18650 20480 18670
rect 20440 18510 20480 18650
rect 20440 18490 20450 18510
rect 20470 18490 20480 18510
rect 20440 18480 20480 18490
rect 20520 18670 20560 18680
rect 20520 18650 20530 18670
rect 20550 18650 20560 18670
rect 20520 18510 20560 18650
rect 20520 18490 20530 18510
rect 20550 18490 20560 18510
rect 20520 18480 20560 18490
rect 20600 18670 20640 18680
rect 20600 18650 20610 18670
rect 20630 18650 20640 18670
rect 20600 18510 20640 18650
rect 20600 18490 20610 18510
rect 20630 18490 20640 18510
rect 20600 18480 20640 18490
rect 20680 18670 20720 18680
rect 20680 18650 20690 18670
rect 20710 18650 20720 18670
rect 20680 18510 20720 18650
rect 20680 18490 20690 18510
rect 20710 18490 20720 18510
rect 20680 18480 20720 18490
rect 20760 18670 20800 18680
rect 20760 18650 20770 18670
rect 20790 18650 20800 18670
rect 20760 18510 20800 18650
rect 20760 18490 20770 18510
rect 20790 18490 20800 18510
rect 20760 18480 20800 18490
rect 20840 18670 20880 18680
rect 20840 18650 20850 18670
rect 20870 18650 20880 18670
rect 20840 18510 20880 18650
rect 20840 18490 20850 18510
rect 20870 18490 20880 18510
rect 20840 18480 20880 18490
rect 20920 18670 20960 18680
rect 20920 18650 20930 18670
rect 20950 18650 20960 18670
rect 20920 18510 20960 18650
rect 20920 18490 20930 18510
rect 20950 18490 20960 18510
rect 20920 18480 20960 18490
rect 0 18430 40 18440
rect 0 18410 10 18430
rect 30 18410 40 18430
rect 0 18270 40 18410
rect 0 18250 10 18270
rect 30 18250 40 18270
rect 0 18240 40 18250
rect 80 18430 120 18440
rect 80 18410 90 18430
rect 110 18410 120 18430
rect 80 18270 120 18410
rect 80 18250 90 18270
rect 110 18250 120 18270
rect 80 18240 120 18250
rect 160 18430 200 18440
rect 160 18410 170 18430
rect 190 18410 200 18430
rect 160 18270 200 18410
rect 160 18250 170 18270
rect 190 18250 200 18270
rect 160 18240 200 18250
rect 240 18430 280 18440
rect 240 18410 250 18430
rect 270 18410 280 18430
rect 240 18270 280 18410
rect 240 18250 250 18270
rect 270 18250 280 18270
rect 240 18240 280 18250
rect 320 18430 360 18440
rect 320 18410 330 18430
rect 350 18410 360 18430
rect 320 18270 360 18410
rect 320 18250 330 18270
rect 350 18250 360 18270
rect 320 18240 360 18250
rect 400 18430 440 18440
rect 400 18410 410 18430
rect 430 18410 440 18430
rect 400 18270 440 18410
rect 400 18250 410 18270
rect 430 18250 440 18270
rect 400 18240 440 18250
rect 480 18430 520 18440
rect 480 18410 490 18430
rect 510 18410 520 18430
rect 480 18270 520 18410
rect 480 18250 490 18270
rect 510 18250 520 18270
rect 480 18240 520 18250
rect 560 18430 600 18440
rect 560 18410 570 18430
rect 590 18410 600 18430
rect 560 18270 600 18410
rect 560 18250 570 18270
rect 590 18250 600 18270
rect 560 18240 600 18250
rect 640 18430 680 18440
rect 640 18410 650 18430
rect 670 18410 680 18430
rect 640 18270 680 18410
rect 640 18250 650 18270
rect 670 18250 680 18270
rect 640 18240 680 18250
rect 720 18430 760 18440
rect 720 18410 730 18430
rect 750 18410 760 18430
rect 720 18270 760 18410
rect 720 18250 730 18270
rect 750 18250 760 18270
rect 720 18240 760 18250
rect 800 18430 840 18440
rect 800 18410 810 18430
rect 830 18410 840 18430
rect 800 18270 840 18410
rect 800 18250 810 18270
rect 830 18250 840 18270
rect 800 18240 840 18250
rect 880 18430 920 18440
rect 880 18410 890 18430
rect 910 18410 920 18430
rect 880 18270 920 18410
rect 880 18250 890 18270
rect 910 18250 920 18270
rect 880 18240 920 18250
rect 960 18430 1000 18440
rect 960 18410 970 18430
rect 990 18410 1000 18430
rect 960 18270 1000 18410
rect 960 18250 970 18270
rect 990 18250 1000 18270
rect 960 18240 1000 18250
rect 1040 18430 1080 18440
rect 1040 18410 1050 18430
rect 1070 18410 1080 18430
rect 1040 18270 1080 18410
rect 1040 18250 1050 18270
rect 1070 18250 1080 18270
rect 1040 18240 1080 18250
rect 1120 18430 1160 18440
rect 1120 18410 1130 18430
rect 1150 18410 1160 18430
rect 1120 18270 1160 18410
rect 1120 18250 1130 18270
rect 1150 18250 1160 18270
rect 1120 18240 1160 18250
rect 1200 18430 1240 18440
rect 1200 18410 1210 18430
rect 1230 18410 1240 18430
rect 1200 18270 1240 18410
rect 1200 18250 1210 18270
rect 1230 18250 1240 18270
rect 1200 18240 1240 18250
rect 1280 18430 1320 18440
rect 1280 18410 1290 18430
rect 1310 18410 1320 18430
rect 1280 18270 1320 18410
rect 1280 18250 1290 18270
rect 1310 18250 1320 18270
rect 1280 18240 1320 18250
rect 1360 18430 1400 18440
rect 1360 18410 1370 18430
rect 1390 18410 1400 18430
rect 1360 18270 1400 18410
rect 1360 18250 1370 18270
rect 1390 18250 1400 18270
rect 1360 18240 1400 18250
rect 1440 18430 1480 18440
rect 1440 18410 1450 18430
rect 1470 18410 1480 18430
rect 1440 18270 1480 18410
rect 1440 18250 1450 18270
rect 1470 18250 1480 18270
rect 1440 18240 1480 18250
rect 1520 18430 1560 18440
rect 1520 18410 1530 18430
rect 1550 18410 1560 18430
rect 1520 18270 1560 18410
rect 1520 18250 1530 18270
rect 1550 18250 1560 18270
rect 1520 18240 1560 18250
rect 1600 18430 1640 18440
rect 1600 18410 1610 18430
rect 1630 18410 1640 18430
rect 1600 18270 1640 18410
rect 1600 18250 1610 18270
rect 1630 18250 1640 18270
rect 1600 18240 1640 18250
rect 1680 18430 1720 18440
rect 1680 18410 1690 18430
rect 1710 18410 1720 18430
rect 1680 18270 1720 18410
rect 1680 18250 1690 18270
rect 1710 18250 1720 18270
rect 1680 18240 1720 18250
rect 1760 18430 1800 18440
rect 1760 18410 1770 18430
rect 1790 18410 1800 18430
rect 1760 18270 1800 18410
rect 1760 18250 1770 18270
rect 1790 18250 1800 18270
rect 1760 18240 1800 18250
rect 1840 18430 1880 18440
rect 1840 18410 1850 18430
rect 1870 18410 1880 18430
rect 1840 18270 1880 18410
rect 1840 18250 1850 18270
rect 1870 18250 1880 18270
rect 1840 18240 1880 18250
rect 1920 18430 1960 18440
rect 1920 18410 1930 18430
rect 1950 18410 1960 18430
rect 1920 18270 1960 18410
rect 1920 18250 1930 18270
rect 1950 18250 1960 18270
rect 1920 18240 1960 18250
rect 2000 18430 2040 18440
rect 2000 18410 2010 18430
rect 2030 18410 2040 18430
rect 2000 18270 2040 18410
rect 2000 18250 2010 18270
rect 2030 18250 2040 18270
rect 2000 18240 2040 18250
rect 2080 18430 2120 18440
rect 2080 18410 2090 18430
rect 2110 18410 2120 18430
rect 2080 18270 2120 18410
rect 2080 18250 2090 18270
rect 2110 18250 2120 18270
rect 2080 18240 2120 18250
rect 2160 18430 2200 18440
rect 2160 18410 2170 18430
rect 2190 18410 2200 18430
rect 2160 18270 2200 18410
rect 2160 18250 2170 18270
rect 2190 18250 2200 18270
rect 2160 18240 2200 18250
rect 2240 18430 2280 18440
rect 2240 18410 2250 18430
rect 2270 18410 2280 18430
rect 2240 18270 2280 18410
rect 2240 18250 2250 18270
rect 2270 18250 2280 18270
rect 2240 18240 2280 18250
rect 2320 18430 2360 18440
rect 2320 18410 2330 18430
rect 2350 18410 2360 18430
rect 2320 18270 2360 18410
rect 2320 18250 2330 18270
rect 2350 18250 2360 18270
rect 2320 18240 2360 18250
rect 2400 18430 2440 18440
rect 2400 18410 2410 18430
rect 2430 18410 2440 18430
rect 2400 18270 2440 18410
rect 2400 18250 2410 18270
rect 2430 18250 2440 18270
rect 2400 18240 2440 18250
rect 2480 18430 2520 18440
rect 2480 18410 2490 18430
rect 2510 18410 2520 18430
rect 2480 18270 2520 18410
rect 2480 18250 2490 18270
rect 2510 18250 2520 18270
rect 2480 18240 2520 18250
rect 2560 18430 2600 18440
rect 2560 18410 2570 18430
rect 2590 18410 2600 18430
rect 2560 18270 2600 18410
rect 2560 18250 2570 18270
rect 2590 18250 2600 18270
rect 2560 18240 2600 18250
rect 2640 18430 2680 18440
rect 2640 18410 2650 18430
rect 2670 18410 2680 18430
rect 2640 18270 2680 18410
rect 2640 18250 2650 18270
rect 2670 18250 2680 18270
rect 2640 18240 2680 18250
rect 2720 18430 2760 18440
rect 2720 18410 2730 18430
rect 2750 18410 2760 18430
rect 2720 18270 2760 18410
rect 2720 18250 2730 18270
rect 2750 18250 2760 18270
rect 2720 18240 2760 18250
rect 2800 18430 2840 18440
rect 2800 18410 2810 18430
rect 2830 18410 2840 18430
rect 2800 18270 2840 18410
rect 2800 18250 2810 18270
rect 2830 18250 2840 18270
rect 2800 18240 2840 18250
rect 2880 18430 2920 18440
rect 2880 18410 2890 18430
rect 2910 18410 2920 18430
rect 2880 18270 2920 18410
rect 2880 18250 2890 18270
rect 2910 18250 2920 18270
rect 2880 18240 2920 18250
rect 2960 18430 3000 18440
rect 2960 18410 2970 18430
rect 2990 18410 3000 18430
rect 2960 18270 3000 18410
rect 2960 18250 2970 18270
rect 2990 18250 3000 18270
rect 2960 18240 3000 18250
rect 3040 18430 3080 18440
rect 3040 18410 3050 18430
rect 3070 18410 3080 18430
rect 3040 18270 3080 18410
rect 3040 18250 3050 18270
rect 3070 18250 3080 18270
rect 3040 18240 3080 18250
rect 3120 18430 3160 18440
rect 3120 18410 3130 18430
rect 3150 18410 3160 18430
rect 3120 18270 3160 18410
rect 3120 18250 3130 18270
rect 3150 18250 3160 18270
rect 3120 18240 3160 18250
rect 3200 18430 3240 18440
rect 3200 18410 3210 18430
rect 3230 18410 3240 18430
rect 3200 18270 3240 18410
rect 3200 18250 3210 18270
rect 3230 18250 3240 18270
rect 3200 18240 3240 18250
rect 3280 18430 3320 18440
rect 3280 18410 3290 18430
rect 3310 18410 3320 18430
rect 3280 18270 3320 18410
rect 3280 18250 3290 18270
rect 3310 18250 3320 18270
rect 3280 18240 3320 18250
rect 3360 18430 3400 18440
rect 3360 18410 3370 18430
rect 3390 18410 3400 18430
rect 3360 18270 3400 18410
rect 3360 18250 3370 18270
rect 3390 18250 3400 18270
rect 3360 18240 3400 18250
rect 3440 18430 3480 18440
rect 3440 18410 3450 18430
rect 3470 18410 3480 18430
rect 3440 18270 3480 18410
rect 3440 18250 3450 18270
rect 3470 18250 3480 18270
rect 3440 18240 3480 18250
rect 3520 18430 3560 18440
rect 3520 18410 3530 18430
rect 3550 18410 3560 18430
rect 3520 18270 3560 18410
rect 3520 18250 3530 18270
rect 3550 18250 3560 18270
rect 3520 18240 3560 18250
rect 3600 18430 3640 18440
rect 3600 18410 3610 18430
rect 3630 18410 3640 18430
rect 3600 18270 3640 18410
rect 3600 18250 3610 18270
rect 3630 18250 3640 18270
rect 3600 18240 3640 18250
rect 3680 18430 3720 18440
rect 3680 18410 3690 18430
rect 3710 18410 3720 18430
rect 3680 18270 3720 18410
rect 3680 18250 3690 18270
rect 3710 18250 3720 18270
rect 3680 18240 3720 18250
rect 3760 18430 3800 18440
rect 3760 18410 3770 18430
rect 3790 18410 3800 18430
rect 3760 18270 3800 18410
rect 3760 18250 3770 18270
rect 3790 18250 3800 18270
rect 3760 18240 3800 18250
rect 3840 18430 3880 18440
rect 3840 18410 3850 18430
rect 3870 18410 3880 18430
rect 3840 18270 3880 18410
rect 3840 18250 3850 18270
rect 3870 18250 3880 18270
rect 3840 18240 3880 18250
rect 3920 18430 3960 18440
rect 3920 18410 3930 18430
rect 3950 18410 3960 18430
rect 3920 18270 3960 18410
rect 3920 18250 3930 18270
rect 3950 18250 3960 18270
rect 3920 18240 3960 18250
rect 4000 18430 4040 18440
rect 4000 18410 4010 18430
rect 4030 18410 4040 18430
rect 4000 18270 4040 18410
rect 4000 18250 4010 18270
rect 4030 18250 4040 18270
rect 4000 18240 4040 18250
rect 4080 18430 4120 18440
rect 4080 18410 4090 18430
rect 4110 18410 4120 18430
rect 4080 18270 4120 18410
rect 4080 18250 4090 18270
rect 4110 18250 4120 18270
rect 4080 18240 4120 18250
rect 4160 18430 4200 18440
rect 4160 18410 4170 18430
rect 4190 18410 4200 18430
rect 4160 18270 4200 18410
rect 4160 18250 4170 18270
rect 4190 18250 4200 18270
rect 4160 18240 4200 18250
rect 4240 18240 4280 18440
rect 4320 18240 4360 18440
rect 4400 18240 4440 18440
rect 4480 18240 4520 18440
rect 4560 18240 4600 18440
rect 4640 18240 4680 18440
rect 4720 18240 4760 18440
rect 4800 18240 4840 18440
rect 4880 18240 4920 18440
rect 4960 18240 5000 18440
rect 5040 18240 5080 18440
rect 5120 18240 5160 18440
rect 5200 18240 5240 18440
rect 5280 18240 5320 18440
rect 5360 18240 5400 18440
rect 5440 18240 5480 18440
rect 5520 18240 5560 18440
rect 5600 18240 5640 18440
rect 5680 18240 5720 18440
rect 5760 18240 5800 18440
rect 5840 18240 5880 18440
rect 5920 18240 5960 18440
rect 6000 18240 6040 18440
rect 6080 18240 6120 18440
rect 6160 18240 6200 18440
rect 6240 18430 6280 18440
rect 6240 18410 6250 18430
rect 6270 18410 6280 18430
rect 6240 18270 6280 18410
rect 6240 18250 6250 18270
rect 6270 18250 6280 18270
rect 6240 18240 6280 18250
rect 6320 18430 6360 18440
rect 6320 18410 6330 18430
rect 6350 18410 6360 18430
rect 6320 18270 6360 18410
rect 6320 18250 6330 18270
rect 6350 18250 6360 18270
rect 6320 18240 6360 18250
rect 6400 18430 6440 18440
rect 6400 18410 6410 18430
rect 6430 18410 6440 18430
rect 6400 18270 6440 18410
rect 6400 18250 6410 18270
rect 6430 18250 6440 18270
rect 6400 18240 6440 18250
rect 6480 18430 6520 18440
rect 6480 18410 6490 18430
rect 6510 18410 6520 18430
rect 6480 18270 6520 18410
rect 6480 18250 6490 18270
rect 6510 18250 6520 18270
rect 6480 18240 6520 18250
rect 6560 18430 6600 18440
rect 6560 18410 6570 18430
rect 6590 18410 6600 18430
rect 6560 18270 6600 18410
rect 6560 18250 6570 18270
rect 6590 18250 6600 18270
rect 6560 18240 6600 18250
rect 6640 18430 6680 18440
rect 6640 18410 6650 18430
rect 6670 18410 6680 18430
rect 6640 18270 6680 18410
rect 6640 18250 6650 18270
rect 6670 18250 6680 18270
rect 6640 18240 6680 18250
rect 6720 18430 6760 18440
rect 6720 18410 6730 18430
rect 6750 18410 6760 18430
rect 6720 18270 6760 18410
rect 6720 18250 6730 18270
rect 6750 18250 6760 18270
rect 6720 18240 6760 18250
rect 6800 18430 6840 18440
rect 6800 18410 6810 18430
rect 6830 18410 6840 18430
rect 6800 18270 6840 18410
rect 6800 18250 6810 18270
rect 6830 18250 6840 18270
rect 6800 18240 6840 18250
rect 6880 18430 6920 18440
rect 6880 18410 6890 18430
rect 6910 18410 6920 18430
rect 6880 18270 6920 18410
rect 6880 18250 6890 18270
rect 6910 18250 6920 18270
rect 6880 18240 6920 18250
rect 6960 18430 7000 18440
rect 6960 18410 6970 18430
rect 6990 18410 7000 18430
rect 6960 18270 7000 18410
rect 6960 18250 6970 18270
rect 6990 18250 7000 18270
rect 6960 18240 7000 18250
rect 7040 18430 7080 18440
rect 7040 18410 7050 18430
rect 7070 18410 7080 18430
rect 7040 18270 7080 18410
rect 7040 18250 7050 18270
rect 7070 18250 7080 18270
rect 7040 18240 7080 18250
rect 7120 18430 7160 18440
rect 7120 18410 7130 18430
rect 7150 18410 7160 18430
rect 7120 18270 7160 18410
rect 7120 18250 7130 18270
rect 7150 18250 7160 18270
rect 7120 18240 7160 18250
rect 7200 18430 7240 18440
rect 7200 18410 7210 18430
rect 7230 18410 7240 18430
rect 7200 18270 7240 18410
rect 7200 18250 7210 18270
rect 7230 18250 7240 18270
rect 7200 18240 7240 18250
rect 7280 18430 7320 18440
rect 7280 18410 7290 18430
rect 7310 18410 7320 18430
rect 7280 18270 7320 18410
rect 7280 18250 7290 18270
rect 7310 18250 7320 18270
rect 7280 18240 7320 18250
rect 7360 18430 7400 18440
rect 7360 18410 7370 18430
rect 7390 18410 7400 18430
rect 7360 18270 7400 18410
rect 7360 18250 7370 18270
rect 7390 18250 7400 18270
rect 7360 18240 7400 18250
rect 7440 18430 7480 18440
rect 7440 18410 7450 18430
rect 7470 18410 7480 18430
rect 7440 18270 7480 18410
rect 7440 18250 7450 18270
rect 7470 18250 7480 18270
rect 7440 18240 7480 18250
rect 7520 18430 7560 18440
rect 7520 18410 7530 18430
rect 7550 18410 7560 18430
rect 7520 18270 7560 18410
rect 7520 18250 7530 18270
rect 7550 18250 7560 18270
rect 7520 18240 7560 18250
rect 7600 18430 7640 18440
rect 7600 18410 7610 18430
rect 7630 18410 7640 18430
rect 7600 18270 7640 18410
rect 7600 18250 7610 18270
rect 7630 18250 7640 18270
rect 7600 18240 7640 18250
rect 7680 18430 7720 18440
rect 7680 18410 7690 18430
rect 7710 18410 7720 18430
rect 7680 18270 7720 18410
rect 7680 18250 7690 18270
rect 7710 18250 7720 18270
rect 7680 18240 7720 18250
rect 7760 18430 7800 18440
rect 7760 18410 7770 18430
rect 7790 18410 7800 18430
rect 7760 18270 7800 18410
rect 7760 18250 7770 18270
rect 7790 18250 7800 18270
rect 7760 18240 7800 18250
rect 7840 18430 7880 18440
rect 7840 18410 7850 18430
rect 7870 18410 7880 18430
rect 7840 18270 7880 18410
rect 7840 18250 7850 18270
rect 7870 18250 7880 18270
rect 7840 18240 7880 18250
rect 7920 18430 7960 18440
rect 7920 18410 7930 18430
rect 7950 18410 7960 18430
rect 7920 18270 7960 18410
rect 7920 18250 7930 18270
rect 7950 18250 7960 18270
rect 7920 18240 7960 18250
rect 8000 18430 8040 18440
rect 8000 18410 8010 18430
rect 8030 18410 8040 18430
rect 8000 18270 8040 18410
rect 8000 18250 8010 18270
rect 8030 18250 8040 18270
rect 8000 18240 8040 18250
rect 8080 18430 8120 18440
rect 8080 18410 8090 18430
rect 8110 18410 8120 18430
rect 8080 18270 8120 18410
rect 8080 18250 8090 18270
rect 8110 18250 8120 18270
rect 8080 18240 8120 18250
rect 8160 18430 8200 18440
rect 8160 18410 8170 18430
rect 8190 18410 8200 18430
rect 8160 18270 8200 18410
rect 8160 18250 8170 18270
rect 8190 18250 8200 18270
rect 8160 18240 8200 18250
rect 8240 18430 8280 18440
rect 8240 18410 8250 18430
rect 8270 18410 8280 18430
rect 8240 18270 8280 18410
rect 8240 18250 8250 18270
rect 8270 18250 8280 18270
rect 8240 18240 8280 18250
rect 8320 18430 8360 18440
rect 8320 18410 8330 18430
rect 8350 18410 8360 18430
rect 8320 18270 8360 18410
rect 8320 18250 8330 18270
rect 8350 18250 8360 18270
rect 8320 18240 8360 18250
rect 8400 18430 8440 18440
rect 8400 18410 8410 18430
rect 8430 18410 8440 18430
rect 8400 18270 8440 18410
rect 8400 18250 8410 18270
rect 8430 18250 8440 18270
rect 8400 18240 8440 18250
rect 8480 18430 8520 18440
rect 8480 18410 8490 18430
rect 8510 18410 8520 18430
rect 8480 18270 8520 18410
rect 8480 18250 8490 18270
rect 8510 18250 8520 18270
rect 8480 18240 8520 18250
rect 8560 18430 8600 18440
rect 8560 18410 8570 18430
rect 8590 18410 8600 18430
rect 8560 18270 8600 18410
rect 8560 18250 8570 18270
rect 8590 18250 8600 18270
rect 8560 18240 8600 18250
rect 8640 18430 8680 18440
rect 8640 18410 8650 18430
rect 8670 18410 8680 18430
rect 8640 18270 8680 18410
rect 8640 18250 8650 18270
rect 8670 18250 8680 18270
rect 8640 18240 8680 18250
rect 8720 18430 8760 18440
rect 8720 18410 8730 18430
rect 8750 18410 8760 18430
rect 8720 18270 8760 18410
rect 8720 18250 8730 18270
rect 8750 18250 8760 18270
rect 8720 18240 8760 18250
rect 8800 18430 8840 18440
rect 8800 18410 8810 18430
rect 8830 18410 8840 18430
rect 8800 18270 8840 18410
rect 8800 18250 8810 18270
rect 8830 18250 8840 18270
rect 8800 18240 8840 18250
rect 8880 18430 8920 18440
rect 8880 18410 8890 18430
rect 8910 18410 8920 18430
rect 8880 18270 8920 18410
rect 8880 18250 8890 18270
rect 8910 18250 8920 18270
rect 8880 18240 8920 18250
rect 8960 18430 9000 18440
rect 8960 18410 8970 18430
rect 8990 18410 9000 18430
rect 8960 18270 9000 18410
rect 8960 18250 8970 18270
rect 8990 18250 9000 18270
rect 8960 18240 9000 18250
rect 9040 18430 9080 18440
rect 9040 18410 9050 18430
rect 9070 18410 9080 18430
rect 9040 18270 9080 18410
rect 9040 18250 9050 18270
rect 9070 18250 9080 18270
rect 9040 18240 9080 18250
rect 9120 18430 9160 18440
rect 9120 18410 9130 18430
rect 9150 18410 9160 18430
rect 9120 18270 9160 18410
rect 9120 18250 9130 18270
rect 9150 18250 9160 18270
rect 9120 18240 9160 18250
rect 9200 18430 9240 18440
rect 9200 18410 9210 18430
rect 9230 18410 9240 18430
rect 9200 18270 9240 18410
rect 9200 18250 9210 18270
rect 9230 18250 9240 18270
rect 9200 18240 9240 18250
rect 9280 18430 9320 18440
rect 9280 18410 9290 18430
rect 9310 18410 9320 18430
rect 9280 18270 9320 18410
rect 9280 18250 9290 18270
rect 9310 18250 9320 18270
rect 9280 18240 9320 18250
rect 9360 18430 9400 18440
rect 9360 18410 9370 18430
rect 9390 18410 9400 18430
rect 9360 18270 9400 18410
rect 9360 18250 9370 18270
rect 9390 18250 9400 18270
rect 9360 18240 9400 18250
rect 9440 18430 9480 18440
rect 9440 18410 9450 18430
rect 9470 18410 9480 18430
rect 9440 18270 9480 18410
rect 9440 18250 9450 18270
rect 9470 18250 9480 18270
rect 9440 18240 9480 18250
rect 9520 18240 9560 18440
rect 9600 18240 9640 18440
rect 9680 18240 9720 18440
rect 9760 18240 9800 18440
rect 9840 18240 9880 18440
rect 9920 18240 9960 18440
rect 10000 18240 10040 18440
rect 10080 18240 10120 18440
rect 10160 18240 10200 18440
rect 10240 18240 10280 18440
rect 10320 18240 10360 18440
rect 10400 18240 10440 18440
rect 10480 18240 10520 18440
rect 10560 18240 10600 18440
rect 10640 18240 10680 18440
rect 10720 18240 10760 18440
rect 10800 18240 10840 18440
rect 10880 18240 10920 18440
rect 10960 18240 11000 18440
rect 11040 18240 11080 18440
rect 11120 18240 11160 18440
rect 11200 18240 11240 18440
rect 11280 18240 11320 18440
rect 11360 18240 11400 18440
rect 11440 18240 11480 18440
rect 11560 18430 11600 18440
rect 11560 18410 11570 18430
rect 11590 18410 11600 18430
rect 11560 18270 11600 18410
rect 11560 18250 11570 18270
rect 11590 18250 11600 18270
rect 11560 18240 11600 18250
rect 11640 18430 11680 18440
rect 11640 18410 11650 18430
rect 11670 18410 11680 18430
rect 11640 18270 11680 18410
rect 11640 18250 11650 18270
rect 11670 18250 11680 18270
rect 11640 18240 11680 18250
rect 11720 18430 11760 18440
rect 11720 18410 11730 18430
rect 11750 18410 11760 18430
rect 11720 18270 11760 18410
rect 11720 18250 11730 18270
rect 11750 18250 11760 18270
rect 11720 18240 11760 18250
rect 11800 18430 11840 18440
rect 11800 18410 11810 18430
rect 11830 18410 11840 18430
rect 11800 18270 11840 18410
rect 11800 18250 11810 18270
rect 11830 18250 11840 18270
rect 11800 18240 11840 18250
rect 11880 18430 11920 18440
rect 11880 18410 11890 18430
rect 11910 18410 11920 18430
rect 11880 18270 11920 18410
rect 11880 18250 11890 18270
rect 11910 18250 11920 18270
rect 11880 18240 11920 18250
rect 11960 18430 12000 18440
rect 11960 18410 11970 18430
rect 11990 18410 12000 18430
rect 11960 18270 12000 18410
rect 11960 18250 11970 18270
rect 11990 18250 12000 18270
rect 11960 18240 12000 18250
rect 12040 18430 12080 18440
rect 12040 18410 12050 18430
rect 12070 18410 12080 18430
rect 12040 18270 12080 18410
rect 12040 18250 12050 18270
rect 12070 18250 12080 18270
rect 12040 18240 12080 18250
rect 12120 18430 12160 18440
rect 12120 18410 12130 18430
rect 12150 18410 12160 18430
rect 12120 18270 12160 18410
rect 12120 18250 12130 18270
rect 12150 18250 12160 18270
rect 12120 18240 12160 18250
rect 12200 18430 12240 18440
rect 12200 18410 12210 18430
rect 12230 18410 12240 18430
rect 12200 18270 12240 18410
rect 12200 18250 12210 18270
rect 12230 18250 12240 18270
rect 12200 18240 12240 18250
rect 12280 18430 12320 18440
rect 12280 18410 12290 18430
rect 12310 18410 12320 18430
rect 12280 18270 12320 18410
rect 12280 18250 12290 18270
rect 12310 18250 12320 18270
rect 12280 18240 12320 18250
rect 12360 18430 12400 18440
rect 12360 18410 12370 18430
rect 12390 18410 12400 18430
rect 12360 18270 12400 18410
rect 12360 18250 12370 18270
rect 12390 18250 12400 18270
rect 12360 18240 12400 18250
rect 12440 18430 12480 18440
rect 12440 18410 12450 18430
rect 12470 18410 12480 18430
rect 12440 18270 12480 18410
rect 12440 18250 12450 18270
rect 12470 18250 12480 18270
rect 12440 18240 12480 18250
rect 12520 18430 12560 18440
rect 12520 18410 12530 18430
rect 12550 18410 12560 18430
rect 12520 18270 12560 18410
rect 12520 18250 12530 18270
rect 12550 18250 12560 18270
rect 12520 18240 12560 18250
rect 12600 18430 12640 18440
rect 12600 18410 12610 18430
rect 12630 18410 12640 18430
rect 12600 18270 12640 18410
rect 12600 18250 12610 18270
rect 12630 18250 12640 18270
rect 12600 18240 12640 18250
rect 12680 18430 12720 18440
rect 12680 18410 12690 18430
rect 12710 18410 12720 18430
rect 12680 18270 12720 18410
rect 12680 18250 12690 18270
rect 12710 18250 12720 18270
rect 12680 18240 12720 18250
rect 12760 18430 12800 18440
rect 12760 18410 12770 18430
rect 12790 18410 12800 18430
rect 12760 18270 12800 18410
rect 12760 18250 12770 18270
rect 12790 18250 12800 18270
rect 12760 18240 12800 18250
rect 12840 18430 12880 18440
rect 12840 18410 12850 18430
rect 12870 18410 12880 18430
rect 12840 18270 12880 18410
rect 12840 18250 12850 18270
rect 12870 18250 12880 18270
rect 12840 18240 12880 18250
rect 12920 18430 12960 18440
rect 12920 18410 12930 18430
rect 12950 18410 12960 18430
rect 12920 18270 12960 18410
rect 12920 18250 12930 18270
rect 12950 18250 12960 18270
rect 12920 18240 12960 18250
rect 13000 18430 13040 18440
rect 13000 18410 13010 18430
rect 13030 18410 13040 18430
rect 13000 18270 13040 18410
rect 13000 18250 13010 18270
rect 13030 18250 13040 18270
rect 13000 18240 13040 18250
rect 13080 18430 13120 18440
rect 13080 18410 13090 18430
rect 13110 18410 13120 18430
rect 13080 18270 13120 18410
rect 13080 18250 13090 18270
rect 13110 18250 13120 18270
rect 13080 18240 13120 18250
rect 13160 18430 13200 18440
rect 13160 18410 13170 18430
rect 13190 18410 13200 18430
rect 13160 18270 13200 18410
rect 13160 18250 13170 18270
rect 13190 18250 13200 18270
rect 13160 18240 13200 18250
rect 13240 18430 13280 18440
rect 13240 18410 13250 18430
rect 13270 18410 13280 18430
rect 13240 18270 13280 18410
rect 13240 18250 13250 18270
rect 13270 18250 13280 18270
rect 13240 18240 13280 18250
rect 13320 18430 13360 18440
rect 13320 18410 13330 18430
rect 13350 18410 13360 18430
rect 13320 18270 13360 18410
rect 13320 18250 13330 18270
rect 13350 18250 13360 18270
rect 13320 18240 13360 18250
rect 13400 18430 13440 18440
rect 13400 18410 13410 18430
rect 13430 18410 13440 18430
rect 13400 18270 13440 18410
rect 13400 18250 13410 18270
rect 13430 18250 13440 18270
rect 13400 18240 13440 18250
rect 13480 18430 13520 18440
rect 13480 18410 13490 18430
rect 13510 18410 13520 18430
rect 13480 18270 13520 18410
rect 13480 18250 13490 18270
rect 13510 18250 13520 18270
rect 13480 18240 13520 18250
rect 13560 18430 13600 18440
rect 13560 18410 13570 18430
rect 13590 18410 13600 18430
rect 13560 18270 13600 18410
rect 13560 18250 13570 18270
rect 13590 18250 13600 18270
rect 13560 18240 13600 18250
rect 13640 18430 13680 18440
rect 13640 18410 13650 18430
rect 13670 18410 13680 18430
rect 13640 18270 13680 18410
rect 13640 18250 13650 18270
rect 13670 18250 13680 18270
rect 13640 18240 13680 18250
rect 13720 18430 13760 18440
rect 13720 18410 13730 18430
rect 13750 18410 13760 18430
rect 13720 18270 13760 18410
rect 13720 18250 13730 18270
rect 13750 18250 13760 18270
rect 13720 18240 13760 18250
rect 13800 18430 13840 18440
rect 13800 18410 13810 18430
rect 13830 18410 13840 18430
rect 13800 18270 13840 18410
rect 13800 18250 13810 18270
rect 13830 18250 13840 18270
rect 13800 18240 13840 18250
rect 13880 18430 13920 18440
rect 13880 18410 13890 18430
rect 13910 18410 13920 18430
rect 13880 18270 13920 18410
rect 13880 18250 13890 18270
rect 13910 18250 13920 18270
rect 13880 18240 13920 18250
rect 13960 18430 14000 18440
rect 13960 18410 13970 18430
rect 13990 18410 14000 18430
rect 13960 18270 14000 18410
rect 13960 18250 13970 18270
rect 13990 18250 14000 18270
rect 13960 18240 14000 18250
rect 14040 18430 14080 18440
rect 14040 18410 14050 18430
rect 14070 18410 14080 18430
rect 14040 18270 14080 18410
rect 14040 18250 14050 18270
rect 14070 18250 14080 18270
rect 14040 18240 14080 18250
rect 14120 18430 14160 18440
rect 14120 18410 14130 18430
rect 14150 18410 14160 18430
rect 14120 18270 14160 18410
rect 14120 18250 14130 18270
rect 14150 18250 14160 18270
rect 14120 18240 14160 18250
rect 14200 18430 14240 18440
rect 14200 18410 14210 18430
rect 14230 18410 14240 18430
rect 14200 18270 14240 18410
rect 14200 18250 14210 18270
rect 14230 18250 14240 18270
rect 14200 18240 14240 18250
rect 14280 18430 14320 18440
rect 14280 18410 14290 18430
rect 14310 18410 14320 18430
rect 14280 18270 14320 18410
rect 14280 18250 14290 18270
rect 14310 18250 14320 18270
rect 14280 18240 14320 18250
rect 14360 18430 14400 18440
rect 14360 18410 14370 18430
rect 14390 18410 14400 18430
rect 14360 18270 14400 18410
rect 14360 18250 14370 18270
rect 14390 18250 14400 18270
rect 14360 18240 14400 18250
rect 14440 18430 14480 18440
rect 14440 18410 14450 18430
rect 14470 18410 14480 18430
rect 14440 18270 14480 18410
rect 14440 18250 14450 18270
rect 14470 18250 14480 18270
rect 14440 18240 14480 18250
rect 14520 18430 14560 18440
rect 14520 18410 14530 18430
rect 14550 18410 14560 18430
rect 14520 18270 14560 18410
rect 14520 18250 14530 18270
rect 14550 18250 14560 18270
rect 14520 18240 14560 18250
rect 14600 18430 14640 18440
rect 14600 18410 14610 18430
rect 14630 18410 14640 18430
rect 14600 18270 14640 18410
rect 14600 18250 14610 18270
rect 14630 18250 14640 18270
rect 14600 18240 14640 18250
rect 14680 18430 14720 18440
rect 14680 18410 14690 18430
rect 14710 18410 14720 18430
rect 14680 18270 14720 18410
rect 14680 18250 14690 18270
rect 14710 18250 14720 18270
rect 14680 18240 14720 18250
rect 14760 18240 14800 18440
rect 14840 18240 14880 18440
rect 14920 18240 14960 18440
rect 15000 18240 15040 18440
rect 15080 18240 15120 18440
rect 15160 18240 15200 18440
rect 15240 18240 15280 18440
rect 15320 18240 15360 18440
rect 15400 18240 15440 18440
rect 15480 18240 15520 18440
rect 15560 18240 15600 18440
rect 15640 18240 15680 18440
rect 15720 18240 15760 18440
rect 15800 18240 15840 18440
rect 15880 18240 15920 18440
rect 15960 18240 16000 18440
rect 16040 18240 16080 18440
rect 16120 18240 16160 18440
rect 16200 18240 16240 18440
rect 16280 18240 16320 18440
rect 16360 18240 16400 18440
rect 16440 18240 16480 18440
rect 16520 18240 16560 18440
rect 16600 18240 16640 18440
rect 16680 18240 16720 18440
rect 16760 18430 16800 18440
rect 16760 18410 16770 18430
rect 16790 18410 16800 18430
rect 16760 18270 16800 18410
rect 16760 18250 16770 18270
rect 16790 18250 16800 18270
rect 16760 18240 16800 18250
rect 16840 18430 16880 18440
rect 16840 18410 16850 18430
rect 16870 18410 16880 18430
rect 16840 18270 16880 18410
rect 16840 18250 16850 18270
rect 16870 18250 16880 18270
rect 16840 18240 16880 18250
rect 16920 18430 16960 18440
rect 16920 18410 16930 18430
rect 16950 18410 16960 18430
rect 16920 18270 16960 18410
rect 16920 18250 16930 18270
rect 16950 18250 16960 18270
rect 16920 18240 16960 18250
rect 17000 18430 17040 18440
rect 17000 18410 17010 18430
rect 17030 18410 17040 18430
rect 17000 18270 17040 18410
rect 17000 18250 17010 18270
rect 17030 18250 17040 18270
rect 17000 18240 17040 18250
rect 17080 18430 17120 18440
rect 17080 18410 17090 18430
rect 17110 18410 17120 18430
rect 17080 18270 17120 18410
rect 17080 18250 17090 18270
rect 17110 18250 17120 18270
rect 17080 18240 17120 18250
rect 17160 18430 17200 18440
rect 17160 18410 17170 18430
rect 17190 18410 17200 18430
rect 17160 18270 17200 18410
rect 17160 18250 17170 18270
rect 17190 18250 17200 18270
rect 17160 18240 17200 18250
rect 17240 18430 17280 18440
rect 17240 18410 17250 18430
rect 17270 18410 17280 18430
rect 17240 18270 17280 18410
rect 17240 18250 17250 18270
rect 17270 18250 17280 18270
rect 17240 18240 17280 18250
rect 17320 18430 17360 18440
rect 17320 18410 17330 18430
rect 17350 18410 17360 18430
rect 17320 18270 17360 18410
rect 17320 18250 17330 18270
rect 17350 18250 17360 18270
rect 17320 18240 17360 18250
rect 17400 18430 17440 18440
rect 17400 18410 17410 18430
rect 17430 18410 17440 18430
rect 17400 18270 17440 18410
rect 17400 18250 17410 18270
rect 17430 18250 17440 18270
rect 17400 18240 17440 18250
rect 17480 18430 17520 18440
rect 17480 18410 17490 18430
rect 17510 18410 17520 18430
rect 17480 18270 17520 18410
rect 17480 18250 17490 18270
rect 17510 18250 17520 18270
rect 17480 18240 17520 18250
rect 17560 18430 17600 18440
rect 17560 18410 17570 18430
rect 17590 18410 17600 18430
rect 17560 18270 17600 18410
rect 17560 18250 17570 18270
rect 17590 18250 17600 18270
rect 17560 18240 17600 18250
rect 17640 18430 17680 18440
rect 17640 18410 17650 18430
rect 17670 18410 17680 18430
rect 17640 18270 17680 18410
rect 17640 18250 17650 18270
rect 17670 18250 17680 18270
rect 17640 18240 17680 18250
rect 17720 18430 17760 18440
rect 17720 18410 17730 18430
rect 17750 18410 17760 18430
rect 17720 18270 17760 18410
rect 17720 18250 17730 18270
rect 17750 18250 17760 18270
rect 17720 18240 17760 18250
rect 17800 18430 17840 18440
rect 17800 18410 17810 18430
rect 17830 18410 17840 18430
rect 17800 18270 17840 18410
rect 17800 18250 17810 18270
rect 17830 18250 17840 18270
rect 17800 18240 17840 18250
rect 17880 18430 17920 18440
rect 17880 18410 17890 18430
rect 17910 18410 17920 18430
rect 17880 18270 17920 18410
rect 17880 18250 17890 18270
rect 17910 18250 17920 18270
rect 17880 18240 17920 18250
rect 17960 18430 18000 18440
rect 17960 18410 17970 18430
rect 17990 18410 18000 18430
rect 17960 18270 18000 18410
rect 17960 18250 17970 18270
rect 17990 18250 18000 18270
rect 17960 18240 18000 18250
rect 18040 18430 18080 18440
rect 18040 18410 18050 18430
rect 18070 18410 18080 18430
rect 18040 18270 18080 18410
rect 18040 18250 18050 18270
rect 18070 18250 18080 18270
rect 18040 18240 18080 18250
rect 18120 18430 18160 18440
rect 18120 18410 18130 18430
rect 18150 18410 18160 18430
rect 18120 18270 18160 18410
rect 18120 18250 18130 18270
rect 18150 18250 18160 18270
rect 18120 18240 18160 18250
rect 18200 18430 18240 18440
rect 18200 18410 18210 18430
rect 18230 18410 18240 18430
rect 18200 18270 18240 18410
rect 18200 18250 18210 18270
rect 18230 18250 18240 18270
rect 18200 18240 18240 18250
rect 18280 18430 18320 18440
rect 18280 18410 18290 18430
rect 18310 18410 18320 18430
rect 18280 18270 18320 18410
rect 18280 18250 18290 18270
rect 18310 18250 18320 18270
rect 18280 18240 18320 18250
rect 18360 18430 18400 18440
rect 18360 18410 18370 18430
rect 18390 18410 18400 18430
rect 18360 18270 18400 18410
rect 18360 18250 18370 18270
rect 18390 18250 18400 18270
rect 18360 18240 18400 18250
rect 18440 18430 18480 18440
rect 18440 18410 18450 18430
rect 18470 18410 18480 18430
rect 18440 18270 18480 18410
rect 18440 18250 18450 18270
rect 18470 18250 18480 18270
rect 18440 18240 18480 18250
rect 18520 18430 18560 18440
rect 18520 18410 18530 18430
rect 18550 18410 18560 18430
rect 18520 18270 18560 18410
rect 18520 18250 18530 18270
rect 18550 18250 18560 18270
rect 18520 18240 18560 18250
rect 18600 18430 18640 18440
rect 18600 18410 18610 18430
rect 18630 18410 18640 18430
rect 18600 18270 18640 18410
rect 18600 18250 18610 18270
rect 18630 18250 18640 18270
rect 18600 18240 18640 18250
rect 18680 18430 18720 18440
rect 18680 18410 18690 18430
rect 18710 18410 18720 18430
rect 18680 18270 18720 18410
rect 18680 18250 18690 18270
rect 18710 18250 18720 18270
rect 18680 18240 18720 18250
rect 18760 18430 18800 18440
rect 18760 18410 18770 18430
rect 18790 18410 18800 18430
rect 18760 18270 18800 18410
rect 18760 18250 18770 18270
rect 18790 18250 18800 18270
rect 18760 18240 18800 18250
rect 18840 18430 18880 18440
rect 18840 18410 18850 18430
rect 18870 18410 18880 18430
rect 18840 18270 18880 18410
rect 18840 18250 18850 18270
rect 18870 18250 18880 18270
rect 18840 18240 18880 18250
rect 18920 18430 18960 18440
rect 18920 18410 18930 18430
rect 18950 18410 18960 18430
rect 18920 18270 18960 18410
rect 18920 18250 18930 18270
rect 18950 18250 18960 18270
rect 18920 18240 18960 18250
rect 19000 18430 19040 18440
rect 19000 18410 19010 18430
rect 19030 18410 19040 18430
rect 19000 18270 19040 18410
rect 19000 18250 19010 18270
rect 19030 18250 19040 18270
rect 19000 18240 19040 18250
rect 19080 18430 19120 18440
rect 19080 18410 19090 18430
rect 19110 18410 19120 18430
rect 19080 18270 19120 18410
rect 19080 18250 19090 18270
rect 19110 18250 19120 18270
rect 19080 18240 19120 18250
rect 19160 18430 19200 18440
rect 19160 18410 19170 18430
rect 19190 18410 19200 18430
rect 19160 18270 19200 18410
rect 19160 18250 19170 18270
rect 19190 18250 19200 18270
rect 19160 18240 19200 18250
rect 19240 18430 19280 18440
rect 19240 18410 19250 18430
rect 19270 18410 19280 18430
rect 19240 18270 19280 18410
rect 19240 18250 19250 18270
rect 19270 18250 19280 18270
rect 19240 18240 19280 18250
rect 19320 18430 19360 18440
rect 19320 18410 19330 18430
rect 19350 18410 19360 18430
rect 19320 18270 19360 18410
rect 19320 18250 19330 18270
rect 19350 18250 19360 18270
rect 19320 18240 19360 18250
rect 19400 18430 19440 18440
rect 19400 18410 19410 18430
rect 19430 18410 19440 18430
rect 19400 18270 19440 18410
rect 19400 18250 19410 18270
rect 19430 18250 19440 18270
rect 19400 18240 19440 18250
rect 19480 18430 19520 18440
rect 19480 18410 19490 18430
rect 19510 18410 19520 18430
rect 19480 18270 19520 18410
rect 19480 18250 19490 18270
rect 19510 18250 19520 18270
rect 19480 18240 19520 18250
rect 19560 18430 19600 18440
rect 19560 18410 19570 18430
rect 19590 18410 19600 18430
rect 19560 18270 19600 18410
rect 19560 18250 19570 18270
rect 19590 18250 19600 18270
rect 19560 18240 19600 18250
rect 19640 18430 19680 18440
rect 19640 18410 19650 18430
rect 19670 18410 19680 18430
rect 19640 18270 19680 18410
rect 19640 18250 19650 18270
rect 19670 18250 19680 18270
rect 19640 18240 19680 18250
rect 19720 18430 19760 18440
rect 19720 18410 19730 18430
rect 19750 18410 19760 18430
rect 19720 18270 19760 18410
rect 19720 18250 19730 18270
rect 19750 18250 19760 18270
rect 19720 18240 19760 18250
rect 19800 18430 19840 18440
rect 19800 18410 19810 18430
rect 19830 18410 19840 18430
rect 19800 18270 19840 18410
rect 19800 18250 19810 18270
rect 19830 18250 19840 18270
rect 19800 18240 19840 18250
rect 19880 18430 19920 18440
rect 19880 18410 19890 18430
rect 19910 18410 19920 18430
rect 19880 18270 19920 18410
rect 19880 18250 19890 18270
rect 19910 18250 19920 18270
rect 19880 18240 19920 18250
rect 19960 18430 20000 18440
rect 19960 18410 19970 18430
rect 19990 18410 20000 18430
rect 19960 18270 20000 18410
rect 19960 18250 19970 18270
rect 19990 18250 20000 18270
rect 19960 18240 20000 18250
rect 20040 18430 20080 18440
rect 20040 18410 20050 18430
rect 20070 18410 20080 18430
rect 20040 18270 20080 18410
rect 20040 18250 20050 18270
rect 20070 18250 20080 18270
rect 20040 18240 20080 18250
rect 20120 18430 20160 18440
rect 20120 18410 20130 18430
rect 20150 18410 20160 18430
rect 20120 18270 20160 18410
rect 20120 18250 20130 18270
rect 20150 18250 20160 18270
rect 20120 18240 20160 18250
rect 20200 18430 20240 18440
rect 20200 18410 20210 18430
rect 20230 18410 20240 18430
rect 20200 18270 20240 18410
rect 20200 18250 20210 18270
rect 20230 18250 20240 18270
rect 20200 18240 20240 18250
rect 20280 18430 20320 18440
rect 20280 18410 20290 18430
rect 20310 18410 20320 18430
rect 20280 18270 20320 18410
rect 20280 18250 20290 18270
rect 20310 18250 20320 18270
rect 20280 18240 20320 18250
rect 20360 18430 20400 18440
rect 20360 18410 20370 18430
rect 20390 18410 20400 18430
rect 20360 18270 20400 18410
rect 20360 18250 20370 18270
rect 20390 18250 20400 18270
rect 20360 18240 20400 18250
rect 20440 18430 20480 18440
rect 20440 18410 20450 18430
rect 20470 18410 20480 18430
rect 20440 18270 20480 18410
rect 20440 18250 20450 18270
rect 20470 18250 20480 18270
rect 20440 18240 20480 18250
rect 20520 18430 20560 18440
rect 20520 18410 20530 18430
rect 20550 18410 20560 18430
rect 20520 18270 20560 18410
rect 20520 18250 20530 18270
rect 20550 18250 20560 18270
rect 20520 18240 20560 18250
rect 20600 18430 20640 18440
rect 20600 18410 20610 18430
rect 20630 18410 20640 18430
rect 20600 18270 20640 18410
rect 20600 18250 20610 18270
rect 20630 18250 20640 18270
rect 20600 18240 20640 18250
rect 20680 18430 20720 18440
rect 20680 18410 20690 18430
rect 20710 18410 20720 18430
rect 20680 18270 20720 18410
rect 20680 18250 20690 18270
rect 20710 18250 20720 18270
rect 20680 18240 20720 18250
rect 20760 18430 20800 18440
rect 20760 18410 20770 18430
rect 20790 18410 20800 18430
rect 20760 18270 20800 18410
rect 20760 18250 20770 18270
rect 20790 18250 20800 18270
rect 20760 18240 20800 18250
rect 20840 18430 20880 18440
rect 20840 18410 20850 18430
rect 20870 18410 20880 18430
rect 20840 18270 20880 18410
rect 20840 18250 20850 18270
rect 20870 18250 20880 18270
rect 20840 18240 20880 18250
rect 20920 18430 20960 18440
rect 20920 18410 20930 18430
rect 20950 18410 20960 18430
rect 20920 18270 20960 18410
rect 20920 18250 20930 18270
rect 20950 18250 20960 18270
rect 20920 18240 20960 18250
rect 0 18190 40 18200
rect 0 18170 10 18190
rect 30 18170 40 18190
rect 0 18030 40 18170
rect 0 18010 10 18030
rect 30 18010 40 18030
rect 0 17870 40 18010
rect 0 17850 10 17870
rect 30 17850 40 17870
rect 0 17710 40 17850
rect 0 17690 10 17710
rect 30 17690 40 17710
rect 0 17550 40 17690
rect 0 17530 10 17550
rect 30 17530 40 17550
rect 0 17390 40 17530
rect 0 17370 10 17390
rect 30 17370 40 17390
rect 0 17230 40 17370
rect 0 17210 10 17230
rect 30 17210 40 17230
rect 0 17200 40 17210
rect 80 18190 120 18200
rect 80 18170 90 18190
rect 110 18170 120 18190
rect 80 18030 120 18170
rect 80 18010 90 18030
rect 110 18010 120 18030
rect 80 17870 120 18010
rect 80 17850 90 17870
rect 110 17850 120 17870
rect 80 17710 120 17850
rect 80 17690 90 17710
rect 110 17690 120 17710
rect 80 17550 120 17690
rect 80 17530 90 17550
rect 110 17530 120 17550
rect 80 17390 120 17530
rect 80 17370 90 17390
rect 110 17370 120 17390
rect 80 17230 120 17370
rect 80 17210 90 17230
rect 110 17210 120 17230
rect 80 17200 120 17210
rect 160 18190 200 18200
rect 160 18170 170 18190
rect 190 18170 200 18190
rect 160 18030 200 18170
rect 160 18010 170 18030
rect 190 18010 200 18030
rect 160 17870 200 18010
rect 160 17850 170 17870
rect 190 17850 200 17870
rect 160 17710 200 17850
rect 160 17690 170 17710
rect 190 17690 200 17710
rect 160 17550 200 17690
rect 160 17530 170 17550
rect 190 17530 200 17550
rect 160 17390 200 17530
rect 160 17370 170 17390
rect 190 17370 200 17390
rect 160 17230 200 17370
rect 160 17210 170 17230
rect 190 17210 200 17230
rect 160 17200 200 17210
rect 240 18190 280 18200
rect 240 18170 250 18190
rect 270 18170 280 18190
rect 240 18030 280 18170
rect 240 18010 250 18030
rect 270 18010 280 18030
rect 240 17870 280 18010
rect 240 17850 250 17870
rect 270 17850 280 17870
rect 240 17710 280 17850
rect 240 17690 250 17710
rect 270 17690 280 17710
rect 240 17550 280 17690
rect 240 17530 250 17550
rect 270 17530 280 17550
rect 240 17390 280 17530
rect 240 17370 250 17390
rect 270 17370 280 17390
rect 240 17230 280 17370
rect 240 17210 250 17230
rect 270 17210 280 17230
rect 240 17200 280 17210
rect 320 18190 360 18200
rect 320 18170 330 18190
rect 350 18170 360 18190
rect 320 18030 360 18170
rect 320 18010 330 18030
rect 350 18010 360 18030
rect 320 17870 360 18010
rect 320 17850 330 17870
rect 350 17850 360 17870
rect 320 17710 360 17850
rect 320 17690 330 17710
rect 350 17690 360 17710
rect 320 17550 360 17690
rect 320 17530 330 17550
rect 350 17530 360 17550
rect 320 17390 360 17530
rect 320 17370 330 17390
rect 350 17370 360 17390
rect 320 17230 360 17370
rect 320 17210 330 17230
rect 350 17210 360 17230
rect 320 17200 360 17210
rect 400 18190 440 18200
rect 400 18170 410 18190
rect 430 18170 440 18190
rect 400 18030 440 18170
rect 400 18010 410 18030
rect 430 18010 440 18030
rect 400 17870 440 18010
rect 400 17850 410 17870
rect 430 17850 440 17870
rect 400 17710 440 17850
rect 400 17690 410 17710
rect 430 17690 440 17710
rect 400 17550 440 17690
rect 400 17530 410 17550
rect 430 17530 440 17550
rect 400 17390 440 17530
rect 400 17370 410 17390
rect 430 17370 440 17390
rect 400 17230 440 17370
rect 400 17210 410 17230
rect 430 17210 440 17230
rect 400 17200 440 17210
rect 480 18190 520 18200
rect 480 18170 490 18190
rect 510 18170 520 18190
rect 480 18030 520 18170
rect 480 18010 490 18030
rect 510 18010 520 18030
rect 480 17870 520 18010
rect 480 17850 490 17870
rect 510 17850 520 17870
rect 480 17710 520 17850
rect 480 17690 490 17710
rect 510 17690 520 17710
rect 480 17550 520 17690
rect 480 17530 490 17550
rect 510 17530 520 17550
rect 480 17390 520 17530
rect 480 17370 490 17390
rect 510 17370 520 17390
rect 480 17230 520 17370
rect 480 17210 490 17230
rect 510 17210 520 17230
rect 480 17200 520 17210
rect 560 18190 600 18200
rect 560 18170 570 18190
rect 590 18170 600 18190
rect 560 18030 600 18170
rect 560 18010 570 18030
rect 590 18010 600 18030
rect 560 17870 600 18010
rect 560 17850 570 17870
rect 590 17850 600 17870
rect 560 17710 600 17850
rect 560 17690 570 17710
rect 590 17690 600 17710
rect 560 17550 600 17690
rect 560 17530 570 17550
rect 590 17530 600 17550
rect 560 17390 600 17530
rect 560 17370 570 17390
rect 590 17370 600 17390
rect 560 17230 600 17370
rect 560 17210 570 17230
rect 590 17210 600 17230
rect 560 17200 600 17210
rect 640 18190 680 18200
rect 640 18170 650 18190
rect 670 18170 680 18190
rect 640 18030 680 18170
rect 640 18010 650 18030
rect 670 18010 680 18030
rect 640 17870 680 18010
rect 640 17850 650 17870
rect 670 17850 680 17870
rect 640 17710 680 17850
rect 640 17690 650 17710
rect 670 17690 680 17710
rect 640 17550 680 17690
rect 640 17530 650 17550
rect 670 17530 680 17550
rect 640 17390 680 17530
rect 640 17370 650 17390
rect 670 17370 680 17390
rect 640 17230 680 17370
rect 640 17210 650 17230
rect 670 17210 680 17230
rect 640 17200 680 17210
rect 720 18190 760 18200
rect 720 18170 730 18190
rect 750 18170 760 18190
rect 720 18030 760 18170
rect 720 18010 730 18030
rect 750 18010 760 18030
rect 720 17870 760 18010
rect 720 17850 730 17870
rect 750 17850 760 17870
rect 720 17710 760 17850
rect 720 17690 730 17710
rect 750 17690 760 17710
rect 720 17550 760 17690
rect 720 17530 730 17550
rect 750 17530 760 17550
rect 720 17390 760 17530
rect 720 17370 730 17390
rect 750 17370 760 17390
rect 720 17230 760 17370
rect 720 17210 730 17230
rect 750 17210 760 17230
rect 720 17200 760 17210
rect 800 18190 840 18200
rect 800 18170 810 18190
rect 830 18170 840 18190
rect 800 18030 840 18170
rect 800 18010 810 18030
rect 830 18010 840 18030
rect 800 17870 840 18010
rect 800 17850 810 17870
rect 830 17850 840 17870
rect 800 17710 840 17850
rect 800 17690 810 17710
rect 830 17690 840 17710
rect 800 17550 840 17690
rect 800 17530 810 17550
rect 830 17530 840 17550
rect 800 17390 840 17530
rect 800 17370 810 17390
rect 830 17370 840 17390
rect 800 17230 840 17370
rect 800 17210 810 17230
rect 830 17210 840 17230
rect 800 17200 840 17210
rect 880 18190 920 18200
rect 880 18170 890 18190
rect 910 18170 920 18190
rect 880 18030 920 18170
rect 880 18010 890 18030
rect 910 18010 920 18030
rect 880 17870 920 18010
rect 880 17850 890 17870
rect 910 17850 920 17870
rect 880 17710 920 17850
rect 880 17690 890 17710
rect 910 17690 920 17710
rect 880 17550 920 17690
rect 880 17530 890 17550
rect 910 17530 920 17550
rect 880 17390 920 17530
rect 880 17370 890 17390
rect 910 17370 920 17390
rect 880 17230 920 17370
rect 880 17210 890 17230
rect 910 17210 920 17230
rect 880 17200 920 17210
rect 960 18190 1000 18200
rect 960 18170 970 18190
rect 990 18170 1000 18190
rect 960 18030 1000 18170
rect 960 18010 970 18030
rect 990 18010 1000 18030
rect 960 17870 1000 18010
rect 960 17850 970 17870
rect 990 17850 1000 17870
rect 960 17710 1000 17850
rect 960 17690 970 17710
rect 990 17690 1000 17710
rect 960 17550 1000 17690
rect 960 17530 970 17550
rect 990 17530 1000 17550
rect 960 17390 1000 17530
rect 960 17370 970 17390
rect 990 17370 1000 17390
rect 960 17230 1000 17370
rect 960 17210 970 17230
rect 990 17210 1000 17230
rect 960 17200 1000 17210
rect 1040 18190 1080 18200
rect 1040 18170 1050 18190
rect 1070 18170 1080 18190
rect 1040 18030 1080 18170
rect 1040 18010 1050 18030
rect 1070 18010 1080 18030
rect 1040 17870 1080 18010
rect 1040 17850 1050 17870
rect 1070 17850 1080 17870
rect 1040 17710 1080 17850
rect 1040 17690 1050 17710
rect 1070 17690 1080 17710
rect 1040 17550 1080 17690
rect 1040 17530 1050 17550
rect 1070 17530 1080 17550
rect 1040 17390 1080 17530
rect 1040 17370 1050 17390
rect 1070 17370 1080 17390
rect 1040 17230 1080 17370
rect 1040 17210 1050 17230
rect 1070 17210 1080 17230
rect 1040 17200 1080 17210
rect 1120 18190 1160 18200
rect 1120 18170 1130 18190
rect 1150 18170 1160 18190
rect 1120 18030 1160 18170
rect 1120 18010 1130 18030
rect 1150 18010 1160 18030
rect 1120 17870 1160 18010
rect 1120 17850 1130 17870
rect 1150 17850 1160 17870
rect 1120 17710 1160 17850
rect 1120 17690 1130 17710
rect 1150 17690 1160 17710
rect 1120 17550 1160 17690
rect 1120 17530 1130 17550
rect 1150 17530 1160 17550
rect 1120 17390 1160 17530
rect 1120 17370 1130 17390
rect 1150 17370 1160 17390
rect 1120 17230 1160 17370
rect 1120 17210 1130 17230
rect 1150 17210 1160 17230
rect 1120 17200 1160 17210
rect 1200 18190 1240 18200
rect 1200 18170 1210 18190
rect 1230 18170 1240 18190
rect 1200 18030 1240 18170
rect 1200 18010 1210 18030
rect 1230 18010 1240 18030
rect 1200 17870 1240 18010
rect 1200 17850 1210 17870
rect 1230 17850 1240 17870
rect 1200 17710 1240 17850
rect 1200 17690 1210 17710
rect 1230 17690 1240 17710
rect 1200 17550 1240 17690
rect 1200 17530 1210 17550
rect 1230 17530 1240 17550
rect 1200 17390 1240 17530
rect 1200 17370 1210 17390
rect 1230 17370 1240 17390
rect 1200 17230 1240 17370
rect 1200 17210 1210 17230
rect 1230 17210 1240 17230
rect 1200 17200 1240 17210
rect 1280 18190 1320 18200
rect 1280 18170 1290 18190
rect 1310 18170 1320 18190
rect 1280 18030 1320 18170
rect 1280 18010 1290 18030
rect 1310 18010 1320 18030
rect 1280 17870 1320 18010
rect 1280 17850 1290 17870
rect 1310 17850 1320 17870
rect 1280 17710 1320 17850
rect 1280 17690 1290 17710
rect 1310 17690 1320 17710
rect 1280 17550 1320 17690
rect 1280 17530 1290 17550
rect 1310 17530 1320 17550
rect 1280 17390 1320 17530
rect 1280 17370 1290 17390
rect 1310 17370 1320 17390
rect 1280 17230 1320 17370
rect 1280 17210 1290 17230
rect 1310 17210 1320 17230
rect 1280 17200 1320 17210
rect 1360 18190 1400 18200
rect 1360 18170 1370 18190
rect 1390 18170 1400 18190
rect 1360 18030 1400 18170
rect 1360 18010 1370 18030
rect 1390 18010 1400 18030
rect 1360 17870 1400 18010
rect 1360 17850 1370 17870
rect 1390 17850 1400 17870
rect 1360 17710 1400 17850
rect 1360 17690 1370 17710
rect 1390 17690 1400 17710
rect 1360 17550 1400 17690
rect 1360 17530 1370 17550
rect 1390 17530 1400 17550
rect 1360 17390 1400 17530
rect 1360 17370 1370 17390
rect 1390 17370 1400 17390
rect 1360 17230 1400 17370
rect 1360 17210 1370 17230
rect 1390 17210 1400 17230
rect 1360 17200 1400 17210
rect 1440 18190 1480 18200
rect 1440 18170 1450 18190
rect 1470 18170 1480 18190
rect 1440 18030 1480 18170
rect 1440 18010 1450 18030
rect 1470 18010 1480 18030
rect 1440 17870 1480 18010
rect 1440 17850 1450 17870
rect 1470 17850 1480 17870
rect 1440 17710 1480 17850
rect 1440 17690 1450 17710
rect 1470 17690 1480 17710
rect 1440 17550 1480 17690
rect 1440 17530 1450 17550
rect 1470 17530 1480 17550
rect 1440 17390 1480 17530
rect 1440 17370 1450 17390
rect 1470 17370 1480 17390
rect 1440 17230 1480 17370
rect 1440 17210 1450 17230
rect 1470 17210 1480 17230
rect 1440 17200 1480 17210
rect 1520 18190 1560 18200
rect 1520 18170 1530 18190
rect 1550 18170 1560 18190
rect 1520 18030 1560 18170
rect 1520 18010 1530 18030
rect 1550 18010 1560 18030
rect 1520 17870 1560 18010
rect 1520 17850 1530 17870
rect 1550 17850 1560 17870
rect 1520 17710 1560 17850
rect 1520 17690 1530 17710
rect 1550 17690 1560 17710
rect 1520 17550 1560 17690
rect 1520 17530 1530 17550
rect 1550 17530 1560 17550
rect 1520 17390 1560 17530
rect 1520 17370 1530 17390
rect 1550 17370 1560 17390
rect 1520 17230 1560 17370
rect 1520 17210 1530 17230
rect 1550 17210 1560 17230
rect 1520 17200 1560 17210
rect 1600 18190 1640 18200
rect 1600 18170 1610 18190
rect 1630 18170 1640 18190
rect 1600 18030 1640 18170
rect 1600 18010 1610 18030
rect 1630 18010 1640 18030
rect 1600 17870 1640 18010
rect 1600 17850 1610 17870
rect 1630 17850 1640 17870
rect 1600 17710 1640 17850
rect 1600 17690 1610 17710
rect 1630 17690 1640 17710
rect 1600 17550 1640 17690
rect 1600 17530 1610 17550
rect 1630 17530 1640 17550
rect 1600 17390 1640 17530
rect 1600 17370 1610 17390
rect 1630 17370 1640 17390
rect 1600 17230 1640 17370
rect 1600 17210 1610 17230
rect 1630 17210 1640 17230
rect 1600 17200 1640 17210
rect 1680 18190 1720 18200
rect 1680 18170 1690 18190
rect 1710 18170 1720 18190
rect 1680 18030 1720 18170
rect 1680 18010 1690 18030
rect 1710 18010 1720 18030
rect 1680 17870 1720 18010
rect 1680 17850 1690 17870
rect 1710 17850 1720 17870
rect 1680 17710 1720 17850
rect 1680 17690 1690 17710
rect 1710 17690 1720 17710
rect 1680 17550 1720 17690
rect 1680 17530 1690 17550
rect 1710 17530 1720 17550
rect 1680 17390 1720 17530
rect 1680 17370 1690 17390
rect 1710 17370 1720 17390
rect 1680 17230 1720 17370
rect 1680 17210 1690 17230
rect 1710 17210 1720 17230
rect 1680 17200 1720 17210
rect 1760 18190 1800 18200
rect 1760 18170 1770 18190
rect 1790 18170 1800 18190
rect 1760 18030 1800 18170
rect 1760 18010 1770 18030
rect 1790 18010 1800 18030
rect 1760 17870 1800 18010
rect 1760 17850 1770 17870
rect 1790 17850 1800 17870
rect 1760 17710 1800 17850
rect 1760 17690 1770 17710
rect 1790 17690 1800 17710
rect 1760 17550 1800 17690
rect 1760 17530 1770 17550
rect 1790 17530 1800 17550
rect 1760 17390 1800 17530
rect 1760 17370 1770 17390
rect 1790 17370 1800 17390
rect 1760 17230 1800 17370
rect 1760 17210 1770 17230
rect 1790 17210 1800 17230
rect 1760 17200 1800 17210
rect 1840 18190 1880 18200
rect 1840 18170 1850 18190
rect 1870 18170 1880 18190
rect 1840 18030 1880 18170
rect 1840 18010 1850 18030
rect 1870 18010 1880 18030
rect 1840 17870 1880 18010
rect 1840 17850 1850 17870
rect 1870 17850 1880 17870
rect 1840 17710 1880 17850
rect 1840 17690 1850 17710
rect 1870 17690 1880 17710
rect 1840 17550 1880 17690
rect 1840 17530 1850 17550
rect 1870 17530 1880 17550
rect 1840 17390 1880 17530
rect 1840 17370 1850 17390
rect 1870 17370 1880 17390
rect 1840 17230 1880 17370
rect 1840 17210 1850 17230
rect 1870 17210 1880 17230
rect 1840 17200 1880 17210
rect 1920 18190 1960 18200
rect 1920 18170 1930 18190
rect 1950 18170 1960 18190
rect 1920 18030 1960 18170
rect 1920 18010 1930 18030
rect 1950 18010 1960 18030
rect 1920 17870 1960 18010
rect 1920 17850 1930 17870
rect 1950 17850 1960 17870
rect 1920 17710 1960 17850
rect 1920 17690 1930 17710
rect 1950 17690 1960 17710
rect 1920 17550 1960 17690
rect 1920 17530 1930 17550
rect 1950 17530 1960 17550
rect 1920 17390 1960 17530
rect 1920 17370 1930 17390
rect 1950 17370 1960 17390
rect 1920 17230 1960 17370
rect 1920 17210 1930 17230
rect 1950 17210 1960 17230
rect 1920 17200 1960 17210
rect 2000 18190 2040 18200
rect 2000 18170 2010 18190
rect 2030 18170 2040 18190
rect 2000 18030 2040 18170
rect 2000 18010 2010 18030
rect 2030 18010 2040 18030
rect 2000 17870 2040 18010
rect 2000 17850 2010 17870
rect 2030 17850 2040 17870
rect 2000 17710 2040 17850
rect 2000 17690 2010 17710
rect 2030 17690 2040 17710
rect 2000 17550 2040 17690
rect 2000 17530 2010 17550
rect 2030 17530 2040 17550
rect 2000 17390 2040 17530
rect 2000 17370 2010 17390
rect 2030 17370 2040 17390
rect 2000 17230 2040 17370
rect 2000 17210 2010 17230
rect 2030 17210 2040 17230
rect 2000 17200 2040 17210
rect 2080 18190 2120 18200
rect 2080 18170 2090 18190
rect 2110 18170 2120 18190
rect 2080 18030 2120 18170
rect 2080 18010 2090 18030
rect 2110 18010 2120 18030
rect 2080 17870 2120 18010
rect 2080 17850 2090 17870
rect 2110 17850 2120 17870
rect 2080 17710 2120 17850
rect 2080 17690 2090 17710
rect 2110 17690 2120 17710
rect 2080 17550 2120 17690
rect 2080 17530 2090 17550
rect 2110 17530 2120 17550
rect 2080 17390 2120 17530
rect 2080 17370 2090 17390
rect 2110 17370 2120 17390
rect 2080 17230 2120 17370
rect 2080 17210 2090 17230
rect 2110 17210 2120 17230
rect 2080 17200 2120 17210
rect 2160 18190 2200 18200
rect 2160 18170 2170 18190
rect 2190 18170 2200 18190
rect 2160 18030 2200 18170
rect 2160 18010 2170 18030
rect 2190 18010 2200 18030
rect 2160 17870 2200 18010
rect 2160 17850 2170 17870
rect 2190 17850 2200 17870
rect 2160 17710 2200 17850
rect 2160 17690 2170 17710
rect 2190 17690 2200 17710
rect 2160 17550 2200 17690
rect 2160 17530 2170 17550
rect 2190 17530 2200 17550
rect 2160 17390 2200 17530
rect 2160 17370 2170 17390
rect 2190 17370 2200 17390
rect 2160 17230 2200 17370
rect 2160 17210 2170 17230
rect 2190 17210 2200 17230
rect 2160 17200 2200 17210
rect 2240 18190 2280 18200
rect 2240 18170 2250 18190
rect 2270 18170 2280 18190
rect 2240 18030 2280 18170
rect 2240 18010 2250 18030
rect 2270 18010 2280 18030
rect 2240 17870 2280 18010
rect 2240 17850 2250 17870
rect 2270 17850 2280 17870
rect 2240 17710 2280 17850
rect 2240 17690 2250 17710
rect 2270 17690 2280 17710
rect 2240 17550 2280 17690
rect 2240 17530 2250 17550
rect 2270 17530 2280 17550
rect 2240 17390 2280 17530
rect 2240 17370 2250 17390
rect 2270 17370 2280 17390
rect 2240 17230 2280 17370
rect 2240 17210 2250 17230
rect 2270 17210 2280 17230
rect 2240 17200 2280 17210
rect 2320 18190 2360 18200
rect 2320 18170 2330 18190
rect 2350 18170 2360 18190
rect 2320 18030 2360 18170
rect 2320 18010 2330 18030
rect 2350 18010 2360 18030
rect 2320 17870 2360 18010
rect 2320 17850 2330 17870
rect 2350 17850 2360 17870
rect 2320 17710 2360 17850
rect 2320 17690 2330 17710
rect 2350 17690 2360 17710
rect 2320 17550 2360 17690
rect 2320 17530 2330 17550
rect 2350 17530 2360 17550
rect 2320 17390 2360 17530
rect 2320 17370 2330 17390
rect 2350 17370 2360 17390
rect 2320 17230 2360 17370
rect 2320 17210 2330 17230
rect 2350 17210 2360 17230
rect 2320 17200 2360 17210
rect 2400 18190 2440 18200
rect 2400 18170 2410 18190
rect 2430 18170 2440 18190
rect 2400 18030 2440 18170
rect 2400 18010 2410 18030
rect 2430 18010 2440 18030
rect 2400 17870 2440 18010
rect 2400 17850 2410 17870
rect 2430 17850 2440 17870
rect 2400 17710 2440 17850
rect 2400 17690 2410 17710
rect 2430 17690 2440 17710
rect 2400 17550 2440 17690
rect 2400 17530 2410 17550
rect 2430 17530 2440 17550
rect 2400 17390 2440 17530
rect 2400 17370 2410 17390
rect 2430 17370 2440 17390
rect 2400 17230 2440 17370
rect 2400 17210 2410 17230
rect 2430 17210 2440 17230
rect 2400 17200 2440 17210
rect 2480 18190 2520 18200
rect 2480 18170 2490 18190
rect 2510 18170 2520 18190
rect 2480 18030 2520 18170
rect 2480 18010 2490 18030
rect 2510 18010 2520 18030
rect 2480 17870 2520 18010
rect 2480 17850 2490 17870
rect 2510 17850 2520 17870
rect 2480 17710 2520 17850
rect 2480 17690 2490 17710
rect 2510 17690 2520 17710
rect 2480 17550 2520 17690
rect 2480 17530 2490 17550
rect 2510 17530 2520 17550
rect 2480 17390 2520 17530
rect 2480 17370 2490 17390
rect 2510 17370 2520 17390
rect 2480 17230 2520 17370
rect 2480 17210 2490 17230
rect 2510 17210 2520 17230
rect 2480 17200 2520 17210
rect 2560 18190 2600 18200
rect 2560 18170 2570 18190
rect 2590 18170 2600 18190
rect 2560 18030 2600 18170
rect 2560 18010 2570 18030
rect 2590 18010 2600 18030
rect 2560 17870 2600 18010
rect 2560 17850 2570 17870
rect 2590 17850 2600 17870
rect 2560 17710 2600 17850
rect 2560 17690 2570 17710
rect 2590 17690 2600 17710
rect 2560 17550 2600 17690
rect 2560 17530 2570 17550
rect 2590 17530 2600 17550
rect 2560 17390 2600 17530
rect 2560 17370 2570 17390
rect 2590 17370 2600 17390
rect 2560 17230 2600 17370
rect 2560 17210 2570 17230
rect 2590 17210 2600 17230
rect 2560 17200 2600 17210
rect 2640 18190 2680 18200
rect 2640 18170 2650 18190
rect 2670 18170 2680 18190
rect 2640 18030 2680 18170
rect 2640 18010 2650 18030
rect 2670 18010 2680 18030
rect 2640 17870 2680 18010
rect 2640 17850 2650 17870
rect 2670 17850 2680 17870
rect 2640 17710 2680 17850
rect 2640 17690 2650 17710
rect 2670 17690 2680 17710
rect 2640 17550 2680 17690
rect 2640 17530 2650 17550
rect 2670 17530 2680 17550
rect 2640 17390 2680 17530
rect 2640 17370 2650 17390
rect 2670 17370 2680 17390
rect 2640 17230 2680 17370
rect 2640 17210 2650 17230
rect 2670 17210 2680 17230
rect 2640 17200 2680 17210
rect 2720 18190 2760 18200
rect 2720 18170 2730 18190
rect 2750 18170 2760 18190
rect 2720 18030 2760 18170
rect 2720 18010 2730 18030
rect 2750 18010 2760 18030
rect 2720 17870 2760 18010
rect 2720 17850 2730 17870
rect 2750 17850 2760 17870
rect 2720 17710 2760 17850
rect 2720 17690 2730 17710
rect 2750 17690 2760 17710
rect 2720 17550 2760 17690
rect 2720 17530 2730 17550
rect 2750 17530 2760 17550
rect 2720 17390 2760 17530
rect 2720 17370 2730 17390
rect 2750 17370 2760 17390
rect 2720 17230 2760 17370
rect 2720 17210 2730 17230
rect 2750 17210 2760 17230
rect 2720 17200 2760 17210
rect 2800 18190 2840 18200
rect 2800 18170 2810 18190
rect 2830 18170 2840 18190
rect 2800 18030 2840 18170
rect 2800 18010 2810 18030
rect 2830 18010 2840 18030
rect 2800 17870 2840 18010
rect 2800 17850 2810 17870
rect 2830 17850 2840 17870
rect 2800 17710 2840 17850
rect 2800 17690 2810 17710
rect 2830 17690 2840 17710
rect 2800 17550 2840 17690
rect 2800 17530 2810 17550
rect 2830 17530 2840 17550
rect 2800 17390 2840 17530
rect 2800 17370 2810 17390
rect 2830 17370 2840 17390
rect 2800 17230 2840 17370
rect 2800 17210 2810 17230
rect 2830 17210 2840 17230
rect 2800 17200 2840 17210
rect 2880 18190 2920 18200
rect 2880 18170 2890 18190
rect 2910 18170 2920 18190
rect 2880 18030 2920 18170
rect 2880 18010 2890 18030
rect 2910 18010 2920 18030
rect 2880 17870 2920 18010
rect 2880 17850 2890 17870
rect 2910 17850 2920 17870
rect 2880 17710 2920 17850
rect 2880 17690 2890 17710
rect 2910 17690 2920 17710
rect 2880 17550 2920 17690
rect 2880 17530 2890 17550
rect 2910 17530 2920 17550
rect 2880 17390 2920 17530
rect 2880 17370 2890 17390
rect 2910 17370 2920 17390
rect 2880 17230 2920 17370
rect 2880 17210 2890 17230
rect 2910 17210 2920 17230
rect 2880 17200 2920 17210
rect 2960 18190 3000 18200
rect 2960 18170 2970 18190
rect 2990 18170 3000 18190
rect 2960 18030 3000 18170
rect 2960 18010 2970 18030
rect 2990 18010 3000 18030
rect 2960 17870 3000 18010
rect 2960 17850 2970 17870
rect 2990 17850 3000 17870
rect 2960 17710 3000 17850
rect 2960 17690 2970 17710
rect 2990 17690 3000 17710
rect 2960 17550 3000 17690
rect 2960 17530 2970 17550
rect 2990 17530 3000 17550
rect 2960 17390 3000 17530
rect 2960 17370 2970 17390
rect 2990 17370 3000 17390
rect 2960 17230 3000 17370
rect 2960 17210 2970 17230
rect 2990 17210 3000 17230
rect 2960 17200 3000 17210
rect 3040 18190 3080 18200
rect 3040 18170 3050 18190
rect 3070 18170 3080 18190
rect 3040 18030 3080 18170
rect 3040 18010 3050 18030
rect 3070 18010 3080 18030
rect 3040 17870 3080 18010
rect 3040 17850 3050 17870
rect 3070 17850 3080 17870
rect 3040 17710 3080 17850
rect 3040 17690 3050 17710
rect 3070 17690 3080 17710
rect 3040 17550 3080 17690
rect 3040 17530 3050 17550
rect 3070 17530 3080 17550
rect 3040 17390 3080 17530
rect 3040 17370 3050 17390
rect 3070 17370 3080 17390
rect 3040 17230 3080 17370
rect 3040 17210 3050 17230
rect 3070 17210 3080 17230
rect 3040 17200 3080 17210
rect 3120 18190 3160 18200
rect 3120 18170 3130 18190
rect 3150 18170 3160 18190
rect 3120 18030 3160 18170
rect 3120 18010 3130 18030
rect 3150 18010 3160 18030
rect 3120 17870 3160 18010
rect 3120 17850 3130 17870
rect 3150 17850 3160 17870
rect 3120 17710 3160 17850
rect 3120 17690 3130 17710
rect 3150 17690 3160 17710
rect 3120 17550 3160 17690
rect 3120 17530 3130 17550
rect 3150 17530 3160 17550
rect 3120 17390 3160 17530
rect 3120 17370 3130 17390
rect 3150 17370 3160 17390
rect 3120 17230 3160 17370
rect 3120 17210 3130 17230
rect 3150 17210 3160 17230
rect 3120 17200 3160 17210
rect 3200 18190 3240 18200
rect 3200 18170 3210 18190
rect 3230 18170 3240 18190
rect 3200 18030 3240 18170
rect 3200 18010 3210 18030
rect 3230 18010 3240 18030
rect 3200 17870 3240 18010
rect 3200 17850 3210 17870
rect 3230 17850 3240 17870
rect 3200 17710 3240 17850
rect 3200 17690 3210 17710
rect 3230 17690 3240 17710
rect 3200 17550 3240 17690
rect 3200 17530 3210 17550
rect 3230 17530 3240 17550
rect 3200 17390 3240 17530
rect 3200 17370 3210 17390
rect 3230 17370 3240 17390
rect 3200 17230 3240 17370
rect 3200 17210 3210 17230
rect 3230 17210 3240 17230
rect 3200 17200 3240 17210
rect 3280 18190 3320 18200
rect 3280 18170 3290 18190
rect 3310 18170 3320 18190
rect 3280 18030 3320 18170
rect 3280 18010 3290 18030
rect 3310 18010 3320 18030
rect 3280 17870 3320 18010
rect 3280 17850 3290 17870
rect 3310 17850 3320 17870
rect 3280 17710 3320 17850
rect 3280 17690 3290 17710
rect 3310 17690 3320 17710
rect 3280 17550 3320 17690
rect 3280 17530 3290 17550
rect 3310 17530 3320 17550
rect 3280 17390 3320 17530
rect 3280 17370 3290 17390
rect 3310 17370 3320 17390
rect 3280 17230 3320 17370
rect 3280 17210 3290 17230
rect 3310 17210 3320 17230
rect 3280 17200 3320 17210
rect 3360 18190 3400 18200
rect 3360 18170 3370 18190
rect 3390 18170 3400 18190
rect 3360 18030 3400 18170
rect 3360 18010 3370 18030
rect 3390 18010 3400 18030
rect 3360 17870 3400 18010
rect 3360 17850 3370 17870
rect 3390 17850 3400 17870
rect 3360 17710 3400 17850
rect 3360 17690 3370 17710
rect 3390 17690 3400 17710
rect 3360 17550 3400 17690
rect 3360 17530 3370 17550
rect 3390 17530 3400 17550
rect 3360 17390 3400 17530
rect 3360 17370 3370 17390
rect 3390 17370 3400 17390
rect 3360 17230 3400 17370
rect 3360 17210 3370 17230
rect 3390 17210 3400 17230
rect 3360 17200 3400 17210
rect 3440 18190 3480 18200
rect 3440 18170 3450 18190
rect 3470 18170 3480 18190
rect 3440 18030 3480 18170
rect 3440 18010 3450 18030
rect 3470 18010 3480 18030
rect 3440 17870 3480 18010
rect 3440 17850 3450 17870
rect 3470 17850 3480 17870
rect 3440 17710 3480 17850
rect 3440 17690 3450 17710
rect 3470 17690 3480 17710
rect 3440 17550 3480 17690
rect 3440 17530 3450 17550
rect 3470 17530 3480 17550
rect 3440 17390 3480 17530
rect 3440 17370 3450 17390
rect 3470 17370 3480 17390
rect 3440 17230 3480 17370
rect 3440 17210 3450 17230
rect 3470 17210 3480 17230
rect 3440 17200 3480 17210
rect 3520 18190 3560 18200
rect 3520 18170 3530 18190
rect 3550 18170 3560 18190
rect 3520 18030 3560 18170
rect 3520 18010 3530 18030
rect 3550 18010 3560 18030
rect 3520 17870 3560 18010
rect 3520 17850 3530 17870
rect 3550 17850 3560 17870
rect 3520 17710 3560 17850
rect 3520 17690 3530 17710
rect 3550 17690 3560 17710
rect 3520 17550 3560 17690
rect 3520 17530 3530 17550
rect 3550 17530 3560 17550
rect 3520 17390 3560 17530
rect 3520 17370 3530 17390
rect 3550 17370 3560 17390
rect 3520 17230 3560 17370
rect 3520 17210 3530 17230
rect 3550 17210 3560 17230
rect 3520 17200 3560 17210
rect 3600 18190 3640 18200
rect 3600 18170 3610 18190
rect 3630 18170 3640 18190
rect 3600 18030 3640 18170
rect 3600 18010 3610 18030
rect 3630 18010 3640 18030
rect 3600 17870 3640 18010
rect 3600 17850 3610 17870
rect 3630 17850 3640 17870
rect 3600 17710 3640 17850
rect 3600 17690 3610 17710
rect 3630 17690 3640 17710
rect 3600 17550 3640 17690
rect 3600 17530 3610 17550
rect 3630 17530 3640 17550
rect 3600 17390 3640 17530
rect 3600 17370 3610 17390
rect 3630 17370 3640 17390
rect 3600 17230 3640 17370
rect 3600 17210 3610 17230
rect 3630 17210 3640 17230
rect 3600 17200 3640 17210
rect 3680 18190 3720 18200
rect 3680 18170 3690 18190
rect 3710 18170 3720 18190
rect 3680 18030 3720 18170
rect 3680 18010 3690 18030
rect 3710 18010 3720 18030
rect 3680 17870 3720 18010
rect 3680 17850 3690 17870
rect 3710 17850 3720 17870
rect 3680 17710 3720 17850
rect 3680 17690 3690 17710
rect 3710 17690 3720 17710
rect 3680 17550 3720 17690
rect 3680 17530 3690 17550
rect 3710 17530 3720 17550
rect 3680 17390 3720 17530
rect 3680 17370 3690 17390
rect 3710 17370 3720 17390
rect 3680 17230 3720 17370
rect 3680 17210 3690 17230
rect 3710 17210 3720 17230
rect 3680 17200 3720 17210
rect 3760 18190 3800 18200
rect 3760 18170 3770 18190
rect 3790 18170 3800 18190
rect 3760 18030 3800 18170
rect 3760 18010 3770 18030
rect 3790 18010 3800 18030
rect 3760 17870 3800 18010
rect 3760 17850 3770 17870
rect 3790 17850 3800 17870
rect 3760 17710 3800 17850
rect 3760 17690 3770 17710
rect 3790 17690 3800 17710
rect 3760 17550 3800 17690
rect 3760 17530 3770 17550
rect 3790 17530 3800 17550
rect 3760 17390 3800 17530
rect 3760 17370 3770 17390
rect 3790 17370 3800 17390
rect 3760 17230 3800 17370
rect 3760 17210 3770 17230
rect 3790 17210 3800 17230
rect 3760 17200 3800 17210
rect 3840 18190 3880 18200
rect 3840 18170 3850 18190
rect 3870 18170 3880 18190
rect 3840 18030 3880 18170
rect 3840 18010 3850 18030
rect 3870 18010 3880 18030
rect 3840 17870 3880 18010
rect 3840 17850 3850 17870
rect 3870 17850 3880 17870
rect 3840 17710 3880 17850
rect 3840 17690 3850 17710
rect 3870 17690 3880 17710
rect 3840 17550 3880 17690
rect 3840 17530 3850 17550
rect 3870 17530 3880 17550
rect 3840 17390 3880 17530
rect 3840 17370 3850 17390
rect 3870 17370 3880 17390
rect 3840 17230 3880 17370
rect 3840 17210 3850 17230
rect 3870 17210 3880 17230
rect 3840 17200 3880 17210
rect 3920 18190 3960 18200
rect 3920 18170 3930 18190
rect 3950 18170 3960 18190
rect 3920 18030 3960 18170
rect 3920 18010 3930 18030
rect 3950 18010 3960 18030
rect 3920 17870 3960 18010
rect 3920 17850 3930 17870
rect 3950 17850 3960 17870
rect 3920 17710 3960 17850
rect 3920 17690 3930 17710
rect 3950 17690 3960 17710
rect 3920 17550 3960 17690
rect 3920 17530 3930 17550
rect 3950 17530 3960 17550
rect 3920 17390 3960 17530
rect 3920 17370 3930 17390
rect 3950 17370 3960 17390
rect 3920 17230 3960 17370
rect 3920 17210 3930 17230
rect 3950 17210 3960 17230
rect 3920 17200 3960 17210
rect 4000 18190 4040 18200
rect 4000 18170 4010 18190
rect 4030 18170 4040 18190
rect 4000 18030 4040 18170
rect 4000 18010 4010 18030
rect 4030 18010 4040 18030
rect 4000 17870 4040 18010
rect 4000 17850 4010 17870
rect 4030 17850 4040 17870
rect 4000 17710 4040 17850
rect 4000 17690 4010 17710
rect 4030 17690 4040 17710
rect 4000 17550 4040 17690
rect 4000 17530 4010 17550
rect 4030 17530 4040 17550
rect 4000 17390 4040 17530
rect 4000 17370 4010 17390
rect 4030 17370 4040 17390
rect 4000 17230 4040 17370
rect 4000 17210 4010 17230
rect 4030 17210 4040 17230
rect 4000 17200 4040 17210
rect 4080 18190 4120 18200
rect 4080 18170 4090 18190
rect 4110 18170 4120 18190
rect 4080 18030 4120 18170
rect 4080 18010 4090 18030
rect 4110 18010 4120 18030
rect 4080 17870 4120 18010
rect 4080 17850 4090 17870
rect 4110 17850 4120 17870
rect 4080 17710 4120 17850
rect 4080 17690 4090 17710
rect 4110 17690 4120 17710
rect 4080 17550 4120 17690
rect 4080 17530 4090 17550
rect 4110 17530 4120 17550
rect 4080 17390 4120 17530
rect 4080 17370 4090 17390
rect 4110 17370 4120 17390
rect 4080 17230 4120 17370
rect 4080 17210 4090 17230
rect 4110 17210 4120 17230
rect 4080 17200 4120 17210
rect 4160 18190 4200 18200
rect 4160 18170 4170 18190
rect 4190 18170 4200 18190
rect 4160 18030 4200 18170
rect 4160 18010 4170 18030
rect 4190 18010 4200 18030
rect 4160 17870 4200 18010
rect 4160 17850 4170 17870
rect 4190 17850 4200 17870
rect 4160 17710 4200 17850
rect 4160 17690 4170 17710
rect 4190 17690 4200 17710
rect 4160 17550 4200 17690
rect 4160 17530 4170 17550
rect 4190 17530 4200 17550
rect 4160 17390 4200 17530
rect 4160 17370 4170 17390
rect 4190 17370 4200 17390
rect 4160 17230 4200 17370
rect 4160 17210 4170 17230
rect 4190 17210 4200 17230
rect 4160 17200 4200 17210
rect 4240 17200 4280 18200
rect 4320 17200 4360 18200
rect 4400 17200 4440 18200
rect 4480 17200 4520 18200
rect 4560 17200 4600 18200
rect 4640 17200 4680 18200
rect 4720 17200 4760 18200
rect 4800 17200 4840 18200
rect 4880 17200 4920 18200
rect 4960 17200 5000 18200
rect 5040 17200 5080 18200
rect 5120 17200 5160 18200
rect 5200 17200 5240 18200
rect 5280 17200 5320 18200
rect 5360 17200 5400 18200
rect 5440 17200 5480 18200
rect 5520 17200 5560 18200
rect 5600 17200 5640 18200
rect 5680 17200 5720 18200
rect 5760 17200 5800 18200
rect 5840 17200 5880 18200
rect 5920 17200 5960 18200
rect 6000 17200 6040 18200
rect 6080 17200 6120 18200
rect 6160 17200 6200 18200
rect 6240 18190 6280 18200
rect 6240 18170 6250 18190
rect 6270 18170 6280 18190
rect 6240 18030 6280 18170
rect 6240 18010 6250 18030
rect 6270 18010 6280 18030
rect 6240 17870 6280 18010
rect 6240 17850 6250 17870
rect 6270 17850 6280 17870
rect 6240 17710 6280 17850
rect 6240 17690 6250 17710
rect 6270 17690 6280 17710
rect 6240 17550 6280 17690
rect 6240 17530 6250 17550
rect 6270 17530 6280 17550
rect 6240 17390 6280 17530
rect 6240 17370 6250 17390
rect 6270 17370 6280 17390
rect 6240 17230 6280 17370
rect 6240 17210 6250 17230
rect 6270 17210 6280 17230
rect 6240 17200 6280 17210
rect 6320 18190 6360 18200
rect 6320 18170 6330 18190
rect 6350 18170 6360 18190
rect 6320 18030 6360 18170
rect 6320 18010 6330 18030
rect 6350 18010 6360 18030
rect 6320 17870 6360 18010
rect 6320 17850 6330 17870
rect 6350 17850 6360 17870
rect 6320 17710 6360 17850
rect 6320 17690 6330 17710
rect 6350 17690 6360 17710
rect 6320 17550 6360 17690
rect 6320 17530 6330 17550
rect 6350 17530 6360 17550
rect 6320 17390 6360 17530
rect 6320 17370 6330 17390
rect 6350 17370 6360 17390
rect 6320 17230 6360 17370
rect 6320 17210 6330 17230
rect 6350 17210 6360 17230
rect 6320 17200 6360 17210
rect 6400 18190 6440 18200
rect 6400 18170 6410 18190
rect 6430 18170 6440 18190
rect 6400 18030 6440 18170
rect 6400 18010 6410 18030
rect 6430 18010 6440 18030
rect 6400 17870 6440 18010
rect 6400 17850 6410 17870
rect 6430 17850 6440 17870
rect 6400 17710 6440 17850
rect 6400 17690 6410 17710
rect 6430 17690 6440 17710
rect 6400 17550 6440 17690
rect 6400 17530 6410 17550
rect 6430 17530 6440 17550
rect 6400 17390 6440 17530
rect 6400 17370 6410 17390
rect 6430 17370 6440 17390
rect 6400 17230 6440 17370
rect 6400 17210 6410 17230
rect 6430 17210 6440 17230
rect 6400 17200 6440 17210
rect 6480 18190 6520 18200
rect 6480 18170 6490 18190
rect 6510 18170 6520 18190
rect 6480 18030 6520 18170
rect 6480 18010 6490 18030
rect 6510 18010 6520 18030
rect 6480 17870 6520 18010
rect 6480 17850 6490 17870
rect 6510 17850 6520 17870
rect 6480 17710 6520 17850
rect 6480 17690 6490 17710
rect 6510 17690 6520 17710
rect 6480 17550 6520 17690
rect 6480 17530 6490 17550
rect 6510 17530 6520 17550
rect 6480 17390 6520 17530
rect 6480 17370 6490 17390
rect 6510 17370 6520 17390
rect 6480 17230 6520 17370
rect 6480 17210 6490 17230
rect 6510 17210 6520 17230
rect 6480 17200 6520 17210
rect 6560 18190 6600 18200
rect 6560 18170 6570 18190
rect 6590 18170 6600 18190
rect 6560 18030 6600 18170
rect 6560 18010 6570 18030
rect 6590 18010 6600 18030
rect 6560 17870 6600 18010
rect 6560 17850 6570 17870
rect 6590 17850 6600 17870
rect 6560 17710 6600 17850
rect 6560 17690 6570 17710
rect 6590 17690 6600 17710
rect 6560 17550 6600 17690
rect 6560 17530 6570 17550
rect 6590 17530 6600 17550
rect 6560 17390 6600 17530
rect 6560 17370 6570 17390
rect 6590 17370 6600 17390
rect 6560 17230 6600 17370
rect 6560 17210 6570 17230
rect 6590 17210 6600 17230
rect 6560 17200 6600 17210
rect 6640 18190 6680 18200
rect 6640 18170 6650 18190
rect 6670 18170 6680 18190
rect 6640 18030 6680 18170
rect 6640 18010 6650 18030
rect 6670 18010 6680 18030
rect 6640 17870 6680 18010
rect 6640 17850 6650 17870
rect 6670 17850 6680 17870
rect 6640 17710 6680 17850
rect 6640 17690 6650 17710
rect 6670 17690 6680 17710
rect 6640 17550 6680 17690
rect 6640 17530 6650 17550
rect 6670 17530 6680 17550
rect 6640 17390 6680 17530
rect 6640 17370 6650 17390
rect 6670 17370 6680 17390
rect 6640 17230 6680 17370
rect 6640 17210 6650 17230
rect 6670 17210 6680 17230
rect 6640 17200 6680 17210
rect 6720 18190 6760 18200
rect 6720 18170 6730 18190
rect 6750 18170 6760 18190
rect 6720 18030 6760 18170
rect 6720 18010 6730 18030
rect 6750 18010 6760 18030
rect 6720 17870 6760 18010
rect 6720 17850 6730 17870
rect 6750 17850 6760 17870
rect 6720 17710 6760 17850
rect 6720 17690 6730 17710
rect 6750 17690 6760 17710
rect 6720 17550 6760 17690
rect 6720 17530 6730 17550
rect 6750 17530 6760 17550
rect 6720 17390 6760 17530
rect 6720 17370 6730 17390
rect 6750 17370 6760 17390
rect 6720 17230 6760 17370
rect 6720 17210 6730 17230
rect 6750 17210 6760 17230
rect 6720 17200 6760 17210
rect 6800 18190 6840 18200
rect 6800 18170 6810 18190
rect 6830 18170 6840 18190
rect 6800 18030 6840 18170
rect 6800 18010 6810 18030
rect 6830 18010 6840 18030
rect 6800 17870 6840 18010
rect 6800 17850 6810 17870
rect 6830 17850 6840 17870
rect 6800 17710 6840 17850
rect 6800 17690 6810 17710
rect 6830 17690 6840 17710
rect 6800 17550 6840 17690
rect 6800 17530 6810 17550
rect 6830 17530 6840 17550
rect 6800 17390 6840 17530
rect 6800 17370 6810 17390
rect 6830 17370 6840 17390
rect 6800 17230 6840 17370
rect 6800 17210 6810 17230
rect 6830 17210 6840 17230
rect 6800 17200 6840 17210
rect 6880 18190 6920 18200
rect 6880 18170 6890 18190
rect 6910 18170 6920 18190
rect 6880 18030 6920 18170
rect 6880 18010 6890 18030
rect 6910 18010 6920 18030
rect 6880 17870 6920 18010
rect 6880 17850 6890 17870
rect 6910 17850 6920 17870
rect 6880 17710 6920 17850
rect 6880 17690 6890 17710
rect 6910 17690 6920 17710
rect 6880 17550 6920 17690
rect 6880 17530 6890 17550
rect 6910 17530 6920 17550
rect 6880 17390 6920 17530
rect 6880 17370 6890 17390
rect 6910 17370 6920 17390
rect 6880 17230 6920 17370
rect 6880 17210 6890 17230
rect 6910 17210 6920 17230
rect 6880 17200 6920 17210
rect 6960 18190 7000 18200
rect 6960 18170 6970 18190
rect 6990 18170 7000 18190
rect 6960 18030 7000 18170
rect 6960 18010 6970 18030
rect 6990 18010 7000 18030
rect 6960 17870 7000 18010
rect 6960 17850 6970 17870
rect 6990 17850 7000 17870
rect 6960 17710 7000 17850
rect 6960 17690 6970 17710
rect 6990 17690 7000 17710
rect 6960 17550 7000 17690
rect 6960 17530 6970 17550
rect 6990 17530 7000 17550
rect 6960 17390 7000 17530
rect 6960 17370 6970 17390
rect 6990 17370 7000 17390
rect 6960 17230 7000 17370
rect 6960 17210 6970 17230
rect 6990 17210 7000 17230
rect 6960 17200 7000 17210
rect 7040 18190 7080 18200
rect 7040 18170 7050 18190
rect 7070 18170 7080 18190
rect 7040 18030 7080 18170
rect 7040 18010 7050 18030
rect 7070 18010 7080 18030
rect 7040 17870 7080 18010
rect 7040 17850 7050 17870
rect 7070 17850 7080 17870
rect 7040 17710 7080 17850
rect 7040 17690 7050 17710
rect 7070 17690 7080 17710
rect 7040 17550 7080 17690
rect 7040 17530 7050 17550
rect 7070 17530 7080 17550
rect 7040 17390 7080 17530
rect 7040 17370 7050 17390
rect 7070 17370 7080 17390
rect 7040 17230 7080 17370
rect 7040 17210 7050 17230
rect 7070 17210 7080 17230
rect 7040 17200 7080 17210
rect 7120 18190 7160 18200
rect 7120 18170 7130 18190
rect 7150 18170 7160 18190
rect 7120 18030 7160 18170
rect 7120 18010 7130 18030
rect 7150 18010 7160 18030
rect 7120 17870 7160 18010
rect 7120 17850 7130 17870
rect 7150 17850 7160 17870
rect 7120 17710 7160 17850
rect 7120 17690 7130 17710
rect 7150 17690 7160 17710
rect 7120 17550 7160 17690
rect 7120 17530 7130 17550
rect 7150 17530 7160 17550
rect 7120 17390 7160 17530
rect 7120 17370 7130 17390
rect 7150 17370 7160 17390
rect 7120 17230 7160 17370
rect 7120 17210 7130 17230
rect 7150 17210 7160 17230
rect 7120 17200 7160 17210
rect 7200 18190 7240 18200
rect 7200 18170 7210 18190
rect 7230 18170 7240 18190
rect 7200 18030 7240 18170
rect 7200 18010 7210 18030
rect 7230 18010 7240 18030
rect 7200 17870 7240 18010
rect 7200 17850 7210 17870
rect 7230 17850 7240 17870
rect 7200 17710 7240 17850
rect 7200 17690 7210 17710
rect 7230 17690 7240 17710
rect 7200 17550 7240 17690
rect 7200 17530 7210 17550
rect 7230 17530 7240 17550
rect 7200 17390 7240 17530
rect 7200 17370 7210 17390
rect 7230 17370 7240 17390
rect 7200 17230 7240 17370
rect 7200 17210 7210 17230
rect 7230 17210 7240 17230
rect 7200 17200 7240 17210
rect 7280 18190 7320 18200
rect 7280 18170 7290 18190
rect 7310 18170 7320 18190
rect 7280 18030 7320 18170
rect 7280 18010 7290 18030
rect 7310 18010 7320 18030
rect 7280 17870 7320 18010
rect 7280 17850 7290 17870
rect 7310 17850 7320 17870
rect 7280 17710 7320 17850
rect 7280 17690 7290 17710
rect 7310 17690 7320 17710
rect 7280 17550 7320 17690
rect 7280 17530 7290 17550
rect 7310 17530 7320 17550
rect 7280 17390 7320 17530
rect 7280 17370 7290 17390
rect 7310 17370 7320 17390
rect 7280 17230 7320 17370
rect 7280 17210 7290 17230
rect 7310 17210 7320 17230
rect 7280 17200 7320 17210
rect 7360 18190 7400 18200
rect 7360 18170 7370 18190
rect 7390 18170 7400 18190
rect 7360 18030 7400 18170
rect 7360 18010 7370 18030
rect 7390 18010 7400 18030
rect 7360 17870 7400 18010
rect 7360 17850 7370 17870
rect 7390 17850 7400 17870
rect 7360 17710 7400 17850
rect 7360 17690 7370 17710
rect 7390 17690 7400 17710
rect 7360 17550 7400 17690
rect 7360 17530 7370 17550
rect 7390 17530 7400 17550
rect 7360 17390 7400 17530
rect 7360 17370 7370 17390
rect 7390 17370 7400 17390
rect 7360 17230 7400 17370
rect 7360 17210 7370 17230
rect 7390 17210 7400 17230
rect 7360 17200 7400 17210
rect 7440 18190 7480 18200
rect 7440 18170 7450 18190
rect 7470 18170 7480 18190
rect 7440 18030 7480 18170
rect 7440 18010 7450 18030
rect 7470 18010 7480 18030
rect 7440 17870 7480 18010
rect 7440 17850 7450 17870
rect 7470 17850 7480 17870
rect 7440 17710 7480 17850
rect 7440 17690 7450 17710
rect 7470 17690 7480 17710
rect 7440 17550 7480 17690
rect 7440 17530 7450 17550
rect 7470 17530 7480 17550
rect 7440 17390 7480 17530
rect 7440 17370 7450 17390
rect 7470 17370 7480 17390
rect 7440 17230 7480 17370
rect 7440 17210 7450 17230
rect 7470 17210 7480 17230
rect 7440 17200 7480 17210
rect 7520 18190 7560 18200
rect 7520 18170 7530 18190
rect 7550 18170 7560 18190
rect 7520 18030 7560 18170
rect 7520 18010 7530 18030
rect 7550 18010 7560 18030
rect 7520 17870 7560 18010
rect 7520 17850 7530 17870
rect 7550 17850 7560 17870
rect 7520 17710 7560 17850
rect 7520 17690 7530 17710
rect 7550 17690 7560 17710
rect 7520 17550 7560 17690
rect 7520 17530 7530 17550
rect 7550 17530 7560 17550
rect 7520 17390 7560 17530
rect 7520 17370 7530 17390
rect 7550 17370 7560 17390
rect 7520 17230 7560 17370
rect 7520 17210 7530 17230
rect 7550 17210 7560 17230
rect 7520 17200 7560 17210
rect 7600 18190 7640 18200
rect 7600 18170 7610 18190
rect 7630 18170 7640 18190
rect 7600 18030 7640 18170
rect 7600 18010 7610 18030
rect 7630 18010 7640 18030
rect 7600 17870 7640 18010
rect 7600 17850 7610 17870
rect 7630 17850 7640 17870
rect 7600 17710 7640 17850
rect 7600 17690 7610 17710
rect 7630 17690 7640 17710
rect 7600 17550 7640 17690
rect 7600 17530 7610 17550
rect 7630 17530 7640 17550
rect 7600 17390 7640 17530
rect 7600 17370 7610 17390
rect 7630 17370 7640 17390
rect 7600 17230 7640 17370
rect 7600 17210 7610 17230
rect 7630 17210 7640 17230
rect 7600 17200 7640 17210
rect 7680 18190 7720 18200
rect 7680 18170 7690 18190
rect 7710 18170 7720 18190
rect 7680 18030 7720 18170
rect 7680 18010 7690 18030
rect 7710 18010 7720 18030
rect 7680 17870 7720 18010
rect 7680 17850 7690 17870
rect 7710 17850 7720 17870
rect 7680 17710 7720 17850
rect 7680 17690 7690 17710
rect 7710 17690 7720 17710
rect 7680 17550 7720 17690
rect 7680 17530 7690 17550
rect 7710 17530 7720 17550
rect 7680 17390 7720 17530
rect 7680 17370 7690 17390
rect 7710 17370 7720 17390
rect 7680 17230 7720 17370
rect 7680 17210 7690 17230
rect 7710 17210 7720 17230
rect 7680 17200 7720 17210
rect 7760 18190 7800 18200
rect 7760 18170 7770 18190
rect 7790 18170 7800 18190
rect 7760 18030 7800 18170
rect 7760 18010 7770 18030
rect 7790 18010 7800 18030
rect 7760 17870 7800 18010
rect 7760 17850 7770 17870
rect 7790 17850 7800 17870
rect 7760 17710 7800 17850
rect 7760 17690 7770 17710
rect 7790 17690 7800 17710
rect 7760 17550 7800 17690
rect 7760 17530 7770 17550
rect 7790 17530 7800 17550
rect 7760 17390 7800 17530
rect 7760 17370 7770 17390
rect 7790 17370 7800 17390
rect 7760 17230 7800 17370
rect 7760 17210 7770 17230
rect 7790 17210 7800 17230
rect 7760 17200 7800 17210
rect 7840 18190 7880 18200
rect 7840 18170 7850 18190
rect 7870 18170 7880 18190
rect 7840 18030 7880 18170
rect 7840 18010 7850 18030
rect 7870 18010 7880 18030
rect 7840 17870 7880 18010
rect 7840 17850 7850 17870
rect 7870 17850 7880 17870
rect 7840 17710 7880 17850
rect 7840 17690 7850 17710
rect 7870 17690 7880 17710
rect 7840 17550 7880 17690
rect 7840 17530 7850 17550
rect 7870 17530 7880 17550
rect 7840 17390 7880 17530
rect 7840 17370 7850 17390
rect 7870 17370 7880 17390
rect 7840 17230 7880 17370
rect 7840 17210 7850 17230
rect 7870 17210 7880 17230
rect 7840 17200 7880 17210
rect 7920 18190 7960 18200
rect 7920 18170 7930 18190
rect 7950 18170 7960 18190
rect 7920 18030 7960 18170
rect 7920 18010 7930 18030
rect 7950 18010 7960 18030
rect 7920 17870 7960 18010
rect 7920 17850 7930 17870
rect 7950 17850 7960 17870
rect 7920 17710 7960 17850
rect 7920 17690 7930 17710
rect 7950 17690 7960 17710
rect 7920 17550 7960 17690
rect 7920 17530 7930 17550
rect 7950 17530 7960 17550
rect 7920 17390 7960 17530
rect 7920 17370 7930 17390
rect 7950 17370 7960 17390
rect 7920 17230 7960 17370
rect 7920 17210 7930 17230
rect 7950 17210 7960 17230
rect 7920 17200 7960 17210
rect 8000 18190 8040 18200
rect 8000 18170 8010 18190
rect 8030 18170 8040 18190
rect 8000 18030 8040 18170
rect 8000 18010 8010 18030
rect 8030 18010 8040 18030
rect 8000 17870 8040 18010
rect 8000 17850 8010 17870
rect 8030 17850 8040 17870
rect 8000 17710 8040 17850
rect 8000 17690 8010 17710
rect 8030 17690 8040 17710
rect 8000 17550 8040 17690
rect 8000 17530 8010 17550
rect 8030 17530 8040 17550
rect 8000 17390 8040 17530
rect 8000 17370 8010 17390
rect 8030 17370 8040 17390
rect 8000 17230 8040 17370
rect 8000 17210 8010 17230
rect 8030 17210 8040 17230
rect 8000 17200 8040 17210
rect 8080 18190 8120 18200
rect 8080 18170 8090 18190
rect 8110 18170 8120 18190
rect 8080 18030 8120 18170
rect 8080 18010 8090 18030
rect 8110 18010 8120 18030
rect 8080 17870 8120 18010
rect 8080 17850 8090 17870
rect 8110 17850 8120 17870
rect 8080 17710 8120 17850
rect 8080 17690 8090 17710
rect 8110 17690 8120 17710
rect 8080 17550 8120 17690
rect 8080 17530 8090 17550
rect 8110 17530 8120 17550
rect 8080 17390 8120 17530
rect 8080 17370 8090 17390
rect 8110 17370 8120 17390
rect 8080 17230 8120 17370
rect 8080 17210 8090 17230
rect 8110 17210 8120 17230
rect 8080 17200 8120 17210
rect 8160 18190 8200 18200
rect 8160 18170 8170 18190
rect 8190 18170 8200 18190
rect 8160 18030 8200 18170
rect 8160 18010 8170 18030
rect 8190 18010 8200 18030
rect 8160 17870 8200 18010
rect 8160 17850 8170 17870
rect 8190 17850 8200 17870
rect 8160 17710 8200 17850
rect 8160 17690 8170 17710
rect 8190 17690 8200 17710
rect 8160 17550 8200 17690
rect 8160 17530 8170 17550
rect 8190 17530 8200 17550
rect 8160 17390 8200 17530
rect 8160 17370 8170 17390
rect 8190 17370 8200 17390
rect 8160 17230 8200 17370
rect 8160 17210 8170 17230
rect 8190 17210 8200 17230
rect 8160 17200 8200 17210
rect 8240 18190 8280 18200
rect 8240 18170 8250 18190
rect 8270 18170 8280 18190
rect 8240 18030 8280 18170
rect 8240 18010 8250 18030
rect 8270 18010 8280 18030
rect 8240 17870 8280 18010
rect 8240 17850 8250 17870
rect 8270 17850 8280 17870
rect 8240 17710 8280 17850
rect 8240 17690 8250 17710
rect 8270 17690 8280 17710
rect 8240 17550 8280 17690
rect 8240 17530 8250 17550
rect 8270 17530 8280 17550
rect 8240 17390 8280 17530
rect 8240 17370 8250 17390
rect 8270 17370 8280 17390
rect 8240 17230 8280 17370
rect 8240 17210 8250 17230
rect 8270 17210 8280 17230
rect 8240 17200 8280 17210
rect 8320 18190 8360 18200
rect 8320 18170 8330 18190
rect 8350 18170 8360 18190
rect 8320 18030 8360 18170
rect 8320 18010 8330 18030
rect 8350 18010 8360 18030
rect 8320 17870 8360 18010
rect 8320 17850 8330 17870
rect 8350 17850 8360 17870
rect 8320 17710 8360 17850
rect 8320 17690 8330 17710
rect 8350 17690 8360 17710
rect 8320 17550 8360 17690
rect 8320 17530 8330 17550
rect 8350 17530 8360 17550
rect 8320 17390 8360 17530
rect 8320 17370 8330 17390
rect 8350 17370 8360 17390
rect 8320 17230 8360 17370
rect 8320 17210 8330 17230
rect 8350 17210 8360 17230
rect 8320 17200 8360 17210
rect 8400 18190 8440 18200
rect 8400 18170 8410 18190
rect 8430 18170 8440 18190
rect 8400 18030 8440 18170
rect 8400 18010 8410 18030
rect 8430 18010 8440 18030
rect 8400 17870 8440 18010
rect 8400 17850 8410 17870
rect 8430 17850 8440 17870
rect 8400 17710 8440 17850
rect 8400 17690 8410 17710
rect 8430 17690 8440 17710
rect 8400 17550 8440 17690
rect 8400 17530 8410 17550
rect 8430 17530 8440 17550
rect 8400 17390 8440 17530
rect 8400 17370 8410 17390
rect 8430 17370 8440 17390
rect 8400 17230 8440 17370
rect 8400 17210 8410 17230
rect 8430 17210 8440 17230
rect 8400 17200 8440 17210
rect 8480 18190 8520 18200
rect 8480 18170 8490 18190
rect 8510 18170 8520 18190
rect 8480 18030 8520 18170
rect 8480 18010 8490 18030
rect 8510 18010 8520 18030
rect 8480 17870 8520 18010
rect 8480 17850 8490 17870
rect 8510 17850 8520 17870
rect 8480 17710 8520 17850
rect 8480 17690 8490 17710
rect 8510 17690 8520 17710
rect 8480 17550 8520 17690
rect 8480 17530 8490 17550
rect 8510 17530 8520 17550
rect 8480 17390 8520 17530
rect 8480 17370 8490 17390
rect 8510 17370 8520 17390
rect 8480 17230 8520 17370
rect 8480 17210 8490 17230
rect 8510 17210 8520 17230
rect 8480 17200 8520 17210
rect 8560 18190 8600 18200
rect 8560 18170 8570 18190
rect 8590 18170 8600 18190
rect 8560 18030 8600 18170
rect 8560 18010 8570 18030
rect 8590 18010 8600 18030
rect 8560 17870 8600 18010
rect 8560 17850 8570 17870
rect 8590 17850 8600 17870
rect 8560 17710 8600 17850
rect 8560 17690 8570 17710
rect 8590 17690 8600 17710
rect 8560 17550 8600 17690
rect 8560 17530 8570 17550
rect 8590 17530 8600 17550
rect 8560 17390 8600 17530
rect 8560 17370 8570 17390
rect 8590 17370 8600 17390
rect 8560 17230 8600 17370
rect 8560 17210 8570 17230
rect 8590 17210 8600 17230
rect 8560 17200 8600 17210
rect 8640 18190 8680 18200
rect 8640 18170 8650 18190
rect 8670 18170 8680 18190
rect 8640 18030 8680 18170
rect 8640 18010 8650 18030
rect 8670 18010 8680 18030
rect 8640 17870 8680 18010
rect 8640 17850 8650 17870
rect 8670 17850 8680 17870
rect 8640 17710 8680 17850
rect 8640 17690 8650 17710
rect 8670 17690 8680 17710
rect 8640 17550 8680 17690
rect 8640 17530 8650 17550
rect 8670 17530 8680 17550
rect 8640 17390 8680 17530
rect 8640 17370 8650 17390
rect 8670 17370 8680 17390
rect 8640 17230 8680 17370
rect 8640 17210 8650 17230
rect 8670 17210 8680 17230
rect 8640 17200 8680 17210
rect 8720 18190 8760 18200
rect 8720 18170 8730 18190
rect 8750 18170 8760 18190
rect 8720 18030 8760 18170
rect 8720 18010 8730 18030
rect 8750 18010 8760 18030
rect 8720 17870 8760 18010
rect 8720 17850 8730 17870
rect 8750 17850 8760 17870
rect 8720 17710 8760 17850
rect 8720 17690 8730 17710
rect 8750 17690 8760 17710
rect 8720 17550 8760 17690
rect 8720 17530 8730 17550
rect 8750 17530 8760 17550
rect 8720 17390 8760 17530
rect 8720 17370 8730 17390
rect 8750 17370 8760 17390
rect 8720 17230 8760 17370
rect 8720 17210 8730 17230
rect 8750 17210 8760 17230
rect 8720 17200 8760 17210
rect 8800 18190 8840 18200
rect 8800 18170 8810 18190
rect 8830 18170 8840 18190
rect 8800 18030 8840 18170
rect 8800 18010 8810 18030
rect 8830 18010 8840 18030
rect 8800 17870 8840 18010
rect 8800 17850 8810 17870
rect 8830 17850 8840 17870
rect 8800 17710 8840 17850
rect 8800 17690 8810 17710
rect 8830 17690 8840 17710
rect 8800 17550 8840 17690
rect 8800 17530 8810 17550
rect 8830 17530 8840 17550
rect 8800 17390 8840 17530
rect 8800 17370 8810 17390
rect 8830 17370 8840 17390
rect 8800 17230 8840 17370
rect 8800 17210 8810 17230
rect 8830 17210 8840 17230
rect 8800 17200 8840 17210
rect 8880 18190 8920 18200
rect 8880 18170 8890 18190
rect 8910 18170 8920 18190
rect 8880 18030 8920 18170
rect 8880 18010 8890 18030
rect 8910 18010 8920 18030
rect 8880 17870 8920 18010
rect 8880 17850 8890 17870
rect 8910 17850 8920 17870
rect 8880 17710 8920 17850
rect 8880 17690 8890 17710
rect 8910 17690 8920 17710
rect 8880 17550 8920 17690
rect 8880 17530 8890 17550
rect 8910 17530 8920 17550
rect 8880 17390 8920 17530
rect 8880 17370 8890 17390
rect 8910 17370 8920 17390
rect 8880 17230 8920 17370
rect 8880 17210 8890 17230
rect 8910 17210 8920 17230
rect 8880 17200 8920 17210
rect 8960 18190 9000 18200
rect 8960 18170 8970 18190
rect 8990 18170 9000 18190
rect 8960 18030 9000 18170
rect 8960 18010 8970 18030
rect 8990 18010 9000 18030
rect 8960 17870 9000 18010
rect 8960 17850 8970 17870
rect 8990 17850 9000 17870
rect 8960 17710 9000 17850
rect 8960 17690 8970 17710
rect 8990 17690 9000 17710
rect 8960 17550 9000 17690
rect 8960 17530 8970 17550
rect 8990 17530 9000 17550
rect 8960 17390 9000 17530
rect 8960 17370 8970 17390
rect 8990 17370 9000 17390
rect 8960 17230 9000 17370
rect 8960 17210 8970 17230
rect 8990 17210 9000 17230
rect 8960 17200 9000 17210
rect 9040 18190 9080 18200
rect 9040 18170 9050 18190
rect 9070 18170 9080 18190
rect 9040 18030 9080 18170
rect 9040 18010 9050 18030
rect 9070 18010 9080 18030
rect 9040 17870 9080 18010
rect 9040 17850 9050 17870
rect 9070 17850 9080 17870
rect 9040 17710 9080 17850
rect 9040 17690 9050 17710
rect 9070 17690 9080 17710
rect 9040 17550 9080 17690
rect 9040 17530 9050 17550
rect 9070 17530 9080 17550
rect 9040 17390 9080 17530
rect 9040 17370 9050 17390
rect 9070 17370 9080 17390
rect 9040 17230 9080 17370
rect 9040 17210 9050 17230
rect 9070 17210 9080 17230
rect 9040 17200 9080 17210
rect 9120 18190 9160 18200
rect 9120 18170 9130 18190
rect 9150 18170 9160 18190
rect 9120 18030 9160 18170
rect 9120 18010 9130 18030
rect 9150 18010 9160 18030
rect 9120 17870 9160 18010
rect 9120 17850 9130 17870
rect 9150 17850 9160 17870
rect 9120 17710 9160 17850
rect 9120 17690 9130 17710
rect 9150 17690 9160 17710
rect 9120 17550 9160 17690
rect 9120 17530 9130 17550
rect 9150 17530 9160 17550
rect 9120 17390 9160 17530
rect 9120 17370 9130 17390
rect 9150 17370 9160 17390
rect 9120 17230 9160 17370
rect 9120 17210 9130 17230
rect 9150 17210 9160 17230
rect 9120 17200 9160 17210
rect 9200 18190 9240 18200
rect 9200 18170 9210 18190
rect 9230 18170 9240 18190
rect 9200 18030 9240 18170
rect 9200 18010 9210 18030
rect 9230 18010 9240 18030
rect 9200 17870 9240 18010
rect 9200 17850 9210 17870
rect 9230 17850 9240 17870
rect 9200 17710 9240 17850
rect 9200 17690 9210 17710
rect 9230 17690 9240 17710
rect 9200 17550 9240 17690
rect 9200 17530 9210 17550
rect 9230 17530 9240 17550
rect 9200 17390 9240 17530
rect 9200 17370 9210 17390
rect 9230 17370 9240 17390
rect 9200 17230 9240 17370
rect 9200 17210 9210 17230
rect 9230 17210 9240 17230
rect 9200 17200 9240 17210
rect 9280 18190 9320 18200
rect 9280 18170 9290 18190
rect 9310 18170 9320 18190
rect 9280 18030 9320 18170
rect 9280 18010 9290 18030
rect 9310 18010 9320 18030
rect 9280 17870 9320 18010
rect 9280 17850 9290 17870
rect 9310 17850 9320 17870
rect 9280 17710 9320 17850
rect 9280 17690 9290 17710
rect 9310 17690 9320 17710
rect 9280 17550 9320 17690
rect 9280 17530 9290 17550
rect 9310 17530 9320 17550
rect 9280 17390 9320 17530
rect 9280 17370 9290 17390
rect 9310 17370 9320 17390
rect 9280 17230 9320 17370
rect 9280 17210 9290 17230
rect 9310 17210 9320 17230
rect 9280 17200 9320 17210
rect 9360 18190 9400 18200
rect 9360 18170 9370 18190
rect 9390 18170 9400 18190
rect 9360 18030 9400 18170
rect 9360 18010 9370 18030
rect 9390 18010 9400 18030
rect 9360 17870 9400 18010
rect 9360 17850 9370 17870
rect 9390 17850 9400 17870
rect 9360 17710 9400 17850
rect 9360 17690 9370 17710
rect 9390 17690 9400 17710
rect 9360 17550 9400 17690
rect 9360 17530 9370 17550
rect 9390 17530 9400 17550
rect 9360 17390 9400 17530
rect 9360 17370 9370 17390
rect 9390 17370 9400 17390
rect 9360 17230 9400 17370
rect 9360 17210 9370 17230
rect 9390 17210 9400 17230
rect 9360 17200 9400 17210
rect 9440 18190 9480 18200
rect 9440 18170 9450 18190
rect 9470 18170 9480 18190
rect 9440 18030 9480 18170
rect 9440 18010 9450 18030
rect 9470 18010 9480 18030
rect 9440 17870 9480 18010
rect 9440 17850 9450 17870
rect 9470 17850 9480 17870
rect 9440 17710 9480 17850
rect 9440 17690 9450 17710
rect 9470 17690 9480 17710
rect 9440 17550 9480 17690
rect 9440 17530 9450 17550
rect 9470 17530 9480 17550
rect 9440 17390 9480 17530
rect 9440 17370 9450 17390
rect 9470 17370 9480 17390
rect 9440 17230 9480 17370
rect 9440 17210 9450 17230
rect 9470 17210 9480 17230
rect 9440 17200 9480 17210
rect 9520 17200 9560 18200
rect 9600 17200 9640 18200
rect 9680 17200 9720 18200
rect 9760 17200 9800 18200
rect 9840 17200 9880 18200
rect 9920 17200 9960 18200
rect 10000 17200 10040 18200
rect 10080 17200 10120 18200
rect 10160 17200 10200 18200
rect 10240 17200 10280 18200
rect 10320 17200 10360 18200
rect 10400 17200 10440 18200
rect 10480 17200 10520 18200
rect 10560 17200 10600 18200
rect 10640 17200 10680 18200
rect 10720 17200 10760 18200
rect 10800 17200 10840 18200
rect 10880 17200 10920 18200
rect 10960 17200 11000 18200
rect 11040 17200 11080 18200
rect 11120 17200 11160 18200
rect 11200 17200 11240 18200
rect 11280 17200 11320 18200
rect 11360 17200 11400 18200
rect 11440 17200 11480 18200
rect 11560 18190 11600 18200
rect 11560 18170 11570 18190
rect 11590 18170 11600 18190
rect 11560 18030 11600 18170
rect 11560 18010 11570 18030
rect 11590 18010 11600 18030
rect 11560 17870 11600 18010
rect 11560 17850 11570 17870
rect 11590 17850 11600 17870
rect 11560 17710 11600 17850
rect 11560 17690 11570 17710
rect 11590 17690 11600 17710
rect 11560 17550 11600 17690
rect 11560 17530 11570 17550
rect 11590 17530 11600 17550
rect 11560 17390 11600 17530
rect 11560 17370 11570 17390
rect 11590 17370 11600 17390
rect 11560 17230 11600 17370
rect 11560 17210 11570 17230
rect 11590 17210 11600 17230
rect 11560 17200 11600 17210
rect 11640 18190 11680 18200
rect 11640 18170 11650 18190
rect 11670 18170 11680 18190
rect 11640 18030 11680 18170
rect 11640 18010 11650 18030
rect 11670 18010 11680 18030
rect 11640 17870 11680 18010
rect 11640 17850 11650 17870
rect 11670 17850 11680 17870
rect 11640 17710 11680 17850
rect 11640 17690 11650 17710
rect 11670 17690 11680 17710
rect 11640 17550 11680 17690
rect 11640 17530 11650 17550
rect 11670 17530 11680 17550
rect 11640 17390 11680 17530
rect 11640 17370 11650 17390
rect 11670 17370 11680 17390
rect 11640 17230 11680 17370
rect 11640 17210 11650 17230
rect 11670 17210 11680 17230
rect 11640 17200 11680 17210
rect 11720 18190 11760 18200
rect 11720 18170 11730 18190
rect 11750 18170 11760 18190
rect 11720 18030 11760 18170
rect 11720 18010 11730 18030
rect 11750 18010 11760 18030
rect 11720 17870 11760 18010
rect 11720 17850 11730 17870
rect 11750 17850 11760 17870
rect 11720 17710 11760 17850
rect 11720 17690 11730 17710
rect 11750 17690 11760 17710
rect 11720 17550 11760 17690
rect 11720 17530 11730 17550
rect 11750 17530 11760 17550
rect 11720 17390 11760 17530
rect 11720 17370 11730 17390
rect 11750 17370 11760 17390
rect 11720 17230 11760 17370
rect 11720 17210 11730 17230
rect 11750 17210 11760 17230
rect 11720 17200 11760 17210
rect 11800 18190 11840 18200
rect 11800 18170 11810 18190
rect 11830 18170 11840 18190
rect 11800 18030 11840 18170
rect 11800 18010 11810 18030
rect 11830 18010 11840 18030
rect 11800 17870 11840 18010
rect 11800 17850 11810 17870
rect 11830 17850 11840 17870
rect 11800 17710 11840 17850
rect 11800 17690 11810 17710
rect 11830 17690 11840 17710
rect 11800 17550 11840 17690
rect 11800 17530 11810 17550
rect 11830 17530 11840 17550
rect 11800 17390 11840 17530
rect 11800 17370 11810 17390
rect 11830 17370 11840 17390
rect 11800 17230 11840 17370
rect 11800 17210 11810 17230
rect 11830 17210 11840 17230
rect 11800 17200 11840 17210
rect 11880 18190 11920 18200
rect 11880 18170 11890 18190
rect 11910 18170 11920 18190
rect 11880 18030 11920 18170
rect 11880 18010 11890 18030
rect 11910 18010 11920 18030
rect 11880 17870 11920 18010
rect 11880 17850 11890 17870
rect 11910 17850 11920 17870
rect 11880 17710 11920 17850
rect 11880 17690 11890 17710
rect 11910 17690 11920 17710
rect 11880 17550 11920 17690
rect 11880 17530 11890 17550
rect 11910 17530 11920 17550
rect 11880 17390 11920 17530
rect 11880 17370 11890 17390
rect 11910 17370 11920 17390
rect 11880 17230 11920 17370
rect 11880 17210 11890 17230
rect 11910 17210 11920 17230
rect 11880 17200 11920 17210
rect 11960 18190 12000 18200
rect 11960 18170 11970 18190
rect 11990 18170 12000 18190
rect 11960 18030 12000 18170
rect 11960 18010 11970 18030
rect 11990 18010 12000 18030
rect 11960 17870 12000 18010
rect 11960 17850 11970 17870
rect 11990 17850 12000 17870
rect 11960 17710 12000 17850
rect 11960 17690 11970 17710
rect 11990 17690 12000 17710
rect 11960 17550 12000 17690
rect 11960 17530 11970 17550
rect 11990 17530 12000 17550
rect 11960 17390 12000 17530
rect 11960 17370 11970 17390
rect 11990 17370 12000 17390
rect 11960 17230 12000 17370
rect 11960 17210 11970 17230
rect 11990 17210 12000 17230
rect 11960 17200 12000 17210
rect 12040 18190 12080 18200
rect 12040 18170 12050 18190
rect 12070 18170 12080 18190
rect 12040 18030 12080 18170
rect 12040 18010 12050 18030
rect 12070 18010 12080 18030
rect 12040 17870 12080 18010
rect 12040 17850 12050 17870
rect 12070 17850 12080 17870
rect 12040 17710 12080 17850
rect 12040 17690 12050 17710
rect 12070 17690 12080 17710
rect 12040 17550 12080 17690
rect 12040 17530 12050 17550
rect 12070 17530 12080 17550
rect 12040 17390 12080 17530
rect 12040 17370 12050 17390
rect 12070 17370 12080 17390
rect 12040 17230 12080 17370
rect 12040 17210 12050 17230
rect 12070 17210 12080 17230
rect 12040 17200 12080 17210
rect 12120 18190 12160 18200
rect 12120 18170 12130 18190
rect 12150 18170 12160 18190
rect 12120 18030 12160 18170
rect 12120 18010 12130 18030
rect 12150 18010 12160 18030
rect 12120 17870 12160 18010
rect 12120 17850 12130 17870
rect 12150 17850 12160 17870
rect 12120 17710 12160 17850
rect 12120 17690 12130 17710
rect 12150 17690 12160 17710
rect 12120 17550 12160 17690
rect 12120 17530 12130 17550
rect 12150 17530 12160 17550
rect 12120 17390 12160 17530
rect 12120 17370 12130 17390
rect 12150 17370 12160 17390
rect 12120 17230 12160 17370
rect 12120 17210 12130 17230
rect 12150 17210 12160 17230
rect 12120 17200 12160 17210
rect 12200 18190 12240 18200
rect 12200 18170 12210 18190
rect 12230 18170 12240 18190
rect 12200 18030 12240 18170
rect 12200 18010 12210 18030
rect 12230 18010 12240 18030
rect 12200 17870 12240 18010
rect 12200 17850 12210 17870
rect 12230 17850 12240 17870
rect 12200 17710 12240 17850
rect 12200 17690 12210 17710
rect 12230 17690 12240 17710
rect 12200 17550 12240 17690
rect 12200 17530 12210 17550
rect 12230 17530 12240 17550
rect 12200 17390 12240 17530
rect 12200 17370 12210 17390
rect 12230 17370 12240 17390
rect 12200 17230 12240 17370
rect 12200 17210 12210 17230
rect 12230 17210 12240 17230
rect 12200 17200 12240 17210
rect 12280 18190 12320 18200
rect 12280 18170 12290 18190
rect 12310 18170 12320 18190
rect 12280 18030 12320 18170
rect 12280 18010 12290 18030
rect 12310 18010 12320 18030
rect 12280 17870 12320 18010
rect 12280 17850 12290 17870
rect 12310 17850 12320 17870
rect 12280 17710 12320 17850
rect 12280 17690 12290 17710
rect 12310 17690 12320 17710
rect 12280 17550 12320 17690
rect 12280 17530 12290 17550
rect 12310 17530 12320 17550
rect 12280 17390 12320 17530
rect 12280 17370 12290 17390
rect 12310 17370 12320 17390
rect 12280 17230 12320 17370
rect 12280 17210 12290 17230
rect 12310 17210 12320 17230
rect 12280 17200 12320 17210
rect 12360 18190 12400 18200
rect 12360 18170 12370 18190
rect 12390 18170 12400 18190
rect 12360 18030 12400 18170
rect 12360 18010 12370 18030
rect 12390 18010 12400 18030
rect 12360 17870 12400 18010
rect 12360 17850 12370 17870
rect 12390 17850 12400 17870
rect 12360 17710 12400 17850
rect 12360 17690 12370 17710
rect 12390 17690 12400 17710
rect 12360 17550 12400 17690
rect 12360 17530 12370 17550
rect 12390 17530 12400 17550
rect 12360 17390 12400 17530
rect 12360 17370 12370 17390
rect 12390 17370 12400 17390
rect 12360 17230 12400 17370
rect 12360 17210 12370 17230
rect 12390 17210 12400 17230
rect 12360 17200 12400 17210
rect 12440 18190 12480 18200
rect 12440 18170 12450 18190
rect 12470 18170 12480 18190
rect 12440 18030 12480 18170
rect 12440 18010 12450 18030
rect 12470 18010 12480 18030
rect 12440 17870 12480 18010
rect 12440 17850 12450 17870
rect 12470 17850 12480 17870
rect 12440 17710 12480 17850
rect 12440 17690 12450 17710
rect 12470 17690 12480 17710
rect 12440 17550 12480 17690
rect 12440 17530 12450 17550
rect 12470 17530 12480 17550
rect 12440 17390 12480 17530
rect 12440 17370 12450 17390
rect 12470 17370 12480 17390
rect 12440 17230 12480 17370
rect 12440 17210 12450 17230
rect 12470 17210 12480 17230
rect 12440 17200 12480 17210
rect 12520 18190 12560 18200
rect 12520 18170 12530 18190
rect 12550 18170 12560 18190
rect 12520 18030 12560 18170
rect 12520 18010 12530 18030
rect 12550 18010 12560 18030
rect 12520 17870 12560 18010
rect 12520 17850 12530 17870
rect 12550 17850 12560 17870
rect 12520 17710 12560 17850
rect 12520 17690 12530 17710
rect 12550 17690 12560 17710
rect 12520 17550 12560 17690
rect 12520 17530 12530 17550
rect 12550 17530 12560 17550
rect 12520 17390 12560 17530
rect 12520 17370 12530 17390
rect 12550 17370 12560 17390
rect 12520 17230 12560 17370
rect 12520 17210 12530 17230
rect 12550 17210 12560 17230
rect 12520 17200 12560 17210
rect 12600 18190 12640 18200
rect 12600 18170 12610 18190
rect 12630 18170 12640 18190
rect 12600 18030 12640 18170
rect 12600 18010 12610 18030
rect 12630 18010 12640 18030
rect 12600 17870 12640 18010
rect 12600 17850 12610 17870
rect 12630 17850 12640 17870
rect 12600 17710 12640 17850
rect 12600 17690 12610 17710
rect 12630 17690 12640 17710
rect 12600 17550 12640 17690
rect 12600 17530 12610 17550
rect 12630 17530 12640 17550
rect 12600 17390 12640 17530
rect 12600 17370 12610 17390
rect 12630 17370 12640 17390
rect 12600 17230 12640 17370
rect 12600 17210 12610 17230
rect 12630 17210 12640 17230
rect 12600 17200 12640 17210
rect 12680 18190 12720 18200
rect 12680 18170 12690 18190
rect 12710 18170 12720 18190
rect 12680 18030 12720 18170
rect 12680 18010 12690 18030
rect 12710 18010 12720 18030
rect 12680 17870 12720 18010
rect 12680 17850 12690 17870
rect 12710 17850 12720 17870
rect 12680 17710 12720 17850
rect 12680 17690 12690 17710
rect 12710 17690 12720 17710
rect 12680 17550 12720 17690
rect 12680 17530 12690 17550
rect 12710 17530 12720 17550
rect 12680 17390 12720 17530
rect 12680 17370 12690 17390
rect 12710 17370 12720 17390
rect 12680 17230 12720 17370
rect 12680 17210 12690 17230
rect 12710 17210 12720 17230
rect 12680 17200 12720 17210
rect 12760 18190 12800 18200
rect 12760 18170 12770 18190
rect 12790 18170 12800 18190
rect 12760 18030 12800 18170
rect 12760 18010 12770 18030
rect 12790 18010 12800 18030
rect 12760 17870 12800 18010
rect 12760 17850 12770 17870
rect 12790 17850 12800 17870
rect 12760 17710 12800 17850
rect 12760 17690 12770 17710
rect 12790 17690 12800 17710
rect 12760 17550 12800 17690
rect 12760 17530 12770 17550
rect 12790 17530 12800 17550
rect 12760 17390 12800 17530
rect 12760 17370 12770 17390
rect 12790 17370 12800 17390
rect 12760 17230 12800 17370
rect 12760 17210 12770 17230
rect 12790 17210 12800 17230
rect 12760 17200 12800 17210
rect 12840 18190 12880 18200
rect 12840 18170 12850 18190
rect 12870 18170 12880 18190
rect 12840 18030 12880 18170
rect 12840 18010 12850 18030
rect 12870 18010 12880 18030
rect 12840 17870 12880 18010
rect 12840 17850 12850 17870
rect 12870 17850 12880 17870
rect 12840 17710 12880 17850
rect 12840 17690 12850 17710
rect 12870 17690 12880 17710
rect 12840 17550 12880 17690
rect 12840 17530 12850 17550
rect 12870 17530 12880 17550
rect 12840 17390 12880 17530
rect 12840 17370 12850 17390
rect 12870 17370 12880 17390
rect 12840 17230 12880 17370
rect 12840 17210 12850 17230
rect 12870 17210 12880 17230
rect 12840 17200 12880 17210
rect 12920 18190 12960 18200
rect 12920 18170 12930 18190
rect 12950 18170 12960 18190
rect 12920 18030 12960 18170
rect 12920 18010 12930 18030
rect 12950 18010 12960 18030
rect 12920 17870 12960 18010
rect 12920 17850 12930 17870
rect 12950 17850 12960 17870
rect 12920 17710 12960 17850
rect 12920 17690 12930 17710
rect 12950 17690 12960 17710
rect 12920 17550 12960 17690
rect 12920 17530 12930 17550
rect 12950 17530 12960 17550
rect 12920 17390 12960 17530
rect 12920 17370 12930 17390
rect 12950 17370 12960 17390
rect 12920 17230 12960 17370
rect 12920 17210 12930 17230
rect 12950 17210 12960 17230
rect 12920 17200 12960 17210
rect 13000 18190 13040 18200
rect 13000 18170 13010 18190
rect 13030 18170 13040 18190
rect 13000 18030 13040 18170
rect 13000 18010 13010 18030
rect 13030 18010 13040 18030
rect 13000 17870 13040 18010
rect 13000 17850 13010 17870
rect 13030 17850 13040 17870
rect 13000 17710 13040 17850
rect 13000 17690 13010 17710
rect 13030 17690 13040 17710
rect 13000 17550 13040 17690
rect 13000 17530 13010 17550
rect 13030 17530 13040 17550
rect 13000 17390 13040 17530
rect 13000 17370 13010 17390
rect 13030 17370 13040 17390
rect 13000 17230 13040 17370
rect 13000 17210 13010 17230
rect 13030 17210 13040 17230
rect 13000 17200 13040 17210
rect 13080 18190 13120 18200
rect 13080 18170 13090 18190
rect 13110 18170 13120 18190
rect 13080 18030 13120 18170
rect 13080 18010 13090 18030
rect 13110 18010 13120 18030
rect 13080 17870 13120 18010
rect 13080 17850 13090 17870
rect 13110 17850 13120 17870
rect 13080 17710 13120 17850
rect 13080 17690 13090 17710
rect 13110 17690 13120 17710
rect 13080 17550 13120 17690
rect 13080 17530 13090 17550
rect 13110 17530 13120 17550
rect 13080 17390 13120 17530
rect 13080 17370 13090 17390
rect 13110 17370 13120 17390
rect 13080 17230 13120 17370
rect 13080 17210 13090 17230
rect 13110 17210 13120 17230
rect 13080 17200 13120 17210
rect 13160 18190 13200 18200
rect 13160 18170 13170 18190
rect 13190 18170 13200 18190
rect 13160 18030 13200 18170
rect 13160 18010 13170 18030
rect 13190 18010 13200 18030
rect 13160 17870 13200 18010
rect 13160 17850 13170 17870
rect 13190 17850 13200 17870
rect 13160 17710 13200 17850
rect 13160 17690 13170 17710
rect 13190 17690 13200 17710
rect 13160 17550 13200 17690
rect 13160 17530 13170 17550
rect 13190 17530 13200 17550
rect 13160 17390 13200 17530
rect 13160 17370 13170 17390
rect 13190 17370 13200 17390
rect 13160 17230 13200 17370
rect 13160 17210 13170 17230
rect 13190 17210 13200 17230
rect 13160 17200 13200 17210
rect 13240 18190 13280 18200
rect 13240 18170 13250 18190
rect 13270 18170 13280 18190
rect 13240 18030 13280 18170
rect 13240 18010 13250 18030
rect 13270 18010 13280 18030
rect 13240 17870 13280 18010
rect 13240 17850 13250 17870
rect 13270 17850 13280 17870
rect 13240 17710 13280 17850
rect 13240 17690 13250 17710
rect 13270 17690 13280 17710
rect 13240 17550 13280 17690
rect 13240 17530 13250 17550
rect 13270 17530 13280 17550
rect 13240 17390 13280 17530
rect 13240 17370 13250 17390
rect 13270 17370 13280 17390
rect 13240 17230 13280 17370
rect 13240 17210 13250 17230
rect 13270 17210 13280 17230
rect 13240 17200 13280 17210
rect 13320 18190 13360 18200
rect 13320 18170 13330 18190
rect 13350 18170 13360 18190
rect 13320 18030 13360 18170
rect 13320 18010 13330 18030
rect 13350 18010 13360 18030
rect 13320 17870 13360 18010
rect 13320 17850 13330 17870
rect 13350 17850 13360 17870
rect 13320 17710 13360 17850
rect 13320 17690 13330 17710
rect 13350 17690 13360 17710
rect 13320 17550 13360 17690
rect 13320 17530 13330 17550
rect 13350 17530 13360 17550
rect 13320 17390 13360 17530
rect 13320 17370 13330 17390
rect 13350 17370 13360 17390
rect 13320 17230 13360 17370
rect 13320 17210 13330 17230
rect 13350 17210 13360 17230
rect 13320 17200 13360 17210
rect 13400 18190 13440 18200
rect 13400 18170 13410 18190
rect 13430 18170 13440 18190
rect 13400 18030 13440 18170
rect 13400 18010 13410 18030
rect 13430 18010 13440 18030
rect 13400 17870 13440 18010
rect 13400 17850 13410 17870
rect 13430 17850 13440 17870
rect 13400 17710 13440 17850
rect 13400 17690 13410 17710
rect 13430 17690 13440 17710
rect 13400 17550 13440 17690
rect 13400 17530 13410 17550
rect 13430 17530 13440 17550
rect 13400 17390 13440 17530
rect 13400 17370 13410 17390
rect 13430 17370 13440 17390
rect 13400 17230 13440 17370
rect 13400 17210 13410 17230
rect 13430 17210 13440 17230
rect 13400 17200 13440 17210
rect 13480 18190 13520 18200
rect 13480 18170 13490 18190
rect 13510 18170 13520 18190
rect 13480 18030 13520 18170
rect 13480 18010 13490 18030
rect 13510 18010 13520 18030
rect 13480 17870 13520 18010
rect 13480 17850 13490 17870
rect 13510 17850 13520 17870
rect 13480 17710 13520 17850
rect 13480 17690 13490 17710
rect 13510 17690 13520 17710
rect 13480 17550 13520 17690
rect 13480 17530 13490 17550
rect 13510 17530 13520 17550
rect 13480 17390 13520 17530
rect 13480 17370 13490 17390
rect 13510 17370 13520 17390
rect 13480 17230 13520 17370
rect 13480 17210 13490 17230
rect 13510 17210 13520 17230
rect 13480 17200 13520 17210
rect 13560 18190 13600 18200
rect 13560 18170 13570 18190
rect 13590 18170 13600 18190
rect 13560 18030 13600 18170
rect 13560 18010 13570 18030
rect 13590 18010 13600 18030
rect 13560 17870 13600 18010
rect 13560 17850 13570 17870
rect 13590 17850 13600 17870
rect 13560 17710 13600 17850
rect 13560 17690 13570 17710
rect 13590 17690 13600 17710
rect 13560 17550 13600 17690
rect 13560 17530 13570 17550
rect 13590 17530 13600 17550
rect 13560 17390 13600 17530
rect 13560 17370 13570 17390
rect 13590 17370 13600 17390
rect 13560 17230 13600 17370
rect 13560 17210 13570 17230
rect 13590 17210 13600 17230
rect 13560 17200 13600 17210
rect 13640 18190 13680 18200
rect 13640 18170 13650 18190
rect 13670 18170 13680 18190
rect 13640 18030 13680 18170
rect 13640 18010 13650 18030
rect 13670 18010 13680 18030
rect 13640 17870 13680 18010
rect 13640 17850 13650 17870
rect 13670 17850 13680 17870
rect 13640 17710 13680 17850
rect 13640 17690 13650 17710
rect 13670 17690 13680 17710
rect 13640 17550 13680 17690
rect 13640 17530 13650 17550
rect 13670 17530 13680 17550
rect 13640 17390 13680 17530
rect 13640 17370 13650 17390
rect 13670 17370 13680 17390
rect 13640 17230 13680 17370
rect 13640 17210 13650 17230
rect 13670 17210 13680 17230
rect 13640 17200 13680 17210
rect 13720 18190 13760 18200
rect 13720 18170 13730 18190
rect 13750 18170 13760 18190
rect 13720 18030 13760 18170
rect 13720 18010 13730 18030
rect 13750 18010 13760 18030
rect 13720 17870 13760 18010
rect 13720 17850 13730 17870
rect 13750 17850 13760 17870
rect 13720 17710 13760 17850
rect 13720 17690 13730 17710
rect 13750 17690 13760 17710
rect 13720 17550 13760 17690
rect 13720 17530 13730 17550
rect 13750 17530 13760 17550
rect 13720 17390 13760 17530
rect 13720 17370 13730 17390
rect 13750 17370 13760 17390
rect 13720 17230 13760 17370
rect 13720 17210 13730 17230
rect 13750 17210 13760 17230
rect 13720 17200 13760 17210
rect 13800 18190 13840 18200
rect 13800 18170 13810 18190
rect 13830 18170 13840 18190
rect 13800 18030 13840 18170
rect 13800 18010 13810 18030
rect 13830 18010 13840 18030
rect 13800 17870 13840 18010
rect 13800 17850 13810 17870
rect 13830 17850 13840 17870
rect 13800 17710 13840 17850
rect 13800 17690 13810 17710
rect 13830 17690 13840 17710
rect 13800 17550 13840 17690
rect 13800 17530 13810 17550
rect 13830 17530 13840 17550
rect 13800 17390 13840 17530
rect 13800 17370 13810 17390
rect 13830 17370 13840 17390
rect 13800 17230 13840 17370
rect 13800 17210 13810 17230
rect 13830 17210 13840 17230
rect 13800 17200 13840 17210
rect 13880 18190 13920 18200
rect 13880 18170 13890 18190
rect 13910 18170 13920 18190
rect 13880 18030 13920 18170
rect 13880 18010 13890 18030
rect 13910 18010 13920 18030
rect 13880 17870 13920 18010
rect 13880 17850 13890 17870
rect 13910 17850 13920 17870
rect 13880 17710 13920 17850
rect 13880 17690 13890 17710
rect 13910 17690 13920 17710
rect 13880 17550 13920 17690
rect 13880 17530 13890 17550
rect 13910 17530 13920 17550
rect 13880 17390 13920 17530
rect 13880 17370 13890 17390
rect 13910 17370 13920 17390
rect 13880 17230 13920 17370
rect 13880 17210 13890 17230
rect 13910 17210 13920 17230
rect 13880 17200 13920 17210
rect 13960 18190 14000 18200
rect 13960 18170 13970 18190
rect 13990 18170 14000 18190
rect 13960 18030 14000 18170
rect 13960 18010 13970 18030
rect 13990 18010 14000 18030
rect 13960 17870 14000 18010
rect 13960 17850 13970 17870
rect 13990 17850 14000 17870
rect 13960 17710 14000 17850
rect 13960 17690 13970 17710
rect 13990 17690 14000 17710
rect 13960 17550 14000 17690
rect 13960 17530 13970 17550
rect 13990 17530 14000 17550
rect 13960 17390 14000 17530
rect 13960 17370 13970 17390
rect 13990 17370 14000 17390
rect 13960 17230 14000 17370
rect 13960 17210 13970 17230
rect 13990 17210 14000 17230
rect 13960 17200 14000 17210
rect 14040 18190 14080 18200
rect 14040 18170 14050 18190
rect 14070 18170 14080 18190
rect 14040 18030 14080 18170
rect 14040 18010 14050 18030
rect 14070 18010 14080 18030
rect 14040 17870 14080 18010
rect 14040 17850 14050 17870
rect 14070 17850 14080 17870
rect 14040 17710 14080 17850
rect 14040 17690 14050 17710
rect 14070 17690 14080 17710
rect 14040 17550 14080 17690
rect 14040 17530 14050 17550
rect 14070 17530 14080 17550
rect 14040 17390 14080 17530
rect 14040 17370 14050 17390
rect 14070 17370 14080 17390
rect 14040 17230 14080 17370
rect 14040 17210 14050 17230
rect 14070 17210 14080 17230
rect 14040 17200 14080 17210
rect 14120 18190 14160 18200
rect 14120 18170 14130 18190
rect 14150 18170 14160 18190
rect 14120 18030 14160 18170
rect 14120 18010 14130 18030
rect 14150 18010 14160 18030
rect 14120 17870 14160 18010
rect 14120 17850 14130 17870
rect 14150 17850 14160 17870
rect 14120 17710 14160 17850
rect 14120 17690 14130 17710
rect 14150 17690 14160 17710
rect 14120 17550 14160 17690
rect 14120 17530 14130 17550
rect 14150 17530 14160 17550
rect 14120 17390 14160 17530
rect 14120 17370 14130 17390
rect 14150 17370 14160 17390
rect 14120 17230 14160 17370
rect 14120 17210 14130 17230
rect 14150 17210 14160 17230
rect 14120 17200 14160 17210
rect 14200 18190 14240 18200
rect 14200 18170 14210 18190
rect 14230 18170 14240 18190
rect 14200 18030 14240 18170
rect 14200 18010 14210 18030
rect 14230 18010 14240 18030
rect 14200 17870 14240 18010
rect 14200 17850 14210 17870
rect 14230 17850 14240 17870
rect 14200 17710 14240 17850
rect 14200 17690 14210 17710
rect 14230 17690 14240 17710
rect 14200 17550 14240 17690
rect 14200 17530 14210 17550
rect 14230 17530 14240 17550
rect 14200 17390 14240 17530
rect 14200 17370 14210 17390
rect 14230 17370 14240 17390
rect 14200 17230 14240 17370
rect 14200 17210 14210 17230
rect 14230 17210 14240 17230
rect 14200 17200 14240 17210
rect 14280 18190 14320 18200
rect 14280 18170 14290 18190
rect 14310 18170 14320 18190
rect 14280 18030 14320 18170
rect 14280 18010 14290 18030
rect 14310 18010 14320 18030
rect 14280 17870 14320 18010
rect 14280 17850 14290 17870
rect 14310 17850 14320 17870
rect 14280 17710 14320 17850
rect 14280 17690 14290 17710
rect 14310 17690 14320 17710
rect 14280 17550 14320 17690
rect 14280 17530 14290 17550
rect 14310 17530 14320 17550
rect 14280 17390 14320 17530
rect 14280 17370 14290 17390
rect 14310 17370 14320 17390
rect 14280 17230 14320 17370
rect 14280 17210 14290 17230
rect 14310 17210 14320 17230
rect 14280 17200 14320 17210
rect 14360 18190 14400 18200
rect 14360 18170 14370 18190
rect 14390 18170 14400 18190
rect 14360 18030 14400 18170
rect 14360 18010 14370 18030
rect 14390 18010 14400 18030
rect 14360 17870 14400 18010
rect 14360 17850 14370 17870
rect 14390 17850 14400 17870
rect 14360 17710 14400 17850
rect 14360 17690 14370 17710
rect 14390 17690 14400 17710
rect 14360 17550 14400 17690
rect 14360 17530 14370 17550
rect 14390 17530 14400 17550
rect 14360 17390 14400 17530
rect 14360 17370 14370 17390
rect 14390 17370 14400 17390
rect 14360 17230 14400 17370
rect 14360 17210 14370 17230
rect 14390 17210 14400 17230
rect 14360 17200 14400 17210
rect 14440 18190 14480 18200
rect 14440 18170 14450 18190
rect 14470 18170 14480 18190
rect 14440 18030 14480 18170
rect 14440 18010 14450 18030
rect 14470 18010 14480 18030
rect 14440 17870 14480 18010
rect 14440 17850 14450 17870
rect 14470 17850 14480 17870
rect 14440 17710 14480 17850
rect 14440 17690 14450 17710
rect 14470 17690 14480 17710
rect 14440 17550 14480 17690
rect 14440 17530 14450 17550
rect 14470 17530 14480 17550
rect 14440 17390 14480 17530
rect 14440 17370 14450 17390
rect 14470 17370 14480 17390
rect 14440 17230 14480 17370
rect 14440 17210 14450 17230
rect 14470 17210 14480 17230
rect 14440 17200 14480 17210
rect 14520 18190 14560 18200
rect 14520 18170 14530 18190
rect 14550 18170 14560 18190
rect 14520 18030 14560 18170
rect 14520 18010 14530 18030
rect 14550 18010 14560 18030
rect 14520 17870 14560 18010
rect 14520 17850 14530 17870
rect 14550 17850 14560 17870
rect 14520 17710 14560 17850
rect 14520 17690 14530 17710
rect 14550 17690 14560 17710
rect 14520 17550 14560 17690
rect 14520 17530 14530 17550
rect 14550 17530 14560 17550
rect 14520 17390 14560 17530
rect 14520 17370 14530 17390
rect 14550 17370 14560 17390
rect 14520 17230 14560 17370
rect 14520 17210 14530 17230
rect 14550 17210 14560 17230
rect 14520 17200 14560 17210
rect 14600 18190 14640 18200
rect 14600 18170 14610 18190
rect 14630 18170 14640 18190
rect 14600 18030 14640 18170
rect 14600 18010 14610 18030
rect 14630 18010 14640 18030
rect 14600 17870 14640 18010
rect 14600 17850 14610 17870
rect 14630 17850 14640 17870
rect 14600 17710 14640 17850
rect 14600 17690 14610 17710
rect 14630 17690 14640 17710
rect 14600 17550 14640 17690
rect 14600 17530 14610 17550
rect 14630 17530 14640 17550
rect 14600 17390 14640 17530
rect 14600 17370 14610 17390
rect 14630 17370 14640 17390
rect 14600 17230 14640 17370
rect 14600 17210 14610 17230
rect 14630 17210 14640 17230
rect 14600 17200 14640 17210
rect 14680 18190 14720 18200
rect 14680 18170 14690 18190
rect 14710 18170 14720 18190
rect 14680 18030 14720 18170
rect 14680 18010 14690 18030
rect 14710 18010 14720 18030
rect 14680 17870 14720 18010
rect 14680 17850 14690 17870
rect 14710 17850 14720 17870
rect 14680 17710 14720 17850
rect 14680 17690 14690 17710
rect 14710 17690 14720 17710
rect 14680 17550 14720 17690
rect 14680 17530 14690 17550
rect 14710 17530 14720 17550
rect 14680 17390 14720 17530
rect 14680 17370 14690 17390
rect 14710 17370 14720 17390
rect 14680 17230 14720 17370
rect 14680 17210 14690 17230
rect 14710 17210 14720 17230
rect 14680 17200 14720 17210
rect 14760 17200 14800 18200
rect 14840 17200 14880 18200
rect 14920 17200 14960 18200
rect 15000 17200 15040 18200
rect 15080 17200 15120 18200
rect 15160 17200 15200 18200
rect 15240 17200 15280 18200
rect 15320 17200 15360 18200
rect 15400 17200 15440 18200
rect 15480 17200 15520 18200
rect 15560 17200 15600 18200
rect 15640 17200 15680 18200
rect 15720 17200 15760 18200
rect 15800 17200 15840 18200
rect 15880 17200 15920 18200
rect 15960 17200 16000 18200
rect 16040 17200 16080 18200
rect 16120 17200 16160 18200
rect 16200 17200 16240 18200
rect 16280 17200 16320 18200
rect 16360 17200 16400 18200
rect 16440 17200 16480 18200
rect 16520 17200 16560 18200
rect 16600 17200 16640 18200
rect 16680 17200 16720 18200
rect 16760 18190 16800 18200
rect 16760 18170 16770 18190
rect 16790 18170 16800 18190
rect 16760 18030 16800 18170
rect 16760 18010 16770 18030
rect 16790 18010 16800 18030
rect 16760 17870 16800 18010
rect 16760 17850 16770 17870
rect 16790 17850 16800 17870
rect 16760 17710 16800 17850
rect 16760 17690 16770 17710
rect 16790 17690 16800 17710
rect 16760 17550 16800 17690
rect 16760 17530 16770 17550
rect 16790 17530 16800 17550
rect 16760 17390 16800 17530
rect 16760 17370 16770 17390
rect 16790 17370 16800 17390
rect 16760 17230 16800 17370
rect 16760 17210 16770 17230
rect 16790 17210 16800 17230
rect 16760 17200 16800 17210
rect 16840 18190 16880 18200
rect 16840 18170 16850 18190
rect 16870 18170 16880 18190
rect 16840 18030 16880 18170
rect 16840 18010 16850 18030
rect 16870 18010 16880 18030
rect 16840 17870 16880 18010
rect 16840 17850 16850 17870
rect 16870 17850 16880 17870
rect 16840 17710 16880 17850
rect 16840 17690 16850 17710
rect 16870 17690 16880 17710
rect 16840 17550 16880 17690
rect 16840 17530 16850 17550
rect 16870 17530 16880 17550
rect 16840 17390 16880 17530
rect 16840 17370 16850 17390
rect 16870 17370 16880 17390
rect 16840 17230 16880 17370
rect 16840 17210 16850 17230
rect 16870 17210 16880 17230
rect 16840 17200 16880 17210
rect 16920 18190 16960 18200
rect 16920 18170 16930 18190
rect 16950 18170 16960 18190
rect 16920 18030 16960 18170
rect 16920 18010 16930 18030
rect 16950 18010 16960 18030
rect 16920 17870 16960 18010
rect 16920 17850 16930 17870
rect 16950 17850 16960 17870
rect 16920 17710 16960 17850
rect 16920 17690 16930 17710
rect 16950 17690 16960 17710
rect 16920 17550 16960 17690
rect 16920 17530 16930 17550
rect 16950 17530 16960 17550
rect 16920 17390 16960 17530
rect 16920 17370 16930 17390
rect 16950 17370 16960 17390
rect 16920 17230 16960 17370
rect 16920 17210 16930 17230
rect 16950 17210 16960 17230
rect 16920 17200 16960 17210
rect 17000 18190 17040 18200
rect 17000 18170 17010 18190
rect 17030 18170 17040 18190
rect 17000 18030 17040 18170
rect 17000 18010 17010 18030
rect 17030 18010 17040 18030
rect 17000 17870 17040 18010
rect 17000 17850 17010 17870
rect 17030 17850 17040 17870
rect 17000 17710 17040 17850
rect 17000 17690 17010 17710
rect 17030 17690 17040 17710
rect 17000 17550 17040 17690
rect 17000 17530 17010 17550
rect 17030 17530 17040 17550
rect 17000 17390 17040 17530
rect 17000 17370 17010 17390
rect 17030 17370 17040 17390
rect 17000 17230 17040 17370
rect 17000 17210 17010 17230
rect 17030 17210 17040 17230
rect 17000 17200 17040 17210
rect 17080 18190 17120 18200
rect 17080 18170 17090 18190
rect 17110 18170 17120 18190
rect 17080 18030 17120 18170
rect 17080 18010 17090 18030
rect 17110 18010 17120 18030
rect 17080 17870 17120 18010
rect 17080 17850 17090 17870
rect 17110 17850 17120 17870
rect 17080 17710 17120 17850
rect 17080 17690 17090 17710
rect 17110 17690 17120 17710
rect 17080 17550 17120 17690
rect 17080 17530 17090 17550
rect 17110 17530 17120 17550
rect 17080 17390 17120 17530
rect 17080 17370 17090 17390
rect 17110 17370 17120 17390
rect 17080 17230 17120 17370
rect 17080 17210 17090 17230
rect 17110 17210 17120 17230
rect 17080 17200 17120 17210
rect 17160 18190 17200 18200
rect 17160 18170 17170 18190
rect 17190 18170 17200 18190
rect 17160 18030 17200 18170
rect 17160 18010 17170 18030
rect 17190 18010 17200 18030
rect 17160 17870 17200 18010
rect 17160 17850 17170 17870
rect 17190 17850 17200 17870
rect 17160 17710 17200 17850
rect 17160 17690 17170 17710
rect 17190 17690 17200 17710
rect 17160 17550 17200 17690
rect 17160 17530 17170 17550
rect 17190 17530 17200 17550
rect 17160 17390 17200 17530
rect 17160 17370 17170 17390
rect 17190 17370 17200 17390
rect 17160 17230 17200 17370
rect 17160 17210 17170 17230
rect 17190 17210 17200 17230
rect 17160 17200 17200 17210
rect 17240 18190 17280 18200
rect 17240 18170 17250 18190
rect 17270 18170 17280 18190
rect 17240 18030 17280 18170
rect 17240 18010 17250 18030
rect 17270 18010 17280 18030
rect 17240 17870 17280 18010
rect 17240 17850 17250 17870
rect 17270 17850 17280 17870
rect 17240 17710 17280 17850
rect 17240 17690 17250 17710
rect 17270 17690 17280 17710
rect 17240 17550 17280 17690
rect 17240 17530 17250 17550
rect 17270 17530 17280 17550
rect 17240 17390 17280 17530
rect 17240 17370 17250 17390
rect 17270 17370 17280 17390
rect 17240 17230 17280 17370
rect 17240 17210 17250 17230
rect 17270 17210 17280 17230
rect 17240 17200 17280 17210
rect 17320 18190 17360 18200
rect 17320 18170 17330 18190
rect 17350 18170 17360 18190
rect 17320 18030 17360 18170
rect 17320 18010 17330 18030
rect 17350 18010 17360 18030
rect 17320 17870 17360 18010
rect 17320 17850 17330 17870
rect 17350 17850 17360 17870
rect 17320 17710 17360 17850
rect 17320 17690 17330 17710
rect 17350 17690 17360 17710
rect 17320 17550 17360 17690
rect 17320 17530 17330 17550
rect 17350 17530 17360 17550
rect 17320 17390 17360 17530
rect 17320 17370 17330 17390
rect 17350 17370 17360 17390
rect 17320 17230 17360 17370
rect 17320 17210 17330 17230
rect 17350 17210 17360 17230
rect 17320 17200 17360 17210
rect 17400 18190 17440 18200
rect 17400 18170 17410 18190
rect 17430 18170 17440 18190
rect 17400 18030 17440 18170
rect 17400 18010 17410 18030
rect 17430 18010 17440 18030
rect 17400 17870 17440 18010
rect 17400 17850 17410 17870
rect 17430 17850 17440 17870
rect 17400 17710 17440 17850
rect 17400 17690 17410 17710
rect 17430 17690 17440 17710
rect 17400 17550 17440 17690
rect 17400 17530 17410 17550
rect 17430 17530 17440 17550
rect 17400 17390 17440 17530
rect 17400 17370 17410 17390
rect 17430 17370 17440 17390
rect 17400 17230 17440 17370
rect 17400 17210 17410 17230
rect 17430 17210 17440 17230
rect 17400 17200 17440 17210
rect 17480 18190 17520 18200
rect 17480 18170 17490 18190
rect 17510 18170 17520 18190
rect 17480 18030 17520 18170
rect 17480 18010 17490 18030
rect 17510 18010 17520 18030
rect 17480 17870 17520 18010
rect 17480 17850 17490 17870
rect 17510 17850 17520 17870
rect 17480 17710 17520 17850
rect 17480 17690 17490 17710
rect 17510 17690 17520 17710
rect 17480 17550 17520 17690
rect 17480 17530 17490 17550
rect 17510 17530 17520 17550
rect 17480 17390 17520 17530
rect 17480 17370 17490 17390
rect 17510 17370 17520 17390
rect 17480 17230 17520 17370
rect 17480 17210 17490 17230
rect 17510 17210 17520 17230
rect 17480 17200 17520 17210
rect 17560 18190 17600 18200
rect 17560 18170 17570 18190
rect 17590 18170 17600 18190
rect 17560 18030 17600 18170
rect 17560 18010 17570 18030
rect 17590 18010 17600 18030
rect 17560 17870 17600 18010
rect 17560 17850 17570 17870
rect 17590 17850 17600 17870
rect 17560 17710 17600 17850
rect 17560 17690 17570 17710
rect 17590 17690 17600 17710
rect 17560 17550 17600 17690
rect 17560 17530 17570 17550
rect 17590 17530 17600 17550
rect 17560 17390 17600 17530
rect 17560 17370 17570 17390
rect 17590 17370 17600 17390
rect 17560 17230 17600 17370
rect 17560 17210 17570 17230
rect 17590 17210 17600 17230
rect 17560 17200 17600 17210
rect 17640 18190 17680 18200
rect 17640 18170 17650 18190
rect 17670 18170 17680 18190
rect 17640 18030 17680 18170
rect 17640 18010 17650 18030
rect 17670 18010 17680 18030
rect 17640 17870 17680 18010
rect 17640 17850 17650 17870
rect 17670 17850 17680 17870
rect 17640 17710 17680 17850
rect 17640 17690 17650 17710
rect 17670 17690 17680 17710
rect 17640 17550 17680 17690
rect 17640 17530 17650 17550
rect 17670 17530 17680 17550
rect 17640 17390 17680 17530
rect 17640 17370 17650 17390
rect 17670 17370 17680 17390
rect 17640 17230 17680 17370
rect 17640 17210 17650 17230
rect 17670 17210 17680 17230
rect 17640 17200 17680 17210
rect 17720 18190 17760 18200
rect 17720 18170 17730 18190
rect 17750 18170 17760 18190
rect 17720 18030 17760 18170
rect 17720 18010 17730 18030
rect 17750 18010 17760 18030
rect 17720 17870 17760 18010
rect 17720 17850 17730 17870
rect 17750 17850 17760 17870
rect 17720 17710 17760 17850
rect 17720 17690 17730 17710
rect 17750 17690 17760 17710
rect 17720 17550 17760 17690
rect 17720 17530 17730 17550
rect 17750 17530 17760 17550
rect 17720 17390 17760 17530
rect 17720 17370 17730 17390
rect 17750 17370 17760 17390
rect 17720 17230 17760 17370
rect 17720 17210 17730 17230
rect 17750 17210 17760 17230
rect 17720 17200 17760 17210
rect 17800 18190 17840 18200
rect 17800 18170 17810 18190
rect 17830 18170 17840 18190
rect 17800 18030 17840 18170
rect 17800 18010 17810 18030
rect 17830 18010 17840 18030
rect 17800 17870 17840 18010
rect 17800 17850 17810 17870
rect 17830 17850 17840 17870
rect 17800 17710 17840 17850
rect 17800 17690 17810 17710
rect 17830 17690 17840 17710
rect 17800 17550 17840 17690
rect 17800 17530 17810 17550
rect 17830 17530 17840 17550
rect 17800 17390 17840 17530
rect 17800 17370 17810 17390
rect 17830 17370 17840 17390
rect 17800 17230 17840 17370
rect 17800 17210 17810 17230
rect 17830 17210 17840 17230
rect 17800 17200 17840 17210
rect 17880 18190 17920 18200
rect 17880 18170 17890 18190
rect 17910 18170 17920 18190
rect 17880 18030 17920 18170
rect 17880 18010 17890 18030
rect 17910 18010 17920 18030
rect 17880 17870 17920 18010
rect 17880 17850 17890 17870
rect 17910 17850 17920 17870
rect 17880 17710 17920 17850
rect 17880 17690 17890 17710
rect 17910 17690 17920 17710
rect 17880 17550 17920 17690
rect 17880 17530 17890 17550
rect 17910 17530 17920 17550
rect 17880 17390 17920 17530
rect 17880 17370 17890 17390
rect 17910 17370 17920 17390
rect 17880 17230 17920 17370
rect 17880 17210 17890 17230
rect 17910 17210 17920 17230
rect 17880 17200 17920 17210
rect 17960 18190 18000 18200
rect 17960 18170 17970 18190
rect 17990 18170 18000 18190
rect 17960 18030 18000 18170
rect 17960 18010 17970 18030
rect 17990 18010 18000 18030
rect 17960 17870 18000 18010
rect 17960 17850 17970 17870
rect 17990 17850 18000 17870
rect 17960 17710 18000 17850
rect 17960 17690 17970 17710
rect 17990 17690 18000 17710
rect 17960 17550 18000 17690
rect 17960 17530 17970 17550
rect 17990 17530 18000 17550
rect 17960 17390 18000 17530
rect 17960 17370 17970 17390
rect 17990 17370 18000 17390
rect 17960 17230 18000 17370
rect 17960 17210 17970 17230
rect 17990 17210 18000 17230
rect 17960 17200 18000 17210
rect 18040 18190 18080 18200
rect 18040 18170 18050 18190
rect 18070 18170 18080 18190
rect 18040 18030 18080 18170
rect 18040 18010 18050 18030
rect 18070 18010 18080 18030
rect 18040 17870 18080 18010
rect 18040 17850 18050 17870
rect 18070 17850 18080 17870
rect 18040 17710 18080 17850
rect 18040 17690 18050 17710
rect 18070 17690 18080 17710
rect 18040 17550 18080 17690
rect 18040 17530 18050 17550
rect 18070 17530 18080 17550
rect 18040 17390 18080 17530
rect 18040 17370 18050 17390
rect 18070 17370 18080 17390
rect 18040 17230 18080 17370
rect 18040 17210 18050 17230
rect 18070 17210 18080 17230
rect 18040 17200 18080 17210
rect 18120 18190 18160 18200
rect 18120 18170 18130 18190
rect 18150 18170 18160 18190
rect 18120 18030 18160 18170
rect 18120 18010 18130 18030
rect 18150 18010 18160 18030
rect 18120 17870 18160 18010
rect 18120 17850 18130 17870
rect 18150 17850 18160 17870
rect 18120 17710 18160 17850
rect 18120 17690 18130 17710
rect 18150 17690 18160 17710
rect 18120 17550 18160 17690
rect 18120 17530 18130 17550
rect 18150 17530 18160 17550
rect 18120 17390 18160 17530
rect 18120 17370 18130 17390
rect 18150 17370 18160 17390
rect 18120 17230 18160 17370
rect 18120 17210 18130 17230
rect 18150 17210 18160 17230
rect 18120 17200 18160 17210
rect 18200 18190 18240 18200
rect 18200 18170 18210 18190
rect 18230 18170 18240 18190
rect 18200 18030 18240 18170
rect 18200 18010 18210 18030
rect 18230 18010 18240 18030
rect 18200 17870 18240 18010
rect 18200 17850 18210 17870
rect 18230 17850 18240 17870
rect 18200 17710 18240 17850
rect 18200 17690 18210 17710
rect 18230 17690 18240 17710
rect 18200 17550 18240 17690
rect 18200 17530 18210 17550
rect 18230 17530 18240 17550
rect 18200 17390 18240 17530
rect 18200 17370 18210 17390
rect 18230 17370 18240 17390
rect 18200 17230 18240 17370
rect 18200 17210 18210 17230
rect 18230 17210 18240 17230
rect 18200 17200 18240 17210
rect 18280 18190 18320 18200
rect 18280 18170 18290 18190
rect 18310 18170 18320 18190
rect 18280 18030 18320 18170
rect 18280 18010 18290 18030
rect 18310 18010 18320 18030
rect 18280 17870 18320 18010
rect 18280 17850 18290 17870
rect 18310 17850 18320 17870
rect 18280 17710 18320 17850
rect 18280 17690 18290 17710
rect 18310 17690 18320 17710
rect 18280 17550 18320 17690
rect 18280 17530 18290 17550
rect 18310 17530 18320 17550
rect 18280 17390 18320 17530
rect 18280 17370 18290 17390
rect 18310 17370 18320 17390
rect 18280 17230 18320 17370
rect 18280 17210 18290 17230
rect 18310 17210 18320 17230
rect 18280 17200 18320 17210
rect 18360 18190 18400 18200
rect 18360 18170 18370 18190
rect 18390 18170 18400 18190
rect 18360 18030 18400 18170
rect 18360 18010 18370 18030
rect 18390 18010 18400 18030
rect 18360 17870 18400 18010
rect 18360 17850 18370 17870
rect 18390 17850 18400 17870
rect 18360 17710 18400 17850
rect 18360 17690 18370 17710
rect 18390 17690 18400 17710
rect 18360 17550 18400 17690
rect 18360 17530 18370 17550
rect 18390 17530 18400 17550
rect 18360 17390 18400 17530
rect 18360 17370 18370 17390
rect 18390 17370 18400 17390
rect 18360 17230 18400 17370
rect 18360 17210 18370 17230
rect 18390 17210 18400 17230
rect 18360 17200 18400 17210
rect 18440 18190 18480 18200
rect 18440 18170 18450 18190
rect 18470 18170 18480 18190
rect 18440 18030 18480 18170
rect 18440 18010 18450 18030
rect 18470 18010 18480 18030
rect 18440 17870 18480 18010
rect 18440 17850 18450 17870
rect 18470 17850 18480 17870
rect 18440 17710 18480 17850
rect 18440 17690 18450 17710
rect 18470 17690 18480 17710
rect 18440 17550 18480 17690
rect 18440 17530 18450 17550
rect 18470 17530 18480 17550
rect 18440 17390 18480 17530
rect 18440 17370 18450 17390
rect 18470 17370 18480 17390
rect 18440 17230 18480 17370
rect 18440 17210 18450 17230
rect 18470 17210 18480 17230
rect 18440 17200 18480 17210
rect 18520 18190 18560 18200
rect 18520 18170 18530 18190
rect 18550 18170 18560 18190
rect 18520 18030 18560 18170
rect 18520 18010 18530 18030
rect 18550 18010 18560 18030
rect 18520 17870 18560 18010
rect 18520 17850 18530 17870
rect 18550 17850 18560 17870
rect 18520 17710 18560 17850
rect 18520 17690 18530 17710
rect 18550 17690 18560 17710
rect 18520 17550 18560 17690
rect 18520 17530 18530 17550
rect 18550 17530 18560 17550
rect 18520 17390 18560 17530
rect 18520 17370 18530 17390
rect 18550 17370 18560 17390
rect 18520 17230 18560 17370
rect 18520 17210 18530 17230
rect 18550 17210 18560 17230
rect 18520 17200 18560 17210
rect 18600 18190 18640 18200
rect 18600 18170 18610 18190
rect 18630 18170 18640 18190
rect 18600 18030 18640 18170
rect 18600 18010 18610 18030
rect 18630 18010 18640 18030
rect 18600 17870 18640 18010
rect 18600 17850 18610 17870
rect 18630 17850 18640 17870
rect 18600 17710 18640 17850
rect 18600 17690 18610 17710
rect 18630 17690 18640 17710
rect 18600 17550 18640 17690
rect 18600 17530 18610 17550
rect 18630 17530 18640 17550
rect 18600 17390 18640 17530
rect 18600 17370 18610 17390
rect 18630 17370 18640 17390
rect 18600 17230 18640 17370
rect 18600 17210 18610 17230
rect 18630 17210 18640 17230
rect 18600 17200 18640 17210
rect 18680 18190 18720 18200
rect 18680 18170 18690 18190
rect 18710 18170 18720 18190
rect 18680 18030 18720 18170
rect 18680 18010 18690 18030
rect 18710 18010 18720 18030
rect 18680 17870 18720 18010
rect 18680 17850 18690 17870
rect 18710 17850 18720 17870
rect 18680 17710 18720 17850
rect 18680 17690 18690 17710
rect 18710 17690 18720 17710
rect 18680 17550 18720 17690
rect 18680 17530 18690 17550
rect 18710 17530 18720 17550
rect 18680 17390 18720 17530
rect 18680 17370 18690 17390
rect 18710 17370 18720 17390
rect 18680 17230 18720 17370
rect 18680 17210 18690 17230
rect 18710 17210 18720 17230
rect 18680 17200 18720 17210
rect 18760 18190 18800 18200
rect 18760 18170 18770 18190
rect 18790 18170 18800 18190
rect 18760 18030 18800 18170
rect 18760 18010 18770 18030
rect 18790 18010 18800 18030
rect 18760 17870 18800 18010
rect 18760 17850 18770 17870
rect 18790 17850 18800 17870
rect 18760 17710 18800 17850
rect 18760 17690 18770 17710
rect 18790 17690 18800 17710
rect 18760 17550 18800 17690
rect 18760 17530 18770 17550
rect 18790 17530 18800 17550
rect 18760 17390 18800 17530
rect 18760 17370 18770 17390
rect 18790 17370 18800 17390
rect 18760 17230 18800 17370
rect 18760 17210 18770 17230
rect 18790 17210 18800 17230
rect 18760 17200 18800 17210
rect 18840 18190 18880 18200
rect 18840 18170 18850 18190
rect 18870 18170 18880 18190
rect 18840 18030 18880 18170
rect 18840 18010 18850 18030
rect 18870 18010 18880 18030
rect 18840 17870 18880 18010
rect 18840 17850 18850 17870
rect 18870 17850 18880 17870
rect 18840 17710 18880 17850
rect 18840 17690 18850 17710
rect 18870 17690 18880 17710
rect 18840 17550 18880 17690
rect 18840 17530 18850 17550
rect 18870 17530 18880 17550
rect 18840 17390 18880 17530
rect 18840 17370 18850 17390
rect 18870 17370 18880 17390
rect 18840 17230 18880 17370
rect 18840 17210 18850 17230
rect 18870 17210 18880 17230
rect 18840 17200 18880 17210
rect 18920 18190 18960 18200
rect 18920 18170 18930 18190
rect 18950 18170 18960 18190
rect 18920 18030 18960 18170
rect 18920 18010 18930 18030
rect 18950 18010 18960 18030
rect 18920 17870 18960 18010
rect 18920 17850 18930 17870
rect 18950 17850 18960 17870
rect 18920 17710 18960 17850
rect 18920 17690 18930 17710
rect 18950 17690 18960 17710
rect 18920 17550 18960 17690
rect 18920 17530 18930 17550
rect 18950 17530 18960 17550
rect 18920 17390 18960 17530
rect 18920 17370 18930 17390
rect 18950 17370 18960 17390
rect 18920 17230 18960 17370
rect 18920 17210 18930 17230
rect 18950 17210 18960 17230
rect 18920 17200 18960 17210
rect 19000 18190 19040 18200
rect 19000 18170 19010 18190
rect 19030 18170 19040 18190
rect 19000 18030 19040 18170
rect 19000 18010 19010 18030
rect 19030 18010 19040 18030
rect 19000 17870 19040 18010
rect 19000 17850 19010 17870
rect 19030 17850 19040 17870
rect 19000 17710 19040 17850
rect 19000 17690 19010 17710
rect 19030 17690 19040 17710
rect 19000 17550 19040 17690
rect 19000 17530 19010 17550
rect 19030 17530 19040 17550
rect 19000 17390 19040 17530
rect 19000 17370 19010 17390
rect 19030 17370 19040 17390
rect 19000 17230 19040 17370
rect 19000 17210 19010 17230
rect 19030 17210 19040 17230
rect 19000 17200 19040 17210
rect 19080 18190 19120 18200
rect 19080 18170 19090 18190
rect 19110 18170 19120 18190
rect 19080 18030 19120 18170
rect 19080 18010 19090 18030
rect 19110 18010 19120 18030
rect 19080 17870 19120 18010
rect 19080 17850 19090 17870
rect 19110 17850 19120 17870
rect 19080 17710 19120 17850
rect 19080 17690 19090 17710
rect 19110 17690 19120 17710
rect 19080 17550 19120 17690
rect 19080 17530 19090 17550
rect 19110 17530 19120 17550
rect 19080 17390 19120 17530
rect 19080 17370 19090 17390
rect 19110 17370 19120 17390
rect 19080 17230 19120 17370
rect 19080 17210 19090 17230
rect 19110 17210 19120 17230
rect 19080 17200 19120 17210
rect 19160 18190 19200 18200
rect 19160 18170 19170 18190
rect 19190 18170 19200 18190
rect 19160 18030 19200 18170
rect 19160 18010 19170 18030
rect 19190 18010 19200 18030
rect 19160 17870 19200 18010
rect 19160 17850 19170 17870
rect 19190 17850 19200 17870
rect 19160 17710 19200 17850
rect 19160 17690 19170 17710
rect 19190 17690 19200 17710
rect 19160 17550 19200 17690
rect 19160 17530 19170 17550
rect 19190 17530 19200 17550
rect 19160 17390 19200 17530
rect 19160 17370 19170 17390
rect 19190 17370 19200 17390
rect 19160 17230 19200 17370
rect 19160 17210 19170 17230
rect 19190 17210 19200 17230
rect 19160 17200 19200 17210
rect 19240 18190 19280 18200
rect 19240 18170 19250 18190
rect 19270 18170 19280 18190
rect 19240 18030 19280 18170
rect 19240 18010 19250 18030
rect 19270 18010 19280 18030
rect 19240 17870 19280 18010
rect 19240 17850 19250 17870
rect 19270 17850 19280 17870
rect 19240 17710 19280 17850
rect 19240 17690 19250 17710
rect 19270 17690 19280 17710
rect 19240 17550 19280 17690
rect 19240 17530 19250 17550
rect 19270 17530 19280 17550
rect 19240 17390 19280 17530
rect 19240 17370 19250 17390
rect 19270 17370 19280 17390
rect 19240 17230 19280 17370
rect 19240 17210 19250 17230
rect 19270 17210 19280 17230
rect 19240 17200 19280 17210
rect 19320 18190 19360 18200
rect 19320 18170 19330 18190
rect 19350 18170 19360 18190
rect 19320 18030 19360 18170
rect 19320 18010 19330 18030
rect 19350 18010 19360 18030
rect 19320 17870 19360 18010
rect 19320 17850 19330 17870
rect 19350 17850 19360 17870
rect 19320 17710 19360 17850
rect 19320 17690 19330 17710
rect 19350 17690 19360 17710
rect 19320 17550 19360 17690
rect 19320 17530 19330 17550
rect 19350 17530 19360 17550
rect 19320 17390 19360 17530
rect 19320 17370 19330 17390
rect 19350 17370 19360 17390
rect 19320 17230 19360 17370
rect 19320 17210 19330 17230
rect 19350 17210 19360 17230
rect 19320 17200 19360 17210
rect 19400 18190 19440 18200
rect 19400 18170 19410 18190
rect 19430 18170 19440 18190
rect 19400 18030 19440 18170
rect 19400 18010 19410 18030
rect 19430 18010 19440 18030
rect 19400 17870 19440 18010
rect 19400 17850 19410 17870
rect 19430 17850 19440 17870
rect 19400 17710 19440 17850
rect 19400 17690 19410 17710
rect 19430 17690 19440 17710
rect 19400 17550 19440 17690
rect 19400 17530 19410 17550
rect 19430 17530 19440 17550
rect 19400 17390 19440 17530
rect 19400 17370 19410 17390
rect 19430 17370 19440 17390
rect 19400 17230 19440 17370
rect 19400 17210 19410 17230
rect 19430 17210 19440 17230
rect 19400 17200 19440 17210
rect 19480 18190 19520 18200
rect 19480 18170 19490 18190
rect 19510 18170 19520 18190
rect 19480 18030 19520 18170
rect 19480 18010 19490 18030
rect 19510 18010 19520 18030
rect 19480 17870 19520 18010
rect 19480 17850 19490 17870
rect 19510 17850 19520 17870
rect 19480 17710 19520 17850
rect 19480 17690 19490 17710
rect 19510 17690 19520 17710
rect 19480 17550 19520 17690
rect 19480 17530 19490 17550
rect 19510 17530 19520 17550
rect 19480 17390 19520 17530
rect 19480 17370 19490 17390
rect 19510 17370 19520 17390
rect 19480 17230 19520 17370
rect 19480 17210 19490 17230
rect 19510 17210 19520 17230
rect 19480 17200 19520 17210
rect 19560 18190 19600 18200
rect 19560 18170 19570 18190
rect 19590 18170 19600 18190
rect 19560 18030 19600 18170
rect 19560 18010 19570 18030
rect 19590 18010 19600 18030
rect 19560 17870 19600 18010
rect 19560 17850 19570 17870
rect 19590 17850 19600 17870
rect 19560 17710 19600 17850
rect 19560 17690 19570 17710
rect 19590 17690 19600 17710
rect 19560 17550 19600 17690
rect 19560 17530 19570 17550
rect 19590 17530 19600 17550
rect 19560 17390 19600 17530
rect 19560 17370 19570 17390
rect 19590 17370 19600 17390
rect 19560 17230 19600 17370
rect 19560 17210 19570 17230
rect 19590 17210 19600 17230
rect 19560 17200 19600 17210
rect 19640 18190 19680 18200
rect 19640 18170 19650 18190
rect 19670 18170 19680 18190
rect 19640 18030 19680 18170
rect 19640 18010 19650 18030
rect 19670 18010 19680 18030
rect 19640 17870 19680 18010
rect 19640 17850 19650 17870
rect 19670 17850 19680 17870
rect 19640 17710 19680 17850
rect 19640 17690 19650 17710
rect 19670 17690 19680 17710
rect 19640 17550 19680 17690
rect 19640 17530 19650 17550
rect 19670 17530 19680 17550
rect 19640 17390 19680 17530
rect 19640 17370 19650 17390
rect 19670 17370 19680 17390
rect 19640 17230 19680 17370
rect 19640 17210 19650 17230
rect 19670 17210 19680 17230
rect 19640 17200 19680 17210
rect 19720 18190 19760 18200
rect 19720 18170 19730 18190
rect 19750 18170 19760 18190
rect 19720 18030 19760 18170
rect 19720 18010 19730 18030
rect 19750 18010 19760 18030
rect 19720 17870 19760 18010
rect 19720 17850 19730 17870
rect 19750 17850 19760 17870
rect 19720 17710 19760 17850
rect 19720 17690 19730 17710
rect 19750 17690 19760 17710
rect 19720 17550 19760 17690
rect 19720 17530 19730 17550
rect 19750 17530 19760 17550
rect 19720 17390 19760 17530
rect 19720 17370 19730 17390
rect 19750 17370 19760 17390
rect 19720 17230 19760 17370
rect 19720 17210 19730 17230
rect 19750 17210 19760 17230
rect 19720 17200 19760 17210
rect 19800 18190 19840 18200
rect 19800 18170 19810 18190
rect 19830 18170 19840 18190
rect 19800 18030 19840 18170
rect 19800 18010 19810 18030
rect 19830 18010 19840 18030
rect 19800 17870 19840 18010
rect 19800 17850 19810 17870
rect 19830 17850 19840 17870
rect 19800 17710 19840 17850
rect 19800 17690 19810 17710
rect 19830 17690 19840 17710
rect 19800 17550 19840 17690
rect 19800 17530 19810 17550
rect 19830 17530 19840 17550
rect 19800 17390 19840 17530
rect 19800 17370 19810 17390
rect 19830 17370 19840 17390
rect 19800 17230 19840 17370
rect 19800 17210 19810 17230
rect 19830 17210 19840 17230
rect 19800 17200 19840 17210
rect 19880 18190 19920 18200
rect 19880 18170 19890 18190
rect 19910 18170 19920 18190
rect 19880 18030 19920 18170
rect 19880 18010 19890 18030
rect 19910 18010 19920 18030
rect 19880 17870 19920 18010
rect 19880 17850 19890 17870
rect 19910 17850 19920 17870
rect 19880 17710 19920 17850
rect 19880 17690 19890 17710
rect 19910 17690 19920 17710
rect 19880 17550 19920 17690
rect 19880 17530 19890 17550
rect 19910 17530 19920 17550
rect 19880 17390 19920 17530
rect 19880 17370 19890 17390
rect 19910 17370 19920 17390
rect 19880 17230 19920 17370
rect 19880 17210 19890 17230
rect 19910 17210 19920 17230
rect 19880 17200 19920 17210
rect 19960 18190 20000 18200
rect 19960 18170 19970 18190
rect 19990 18170 20000 18190
rect 19960 18030 20000 18170
rect 19960 18010 19970 18030
rect 19990 18010 20000 18030
rect 19960 17870 20000 18010
rect 19960 17850 19970 17870
rect 19990 17850 20000 17870
rect 19960 17710 20000 17850
rect 19960 17690 19970 17710
rect 19990 17690 20000 17710
rect 19960 17550 20000 17690
rect 19960 17530 19970 17550
rect 19990 17530 20000 17550
rect 19960 17390 20000 17530
rect 19960 17370 19970 17390
rect 19990 17370 20000 17390
rect 19960 17230 20000 17370
rect 19960 17210 19970 17230
rect 19990 17210 20000 17230
rect 19960 17200 20000 17210
rect 20040 18190 20080 18200
rect 20040 18170 20050 18190
rect 20070 18170 20080 18190
rect 20040 18030 20080 18170
rect 20040 18010 20050 18030
rect 20070 18010 20080 18030
rect 20040 17870 20080 18010
rect 20040 17850 20050 17870
rect 20070 17850 20080 17870
rect 20040 17710 20080 17850
rect 20040 17690 20050 17710
rect 20070 17690 20080 17710
rect 20040 17550 20080 17690
rect 20040 17530 20050 17550
rect 20070 17530 20080 17550
rect 20040 17390 20080 17530
rect 20040 17370 20050 17390
rect 20070 17370 20080 17390
rect 20040 17230 20080 17370
rect 20040 17210 20050 17230
rect 20070 17210 20080 17230
rect 20040 17200 20080 17210
rect 20120 18190 20160 18200
rect 20120 18170 20130 18190
rect 20150 18170 20160 18190
rect 20120 18030 20160 18170
rect 20120 18010 20130 18030
rect 20150 18010 20160 18030
rect 20120 17870 20160 18010
rect 20120 17850 20130 17870
rect 20150 17850 20160 17870
rect 20120 17710 20160 17850
rect 20120 17690 20130 17710
rect 20150 17690 20160 17710
rect 20120 17550 20160 17690
rect 20120 17530 20130 17550
rect 20150 17530 20160 17550
rect 20120 17390 20160 17530
rect 20120 17370 20130 17390
rect 20150 17370 20160 17390
rect 20120 17230 20160 17370
rect 20120 17210 20130 17230
rect 20150 17210 20160 17230
rect 20120 17200 20160 17210
rect 20200 18190 20240 18200
rect 20200 18170 20210 18190
rect 20230 18170 20240 18190
rect 20200 18030 20240 18170
rect 20200 18010 20210 18030
rect 20230 18010 20240 18030
rect 20200 17870 20240 18010
rect 20200 17850 20210 17870
rect 20230 17850 20240 17870
rect 20200 17710 20240 17850
rect 20200 17690 20210 17710
rect 20230 17690 20240 17710
rect 20200 17550 20240 17690
rect 20200 17530 20210 17550
rect 20230 17530 20240 17550
rect 20200 17390 20240 17530
rect 20200 17370 20210 17390
rect 20230 17370 20240 17390
rect 20200 17230 20240 17370
rect 20200 17210 20210 17230
rect 20230 17210 20240 17230
rect 20200 17200 20240 17210
rect 20280 18190 20320 18200
rect 20280 18170 20290 18190
rect 20310 18170 20320 18190
rect 20280 18030 20320 18170
rect 20280 18010 20290 18030
rect 20310 18010 20320 18030
rect 20280 17870 20320 18010
rect 20280 17850 20290 17870
rect 20310 17850 20320 17870
rect 20280 17710 20320 17850
rect 20280 17690 20290 17710
rect 20310 17690 20320 17710
rect 20280 17550 20320 17690
rect 20280 17530 20290 17550
rect 20310 17530 20320 17550
rect 20280 17390 20320 17530
rect 20280 17370 20290 17390
rect 20310 17370 20320 17390
rect 20280 17230 20320 17370
rect 20280 17210 20290 17230
rect 20310 17210 20320 17230
rect 20280 17200 20320 17210
rect 20360 18190 20400 18200
rect 20360 18170 20370 18190
rect 20390 18170 20400 18190
rect 20360 18030 20400 18170
rect 20360 18010 20370 18030
rect 20390 18010 20400 18030
rect 20360 17870 20400 18010
rect 20360 17850 20370 17870
rect 20390 17850 20400 17870
rect 20360 17710 20400 17850
rect 20360 17690 20370 17710
rect 20390 17690 20400 17710
rect 20360 17550 20400 17690
rect 20360 17530 20370 17550
rect 20390 17530 20400 17550
rect 20360 17390 20400 17530
rect 20360 17370 20370 17390
rect 20390 17370 20400 17390
rect 20360 17230 20400 17370
rect 20360 17210 20370 17230
rect 20390 17210 20400 17230
rect 20360 17200 20400 17210
rect 20440 18190 20480 18200
rect 20440 18170 20450 18190
rect 20470 18170 20480 18190
rect 20440 18030 20480 18170
rect 20440 18010 20450 18030
rect 20470 18010 20480 18030
rect 20440 17870 20480 18010
rect 20440 17850 20450 17870
rect 20470 17850 20480 17870
rect 20440 17710 20480 17850
rect 20440 17690 20450 17710
rect 20470 17690 20480 17710
rect 20440 17550 20480 17690
rect 20440 17530 20450 17550
rect 20470 17530 20480 17550
rect 20440 17390 20480 17530
rect 20440 17370 20450 17390
rect 20470 17370 20480 17390
rect 20440 17230 20480 17370
rect 20440 17210 20450 17230
rect 20470 17210 20480 17230
rect 20440 17200 20480 17210
rect 20520 18190 20560 18200
rect 20520 18170 20530 18190
rect 20550 18170 20560 18190
rect 20520 18030 20560 18170
rect 20520 18010 20530 18030
rect 20550 18010 20560 18030
rect 20520 17870 20560 18010
rect 20520 17850 20530 17870
rect 20550 17850 20560 17870
rect 20520 17710 20560 17850
rect 20520 17690 20530 17710
rect 20550 17690 20560 17710
rect 20520 17550 20560 17690
rect 20520 17530 20530 17550
rect 20550 17530 20560 17550
rect 20520 17390 20560 17530
rect 20520 17370 20530 17390
rect 20550 17370 20560 17390
rect 20520 17230 20560 17370
rect 20520 17210 20530 17230
rect 20550 17210 20560 17230
rect 20520 17200 20560 17210
rect 20600 18190 20640 18200
rect 20600 18170 20610 18190
rect 20630 18170 20640 18190
rect 20600 18030 20640 18170
rect 20600 18010 20610 18030
rect 20630 18010 20640 18030
rect 20600 17870 20640 18010
rect 20600 17850 20610 17870
rect 20630 17850 20640 17870
rect 20600 17710 20640 17850
rect 20600 17690 20610 17710
rect 20630 17690 20640 17710
rect 20600 17550 20640 17690
rect 20600 17530 20610 17550
rect 20630 17530 20640 17550
rect 20600 17390 20640 17530
rect 20600 17370 20610 17390
rect 20630 17370 20640 17390
rect 20600 17230 20640 17370
rect 20600 17210 20610 17230
rect 20630 17210 20640 17230
rect 20600 17200 20640 17210
rect 20680 18190 20720 18200
rect 20680 18170 20690 18190
rect 20710 18170 20720 18190
rect 20680 18030 20720 18170
rect 20680 18010 20690 18030
rect 20710 18010 20720 18030
rect 20680 17870 20720 18010
rect 20680 17850 20690 17870
rect 20710 17850 20720 17870
rect 20680 17710 20720 17850
rect 20680 17690 20690 17710
rect 20710 17690 20720 17710
rect 20680 17550 20720 17690
rect 20680 17530 20690 17550
rect 20710 17530 20720 17550
rect 20680 17390 20720 17530
rect 20680 17370 20690 17390
rect 20710 17370 20720 17390
rect 20680 17230 20720 17370
rect 20680 17210 20690 17230
rect 20710 17210 20720 17230
rect 20680 17200 20720 17210
rect 20760 18190 20800 18200
rect 20760 18170 20770 18190
rect 20790 18170 20800 18190
rect 20760 18030 20800 18170
rect 20760 18010 20770 18030
rect 20790 18010 20800 18030
rect 20760 17870 20800 18010
rect 20760 17850 20770 17870
rect 20790 17850 20800 17870
rect 20760 17710 20800 17850
rect 20760 17690 20770 17710
rect 20790 17690 20800 17710
rect 20760 17550 20800 17690
rect 20760 17530 20770 17550
rect 20790 17530 20800 17550
rect 20760 17390 20800 17530
rect 20760 17370 20770 17390
rect 20790 17370 20800 17390
rect 20760 17230 20800 17370
rect 20760 17210 20770 17230
rect 20790 17210 20800 17230
rect 20760 17200 20800 17210
rect 20840 18190 20880 18200
rect 20840 18170 20850 18190
rect 20870 18170 20880 18190
rect 20840 18030 20880 18170
rect 20840 18010 20850 18030
rect 20870 18010 20880 18030
rect 20840 17870 20880 18010
rect 20840 17850 20850 17870
rect 20870 17850 20880 17870
rect 20840 17710 20880 17850
rect 20840 17690 20850 17710
rect 20870 17690 20880 17710
rect 20840 17550 20880 17690
rect 20840 17530 20850 17550
rect 20870 17530 20880 17550
rect 20840 17390 20880 17530
rect 20840 17370 20850 17390
rect 20870 17370 20880 17390
rect 20840 17230 20880 17370
rect 20840 17210 20850 17230
rect 20870 17210 20880 17230
rect 20840 17200 20880 17210
rect 20920 18190 20960 18200
rect 20920 18170 20930 18190
rect 20950 18170 20960 18190
rect 20920 18030 20960 18170
rect 20920 18010 20930 18030
rect 20950 18010 20960 18030
rect 20920 17870 20960 18010
rect 20920 17850 20930 17870
rect 20950 17850 20960 17870
rect 20920 17710 20960 17850
rect 20920 17690 20930 17710
rect 20950 17690 20960 17710
rect 20920 17550 20960 17690
rect 20920 17530 20930 17550
rect 20950 17530 20960 17550
rect 20920 17390 20960 17530
rect 20920 17370 20930 17390
rect 20950 17370 20960 17390
rect 20920 17230 20960 17370
rect 20920 17210 20930 17230
rect 20950 17210 20960 17230
rect 20920 17200 20960 17210
rect 0 17150 40 17160
rect 0 17130 10 17150
rect 30 17130 40 17150
rect 0 16990 40 17130
rect 0 16970 10 16990
rect 30 16970 40 16990
rect 0 16960 40 16970
rect 80 17150 120 17160
rect 80 17130 90 17150
rect 110 17130 120 17150
rect 80 16990 120 17130
rect 80 16970 90 16990
rect 110 16970 120 16990
rect 80 16960 120 16970
rect 160 17150 200 17160
rect 160 17130 170 17150
rect 190 17130 200 17150
rect 160 16990 200 17130
rect 160 16970 170 16990
rect 190 16970 200 16990
rect 160 16960 200 16970
rect 240 17150 280 17160
rect 240 17130 250 17150
rect 270 17130 280 17150
rect 240 16990 280 17130
rect 240 16970 250 16990
rect 270 16970 280 16990
rect 240 16960 280 16970
rect 320 17150 360 17160
rect 320 17130 330 17150
rect 350 17130 360 17150
rect 320 16990 360 17130
rect 320 16970 330 16990
rect 350 16970 360 16990
rect 320 16960 360 16970
rect 400 17150 440 17160
rect 400 17130 410 17150
rect 430 17130 440 17150
rect 400 16990 440 17130
rect 400 16970 410 16990
rect 430 16970 440 16990
rect 400 16960 440 16970
rect 480 17150 520 17160
rect 480 17130 490 17150
rect 510 17130 520 17150
rect 480 16990 520 17130
rect 480 16970 490 16990
rect 510 16970 520 16990
rect 480 16960 520 16970
rect 560 17150 600 17160
rect 560 17130 570 17150
rect 590 17130 600 17150
rect 560 16990 600 17130
rect 560 16970 570 16990
rect 590 16970 600 16990
rect 560 16960 600 16970
rect 640 17150 680 17160
rect 640 17130 650 17150
rect 670 17130 680 17150
rect 640 16990 680 17130
rect 640 16970 650 16990
rect 670 16970 680 16990
rect 640 16960 680 16970
rect 720 17150 760 17160
rect 720 17130 730 17150
rect 750 17130 760 17150
rect 720 16990 760 17130
rect 720 16970 730 16990
rect 750 16970 760 16990
rect 720 16960 760 16970
rect 800 17150 840 17160
rect 800 17130 810 17150
rect 830 17130 840 17150
rect 800 16990 840 17130
rect 800 16970 810 16990
rect 830 16970 840 16990
rect 800 16960 840 16970
rect 880 17150 920 17160
rect 880 17130 890 17150
rect 910 17130 920 17150
rect 880 16990 920 17130
rect 880 16970 890 16990
rect 910 16970 920 16990
rect 880 16960 920 16970
rect 960 17150 1000 17160
rect 960 17130 970 17150
rect 990 17130 1000 17150
rect 960 16990 1000 17130
rect 960 16970 970 16990
rect 990 16970 1000 16990
rect 960 16960 1000 16970
rect 1040 17150 1080 17160
rect 1040 17130 1050 17150
rect 1070 17130 1080 17150
rect 1040 16990 1080 17130
rect 1040 16970 1050 16990
rect 1070 16970 1080 16990
rect 1040 16960 1080 16970
rect 1120 17150 1160 17160
rect 1120 17130 1130 17150
rect 1150 17130 1160 17150
rect 1120 16990 1160 17130
rect 1120 16970 1130 16990
rect 1150 16970 1160 16990
rect 1120 16960 1160 16970
rect 1200 17150 1240 17160
rect 1200 17130 1210 17150
rect 1230 17130 1240 17150
rect 1200 16990 1240 17130
rect 1200 16970 1210 16990
rect 1230 16970 1240 16990
rect 1200 16960 1240 16970
rect 1280 17150 1320 17160
rect 1280 17130 1290 17150
rect 1310 17130 1320 17150
rect 1280 16990 1320 17130
rect 1280 16970 1290 16990
rect 1310 16970 1320 16990
rect 1280 16960 1320 16970
rect 1360 17150 1400 17160
rect 1360 17130 1370 17150
rect 1390 17130 1400 17150
rect 1360 16990 1400 17130
rect 1360 16970 1370 16990
rect 1390 16970 1400 16990
rect 1360 16960 1400 16970
rect 1440 17150 1480 17160
rect 1440 17130 1450 17150
rect 1470 17130 1480 17150
rect 1440 16990 1480 17130
rect 1440 16970 1450 16990
rect 1470 16970 1480 16990
rect 1440 16960 1480 16970
rect 1520 17150 1560 17160
rect 1520 17130 1530 17150
rect 1550 17130 1560 17150
rect 1520 16990 1560 17130
rect 1520 16970 1530 16990
rect 1550 16970 1560 16990
rect 1520 16960 1560 16970
rect 1600 17150 1640 17160
rect 1600 17130 1610 17150
rect 1630 17130 1640 17150
rect 1600 16990 1640 17130
rect 1600 16970 1610 16990
rect 1630 16970 1640 16990
rect 1600 16960 1640 16970
rect 1680 17150 1720 17160
rect 1680 17130 1690 17150
rect 1710 17130 1720 17150
rect 1680 16990 1720 17130
rect 1680 16970 1690 16990
rect 1710 16970 1720 16990
rect 1680 16960 1720 16970
rect 1760 17150 1800 17160
rect 1760 17130 1770 17150
rect 1790 17130 1800 17150
rect 1760 16990 1800 17130
rect 1760 16970 1770 16990
rect 1790 16970 1800 16990
rect 1760 16960 1800 16970
rect 1840 17150 1880 17160
rect 1840 17130 1850 17150
rect 1870 17130 1880 17150
rect 1840 16990 1880 17130
rect 1840 16970 1850 16990
rect 1870 16970 1880 16990
rect 1840 16960 1880 16970
rect 1920 17150 1960 17160
rect 1920 17130 1930 17150
rect 1950 17130 1960 17150
rect 1920 16990 1960 17130
rect 1920 16970 1930 16990
rect 1950 16970 1960 16990
rect 1920 16960 1960 16970
rect 2000 17150 2040 17160
rect 2000 17130 2010 17150
rect 2030 17130 2040 17150
rect 2000 16990 2040 17130
rect 2000 16970 2010 16990
rect 2030 16970 2040 16990
rect 2000 16960 2040 16970
rect 2080 17150 2120 17160
rect 2080 17130 2090 17150
rect 2110 17130 2120 17150
rect 2080 16990 2120 17130
rect 2080 16970 2090 16990
rect 2110 16970 2120 16990
rect 2080 16960 2120 16970
rect 2160 17150 2200 17160
rect 2160 17130 2170 17150
rect 2190 17130 2200 17150
rect 2160 16990 2200 17130
rect 2160 16970 2170 16990
rect 2190 16970 2200 16990
rect 2160 16960 2200 16970
rect 2240 17150 2280 17160
rect 2240 17130 2250 17150
rect 2270 17130 2280 17150
rect 2240 16990 2280 17130
rect 2240 16970 2250 16990
rect 2270 16970 2280 16990
rect 2240 16960 2280 16970
rect 2320 17150 2360 17160
rect 2320 17130 2330 17150
rect 2350 17130 2360 17150
rect 2320 16990 2360 17130
rect 2320 16970 2330 16990
rect 2350 16970 2360 16990
rect 2320 16960 2360 16970
rect 2400 17150 2440 17160
rect 2400 17130 2410 17150
rect 2430 17130 2440 17150
rect 2400 16990 2440 17130
rect 2400 16970 2410 16990
rect 2430 16970 2440 16990
rect 2400 16960 2440 16970
rect 2480 17150 2520 17160
rect 2480 17130 2490 17150
rect 2510 17130 2520 17150
rect 2480 16990 2520 17130
rect 2480 16970 2490 16990
rect 2510 16970 2520 16990
rect 2480 16960 2520 16970
rect 2560 17150 2600 17160
rect 2560 17130 2570 17150
rect 2590 17130 2600 17150
rect 2560 16990 2600 17130
rect 2560 16970 2570 16990
rect 2590 16970 2600 16990
rect 2560 16960 2600 16970
rect 2640 17150 2680 17160
rect 2640 17130 2650 17150
rect 2670 17130 2680 17150
rect 2640 16990 2680 17130
rect 2640 16970 2650 16990
rect 2670 16970 2680 16990
rect 2640 16960 2680 16970
rect 2720 17150 2760 17160
rect 2720 17130 2730 17150
rect 2750 17130 2760 17150
rect 2720 16990 2760 17130
rect 2720 16970 2730 16990
rect 2750 16970 2760 16990
rect 2720 16960 2760 16970
rect 2800 17150 2840 17160
rect 2800 17130 2810 17150
rect 2830 17130 2840 17150
rect 2800 16990 2840 17130
rect 2800 16970 2810 16990
rect 2830 16970 2840 16990
rect 2800 16960 2840 16970
rect 2880 17150 2920 17160
rect 2880 17130 2890 17150
rect 2910 17130 2920 17150
rect 2880 16990 2920 17130
rect 2880 16970 2890 16990
rect 2910 16970 2920 16990
rect 2880 16960 2920 16970
rect 2960 17150 3000 17160
rect 2960 17130 2970 17150
rect 2990 17130 3000 17150
rect 2960 16990 3000 17130
rect 2960 16970 2970 16990
rect 2990 16970 3000 16990
rect 2960 16960 3000 16970
rect 3040 17150 3080 17160
rect 3040 17130 3050 17150
rect 3070 17130 3080 17150
rect 3040 16990 3080 17130
rect 3040 16970 3050 16990
rect 3070 16970 3080 16990
rect 3040 16960 3080 16970
rect 3120 17150 3160 17160
rect 3120 17130 3130 17150
rect 3150 17130 3160 17150
rect 3120 16990 3160 17130
rect 3120 16970 3130 16990
rect 3150 16970 3160 16990
rect 3120 16960 3160 16970
rect 3200 17150 3240 17160
rect 3200 17130 3210 17150
rect 3230 17130 3240 17150
rect 3200 16990 3240 17130
rect 3200 16970 3210 16990
rect 3230 16970 3240 16990
rect 3200 16960 3240 16970
rect 3280 17150 3320 17160
rect 3280 17130 3290 17150
rect 3310 17130 3320 17150
rect 3280 16990 3320 17130
rect 3280 16970 3290 16990
rect 3310 16970 3320 16990
rect 3280 16960 3320 16970
rect 3360 17150 3400 17160
rect 3360 17130 3370 17150
rect 3390 17130 3400 17150
rect 3360 16990 3400 17130
rect 3360 16970 3370 16990
rect 3390 16970 3400 16990
rect 3360 16960 3400 16970
rect 3440 17150 3480 17160
rect 3440 17130 3450 17150
rect 3470 17130 3480 17150
rect 3440 16990 3480 17130
rect 3440 16970 3450 16990
rect 3470 16970 3480 16990
rect 3440 16960 3480 16970
rect 3520 17150 3560 17160
rect 3520 17130 3530 17150
rect 3550 17130 3560 17150
rect 3520 16990 3560 17130
rect 3520 16970 3530 16990
rect 3550 16970 3560 16990
rect 3520 16960 3560 16970
rect 3600 17150 3640 17160
rect 3600 17130 3610 17150
rect 3630 17130 3640 17150
rect 3600 16990 3640 17130
rect 3600 16970 3610 16990
rect 3630 16970 3640 16990
rect 3600 16960 3640 16970
rect 3680 17150 3720 17160
rect 3680 17130 3690 17150
rect 3710 17130 3720 17150
rect 3680 16990 3720 17130
rect 3680 16970 3690 16990
rect 3710 16970 3720 16990
rect 3680 16960 3720 16970
rect 3760 17150 3800 17160
rect 3760 17130 3770 17150
rect 3790 17130 3800 17150
rect 3760 16990 3800 17130
rect 3760 16970 3770 16990
rect 3790 16970 3800 16990
rect 3760 16960 3800 16970
rect 3840 17150 3880 17160
rect 3840 17130 3850 17150
rect 3870 17130 3880 17150
rect 3840 16990 3880 17130
rect 3840 16970 3850 16990
rect 3870 16970 3880 16990
rect 3840 16960 3880 16970
rect 3920 17150 3960 17160
rect 3920 17130 3930 17150
rect 3950 17130 3960 17150
rect 3920 16990 3960 17130
rect 3920 16970 3930 16990
rect 3950 16970 3960 16990
rect 3920 16960 3960 16970
rect 4000 17150 4040 17160
rect 4000 17130 4010 17150
rect 4030 17130 4040 17150
rect 4000 16990 4040 17130
rect 4000 16970 4010 16990
rect 4030 16970 4040 16990
rect 4000 16960 4040 16970
rect 4080 17150 4120 17160
rect 4080 17130 4090 17150
rect 4110 17130 4120 17150
rect 4080 16990 4120 17130
rect 4080 16970 4090 16990
rect 4110 16970 4120 16990
rect 4080 16960 4120 16970
rect 4160 17150 4200 17160
rect 4160 17130 4170 17150
rect 4190 17130 4200 17150
rect 4160 16990 4200 17130
rect 4160 16970 4170 16990
rect 4190 16970 4200 16990
rect 4160 16960 4200 16970
rect 4240 16960 4280 17160
rect 4320 16960 4360 17160
rect 4400 16960 4440 17160
rect 4480 16960 4520 17160
rect 4560 16960 4600 17160
rect 4640 16960 4680 17160
rect 4720 16960 4760 17160
rect 4800 16960 4840 17160
rect 4880 16960 4920 17160
rect 4960 16960 5000 17160
rect 5040 16960 5080 17160
rect 5120 16960 5160 17160
rect 5200 16960 5240 17160
rect 5280 16960 5320 17160
rect 5360 16960 5400 17160
rect 5440 16960 5480 17160
rect 5520 16960 5560 17160
rect 5600 16960 5640 17160
rect 5680 16960 5720 17160
rect 5760 16960 5800 17160
rect 5840 16960 5880 17160
rect 5920 16960 5960 17160
rect 6000 16960 6040 17160
rect 6080 16960 6120 17160
rect 6160 16960 6200 17160
rect 6240 17150 6280 17160
rect 6240 17130 6250 17150
rect 6270 17130 6280 17150
rect 6240 16990 6280 17130
rect 6240 16970 6250 16990
rect 6270 16970 6280 16990
rect 6240 16960 6280 16970
rect 6320 17150 6360 17160
rect 6320 17130 6330 17150
rect 6350 17130 6360 17150
rect 6320 16990 6360 17130
rect 6320 16970 6330 16990
rect 6350 16970 6360 16990
rect 6320 16960 6360 16970
rect 6400 17150 6440 17160
rect 6400 17130 6410 17150
rect 6430 17130 6440 17150
rect 6400 16990 6440 17130
rect 6400 16970 6410 16990
rect 6430 16970 6440 16990
rect 6400 16960 6440 16970
rect 6480 17150 6520 17160
rect 6480 17130 6490 17150
rect 6510 17130 6520 17150
rect 6480 16990 6520 17130
rect 6480 16970 6490 16990
rect 6510 16970 6520 16990
rect 6480 16960 6520 16970
rect 6560 17150 6600 17160
rect 6560 17130 6570 17150
rect 6590 17130 6600 17150
rect 6560 16990 6600 17130
rect 6560 16970 6570 16990
rect 6590 16970 6600 16990
rect 6560 16960 6600 16970
rect 6640 17150 6680 17160
rect 6640 17130 6650 17150
rect 6670 17130 6680 17150
rect 6640 16990 6680 17130
rect 6640 16970 6650 16990
rect 6670 16970 6680 16990
rect 6640 16960 6680 16970
rect 6720 17150 6760 17160
rect 6720 17130 6730 17150
rect 6750 17130 6760 17150
rect 6720 16990 6760 17130
rect 6720 16970 6730 16990
rect 6750 16970 6760 16990
rect 6720 16960 6760 16970
rect 6800 17150 6840 17160
rect 6800 17130 6810 17150
rect 6830 17130 6840 17150
rect 6800 16990 6840 17130
rect 6800 16970 6810 16990
rect 6830 16970 6840 16990
rect 6800 16960 6840 16970
rect 6880 17150 6920 17160
rect 6880 17130 6890 17150
rect 6910 17130 6920 17150
rect 6880 16990 6920 17130
rect 6880 16970 6890 16990
rect 6910 16970 6920 16990
rect 6880 16960 6920 16970
rect 6960 17150 7000 17160
rect 6960 17130 6970 17150
rect 6990 17130 7000 17150
rect 6960 16990 7000 17130
rect 6960 16970 6970 16990
rect 6990 16970 7000 16990
rect 6960 16960 7000 16970
rect 7040 17150 7080 17160
rect 7040 17130 7050 17150
rect 7070 17130 7080 17150
rect 7040 16990 7080 17130
rect 7040 16970 7050 16990
rect 7070 16970 7080 16990
rect 7040 16960 7080 16970
rect 7120 17150 7160 17160
rect 7120 17130 7130 17150
rect 7150 17130 7160 17150
rect 7120 16990 7160 17130
rect 7120 16970 7130 16990
rect 7150 16970 7160 16990
rect 7120 16960 7160 16970
rect 7200 17150 7240 17160
rect 7200 17130 7210 17150
rect 7230 17130 7240 17150
rect 7200 16990 7240 17130
rect 7200 16970 7210 16990
rect 7230 16970 7240 16990
rect 7200 16960 7240 16970
rect 7280 17150 7320 17160
rect 7280 17130 7290 17150
rect 7310 17130 7320 17150
rect 7280 16990 7320 17130
rect 7280 16970 7290 16990
rect 7310 16970 7320 16990
rect 7280 16960 7320 16970
rect 7360 17150 7400 17160
rect 7360 17130 7370 17150
rect 7390 17130 7400 17150
rect 7360 16990 7400 17130
rect 7360 16970 7370 16990
rect 7390 16970 7400 16990
rect 7360 16960 7400 16970
rect 7440 17150 7480 17160
rect 7440 17130 7450 17150
rect 7470 17130 7480 17150
rect 7440 16990 7480 17130
rect 7440 16970 7450 16990
rect 7470 16970 7480 16990
rect 7440 16960 7480 16970
rect 7520 17150 7560 17160
rect 7520 17130 7530 17150
rect 7550 17130 7560 17150
rect 7520 16990 7560 17130
rect 7520 16970 7530 16990
rect 7550 16970 7560 16990
rect 7520 16960 7560 16970
rect 7600 17150 7640 17160
rect 7600 17130 7610 17150
rect 7630 17130 7640 17150
rect 7600 16990 7640 17130
rect 7600 16970 7610 16990
rect 7630 16970 7640 16990
rect 7600 16960 7640 16970
rect 7680 17150 7720 17160
rect 7680 17130 7690 17150
rect 7710 17130 7720 17150
rect 7680 16990 7720 17130
rect 7680 16970 7690 16990
rect 7710 16970 7720 16990
rect 7680 16960 7720 16970
rect 7760 17150 7800 17160
rect 7760 17130 7770 17150
rect 7790 17130 7800 17150
rect 7760 16990 7800 17130
rect 7760 16970 7770 16990
rect 7790 16970 7800 16990
rect 7760 16960 7800 16970
rect 7840 17150 7880 17160
rect 7840 17130 7850 17150
rect 7870 17130 7880 17150
rect 7840 16990 7880 17130
rect 7840 16970 7850 16990
rect 7870 16970 7880 16990
rect 7840 16960 7880 16970
rect 7920 17150 7960 17160
rect 7920 17130 7930 17150
rect 7950 17130 7960 17150
rect 7920 16990 7960 17130
rect 7920 16970 7930 16990
rect 7950 16970 7960 16990
rect 7920 16960 7960 16970
rect 8000 17150 8040 17160
rect 8000 17130 8010 17150
rect 8030 17130 8040 17150
rect 8000 16990 8040 17130
rect 8000 16970 8010 16990
rect 8030 16970 8040 16990
rect 8000 16960 8040 16970
rect 8080 17150 8120 17160
rect 8080 17130 8090 17150
rect 8110 17130 8120 17150
rect 8080 16990 8120 17130
rect 8080 16970 8090 16990
rect 8110 16970 8120 16990
rect 8080 16960 8120 16970
rect 8160 17150 8200 17160
rect 8160 17130 8170 17150
rect 8190 17130 8200 17150
rect 8160 16990 8200 17130
rect 8160 16970 8170 16990
rect 8190 16970 8200 16990
rect 8160 16960 8200 16970
rect 8240 17150 8280 17160
rect 8240 17130 8250 17150
rect 8270 17130 8280 17150
rect 8240 16990 8280 17130
rect 8240 16970 8250 16990
rect 8270 16970 8280 16990
rect 8240 16960 8280 16970
rect 8320 17150 8360 17160
rect 8320 17130 8330 17150
rect 8350 17130 8360 17150
rect 8320 16990 8360 17130
rect 8320 16970 8330 16990
rect 8350 16970 8360 16990
rect 8320 16960 8360 16970
rect 8400 17150 8440 17160
rect 8400 17130 8410 17150
rect 8430 17130 8440 17150
rect 8400 16990 8440 17130
rect 8400 16970 8410 16990
rect 8430 16970 8440 16990
rect 8400 16960 8440 16970
rect 8480 17150 8520 17160
rect 8480 17130 8490 17150
rect 8510 17130 8520 17150
rect 8480 16990 8520 17130
rect 8480 16970 8490 16990
rect 8510 16970 8520 16990
rect 8480 16960 8520 16970
rect 8560 17150 8600 17160
rect 8560 17130 8570 17150
rect 8590 17130 8600 17150
rect 8560 16990 8600 17130
rect 8560 16970 8570 16990
rect 8590 16970 8600 16990
rect 8560 16960 8600 16970
rect 8640 17150 8680 17160
rect 8640 17130 8650 17150
rect 8670 17130 8680 17150
rect 8640 16990 8680 17130
rect 8640 16970 8650 16990
rect 8670 16970 8680 16990
rect 8640 16960 8680 16970
rect 8720 17150 8760 17160
rect 8720 17130 8730 17150
rect 8750 17130 8760 17150
rect 8720 16990 8760 17130
rect 8720 16970 8730 16990
rect 8750 16970 8760 16990
rect 8720 16960 8760 16970
rect 8800 17150 8840 17160
rect 8800 17130 8810 17150
rect 8830 17130 8840 17150
rect 8800 16990 8840 17130
rect 8800 16970 8810 16990
rect 8830 16970 8840 16990
rect 8800 16960 8840 16970
rect 8880 17150 8920 17160
rect 8880 17130 8890 17150
rect 8910 17130 8920 17150
rect 8880 16990 8920 17130
rect 8880 16970 8890 16990
rect 8910 16970 8920 16990
rect 8880 16960 8920 16970
rect 8960 17150 9000 17160
rect 8960 17130 8970 17150
rect 8990 17130 9000 17150
rect 8960 16990 9000 17130
rect 8960 16970 8970 16990
rect 8990 16970 9000 16990
rect 8960 16960 9000 16970
rect 9040 17150 9080 17160
rect 9040 17130 9050 17150
rect 9070 17130 9080 17150
rect 9040 16990 9080 17130
rect 9040 16970 9050 16990
rect 9070 16970 9080 16990
rect 9040 16960 9080 16970
rect 9120 17150 9160 17160
rect 9120 17130 9130 17150
rect 9150 17130 9160 17150
rect 9120 16990 9160 17130
rect 9120 16970 9130 16990
rect 9150 16970 9160 16990
rect 9120 16960 9160 16970
rect 9200 17150 9240 17160
rect 9200 17130 9210 17150
rect 9230 17130 9240 17150
rect 9200 16990 9240 17130
rect 9200 16970 9210 16990
rect 9230 16970 9240 16990
rect 9200 16960 9240 16970
rect 9280 17150 9320 17160
rect 9280 17130 9290 17150
rect 9310 17130 9320 17150
rect 9280 16990 9320 17130
rect 9280 16970 9290 16990
rect 9310 16970 9320 16990
rect 9280 16960 9320 16970
rect 9360 17150 9400 17160
rect 9360 17130 9370 17150
rect 9390 17130 9400 17150
rect 9360 16990 9400 17130
rect 9360 16970 9370 16990
rect 9390 16970 9400 16990
rect 9360 16960 9400 16970
rect 9440 17150 9480 17160
rect 9440 17130 9450 17150
rect 9470 17130 9480 17150
rect 9440 16990 9480 17130
rect 9440 16970 9450 16990
rect 9470 16970 9480 16990
rect 9440 16960 9480 16970
rect 9520 16960 9560 17160
rect 9600 16960 9640 17160
rect 9680 16960 9720 17160
rect 9760 16960 9800 17160
rect 9840 16960 9880 17160
rect 9920 16960 9960 17160
rect 10000 16960 10040 17160
rect 10080 16960 10120 17160
rect 10160 16960 10200 17160
rect 10240 16960 10280 17160
rect 10320 16960 10360 17160
rect 10400 16960 10440 17160
rect 10480 16960 10520 17160
rect 10560 16960 10600 17160
rect 10640 16960 10680 17160
rect 10720 16960 10760 17160
rect 10800 16960 10840 17160
rect 10880 16960 10920 17160
rect 10960 16960 11000 17160
rect 11040 16960 11080 17160
rect 11120 16960 11160 17160
rect 11200 16960 11240 17160
rect 11280 16960 11320 17160
rect 11360 16960 11400 17160
rect 11440 16960 11480 17160
rect 11560 17150 11600 17160
rect 11560 17130 11570 17150
rect 11590 17130 11600 17150
rect 11560 16990 11600 17130
rect 11560 16970 11570 16990
rect 11590 16970 11600 16990
rect 11560 16960 11600 16970
rect 11640 17150 11680 17160
rect 11640 17130 11650 17150
rect 11670 17130 11680 17150
rect 11640 16990 11680 17130
rect 11640 16970 11650 16990
rect 11670 16970 11680 16990
rect 11640 16960 11680 16970
rect 11720 17150 11760 17160
rect 11720 17130 11730 17150
rect 11750 17130 11760 17150
rect 11720 16990 11760 17130
rect 11720 16970 11730 16990
rect 11750 16970 11760 16990
rect 11720 16960 11760 16970
rect 11800 17150 11840 17160
rect 11800 17130 11810 17150
rect 11830 17130 11840 17150
rect 11800 16990 11840 17130
rect 11800 16970 11810 16990
rect 11830 16970 11840 16990
rect 11800 16960 11840 16970
rect 11880 17150 11920 17160
rect 11880 17130 11890 17150
rect 11910 17130 11920 17150
rect 11880 16990 11920 17130
rect 11880 16970 11890 16990
rect 11910 16970 11920 16990
rect 11880 16960 11920 16970
rect 11960 17150 12000 17160
rect 11960 17130 11970 17150
rect 11990 17130 12000 17150
rect 11960 16990 12000 17130
rect 11960 16970 11970 16990
rect 11990 16970 12000 16990
rect 11960 16960 12000 16970
rect 12040 17150 12080 17160
rect 12040 17130 12050 17150
rect 12070 17130 12080 17150
rect 12040 16990 12080 17130
rect 12040 16970 12050 16990
rect 12070 16970 12080 16990
rect 12040 16960 12080 16970
rect 12120 17150 12160 17160
rect 12120 17130 12130 17150
rect 12150 17130 12160 17150
rect 12120 16990 12160 17130
rect 12120 16970 12130 16990
rect 12150 16970 12160 16990
rect 12120 16960 12160 16970
rect 12200 17150 12240 17160
rect 12200 17130 12210 17150
rect 12230 17130 12240 17150
rect 12200 16990 12240 17130
rect 12200 16970 12210 16990
rect 12230 16970 12240 16990
rect 12200 16960 12240 16970
rect 12280 17150 12320 17160
rect 12280 17130 12290 17150
rect 12310 17130 12320 17150
rect 12280 16990 12320 17130
rect 12280 16970 12290 16990
rect 12310 16970 12320 16990
rect 12280 16960 12320 16970
rect 12360 17150 12400 17160
rect 12360 17130 12370 17150
rect 12390 17130 12400 17150
rect 12360 16990 12400 17130
rect 12360 16970 12370 16990
rect 12390 16970 12400 16990
rect 12360 16960 12400 16970
rect 12440 17150 12480 17160
rect 12440 17130 12450 17150
rect 12470 17130 12480 17150
rect 12440 16990 12480 17130
rect 12440 16970 12450 16990
rect 12470 16970 12480 16990
rect 12440 16960 12480 16970
rect 12520 17150 12560 17160
rect 12520 17130 12530 17150
rect 12550 17130 12560 17150
rect 12520 16990 12560 17130
rect 12520 16970 12530 16990
rect 12550 16970 12560 16990
rect 12520 16960 12560 16970
rect 12600 17150 12640 17160
rect 12600 17130 12610 17150
rect 12630 17130 12640 17150
rect 12600 16990 12640 17130
rect 12600 16970 12610 16990
rect 12630 16970 12640 16990
rect 12600 16960 12640 16970
rect 12680 17150 12720 17160
rect 12680 17130 12690 17150
rect 12710 17130 12720 17150
rect 12680 16990 12720 17130
rect 12680 16970 12690 16990
rect 12710 16970 12720 16990
rect 12680 16960 12720 16970
rect 12760 17150 12800 17160
rect 12760 17130 12770 17150
rect 12790 17130 12800 17150
rect 12760 16990 12800 17130
rect 12760 16970 12770 16990
rect 12790 16970 12800 16990
rect 12760 16960 12800 16970
rect 12840 17150 12880 17160
rect 12840 17130 12850 17150
rect 12870 17130 12880 17150
rect 12840 16990 12880 17130
rect 12840 16970 12850 16990
rect 12870 16970 12880 16990
rect 12840 16960 12880 16970
rect 12920 17150 12960 17160
rect 12920 17130 12930 17150
rect 12950 17130 12960 17150
rect 12920 16990 12960 17130
rect 12920 16970 12930 16990
rect 12950 16970 12960 16990
rect 12920 16960 12960 16970
rect 13000 17150 13040 17160
rect 13000 17130 13010 17150
rect 13030 17130 13040 17150
rect 13000 16990 13040 17130
rect 13000 16970 13010 16990
rect 13030 16970 13040 16990
rect 13000 16960 13040 16970
rect 13080 17150 13120 17160
rect 13080 17130 13090 17150
rect 13110 17130 13120 17150
rect 13080 16990 13120 17130
rect 13080 16970 13090 16990
rect 13110 16970 13120 16990
rect 13080 16960 13120 16970
rect 13160 17150 13200 17160
rect 13160 17130 13170 17150
rect 13190 17130 13200 17150
rect 13160 16990 13200 17130
rect 13160 16970 13170 16990
rect 13190 16970 13200 16990
rect 13160 16960 13200 16970
rect 13240 17150 13280 17160
rect 13240 17130 13250 17150
rect 13270 17130 13280 17150
rect 13240 16990 13280 17130
rect 13240 16970 13250 16990
rect 13270 16970 13280 16990
rect 13240 16960 13280 16970
rect 13320 17150 13360 17160
rect 13320 17130 13330 17150
rect 13350 17130 13360 17150
rect 13320 16990 13360 17130
rect 13320 16970 13330 16990
rect 13350 16970 13360 16990
rect 13320 16960 13360 16970
rect 13400 17150 13440 17160
rect 13400 17130 13410 17150
rect 13430 17130 13440 17150
rect 13400 16990 13440 17130
rect 13400 16970 13410 16990
rect 13430 16970 13440 16990
rect 13400 16960 13440 16970
rect 13480 17150 13520 17160
rect 13480 17130 13490 17150
rect 13510 17130 13520 17150
rect 13480 16990 13520 17130
rect 13480 16970 13490 16990
rect 13510 16970 13520 16990
rect 13480 16960 13520 16970
rect 13560 17150 13600 17160
rect 13560 17130 13570 17150
rect 13590 17130 13600 17150
rect 13560 16990 13600 17130
rect 13560 16970 13570 16990
rect 13590 16970 13600 16990
rect 13560 16960 13600 16970
rect 13640 17150 13680 17160
rect 13640 17130 13650 17150
rect 13670 17130 13680 17150
rect 13640 16990 13680 17130
rect 13640 16970 13650 16990
rect 13670 16970 13680 16990
rect 13640 16960 13680 16970
rect 13720 17150 13760 17160
rect 13720 17130 13730 17150
rect 13750 17130 13760 17150
rect 13720 16990 13760 17130
rect 13720 16970 13730 16990
rect 13750 16970 13760 16990
rect 13720 16960 13760 16970
rect 13800 17150 13840 17160
rect 13800 17130 13810 17150
rect 13830 17130 13840 17150
rect 13800 16990 13840 17130
rect 13800 16970 13810 16990
rect 13830 16970 13840 16990
rect 13800 16960 13840 16970
rect 13880 17150 13920 17160
rect 13880 17130 13890 17150
rect 13910 17130 13920 17150
rect 13880 16990 13920 17130
rect 13880 16970 13890 16990
rect 13910 16970 13920 16990
rect 13880 16960 13920 16970
rect 13960 17150 14000 17160
rect 13960 17130 13970 17150
rect 13990 17130 14000 17150
rect 13960 16990 14000 17130
rect 13960 16970 13970 16990
rect 13990 16970 14000 16990
rect 13960 16960 14000 16970
rect 14040 17150 14080 17160
rect 14040 17130 14050 17150
rect 14070 17130 14080 17150
rect 14040 16990 14080 17130
rect 14040 16970 14050 16990
rect 14070 16970 14080 16990
rect 14040 16960 14080 16970
rect 14120 17150 14160 17160
rect 14120 17130 14130 17150
rect 14150 17130 14160 17150
rect 14120 16990 14160 17130
rect 14120 16970 14130 16990
rect 14150 16970 14160 16990
rect 14120 16960 14160 16970
rect 14200 17150 14240 17160
rect 14200 17130 14210 17150
rect 14230 17130 14240 17150
rect 14200 16990 14240 17130
rect 14200 16970 14210 16990
rect 14230 16970 14240 16990
rect 14200 16960 14240 16970
rect 14280 17150 14320 17160
rect 14280 17130 14290 17150
rect 14310 17130 14320 17150
rect 14280 16990 14320 17130
rect 14280 16970 14290 16990
rect 14310 16970 14320 16990
rect 14280 16960 14320 16970
rect 14360 17150 14400 17160
rect 14360 17130 14370 17150
rect 14390 17130 14400 17150
rect 14360 16990 14400 17130
rect 14360 16970 14370 16990
rect 14390 16970 14400 16990
rect 14360 16960 14400 16970
rect 14440 17150 14480 17160
rect 14440 17130 14450 17150
rect 14470 17130 14480 17150
rect 14440 16990 14480 17130
rect 14440 16970 14450 16990
rect 14470 16970 14480 16990
rect 14440 16960 14480 16970
rect 14520 17150 14560 17160
rect 14520 17130 14530 17150
rect 14550 17130 14560 17150
rect 14520 16990 14560 17130
rect 14520 16970 14530 16990
rect 14550 16970 14560 16990
rect 14520 16960 14560 16970
rect 14600 17150 14640 17160
rect 14600 17130 14610 17150
rect 14630 17130 14640 17150
rect 14600 16990 14640 17130
rect 14600 16970 14610 16990
rect 14630 16970 14640 16990
rect 14600 16960 14640 16970
rect 14680 17150 14720 17160
rect 14680 17130 14690 17150
rect 14710 17130 14720 17150
rect 14680 16990 14720 17130
rect 14680 16970 14690 16990
rect 14710 16970 14720 16990
rect 14680 16960 14720 16970
rect 14760 16960 14800 17160
rect 14840 16960 14880 17160
rect 14920 16960 14960 17160
rect 15000 16960 15040 17160
rect 15080 16960 15120 17160
rect 15160 16960 15200 17160
rect 15240 16960 15280 17160
rect 15320 16960 15360 17160
rect 15400 16960 15440 17160
rect 15480 16960 15520 17160
rect 15560 16960 15600 17160
rect 15640 16960 15680 17160
rect 15720 16960 15760 17160
rect 15800 16960 15840 17160
rect 15880 16960 15920 17160
rect 15960 16960 16000 17160
rect 16040 16960 16080 17160
rect 16120 16960 16160 17160
rect 16200 16960 16240 17160
rect 16280 16960 16320 17160
rect 16360 16960 16400 17160
rect 16440 16960 16480 17160
rect 16520 16960 16560 17160
rect 16600 16960 16640 17160
rect 16680 16960 16720 17160
rect 16760 17150 16800 17160
rect 16760 17130 16770 17150
rect 16790 17130 16800 17150
rect 16760 16990 16800 17130
rect 16760 16970 16770 16990
rect 16790 16970 16800 16990
rect 16760 16960 16800 16970
rect 16840 17150 16880 17160
rect 16840 17130 16850 17150
rect 16870 17130 16880 17150
rect 16840 16990 16880 17130
rect 16840 16970 16850 16990
rect 16870 16970 16880 16990
rect 16840 16960 16880 16970
rect 16920 17150 16960 17160
rect 16920 17130 16930 17150
rect 16950 17130 16960 17150
rect 16920 16990 16960 17130
rect 16920 16970 16930 16990
rect 16950 16970 16960 16990
rect 16920 16960 16960 16970
rect 17000 17150 17040 17160
rect 17000 17130 17010 17150
rect 17030 17130 17040 17150
rect 17000 16990 17040 17130
rect 17000 16970 17010 16990
rect 17030 16970 17040 16990
rect 17000 16960 17040 16970
rect 17080 17150 17120 17160
rect 17080 17130 17090 17150
rect 17110 17130 17120 17150
rect 17080 16990 17120 17130
rect 17080 16970 17090 16990
rect 17110 16970 17120 16990
rect 17080 16960 17120 16970
rect 17160 17150 17200 17160
rect 17160 17130 17170 17150
rect 17190 17130 17200 17150
rect 17160 16990 17200 17130
rect 17160 16970 17170 16990
rect 17190 16970 17200 16990
rect 17160 16960 17200 16970
rect 17240 17150 17280 17160
rect 17240 17130 17250 17150
rect 17270 17130 17280 17150
rect 17240 16990 17280 17130
rect 17240 16970 17250 16990
rect 17270 16970 17280 16990
rect 17240 16960 17280 16970
rect 17320 17150 17360 17160
rect 17320 17130 17330 17150
rect 17350 17130 17360 17150
rect 17320 16990 17360 17130
rect 17320 16970 17330 16990
rect 17350 16970 17360 16990
rect 17320 16960 17360 16970
rect 17400 17150 17440 17160
rect 17400 17130 17410 17150
rect 17430 17130 17440 17150
rect 17400 16990 17440 17130
rect 17400 16970 17410 16990
rect 17430 16970 17440 16990
rect 17400 16960 17440 16970
rect 17480 17150 17520 17160
rect 17480 17130 17490 17150
rect 17510 17130 17520 17150
rect 17480 16990 17520 17130
rect 17480 16970 17490 16990
rect 17510 16970 17520 16990
rect 17480 16960 17520 16970
rect 17560 17150 17600 17160
rect 17560 17130 17570 17150
rect 17590 17130 17600 17150
rect 17560 16990 17600 17130
rect 17560 16970 17570 16990
rect 17590 16970 17600 16990
rect 17560 16960 17600 16970
rect 17640 17150 17680 17160
rect 17640 17130 17650 17150
rect 17670 17130 17680 17150
rect 17640 16990 17680 17130
rect 17640 16970 17650 16990
rect 17670 16970 17680 16990
rect 17640 16960 17680 16970
rect 17720 17150 17760 17160
rect 17720 17130 17730 17150
rect 17750 17130 17760 17150
rect 17720 16990 17760 17130
rect 17720 16970 17730 16990
rect 17750 16970 17760 16990
rect 17720 16960 17760 16970
rect 17800 17150 17840 17160
rect 17800 17130 17810 17150
rect 17830 17130 17840 17150
rect 17800 16990 17840 17130
rect 17800 16970 17810 16990
rect 17830 16970 17840 16990
rect 17800 16960 17840 16970
rect 17880 17150 17920 17160
rect 17880 17130 17890 17150
rect 17910 17130 17920 17150
rect 17880 16990 17920 17130
rect 17880 16970 17890 16990
rect 17910 16970 17920 16990
rect 17880 16960 17920 16970
rect 17960 17150 18000 17160
rect 17960 17130 17970 17150
rect 17990 17130 18000 17150
rect 17960 16990 18000 17130
rect 17960 16970 17970 16990
rect 17990 16970 18000 16990
rect 17960 16960 18000 16970
rect 18040 17150 18080 17160
rect 18040 17130 18050 17150
rect 18070 17130 18080 17150
rect 18040 16990 18080 17130
rect 18040 16970 18050 16990
rect 18070 16970 18080 16990
rect 18040 16960 18080 16970
rect 18120 17150 18160 17160
rect 18120 17130 18130 17150
rect 18150 17130 18160 17150
rect 18120 16990 18160 17130
rect 18120 16970 18130 16990
rect 18150 16970 18160 16990
rect 18120 16960 18160 16970
rect 18200 17150 18240 17160
rect 18200 17130 18210 17150
rect 18230 17130 18240 17150
rect 18200 16990 18240 17130
rect 18200 16970 18210 16990
rect 18230 16970 18240 16990
rect 18200 16960 18240 16970
rect 18280 17150 18320 17160
rect 18280 17130 18290 17150
rect 18310 17130 18320 17150
rect 18280 16990 18320 17130
rect 18280 16970 18290 16990
rect 18310 16970 18320 16990
rect 18280 16960 18320 16970
rect 18360 17150 18400 17160
rect 18360 17130 18370 17150
rect 18390 17130 18400 17150
rect 18360 16990 18400 17130
rect 18360 16970 18370 16990
rect 18390 16970 18400 16990
rect 18360 16960 18400 16970
rect 18440 17150 18480 17160
rect 18440 17130 18450 17150
rect 18470 17130 18480 17150
rect 18440 16990 18480 17130
rect 18440 16970 18450 16990
rect 18470 16970 18480 16990
rect 18440 16960 18480 16970
rect 18520 17150 18560 17160
rect 18520 17130 18530 17150
rect 18550 17130 18560 17150
rect 18520 16990 18560 17130
rect 18520 16970 18530 16990
rect 18550 16970 18560 16990
rect 18520 16960 18560 16970
rect 18600 17150 18640 17160
rect 18600 17130 18610 17150
rect 18630 17130 18640 17150
rect 18600 16990 18640 17130
rect 18600 16970 18610 16990
rect 18630 16970 18640 16990
rect 18600 16960 18640 16970
rect 18680 17150 18720 17160
rect 18680 17130 18690 17150
rect 18710 17130 18720 17150
rect 18680 16990 18720 17130
rect 18680 16970 18690 16990
rect 18710 16970 18720 16990
rect 18680 16960 18720 16970
rect 18760 17150 18800 17160
rect 18760 17130 18770 17150
rect 18790 17130 18800 17150
rect 18760 16990 18800 17130
rect 18760 16970 18770 16990
rect 18790 16970 18800 16990
rect 18760 16960 18800 16970
rect 18840 17150 18880 17160
rect 18840 17130 18850 17150
rect 18870 17130 18880 17150
rect 18840 16990 18880 17130
rect 18840 16970 18850 16990
rect 18870 16970 18880 16990
rect 18840 16960 18880 16970
rect 18920 17150 18960 17160
rect 18920 17130 18930 17150
rect 18950 17130 18960 17150
rect 18920 16990 18960 17130
rect 18920 16970 18930 16990
rect 18950 16970 18960 16990
rect 18920 16960 18960 16970
rect 19000 17150 19040 17160
rect 19000 17130 19010 17150
rect 19030 17130 19040 17150
rect 19000 16990 19040 17130
rect 19000 16970 19010 16990
rect 19030 16970 19040 16990
rect 19000 16960 19040 16970
rect 19080 17150 19120 17160
rect 19080 17130 19090 17150
rect 19110 17130 19120 17150
rect 19080 16990 19120 17130
rect 19080 16970 19090 16990
rect 19110 16970 19120 16990
rect 19080 16960 19120 16970
rect 19160 17150 19200 17160
rect 19160 17130 19170 17150
rect 19190 17130 19200 17150
rect 19160 16990 19200 17130
rect 19160 16970 19170 16990
rect 19190 16970 19200 16990
rect 19160 16960 19200 16970
rect 19240 17150 19280 17160
rect 19240 17130 19250 17150
rect 19270 17130 19280 17150
rect 19240 16990 19280 17130
rect 19240 16970 19250 16990
rect 19270 16970 19280 16990
rect 19240 16960 19280 16970
rect 19320 17150 19360 17160
rect 19320 17130 19330 17150
rect 19350 17130 19360 17150
rect 19320 16990 19360 17130
rect 19320 16970 19330 16990
rect 19350 16970 19360 16990
rect 19320 16960 19360 16970
rect 19400 17150 19440 17160
rect 19400 17130 19410 17150
rect 19430 17130 19440 17150
rect 19400 16990 19440 17130
rect 19400 16970 19410 16990
rect 19430 16970 19440 16990
rect 19400 16960 19440 16970
rect 19480 17150 19520 17160
rect 19480 17130 19490 17150
rect 19510 17130 19520 17150
rect 19480 16990 19520 17130
rect 19480 16970 19490 16990
rect 19510 16970 19520 16990
rect 19480 16960 19520 16970
rect 19560 17150 19600 17160
rect 19560 17130 19570 17150
rect 19590 17130 19600 17150
rect 19560 16990 19600 17130
rect 19560 16970 19570 16990
rect 19590 16970 19600 16990
rect 19560 16960 19600 16970
rect 19640 17150 19680 17160
rect 19640 17130 19650 17150
rect 19670 17130 19680 17150
rect 19640 16990 19680 17130
rect 19640 16970 19650 16990
rect 19670 16970 19680 16990
rect 19640 16960 19680 16970
rect 19720 17150 19760 17160
rect 19720 17130 19730 17150
rect 19750 17130 19760 17150
rect 19720 16990 19760 17130
rect 19720 16970 19730 16990
rect 19750 16970 19760 16990
rect 19720 16960 19760 16970
rect 19800 17150 19840 17160
rect 19800 17130 19810 17150
rect 19830 17130 19840 17150
rect 19800 16990 19840 17130
rect 19800 16970 19810 16990
rect 19830 16970 19840 16990
rect 19800 16960 19840 16970
rect 19880 17150 19920 17160
rect 19880 17130 19890 17150
rect 19910 17130 19920 17150
rect 19880 16990 19920 17130
rect 19880 16970 19890 16990
rect 19910 16970 19920 16990
rect 19880 16960 19920 16970
rect 19960 17150 20000 17160
rect 19960 17130 19970 17150
rect 19990 17130 20000 17150
rect 19960 16990 20000 17130
rect 19960 16970 19970 16990
rect 19990 16970 20000 16990
rect 19960 16960 20000 16970
rect 20040 17150 20080 17160
rect 20040 17130 20050 17150
rect 20070 17130 20080 17150
rect 20040 16990 20080 17130
rect 20040 16970 20050 16990
rect 20070 16970 20080 16990
rect 20040 16960 20080 16970
rect 20120 17150 20160 17160
rect 20120 17130 20130 17150
rect 20150 17130 20160 17150
rect 20120 16990 20160 17130
rect 20120 16970 20130 16990
rect 20150 16970 20160 16990
rect 20120 16960 20160 16970
rect 20200 17150 20240 17160
rect 20200 17130 20210 17150
rect 20230 17130 20240 17150
rect 20200 16990 20240 17130
rect 20200 16970 20210 16990
rect 20230 16970 20240 16990
rect 20200 16960 20240 16970
rect 20280 17150 20320 17160
rect 20280 17130 20290 17150
rect 20310 17130 20320 17150
rect 20280 16990 20320 17130
rect 20280 16970 20290 16990
rect 20310 16970 20320 16990
rect 20280 16960 20320 16970
rect 20360 17150 20400 17160
rect 20360 17130 20370 17150
rect 20390 17130 20400 17150
rect 20360 16990 20400 17130
rect 20360 16970 20370 16990
rect 20390 16970 20400 16990
rect 20360 16960 20400 16970
rect 20440 17150 20480 17160
rect 20440 17130 20450 17150
rect 20470 17130 20480 17150
rect 20440 16990 20480 17130
rect 20440 16970 20450 16990
rect 20470 16970 20480 16990
rect 20440 16960 20480 16970
rect 20520 17150 20560 17160
rect 20520 17130 20530 17150
rect 20550 17130 20560 17150
rect 20520 16990 20560 17130
rect 20520 16970 20530 16990
rect 20550 16970 20560 16990
rect 20520 16960 20560 16970
rect 20600 17150 20640 17160
rect 20600 17130 20610 17150
rect 20630 17130 20640 17150
rect 20600 16990 20640 17130
rect 20600 16970 20610 16990
rect 20630 16970 20640 16990
rect 20600 16960 20640 16970
rect 20680 17150 20720 17160
rect 20680 17130 20690 17150
rect 20710 17130 20720 17150
rect 20680 16990 20720 17130
rect 20680 16970 20690 16990
rect 20710 16970 20720 16990
rect 20680 16960 20720 16970
rect 20760 17150 20800 17160
rect 20760 17130 20770 17150
rect 20790 17130 20800 17150
rect 20760 16990 20800 17130
rect 20760 16970 20770 16990
rect 20790 16970 20800 16990
rect 20760 16960 20800 16970
rect 20840 17150 20880 17160
rect 20840 17130 20850 17150
rect 20870 17130 20880 17150
rect 20840 16990 20880 17130
rect 20840 16970 20850 16990
rect 20870 16970 20880 16990
rect 20840 16960 20880 16970
rect 20920 17150 20960 17160
rect 20920 17130 20930 17150
rect 20950 17130 20960 17150
rect 20920 16990 20960 17130
rect 20920 16970 20930 16990
rect 20950 16970 20960 16990
rect 20920 16960 20960 16970
rect 0 16910 40 16920
rect 0 16890 10 16910
rect 30 16890 40 16910
rect 0 16750 40 16890
rect 0 16730 10 16750
rect 30 16730 40 16750
rect 0 16720 40 16730
rect 80 16910 120 16920
rect 80 16890 90 16910
rect 110 16890 120 16910
rect 80 16750 120 16890
rect 80 16730 90 16750
rect 110 16730 120 16750
rect 80 16720 120 16730
rect 160 16910 200 16920
rect 160 16890 170 16910
rect 190 16890 200 16910
rect 160 16750 200 16890
rect 160 16730 170 16750
rect 190 16730 200 16750
rect 160 16720 200 16730
rect 240 16910 280 16920
rect 240 16890 250 16910
rect 270 16890 280 16910
rect 240 16750 280 16890
rect 240 16730 250 16750
rect 270 16730 280 16750
rect 240 16720 280 16730
rect 320 16910 360 16920
rect 320 16890 330 16910
rect 350 16890 360 16910
rect 320 16750 360 16890
rect 320 16730 330 16750
rect 350 16730 360 16750
rect 320 16720 360 16730
rect 400 16910 440 16920
rect 400 16890 410 16910
rect 430 16890 440 16910
rect 400 16750 440 16890
rect 400 16730 410 16750
rect 430 16730 440 16750
rect 400 16720 440 16730
rect 480 16910 520 16920
rect 480 16890 490 16910
rect 510 16890 520 16910
rect 480 16750 520 16890
rect 480 16730 490 16750
rect 510 16730 520 16750
rect 480 16720 520 16730
rect 560 16910 600 16920
rect 560 16890 570 16910
rect 590 16890 600 16910
rect 560 16750 600 16890
rect 560 16730 570 16750
rect 590 16730 600 16750
rect 560 16720 600 16730
rect 640 16910 680 16920
rect 640 16890 650 16910
rect 670 16890 680 16910
rect 640 16750 680 16890
rect 640 16730 650 16750
rect 670 16730 680 16750
rect 640 16720 680 16730
rect 720 16910 760 16920
rect 720 16890 730 16910
rect 750 16890 760 16910
rect 720 16750 760 16890
rect 720 16730 730 16750
rect 750 16730 760 16750
rect 720 16720 760 16730
rect 800 16910 840 16920
rect 800 16890 810 16910
rect 830 16890 840 16910
rect 800 16750 840 16890
rect 800 16730 810 16750
rect 830 16730 840 16750
rect 800 16720 840 16730
rect 880 16910 920 16920
rect 880 16890 890 16910
rect 910 16890 920 16910
rect 880 16750 920 16890
rect 880 16730 890 16750
rect 910 16730 920 16750
rect 880 16720 920 16730
rect 960 16910 1000 16920
rect 960 16890 970 16910
rect 990 16890 1000 16910
rect 960 16750 1000 16890
rect 960 16730 970 16750
rect 990 16730 1000 16750
rect 960 16720 1000 16730
rect 1040 16910 1080 16920
rect 1040 16890 1050 16910
rect 1070 16890 1080 16910
rect 1040 16750 1080 16890
rect 1040 16730 1050 16750
rect 1070 16730 1080 16750
rect 1040 16720 1080 16730
rect 1120 16910 1160 16920
rect 1120 16890 1130 16910
rect 1150 16890 1160 16910
rect 1120 16750 1160 16890
rect 1120 16730 1130 16750
rect 1150 16730 1160 16750
rect 1120 16720 1160 16730
rect 1200 16910 1240 16920
rect 1200 16890 1210 16910
rect 1230 16890 1240 16910
rect 1200 16750 1240 16890
rect 1200 16730 1210 16750
rect 1230 16730 1240 16750
rect 1200 16720 1240 16730
rect 1280 16910 1320 16920
rect 1280 16890 1290 16910
rect 1310 16890 1320 16910
rect 1280 16750 1320 16890
rect 1280 16730 1290 16750
rect 1310 16730 1320 16750
rect 1280 16720 1320 16730
rect 1360 16910 1400 16920
rect 1360 16890 1370 16910
rect 1390 16890 1400 16910
rect 1360 16750 1400 16890
rect 1360 16730 1370 16750
rect 1390 16730 1400 16750
rect 1360 16720 1400 16730
rect 1440 16910 1480 16920
rect 1440 16890 1450 16910
rect 1470 16890 1480 16910
rect 1440 16750 1480 16890
rect 1440 16730 1450 16750
rect 1470 16730 1480 16750
rect 1440 16720 1480 16730
rect 1520 16910 1560 16920
rect 1520 16890 1530 16910
rect 1550 16890 1560 16910
rect 1520 16750 1560 16890
rect 1520 16730 1530 16750
rect 1550 16730 1560 16750
rect 1520 16720 1560 16730
rect 1600 16910 1640 16920
rect 1600 16890 1610 16910
rect 1630 16890 1640 16910
rect 1600 16750 1640 16890
rect 1600 16730 1610 16750
rect 1630 16730 1640 16750
rect 1600 16720 1640 16730
rect 1680 16910 1720 16920
rect 1680 16890 1690 16910
rect 1710 16890 1720 16910
rect 1680 16750 1720 16890
rect 1680 16730 1690 16750
rect 1710 16730 1720 16750
rect 1680 16720 1720 16730
rect 1760 16910 1800 16920
rect 1760 16890 1770 16910
rect 1790 16890 1800 16910
rect 1760 16750 1800 16890
rect 1760 16730 1770 16750
rect 1790 16730 1800 16750
rect 1760 16720 1800 16730
rect 1840 16910 1880 16920
rect 1840 16890 1850 16910
rect 1870 16890 1880 16910
rect 1840 16750 1880 16890
rect 1840 16730 1850 16750
rect 1870 16730 1880 16750
rect 1840 16720 1880 16730
rect 1920 16910 1960 16920
rect 1920 16890 1930 16910
rect 1950 16890 1960 16910
rect 1920 16750 1960 16890
rect 1920 16730 1930 16750
rect 1950 16730 1960 16750
rect 1920 16720 1960 16730
rect 2000 16910 2040 16920
rect 2000 16890 2010 16910
rect 2030 16890 2040 16910
rect 2000 16750 2040 16890
rect 2000 16730 2010 16750
rect 2030 16730 2040 16750
rect 2000 16720 2040 16730
rect 2080 16910 2120 16920
rect 2080 16890 2090 16910
rect 2110 16890 2120 16910
rect 2080 16750 2120 16890
rect 2080 16730 2090 16750
rect 2110 16730 2120 16750
rect 2080 16720 2120 16730
rect 2160 16910 2200 16920
rect 2160 16890 2170 16910
rect 2190 16890 2200 16910
rect 2160 16750 2200 16890
rect 2160 16730 2170 16750
rect 2190 16730 2200 16750
rect 2160 16720 2200 16730
rect 2240 16910 2280 16920
rect 2240 16890 2250 16910
rect 2270 16890 2280 16910
rect 2240 16750 2280 16890
rect 2240 16730 2250 16750
rect 2270 16730 2280 16750
rect 2240 16720 2280 16730
rect 2320 16910 2360 16920
rect 2320 16890 2330 16910
rect 2350 16890 2360 16910
rect 2320 16750 2360 16890
rect 2320 16730 2330 16750
rect 2350 16730 2360 16750
rect 2320 16720 2360 16730
rect 2400 16910 2440 16920
rect 2400 16890 2410 16910
rect 2430 16890 2440 16910
rect 2400 16750 2440 16890
rect 2400 16730 2410 16750
rect 2430 16730 2440 16750
rect 2400 16720 2440 16730
rect 2480 16910 2520 16920
rect 2480 16890 2490 16910
rect 2510 16890 2520 16910
rect 2480 16750 2520 16890
rect 2480 16730 2490 16750
rect 2510 16730 2520 16750
rect 2480 16720 2520 16730
rect 2560 16910 2600 16920
rect 2560 16890 2570 16910
rect 2590 16890 2600 16910
rect 2560 16750 2600 16890
rect 2560 16730 2570 16750
rect 2590 16730 2600 16750
rect 2560 16720 2600 16730
rect 2640 16910 2680 16920
rect 2640 16890 2650 16910
rect 2670 16890 2680 16910
rect 2640 16750 2680 16890
rect 2640 16730 2650 16750
rect 2670 16730 2680 16750
rect 2640 16720 2680 16730
rect 2720 16910 2760 16920
rect 2720 16890 2730 16910
rect 2750 16890 2760 16910
rect 2720 16750 2760 16890
rect 2720 16730 2730 16750
rect 2750 16730 2760 16750
rect 2720 16720 2760 16730
rect 2800 16910 2840 16920
rect 2800 16890 2810 16910
rect 2830 16890 2840 16910
rect 2800 16750 2840 16890
rect 2800 16730 2810 16750
rect 2830 16730 2840 16750
rect 2800 16720 2840 16730
rect 2880 16910 2920 16920
rect 2880 16890 2890 16910
rect 2910 16890 2920 16910
rect 2880 16750 2920 16890
rect 2880 16730 2890 16750
rect 2910 16730 2920 16750
rect 2880 16720 2920 16730
rect 2960 16910 3000 16920
rect 2960 16890 2970 16910
rect 2990 16890 3000 16910
rect 2960 16750 3000 16890
rect 2960 16730 2970 16750
rect 2990 16730 3000 16750
rect 2960 16720 3000 16730
rect 3040 16910 3080 16920
rect 3040 16890 3050 16910
rect 3070 16890 3080 16910
rect 3040 16750 3080 16890
rect 3040 16730 3050 16750
rect 3070 16730 3080 16750
rect 3040 16720 3080 16730
rect 3120 16910 3160 16920
rect 3120 16890 3130 16910
rect 3150 16890 3160 16910
rect 3120 16750 3160 16890
rect 3120 16730 3130 16750
rect 3150 16730 3160 16750
rect 3120 16720 3160 16730
rect 3200 16910 3240 16920
rect 3200 16890 3210 16910
rect 3230 16890 3240 16910
rect 3200 16750 3240 16890
rect 3200 16730 3210 16750
rect 3230 16730 3240 16750
rect 3200 16720 3240 16730
rect 3280 16910 3320 16920
rect 3280 16890 3290 16910
rect 3310 16890 3320 16910
rect 3280 16750 3320 16890
rect 3280 16730 3290 16750
rect 3310 16730 3320 16750
rect 3280 16720 3320 16730
rect 3360 16910 3400 16920
rect 3360 16890 3370 16910
rect 3390 16890 3400 16910
rect 3360 16750 3400 16890
rect 3360 16730 3370 16750
rect 3390 16730 3400 16750
rect 3360 16720 3400 16730
rect 3440 16910 3480 16920
rect 3440 16890 3450 16910
rect 3470 16890 3480 16910
rect 3440 16750 3480 16890
rect 3440 16730 3450 16750
rect 3470 16730 3480 16750
rect 3440 16720 3480 16730
rect 3520 16910 3560 16920
rect 3520 16890 3530 16910
rect 3550 16890 3560 16910
rect 3520 16750 3560 16890
rect 3520 16730 3530 16750
rect 3550 16730 3560 16750
rect 3520 16720 3560 16730
rect 3600 16910 3640 16920
rect 3600 16890 3610 16910
rect 3630 16890 3640 16910
rect 3600 16750 3640 16890
rect 3600 16730 3610 16750
rect 3630 16730 3640 16750
rect 3600 16720 3640 16730
rect 3680 16910 3720 16920
rect 3680 16890 3690 16910
rect 3710 16890 3720 16910
rect 3680 16750 3720 16890
rect 3680 16730 3690 16750
rect 3710 16730 3720 16750
rect 3680 16720 3720 16730
rect 3760 16910 3800 16920
rect 3760 16890 3770 16910
rect 3790 16890 3800 16910
rect 3760 16750 3800 16890
rect 3760 16730 3770 16750
rect 3790 16730 3800 16750
rect 3760 16720 3800 16730
rect 3840 16910 3880 16920
rect 3840 16890 3850 16910
rect 3870 16890 3880 16910
rect 3840 16750 3880 16890
rect 3840 16730 3850 16750
rect 3870 16730 3880 16750
rect 3840 16720 3880 16730
rect 3920 16910 3960 16920
rect 3920 16890 3930 16910
rect 3950 16890 3960 16910
rect 3920 16750 3960 16890
rect 3920 16730 3930 16750
rect 3950 16730 3960 16750
rect 3920 16720 3960 16730
rect 4000 16910 4040 16920
rect 4000 16890 4010 16910
rect 4030 16890 4040 16910
rect 4000 16750 4040 16890
rect 4000 16730 4010 16750
rect 4030 16730 4040 16750
rect 4000 16720 4040 16730
rect 4080 16910 4120 16920
rect 4080 16890 4090 16910
rect 4110 16890 4120 16910
rect 4080 16750 4120 16890
rect 4080 16730 4090 16750
rect 4110 16730 4120 16750
rect 4080 16720 4120 16730
rect 4160 16910 4200 16920
rect 4160 16890 4170 16910
rect 4190 16890 4200 16910
rect 4160 16750 4200 16890
rect 4160 16730 4170 16750
rect 4190 16730 4200 16750
rect 4160 16720 4200 16730
rect 4240 16720 4280 16920
rect 4320 16720 4360 16920
rect 4400 16720 4440 16920
rect 4480 16720 4520 16920
rect 4560 16720 4600 16920
rect 4640 16720 4680 16920
rect 4720 16720 4760 16920
rect 4800 16720 4840 16920
rect 4880 16720 4920 16920
rect 4960 16720 5000 16920
rect 5040 16720 5080 16920
rect 5120 16720 5160 16920
rect 5200 16720 5240 16920
rect 5280 16720 5320 16920
rect 5360 16720 5400 16920
rect 5440 16720 5480 16920
rect 5520 16720 5560 16920
rect 5600 16720 5640 16920
rect 5680 16720 5720 16920
rect 5760 16720 5800 16920
rect 5840 16720 5880 16920
rect 5920 16720 5960 16920
rect 6000 16720 6040 16920
rect 6080 16720 6120 16920
rect 6160 16720 6200 16920
rect 6240 16910 6280 16920
rect 6240 16890 6250 16910
rect 6270 16890 6280 16910
rect 6240 16750 6280 16890
rect 6240 16730 6250 16750
rect 6270 16730 6280 16750
rect 6240 16720 6280 16730
rect 6320 16910 6360 16920
rect 6320 16890 6330 16910
rect 6350 16890 6360 16910
rect 6320 16750 6360 16890
rect 6320 16730 6330 16750
rect 6350 16730 6360 16750
rect 6320 16720 6360 16730
rect 6400 16910 6440 16920
rect 6400 16890 6410 16910
rect 6430 16890 6440 16910
rect 6400 16750 6440 16890
rect 6400 16730 6410 16750
rect 6430 16730 6440 16750
rect 6400 16720 6440 16730
rect 6480 16910 6520 16920
rect 6480 16890 6490 16910
rect 6510 16890 6520 16910
rect 6480 16750 6520 16890
rect 6480 16730 6490 16750
rect 6510 16730 6520 16750
rect 6480 16720 6520 16730
rect 6560 16910 6600 16920
rect 6560 16890 6570 16910
rect 6590 16890 6600 16910
rect 6560 16750 6600 16890
rect 6560 16730 6570 16750
rect 6590 16730 6600 16750
rect 6560 16720 6600 16730
rect 6640 16910 6680 16920
rect 6640 16890 6650 16910
rect 6670 16890 6680 16910
rect 6640 16750 6680 16890
rect 6640 16730 6650 16750
rect 6670 16730 6680 16750
rect 6640 16720 6680 16730
rect 6720 16910 6760 16920
rect 6720 16890 6730 16910
rect 6750 16890 6760 16910
rect 6720 16750 6760 16890
rect 6720 16730 6730 16750
rect 6750 16730 6760 16750
rect 6720 16720 6760 16730
rect 6800 16910 6840 16920
rect 6800 16890 6810 16910
rect 6830 16890 6840 16910
rect 6800 16750 6840 16890
rect 6800 16730 6810 16750
rect 6830 16730 6840 16750
rect 6800 16720 6840 16730
rect 6880 16910 6920 16920
rect 6880 16890 6890 16910
rect 6910 16890 6920 16910
rect 6880 16750 6920 16890
rect 6880 16730 6890 16750
rect 6910 16730 6920 16750
rect 6880 16720 6920 16730
rect 6960 16910 7000 16920
rect 6960 16890 6970 16910
rect 6990 16890 7000 16910
rect 6960 16750 7000 16890
rect 6960 16730 6970 16750
rect 6990 16730 7000 16750
rect 6960 16720 7000 16730
rect 7040 16910 7080 16920
rect 7040 16890 7050 16910
rect 7070 16890 7080 16910
rect 7040 16750 7080 16890
rect 7040 16730 7050 16750
rect 7070 16730 7080 16750
rect 7040 16720 7080 16730
rect 7120 16910 7160 16920
rect 7120 16890 7130 16910
rect 7150 16890 7160 16910
rect 7120 16750 7160 16890
rect 7120 16730 7130 16750
rect 7150 16730 7160 16750
rect 7120 16720 7160 16730
rect 7200 16910 7240 16920
rect 7200 16890 7210 16910
rect 7230 16890 7240 16910
rect 7200 16750 7240 16890
rect 7200 16730 7210 16750
rect 7230 16730 7240 16750
rect 7200 16720 7240 16730
rect 7280 16910 7320 16920
rect 7280 16890 7290 16910
rect 7310 16890 7320 16910
rect 7280 16750 7320 16890
rect 7280 16730 7290 16750
rect 7310 16730 7320 16750
rect 7280 16720 7320 16730
rect 7360 16910 7400 16920
rect 7360 16890 7370 16910
rect 7390 16890 7400 16910
rect 7360 16750 7400 16890
rect 7360 16730 7370 16750
rect 7390 16730 7400 16750
rect 7360 16720 7400 16730
rect 7440 16910 7480 16920
rect 7440 16890 7450 16910
rect 7470 16890 7480 16910
rect 7440 16750 7480 16890
rect 7440 16730 7450 16750
rect 7470 16730 7480 16750
rect 7440 16720 7480 16730
rect 7520 16910 7560 16920
rect 7520 16890 7530 16910
rect 7550 16890 7560 16910
rect 7520 16750 7560 16890
rect 7520 16730 7530 16750
rect 7550 16730 7560 16750
rect 7520 16720 7560 16730
rect 7600 16910 7640 16920
rect 7600 16890 7610 16910
rect 7630 16890 7640 16910
rect 7600 16750 7640 16890
rect 7600 16730 7610 16750
rect 7630 16730 7640 16750
rect 7600 16720 7640 16730
rect 7680 16910 7720 16920
rect 7680 16890 7690 16910
rect 7710 16890 7720 16910
rect 7680 16750 7720 16890
rect 7680 16730 7690 16750
rect 7710 16730 7720 16750
rect 7680 16720 7720 16730
rect 7760 16910 7800 16920
rect 7760 16890 7770 16910
rect 7790 16890 7800 16910
rect 7760 16750 7800 16890
rect 7760 16730 7770 16750
rect 7790 16730 7800 16750
rect 7760 16720 7800 16730
rect 7840 16910 7880 16920
rect 7840 16890 7850 16910
rect 7870 16890 7880 16910
rect 7840 16750 7880 16890
rect 7840 16730 7850 16750
rect 7870 16730 7880 16750
rect 7840 16720 7880 16730
rect 7920 16910 7960 16920
rect 7920 16890 7930 16910
rect 7950 16890 7960 16910
rect 7920 16750 7960 16890
rect 7920 16730 7930 16750
rect 7950 16730 7960 16750
rect 7920 16720 7960 16730
rect 8000 16910 8040 16920
rect 8000 16890 8010 16910
rect 8030 16890 8040 16910
rect 8000 16750 8040 16890
rect 8000 16730 8010 16750
rect 8030 16730 8040 16750
rect 8000 16720 8040 16730
rect 8080 16910 8120 16920
rect 8080 16890 8090 16910
rect 8110 16890 8120 16910
rect 8080 16750 8120 16890
rect 8080 16730 8090 16750
rect 8110 16730 8120 16750
rect 8080 16720 8120 16730
rect 8160 16910 8200 16920
rect 8160 16890 8170 16910
rect 8190 16890 8200 16910
rect 8160 16750 8200 16890
rect 8160 16730 8170 16750
rect 8190 16730 8200 16750
rect 8160 16720 8200 16730
rect 8240 16910 8280 16920
rect 8240 16890 8250 16910
rect 8270 16890 8280 16910
rect 8240 16750 8280 16890
rect 8240 16730 8250 16750
rect 8270 16730 8280 16750
rect 8240 16720 8280 16730
rect 8320 16910 8360 16920
rect 8320 16890 8330 16910
rect 8350 16890 8360 16910
rect 8320 16750 8360 16890
rect 8320 16730 8330 16750
rect 8350 16730 8360 16750
rect 8320 16720 8360 16730
rect 8400 16910 8440 16920
rect 8400 16890 8410 16910
rect 8430 16890 8440 16910
rect 8400 16750 8440 16890
rect 8400 16730 8410 16750
rect 8430 16730 8440 16750
rect 8400 16720 8440 16730
rect 8480 16910 8520 16920
rect 8480 16890 8490 16910
rect 8510 16890 8520 16910
rect 8480 16750 8520 16890
rect 8480 16730 8490 16750
rect 8510 16730 8520 16750
rect 8480 16720 8520 16730
rect 8560 16910 8600 16920
rect 8560 16890 8570 16910
rect 8590 16890 8600 16910
rect 8560 16750 8600 16890
rect 8560 16730 8570 16750
rect 8590 16730 8600 16750
rect 8560 16720 8600 16730
rect 8640 16910 8680 16920
rect 8640 16890 8650 16910
rect 8670 16890 8680 16910
rect 8640 16750 8680 16890
rect 8640 16730 8650 16750
rect 8670 16730 8680 16750
rect 8640 16720 8680 16730
rect 8720 16910 8760 16920
rect 8720 16890 8730 16910
rect 8750 16890 8760 16910
rect 8720 16750 8760 16890
rect 8720 16730 8730 16750
rect 8750 16730 8760 16750
rect 8720 16720 8760 16730
rect 8800 16910 8840 16920
rect 8800 16890 8810 16910
rect 8830 16890 8840 16910
rect 8800 16750 8840 16890
rect 8800 16730 8810 16750
rect 8830 16730 8840 16750
rect 8800 16720 8840 16730
rect 8880 16910 8920 16920
rect 8880 16890 8890 16910
rect 8910 16890 8920 16910
rect 8880 16750 8920 16890
rect 8880 16730 8890 16750
rect 8910 16730 8920 16750
rect 8880 16720 8920 16730
rect 8960 16910 9000 16920
rect 8960 16890 8970 16910
rect 8990 16890 9000 16910
rect 8960 16750 9000 16890
rect 8960 16730 8970 16750
rect 8990 16730 9000 16750
rect 8960 16720 9000 16730
rect 9040 16910 9080 16920
rect 9040 16890 9050 16910
rect 9070 16890 9080 16910
rect 9040 16750 9080 16890
rect 9040 16730 9050 16750
rect 9070 16730 9080 16750
rect 9040 16720 9080 16730
rect 9120 16910 9160 16920
rect 9120 16890 9130 16910
rect 9150 16890 9160 16910
rect 9120 16750 9160 16890
rect 9120 16730 9130 16750
rect 9150 16730 9160 16750
rect 9120 16720 9160 16730
rect 9200 16910 9240 16920
rect 9200 16890 9210 16910
rect 9230 16890 9240 16910
rect 9200 16750 9240 16890
rect 9200 16730 9210 16750
rect 9230 16730 9240 16750
rect 9200 16720 9240 16730
rect 9280 16910 9320 16920
rect 9280 16890 9290 16910
rect 9310 16890 9320 16910
rect 9280 16750 9320 16890
rect 9280 16730 9290 16750
rect 9310 16730 9320 16750
rect 9280 16720 9320 16730
rect 9360 16910 9400 16920
rect 9360 16890 9370 16910
rect 9390 16890 9400 16910
rect 9360 16750 9400 16890
rect 9360 16730 9370 16750
rect 9390 16730 9400 16750
rect 9360 16720 9400 16730
rect 9440 16910 9480 16920
rect 9440 16890 9450 16910
rect 9470 16890 9480 16910
rect 9440 16750 9480 16890
rect 9440 16730 9450 16750
rect 9470 16730 9480 16750
rect 9440 16720 9480 16730
rect 9520 16720 9560 16920
rect 9600 16720 9640 16920
rect 9680 16720 9720 16920
rect 9760 16720 9800 16920
rect 9840 16720 9880 16920
rect 9920 16720 9960 16920
rect 10000 16720 10040 16920
rect 10080 16720 10120 16920
rect 10160 16720 10200 16920
rect 10240 16720 10280 16920
rect 10320 16720 10360 16920
rect 10400 16720 10440 16920
rect 10480 16720 10520 16920
rect 10560 16720 10600 16920
rect 10640 16720 10680 16920
rect 10720 16720 10760 16920
rect 10800 16720 10840 16920
rect 10880 16720 10920 16920
rect 10960 16720 11000 16920
rect 11040 16720 11080 16920
rect 11120 16720 11160 16920
rect 11200 16720 11240 16920
rect 11280 16720 11320 16920
rect 11360 16720 11400 16920
rect 11440 16720 11480 16920
rect 11560 16910 11600 16920
rect 11560 16890 11570 16910
rect 11590 16890 11600 16910
rect 11560 16750 11600 16890
rect 11560 16730 11570 16750
rect 11590 16730 11600 16750
rect 11560 16720 11600 16730
rect 11640 16910 11680 16920
rect 11640 16890 11650 16910
rect 11670 16890 11680 16910
rect 11640 16750 11680 16890
rect 11640 16730 11650 16750
rect 11670 16730 11680 16750
rect 11640 16720 11680 16730
rect 11720 16910 11760 16920
rect 11720 16890 11730 16910
rect 11750 16890 11760 16910
rect 11720 16750 11760 16890
rect 11720 16730 11730 16750
rect 11750 16730 11760 16750
rect 11720 16720 11760 16730
rect 11800 16910 11840 16920
rect 11800 16890 11810 16910
rect 11830 16890 11840 16910
rect 11800 16750 11840 16890
rect 11800 16730 11810 16750
rect 11830 16730 11840 16750
rect 11800 16720 11840 16730
rect 11880 16910 11920 16920
rect 11880 16890 11890 16910
rect 11910 16890 11920 16910
rect 11880 16750 11920 16890
rect 11880 16730 11890 16750
rect 11910 16730 11920 16750
rect 11880 16720 11920 16730
rect 11960 16910 12000 16920
rect 11960 16890 11970 16910
rect 11990 16890 12000 16910
rect 11960 16750 12000 16890
rect 11960 16730 11970 16750
rect 11990 16730 12000 16750
rect 11960 16720 12000 16730
rect 12040 16910 12080 16920
rect 12040 16890 12050 16910
rect 12070 16890 12080 16910
rect 12040 16750 12080 16890
rect 12040 16730 12050 16750
rect 12070 16730 12080 16750
rect 12040 16720 12080 16730
rect 12120 16910 12160 16920
rect 12120 16890 12130 16910
rect 12150 16890 12160 16910
rect 12120 16750 12160 16890
rect 12120 16730 12130 16750
rect 12150 16730 12160 16750
rect 12120 16720 12160 16730
rect 12200 16910 12240 16920
rect 12200 16890 12210 16910
rect 12230 16890 12240 16910
rect 12200 16750 12240 16890
rect 12200 16730 12210 16750
rect 12230 16730 12240 16750
rect 12200 16720 12240 16730
rect 12280 16910 12320 16920
rect 12280 16890 12290 16910
rect 12310 16890 12320 16910
rect 12280 16750 12320 16890
rect 12280 16730 12290 16750
rect 12310 16730 12320 16750
rect 12280 16720 12320 16730
rect 12360 16910 12400 16920
rect 12360 16890 12370 16910
rect 12390 16890 12400 16910
rect 12360 16750 12400 16890
rect 12360 16730 12370 16750
rect 12390 16730 12400 16750
rect 12360 16720 12400 16730
rect 12440 16910 12480 16920
rect 12440 16890 12450 16910
rect 12470 16890 12480 16910
rect 12440 16750 12480 16890
rect 12440 16730 12450 16750
rect 12470 16730 12480 16750
rect 12440 16720 12480 16730
rect 12520 16910 12560 16920
rect 12520 16890 12530 16910
rect 12550 16890 12560 16910
rect 12520 16750 12560 16890
rect 12520 16730 12530 16750
rect 12550 16730 12560 16750
rect 12520 16720 12560 16730
rect 12600 16910 12640 16920
rect 12600 16890 12610 16910
rect 12630 16890 12640 16910
rect 12600 16750 12640 16890
rect 12600 16730 12610 16750
rect 12630 16730 12640 16750
rect 12600 16720 12640 16730
rect 12680 16910 12720 16920
rect 12680 16890 12690 16910
rect 12710 16890 12720 16910
rect 12680 16750 12720 16890
rect 12680 16730 12690 16750
rect 12710 16730 12720 16750
rect 12680 16720 12720 16730
rect 12760 16910 12800 16920
rect 12760 16890 12770 16910
rect 12790 16890 12800 16910
rect 12760 16750 12800 16890
rect 12760 16730 12770 16750
rect 12790 16730 12800 16750
rect 12760 16720 12800 16730
rect 12840 16910 12880 16920
rect 12840 16890 12850 16910
rect 12870 16890 12880 16910
rect 12840 16750 12880 16890
rect 12840 16730 12850 16750
rect 12870 16730 12880 16750
rect 12840 16720 12880 16730
rect 12920 16910 12960 16920
rect 12920 16890 12930 16910
rect 12950 16890 12960 16910
rect 12920 16750 12960 16890
rect 12920 16730 12930 16750
rect 12950 16730 12960 16750
rect 12920 16720 12960 16730
rect 13000 16910 13040 16920
rect 13000 16890 13010 16910
rect 13030 16890 13040 16910
rect 13000 16750 13040 16890
rect 13000 16730 13010 16750
rect 13030 16730 13040 16750
rect 13000 16720 13040 16730
rect 13080 16910 13120 16920
rect 13080 16890 13090 16910
rect 13110 16890 13120 16910
rect 13080 16750 13120 16890
rect 13080 16730 13090 16750
rect 13110 16730 13120 16750
rect 13080 16720 13120 16730
rect 13160 16910 13200 16920
rect 13160 16890 13170 16910
rect 13190 16890 13200 16910
rect 13160 16750 13200 16890
rect 13160 16730 13170 16750
rect 13190 16730 13200 16750
rect 13160 16720 13200 16730
rect 13240 16910 13280 16920
rect 13240 16890 13250 16910
rect 13270 16890 13280 16910
rect 13240 16750 13280 16890
rect 13240 16730 13250 16750
rect 13270 16730 13280 16750
rect 13240 16720 13280 16730
rect 13320 16910 13360 16920
rect 13320 16890 13330 16910
rect 13350 16890 13360 16910
rect 13320 16750 13360 16890
rect 13320 16730 13330 16750
rect 13350 16730 13360 16750
rect 13320 16720 13360 16730
rect 13400 16910 13440 16920
rect 13400 16890 13410 16910
rect 13430 16890 13440 16910
rect 13400 16750 13440 16890
rect 13400 16730 13410 16750
rect 13430 16730 13440 16750
rect 13400 16720 13440 16730
rect 13480 16910 13520 16920
rect 13480 16890 13490 16910
rect 13510 16890 13520 16910
rect 13480 16750 13520 16890
rect 13480 16730 13490 16750
rect 13510 16730 13520 16750
rect 13480 16720 13520 16730
rect 13560 16910 13600 16920
rect 13560 16890 13570 16910
rect 13590 16890 13600 16910
rect 13560 16750 13600 16890
rect 13560 16730 13570 16750
rect 13590 16730 13600 16750
rect 13560 16720 13600 16730
rect 13640 16910 13680 16920
rect 13640 16890 13650 16910
rect 13670 16890 13680 16910
rect 13640 16750 13680 16890
rect 13640 16730 13650 16750
rect 13670 16730 13680 16750
rect 13640 16720 13680 16730
rect 13720 16910 13760 16920
rect 13720 16890 13730 16910
rect 13750 16890 13760 16910
rect 13720 16750 13760 16890
rect 13720 16730 13730 16750
rect 13750 16730 13760 16750
rect 13720 16720 13760 16730
rect 13800 16910 13840 16920
rect 13800 16890 13810 16910
rect 13830 16890 13840 16910
rect 13800 16750 13840 16890
rect 13800 16730 13810 16750
rect 13830 16730 13840 16750
rect 13800 16720 13840 16730
rect 13880 16910 13920 16920
rect 13880 16890 13890 16910
rect 13910 16890 13920 16910
rect 13880 16750 13920 16890
rect 13880 16730 13890 16750
rect 13910 16730 13920 16750
rect 13880 16720 13920 16730
rect 13960 16910 14000 16920
rect 13960 16890 13970 16910
rect 13990 16890 14000 16910
rect 13960 16750 14000 16890
rect 13960 16730 13970 16750
rect 13990 16730 14000 16750
rect 13960 16720 14000 16730
rect 14040 16910 14080 16920
rect 14040 16890 14050 16910
rect 14070 16890 14080 16910
rect 14040 16750 14080 16890
rect 14040 16730 14050 16750
rect 14070 16730 14080 16750
rect 14040 16720 14080 16730
rect 14120 16910 14160 16920
rect 14120 16890 14130 16910
rect 14150 16890 14160 16910
rect 14120 16750 14160 16890
rect 14120 16730 14130 16750
rect 14150 16730 14160 16750
rect 14120 16720 14160 16730
rect 14200 16910 14240 16920
rect 14200 16890 14210 16910
rect 14230 16890 14240 16910
rect 14200 16750 14240 16890
rect 14200 16730 14210 16750
rect 14230 16730 14240 16750
rect 14200 16720 14240 16730
rect 14280 16910 14320 16920
rect 14280 16890 14290 16910
rect 14310 16890 14320 16910
rect 14280 16750 14320 16890
rect 14280 16730 14290 16750
rect 14310 16730 14320 16750
rect 14280 16720 14320 16730
rect 14360 16910 14400 16920
rect 14360 16890 14370 16910
rect 14390 16890 14400 16910
rect 14360 16750 14400 16890
rect 14360 16730 14370 16750
rect 14390 16730 14400 16750
rect 14360 16720 14400 16730
rect 14440 16910 14480 16920
rect 14440 16890 14450 16910
rect 14470 16890 14480 16910
rect 14440 16750 14480 16890
rect 14440 16730 14450 16750
rect 14470 16730 14480 16750
rect 14440 16720 14480 16730
rect 14520 16910 14560 16920
rect 14520 16890 14530 16910
rect 14550 16890 14560 16910
rect 14520 16750 14560 16890
rect 14520 16730 14530 16750
rect 14550 16730 14560 16750
rect 14520 16720 14560 16730
rect 14600 16910 14640 16920
rect 14600 16890 14610 16910
rect 14630 16890 14640 16910
rect 14600 16750 14640 16890
rect 14600 16730 14610 16750
rect 14630 16730 14640 16750
rect 14600 16720 14640 16730
rect 14680 16910 14720 16920
rect 14680 16890 14690 16910
rect 14710 16890 14720 16910
rect 14680 16750 14720 16890
rect 14680 16730 14690 16750
rect 14710 16730 14720 16750
rect 14680 16720 14720 16730
rect 14760 16720 14800 16920
rect 14840 16720 14880 16920
rect 14920 16720 14960 16920
rect 15000 16720 15040 16920
rect 15080 16720 15120 16920
rect 15160 16720 15200 16920
rect 15240 16720 15280 16920
rect 15320 16720 15360 16920
rect 15400 16720 15440 16920
rect 15480 16720 15520 16920
rect 15560 16720 15600 16920
rect 15640 16720 15680 16920
rect 15720 16720 15760 16920
rect 15800 16720 15840 16920
rect 15880 16720 15920 16920
rect 15960 16720 16000 16920
rect 16040 16720 16080 16920
rect 16120 16720 16160 16920
rect 16200 16720 16240 16920
rect 16280 16720 16320 16920
rect 16360 16720 16400 16920
rect 16440 16720 16480 16920
rect 16520 16720 16560 16920
rect 16600 16720 16640 16920
rect 16680 16720 16720 16920
rect 16760 16910 16800 16920
rect 16760 16890 16770 16910
rect 16790 16890 16800 16910
rect 16760 16750 16800 16890
rect 16760 16730 16770 16750
rect 16790 16730 16800 16750
rect 16760 16720 16800 16730
rect 16840 16910 16880 16920
rect 16840 16890 16850 16910
rect 16870 16890 16880 16910
rect 16840 16750 16880 16890
rect 16840 16730 16850 16750
rect 16870 16730 16880 16750
rect 16840 16720 16880 16730
rect 16920 16910 16960 16920
rect 16920 16890 16930 16910
rect 16950 16890 16960 16910
rect 16920 16750 16960 16890
rect 16920 16730 16930 16750
rect 16950 16730 16960 16750
rect 16920 16720 16960 16730
rect 17000 16910 17040 16920
rect 17000 16890 17010 16910
rect 17030 16890 17040 16910
rect 17000 16750 17040 16890
rect 17000 16730 17010 16750
rect 17030 16730 17040 16750
rect 17000 16720 17040 16730
rect 17080 16910 17120 16920
rect 17080 16890 17090 16910
rect 17110 16890 17120 16910
rect 17080 16750 17120 16890
rect 17080 16730 17090 16750
rect 17110 16730 17120 16750
rect 17080 16720 17120 16730
rect 17160 16910 17200 16920
rect 17160 16890 17170 16910
rect 17190 16890 17200 16910
rect 17160 16750 17200 16890
rect 17160 16730 17170 16750
rect 17190 16730 17200 16750
rect 17160 16720 17200 16730
rect 17240 16910 17280 16920
rect 17240 16890 17250 16910
rect 17270 16890 17280 16910
rect 17240 16750 17280 16890
rect 17240 16730 17250 16750
rect 17270 16730 17280 16750
rect 17240 16720 17280 16730
rect 17320 16910 17360 16920
rect 17320 16890 17330 16910
rect 17350 16890 17360 16910
rect 17320 16750 17360 16890
rect 17320 16730 17330 16750
rect 17350 16730 17360 16750
rect 17320 16720 17360 16730
rect 17400 16910 17440 16920
rect 17400 16890 17410 16910
rect 17430 16890 17440 16910
rect 17400 16750 17440 16890
rect 17400 16730 17410 16750
rect 17430 16730 17440 16750
rect 17400 16720 17440 16730
rect 17480 16910 17520 16920
rect 17480 16890 17490 16910
rect 17510 16890 17520 16910
rect 17480 16750 17520 16890
rect 17480 16730 17490 16750
rect 17510 16730 17520 16750
rect 17480 16720 17520 16730
rect 17560 16910 17600 16920
rect 17560 16890 17570 16910
rect 17590 16890 17600 16910
rect 17560 16750 17600 16890
rect 17560 16730 17570 16750
rect 17590 16730 17600 16750
rect 17560 16720 17600 16730
rect 17640 16910 17680 16920
rect 17640 16890 17650 16910
rect 17670 16890 17680 16910
rect 17640 16750 17680 16890
rect 17640 16730 17650 16750
rect 17670 16730 17680 16750
rect 17640 16720 17680 16730
rect 17720 16910 17760 16920
rect 17720 16890 17730 16910
rect 17750 16890 17760 16910
rect 17720 16750 17760 16890
rect 17720 16730 17730 16750
rect 17750 16730 17760 16750
rect 17720 16720 17760 16730
rect 17800 16910 17840 16920
rect 17800 16890 17810 16910
rect 17830 16890 17840 16910
rect 17800 16750 17840 16890
rect 17800 16730 17810 16750
rect 17830 16730 17840 16750
rect 17800 16720 17840 16730
rect 17880 16910 17920 16920
rect 17880 16890 17890 16910
rect 17910 16890 17920 16910
rect 17880 16750 17920 16890
rect 17880 16730 17890 16750
rect 17910 16730 17920 16750
rect 17880 16720 17920 16730
rect 17960 16910 18000 16920
rect 17960 16890 17970 16910
rect 17990 16890 18000 16910
rect 17960 16750 18000 16890
rect 17960 16730 17970 16750
rect 17990 16730 18000 16750
rect 17960 16720 18000 16730
rect 18040 16910 18080 16920
rect 18040 16890 18050 16910
rect 18070 16890 18080 16910
rect 18040 16750 18080 16890
rect 18040 16730 18050 16750
rect 18070 16730 18080 16750
rect 18040 16720 18080 16730
rect 18120 16910 18160 16920
rect 18120 16890 18130 16910
rect 18150 16890 18160 16910
rect 18120 16750 18160 16890
rect 18120 16730 18130 16750
rect 18150 16730 18160 16750
rect 18120 16720 18160 16730
rect 18200 16910 18240 16920
rect 18200 16890 18210 16910
rect 18230 16890 18240 16910
rect 18200 16750 18240 16890
rect 18200 16730 18210 16750
rect 18230 16730 18240 16750
rect 18200 16720 18240 16730
rect 18280 16910 18320 16920
rect 18280 16890 18290 16910
rect 18310 16890 18320 16910
rect 18280 16750 18320 16890
rect 18280 16730 18290 16750
rect 18310 16730 18320 16750
rect 18280 16720 18320 16730
rect 18360 16910 18400 16920
rect 18360 16890 18370 16910
rect 18390 16890 18400 16910
rect 18360 16750 18400 16890
rect 18360 16730 18370 16750
rect 18390 16730 18400 16750
rect 18360 16720 18400 16730
rect 18440 16910 18480 16920
rect 18440 16890 18450 16910
rect 18470 16890 18480 16910
rect 18440 16750 18480 16890
rect 18440 16730 18450 16750
rect 18470 16730 18480 16750
rect 18440 16720 18480 16730
rect 18520 16910 18560 16920
rect 18520 16890 18530 16910
rect 18550 16890 18560 16910
rect 18520 16750 18560 16890
rect 18520 16730 18530 16750
rect 18550 16730 18560 16750
rect 18520 16720 18560 16730
rect 18600 16910 18640 16920
rect 18600 16890 18610 16910
rect 18630 16890 18640 16910
rect 18600 16750 18640 16890
rect 18600 16730 18610 16750
rect 18630 16730 18640 16750
rect 18600 16720 18640 16730
rect 18680 16910 18720 16920
rect 18680 16890 18690 16910
rect 18710 16890 18720 16910
rect 18680 16750 18720 16890
rect 18680 16730 18690 16750
rect 18710 16730 18720 16750
rect 18680 16720 18720 16730
rect 18760 16910 18800 16920
rect 18760 16890 18770 16910
rect 18790 16890 18800 16910
rect 18760 16750 18800 16890
rect 18760 16730 18770 16750
rect 18790 16730 18800 16750
rect 18760 16720 18800 16730
rect 18840 16910 18880 16920
rect 18840 16890 18850 16910
rect 18870 16890 18880 16910
rect 18840 16750 18880 16890
rect 18840 16730 18850 16750
rect 18870 16730 18880 16750
rect 18840 16720 18880 16730
rect 18920 16910 18960 16920
rect 18920 16890 18930 16910
rect 18950 16890 18960 16910
rect 18920 16750 18960 16890
rect 18920 16730 18930 16750
rect 18950 16730 18960 16750
rect 18920 16720 18960 16730
rect 19000 16910 19040 16920
rect 19000 16890 19010 16910
rect 19030 16890 19040 16910
rect 19000 16750 19040 16890
rect 19000 16730 19010 16750
rect 19030 16730 19040 16750
rect 19000 16720 19040 16730
rect 19080 16910 19120 16920
rect 19080 16890 19090 16910
rect 19110 16890 19120 16910
rect 19080 16750 19120 16890
rect 19080 16730 19090 16750
rect 19110 16730 19120 16750
rect 19080 16720 19120 16730
rect 19160 16910 19200 16920
rect 19160 16890 19170 16910
rect 19190 16890 19200 16910
rect 19160 16750 19200 16890
rect 19160 16730 19170 16750
rect 19190 16730 19200 16750
rect 19160 16720 19200 16730
rect 19240 16910 19280 16920
rect 19240 16890 19250 16910
rect 19270 16890 19280 16910
rect 19240 16750 19280 16890
rect 19240 16730 19250 16750
rect 19270 16730 19280 16750
rect 19240 16720 19280 16730
rect 19320 16910 19360 16920
rect 19320 16890 19330 16910
rect 19350 16890 19360 16910
rect 19320 16750 19360 16890
rect 19320 16730 19330 16750
rect 19350 16730 19360 16750
rect 19320 16720 19360 16730
rect 19400 16910 19440 16920
rect 19400 16890 19410 16910
rect 19430 16890 19440 16910
rect 19400 16750 19440 16890
rect 19400 16730 19410 16750
rect 19430 16730 19440 16750
rect 19400 16720 19440 16730
rect 19480 16910 19520 16920
rect 19480 16890 19490 16910
rect 19510 16890 19520 16910
rect 19480 16750 19520 16890
rect 19480 16730 19490 16750
rect 19510 16730 19520 16750
rect 19480 16720 19520 16730
rect 19560 16910 19600 16920
rect 19560 16890 19570 16910
rect 19590 16890 19600 16910
rect 19560 16750 19600 16890
rect 19560 16730 19570 16750
rect 19590 16730 19600 16750
rect 19560 16720 19600 16730
rect 19640 16910 19680 16920
rect 19640 16890 19650 16910
rect 19670 16890 19680 16910
rect 19640 16750 19680 16890
rect 19640 16730 19650 16750
rect 19670 16730 19680 16750
rect 19640 16720 19680 16730
rect 19720 16910 19760 16920
rect 19720 16890 19730 16910
rect 19750 16890 19760 16910
rect 19720 16750 19760 16890
rect 19720 16730 19730 16750
rect 19750 16730 19760 16750
rect 19720 16720 19760 16730
rect 19800 16910 19840 16920
rect 19800 16890 19810 16910
rect 19830 16890 19840 16910
rect 19800 16750 19840 16890
rect 19800 16730 19810 16750
rect 19830 16730 19840 16750
rect 19800 16720 19840 16730
rect 19880 16910 19920 16920
rect 19880 16890 19890 16910
rect 19910 16890 19920 16910
rect 19880 16750 19920 16890
rect 19880 16730 19890 16750
rect 19910 16730 19920 16750
rect 19880 16720 19920 16730
rect 19960 16910 20000 16920
rect 19960 16890 19970 16910
rect 19990 16890 20000 16910
rect 19960 16750 20000 16890
rect 19960 16730 19970 16750
rect 19990 16730 20000 16750
rect 19960 16720 20000 16730
rect 20040 16910 20080 16920
rect 20040 16890 20050 16910
rect 20070 16890 20080 16910
rect 20040 16750 20080 16890
rect 20040 16730 20050 16750
rect 20070 16730 20080 16750
rect 20040 16720 20080 16730
rect 20120 16910 20160 16920
rect 20120 16890 20130 16910
rect 20150 16890 20160 16910
rect 20120 16750 20160 16890
rect 20120 16730 20130 16750
rect 20150 16730 20160 16750
rect 20120 16720 20160 16730
rect 20200 16910 20240 16920
rect 20200 16890 20210 16910
rect 20230 16890 20240 16910
rect 20200 16750 20240 16890
rect 20200 16730 20210 16750
rect 20230 16730 20240 16750
rect 20200 16720 20240 16730
rect 20280 16910 20320 16920
rect 20280 16890 20290 16910
rect 20310 16890 20320 16910
rect 20280 16750 20320 16890
rect 20280 16730 20290 16750
rect 20310 16730 20320 16750
rect 20280 16720 20320 16730
rect 20360 16910 20400 16920
rect 20360 16890 20370 16910
rect 20390 16890 20400 16910
rect 20360 16750 20400 16890
rect 20360 16730 20370 16750
rect 20390 16730 20400 16750
rect 20360 16720 20400 16730
rect 20440 16910 20480 16920
rect 20440 16890 20450 16910
rect 20470 16890 20480 16910
rect 20440 16750 20480 16890
rect 20440 16730 20450 16750
rect 20470 16730 20480 16750
rect 20440 16720 20480 16730
rect 20520 16910 20560 16920
rect 20520 16890 20530 16910
rect 20550 16890 20560 16910
rect 20520 16750 20560 16890
rect 20520 16730 20530 16750
rect 20550 16730 20560 16750
rect 20520 16720 20560 16730
rect 20600 16910 20640 16920
rect 20600 16890 20610 16910
rect 20630 16890 20640 16910
rect 20600 16750 20640 16890
rect 20600 16730 20610 16750
rect 20630 16730 20640 16750
rect 20600 16720 20640 16730
rect 20680 16910 20720 16920
rect 20680 16890 20690 16910
rect 20710 16890 20720 16910
rect 20680 16750 20720 16890
rect 20680 16730 20690 16750
rect 20710 16730 20720 16750
rect 20680 16720 20720 16730
rect 20760 16910 20800 16920
rect 20760 16890 20770 16910
rect 20790 16890 20800 16910
rect 20760 16750 20800 16890
rect 20760 16730 20770 16750
rect 20790 16730 20800 16750
rect 20760 16720 20800 16730
rect 20840 16910 20880 16920
rect 20840 16890 20850 16910
rect 20870 16890 20880 16910
rect 20840 16750 20880 16890
rect 20840 16730 20850 16750
rect 20870 16730 20880 16750
rect 20840 16720 20880 16730
rect 20920 16910 20960 16920
rect 20920 16890 20930 16910
rect 20950 16890 20960 16910
rect 20920 16750 20960 16890
rect 20920 16730 20930 16750
rect 20950 16730 20960 16750
rect 20920 16720 20960 16730
rect 0 16670 40 16680
rect 0 16650 10 16670
rect 30 16650 40 16670
rect 0 16510 40 16650
rect 0 16490 10 16510
rect 30 16490 40 16510
rect 0 16480 40 16490
rect 80 16670 120 16680
rect 80 16650 90 16670
rect 110 16650 120 16670
rect 80 16510 120 16650
rect 80 16490 90 16510
rect 110 16490 120 16510
rect 80 16480 120 16490
rect 160 16670 200 16680
rect 160 16650 170 16670
rect 190 16650 200 16670
rect 160 16510 200 16650
rect 160 16490 170 16510
rect 190 16490 200 16510
rect 160 16480 200 16490
rect 240 16670 280 16680
rect 240 16650 250 16670
rect 270 16650 280 16670
rect 240 16510 280 16650
rect 240 16490 250 16510
rect 270 16490 280 16510
rect 240 16480 280 16490
rect 320 16670 360 16680
rect 320 16650 330 16670
rect 350 16650 360 16670
rect 320 16510 360 16650
rect 320 16490 330 16510
rect 350 16490 360 16510
rect 320 16480 360 16490
rect 400 16670 440 16680
rect 400 16650 410 16670
rect 430 16650 440 16670
rect 400 16510 440 16650
rect 400 16490 410 16510
rect 430 16490 440 16510
rect 400 16480 440 16490
rect 480 16670 520 16680
rect 480 16650 490 16670
rect 510 16650 520 16670
rect 480 16510 520 16650
rect 480 16490 490 16510
rect 510 16490 520 16510
rect 480 16480 520 16490
rect 560 16670 600 16680
rect 560 16650 570 16670
rect 590 16650 600 16670
rect 560 16510 600 16650
rect 560 16490 570 16510
rect 590 16490 600 16510
rect 560 16480 600 16490
rect 640 16670 680 16680
rect 640 16650 650 16670
rect 670 16650 680 16670
rect 640 16510 680 16650
rect 640 16490 650 16510
rect 670 16490 680 16510
rect 640 16480 680 16490
rect 720 16670 760 16680
rect 720 16650 730 16670
rect 750 16650 760 16670
rect 720 16510 760 16650
rect 720 16490 730 16510
rect 750 16490 760 16510
rect 720 16480 760 16490
rect 800 16670 840 16680
rect 800 16650 810 16670
rect 830 16650 840 16670
rect 800 16510 840 16650
rect 800 16490 810 16510
rect 830 16490 840 16510
rect 800 16480 840 16490
rect 880 16670 920 16680
rect 880 16650 890 16670
rect 910 16650 920 16670
rect 880 16510 920 16650
rect 880 16490 890 16510
rect 910 16490 920 16510
rect 880 16480 920 16490
rect 960 16670 1000 16680
rect 960 16650 970 16670
rect 990 16650 1000 16670
rect 960 16510 1000 16650
rect 960 16490 970 16510
rect 990 16490 1000 16510
rect 960 16480 1000 16490
rect 1040 16670 1080 16680
rect 1040 16650 1050 16670
rect 1070 16650 1080 16670
rect 1040 16510 1080 16650
rect 1040 16490 1050 16510
rect 1070 16490 1080 16510
rect 1040 16480 1080 16490
rect 1120 16670 1160 16680
rect 1120 16650 1130 16670
rect 1150 16650 1160 16670
rect 1120 16510 1160 16650
rect 1120 16490 1130 16510
rect 1150 16490 1160 16510
rect 1120 16480 1160 16490
rect 1200 16670 1240 16680
rect 1200 16650 1210 16670
rect 1230 16650 1240 16670
rect 1200 16510 1240 16650
rect 1200 16490 1210 16510
rect 1230 16490 1240 16510
rect 1200 16480 1240 16490
rect 1280 16670 1320 16680
rect 1280 16650 1290 16670
rect 1310 16650 1320 16670
rect 1280 16510 1320 16650
rect 1280 16490 1290 16510
rect 1310 16490 1320 16510
rect 1280 16480 1320 16490
rect 1360 16670 1400 16680
rect 1360 16650 1370 16670
rect 1390 16650 1400 16670
rect 1360 16510 1400 16650
rect 1360 16490 1370 16510
rect 1390 16490 1400 16510
rect 1360 16480 1400 16490
rect 1440 16670 1480 16680
rect 1440 16650 1450 16670
rect 1470 16650 1480 16670
rect 1440 16510 1480 16650
rect 1440 16490 1450 16510
rect 1470 16490 1480 16510
rect 1440 16480 1480 16490
rect 1520 16670 1560 16680
rect 1520 16650 1530 16670
rect 1550 16650 1560 16670
rect 1520 16510 1560 16650
rect 1520 16490 1530 16510
rect 1550 16490 1560 16510
rect 1520 16480 1560 16490
rect 1600 16670 1640 16680
rect 1600 16650 1610 16670
rect 1630 16650 1640 16670
rect 1600 16510 1640 16650
rect 1600 16490 1610 16510
rect 1630 16490 1640 16510
rect 1600 16480 1640 16490
rect 1680 16670 1720 16680
rect 1680 16650 1690 16670
rect 1710 16650 1720 16670
rect 1680 16510 1720 16650
rect 1680 16490 1690 16510
rect 1710 16490 1720 16510
rect 1680 16480 1720 16490
rect 1760 16670 1800 16680
rect 1760 16650 1770 16670
rect 1790 16650 1800 16670
rect 1760 16510 1800 16650
rect 1760 16490 1770 16510
rect 1790 16490 1800 16510
rect 1760 16480 1800 16490
rect 1840 16670 1880 16680
rect 1840 16650 1850 16670
rect 1870 16650 1880 16670
rect 1840 16510 1880 16650
rect 1840 16490 1850 16510
rect 1870 16490 1880 16510
rect 1840 16480 1880 16490
rect 1920 16670 1960 16680
rect 1920 16650 1930 16670
rect 1950 16650 1960 16670
rect 1920 16510 1960 16650
rect 1920 16490 1930 16510
rect 1950 16490 1960 16510
rect 1920 16480 1960 16490
rect 2000 16670 2040 16680
rect 2000 16650 2010 16670
rect 2030 16650 2040 16670
rect 2000 16510 2040 16650
rect 2000 16490 2010 16510
rect 2030 16490 2040 16510
rect 2000 16480 2040 16490
rect 2080 16670 2120 16680
rect 2080 16650 2090 16670
rect 2110 16650 2120 16670
rect 2080 16510 2120 16650
rect 2080 16490 2090 16510
rect 2110 16490 2120 16510
rect 2080 16480 2120 16490
rect 2160 16670 2200 16680
rect 2160 16650 2170 16670
rect 2190 16650 2200 16670
rect 2160 16510 2200 16650
rect 2160 16490 2170 16510
rect 2190 16490 2200 16510
rect 2160 16480 2200 16490
rect 2240 16670 2280 16680
rect 2240 16650 2250 16670
rect 2270 16650 2280 16670
rect 2240 16510 2280 16650
rect 2240 16490 2250 16510
rect 2270 16490 2280 16510
rect 2240 16480 2280 16490
rect 2320 16670 2360 16680
rect 2320 16650 2330 16670
rect 2350 16650 2360 16670
rect 2320 16510 2360 16650
rect 2320 16490 2330 16510
rect 2350 16490 2360 16510
rect 2320 16480 2360 16490
rect 2400 16670 2440 16680
rect 2400 16650 2410 16670
rect 2430 16650 2440 16670
rect 2400 16510 2440 16650
rect 2400 16490 2410 16510
rect 2430 16490 2440 16510
rect 2400 16480 2440 16490
rect 2480 16670 2520 16680
rect 2480 16650 2490 16670
rect 2510 16650 2520 16670
rect 2480 16510 2520 16650
rect 2480 16490 2490 16510
rect 2510 16490 2520 16510
rect 2480 16480 2520 16490
rect 2560 16670 2600 16680
rect 2560 16650 2570 16670
rect 2590 16650 2600 16670
rect 2560 16510 2600 16650
rect 2560 16490 2570 16510
rect 2590 16490 2600 16510
rect 2560 16480 2600 16490
rect 2640 16670 2680 16680
rect 2640 16650 2650 16670
rect 2670 16650 2680 16670
rect 2640 16510 2680 16650
rect 2640 16490 2650 16510
rect 2670 16490 2680 16510
rect 2640 16480 2680 16490
rect 2720 16670 2760 16680
rect 2720 16650 2730 16670
rect 2750 16650 2760 16670
rect 2720 16510 2760 16650
rect 2720 16490 2730 16510
rect 2750 16490 2760 16510
rect 2720 16480 2760 16490
rect 2800 16670 2840 16680
rect 2800 16650 2810 16670
rect 2830 16650 2840 16670
rect 2800 16510 2840 16650
rect 2800 16490 2810 16510
rect 2830 16490 2840 16510
rect 2800 16480 2840 16490
rect 2880 16670 2920 16680
rect 2880 16650 2890 16670
rect 2910 16650 2920 16670
rect 2880 16510 2920 16650
rect 2880 16490 2890 16510
rect 2910 16490 2920 16510
rect 2880 16480 2920 16490
rect 2960 16670 3000 16680
rect 2960 16650 2970 16670
rect 2990 16650 3000 16670
rect 2960 16510 3000 16650
rect 2960 16490 2970 16510
rect 2990 16490 3000 16510
rect 2960 16480 3000 16490
rect 3040 16670 3080 16680
rect 3040 16650 3050 16670
rect 3070 16650 3080 16670
rect 3040 16510 3080 16650
rect 3040 16490 3050 16510
rect 3070 16490 3080 16510
rect 3040 16480 3080 16490
rect 3120 16670 3160 16680
rect 3120 16650 3130 16670
rect 3150 16650 3160 16670
rect 3120 16510 3160 16650
rect 3120 16490 3130 16510
rect 3150 16490 3160 16510
rect 3120 16480 3160 16490
rect 3200 16670 3240 16680
rect 3200 16650 3210 16670
rect 3230 16650 3240 16670
rect 3200 16510 3240 16650
rect 3200 16490 3210 16510
rect 3230 16490 3240 16510
rect 3200 16480 3240 16490
rect 3280 16670 3320 16680
rect 3280 16650 3290 16670
rect 3310 16650 3320 16670
rect 3280 16510 3320 16650
rect 3280 16490 3290 16510
rect 3310 16490 3320 16510
rect 3280 16480 3320 16490
rect 3360 16670 3400 16680
rect 3360 16650 3370 16670
rect 3390 16650 3400 16670
rect 3360 16510 3400 16650
rect 3360 16490 3370 16510
rect 3390 16490 3400 16510
rect 3360 16480 3400 16490
rect 3440 16670 3480 16680
rect 3440 16650 3450 16670
rect 3470 16650 3480 16670
rect 3440 16510 3480 16650
rect 3440 16490 3450 16510
rect 3470 16490 3480 16510
rect 3440 16480 3480 16490
rect 3520 16670 3560 16680
rect 3520 16650 3530 16670
rect 3550 16650 3560 16670
rect 3520 16510 3560 16650
rect 3520 16490 3530 16510
rect 3550 16490 3560 16510
rect 3520 16480 3560 16490
rect 3600 16670 3640 16680
rect 3600 16650 3610 16670
rect 3630 16650 3640 16670
rect 3600 16510 3640 16650
rect 3600 16490 3610 16510
rect 3630 16490 3640 16510
rect 3600 16480 3640 16490
rect 3680 16670 3720 16680
rect 3680 16650 3690 16670
rect 3710 16650 3720 16670
rect 3680 16510 3720 16650
rect 3680 16490 3690 16510
rect 3710 16490 3720 16510
rect 3680 16480 3720 16490
rect 3760 16670 3800 16680
rect 3760 16650 3770 16670
rect 3790 16650 3800 16670
rect 3760 16510 3800 16650
rect 3760 16490 3770 16510
rect 3790 16490 3800 16510
rect 3760 16480 3800 16490
rect 3840 16670 3880 16680
rect 3840 16650 3850 16670
rect 3870 16650 3880 16670
rect 3840 16510 3880 16650
rect 3840 16490 3850 16510
rect 3870 16490 3880 16510
rect 3840 16480 3880 16490
rect 3920 16670 3960 16680
rect 3920 16650 3930 16670
rect 3950 16650 3960 16670
rect 3920 16510 3960 16650
rect 3920 16490 3930 16510
rect 3950 16490 3960 16510
rect 3920 16480 3960 16490
rect 4000 16670 4040 16680
rect 4000 16650 4010 16670
rect 4030 16650 4040 16670
rect 4000 16510 4040 16650
rect 4000 16490 4010 16510
rect 4030 16490 4040 16510
rect 4000 16480 4040 16490
rect 4080 16670 4120 16680
rect 4080 16650 4090 16670
rect 4110 16650 4120 16670
rect 4080 16510 4120 16650
rect 4080 16490 4090 16510
rect 4110 16490 4120 16510
rect 4080 16480 4120 16490
rect 4160 16670 4200 16680
rect 4160 16650 4170 16670
rect 4190 16650 4200 16670
rect 4160 16510 4200 16650
rect 4160 16490 4170 16510
rect 4190 16490 4200 16510
rect 4160 16480 4200 16490
rect 4240 16480 4280 16680
rect 4320 16480 4360 16680
rect 4400 16480 4440 16680
rect 4480 16480 4520 16680
rect 4560 16480 4600 16680
rect 4640 16480 4680 16680
rect 4720 16480 4760 16680
rect 4800 16480 4840 16680
rect 4880 16480 4920 16680
rect 4960 16480 5000 16680
rect 5040 16480 5080 16680
rect 5120 16480 5160 16680
rect 5200 16480 5240 16680
rect 5280 16480 5320 16680
rect 5360 16480 5400 16680
rect 5440 16480 5480 16680
rect 5520 16480 5560 16680
rect 5600 16480 5640 16680
rect 5680 16480 5720 16680
rect 5760 16480 5800 16680
rect 5840 16480 5880 16680
rect 5920 16480 5960 16680
rect 6000 16480 6040 16680
rect 6080 16480 6120 16680
rect 6160 16480 6200 16680
rect 6240 16670 6280 16680
rect 6240 16650 6250 16670
rect 6270 16650 6280 16670
rect 6240 16510 6280 16650
rect 6240 16490 6250 16510
rect 6270 16490 6280 16510
rect 6240 16480 6280 16490
rect 6320 16670 6360 16680
rect 6320 16650 6330 16670
rect 6350 16650 6360 16670
rect 6320 16510 6360 16650
rect 6320 16490 6330 16510
rect 6350 16490 6360 16510
rect 6320 16480 6360 16490
rect 6400 16670 6440 16680
rect 6400 16650 6410 16670
rect 6430 16650 6440 16670
rect 6400 16510 6440 16650
rect 6400 16490 6410 16510
rect 6430 16490 6440 16510
rect 6400 16480 6440 16490
rect 6480 16670 6520 16680
rect 6480 16650 6490 16670
rect 6510 16650 6520 16670
rect 6480 16510 6520 16650
rect 6480 16490 6490 16510
rect 6510 16490 6520 16510
rect 6480 16480 6520 16490
rect 6560 16670 6600 16680
rect 6560 16650 6570 16670
rect 6590 16650 6600 16670
rect 6560 16510 6600 16650
rect 6560 16490 6570 16510
rect 6590 16490 6600 16510
rect 6560 16480 6600 16490
rect 6640 16670 6680 16680
rect 6640 16650 6650 16670
rect 6670 16650 6680 16670
rect 6640 16510 6680 16650
rect 6640 16490 6650 16510
rect 6670 16490 6680 16510
rect 6640 16480 6680 16490
rect 6720 16670 6760 16680
rect 6720 16650 6730 16670
rect 6750 16650 6760 16670
rect 6720 16510 6760 16650
rect 6720 16490 6730 16510
rect 6750 16490 6760 16510
rect 6720 16480 6760 16490
rect 6800 16670 6840 16680
rect 6800 16650 6810 16670
rect 6830 16650 6840 16670
rect 6800 16510 6840 16650
rect 6800 16490 6810 16510
rect 6830 16490 6840 16510
rect 6800 16480 6840 16490
rect 6880 16670 6920 16680
rect 6880 16650 6890 16670
rect 6910 16650 6920 16670
rect 6880 16510 6920 16650
rect 6880 16490 6890 16510
rect 6910 16490 6920 16510
rect 6880 16480 6920 16490
rect 6960 16670 7000 16680
rect 6960 16650 6970 16670
rect 6990 16650 7000 16670
rect 6960 16510 7000 16650
rect 6960 16490 6970 16510
rect 6990 16490 7000 16510
rect 6960 16480 7000 16490
rect 7040 16670 7080 16680
rect 7040 16650 7050 16670
rect 7070 16650 7080 16670
rect 7040 16510 7080 16650
rect 7040 16490 7050 16510
rect 7070 16490 7080 16510
rect 7040 16480 7080 16490
rect 7120 16670 7160 16680
rect 7120 16650 7130 16670
rect 7150 16650 7160 16670
rect 7120 16510 7160 16650
rect 7120 16490 7130 16510
rect 7150 16490 7160 16510
rect 7120 16480 7160 16490
rect 7200 16670 7240 16680
rect 7200 16650 7210 16670
rect 7230 16650 7240 16670
rect 7200 16510 7240 16650
rect 7200 16490 7210 16510
rect 7230 16490 7240 16510
rect 7200 16480 7240 16490
rect 7280 16670 7320 16680
rect 7280 16650 7290 16670
rect 7310 16650 7320 16670
rect 7280 16510 7320 16650
rect 7280 16490 7290 16510
rect 7310 16490 7320 16510
rect 7280 16480 7320 16490
rect 7360 16670 7400 16680
rect 7360 16650 7370 16670
rect 7390 16650 7400 16670
rect 7360 16510 7400 16650
rect 7360 16490 7370 16510
rect 7390 16490 7400 16510
rect 7360 16480 7400 16490
rect 7440 16670 7480 16680
rect 7440 16650 7450 16670
rect 7470 16650 7480 16670
rect 7440 16510 7480 16650
rect 7440 16490 7450 16510
rect 7470 16490 7480 16510
rect 7440 16480 7480 16490
rect 7520 16670 7560 16680
rect 7520 16650 7530 16670
rect 7550 16650 7560 16670
rect 7520 16510 7560 16650
rect 7520 16490 7530 16510
rect 7550 16490 7560 16510
rect 7520 16480 7560 16490
rect 7600 16670 7640 16680
rect 7600 16650 7610 16670
rect 7630 16650 7640 16670
rect 7600 16510 7640 16650
rect 7600 16490 7610 16510
rect 7630 16490 7640 16510
rect 7600 16480 7640 16490
rect 7680 16670 7720 16680
rect 7680 16650 7690 16670
rect 7710 16650 7720 16670
rect 7680 16510 7720 16650
rect 7680 16490 7690 16510
rect 7710 16490 7720 16510
rect 7680 16480 7720 16490
rect 7760 16670 7800 16680
rect 7760 16650 7770 16670
rect 7790 16650 7800 16670
rect 7760 16510 7800 16650
rect 7760 16490 7770 16510
rect 7790 16490 7800 16510
rect 7760 16480 7800 16490
rect 7840 16670 7880 16680
rect 7840 16650 7850 16670
rect 7870 16650 7880 16670
rect 7840 16510 7880 16650
rect 7840 16490 7850 16510
rect 7870 16490 7880 16510
rect 7840 16480 7880 16490
rect 7920 16670 7960 16680
rect 7920 16650 7930 16670
rect 7950 16650 7960 16670
rect 7920 16510 7960 16650
rect 7920 16490 7930 16510
rect 7950 16490 7960 16510
rect 7920 16480 7960 16490
rect 8000 16670 8040 16680
rect 8000 16650 8010 16670
rect 8030 16650 8040 16670
rect 8000 16510 8040 16650
rect 8000 16490 8010 16510
rect 8030 16490 8040 16510
rect 8000 16480 8040 16490
rect 8080 16670 8120 16680
rect 8080 16650 8090 16670
rect 8110 16650 8120 16670
rect 8080 16510 8120 16650
rect 8080 16490 8090 16510
rect 8110 16490 8120 16510
rect 8080 16480 8120 16490
rect 8160 16670 8200 16680
rect 8160 16650 8170 16670
rect 8190 16650 8200 16670
rect 8160 16510 8200 16650
rect 8160 16490 8170 16510
rect 8190 16490 8200 16510
rect 8160 16480 8200 16490
rect 8240 16670 8280 16680
rect 8240 16650 8250 16670
rect 8270 16650 8280 16670
rect 8240 16510 8280 16650
rect 8240 16490 8250 16510
rect 8270 16490 8280 16510
rect 8240 16480 8280 16490
rect 8320 16670 8360 16680
rect 8320 16650 8330 16670
rect 8350 16650 8360 16670
rect 8320 16510 8360 16650
rect 8320 16490 8330 16510
rect 8350 16490 8360 16510
rect 8320 16480 8360 16490
rect 8400 16670 8440 16680
rect 8400 16650 8410 16670
rect 8430 16650 8440 16670
rect 8400 16510 8440 16650
rect 8400 16490 8410 16510
rect 8430 16490 8440 16510
rect 8400 16480 8440 16490
rect 8480 16670 8520 16680
rect 8480 16650 8490 16670
rect 8510 16650 8520 16670
rect 8480 16510 8520 16650
rect 8480 16490 8490 16510
rect 8510 16490 8520 16510
rect 8480 16480 8520 16490
rect 8560 16670 8600 16680
rect 8560 16650 8570 16670
rect 8590 16650 8600 16670
rect 8560 16510 8600 16650
rect 8560 16490 8570 16510
rect 8590 16490 8600 16510
rect 8560 16480 8600 16490
rect 8640 16670 8680 16680
rect 8640 16650 8650 16670
rect 8670 16650 8680 16670
rect 8640 16510 8680 16650
rect 8640 16490 8650 16510
rect 8670 16490 8680 16510
rect 8640 16480 8680 16490
rect 8720 16670 8760 16680
rect 8720 16650 8730 16670
rect 8750 16650 8760 16670
rect 8720 16510 8760 16650
rect 8720 16490 8730 16510
rect 8750 16490 8760 16510
rect 8720 16480 8760 16490
rect 8800 16670 8840 16680
rect 8800 16650 8810 16670
rect 8830 16650 8840 16670
rect 8800 16510 8840 16650
rect 8800 16490 8810 16510
rect 8830 16490 8840 16510
rect 8800 16480 8840 16490
rect 8880 16670 8920 16680
rect 8880 16650 8890 16670
rect 8910 16650 8920 16670
rect 8880 16510 8920 16650
rect 8880 16490 8890 16510
rect 8910 16490 8920 16510
rect 8880 16480 8920 16490
rect 8960 16670 9000 16680
rect 8960 16650 8970 16670
rect 8990 16650 9000 16670
rect 8960 16510 9000 16650
rect 8960 16490 8970 16510
rect 8990 16490 9000 16510
rect 8960 16480 9000 16490
rect 9040 16670 9080 16680
rect 9040 16650 9050 16670
rect 9070 16650 9080 16670
rect 9040 16510 9080 16650
rect 9040 16490 9050 16510
rect 9070 16490 9080 16510
rect 9040 16480 9080 16490
rect 9120 16670 9160 16680
rect 9120 16650 9130 16670
rect 9150 16650 9160 16670
rect 9120 16510 9160 16650
rect 9120 16490 9130 16510
rect 9150 16490 9160 16510
rect 9120 16480 9160 16490
rect 9200 16670 9240 16680
rect 9200 16650 9210 16670
rect 9230 16650 9240 16670
rect 9200 16510 9240 16650
rect 9200 16490 9210 16510
rect 9230 16490 9240 16510
rect 9200 16480 9240 16490
rect 9280 16670 9320 16680
rect 9280 16650 9290 16670
rect 9310 16650 9320 16670
rect 9280 16510 9320 16650
rect 9280 16490 9290 16510
rect 9310 16490 9320 16510
rect 9280 16480 9320 16490
rect 9360 16670 9400 16680
rect 9360 16650 9370 16670
rect 9390 16650 9400 16670
rect 9360 16510 9400 16650
rect 9360 16490 9370 16510
rect 9390 16490 9400 16510
rect 9360 16480 9400 16490
rect 9440 16670 9480 16680
rect 9440 16650 9450 16670
rect 9470 16650 9480 16670
rect 9440 16510 9480 16650
rect 9440 16490 9450 16510
rect 9470 16490 9480 16510
rect 9440 16480 9480 16490
rect 9520 16480 9560 16680
rect 9600 16480 9640 16680
rect 9680 16480 9720 16680
rect 9760 16480 9800 16680
rect 9840 16480 9880 16680
rect 9920 16480 9960 16680
rect 10000 16480 10040 16680
rect 10080 16480 10120 16680
rect 10160 16480 10200 16680
rect 10240 16480 10280 16680
rect 10320 16480 10360 16680
rect 10400 16480 10440 16680
rect 10480 16480 10520 16680
rect 10560 16480 10600 16680
rect 10640 16480 10680 16680
rect 10720 16480 10760 16680
rect 10800 16480 10840 16680
rect 10880 16480 10920 16680
rect 10960 16480 11000 16680
rect 11040 16480 11080 16680
rect 11120 16480 11160 16680
rect 11200 16480 11240 16680
rect 11280 16480 11320 16680
rect 11360 16480 11400 16680
rect 11440 16480 11480 16680
rect 11560 16670 11600 16680
rect 11560 16650 11570 16670
rect 11590 16650 11600 16670
rect 11560 16510 11600 16650
rect 11560 16490 11570 16510
rect 11590 16490 11600 16510
rect 11560 16480 11600 16490
rect 11640 16670 11680 16680
rect 11640 16650 11650 16670
rect 11670 16650 11680 16670
rect 11640 16510 11680 16650
rect 11640 16490 11650 16510
rect 11670 16490 11680 16510
rect 11640 16480 11680 16490
rect 11720 16670 11760 16680
rect 11720 16650 11730 16670
rect 11750 16650 11760 16670
rect 11720 16510 11760 16650
rect 11720 16490 11730 16510
rect 11750 16490 11760 16510
rect 11720 16480 11760 16490
rect 11800 16670 11840 16680
rect 11800 16650 11810 16670
rect 11830 16650 11840 16670
rect 11800 16510 11840 16650
rect 11800 16490 11810 16510
rect 11830 16490 11840 16510
rect 11800 16480 11840 16490
rect 11880 16670 11920 16680
rect 11880 16650 11890 16670
rect 11910 16650 11920 16670
rect 11880 16510 11920 16650
rect 11880 16490 11890 16510
rect 11910 16490 11920 16510
rect 11880 16480 11920 16490
rect 11960 16670 12000 16680
rect 11960 16650 11970 16670
rect 11990 16650 12000 16670
rect 11960 16510 12000 16650
rect 11960 16490 11970 16510
rect 11990 16490 12000 16510
rect 11960 16480 12000 16490
rect 12040 16670 12080 16680
rect 12040 16650 12050 16670
rect 12070 16650 12080 16670
rect 12040 16510 12080 16650
rect 12040 16490 12050 16510
rect 12070 16490 12080 16510
rect 12040 16480 12080 16490
rect 12120 16670 12160 16680
rect 12120 16650 12130 16670
rect 12150 16650 12160 16670
rect 12120 16510 12160 16650
rect 12120 16490 12130 16510
rect 12150 16490 12160 16510
rect 12120 16480 12160 16490
rect 12200 16670 12240 16680
rect 12200 16650 12210 16670
rect 12230 16650 12240 16670
rect 12200 16510 12240 16650
rect 12200 16490 12210 16510
rect 12230 16490 12240 16510
rect 12200 16480 12240 16490
rect 12280 16670 12320 16680
rect 12280 16650 12290 16670
rect 12310 16650 12320 16670
rect 12280 16510 12320 16650
rect 12280 16490 12290 16510
rect 12310 16490 12320 16510
rect 12280 16480 12320 16490
rect 12360 16670 12400 16680
rect 12360 16650 12370 16670
rect 12390 16650 12400 16670
rect 12360 16510 12400 16650
rect 12360 16490 12370 16510
rect 12390 16490 12400 16510
rect 12360 16480 12400 16490
rect 12440 16670 12480 16680
rect 12440 16650 12450 16670
rect 12470 16650 12480 16670
rect 12440 16510 12480 16650
rect 12440 16490 12450 16510
rect 12470 16490 12480 16510
rect 12440 16480 12480 16490
rect 12520 16670 12560 16680
rect 12520 16650 12530 16670
rect 12550 16650 12560 16670
rect 12520 16510 12560 16650
rect 12520 16490 12530 16510
rect 12550 16490 12560 16510
rect 12520 16480 12560 16490
rect 12600 16670 12640 16680
rect 12600 16650 12610 16670
rect 12630 16650 12640 16670
rect 12600 16510 12640 16650
rect 12600 16490 12610 16510
rect 12630 16490 12640 16510
rect 12600 16480 12640 16490
rect 12680 16670 12720 16680
rect 12680 16650 12690 16670
rect 12710 16650 12720 16670
rect 12680 16510 12720 16650
rect 12680 16490 12690 16510
rect 12710 16490 12720 16510
rect 12680 16480 12720 16490
rect 12760 16670 12800 16680
rect 12760 16650 12770 16670
rect 12790 16650 12800 16670
rect 12760 16510 12800 16650
rect 12760 16490 12770 16510
rect 12790 16490 12800 16510
rect 12760 16480 12800 16490
rect 12840 16670 12880 16680
rect 12840 16650 12850 16670
rect 12870 16650 12880 16670
rect 12840 16510 12880 16650
rect 12840 16490 12850 16510
rect 12870 16490 12880 16510
rect 12840 16480 12880 16490
rect 12920 16670 12960 16680
rect 12920 16650 12930 16670
rect 12950 16650 12960 16670
rect 12920 16510 12960 16650
rect 12920 16490 12930 16510
rect 12950 16490 12960 16510
rect 12920 16480 12960 16490
rect 13000 16670 13040 16680
rect 13000 16650 13010 16670
rect 13030 16650 13040 16670
rect 13000 16510 13040 16650
rect 13000 16490 13010 16510
rect 13030 16490 13040 16510
rect 13000 16480 13040 16490
rect 13080 16670 13120 16680
rect 13080 16650 13090 16670
rect 13110 16650 13120 16670
rect 13080 16510 13120 16650
rect 13080 16490 13090 16510
rect 13110 16490 13120 16510
rect 13080 16480 13120 16490
rect 13160 16670 13200 16680
rect 13160 16650 13170 16670
rect 13190 16650 13200 16670
rect 13160 16510 13200 16650
rect 13160 16490 13170 16510
rect 13190 16490 13200 16510
rect 13160 16480 13200 16490
rect 13240 16670 13280 16680
rect 13240 16650 13250 16670
rect 13270 16650 13280 16670
rect 13240 16510 13280 16650
rect 13240 16490 13250 16510
rect 13270 16490 13280 16510
rect 13240 16480 13280 16490
rect 13320 16670 13360 16680
rect 13320 16650 13330 16670
rect 13350 16650 13360 16670
rect 13320 16510 13360 16650
rect 13320 16490 13330 16510
rect 13350 16490 13360 16510
rect 13320 16480 13360 16490
rect 13400 16670 13440 16680
rect 13400 16650 13410 16670
rect 13430 16650 13440 16670
rect 13400 16510 13440 16650
rect 13400 16490 13410 16510
rect 13430 16490 13440 16510
rect 13400 16480 13440 16490
rect 13480 16670 13520 16680
rect 13480 16650 13490 16670
rect 13510 16650 13520 16670
rect 13480 16510 13520 16650
rect 13480 16490 13490 16510
rect 13510 16490 13520 16510
rect 13480 16480 13520 16490
rect 13560 16670 13600 16680
rect 13560 16650 13570 16670
rect 13590 16650 13600 16670
rect 13560 16510 13600 16650
rect 13560 16490 13570 16510
rect 13590 16490 13600 16510
rect 13560 16480 13600 16490
rect 13640 16670 13680 16680
rect 13640 16650 13650 16670
rect 13670 16650 13680 16670
rect 13640 16510 13680 16650
rect 13640 16490 13650 16510
rect 13670 16490 13680 16510
rect 13640 16480 13680 16490
rect 13720 16670 13760 16680
rect 13720 16650 13730 16670
rect 13750 16650 13760 16670
rect 13720 16510 13760 16650
rect 13720 16490 13730 16510
rect 13750 16490 13760 16510
rect 13720 16480 13760 16490
rect 13800 16670 13840 16680
rect 13800 16650 13810 16670
rect 13830 16650 13840 16670
rect 13800 16510 13840 16650
rect 13800 16490 13810 16510
rect 13830 16490 13840 16510
rect 13800 16480 13840 16490
rect 13880 16670 13920 16680
rect 13880 16650 13890 16670
rect 13910 16650 13920 16670
rect 13880 16510 13920 16650
rect 13880 16490 13890 16510
rect 13910 16490 13920 16510
rect 13880 16480 13920 16490
rect 13960 16670 14000 16680
rect 13960 16650 13970 16670
rect 13990 16650 14000 16670
rect 13960 16510 14000 16650
rect 13960 16490 13970 16510
rect 13990 16490 14000 16510
rect 13960 16480 14000 16490
rect 14040 16670 14080 16680
rect 14040 16650 14050 16670
rect 14070 16650 14080 16670
rect 14040 16510 14080 16650
rect 14040 16490 14050 16510
rect 14070 16490 14080 16510
rect 14040 16480 14080 16490
rect 14120 16670 14160 16680
rect 14120 16650 14130 16670
rect 14150 16650 14160 16670
rect 14120 16510 14160 16650
rect 14120 16490 14130 16510
rect 14150 16490 14160 16510
rect 14120 16480 14160 16490
rect 14200 16670 14240 16680
rect 14200 16650 14210 16670
rect 14230 16650 14240 16670
rect 14200 16510 14240 16650
rect 14200 16490 14210 16510
rect 14230 16490 14240 16510
rect 14200 16480 14240 16490
rect 14280 16670 14320 16680
rect 14280 16650 14290 16670
rect 14310 16650 14320 16670
rect 14280 16510 14320 16650
rect 14280 16490 14290 16510
rect 14310 16490 14320 16510
rect 14280 16480 14320 16490
rect 14360 16670 14400 16680
rect 14360 16650 14370 16670
rect 14390 16650 14400 16670
rect 14360 16510 14400 16650
rect 14360 16490 14370 16510
rect 14390 16490 14400 16510
rect 14360 16480 14400 16490
rect 14440 16670 14480 16680
rect 14440 16650 14450 16670
rect 14470 16650 14480 16670
rect 14440 16510 14480 16650
rect 14440 16490 14450 16510
rect 14470 16490 14480 16510
rect 14440 16480 14480 16490
rect 14520 16670 14560 16680
rect 14520 16650 14530 16670
rect 14550 16650 14560 16670
rect 14520 16510 14560 16650
rect 14520 16490 14530 16510
rect 14550 16490 14560 16510
rect 14520 16480 14560 16490
rect 14600 16670 14640 16680
rect 14600 16650 14610 16670
rect 14630 16650 14640 16670
rect 14600 16510 14640 16650
rect 14600 16490 14610 16510
rect 14630 16490 14640 16510
rect 14600 16480 14640 16490
rect 14680 16670 14720 16680
rect 14680 16650 14690 16670
rect 14710 16650 14720 16670
rect 14680 16510 14720 16650
rect 14680 16490 14690 16510
rect 14710 16490 14720 16510
rect 14680 16480 14720 16490
rect 14760 16480 14800 16680
rect 14840 16480 14880 16680
rect 14920 16480 14960 16680
rect 15000 16480 15040 16680
rect 15080 16480 15120 16680
rect 15160 16480 15200 16680
rect 15240 16480 15280 16680
rect 15320 16480 15360 16680
rect 15400 16480 15440 16680
rect 15480 16480 15520 16680
rect 15560 16480 15600 16680
rect 15640 16480 15680 16680
rect 15720 16480 15760 16680
rect 15800 16480 15840 16680
rect 15880 16480 15920 16680
rect 15960 16480 16000 16680
rect 16040 16480 16080 16680
rect 16120 16480 16160 16680
rect 16200 16480 16240 16680
rect 16280 16480 16320 16680
rect 16360 16480 16400 16680
rect 16440 16480 16480 16680
rect 16520 16480 16560 16680
rect 16600 16480 16640 16680
rect 16680 16480 16720 16680
rect 16760 16670 16800 16680
rect 16760 16650 16770 16670
rect 16790 16650 16800 16670
rect 16760 16510 16800 16650
rect 16760 16490 16770 16510
rect 16790 16490 16800 16510
rect 16760 16480 16800 16490
rect 16840 16670 16880 16680
rect 16840 16650 16850 16670
rect 16870 16650 16880 16670
rect 16840 16510 16880 16650
rect 16840 16490 16850 16510
rect 16870 16490 16880 16510
rect 16840 16480 16880 16490
rect 16920 16670 16960 16680
rect 16920 16650 16930 16670
rect 16950 16650 16960 16670
rect 16920 16510 16960 16650
rect 16920 16490 16930 16510
rect 16950 16490 16960 16510
rect 16920 16480 16960 16490
rect 17000 16670 17040 16680
rect 17000 16650 17010 16670
rect 17030 16650 17040 16670
rect 17000 16510 17040 16650
rect 17000 16490 17010 16510
rect 17030 16490 17040 16510
rect 17000 16480 17040 16490
rect 17080 16670 17120 16680
rect 17080 16650 17090 16670
rect 17110 16650 17120 16670
rect 17080 16510 17120 16650
rect 17080 16490 17090 16510
rect 17110 16490 17120 16510
rect 17080 16480 17120 16490
rect 17160 16670 17200 16680
rect 17160 16650 17170 16670
rect 17190 16650 17200 16670
rect 17160 16510 17200 16650
rect 17160 16490 17170 16510
rect 17190 16490 17200 16510
rect 17160 16480 17200 16490
rect 17240 16670 17280 16680
rect 17240 16650 17250 16670
rect 17270 16650 17280 16670
rect 17240 16510 17280 16650
rect 17240 16490 17250 16510
rect 17270 16490 17280 16510
rect 17240 16480 17280 16490
rect 17320 16670 17360 16680
rect 17320 16650 17330 16670
rect 17350 16650 17360 16670
rect 17320 16510 17360 16650
rect 17320 16490 17330 16510
rect 17350 16490 17360 16510
rect 17320 16480 17360 16490
rect 17400 16670 17440 16680
rect 17400 16650 17410 16670
rect 17430 16650 17440 16670
rect 17400 16510 17440 16650
rect 17400 16490 17410 16510
rect 17430 16490 17440 16510
rect 17400 16480 17440 16490
rect 17480 16670 17520 16680
rect 17480 16650 17490 16670
rect 17510 16650 17520 16670
rect 17480 16510 17520 16650
rect 17480 16490 17490 16510
rect 17510 16490 17520 16510
rect 17480 16480 17520 16490
rect 17560 16670 17600 16680
rect 17560 16650 17570 16670
rect 17590 16650 17600 16670
rect 17560 16510 17600 16650
rect 17560 16490 17570 16510
rect 17590 16490 17600 16510
rect 17560 16480 17600 16490
rect 17640 16670 17680 16680
rect 17640 16650 17650 16670
rect 17670 16650 17680 16670
rect 17640 16510 17680 16650
rect 17640 16490 17650 16510
rect 17670 16490 17680 16510
rect 17640 16480 17680 16490
rect 17720 16670 17760 16680
rect 17720 16650 17730 16670
rect 17750 16650 17760 16670
rect 17720 16510 17760 16650
rect 17720 16490 17730 16510
rect 17750 16490 17760 16510
rect 17720 16480 17760 16490
rect 17800 16670 17840 16680
rect 17800 16650 17810 16670
rect 17830 16650 17840 16670
rect 17800 16510 17840 16650
rect 17800 16490 17810 16510
rect 17830 16490 17840 16510
rect 17800 16480 17840 16490
rect 17880 16670 17920 16680
rect 17880 16650 17890 16670
rect 17910 16650 17920 16670
rect 17880 16510 17920 16650
rect 17880 16490 17890 16510
rect 17910 16490 17920 16510
rect 17880 16480 17920 16490
rect 17960 16670 18000 16680
rect 17960 16650 17970 16670
rect 17990 16650 18000 16670
rect 17960 16510 18000 16650
rect 17960 16490 17970 16510
rect 17990 16490 18000 16510
rect 17960 16480 18000 16490
rect 18040 16670 18080 16680
rect 18040 16650 18050 16670
rect 18070 16650 18080 16670
rect 18040 16510 18080 16650
rect 18040 16490 18050 16510
rect 18070 16490 18080 16510
rect 18040 16480 18080 16490
rect 18120 16670 18160 16680
rect 18120 16650 18130 16670
rect 18150 16650 18160 16670
rect 18120 16510 18160 16650
rect 18120 16490 18130 16510
rect 18150 16490 18160 16510
rect 18120 16480 18160 16490
rect 18200 16670 18240 16680
rect 18200 16650 18210 16670
rect 18230 16650 18240 16670
rect 18200 16510 18240 16650
rect 18200 16490 18210 16510
rect 18230 16490 18240 16510
rect 18200 16480 18240 16490
rect 18280 16670 18320 16680
rect 18280 16650 18290 16670
rect 18310 16650 18320 16670
rect 18280 16510 18320 16650
rect 18280 16490 18290 16510
rect 18310 16490 18320 16510
rect 18280 16480 18320 16490
rect 18360 16670 18400 16680
rect 18360 16650 18370 16670
rect 18390 16650 18400 16670
rect 18360 16510 18400 16650
rect 18360 16490 18370 16510
rect 18390 16490 18400 16510
rect 18360 16480 18400 16490
rect 18440 16670 18480 16680
rect 18440 16650 18450 16670
rect 18470 16650 18480 16670
rect 18440 16510 18480 16650
rect 18440 16490 18450 16510
rect 18470 16490 18480 16510
rect 18440 16480 18480 16490
rect 18520 16670 18560 16680
rect 18520 16650 18530 16670
rect 18550 16650 18560 16670
rect 18520 16510 18560 16650
rect 18520 16490 18530 16510
rect 18550 16490 18560 16510
rect 18520 16480 18560 16490
rect 18600 16670 18640 16680
rect 18600 16650 18610 16670
rect 18630 16650 18640 16670
rect 18600 16510 18640 16650
rect 18600 16490 18610 16510
rect 18630 16490 18640 16510
rect 18600 16480 18640 16490
rect 18680 16670 18720 16680
rect 18680 16650 18690 16670
rect 18710 16650 18720 16670
rect 18680 16510 18720 16650
rect 18680 16490 18690 16510
rect 18710 16490 18720 16510
rect 18680 16480 18720 16490
rect 18760 16670 18800 16680
rect 18760 16650 18770 16670
rect 18790 16650 18800 16670
rect 18760 16510 18800 16650
rect 18760 16490 18770 16510
rect 18790 16490 18800 16510
rect 18760 16480 18800 16490
rect 18840 16670 18880 16680
rect 18840 16650 18850 16670
rect 18870 16650 18880 16670
rect 18840 16510 18880 16650
rect 18840 16490 18850 16510
rect 18870 16490 18880 16510
rect 18840 16480 18880 16490
rect 18920 16670 18960 16680
rect 18920 16650 18930 16670
rect 18950 16650 18960 16670
rect 18920 16510 18960 16650
rect 18920 16490 18930 16510
rect 18950 16490 18960 16510
rect 18920 16480 18960 16490
rect 19000 16670 19040 16680
rect 19000 16650 19010 16670
rect 19030 16650 19040 16670
rect 19000 16510 19040 16650
rect 19000 16490 19010 16510
rect 19030 16490 19040 16510
rect 19000 16480 19040 16490
rect 19080 16670 19120 16680
rect 19080 16650 19090 16670
rect 19110 16650 19120 16670
rect 19080 16510 19120 16650
rect 19080 16490 19090 16510
rect 19110 16490 19120 16510
rect 19080 16480 19120 16490
rect 19160 16670 19200 16680
rect 19160 16650 19170 16670
rect 19190 16650 19200 16670
rect 19160 16510 19200 16650
rect 19160 16490 19170 16510
rect 19190 16490 19200 16510
rect 19160 16480 19200 16490
rect 19240 16670 19280 16680
rect 19240 16650 19250 16670
rect 19270 16650 19280 16670
rect 19240 16510 19280 16650
rect 19240 16490 19250 16510
rect 19270 16490 19280 16510
rect 19240 16480 19280 16490
rect 19320 16670 19360 16680
rect 19320 16650 19330 16670
rect 19350 16650 19360 16670
rect 19320 16510 19360 16650
rect 19320 16490 19330 16510
rect 19350 16490 19360 16510
rect 19320 16480 19360 16490
rect 19400 16670 19440 16680
rect 19400 16650 19410 16670
rect 19430 16650 19440 16670
rect 19400 16510 19440 16650
rect 19400 16490 19410 16510
rect 19430 16490 19440 16510
rect 19400 16480 19440 16490
rect 19480 16670 19520 16680
rect 19480 16650 19490 16670
rect 19510 16650 19520 16670
rect 19480 16510 19520 16650
rect 19480 16490 19490 16510
rect 19510 16490 19520 16510
rect 19480 16480 19520 16490
rect 19560 16670 19600 16680
rect 19560 16650 19570 16670
rect 19590 16650 19600 16670
rect 19560 16510 19600 16650
rect 19560 16490 19570 16510
rect 19590 16490 19600 16510
rect 19560 16480 19600 16490
rect 19640 16670 19680 16680
rect 19640 16650 19650 16670
rect 19670 16650 19680 16670
rect 19640 16510 19680 16650
rect 19640 16490 19650 16510
rect 19670 16490 19680 16510
rect 19640 16480 19680 16490
rect 19720 16670 19760 16680
rect 19720 16650 19730 16670
rect 19750 16650 19760 16670
rect 19720 16510 19760 16650
rect 19720 16490 19730 16510
rect 19750 16490 19760 16510
rect 19720 16480 19760 16490
rect 19800 16670 19840 16680
rect 19800 16650 19810 16670
rect 19830 16650 19840 16670
rect 19800 16510 19840 16650
rect 19800 16490 19810 16510
rect 19830 16490 19840 16510
rect 19800 16480 19840 16490
rect 19880 16670 19920 16680
rect 19880 16650 19890 16670
rect 19910 16650 19920 16670
rect 19880 16510 19920 16650
rect 19880 16490 19890 16510
rect 19910 16490 19920 16510
rect 19880 16480 19920 16490
rect 19960 16670 20000 16680
rect 19960 16650 19970 16670
rect 19990 16650 20000 16670
rect 19960 16510 20000 16650
rect 19960 16490 19970 16510
rect 19990 16490 20000 16510
rect 19960 16480 20000 16490
rect 20040 16670 20080 16680
rect 20040 16650 20050 16670
rect 20070 16650 20080 16670
rect 20040 16510 20080 16650
rect 20040 16490 20050 16510
rect 20070 16490 20080 16510
rect 20040 16480 20080 16490
rect 20120 16670 20160 16680
rect 20120 16650 20130 16670
rect 20150 16650 20160 16670
rect 20120 16510 20160 16650
rect 20120 16490 20130 16510
rect 20150 16490 20160 16510
rect 20120 16480 20160 16490
rect 20200 16670 20240 16680
rect 20200 16650 20210 16670
rect 20230 16650 20240 16670
rect 20200 16510 20240 16650
rect 20200 16490 20210 16510
rect 20230 16490 20240 16510
rect 20200 16480 20240 16490
rect 20280 16670 20320 16680
rect 20280 16650 20290 16670
rect 20310 16650 20320 16670
rect 20280 16510 20320 16650
rect 20280 16490 20290 16510
rect 20310 16490 20320 16510
rect 20280 16480 20320 16490
rect 20360 16670 20400 16680
rect 20360 16650 20370 16670
rect 20390 16650 20400 16670
rect 20360 16510 20400 16650
rect 20360 16490 20370 16510
rect 20390 16490 20400 16510
rect 20360 16480 20400 16490
rect 20440 16670 20480 16680
rect 20440 16650 20450 16670
rect 20470 16650 20480 16670
rect 20440 16510 20480 16650
rect 20440 16490 20450 16510
rect 20470 16490 20480 16510
rect 20440 16480 20480 16490
rect 20520 16670 20560 16680
rect 20520 16650 20530 16670
rect 20550 16650 20560 16670
rect 20520 16510 20560 16650
rect 20520 16490 20530 16510
rect 20550 16490 20560 16510
rect 20520 16480 20560 16490
rect 20600 16670 20640 16680
rect 20600 16650 20610 16670
rect 20630 16650 20640 16670
rect 20600 16510 20640 16650
rect 20600 16490 20610 16510
rect 20630 16490 20640 16510
rect 20600 16480 20640 16490
rect 20680 16670 20720 16680
rect 20680 16650 20690 16670
rect 20710 16650 20720 16670
rect 20680 16510 20720 16650
rect 20680 16490 20690 16510
rect 20710 16490 20720 16510
rect 20680 16480 20720 16490
rect 20760 16670 20800 16680
rect 20760 16650 20770 16670
rect 20790 16650 20800 16670
rect 20760 16510 20800 16650
rect 20760 16490 20770 16510
rect 20790 16490 20800 16510
rect 20760 16480 20800 16490
rect 20840 16670 20880 16680
rect 20840 16650 20850 16670
rect 20870 16650 20880 16670
rect 20840 16510 20880 16650
rect 20840 16490 20850 16510
rect 20870 16490 20880 16510
rect 20840 16480 20880 16490
rect 20920 16670 20960 16680
rect 20920 16650 20930 16670
rect 20950 16650 20960 16670
rect 20920 16510 20960 16650
rect 20920 16490 20930 16510
rect 20950 16490 20960 16510
rect 20920 16480 20960 16490
rect 0 16430 40 16440
rect 0 16410 10 16430
rect 30 16410 40 16430
rect 0 16270 40 16410
rect 0 16250 10 16270
rect 30 16250 40 16270
rect 0 16240 40 16250
rect 80 16430 120 16440
rect 80 16410 90 16430
rect 110 16410 120 16430
rect 80 16270 120 16410
rect 80 16250 90 16270
rect 110 16250 120 16270
rect 80 16240 120 16250
rect 160 16430 200 16440
rect 160 16410 170 16430
rect 190 16410 200 16430
rect 160 16270 200 16410
rect 160 16250 170 16270
rect 190 16250 200 16270
rect 160 16240 200 16250
rect 240 16430 280 16440
rect 240 16410 250 16430
rect 270 16410 280 16430
rect 240 16270 280 16410
rect 240 16250 250 16270
rect 270 16250 280 16270
rect 240 16240 280 16250
rect 320 16430 360 16440
rect 320 16410 330 16430
rect 350 16410 360 16430
rect 320 16270 360 16410
rect 320 16250 330 16270
rect 350 16250 360 16270
rect 320 16240 360 16250
rect 400 16430 440 16440
rect 400 16410 410 16430
rect 430 16410 440 16430
rect 400 16270 440 16410
rect 400 16250 410 16270
rect 430 16250 440 16270
rect 400 16240 440 16250
rect 480 16430 520 16440
rect 480 16410 490 16430
rect 510 16410 520 16430
rect 480 16270 520 16410
rect 480 16250 490 16270
rect 510 16250 520 16270
rect 480 16240 520 16250
rect 560 16430 600 16440
rect 560 16410 570 16430
rect 590 16410 600 16430
rect 560 16270 600 16410
rect 560 16250 570 16270
rect 590 16250 600 16270
rect 560 16240 600 16250
rect 640 16430 680 16440
rect 640 16410 650 16430
rect 670 16410 680 16430
rect 640 16270 680 16410
rect 640 16250 650 16270
rect 670 16250 680 16270
rect 640 16240 680 16250
rect 720 16430 760 16440
rect 720 16410 730 16430
rect 750 16410 760 16430
rect 720 16270 760 16410
rect 720 16250 730 16270
rect 750 16250 760 16270
rect 720 16240 760 16250
rect 800 16430 840 16440
rect 800 16410 810 16430
rect 830 16410 840 16430
rect 800 16270 840 16410
rect 800 16250 810 16270
rect 830 16250 840 16270
rect 800 16240 840 16250
rect 880 16430 920 16440
rect 880 16410 890 16430
rect 910 16410 920 16430
rect 880 16270 920 16410
rect 880 16250 890 16270
rect 910 16250 920 16270
rect 880 16240 920 16250
rect 960 16430 1000 16440
rect 960 16410 970 16430
rect 990 16410 1000 16430
rect 960 16270 1000 16410
rect 960 16250 970 16270
rect 990 16250 1000 16270
rect 960 16240 1000 16250
rect 1040 16430 1080 16440
rect 1040 16410 1050 16430
rect 1070 16410 1080 16430
rect 1040 16270 1080 16410
rect 1040 16250 1050 16270
rect 1070 16250 1080 16270
rect 1040 16240 1080 16250
rect 1120 16430 1160 16440
rect 1120 16410 1130 16430
rect 1150 16410 1160 16430
rect 1120 16270 1160 16410
rect 1120 16250 1130 16270
rect 1150 16250 1160 16270
rect 1120 16240 1160 16250
rect 1200 16430 1240 16440
rect 1200 16410 1210 16430
rect 1230 16410 1240 16430
rect 1200 16270 1240 16410
rect 1200 16250 1210 16270
rect 1230 16250 1240 16270
rect 1200 16240 1240 16250
rect 1280 16430 1320 16440
rect 1280 16410 1290 16430
rect 1310 16410 1320 16430
rect 1280 16270 1320 16410
rect 1280 16250 1290 16270
rect 1310 16250 1320 16270
rect 1280 16240 1320 16250
rect 1360 16430 1400 16440
rect 1360 16410 1370 16430
rect 1390 16410 1400 16430
rect 1360 16270 1400 16410
rect 1360 16250 1370 16270
rect 1390 16250 1400 16270
rect 1360 16240 1400 16250
rect 1440 16430 1480 16440
rect 1440 16410 1450 16430
rect 1470 16410 1480 16430
rect 1440 16270 1480 16410
rect 1440 16250 1450 16270
rect 1470 16250 1480 16270
rect 1440 16240 1480 16250
rect 1520 16430 1560 16440
rect 1520 16410 1530 16430
rect 1550 16410 1560 16430
rect 1520 16270 1560 16410
rect 1520 16250 1530 16270
rect 1550 16250 1560 16270
rect 1520 16240 1560 16250
rect 1600 16430 1640 16440
rect 1600 16410 1610 16430
rect 1630 16410 1640 16430
rect 1600 16270 1640 16410
rect 1600 16250 1610 16270
rect 1630 16250 1640 16270
rect 1600 16240 1640 16250
rect 1680 16430 1720 16440
rect 1680 16410 1690 16430
rect 1710 16410 1720 16430
rect 1680 16270 1720 16410
rect 1680 16250 1690 16270
rect 1710 16250 1720 16270
rect 1680 16240 1720 16250
rect 1760 16430 1800 16440
rect 1760 16410 1770 16430
rect 1790 16410 1800 16430
rect 1760 16270 1800 16410
rect 1760 16250 1770 16270
rect 1790 16250 1800 16270
rect 1760 16240 1800 16250
rect 1840 16430 1880 16440
rect 1840 16410 1850 16430
rect 1870 16410 1880 16430
rect 1840 16270 1880 16410
rect 1840 16250 1850 16270
rect 1870 16250 1880 16270
rect 1840 16240 1880 16250
rect 1920 16430 1960 16440
rect 1920 16410 1930 16430
rect 1950 16410 1960 16430
rect 1920 16270 1960 16410
rect 1920 16250 1930 16270
rect 1950 16250 1960 16270
rect 1920 16240 1960 16250
rect 2000 16430 2040 16440
rect 2000 16410 2010 16430
rect 2030 16410 2040 16430
rect 2000 16270 2040 16410
rect 2000 16250 2010 16270
rect 2030 16250 2040 16270
rect 2000 16240 2040 16250
rect 2080 16430 2120 16440
rect 2080 16410 2090 16430
rect 2110 16410 2120 16430
rect 2080 16270 2120 16410
rect 2080 16250 2090 16270
rect 2110 16250 2120 16270
rect 2080 16240 2120 16250
rect 2160 16430 2200 16440
rect 2160 16410 2170 16430
rect 2190 16410 2200 16430
rect 2160 16270 2200 16410
rect 2160 16250 2170 16270
rect 2190 16250 2200 16270
rect 2160 16240 2200 16250
rect 2240 16430 2280 16440
rect 2240 16410 2250 16430
rect 2270 16410 2280 16430
rect 2240 16270 2280 16410
rect 2240 16250 2250 16270
rect 2270 16250 2280 16270
rect 2240 16240 2280 16250
rect 2320 16430 2360 16440
rect 2320 16410 2330 16430
rect 2350 16410 2360 16430
rect 2320 16270 2360 16410
rect 2320 16250 2330 16270
rect 2350 16250 2360 16270
rect 2320 16240 2360 16250
rect 2400 16430 2440 16440
rect 2400 16410 2410 16430
rect 2430 16410 2440 16430
rect 2400 16270 2440 16410
rect 2400 16250 2410 16270
rect 2430 16250 2440 16270
rect 2400 16240 2440 16250
rect 2480 16430 2520 16440
rect 2480 16410 2490 16430
rect 2510 16410 2520 16430
rect 2480 16270 2520 16410
rect 2480 16250 2490 16270
rect 2510 16250 2520 16270
rect 2480 16240 2520 16250
rect 2560 16430 2600 16440
rect 2560 16410 2570 16430
rect 2590 16410 2600 16430
rect 2560 16270 2600 16410
rect 2560 16250 2570 16270
rect 2590 16250 2600 16270
rect 2560 16240 2600 16250
rect 2640 16430 2680 16440
rect 2640 16410 2650 16430
rect 2670 16410 2680 16430
rect 2640 16270 2680 16410
rect 2640 16250 2650 16270
rect 2670 16250 2680 16270
rect 2640 16240 2680 16250
rect 2720 16430 2760 16440
rect 2720 16410 2730 16430
rect 2750 16410 2760 16430
rect 2720 16270 2760 16410
rect 2720 16250 2730 16270
rect 2750 16250 2760 16270
rect 2720 16240 2760 16250
rect 2800 16430 2840 16440
rect 2800 16410 2810 16430
rect 2830 16410 2840 16430
rect 2800 16270 2840 16410
rect 2800 16250 2810 16270
rect 2830 16250 2840 16270
rect 2800 16240 2840 16250
rect 2880 16430 2920 16440
rect 2880 16410 2890 16430
rect 2910 16410 2920 16430
rect 2880 16270 2920 16410
rect 2880 16250 2890 16270
rect 2910 16250 2920 16270
rect 2880 16240 2920 16250
rect 2960 16430 3000 16440
rect 2960 16410 2970 16430
rect 2990 16410 3000 16430
rect 2960 16270 3000 16410
rect 2960 16250 2970 16270
rect 2990 16250 3000 16270
rect 2960 16240 3000 16250
rect 3040 16430 3080 16440
rect 3040 16410 3050 16430
rect 3070 16410 3080 16430
rect 3040 16270 3080 16410
rect 3040 16250 3050 16270
rect 3070 16250 3080 16270
rect 3040 16240 3080 16250
rect 3120 16430 3160 16440
rect 3120 16410 3130 16430
rect 3150 16410 3160 16430
rect 3120 16270 3160 16410
rect 3120 16250 3130 16270
rect 3150 16250 3160 16270
rect 3120 16240 3160 16250
rect 3200 16430 3240 16440
rect 3200 16410 3210 16430
rect 3230 16410 3240 16430
rect 3200 16270 3240 16410
rect 3200 16250 3210 16270
rect 3230 16250 3240 16270
rect 3200 16240 3240 16250
rect 3280 16430 3320 16440
rect 3280 16410 3290 16430
rect 3310 16410 3320 16430
rect 3280 16270 3320 16410
rect 3280 16250 3290 16270
rect 3310 16250 3320 16270
rect 3280 16240 3320 16250
rect 3360 16430 3400 16440
rect 3360 16410 3370 16430
rect 3390 16410 3400 16430
rect 3360 16270 3400 16410
rect 3360 16250 3370 16270
rect 3390 16250 3400 16270
rect 3360 16240 3400 16250
rect 3440 16430 3480 16440
rect 3440 16410 3450 16430
rect 3470 16410 3480 16430
rect 3440 16270 3480 16410
rect 3440 16250 3450 16270
rect 3470 16250 3480 16270
rect 3440 16240 3480 16250
rect 3520 16430 3560 16440
rect 3520 16410 3530 16430
rect 3550 16410 3560 16430
rect 3520 16270 3560 16410
rect 3520 16250 3530 16270
rect 3550 16250 3560 16270
rect 3520 16240 3560 16250
rect 3600 16430 3640 16440
rect 3600 16410 3610 16430
rect 3630 16410 3640 16430
rect 3600 16270 3640 16410
rect 3600 16250 3610 16270
rect 3630 16250 3640 16270
rect 3600 16240 3640 16250
rect 3680 16430 3720 16440
rect 3680 16410 3690 16430
rect 3710 16410 3720 16430
rect 3680 16270 3720 16410
rect 3680 16250 3690 16270
rect 3710 16250 3720 16270
rect 3680 16240 3720 16250
rect 3760 16430 3800 16440
rect 3760 16410 3770 16430
rect 3790 16410 3800 16430
rect 3760 16270 3800 16410
rect 3760 16250 3770 16270
rect 3790 16250 3800 16270
rect 3760 16240 3800 16250
rect 3840 16430 3880 16440
rect 3840 16410 3850 16430
rect 3870 16410 3880 16430
rect 3840 16270 3880 16410
rect 3840 16250 3850 16270
rect 3870 16250 3880 16270
rect 3840 16240 3880 16250
rect 3920 16430 3960 16440
rect 3920 16410 3930 16430
rect 3950 16410 3960 16430
rect 3920 16270 3960 16410
rect 3920 16250 3930 16270
rect 3950 16250 3960 16270
rect 3920 16240 3960 16250
rect 4000 16430 4040 16440
rect 4000 16410 4010 16430
rect 4030 16410 4040 16430
rect 4000 16270 4040 16410
rect 4000 16250 4010 16270
rect 4030 16250 4040 16270
rect 4000 16240 4040 16250
rect 4080 16430 4120 16440
rect 4080 16410 4090 16430
rect 4110 16410 4120 16430
rect 4080 16270 4120 16410
rect 4080 16250 4090 16270
rect 4110 16250 4120 16270
rect 4080 16240 4120 16250
rect 4160 16430 4200 16440
rect 4160 16410 4170 16430
rect 4190 16410 4200 16430
rect 4160 16270 4200 16410
rect 4160 16250 4170 16270
rect 4190 16250 4200 16270
rect 4160 16240 4200 16250
rect 4240 16240 4280 16440
rect 4320 16240 4360 16440
rect 4400 16240 4440 16440
rect 4480 16240 4520 16440
rect 4560 16240 4600 16440
rect 4640 16240 4680 16440
rect 4720 16240 4760 16440
rect 4800 16240 4840 16440
rect 4880 16240 4920 16440
rect 4960 16240 5000 16440
rect 5040 16240 5080 16440
rect 5120 16240 5160 16440
rect 5200 16240 5240 16440
rect 5280 16240 5320 16440
rect 5360 16240 5400 16440
rect 5440 16240 5480 16440
rect 5520 16240 5560 16440
rect 5600 16240 5640 16440
rect 5680 16240 5720 16440
rect 5760 16240 5800 16440
rect 5840 16240 5880 16440
rect 5920 16240 5960 16440
rect 6000 16240 6040 16440
rect 6080 16240 6120 16440
rect 6160 16240 6200 16440
rect 6240 16430 6280 16440
rect 6240 16410 6250 16430
rect 6270 16410 6280 16430
rect 6240 16270 6280 16410
rect 6240 16250 6250 16270
rect 6270 16250 6280 16270
rect 6240 16240 6280 16250
rect 6320 16430 6360 16440
rect 6320 16410 6330 16430
rect 6350 16410 6360 16430
rect 6320 16270 6360 16410
rect 6320 16250 6330 16270
rect 6350 16250 6360 16270
rect 6320 16240 6360 16250
rect 6400 16430 6440 16440
rect 6400 16410 6410 16430
rect 6430 16410 6440 16430
rect 6400 16270 6440 16410
rect 6400 16250 6410 16270
rect 6430 16250 6440 16270
rect 6400 16240 6440 16250
rect 6480 16430 6520 16440
rect 6480 16410 6490 16430
rect 6510 16410 6520 16430
rect 6480 16270 6520 16410
rect 6480 16250 6490 16270
rect 6510 16250 6520 16270
rect 6480 16240 6520 16250
rect 6560 16430 6600 16440
rect 6560 16410 6570 16430
rect 6590 16410 6600 16430
rect 6560 16270 6600 16410
rect 6560 16250 6570 16270
rect 6590 16250 6600 16270
rect 6560 16240 6600 16250
rect 6640 16430 6680 16440
rect 6640 16410 6650 16430
rect 6670 16410 6680 16430
rect 6640 16270 6680 16410
rect 6640 16250 6650 16270
rect 6670 16250 6680 16270
rect 6640 16240 6680 16250
rect 6720 16430 6760 16440
rect 6720 16410 6730 16430
rect 6750 16410 6760 16430
rect 6720 16270 6760 16410
rect 6720 16250 6730 16270
rect 6750 16250 6760 16270
rect 6720 16240 6760 16250
rect 6800 16430 6840 16440
rect 6800 16410 6810 16430
rect 6830 16410 6840 16430
rect 6800 16270 6840 16410
rect 6800 16250 6810 16270
rect 6830 16250 6840 16270
rect 6800 16240 6840 16250
rect 6880 16430 6920 16440
rect 6880 16410 6890 16430
rect 6910 16410 6920 16430
rect 6880 16270 6920 16410
rect 6880 16250 6890 16270
rect 6910 16250 6920 16270
rect 6880 16240 6920 16250
rect 6960 16430 7000 16440
rect 6960 16410 6970 16430
rect 6990 16410 7000 16430
rect 6960 16270 7000 16410
rect 6960 16250 6970 16270
rect 6990 16250 7000 16270
rect 6960 16240 7000 16250
rect 7040 16430 7080 16440
rect 7040 16410 7050 16430
rect 7070 16410 7080 16430
rect 7040 16270 7080 16410
rect 7040 16250 7050 16270
rect 7070 16250 7080 16270
rect 7040 16240 7080 16250
rect 7120 16430 7160 16440
rect 7120 16410 7130 16430
rect 7150 16410 7160 16430
rect 7120 16270 7160 16410
rect 7120 16250 7130 16270
rect 7150 16250 7160 16270
rect 7120 16240 7160 16250
rect 7200 16430 7240 16440
rect 7200 16410 7210 16430
rect 7230 16410 7240 16430
rect 7200 16270 7240 16410
rect 7200 16250 7210 16270
rect 7230 16250 7240 16270
rect 7200 16240 7240 16250
rect 7280 16430 7320 16440
rect 7280 16410 7290 16430
rect 7310 16410 7320 16430
rect 7280 16270 7320 16410
rect 7280 16250 7290 16270
rect 7310 16250 7320 16270
rect 7280 16240 7320 16250
rect 7360 16430 7400 16440
rect 7360 16410 7370 16430
rect 7390 16410 7400 16430
rect 7360 16270 7400 16410
rect 7360 16250 7370 16270
rect 7390 16250 7400 16270
rect 7360 16240 7400 16250
rect 7440 16430 7480 16440
rect 7440 16410 7450 16430
rect 7470 16410 7480 16430
rect 7440 16270 7480 16410
rect 7440 16250 7450 16270
rect 7470 16250 7480 16270
rect 7440 16240 7480 16250
rect 7520 16430 7560 16440
rect 7520 16410 7530 16430
rect 7550 16410 7560 16430
rect 7520 16270 7560 16410
rect 7520 16250 7530 16270
rect 7550 16250 7560 16270
rect 7520 16240 7560 16250
rect 7600 16430 7640 16440
rect 7600 16410 7610 16430
rect 7630 16410 7640 16430
rect 7600 16270 7640 16410
rect 7600 16250 7610 16270
rect 7630 16250 7640 16270
rect 7600 16240 7640 16250
rect 7680 16430 7720 16440
rect 7680 16410 7690 16430
rect 7710 16410 7720 16430
rect 7680 16270 7720 16410
rect 7680 16250 7690 16270
rect 7710 16250 7720 16270
rect 7680 16240 7720 16250
rect 7760 16430 7800 16440
rect 7760 16410 7770 16430
rect 7790 16410 7800 16430
rect 7760 16270 7800 16410
rect 7760 16250 7770 16270
rect 7790 16250 7800 16270
rect 7760 16240 7800 16250
rect 7840 16430 7880 16440
rect 7840 16410 7850 16430
rect 7870 16410 7880 16430
rect 7840 16270 7880 16410
rect 7840 16250 7850 16270
rect 7870 16250 7880 16270
rect 7840 16240 7880 16250
rect 7920 16430 7960 16440
rect 7920 16410 7930 16430
rect 7950 16410 7960 16430
rect 7920 16270 7960 16410
rect 7920 16250 7930 16270
rect 7950 16250 7960 16270
rect 7920 16240 7960 16250
rect 8000 16430 8040 16440
rect 8000 16410 8010 16430
rect 8030 16410 8040 16430
rect 8000 16270 8040 16410
rect 8000 16250 8010 16270
rect 8030 16250 8040 16270
rect 8000 16240 8040 16250
rect 8080 16430 8120 16440
rect 8080 16410 8090 16430
rect 8110 16410 8120 16430
rect 8080 16270 8120 16410
rect 8080 16250 8090 16270
rect 8110 16250 8120 16270
rect 8080 16240 8120 16250
rect 8160 16430 8200 16440
rect 8160 16410 8170 16430
rect 8190 16410 8200 16430
rect 8160 16270 8200 16410
rect 8160 16250 8170 16270
rect 8190 16250 8200 16270
rect 8160 16240 8200 16250
rect 8240 16430 8280 16440
rect 8240 16410 8250 16430
rect 8270 16410 8280 16430
rect 8240 16270 8280 16410
rect 8240 16250 8250 16270
rect 8270 16250 8280 16270
rect 8240 16240 8280 16250
rect 8320 16430 8360 16440
rect 8320 16410 8330 16430
rect 8350 16410 8360 16430
rect 8320 16270 8360 16410
rect 8320 16250 8330 16270
rect 8350 16250 8360 16270
rect 8320 16240 8360 16250
rect 8400 16430 8440 16440
rect 8400 16410 8410 16430
rect 8430 16410 8440 16430
rect 8400 16270 8440 16410
rect 8400 16250 8410 16270
rect 8430 16250 8440 16270
rect 8400 16240 8440 16250
rect 8480 16430 8520 16440
rect 8480 16410 8490 16430
rect 8510 16410 8520 16430
rect 8480 16270 8520 16410
rect 8480 16250 8490 16270
rect 8510 16250 8520 16270
rect 8480 16240 8520 16250
rect 8560 16430 8600 16440
rect 8560 16410 8570 16430
rect 8590 16410 8600 16430
rect 8560 16270 8600 16410
rect 8560 16250 8570 16270
rect 8590 16250 8600 16270
rect 8560 16240 8600 16250
rect 8640 16430 8680 16440
rect 8640 16410 8650 16430
rect 8670 16410 8680 16430
rect 8640 16270 8680 16410
rect 8640 16250 8650 16270
rect 8670 16250 8680 16270
rect 8640 16240 8680 16250
rect 8720 16430 8760 16440
rect 8720 16410 8730 16430
rect 8750 16410 8760 16430
rect 8720 16270 8760 16410
rect 8720 16250 8730 16270
rect 8750 16250 8760 16270
rect 8720 16240 8760 16250
rect 8800 16430 8840 16440
rect 8800 16410 8810 16430
rect 8830 16410 8840 16430
rect 8800 16270 8840 16410
rect 8800 16250 8810 16270
rect 8830 16250 8840 16270
rect 8800 16240 8840 16250
rect 8880 16430 8920 16440
rect 8880 16410 8890 16430
rect 8910 16410 8920 16430
rect 8880 16270 8920 16410
rect 8880 16250 8890 16270
rect 8910 16250 8920 16270
rect 8880 16240 8920 16250
rect 8960 16430 9000 16440
rect 8960 16410 8970 16430
rect 8990 16410 9000 16430
rect 8960 16270 9000 16410
rect 8960 16250 8970 16270
rect 8990 16250 9000 16270
rect 8960 16240 9000 16250
rect 9040 16430 9080 16440
rect 9040 16410 9050 16430
rect 9070 16410 9080 16430
rect 9040 16270 9080 16410
rect 9040 16250 9050 16270
rect 9070 16250 9080 16270
rect 9040 16240 9080 16250
rect 9120 16430 9160 16440
rect 9120 16410 9130 16430
rect 9150 16410 9160 16430
rect 9120 16270 9160 16410
rect 9120 16250 9130 16270
rect 9150 16250 9160 16270
rect 9120 16240 9160 16250
rect 9200 16430 9240 16440
rect 9200 16410 9210 16430
rect 9230 16410 9240 16430
rect 9200 16270 9240 16410
rect 9200 16250 9210 16270
rect 9230 16250 9240 16270
rect 9200 16240 9240 16250
rect 9280 16430 9320 16440
rect 9280 16410 9290 16430
rect 9310 16410 9320 16430
rect 9280 16270 9320 16410
rect 9280 16250 9290 16270
rect 9310 16250 9320 16270
rect 9280 16240 9320 16250
rect 9360 16430 9400 16440
rect 9360 16410 9370 16430
rect 9390 16410 9400 16430
rect 9360 16270 9400 16410
rect 9360 16250 9370 16270
rect 9390 16250 9400 16270
rect 9360 16240 9400 16250
rect 9440 16430 9480 16440
rect 9440 16410 9450 16430
rect 9470 16410 9480 16430
rect 9440 16270 9480 16410
rect 9440 16250 9450 16270
rect 9470 16250 9480 16270
rect 9440 16240 9480 16250
rect 9520 16240 9560 16440
rect 9600 16240 9640 16440
rect 9680 16240 9720 16440
rect 9760 16240 9800 16440
rect 9840 16240 9880 16440
rect 9920 16240 9960 16440
rect 10000 16240 10040 16440
rect 10080 16240 10120 16440
rect 10160 16240 10200 16440
rect 10240 16240 10280 16440
rect 10320 16240 10360 16440
rect 10400 16240 10440 16440
rect 10480 16240 10520 16440
rect 10560 16240 10600 16440
rect 10640 16240 10680 16440
rect 10720 16240 10760 16440
rect 10800 16240 10840 16440
rect 10880 16240 10920 16440
rect 10960 16240 11000 16440
rect 11040 16240 11080 16440
rect 11120 16240 11160 16440
rect 11200 16240 11240 16440
rect 11280 16240 11320 16440
rect 11360 16240 11400 16440
rect 11440 16240 11480 16440
rect 11560 16430 11600 16440
rect 11560 16410 11570 16430
rect 11590 16410 11600 16430
rect 11560 16270 11600 16410
rect 11560 16250 11570 16270
rect 11590 16250 11600 16270
rect 11560 16240 11600 16250
rect 11640 16430 11680 16440
rect 11640 16410 11650 16430
rect 11670 16410 11680 16430
rect 11640 16270 11680 16410
rect 11640 16250 11650 16270
rect 11670 16250 11680 16270
rect 11640 16240 11680 16250
rect 11720 16430 11760 16440
rect 11720 16410 11730 16430
rect 11750 16410 11760 16430
rect 11720 16270 11760 16410
rect 11720 16250 11730 16270
rect 11750 16250 11760 16270
rect 11720 16240 11760 16250
rect 11800 16430 11840 16440
rect 11800 16410 11810 16430
rect 11830 16410 11840 16430
rect 11800 16270 11840 16410
rect 11800 16250 11810 16270
rect 11830 16250 11840 16270
rect 11800 16240 11840 16250
rect 11880 16430 11920 16440
rect 11880 16410 11890 16430
rect 11910 16410 11920 16430
rect 11880 16270 11920 16410
rect 11880 16250 11890 16270
rect 11910 16250 11920 16270
rect 11880 16240 11920 16250
rect 11960 16430 12000 16440
rect 11960 16410 11970 16430
rect 11990 16410 12000 16430
rect 11960 16270 12000 16410
rect 11960 16250 11970 16270
rect 11990 16250 12000 16270
rect 11960 16240 12000 16250
rect 12040 16430 12080 16440
rect 12040 16410 12050 16430
rect 12070 16410 12080 16430
rect 12040 16270 12080 16410
rect 12040 16250 12050 16270
rect 12070 16250 12080 16270
rect 12040 16240 12080 16250
rect 12120 16430 12160 16440
rect 12120 16410 12130 16430
rect 12150 16410 12160 16430
rect 12120 16270 12160 16410
rect 12120 16250 12130 16270
rect 12150 16250 12160 16270
rect 12120 16240 12160 16250
rect 12200 16430 12240 16440
rect 12200 16410 12210 16430
rect 12230 16410 12240 16430
rect 12200 16270 12240 16410
rect 12200 16250 12210 16270
rect 12230 16250 12240 16270
rect 12200 16240 12240 16250
rect 12280 16430 12320 16440
rect 12280 16410 12290 16430
rect 12310 16410 12320 16430
rect 12280 16270 12320 16410
rect 12280 16250 12290 16270
rect 12310 16250 12320 16270
rect 12280 16240 12320 16250
rect 12360 16430 12400 16440
rect 12360 16410 12370 16430
rect 12390 16410 12400 16430
rect 12360 16270 12400 16410
rect 12360 16250 12370 16270
rect 12390 16250 12400 16270
rect 12360 16240 12400 16250
rect 12440 16430 12480 16440
rect 12440 16410 12450 16430
rect 12470 16410 12480 16430
rect 12440 16270 12480 16410
rect 12440 16250 12450 16270
rect 12470 16250 12480 16270
rect 12440 16240 12480 16250
rect 12520 16430 12560 16440
rect 12520 16410 12530 16430
rect 12550 16410 12560 16430
rect 12520 16270 12560 16410
rect 12520 16250 12530 16270
rect 12550 16250 12560 16270
rect 12520 16240 12560 16250
rect 12600 16430 12640 16440
rect 12600 16410 12610 16430
rect 12630 16410 12640 16430
rect 12600 16270 12640 16410
rect 12600 16250 12610 16270
rect 12630 16250 12640 16270
rect 12600 16240 12640 16250
rect 12680 16430 12720 16440
rect 12680 16410 12690 16430
rect 12710 16410 12720 16430
rect 12680 16270 12720 16410
rect 12680 16250 12690 16270
rect 12710 16250 12720 16270
rect 12680 16240 12720 16250
rect 12760 16430 12800 16440
rect 12760 16410 12770 16430
rect 12790 16410 12800 16430
rect 12760 16270 12800 16410
rect 12760 16250 12770 16270
rect 12790 16250 12800 16270
rect 12760 16240 12800 16250
rect 12840 16430 12880 16440
rect 12840 16410 12850 16430
rect 12870 16410 12880 16430
rect 12840 16270 12880 16410
rect 12840 16250 12850 16270
rect 12870 16250 12880 16270
rect 12840 16240 12880 16250
rect 12920 16430 12960 16440
rect 12920 16410 12930 16430
rect 12950 16410 12960 16430
rect 12920 16270 12960 16410
rect 12920 16250 12930 16270
rect 12950 16250 12960 16270
rect 12920 16240 12960 16250
rect 13000 16430 13040 16440
rect 13000 16410 13010 16430
rect 13030 16410 13040 16430
rect 13000 16270 13040 16410
rect 13000 16250 13010 16270
rect 13030 16250 13040 16270
rect 13000 16240 13040 16250
rect 13080 16430 13120 16440
rect 13080 16410 13090 16430
rect 13110 16410 13120 16430
rect 13080 16270 13120 16410
rect 13080 16250 13090 16270
rect 13110 16250 13120 16270
rect 13080 16240 13120 16250
rect 13160 16430 13200 16440
rect 13160 16410 13170 16430
rect 13190 16410 13200 16430
rect 13160 16270 13200 16410
rect 13160 16250 13170 16270
rect 13190 16250 13200 16270
rect 13160 16240 13200 16250
rect 13240 16430 13280 16440
rect 13240 16410 13250 16430
rect 13270 16410 13280 16430
rect 13240 16270 13280 16410
rect 13240 16250 13250 16270
rect 13270 16250 13280 16270
rect 13240 16240 13280 16250
rect 13320 16430 13360 16440
rect 13320 16410 13330 16430
rect 13350 16410 13360 16430
rect 13320 16270 13360 16410
rect 13320 16250 13330 16270
rect 13350 16250 13360 16270
rect 13320 16240 13360 16250
rect 13400 16430 13440 16440
rect 13400 16410 13410 16430
rect 13430 16410 13440 16430
rect 13400 16270 13440 16410
rect 13400 16250 13410 16270
rect 13430 16250 13440 16270
rect 13400 16240 13440 16250
rect 13480 16430 13520 16440
rect 13480 16410 13490 16430
rect 13510 16410 13520 16430
rect 13480 16270 13520 16410
rect 13480 16250 13490 16270
rect 13510 16250 13520 16270
rect 13480 16240 13520 16250
rect 13560 16430 13600 16440
rect 13560 16410 13570 16430
rect 13590 16410 13600 16430
rect 13560 16270 13600 16410
rect 13560 16250 13570 16270
rect 13590 16250 13600 16270
rect 13560 16240 13600 16250
rect 13640 16430 13680 16440
rect 13640 16410 13650 16430
rect 13670 16410 13680 16430
rect 13640 16270 13680 16410
rect 13640 16250 13650 16270
rect 13670 16250 13680 16270
rect 13640 16240 13680 16250
rect 13720 16430 13760 16440
rect 13720 16410 13730 16430
rect 13750 16410 13760 16430
rect 13720 16270 13760 16410
rect 13720 16250 13730 16270
rect 13750 16250 13760 16270
rect 13720 16240 13760 16250
rect 13800 16430 13840 16440
rect 13800 16410 13810 16430
rect 13830 16410 13840 16430
rect 13800 16270 13840 16410
rect 13800 16250 13810 16270
rect 13830 16250 13840 16270
rect 13800 16240 13840 16250
rect 13880 16430 13920 16440
rect 13880 16410 13890 16430
rect 13910 16410 13920 16430
rect 13880 16270 13920 16410
rect 13880 16250 13890 16270
rect 13910 16250 13920 16270
rect 13880 16240 13920 16250
rect 13960 16430 14000 16440
rect 13960 16410 13970 16430
rect 13990 16410 14000 16430
rect 13960 16270 14000 16410
rect 13960 16250 13970 16270
rect 13990 16250 14000 16270
rect 13960 16240 14000 16250
rect 14040 16430 14080 16440
rect 14040 16410 14050 16430
rect 14070 16410 14080 16430
rect 14040 16270 14080 16410
rect 14040 16250 14050 16270
rect 14070 16250 14080 16270
rect 14040 16240 14080 16250
rect 14120 16430 14160 16440
rect 14120 16410 14130 16430
rect 14150 16410 14160 16430
rect 14120 16270 14160 16410
rect 14120 16250 14130 16270
rect 14150 16250 14160 16270
rect 14120 16240 14160 16250
rect 14200 16430 14240 16440
rect 14200 16410 14210 16430
rect 14230 16410 14240 16430
rect 14200 16270 14240 16410
rect 14200 16250 14210 16270
rect 14230 16250 14240 16270
rect 14200 16240 14240 16250
rect 14280 16430 14320 16440
rect 14280 16410 14290 16430
rect 14310 16410 14320 16430
rect 14280 16270 14320 16410
rect 14280 16250 14290 16270
rect 14310 16250 14320 16270
rect 14280 16240 14320 16250
rect 14360 16430 14400 16440
rect 14360 16410 14370 16430
rect 14390 16410 14400 16430
rect 14360 16270 14400 16410
rect 14360 16250 14370 16270
rect 14390 16250 14400 16270
rect 14360 16240 14400 16250
rect 14440 16430 14480 16440
rect 14440 16410 14450 16430
rect 14470 16410 14480 16430
rect 14440 16270 14480 16410
rect 14440 16250 14450 16270
rect 14470 16250 14480 16270
rect 14440 16240 14480 16250
rect 14520 16430 14560 16440
rect 14520 16410 14530 16430
rect 14550 16410 14560 16430
rect 14520 16270 14560 16410
rect 14520 16250 14530 16270
rect 14550 16250 14560 16270
rect 14520 16240 14560 16250
rect 14600 16430 14640 16440
rect 14600 16410 14610 16430
rect 14630 16410 14640 16430
rect 14600 16270 14640 16410
rect 14600 16250 14610 16270
rect 14630 16250 14640 16270
rect 14600 16240 14640 16250
rect 14680 16430 14720 16440
rect 14680 16410 14690 16430
rect 14710 16410 14720 16430
rect 14680 16270 14720 16410
rect 14680 16250 14690 16270
rect 14710 16250 14720 16270
rect 14680 16240 14720 16250
rect 14760 16240 14800 16440
rect 14840 16240 14880 16440
rect 14920 16240 14960 16440
rect 15000 16240 15040 16440
rect 15080 16240 15120 16440
rect 15160 16240 15200 16440
rect 15240 16240 15280 16440
rect 15320 16240 15360 16440
rect 15400 16240 15440 16440
rect 15480 16240 15520 16440
rect 15560 16240 15600 16440
rect 15640 16240 15680 16440
rect 15720 16240 15760 16440
rect 15800 16240 15840 16440
rect 15880 16240 15920 16440
rect 15960 16240 16000 16440
rect 16040 16240 16080 16440
rect 16120 16240 16160 16440
rect 16200 16240 16240 16440
rect 16280 16240 16320 16440
rect 16360 16240 16400 16440
rect 16440 16240 16480 16440
rect 16520 16240 16560 16440
rect 16600 16240 16640 16440
rect 16680 16240 16720 16440
rect 16760 16430 16800 16440
rect 16760 16410 16770 16430
rect 16790 16410 16800 16430
rect 16760 16270 16800 16410
rect 16760 16250 16770 16270
rect 16790 16250 16800 16270
rect 16760 16240 16800 16250
rect 16840 16430 16880 16440
rect 16840 16410 16850 16430
rect 16870 16410 16880 16430
rect 16840 16270 16880 16410
rect 16840 16250 16850 16270
rect 16870 16250 16880 16270
rect 16840 16240 16880 16250
rect 16920 16430 16960 16440
rect 16920 16410 16930 16430
rect 16950 16410 16960 16430
rect 16920 16270 16960 16410
rect 16920 16250 16930 16270
rect 16950 16250 16960 16270
rect 16920 16240 16960 16250
rect 17000 16430 17040 16440
rect 17000 16410 17010 16430
rect 17030 16410 17040 16430
rect 17000 16270 17040 16410
rect 17000 16250 17010 16270
rect 17030 16250 17040 16270
rect 17000 16240 17040 16250
rect 17080 16430 17120 16440
rect 17080 16410 17090 16430
rect 17110 16410 17120 16430
rect 17080 16270 17120 16410
rect 17080 16250 17090 16270
rect 17110 16250 17120 16270
rect 17080 16240 17120 16250
rect 17160 16430 17200 16440
rect 17160 16410 17170 16430
rect 17190 16410 17200 16430
rect 17160 16270 17200 16410
rect 17160 16250 17170 16270
rect 17190 16250 17200 16270
rect 17160 16240 17200 16250
rect 17240 16430 17280 16440
rect 17240 16410 17250 16430
rect 17270 16410 17280 16430
rect 17240 16270 17280 16410
rect 17240 16250 17250 16270
rect 17270 16250 17280 16270
rect 17240 16240 17280 16250
rect 17320 16430 17360 16440
rect 17320 16410 17330 16430
rect 17350 16410 17360 16430
rect 17320 16270 17360 16410
rect 17320 16250 17330 16270
rect 17350 16250 17360 16270
rect 17320 16240 17360 16250
rect 17400 16430 17440 16440
rect 17400 16410 17410 16430
rect 17430 16410 17440 16430
rect 17400 16270 17440 16410
rect 17400 16250 17410 16270
rect 17430 16250 17440 16270
rect 17400 16240 17440 16250
rect 17480 16430 17520 16440
rect 17480 16410 17490 16430
rect 17510 16410 17520 16430
rect 17480 16270 17520 16410
rect 17480 16250 17490 16270
rect 17510 16250 17520 16270
rect 17480 16240 17520 16250
rect 17560 16430 17600 16440
rect 17560 16410 17570 16430
rect 17590 16410 17600 16430
rect 17560 16270 17600 16410
rect 17560 16250 17570 16270
rect 17590 16250 17600 16270
rect 17560 16240 17600 16250
rect 17640 16430 17680 16440
rect 17640 16410 17650 16430
rect 17670 16410 17680 16430
rect 17640 16270 17680 16410
rect 17640 16250 17650 16270
rect 17670 16250 17680 16270
rect 17640 16240 17680 16250
rect 17720 16430 17760 16440
rect 17720 16410 17730 16430
rect 17750 16410 17760 16430
rect 17720 16270 17760 16410
rect 17720 16250 17730 16270
rect 17750 16250 17760 16270
rect 17720 16240 17760 16250
rect 17800 16430 17840 16440
rect 17800 16410 17810 16430
rect 17830 16410 17840 16430
rect 17800 16270 17840 16410
rect 17800 16250 17810 16270
rect 17830 16250 17840 16270
rect 17800 16240 17840 16250
rect 17880 16430 17920 16440
rect 17880 16410 17890 16430
rect 17910 16410 17920 16430
rect 17880 16270 17920 16410
rect 17880 16250 17890 16270
rect 17910 16250 17920 16270
rect 17880 16240 17920 16250
rect 17960 16430 18000 16440
rect 17960 16410 17970 16430
rect 17990 16410 18000 16430
rect 17960 16270 18000 16410
rect 17960 16250 17970 16270
rect 17990 16250 18000 16270
rect 17960 16240 18000 16250
rect 18040 16430 18080 16440
rect 18040 16410 18050 16430
rect 18070 16410 18080 16430
rect 18040 16270 18080 16410
rect 18040 16250 18050 16270
rect 18070 16250 18080 16270
rect 18040 16240 18080 16250
rect 18120 16430 18160 16440
rect 18120 16410 18130 16430
rect 18150 16410 18160 16430
rect 18120 16270 18160 16410
rect 18120 16250 18130 16270
rect 18150 16250 18160 16270
rect 18120 16240 18160 16250
rect 18200 16430 18240 16440
rect 18200 16410 18210 16430
rect 18230 16410 18240 16430
rect 18200 16270 18240 16410
rect 18200 16250 18210 16270
rect 18230 16250 18240 16270
rect 18200 16240 18240 16250
rect 18280 16430 18320 16440
rect 18280 16410 18290 16430
rect 18310 16410 18320 16430
rect 18280 16270 18320 16410
rect 18280 16250 18290 16270
rect 18310 16250 18320 16270
rect 18280 16240 18320 16250
rect 18360 16430 18400 16440
rect 18360 16410 18370 16430
rect 18390 16410 18400 16430
rect 18360 16270 18400 16410
rect 18360 16250 18370 16270
rect 18390 16250 18400 16270
rect 18360 16240 18400 16250
rect 18440 16430 18480 16440
rect 18440 16410 18450 16430
rect 18470 16410 18480 16430
rect 18440 16270 18480 16410
rect 18440 16250 18450 16270
rect 18470 16250 18480 16270
rect 18440 16240 18480 16250
rect 18520 16430 18560 16440
rect 18520 16410 18530 16430
rect 18550 16410 18560 16430
rect 18520 16270 18560 16410
rect 18520 16250 18530 16270
rect 18550 16250 18560 16270
rect 18520 16240 18560 16250
rect 18600 16430 18640 16440
rect 18600 16410 18610 16430
rect 18630 16410 18640 16430
rect 18600 16270 18640 16410
rect 18600 16250 18610 16270
rect 18630 16250 18640 16270
rect 18600 16240 18640 16250
rect 18680 16430 18720 16440
rect 18680 16410 18690 16430
rect 18710 16410 18720 16430
rect 18680 16270 18720 16410
rect 18680 16250 18690 16270
rect 18710 16250 18720 16270
rect 18680 16240 18720 16250
rect 18760 16430 18800 16440
rect 18760 16410 18770 16430
rect 18790 16410 18800 16430
rect 18760 16270 18800 16410
rect 18760 16250 18770 16270
rect 18790 16250 18800 16270
rect 18760 16240 18800 16250
rect 18840 16430 18880 16440
rect 18840 16410 18850 16430
rect 18870 16410 18880 16430
rect 18840 16270 18880 16410
rect 18840 16250 18850 16270
rect 18870 16250 18880 16270
rect 18840 16240 18880 16250
rect 18920 16430 18960 16440
rect 18920 16410 18930 16430
rect 18950 16410 18960 16430
rect 18920 16270 18960 16410
rect 18920 16250 18930 16270
rect 18950 16250 18960 16270
rect 18920 16240 18960 16250
rect 19000 16430 19040 16440
rect 19000 16410 19010 16430
rect 19030 16410 19040 16430
rect 19000 16270 19040 16410
rect 19000 16250 19010 16270
rect 19030 16250 19040 16270
rect 19000 16240 19040 16250
rect 19080 16430 19120 16440
rect 19080 16410 19090 16430
rect 19110 16410 19120 16430
rect 19080 16270 19120 16410
rect 19080 16250 19090 16270
rect 19110 16250 19120 16270
rect 19080 16240 19120 16250
rect 19160 16430 19200 16440
rect 19160 16410 19170 16430
rect 19190 16410 19200 16430
rect 19160 16270 19200 16410
rect 19160 16250 19170 16270
rect 19190 16250 19200 16270
rect 19160 16240 19200 16250
rect 19240 16430 19280 16440
rect 19240 16410 19250 16430
rect 19270 16410 19280 16430
rect 19240 16270 19280 16410
rect 19240 16250 19250 16270
rect 19270 16250 19280 16270
rect 19240 16240 19280 16250
rect 19320 16430 19360 16440
rect 19320 16410 19330 16430
rect 19350 16410 19360 16430
rect 19320 16270 19360 16410
rect 19320 16250 19330 16270
rect 19350 16250 19360 16270
rect 19320 16240 19360 16250
rect 19400 16430 19440 16440
rect 19400 16410 19410 16430
rect 19430 16410 19440 16430
rect 19400 16270 19440 16410
rect 19400 16250 19410 16270
rect 19430 16250 19440 16270
rect 19400 16240 19440 16250
rect 19480 16430 19520 16440
rect 19480 16410 19490 16430
rect 19510 16410 19520 16430
rect 19480 16270 19520 16410
rect 19480 16250 19490 16270
rect 19510 16250 19520 16270
rect 19480 16240 19520 16250
rect 19560 16430 19600 16440
rect 19560 16410 19570 16430
rect 19590 16410 19600 16430
rect 19560 16270 19600 16410
rect 19560 16250 19570 16270
rect 19590 16250 19600 16270
rect 19560 16240 19600 16250
rect 19640 16430 19680 16440
rect 19640 16410 19650 16430
rect 19670 16410 19680 16430
rect 19640 16270 19680 16410
rect 19640 16250 19650 16270
rect 19670 16250 19680 16270
rect 19640 16240 19680 16250
rect 19720 16430 19760 16440
rect 19720 16410 19730 16430
rect 19750 16410 19760 16430
rect 19720 16270 19760 16410
rect 19720 16250 19730 16270
rect 19750 16250 19760 16270
rect 19720 16240 19760 16250
rect 19800 16430 19840 16440
rect 19800 16410 19810 16430
rect 19830 16410 19840 16430
rect 19800 16270 19840 16410
rect 19800 16250 19810 16270
rect 19830 16250 19840 16270
rect 19800 16240 19840 16250
rect 19880 16430 19920 16440
rect 19880 16410 19890 16430
rect 19910 16410 19920 16430
rect 19880 16270 19920 16410
rect 19880 16250 19890 16270
rect 19910 16250 19920 16270
rect 19880 16240 19920 16250
rect 19960 16430 20000 16440
rect 19960 16410 19970 16430
rect 19990 16410 20000 16430
rect 19960 16270 20000 16410
rect 19960 16250 19970 16270
rect 19990 16250 20000 16270
rect 19960 16240 20000 16250
rect 20040 16430 20080 16440
rect 20040 16410 20050 16430
rect 20070 16410 20080 16430
rect 20040 16270 20080 16410
rect 20040 16250 20050 16270
rect 20070 16250 20080 16270
rect 20040 16240 20080 16250
rect 20120 16430 20160 16440
rect 20120 16410 20130 16430
rect 20150 16410 20160 16430
rect 20120 16270 20160 16410
rect 20120 16250 20130 16270
rect 20150 16250 20160 16270
rect 20120 16240 20160 16250
rect 20200 16430 20240 16440
rect 20200 16410 20210 16430
rect 20230 16410 20240 16430
rect 20200 16270 20240 16410
rect 20200 16250 20210 16270
rect 20230 16250 20240 16270
rect 20200 16240 20240 16250
rect 20280 16430 20320 16440
rect 20280 16410 20290 16430
rect 20310 16410 20320 16430
rect 20280 16270 20320 16410
rect 20280 16250 20290 16270
rect 20310 16250 20320 16270
rect 20280 16240 20320 16250
rect 20360 16430 20400 16440
rect 20360 16410 20370 16430
rect 20390 16410 20400 16430
rect 20360 16270 20400 16410
rect 20360 16250 20370 16270
rect 20390 16250 20400 16270
rect 20360 16240 20400 16250
rect 20440 16430 20480 16440
rect 20440 16410 20450 16430
rect 20470 16410 20480 16430
rect 20440 16270 20480 16410
rect 20440 16250 20450 16270
rect 20470 16250 20480 16270
rect 20440 16240 20480 16250
rect 20520 16430 20560 16440
rect 20520 16410 20530 16430
rect 20550 16410 20560 16430
rect 20520 16270 20560 16410
rect 20520 16250 20530 16270
rect 20550 16250 20560 16270
rect 20520 16240 20560 16250
rect 20600 16430 20640 16440
rect 20600 16410 20610 16430
rect 20630 16410 20640 16430
rect 20600 16270 20640 16410
rect 20600 16250 20610 16270
rect 20630 16250 20640 16270
rect 20600 16240 20640 16250
rect 20680 16430 20720 16440
rect 20680 16410 20690 16430
rect 20710 16410 20720 16430
rect 20680 16270 20720 16410
rect 20680 16250 20690 16270
rect 20710 16250 20720 16270
rect 20680 16240 20720 16250
rect 20760 16430 20800 16440
rect 20760 16410 20770 16430
rect 20790 16410 20800 16430
rect 20760 16270 20800 16410
rect 20760 16250 20770 16270
rect 20790 16250 20800 16270
rect 20760 16240 20800 16250
rect 20840 16430 20880 16440
rect 20840 16410 20850 16430
rect 20870 16410 20880 16430
rect 20840 16270 20880 16410
rect 20840 16250 20850 16270
rect 20870 16250 20880 16270
rect 20840 16240 20880 16250
rect 20920 16430 20960 16440
rect 20920 16410 20930 16430
rect 20950 16410 20960 16430
rect 20920 16270 20960 16410
rect 20920 16250 20930 16270
rect 20950 16250 20960 16270
rect 20920 16240 20960 16250
rect 0 16190 40 16200
rect 0 16170 10 16190
rect 30 16170 40 16190
rect 0 16030 40 16170
rect 0 16010 10 16030
rect 30 16010 40 16030
rect 0 15870 40 16010
rect 0 15850 10 15870
rect 30 15850 40 15870
rect 0 15710 40 15850
rect 0 15690 10 15710
rect 30 15690 40 15710
rect 0 15550 40 15690
rect 0 15530 10 15550
rect 30 15530 40 15550
rect 0 15390 40 15530
rect 0 15370 10 15390
rect 30 15370 40 15390
rect 0 15230 40 15370
rect 0 15210 10 15230
rect 30 15210 40 15230
rect 0 15200 40 15210
rect 80 16190 120 16200
rect 80 16170 90 16190
rect 110 16170 120 16190
rect 80 16030 120 16170
rect 80 16010 90 16030
rect 110 16010 120 16030
rect 80 15870 120 16010
rect 80 15850 90 15870
rect 110 15850 120 15870
rect 80 15710 120 15850
rect 80 15690 90 15710
rect 110 15690 120 15710
rect 80 15550 120 15690
rect 80 15530 90 15550
rect 110 15530 120 15550
rect 80 15390 120 15530
rect 80 15370 90 15390
rect 110 15370 120 15390
rect 80 15230 120 15370
rect 80 15210 90 15230
rect 110 15210 120 15230
rect 80 15200 120 15210
rect 160 16190 200 16200
rect 160 16170 170 16190
rect 190 16170 200 16190
rect 160 16030 200 16170
rect 160 16010 170 16030
rect 190 16010 200 16030
rect 160 15870 200 16010
rect 160 15850 170 15870
rect 190 15850 200 15870
rect 160 15710 200 15850
rect 160 15690 170 15710
rect 190 15690 200 15710
rect 160 15550 200 15690
rect 160 15530 170 15550
rect 190 15530 200 15550
rect 160 15390 200 15530
rect 160 15370 170 15390
rect 190 15370 200 15390
rect 160 15230 200 15370
rect 160 15210 170 15230
rect 190 15210 200 15230
rect 160 15200 200 15210
rect 240 16190 280 16200
rect 240 16170 250 16190
rect 270 16170 280 16190
rect 240 16030 280 16170
rect 240 16010 250 16030
rect 270 16010 280 16030
rect 240 15870 280 16010
rect 240 15850 250 15870
rect 270 15850 280 15870
rect 240 15710 280 15850
rect 240 15690 250 15710
rect 270 15690 280 15710
rect 240 15550 280 15690
rect 240 15530 250 15550
rect 270 15530 280 15550
rect 240 15390 280 15530
rect 240 15370 250 15390
rect 270 15370 280 15390
rect 240 15230 280 15370
rect 240 15210 250 15230
rect 270 15210 280 15230
rect 240 15200 280 15210
rect 320 16190 360 16200
rect 320 16170 330 16190
rect 350 16170 360 16190
rect 320 16030 360 16170
rect 320 16010 330 16030
rect 350 16010 360 16030
rect 320 15870 360 16010
rect 320 15850 330 15870
rect 350 15850 360 15870
rect 320 15710 360 15850
rect 320 15690 330 15710
rect 350 15690 360 15710
rect 320 15550 360 15690
rect 320 15530 330 15550
rect 350 15530 360 15550
rect 320 15390 360 15530
rect 320 15370 330 15390
rect 350 15370 360 15390
rect 320 15230 360 15370
rect 320 15210 330 15230
rect 350 15210 360 15230
rect 320 15200 360 15210
rect 400 16190 440 16200
rect 400 16170 410 16190
rect 430 16170 440 16190
rect 400 16030 440 16170
rect 400 16010 410 16030
rect 430 16010 440 16030
rect 400 15870 440 16010
rect 400 15850 410 15870
rect 430 15850 440 15870
rect 400 15710 440 15850
rect 400 15690 410 15710
rect 430 15690 440 15710
rect 400 15550 440 15690
rect 400 15530 410 15550
rect 430 15530 440 15550
rect 400 15390 440 15530
rect 400 15370 410 15390
rect 430 15370 440 15390
rect 400 15230 440 15370
rect 400 15210 410 15230
rect 430 15210 440 15230
rect 400 15200 440 15210
rect 480 16190 520 16200
rect 480 16170 490 16190
rect 510 16170 520 16190
rect 480 16030 520 16170
rect 480 16010 490 16030
rect 510 16010 520 16030
rect 480 15870 520 16010
rect 480 15850 490 15870
rect 510 15850 520 15870
rect 480 15710 520 15850
rect 480 15690 490 15710
rect 510 15690 520 15710
rect 480 15550 520 15690
rect 480 15530 490 15550
rect 510 15530 520 15550
rect 480 15390 520 15530
rect 480 15370 490 15390
rect 510 15370 520 15390
rect 480 15230 520 15370
rect 480 15210 490 15230
rect 510 15210 520 15230
rect 480 15200 520 15210
rect 560 16190 600 16200
rect 560 16170 570 16190
rect 590 16170 600 16190
rect 560 16030 600 16170
rect 560 16010 570 16030
rect 590 16010 600 16030
rect 560 15870 600 16010
rect 560 15850 570 15870
rect 590 15850 600 15870
rect 560 15710 600 15850
rect 560 15690 570 15710
rect 590 15690 600 15710
rect 560 15550 600 15690
rect 560 15530 570 15550
rect 590 15530 600 15550
rect 560 15390 600 15530
rect 560 15370 570 15390
rect 590 15370 600 15390
rect 560 15230 600 15370
rect 560 15210 570 15230
rect 590 15210 600 15230
rect 560 15200 600 15210
rect 640 16190 680 16200
rect 640 16170 650 16190
rect 670 16170 680 16190
rect 640 16030 680 16170
rect 640 16010 650 16030
rect 670 16010 680 16030
rect 640 15870 680 16010
rect 640 15850 650 15870
rect 670 15850 680 15870
rect 640 15710 680 15850
rect 640 15690 650 15710
rect 670 15690 680 15710
rect 640 15550 680 15690
rect 640 15530 650 15550
rect 670 15530 680 15550
rect 640 15390 680 15530
rect 640 15370 650 15390
rect 670 15370 680 15390
rect 640 15230 680 15370
rect 640 15210 650 15230
rect 670 15210 680 15230
rect 640 15200 680 15210
rect 720 16190 760 16200
rect 720 16170 730 16190
rect 750 16170 760 16190
rect 720 16030 760 16170
rect 720 16010 730 16030
rect 750 16010 760 16030
rect 720 15870 760 16010
rect 720 15850 730 15870
rect 750 15850 760 15870
rect 720 15710 760 15850
rect 720 15690 730 15710
rect 750 15690 760 15710
rect 720 15550 760 15690
rect 720 15530 730 15550
rect 750 15530 760 15550
rect 720 15390 760 15530
rect 720 15370 730 15390
rect 750 15370 760 15390
rect 720 15230 760 15370
rect 720 15210 730 15230
rect 750 15210 760 15230
rect 720 15200 760 15210
rect 800 16190 840 16200
rect 800 16170 810 16190
rect 830 16170 840 16190
rect 800 16030 840 16170
rect 800 16010 810 16030
rect 830 16010 840 16030
rect 800 15870 840 16010
rect 800 15850 810 15870
rect 830 15850 840 15870
rect 800 15710 840 15850
rect 800 15690 810 15710
rect 830 15690 840 15710
rect 800 15550 840 15690
rect 800 15530 810 15550
rect 830 15530 840 15550
rect 800 15390 840 15530
rect 800 15370 810 15390
rect 830 15370 840 15390
rect 800 15230 840 15370
rect 800 15210 810 15230
rect 830 15210 840 15230
rect 800 15200 840 15210
rect 880 16190 920 16200
rect 880 16170 890 16190
rect 910 16170 920 16190
rect 880 16030 920 16170
rect 880 16010 890 16030
rect 910 16010 920 16030
rect 880 15870 920 16010
rect 880 15850 890 15870
rect 910 15850 920 15870
rect 880 15710 920 15850
rect 880 15690 890 15710
rect 910 15690 920 15710
rect 880 15550 920 15690
rect 880 15530 890 15550
rect 910 15530 920 15550
rect 880 15390 920 15530
rect 880 15370 890 15390
rect 910 15370 920 15390
rect 880 15230 920 15370
rect 880 15210 890 15230
rect 910 15210 920 15230
rect 880 15200 920 15210
rect 960 16190 1000 16200
rect 960 16170 970 16190
rect 990 16170 1000 16190
rect 960 16030 1000 16170
rect 960 16010 970 16030
rect 990 16010 1000 16030
rect 960 15870 1000 16010
rect 960 15850 970 15870
rect 990 15850 1000 15870
rect 960 15710 1000 15850
rect 960 15690 970 15710
rect 990 15690 1000 15710
rect 960 15550 1000 15690
rect 960 15530 970 15550
rect 990 15530 1000 15550
rect 960 15390 1000 15530
rect 960 15370 970 15390
rect 990 15370 1000 15390
rect 960 15230 1000 15370
rect 960 15210 970 15230
rect 990 15210 1000 15230
rect 960 15200 1000 15210
rect 1040 16190 1080 16200
rect 1040 16170 1050 16190
rect 1070 16170 1080 16190
rect 1040 16030 1080 16170
rect 1040 16010 1050 16030
rect 1070 16010 1080 16030
rect 1040 15870 1080 16010
rect 1040 15850 1050 15870
rect 1070 15850 1080 15870
rect 1040 15710 1080 15850
rect 1040 15690 1050 15710
rect 1070 15690 1080 15710
rect 1040 15550 1080 15690
rect 1040 15530 1050 15550
rect 1070 15530 1080 15550
rect 1040 15390 1080 15530
rect 1040 15370 1050 15390
rect 1070 15370 1080 15390
rect 1040 15230 1080 15370
rect 1040 15210 1050 15230
rect 1070 15210 1080 15230
rect 1040 15200 1080 15210
rect 1120 16190 1160 16200
rect 1120 16170 1130 16190
rect 1150 16170 1160 16190
rect 1120 16030 1160 16170
rect 1120 16010 1130 16030
rect 1150 16010 1160 16030
rect 1120 15870 1160 16010
rect 1120 15850 1130 15870
rect 1150 15850 1160 15870
rect 1120 15710 1160 15850
rect 1120 15690 1130 15710
rect 1150 15690 1160 15710
rect 1120 15550 1160 15690
rect 1120 15530 1130 15550
rect 1150 15530 1160 15550
rect 1120 15390 1160 15530
rect 1120 15370 1130 15390
rect 1150 15370 1160 15390
rect 1120 15230 1160 15370
rect 1120 15210 1130 15230
rect 1150 15210 1160 15230
rect 1120 15200 1160 15210
rect 1200 16190 1240 16200
rect 1200 16170 1210 16190
rect 1230 16170 1240 16190
rect 1200 16030 1240 16170
rect 1200 16010 1210 16030
rect 1230 16010 1240 16030
rect 1200 15870 1240 16010
rect 1200 15850 1210 15870
rect 1230 15850 1240 15870
rect 1200 15710 1240 15850
rect 1200 15690 1210 15710
rect 1230 15690 1240 15710
rect 1200 15550 1240 15690
rect 1200 15530 1210 15550
rect 1230 15530 1240 15550
rect 1200 15390 1240 15530
rect 1200 15370 1210 15390
rect 1230 15370 1240 15390
rect 1200 15230 1240 15370
rect 1200 15210 1210 15230
rect 1230 15210 1240 15230
rect 1200 15200 1240 15210
rect 1280 16190 1320 16200
rect 1280 16170 1290 16190
rect 1310 16170 1320 16190
rect 1280 16030 1320 16170
rect 1280 16010 1290 16030
rect 1310 16010 1320 16030
rect 1280 15870 1320 16010
rect 1280 15850 1290 15870
rect 1310 15850 1320 15870
rect 1280 15710 1320 15850
rect 1280 15690 1290 15710
rect 1310 15690 1320 15710
rect 1280 15550 1320 15690
rect 1280 15530 1290 15550
rect 1310 15530 1320 15550
rect 1280 15390 1320 15530
rect 1280 15370 1290 15390
rect 1310 15370 1320 15390
rect 1280 15230 1320 15370
rect 1280 15210 1290 15230
rect 1310 15210 1320 15230
rect 1280 15200 1320 15210
rect 1360 16190 1400 16200
rect 1360 16170 1370 16190
rect 1390 16170 1400 16190
rect 1360 16030 1400 16170
rect 1360 16010 1370 16030
rect 1390 16010 1400 16030
rect 1360 15870 1400 16010
rect 1360 15850 1370 15870
rect 1390 15850 1400 15870
rect 1360 15710 1400 15850
rect 1360 15690 1370 15710
rect 1390 15690 1400 15710
rect 1360 15550 1400 15690
rect 1360 15530 1370 15550
rect 1390 15530 1400 15550
rect 1360 15390 1400 15530
rect 1360 15370 1370 15390
rect 1390 15370 1400 15390
rect 1360 15230 1400 15370
rect 1360 15210 1370 15230
rect 1390 15210 1400 15230
rect 1360 15200 1400 15210
rect 1440 16190 1480 16200
rect 1440 16170 1450 16190
rect 1470 16170 1480 16190
rect 1440 16030 1480 16170
rect 1440 16010 1450 16030
rect 1470 16010 1480 16030
rect 1440 15870 1480 16010
rect 1440 15850 1450 15870
rect 1470 15850 1480 15870
rect 1440 15710 1480 15850
rect 1440 15690 1450 15710
rect 1470 15690 1480 15710
rect 1440 15550 1480 15690
rect 1440 15530 1450 15550
rect 1470 15530 1480 15550
rect 1440 15390 1480 15530
rect 1440 15370 1450 15390
rect 1470 15370 1480 15390
rect 1440 15230 1480 15370
rect 1440 15210 1450 15230
rect 1470 15210 1480 15230
rect 1440 15200 1480 15210
rect 1520 16190 1560 16200
rect 1520 16170 1530 16190
rect 1550 16170 1560 16190
rect 1520 16030 1560 16170
rect 1520 16010 1530 16030
rect 1550 16010 1560 16030
rect 1520 15870 1560 16010
rect 1520 15850 1530 15870
rect 1550 15850 1560 15870
rect 1520 15710 1560 15850
rect 1520 15690 1530 15710
rect 1550 15690 1560 15710
rect 1520 15550 1560 15690
rect 1520 15530 1530 15550
rect 1550 15530 1560 15550
rect 1520 15390 1560 15530
rect 1520 15370 1530 15390
rect 1550 15370 1560 15390
rect 1520 15230 1560 15370
rect 1520 15210 1530 15230
rect 1550 15210 1560 15230
rect 1520 15200 1560 15210
rect 1600 16190 1640 16200
rect 1600 16170 1610 16190
rect 1630 16170 1640 16190
rect 1600 16030 1640 16170
rect 1600 16010 1610 16030
rect 1630 16010 1640 16030
rect 1600 15870 1640 16010
rect 1600 15850 1610 15870
rect 1630 15850 1640 15870
rect 1600 15710 1640 15850
rect 1600 15690 1610 15710
rect 1630 15690 1640 15710
rect 1600 15550 1640 15690
rect 1600 15530 1610 15550
rect 1630 15530 1640 15550
rect 1600 15390 1640 15530
rect 1600 15370 1610 15390
rect 1630 15370 1640 15390
rect 1600 15230 1640 15370
rect 1600 15210 1610 15230
rect 1630 15210 1640 15230
rect 1600 15200 1640 15210
rect 1680 16190 1720 16200
rect 1680 16170 1690 16190
rect 1710 16170 1720 16190
rect 1680 16030 1720 16170
rect 1680 16010 1690 16030
rect 1710 16010 1720 16030
rect 1680 15870 1720 16010
rect 1680 15850 1690 15870
rect 1710 15850 1720 15870
rect 1680 15710 1720 15850
rect 1680 15690 1690 15710
rect 1710 15690 1720 15710
rect 1680 15550 1720 15690
rect 1680 15530 1690 15550
rect 1710 15530 1720 15550
rect 1680 15390 1720 15530
rect 1680 15370 1690 15390
rect 1710 15370 1720 15390
rect 1680 15230 1720 15370
rect 1680 15210 1690 15230
rect 1710 15210 1720 15230
rect 1680 15200 1720 15210
rect 1760 16190 1800 16200
rect 1760 16170 1770 16190
rect 1790 16170 1800 16190
rect 1760 16030 1800 16170
rect 1760 16010 1770 16030
rect 1790 16010 1800 16030
rect 1760 15870 1800 16010
rect 1760 15850 1770 15870
rect 1790 15850 1800 15870
rect 1760 15710 1800 15850
rect 1760 15690 1770 15710
rect 1790 15690 1800 15710
rect 1760 15550 1800 15690
rect 1760 15530 1770 15550
rect 1790 15530 1800 15550
rect 1760 15390 1800 15530
rect 1760 15370 1770 15390
rect 1790 15370 1800 15390
rect 1760 15230 1800 15370
rect 1760 15210 1770 15230
rect 1790 15210 1800 15230
rect 1760 15200 1800 15210
rect 1840 16190 1880 16200
rect 1840 16170 1850 16190
rect 1870 16170 1880 16190
rect 1840 16030 1880 16170
rect 1840 16010 1850 16030
rect 1870 16010 1880 16030
rect 1840 15870 1880 16010
rect 1840 15850 1850 15870
rect 1870 15850 1880 15870
rect 1840 15710 1880 15850
rect 1840 15690 1850 15710
rect 1870 15690 1880 15710
rect 1840 15550 1880 15690
rect 1840 15530 1850 15550
rect 1870 15530 1880 15550
rect 1840 15390 1880 15530
rect 1840 15370 1850 15390
rect 1870 15370 1880 15390
rect 1840 15230 1880 15370
rect 1840 15210 1850 15230
rect 1870 15210 1880 15230
rect 1840 15200 1880 15210
rect 1920 16190 1960 16200
rect 1920 16170 1930 16190
rect 1950 16170 1960 16190
rect 1920 16030 1960 16170
rect 1920 16010 1930 16030
rect 1950 16010 1960 16030
rect 1920 15870 1960 16010
rect 1920 15850 1930 15870
rect 1950 15850 1960 15870
rect 1920 15710 1960 15850
rect 1920 15690 1930 15710
rect 1950 15690 1960 15710
rect 1920 15550 1960 15690
rect 1920 15530 1930 15550
rect 1950 15530 1960 15550
rect 1920 15390 1960 15530
rect 1920 15370 1930 15390
rect 1950 15370 1960 15390
rect 1920 15230 1960 15370
rect 1920 15210 1930 15230
rect 1950 15210 1960 15230
rect 1920 15200 1960 15210
rect 2000 16190 2040 16200
rect 2000 16170 2010 16190
rect 2030 16170 2040 16190
rect 2000 16030 2040 16170
rect 2000 16010 2010 16030
rect 2030 16010 2040 16030
rect 2000 15870 2040 16010
rect 2000 15850 2010 15870
rect 2030 15850 2040 15870
rect 2000 15710 2040 15850
rect 2000 15690 2010 15710
rect 2030 15690 2040 15710
rect 2000 15550 2040 15690
rect 2000 15530 2010 15550
rect 2030 15530 2040 15550
rect 2000 15390 2040 15530
rect 2000 15370 2010 15390
rect 2030 15370 2040 15390
rect 2000 15230 2040 15370
rect 2000 15210 2010 15230
rect 2030 15210 2040 15230
rect 2000 15200 2040 15210
rect 2080 16190 2120 16200
rect 2080 16170 2090 16190
rect 2110 16170 2120 16190
rect 2080 16030 2120 16170
rect 2080 16010 2090 16030
rect 2110 16010 2120 16030
rect 2080 15870 2120 16010
rect 2080 15850 2090 15870
rect 2110 15850 2120 15870
rect 2080 15710 2120 15850
rect 2080 15690 2090 15710
rect 2110 15690 2120 15710
rect 2080 15550 2120 15690
rect 2080 15530 2090 15550
rect 2110 15530 2120 15550
rect 2080 15390 2120 15530
rect 2080 15370 2090 15390
rect 2110 15370 2120 15390
rect 2080 15230 2120 15370
rect 2080 15210 2090 15230
rect 2110 15210 2120 15230
rect 2080 15200 2120 15210
rect 2160 16190 2200 16200
rect 2160 16170 2170 16190
rect 2190 16170 2200 16190
rect 2160 16030 2200 16170
rect 2160 16010 2170 16030
rect 2190 16010 2200 16030
rect 2160 15870 2200 16010
rect 2160 15850 2170 15870
rect 2190 15850 2200 15870
rect 2160 15710 2200 15850
rect 2160 15690 2170 15710
rect 2190 15690 2200 15710
rect 2160 15550 2200 15690
rect 2160 15530 2170 15550
rect 2190 15530 2200 15550
rect 2160 15390 2200 15530
rect 2160 15370 2170 15390
rect 2190 15370 2200 15390
rect 2160 15230 2200 15370
rect 2160 15210 2170 15230
rect 2190 15210 2200 15230
rect 2160 15200 2200 15210
rect 2240 16190 2280 16200
rect 2240 16170 2250 16190
rect 2270 16170 2280 16190
rect 2240 16030 2280 16170
rect 2240 16010 2250 16030
rect 2270 16010 2280 16030
rect 2240 15870 2280 16010
rect 2240 15850 2250 15870
rect 2270 15850 2280 15870
rect 2240 15710 2280 15850
rect 2240 15690 2250 15710
rect 2270 15690 2280 15710
rect 2240 15550 2280 15690
rect 2240 15530 2250 15550
rect 2270 15530 2280 15550
rect 2240 15390 2280 15530
rect 2240 15370 2250 15390
rect 2270 15370 2280 15390
rect 2240 15230 2280 15370
rect 2240 15210 2250 15230
rect 2270 15210 2280 15230
rect 2240 15200 2280 15210
rect 2320 16190 2360 16200
rect 2320 16170 2330 16190
rect 2350 16170 2360 16190
rect 2320 16030 2360 16170
rect 2320 16010 2330 16030
rect 2350 16010 2360 16030
rect 2320 15870 2360 16010
rect 2320 15850 2330 15870
rect 2350 15850 2360 15870
rect 2320 15710 2360 15850
rect 2320 15690 2330 15710
rect 2350 15690 2360 15710
rect 2320 15550 2360 15690
rect 2320 15530 2330 15550
rect 2350 15530 2360 15550
rect 2320 15390 2360 15530
rect 2320 15370 2330 15390
rect 2350 15370 2360 15390
rect 2320 15230 2360 15370
rect 2320 15210 2330 15230
rect 2350 15210 2360 15230
rect 2320 15200 2360 15210
rect 2400 16190 2440 16200
rect 2400 16170 2410 16190
rect 2430 16170 2440 16190
rect 2400 16030 2440 16170
rect 2400 16010 2410 16030
rect 2430 16010 2440 16030
rect 2400 15870 2440 16010
rect 2400 15850 2410 15870
rect 2430 15850 2440 15870
rect 2400 15710 2440 15850
rect 2400 15690 2410 15710
rect 2430 15690 2440 15710
rect 2400 15550 2440 15690
rect 2400 15530 2410 15550
rect 2430 15530 2440 15550
rect 2400 15390 2440 15530
rect 2400 15370 2410 15390
rect 2430 15370 2440 15390
rect 2400 15230 2440 15370
rect 2400 15210 2410 15230
rect 2430 15210 2440 15230
rect 2400 15200 2440 15210
rect 2480 16190 2520 16200
rect 2480 16170 2490 16190
rect 2510 16170 2520 16190
rect 2480 16030 2520 16170
rect 2480 16010 2490 16030
rect 2510 16010 2520 16030
rect 2480 15870 2520 16010
rect 2480 15850 2490 15870
rect 2510 15850 2520 15870
rect 2480 15710 2520 15850
rect 2480 15690 2490 15710
rect 2510 15690 2520 15710
rect 2480 15550 2520 15690
rect 2480 15530 2490 15550
rect 2510 15530 2520 15550
rect 2480 15390 2520 15530
rect 2480 15370 2490 15390
rect 2510 15370 2520 15390
rect 2480 15230 2520 15370
rect 2480 15210 2490 15230
rect 2510 15210 2520 15230
rect 2480 15200 2520 15210
rect 2560 16190 2600 16200
rect 2560 16170 2570 16190
rect 2590 16170 2600 16190
rect 2560 16030 2600 16170
rect 2560 16010 2570 16030
rect 2590 16010 2600 16030
rect 2560 15870 2600 16010
rect 2560 15850 2570 15870
rect 2590 15850 2600 15870
rect 2560 15710 2600 15850
rect 2560 15690 2570 15710
rect 2590 15690 2600 15710
rect 2560 15550 2600 15690
rect 2560 15530 2570 15550
rect 2590 15530 2600 15550
rect 2560 15390 2600 15530
rect 2560 15370 2570 15390
rect 2590 15370 2600 15390
rect 2560 15230 2600 15370
rect 2560 15210 2570 15230
rect 2590 15210 2600 15230
rect 2560 15200 2600 15210
rect 2640 16190 2680 16200
rect 2640 16170 2650 16190
rect 2670 16170 2680 16190
rect 2640 16030 2680 16170
rect 2640 16010 2650 16030
rect 2670 16010 2680 16030
rect 2640 15870 2680 16010
rect 2640 15850 2650 15870
rect 2670 15850 2680 15870
rect 2640 15710 2680 15850
rect 2640 15690 2650 15710
rect 2670 15690 2680 15710
rect 2640 15550 2680 15690
rect 2640 15530 2650 15550
rect 2670 15530 2680 15550
rect 2640 15390 2680 15530
rect 2640 15370 2650 15390
rect 2670 15370 2680 15390
rect 2640 15230 2680 15370
rect 2640 15210 2650 15230
rect 2670 15210 2680 15230
rect 2640 15200 2680 15210
rect 2720 16190 2760 16200
rect 2720 16170 2730 16190
rect 2750 16170 2760 16190
rect 2720 16030 2760 16170
rect 2720 16010 2730 16030
rect 2750 16010 2760 16030
rect 2720 15870 2760 16010
rect 2720 15850 2730 15870
rect 2750 15850 2760 15870
rect 2720 15710 2760 15850
rect 2720 15690 2730 15710
rect 2750 15690 2760 15710
rect 2720 15550 2760 15690
rect 2720 15530 2730 15550
rect 2750 15530 2760 15550
rect 2720 15390 2760 15530
rect 2720 15370 2730 15390
rect 2750 15370 2760 15390
rect 2720 15230 2760 15370
rect 2720 15210 2730 15230
rect 2750 15210 2760 15230
rect 2720 15200 2760 15210
rect 2800 16190 2840 16200
rect 2800 16170 2810 16190
rect 2830 16170 2840 16190
rect 2800 16030 2840 16170
rect 2800 16010 2810 16030
rect 2830 16010 2840 16030
rect 2800 15870 2840 16010
rect 2800 15850 2810 15870
rect 2830 15850 2840 15870
rect 2800 15710 2840 15850
rect 2800 15690 2810 15710
rect 2830 15690 2840 15710
rect 2800 15550 2840 15690
rect 2800 15530 2810 15550
rect 2830 15530 2840 15550
rect 2800 15390 2840 15530
rect 2800 15370 2810 15390
rect 2830 15370 2840 15390
rect 2800 15230 2840 15370
rect 2800 15210 2810 15230
rect 2830 15210 2840 15230
rect 2800 15200 2840 15210
rect 2880 16190 2920 16200
rect 2880 16170 2890 16190
rect 2910 16170 2920 16190
rect 2880 16030 2920 16170
rect 2880 16010 2890 16030
rect 2910 16010 2920 16030
rect 2880 15870 2920 16010
rect 2880 15850 2890 15870
rect 2910 15850 2920 15870
rect 2880 15710 2920 15850
rect 2880 15690 2890 15710
rect 2910 15690 2920 15710
rect 2880 15550 2920 15690
rect 2880 15530 2890 15550
rect 2910 15530 2920 15550
rect 2880 15390 2920 15530
rect 2880 15370 2890 15390
rect 2910 15370 2920 15390
rect 2880 15230 2920 15370
rect 2880 15210 2890 15230
rect 2910 15210 2920 15230
rect 2880 15200 2920 15210
rect 2960 16190 3000 16200
rect 2960 16170 2970 16190
rect 2990 16170 3000 16190
rect 2960 16030 3000 16170
rect 2960 16010 2970 16030
rect 2990 16010 3000 16030
rect 2960 15870 3000 16010
rect 2960 15850 2970 15870
rect 2990 15850 3000 15870
rect 2960 15710 3000 15850
rect 2960 15690 2970 15710
rect 2990 15690 3000 15710
rect 2960 15550 3000 15690
rect 2960 15530 2970 15550
rect 2990 15530 3000 15550
rect 2960 15390 3000 15530
rect 2960 15370 2970 15390
rect 2990 15370 3000 15390
rect 2960 15230 3000 15370
rect 2960 15210 2970 15230
rect 2990 15210 3000 15230
rect 2960 15200 3000 15210
rect 3040 16190 3080 16200
rect 3040 16170 3050 16190
rect 3070 16170 3080 16190
rect 3040 16030 3080 16170
rect 3040 16010 3050 16030
rect 3070 16010 3080 16030
rect 3040 15870 3080 16010
rect 3040 15850 3050 15870
rect 3070 15850 3080 15870
rect 3040 15710 3080 15850
rect 3040 15690 3050 15710
rect 3070 15690 3080 15710
rect 3040 15550 3080 15690
rect 3040 15530 3050 15550
rect 3070 15530 3080 15550
rect 3040 15390 3080 15530
rect 3040 15370 3050 15390
rect 3070 15370 3080 15390
rect 3040 15230 3080 15370
rect 3040 15210 3050 15230
rect 3070 15210 3080 15230
rect 3040 15200 3080 15210
rect 3120 16190 3160 16200
rect 3120 16170 3130 16190
rect 3150 16170 3160 16190
rect 3120 16030 3160 16170
rect 3120 16010 3130 16030
rect 3150 16010 3160 16030
rect 3120 15870 3160 16010
rect 3120 15850 3130 15870
rect 3150 15850 3160 15870
rect 3120 15710 3160 15850
rect 3120 15690 3130 15710
rect 3150 15690 3160 15710
rect 3120 15550 3160 15690
rect 3120 15530 3130 15550
rect 3150 15530 3160 15550
rect 3120 15390 3160 15530
rect 3120 15370 3130 15390
rect 3150 15370 3160 15390
rect 3120 15230 3160 15370
rect 3120 15210 3130 15230
rect 3150 15210 3160 15230
rect 3120 15200 3160 15210
rect 3200 16190 3240 16200
rect 3200 16170 3210 16190
rect 3230 16170 3240 16190
rect 3200 16030 3240 16170
rect 3200 16010 3210 16030
rect 3230 16010 3240 16030
rect 3200 15870 3240 16010
rect 3200 15850 3210 15870
rect 3230 15850 3240 15870
rect 3200 15710 3240 15850
rect 3200 15690 3210 15710
rect 3230 15690 3240 15710
rect 3200 15550 3240 15690
rect 3200 15530 3210 15550
rect 3230 15530 3240 15550
rect 3200 15390 3240 15530
rect 3200 15370 3210 15390
rect 3230 15370 3240 15390
rect 3200 15230 3240 15370
rect 3200 15210 3210 15230
rect 3230 15210 3240 15230
rect 3200 15200 3240 15210
rect 3280 16190 3320 16200
rect 3280 16170 3290 16190
rect 3310 16170 3320 16190
rect 3280 16030 3320 16170
rect 3280 16010 3290 16030
rect 3310 16010 3320 16030
rect 3280 15870 3320 16010
rect 3280 15850 3290 15870
rect 3310 15850 3320 15870
rect 3280 15710 3320 15850
rect 3280 15690 3290 15710
rect 3310 15690 3320 15710
rect 3280 15550 3320 15690
rect 3280 15530 3290 15550
rect 3310 15530 3320 15550
rect 3280 15390 3320 15530
rect 3280 15370 3290 15390
rect 3310 15370 3320 15390
rect 3280 15230 3320 15370
rect 3280 15210 3290 15230
rect 3310 15210 3320 15230
rect 3280 15200 3320 15210
rect 3360 16190 3400 16200
rect 3360 16170 3370 16190
rect 3390 16170 3400 16190
rect 3360 16030 3400 16170
rect 3360 16010 3370 16030
rect 3390 16010 3400 16030
rect 3360 15870 3400 16010
rect 3360 15850 3370 15870
rect 3390 15850 3400 15870
rect 3360 15710 3400 15850
rect 3360 15690 3370 15710
rect 3390 15690 3400 15710
rect 3360 15550 3400 15690
rect 3360 15530 3370 15550
rect 3390 15530 3400 15550
rect 3360 15390 3400 15530
rect 3360 15370 3370 15390
rect 3390 15370 3400 15390
rect 3360 15230 3400 15370
rect 3360 15210 3370 15230
rect 3390 15210 3400 15230
rect 3360 15200 3400 15210
rect 3440 16190 3480 16200
rect 3440 16170 3450 16190
rect 3470 16170 3480 16190
rect 3440 16030 3480 16170
rect 3440 16010 3450 16030
rect 3470 16010 3480 16030
rect 3440 15870 3480 16010
rect 3440 15850 3450 15870
rect 3470 15850 3480 15870
rect 3440 15710 3480 15850
rect 3440 15690 3450 15710
rect 3470 15690 3480 15710
rect 3440 15550 3480 15690
rect 3440 15530 3450 15550
rect 3470 15530 3480 15550
rect 3440 15390 3480 15530
rect 3440 15370 3450 15390
rect 3470 15370 3480 15390
rect 3440 15230 3480 15370
rect 3440 15210 3450 15230
rect 3470 15210 3480 15230
rect 3440 15200 3480 15210
rect 3520 16190 3560 16200
rect 3520 16170 3530 16190
rect 3550 16170 3560 16190
rect 3520 16030 3560 16170
rect 3520 16010 3530 16030
rect 3550 16010 3560 16030
rect 3520 15870 3560 16010
rect 3520 15850 3530 15870
rect 3550 15850 3560 15870
rect 3520 15710 3560 15850
rect 3520 15690 3530 15710
rect 3550 15690 3560 15710
rect 3520 15550 3560 15690
rect 3520 15530 3530 15550
rect 3550 15530 3560 15550
rect 3520 15390 3560 15530
rect 3520 15370 3530 15390
rect 3550 15370 3560 15390
rect 3520 15230 3560 15370
rect 3520 15210 3530 15230
rect 3550 15210 3560 15230
rect 3520 15200 3560 15210
rect 3600 16190 3640 16200
rect 3600 16170 3610 16190
rect 3630 16170 3640 16190
rect 3600 16030 3640 16170
rect 3600 16010 3610 16030
rect 3630 16010 3640 16030
rect 3600 15870 3640 16010
rect 3600 15850 3610 15870
rect 3630 15850 3640 15870
rect 3600 15710 3640 15850
rect 3600 15690 3610 15710
rect 3630 15690 3640 15710
rect 3600 15550 3640 15690
rect 3600 15530 3610 15550
rect 3630 15530 3640 15550
rect 3600 15390 3640 15530
rect 3600 15370 3610 15390
rect 3630 15370 3640 15390
rect 3600 15230 3640 15370
rect 3600 15210 3610 15230
rect 3630 15210 3640 15230
rect 3600 15200 3640 15210
rect 3680 16190 3720 16200
rect 3680 16170 3690 16190
rect 3710 16170 3720 16190
rect 3680 16030 3720 16170
rect 3680 16010 3690 16030
rect 3710 16010 3720 16030
rect 3680 15870 3720 16010
rect 3680 15850 3690 15870
rect 3710 15850 3720 15870
rect 3680 15710 3720 15850
rect 3680 15690 3690 15710
rect 3710 15690 3720 15710
rect 3680 15550 3720 15690
rect 3680 15530 3690 15550
rect 3710 15530 3720 15550
rect 3680 15390 3720 15530
rect 3680 15370 3690 15390
rect 3710 15370 3720 15390
rect 3680 15230 3720 15370
rect 3680 15210 3690 15230
rect 3710 15210 3720 15230
rect 3680 15200 3720 15210
rect 3760 16190 3800 16200
rect 3760 16170 3770 16190
rect 3790 16170 3800 16190
rect 3760 16030 3800 16170
rect 3760 16010 3770 16030
rect 3790 16010 3800 16030
rect 3760 15870 3800 16010
rect 3760 15850 3770 15870
rect 3790 15850 3800 15870
rect 3760 15710 3800 15850
rect 3760 15690 3770 15710
rect 3790 15690 3800 15710
rect 3760 15550 3800 15690
rect 3760 15530 3770 15550
rect 3790 15530 3800 15550
rect 3760 15390 3800 15530
rect 3760 15370 3770 15390
rect 3790 15370 3800 15390
rect 3760 15230 3800 15370
rect 3760 15210 3770 15230
rect 3790 15210 3800 15230
rect 3760 15200 3800 15210
rect 3840 16190 3880 16200
rect 3840 16170 3850 16190
rect 3870 16170 3880 16190
rect 3840 16030 3880 16170
rect 3840 16010 3850 16030
rect 3870 16010 3880 16030
rect 3840 15870 3880 16010
rect 3840 15850 3850 15870
rect 3870 15850 3880 15870
rect 3840 15710 3880 15850
rect 3840 15690 3850 15710
rect 3870 15690 3880 15710
rect 3840 15550 3880 15690
rect 3840 15530 3850 15550
rect 3870 15530 3880 15550
rect 3840 15390 3880 15530
rect 3840 15370 3850 15390
rect 3870 15370 3880 15390
rect 3840 15230 3880 15370
rect 3840 15210 3850 15230
rect 3870 15210 3880 15230
rect 3840 15200 3880 15210
rect 3920 16190 3960 16200
rect 3920 16170 3930 16190
rect 3950 16170 3960 16190
rect 3920 16030 3960 16170
rect 3920 16010 3930 16030
rect 3950 16010 3960 16030
rect 3920 15870 3960 16010
rect 3920 15850 3930 15870
rect 3950 15850 3960 15870
rect 3920 15710 3960 15850
rect 3920 15690 3930 15710
rect 3950 15690 3960 15710
rect 3920 15550 3960 15690
rect 3920 15530 3930 15550
rect 3950 15530 3960 15550
rect 3920 15390 3960 15530
rect 3920 15370 3930 15390
rect 3950 15370 3960 15390
rect 3920 15230 3960 15370
rect 3920 15210 3930 15230
rect 3950 15210 3960 15230
rect 3920 15200 3960 15210
rect 4000 16190 4040 16200
rect 4000 16170 4010 16190
rect 4030 16170 4040 16190
rect 4000 16030 4040 16170
rect 4000 16010 4010 16030
rect 4030 16010 4040 16030
rect 4000 15870 4040 16010
rect 4000 15850 4010 15870
rect 4030 15850 4040 15870
rect 4000 15710 4040 15850
rect 4000 15690 4010 15710
rect 4030 15690 4040 15710
rect 4000 15550 4040 15690
rect 4000 15530 4010 15550
rect 4030 15530 4040 15550
rect 4000 15390 4040 15530
rect 4000 15370 4010 15390
rect 4030 15370 4040 15390
rect 4000 15230 4040 15370
rect 4000 15210 4010 15230
rect 4030 15210 4040 15230
rect 4000 15200 4040 15210
rect 4080 16190 4120 16200
rect 4080 16170 4090 16190
rect 4110 16170 4120 16190
rect 4080 16030 4120 16170
rect 4080 16010 4090 16030
rect 4110 16010 4120 16030
rect 4080 15870 4120 16010
rect 4080 15850 4090 15870
rect 4110 15850 4120 15870
rect 4080 15710 4120 15850
rect 4080 15690 4090 15710
rect 4110 15690 4120 15710
rect 4080 15550 4120 15690
rect 4080 15530 4090 15550
rect 4110 15530 4120 15550
rect 4080 15390 4120 15530
rect 4080 15370 4090 15390
rect 4110 15370 4120 15390
rect 4080 15230 4120 15370
rect 4080 15210 4090 15230
rect 4110 15210 4120 15230
rect 4080 15200 4120 15210
rect 4160 16190 4200 16200
rect 4160 16170 4170 16190
rect 4190 16170 4200 16190
rect 4160 16030 4200 16170
rect 4160 16010 4170 16030
rect 4190 16010 4200 16030
rect 4160 15870 4200 16010
rect 4160 15850 4170 15870
rect 4190 15850 4200 15870
rect 4160 15710 4200 15850
rect 4160 15690 4170 15710
rect 4190 15690 4200 15710
rect 4160 15550 4200 15690
rect 4160 15530 4170 15550
rect 4190 15530 4200 15550
rect 4160 15390 4200 15530
rect 4160 15370 4170 15390
rect 4190 15370 4200 15390
rect 4160 15230 4200 15370
rect 4160 15210 4170 15230
rect 4190 15210 4200 15230
rect 4160 15200 4200 15210
rect 4240 15200 4280 16200
rect 4320 15200 4360 16200
rect 4400 15200 4440 16200
rect 4480 15200 4520 16200
rect 4560 15200 4600 16200
rect 4640 15200 4680 16200
rect 4720 15200 4760 16200
rect 4800 15200 4840 16200
rect 4880 15200 4920 16200
rect 4960 15200 5000 16200
rect 5040 15200 5080 16200
rect 5120 15200 5160 16200
rect 5200 15200 5240 16200
rect 5280 15200 5320 16200
rect 5360 15200 5400 16200
rect 5440 15200 5480 16200
rect 5520 15200 5560 16200
rect 5600 15200 5640 16200
rect 5680 15200 5720 16200
rect 5760 15200 5800 16200
rect 5840 15200 5880 16200
rect 5920 15200 5960 16200
rect 6000 15200 6040 16200
rect 6080 15200 6120 16200
rect 6160 15200 6200 16200
rect 6240 16190 6280 16200
rect 6240 16170 6250 16190
rect 6270 16170 6280 16190
rect 6240 16030 6280 16170
rect 6240 16010 6250 16030
rect 6270 16010 6280 16030
rect 6240 15870 6280 16010
rect 6240 15850 6250 15870
rect 6270 15850 6280 15870
rect 6240 15710 6280 15850
rect 6240 15690 6250 15710
rect 6270 15690 6280 15710
rect 6240 15550 6280 15690
rect 6240 15530 6250 15550
rect 6270 15530 6280 15550
rect 6240 15390 6280 15530
rect 6240 15370 6250 15390
rect 6270 15370 6280 15390
rect 6240 15230 6280 15370
rect 6240 15210 6250 15230
rect 6270 15210 6280 15230
rect 6240 15200 6280 15210
rect 6320 16190 6360 16200
rect 6320 16170 6330 16190
rect 6350 16170 6360 16190
rect 6320 16030 6360 16170
rect 6320 16010 6330 16030
rect 6350 16010 6360 16030
rect 6320 15870 6360 16010
rect 6320 15850 6330 15870
rect 6350 15850 6360 15870
rect 6320 15710 6360 15850
rect 6320 15690 6330 15710
rect 6350 15690 6360 15710
rect 6320 15550 6360 15690
rect 6320 15530 6330 15550
rect 6350 15530 6360 15550
rect 6320 15390 6360 15530
rect 6320 15370 6330 15390
rect 6350 15370 6360 15390
rect 6320 15230 6360 15370
rect 6320 15210 6330 15230
rect 6350 15210 6360 15230
rect 6320 15200 6360 15210
rect 6400 16190 6440 16200
rect 6400 16170 6410 16190
rect 6430 16170 6440 16190
rect 6400 16030 6440 16170
rect 6400 16010 6410 16030
rect 6430 16010 6440 16030
rect 6400 15870 6440 16010
rect 6400 15850 6410 15870
rect 6430 15850 6440 15870
rect 6400 15710 6440 15850
rect 6400 15690 6410 15710
rect 6430 15690 6440 15710
rect 6400 15550 6440 15690
rect 6400 15530 6410 15550
rect 6430 15530 6440 15550
rect 6400 15390 6440 15530
rect 6400 15370 6410 15390
rect 6430 15370 6440 15390
rect 6400 15230 6440 15370
rect 6400 15210 6410 15230
rect 6430 15210 6440 15230
rect 6400 15200 6440 15210
rect 6480 16190 6520 16200
rect 6480 16170 6490 16190
rect 6510 16170 6520 16190
rect 6480 16030 6520 16170
rect 6480 16010 6490 16030
rect 6510 16010 6520 16030
rect 6480 15870 6520 16010
rect 6480 15850 6490 15870
rect 6510 15850 6520 15870
rect 6480 15710 6520 15850
rect 6480 15690 6490 15710
rect 6510 15690 6520 15710
rect 6480 15550 6520 15690
rect 6480 15530 6490 15550
rect 6510 15530 6520 15550
rect 6480 15390 6520 15530
rect 6480 15370 6490 15390
rect 6510 15370 6520 15390
rect 6480 15230 6520 15370
rect 6480 15210 6490 15230
rect 6510 15210 6520 15230
rect 6480 15200 6520 15210
rect 6560 16190 6600 16200
rect 6560 16170 6570 16190
rect 6590 16170 6600 16190
rect 6560 16030 6600 16170
rect 6560 16010 6570 16030
rect 6590 16010 6600 16030
rect 6560 15870 6600 16010
rect 6560 15850 6570 15870
rect 6590 15850 6600 15870
rect 6560 15710 6600 15850
rect 6560 15690 6570 15710
rect 6590 15690 6600 15710
rect 6560 15550 6600 15690
rect 6560 15530 6570 15550
rect 6590 15530 6600 15550
rect 6560 15390 6600 15530
rect 6560 15370 6570 15390
rect 6590 15370 6600 15390
rect 6560 15230 6600 15370
rect 6560 15210 6570 15230
rect 6590 15210 6600 15230
rect 6560 15200 6600 15210
rect 6640 16190 6680 16200
rect 6640 16170 6650 16190
rect 6670 16170 6680 16190
rect 6640 16030 6680 16170
rect 6640 16010 6650 16030
rect 6670 16010 6680 16030
rect 6640 15870 6680 16010
rect 6640 15850 6650 15870
rect 6670 15850 6680 15870
rect 6640 15710 6680 15850
rect 6640 15690 6650 15710
rect 6670 15690 6680 15710
rect 6640 15550 6680 15690
rect 6640 15530 6650 15550
rect 6670 15530 6680 15550
rect 6640 15390 6680 15530
rect 6640 15370 6650 15390
rect 6670 15370 6680 15390
rect 6640 15230 6680 15370
rect 6640 15210 6650 15230
rect 6670 15210 6680 15230
rect 6640 15200 6680 15210
rect 6720 16190 6760 16200
rect 6720 16170 6730 16190
rect 6750 16170 6760 16190
rect 6720 16030 6760 16170
rect 6720 16010 6730 16030
rect 6750 16010 6760 16030
rect 6720 15870 6760 16010
rect 6720 15850 6730 15870
rect 6750 15850 6760 15870
rect 6720 15710 6760 15850
rect 6720 15690 6730 15710
rect 6750 15690 6760 15710
rect 6720 15550 6760 15690
rect 6720 15530 6730 15550
rect 6750 15530 6760 15550
rect 6720 15390 6760 15530
rect 6720 15370 6730 15390
rect 6750 15370 6760 15390
rect 6720 15230 6760 15370
rect 6720 15210 6730 15230
rect 6750 15210 6760 15230
rect 6720 15200 6760 15210
rect 6800 16190 6840 16200
rect 6800 16170 6810 16190
rect 6830 16170 6840 16190
rect 6800 16030 6840 16170
rect 6800 16010 6810 16030
rect 6830 16010 6840 16030
rect 6800 15870 6840 16010
rect 6800 15850 6810 15870
rect 6830 15850 6840 15870
rect 6800 15710 6840 15850
rect 6800 15690 6810 15710
rect 6830 15690 6840 15710
rect 6800 15550 6840 15690
rect 6800 15530 6810 15550
rect 6830 15530 6840 15550
rect 6800 15390 6840 15530
rect 6800 15370 6810 15390
rect 6830 15370 6840 15390
rect 6800 15230 6840 15370
rect 6800 15210 6810 15230
rect 6830 15210 6840 15230
rect 6800 15200 6840 15210
rect 6880 16190 6920 16200
rect 6880 16170 6890 16190
rect 6910 16170 6920 16190
rect 6880 16030 6920 16170
rect 6880 16010 6890 16030
rect 6910 16010 6920 16030
rect 6880 15870 6920 16010
rect 6880 15850 6890 15870
rect 6910 15850 6920 15870
rect 6880 15710 6920 15850
rect 6880 15690 6890 15710
rect 6910 15690 6920 15710
rect 6880 15550 6920 15690
rect 6880 15530 6890 15550
rect 6910 15530 6920 15550
rect 6880 15390 6920 15530
rect 6880 15370 6890 15390
rect 6910 15370 6920 15390
rect 6880 15230 6920 15370
rect 6880 15210 6890 15230
rect 6910 15210 6920 15230
rect 6880 15200 6920 15210
rect 6960 16190 7000 16200
rect 6960 16170 6970 16190
rect 6990 16170 7000 16190
rect 6960 16030 7000 16170
rect 6960 16010 6970 16030
rect 6990 16010 7000 16030
rect 6960 15870 7000 16010
rect 6960 15850 6970 15870
rect 6990 15850 7000 15870
rect 6960 15710 7000 15850
rect 6960 15690 6970 15710
rect 6990 15690 7000 15710
rect 6960 15550 7000 15690
rect 6960 15530 6970 15550
rect 6990 15530 7000 15550
rect 6960 15390 7000 15530
rect 6960 15370 6970 15390
rect 6990 15370 7000 15390
rect 6960 15230 7000 15370
rect 6960 15210 6970 15230
rect 6990 15210 7000 15230
rect 6960 15200 7000 15210
rect 7040 16190 7080 16200
rect 7040 16170 7050 16190
rect 7070 16170 7080 16190
rect 7040 16030 7080 16170
rect 7040 16010 7050 16030
rect 7070 16010 7080 16030
rect 7040 15870 7080 16010
rect 7040 15850 7050 15870
rect 7070 15850 7080 15870
rect 7040 15710 7080 15850
rect 7040 15690 7050 15710
rect 7070 15690 7080 15710
rect 7040 15550 7080 15690
rect 7040 15530 7050 15550
rect 7070 15530 7080 15550
rect 7040 15390 7080 15530
rect 7040 15370 7050 15390
rect 7070 15370 7080 15390
rect 7040 15230 7080 15370
rect 7040 15210 7050 15230
rect 7070 15210 7080 15230
rect 7040 15200 7080 15210
rect 7120 16190 7160 16200
rect 7120 16170 7130 16190
rect 7150 16170 7160 16190
rect 7120 16030 7160 16170
rect 7120 16010 7130 16030
rect 7150 16010 7160 16030
rect 7120 15870 7160 16010
rect 7120 15850 7130 15870
rect 7150 15850 7160 15870
rect 7120 15710 7160 15850
rect 7120 15690 7130 15710
rect 7150 15690 7160 15710
rect 7120 15550 7160 15690
rect 7120 15530 7130 15550
rect 7150 15530 7160 15550
rect 7120 15390 7160 15530
rect 7120 15370 7130 15390
rect 7150 15370 7160 15390
rect 7120 15230 7160 15370
rect 7120 15210 7130 15230
rect 7150 15210 7160 15230
rect 7120 15200 7160 15210
rect 7200 16190 7240 16200
rect 7200 16170 7210 16190
rect 7230 16170 7240 16190
rect 7200 16030 7240 16170
rect 7200 16010 7210 16030
rect 7230 16010 7240 16030
rect 7200 15870 7240 16010
rect 7200 15850 7210 15870
rect 7230 15850 7240 15870
rect 7200 15710 7240 15850
rect 7200 15690 7210 15710
rect 7230 15690 7240 15710
rect 7200 15550 7240 15690
rect 7200 15530 7210 15550
rect 7230 15530 7240 15550
rect 7200 15390 7240 15530
rect 7200 15370 7210 15390
rect 7230 15370 7240 15390
rect 7200 15230 7240 15370
rect 7200 15210 7210 15230
rect 7230 15210 7240 15230
rect 7200 15200 7240 15210
rect 7280 16190 7320 16200
rect 7280 16170 7290 16190
rect 7310 16170 7320 16190
rect 7280 16030 7320 16170
rect 7280 16010 7290 16030
rect 7310 16010 7320 16030
rect 7280 15870 7320 16010
rect 7280 15850 7290 15870
rect 7310 15850 7320 15870
rect 7280 15710 7320 15850
rect 7280 15690 7290 15710
rect 7310 15690 7320 15710
rect 7280 15550 7320 15690
rect 7280 15530 7290 15550
rect 7310 15530 7320 15550
rect 7280 15390 7320 15530
rect 7280 15370 7290 15390
rect 7310 15370 7320 15390
rect 7280 15230 7320 15370
rect 7280 15210 7290 15230
rect 7310 15210 7320 15230
rect 7280 15200 7320 15210
rect 7360 16190 7400 16200
rect 7360 16170 7370 16190
rect 7390 16170 7400 16190
rect 7360 16030 7400 16170
rect 7360 16010 7370 16030
rect 7390 16010 7400 16030
rect 7360 15870 7400 16010
rect 7360 15850 7370 15870
rect 7390 15850 7400 15870
rect 7360 15710 7400 15850
rect 7360 15690 7370 15710
rect 7390 15690 7400 15710
rect 7360 15550 7400 15690
rect 7360 15530 7370 15550
rect 7390 15530 7400 15550
rect 7360 15390 7400 15530
rect 7360 15370 7370 15390
rect 7390 15370 7400 15390
rect 7360 15230 7400 15370
rect 7360 15210 7370 15230
rect 7390 15210 7400 15230
rect 7360 15200 7400 15210
rect 7440 16190 7480 16200
rect 7440 16170 7450 16190
rect 7470 16170 7480 16190
rect 7440 16030 7480 16170
rect 7440 16010 7450 16030
rect 7470 16010 7480 16030
rect 7440 15870 7480 16010
rect 7440 15850 7450 15870
rect 7470 15850 7480 15870
rect 7440 15710 7480 15850
rect 7440 15690 7450 15710
rect 7470 15690 7480 15710
rect 7440 15550 7480 15690
rect 7440 15530 7450 15550
rect 7470 15530 7480 15550
rect 7440 15390 7480 15530
rect 7440 15370 7450 15390
rect 7470 15370 7480 15390
rect 7440 15230 7480 15370
rect 7440 15210 7450 15230
rect 7470 15210 7480 15230
rect 7440 15200 7480 15210
rect 7520 16190 7560 16200
rect 7520 16170 7530 16190
rect 7550 16170 7560 16190
rect 7520 16030 7560 16170
rect 7520 16010 7530 16030
rect 7550 16010 7560 16030
rect 7520 15870 7560 16010
rect 7520 15850 7530 15870
rect 7550 15850 7560 15870
rect 7520 15710 7560 15850
rect 7520 15690 7530 15710
rect 7550 15690 7560 15710
rect 7520 15550 7560 15690
rect 7520 15530 7530 15550
rect 7550 15530 7560 15550
rect 7520 15390 7560 15530
rect 7520 15370 7530 15390
rect 7550 15370 7560 15390
rect 7520 15230 7560 15370
rect 7520 15210 7530 15230
rect 7550 15210 7560 15230
rect 7520 15200 7560 15210
rect 7600 16190 7640 16200
rect 7600 16170 7610 16190
rect 7630 16170 7640 16190
rect 7600 16030 7640 16170
rect 7600 16010 7610 16030
rect 7630 16010 7640 16030
rect 7600 15870 7640 16010
rect 7600 15850 7610 15870
rect 7630 15850 7640 15870
rect 7600 15710 7640 15850
rect 7600 15690 7610 15710
rect 7630 15690 7640 15710
rect 7600 15550 7640 15690
rect 7600 15530 7610 15550
rect 7630 15530 7640 15550
rect 7600 15390 7640 15530
rect 7600 15370 7610 15390
rect 7630 15370 7640 15390
rect 7600 15230 7640 15370
rect 7600 15210 7610 15230
rect 7630 15210 7640 15230
rect 7600 15200 7640 15210
rect 7680 16190 7720 16200
rect 7680 16170 7690 16190
rect 7710 16170 7720 16190
rect 7680 16030 7720 16170
rect 7680 16010 7690 16030
rect 7710 16010 7720 16030
rect 7680 15870 7720 16010
rect 7680 15850 7690 15870
rect 7710 15850 7720 15870
rect 7680 15710 7720 15850
rect 7680 15690 7690 15710
rect 7710 15690 7720 15710
rect 7680 15550 7720 15690
rect 7680 15530 7690 15550
rect 7710 15530 7720 15550
rect 7680 15390 7720 15530
rect 7680 15370 7690 15390
rect 7710 15370 7720 15390
rect 7680 15230 7720 15370
rect 7680 15210 7690 15230
rect 7710 15210 7720 15230
rect 7680 15200 7720 15210
rect 7760 16190 7800 16200
rect 7760 16170 7770 16190
rect 7790 16170 7800 16190
rect 7760 16030 7800 16170
rect 7760 16010 7770 16030
rect 7790 16010 7800 16030
rect 7760 15870 7800 16010
rect 7760 15850 7770 15870
rect 7790 15850 7800 15870
rect 7760 15710 7800 15850
rect 7760 15690 7770 15710
rect 7790 15690 7800 15710
rect 7760 15550 7800 15690
rect 7760 15530 7770 15550
rect 7790 15530 7800 15550
rect 7760 15390 7800 15530
rect 7760 15370 7770 15390
rect 7790 15370 7800 15390
rect 7760 15230 7800 15370
rect 7760 15210 7770 15230
rect 7790 15210 7800 15230
rect 7760 15200 7800 15210
rect 7840 16190 7880 16200
rect 7840 16170 7850 16190
rect 7870 16170 7880 16190
rect 7840 16030 7880 16170
rect 7840 16010 7850 16030
rect 7870 16010 7880 16030
rect 7840 15870 7880 16010
rect 7840 15850 7850 15870
rect 7870 15850 7880 15870
rect 7840 15710 7880 15850
rect 7840 15690 7850 15710
rect 7870 15690 7880 15710
rect 7840 15550 7880 15690
rect 7840 15530 7850 15550
rect 7870 15530 7880 15550
rect 7840 15390 7880 15530
rect 7840 15370 7850 15390
rect 7870 15370 7880 15390
rect 7840 15230 7880 15370
rect 7840 15210 7850 15230
rect 7870 15210 7880 15230
rect 7840 15200 7880 15210
rect 7920 16190 7960 16200
rect 7920 16170 7930 16190
rect 7950 16170 7960 16190
rect 7920 16030 7960 16170
rect 7920 16010 7930 16030
rect 7950 16010 7960 16030
rect 7920 15870 7960 16010
rect 7920 15850 7930 15870
rect 7950 15850 7960 15870
rect 7920 15710 7960 15850
rect 7920 15690 7930 15710
rect 7950 15690 7960 15710
rect 7920 15550 7960 15690
rect 7920 15530 7930 15550
rect 7950 15530 7960 15550
rect 7920 15390 7960 15530
rect 7920 15370 7930 15390
rect 7950 15370 7960 15390
rect 7920 15230 7960 15370
rect 7920 15210 7930 15230
rect 7950 15210 7960 15230
rect 7920 15200 7960 15210
rect 8000 16190 8040 16200
rect 8000 16170 8010 16190
rect 8030 16170 8040 16190
rect 8000 16030 8040 16170
rect 8000 16010 8010 16030
rect 8030 16010 8040 16030
rect 8000 15870 8040 16010
rect 8000 15850 8010 15870
rect 8030 15850 8040 15870
rect 8000 15710 8040 15850
rect 8000 15690 8010 15710
rect 8030 15690 8040 15710
rect 8000 15550 8040 15690
rect 8000 15530 8010 15550
rect 8030 15530 8040 15550
rect 8000 15390 8040 15530
rect 8000 15370 8010 15390
rect 8030 15370 8040 15390
rect 8000 15230 8040 15370
rect 8000 15210 8010 15230
rect 8030 15210 8040 15230
rect 8000 15200 8040 15210
rect 8080 16190 8120 16200
rect 8080 16170 8090 16190
rect 8110 16170 8120 16190
rect 8080 16030 8120 16170
rect 8080 16010 8090 16030
rect 8110 16010 8120 16030
rect 8080 15870 8120 16010
rect 8080 15850 8090 15870
rect 8110 15850 8120 15870
rect 8080 15710 8120 15850
rect 8080 15690 8090 15710
rect 8110 15690 8120 15710
rect 8080 15550 8120 15690
rect 8080 15530 8090 15550
rect 8110 15530 8120 15550
rect 8080 15390 8120 15530
rect 8080 15370 8090 15390
rect 8110 15370 8120 15390
rect 8080 15230 8120 15370
rect 8080 15210 8090 15230
rect 8110 15210 8120 15230
rect 8080 15200 8120 15210
rect 8160 16190 8200 16200
rect 8160 16170 8170 16190
rect 8190 16170 8200 16190
rect 8160 16030 8200 16170
rect 8160 16010 8170 16030
rect 8190 16010 8200 16030
rect 8160 15870 8200 16010
rect 8160 15850 8170 15870
rect 8190 15850 8200 15870
rect 8160 15710 8200 15850
rect 8160 15690 8170 15710
rect 8190 15690 8200 15710
rect 8160 15550 8200 15690
rect 8160 15530 8170 15550
rect 8190 15530 8200 15550
rect 8160 15390 8200 15530
rect 8160 15370 8170 15390
rect 8190 15370 8200 15390
rect 8160 15230 8200 15370
rect 8160 15210 8170 15230
rect 8190 15210 8200 15230
rect 8160 15200 8200 15210
rect 8240 16190 8280 16200
rect 8240 16170 8250 16190
rect 8270 16170 8280 16190
rect 8240 16030 8280 16170
rect 8240 16010 8250 16030
rect 8270 16010 8280 16030
rect 8240 15870 8280 16010
rect 8240 15850 8250 15870
rect 8270 15850 8280 15870
rect 8240 15710 8280 15850
rect 8240 15690 8250 15710
rect 8270 15690 8280 15710
rect 8240 15550 8280 15690
rect 8240 15530 8250 15550
rect 8270 15530 8280 15550
rect 8240 15390 8280 15530
rect 8240 15370 8250 15390
rect 8270 15370 8280 15390
rect 8240 15230 8280 15370
rect 8240 15210 8250 15230
rect 8270 15210 8280 15230
rect 8240 15200 8280 15210
rect 8320 16190 8360 16200
rect 8320 16170 8330 16190
rect 8350 16170 8360 16190
rect 8320 16030 8360 16170
rect 8320 16010 8330 16030
rect 8350 16010 8360 16030
rect 8320 15870 8360 16010
rect 8320 15850 8330 15870
rect 8350 15850 8360 15870
rect 8320 15710 8360 15850
rect 8320 15690 8330 15710
rect 8350 15690 8360 15710
rect 8320 15550 8360 15690
rect 8320 15530 8330 15550
rect 8350 15530 8360 15550
rect 8320 15390 8360 15530
rect 8320 15370 8330 15390
rect 8350 15370 8360 15390
rect 8320 15230 8360 15370
rect 8320 15210 8330 15230
rect 8350 15210 8360 15230
rect 8320 15200 8360 15210
rect 8400 16190 8440 16200
rect 8400 16170 8410 16190
rect 8430 16170 8440 16190
rect 8400 16030 8440 16170
rect 8400 16010 8410 16030
rect 8430 16010 8440 16030
rect 8400 15870 8440 16010
rect 8400 15850 8410 15870
rect 8430 15850 8440 15870
rect 8400 15710 8440 15850
rect 8400 15690 8410 15710
rect 8430 15690 8440 15710
rect 8400 15550 8440 15690
rect 8400 15530 8410 15550
rect 8430 15530 8440 15550
rect 8400 15390 8440 15530
rect 8400 15370 8410 15390
rect 8430 15370 8440 15390
rect 8400 15230 8440 15370
rect 8400 15210 8410 15230
rect 8430 15210 8440 15230
rect 8400 15200 8440 15210
rect 8480 16190 8520 16200
rect 8480 16170 8490 16190
rect 8510 16170 8520 16190
rect 8480 16030 8520 16170
rect 8480 16010 8490 16030
rect 8510 16010 8520 16030
rect 8480 15870 8520 16010
rect 8480 15850 8490 15870
rect 8510 15850 8520 15870
rect 8480 15710 8520 15850
rect 8480 15690 8490 15710
rect 8510 15690 8520 15710
rect 8480 15550 8520 15690
rect 8480 15530 8490 15550
rect 8510 15530 8520 15550
rect 8480 15390 8520 15530
rect 8480 15370 8490 15390
rect 8510 15370 8520 15390
rect 8480 15230 8520 15370
rect 8480 15210 8490 15230
rect 8510 15210 8520 15230
rect 8480 15200 8520 15210
rect 8560 16190 8600 16200
rect 8560 16170 8570 16190
rect 8590 16170 8600 16190
rect 8560 16030 8600 16170
rect 8560 16010 8570 16030
rect 8590 16010 8600 16030
rect 8560 15870 8600 16010
rect 8560 15850 8570 15870
rect 8590 15850 8600 15870
rect 8560 15710 8600 15850
rect 8560 15690 8570 15710
rect 8590 15690 8600 15710
rect 8560 15550 8600 15690
rect 8560 15530 8570 15550
rect 8590 15530 8600 15550
rect 8560 15390 8600 15530
rect 8560 15370 8570 15390
rect 8590 15370 8600 15390
rect 8560 15230 8600 15370
rect 8560 15210 8570 15230
rect 8590 15210 8600 15230
rect 8560 15200 8600 15210
rect 8640 16190 8680 16200
rect 8640 16170 8650 16190
rect 8670 16170 8680 16190
rect 8640 16030 8680 16170
rect 8640 16010 8650 16030
rect 8670 16010 8680 16030
rect 8640 15870 8680 16010
rect 8640 15850 8650 15870
rect 8670 15850 8680 15870
rect 8640 15710 8680 15850
rect 8640 15690 8650 15710
rect 8670 15690 8680 15710
rect 8640 15550 8680 15690
rect 8640 15530 8650 15550
rect 8670 15530 8680 15550
rect 8640 15390 8680 15530
rect 8640 15370 8650 15390
rect 8670 15370 8680 15390
rect 8640 15230 8680 15370
rect 8640 15210 8650 15230
rect 8670 15210 8680 15230
rect 8640 15200 8680 15210
rect 8720 16190 8760 16200
rect 8720 16170 8730 16190
rect 8750 16170 8760 16190
rect 8720 16030 8760 16170
rect 8720 16010 8730 16030
rect 8750 16010 8760 16030
rect 8720 15870 8760 16010
rect 8720 15850 8730 15870
rect 8750 15850 8760 15870
rect 8720 15710 8760 15850
rect 8720 15690 8730 15710
rect 8750 15690 8760 15710
rect 8720 15550 8760 15690
rect 8720 15530 8730 15550
rect 8750 15530 8760 15550
rect 8720 15390 8760 15530
rect 8720 15370 8730 15390
rect 8750 15370 8760 15390
rect 8720 15230 8760 15370
rect 8720 15210 8730 15230
rect 8750 15210 8760 15230
rect 8720 15200 8760 15210
rect 8800 16190 8840 16200
rect 8800 16170 8810 16190
rect 8830 16170 8840 16190
rect 8800 16030 8840 16170
rect 8800 16010 8810 16030
rect 8830 16010 8840 16030
rect 8800 15870 8840 16010
rect 8800 15850 8810 15870
rect 8830 15850 8840 15870
rect 8800 15710 8840 15850
rect 8800 15690 8810 15710
rect 8830 15690 8840 15710
rect 8800 15550 8840 15690
rect 8800 15530 8810 15550
rect 8830 15530 8840 15550
rect 8800 15390 8840 15530
rect 8800 15370 8810 15390
rect 8830 15370 8840 15390
rect 8800 15230 8840 15370
rect 8800 15210 8810 15230
rect 8830 15210 8840 15230
rect 8800 15200 8840 15210
rect 8880 16190 8920 16200
rect 8880 16170 8890 16190
rect 8910 16170 8920 16190
rect 8880 16030 8920 16170
rect 8880 16010 8890 16030
rect 8910 16010 8920 16030
rect 8880 15870 8920 16010
rect 8880 15850 8890 15870
rect 8910 15850 8920 15870
rect 8880 15710 8920 15850
rect 8880 15690 8890 15710
rect 8910 15690 8920 15710
rect 8880 15550 8920 15690
rect 8880 15530 8890 15550
rect 8910 15530 8920 15550
rect 8880 15390 8920 15530
rect 8880 15370 8890 15390
rect 8910 15370 8920 15390
rect 8880 15230 8920 15370
rect 8880 15210 8890 15230
rect 8910 15210 8920 15230
rect 8880 15200 8920 15210
rect 8960 16190 9000 16200
rect 8960 16170 8970 16190
rect 8990 16170 9000 16190
rect 8960 16030 9000 16170
rect 8960 16010 8970 16030
rect 8990 16010 9000 16030
rect 8960 15870 9000 16010
rect 8960 15850 8970 15870
rect 8990 15850 9000 15870
rect 8960 15710 9000 15850
rect 8960 15690 8970 15710
rect 8990 15690 9000 15710
rect 8960 15550 9000 15690
rect 8960 15530 8970 15550
rect 8990 15530 9000 15550
rect 8960 15390 9000 15530
rect 8960 15370 8970 15390
rect 8990 15370 9000 15390
rect 8960 15230 9000 15370
rect 8960 15210 8970 15230
rect 8990 15210 9000 15230
rect 8960 15200 9000 15210
rect 9040 16190 9080 16200
rect 9040 16170 9050 16190
rect 9070 16170 9080 16190
rect 9040 16030 9080 16170
rect 9040 16010 9050 16030
rect 9070 16010 9080 16030
rect 9040 15870 9080 16010
rect 9040 15850 9050 15870
rect 9070 15850 9080 15870
rect 9040 15710 9080 15850
rect 9040 15690 9050 15710
rect 9070 15690 9080 15710
rect 9040 15550 9080 15690
rect 9040 15530 9050 15550
rect 9070 15530 9080 15550
rect 9040 15390 9080 15530
rect 9040 15370 9050 15390
rect 9070 15370 9080 15390
rect 9040 15230 9080 15370
rect 9040 15210 9050 15230
rect 9070 15210 9080 15230
rect 9040 15200 9080 15210
rect 9120 16190 9160 16200
rect 9120 16170 9130 16190
rect 9150 16170 9160 16190
rect 9120 16030 9160 16170
rect 9120 16010 9130 16030
rect 9150 16010 9160 16030
rect 9120 15870 9160 16010
rect 9120 15850 9130 15870
rect 9150 15850 9160 15870
rect 9120 15710 9160 15850
rect 9120 15690 9130 15710
rect 9150 15690 9160 15710
rect 9120 15550 9160 15690
rect 9120 15530 9130 15550
rect 9150 15530 9160 15550
rect 9120 15390 9160 15530
rect 9120 15370 9130 15390
rect 9150 15370 9160 15390
rect 9120 15230 9160 15370
rect 9120 15210 9130 15230
rect 9150 15210 9160 15230
rect 9120 15200 9160 15210
rect 9200 16190 9240 16200
rect 9200 16170 9210 16190
rect 9230 16170 9240 16190
rect 9200 16030 9240 16170
rect 9200 16010 9210 16030
rect 9230 16010 9240 16030
rect 9200 15870 9240 16010
rect 9200 15850 9210 15870
rect 9230 15850 9240 15870
rect 9200 15710 9240 15850
rect 9200 15690 9210 15710
rect 9230 15690 9240 15710
rect 9200 15550 9240 15690
rect 9200 15530 9210 15550
rect 9230 15530 9240 15550
rect 9200 15390 9240 15530
rect 9200 15370 9210 15390
rect 9230 15370 9240 15390
rect 9200 15230 9240 15370
rect 9200 15210 9210 15230
rect 9230 15210 9240 15230
rect 9200 15200 9240 15210
rect 9280 16190 9320 16200
rect 9280 16170 9290 16190
rect 9310 16170 9320 16190
rect 9280 16030 9320 16170
rect 9280 16010 9290 16030
rect 9310 16010 9320 16030
rect 9280 15870 9320 16010
rect 9280 15850 9290 15870
rect 9310 15850 9320 15870
rect 9280 15710 9320 15850
rect 9280 15690 9290 15710
rect 9310 15690 9320 15710
rect 9280 15550 9320 15690
rect 9280 15530 9290 15550
rect 9310 15530 9320 15550
rect 9280 15390 9320 15530
rect 9280 15370 9290 15390
rect 9310 15370 9320 15390
rect 9280 15230 9320 15370
rect 9280 15210 9290 15230
rect 9310 15210 9320 15230
rect 9280 15200 9320 15210
rect 9360 16190 9400 16200
rect 9360 16170 9370 16190
rect 9390 16170 9400 16190
rect 9360 16030 9400 16170
rect 9360 16010 9370 16030
rect 9390 16010 9400 16030
rect 9360 15870 9400 16010
rect 9360 15850 9370 15870
rect 9390 15850 9400 15870
rect 9360 15710 9400 15850
rect 9360 15690 9370 15710
rect 9390 15690 9400 15710
rect 9360 15550 9400 15690
rect 9360 15530 9370 15550
rect 9390 15530 9400 15550
rect 9360 15390 9400 15530
rect 9360 15370 9370 15390
rect 9390 15370 9400 15390
rect 9360 15230 9400 15370
rect 9360 15210 9370 15230
rect 9390 15210 9400 15230
rect 9360 15200 9400 15210
rect 9440 16190 9480 16200
rect 9440 16170 9450 16190
rect 9470 16170 9480 16190
rect 9440 16030 9480 16170
rect 9440 16010 9450 16030
rect 9470 16010 9480 16030
rect 9440 15870 9480 16010
rect 9440 15850 9450 15870
rect 9470 15850 9480 15870
rect 9440 15710 9480 15850
rect 9440 15690 9450 15710
rect 9470 15690 9480 15710
rect 9440 15550 9480 15690
rect 9440 15530 9450 15550
rect 9470 15530 9480 15550
rect 9440 15390 9480 15530
rect 9440 15370 9450 15390
rect 9470 15370 9480 15390
rect 9440 15230 9480 15370
rect 9440 15210 9450 15230
rect 9470 15210 9480 15230
rect 9440 15200 9480 15210
rect 9520 15200 9560 16200
rect 9600 15200 9640 16200
rect 9680 15200 9720 16200
rect 9760 15200 9800 16200
rect 9840 15200 9880 16200
rect 9920 15200 9960 16200
rect 10000 15200 10040 16200
rect 10080 15200 10120 16200
rect 10160 15200 10200 16200
rect 10240 15200 10280 16200
rect 10320 15200 10360 16200
rect 10400 15200 10440 16200
rect 10480 15200 10520 16200
rect 10560 15200 10600 16200
rect 10640 15200 10680 16200
rect 10720 15200 10760 16200
rect 10800 15200 10840 16200
rect 10880 15200 10920 16200
rect 10960 15200 11000 16200
rect 11040 15200 11080 16200
rect 11120 15200 11160 16200
rect 11200 15200 11240 16200
rect 11280 15200 11320 16200
rect 11360 15200 11400 16200
rect 11440 15200 11480 16200
rect 11560 16190 11600 16200
rect 11560 16170 11570 16190
rect 11590 16170 11600 16190
rect 11560 16030 11600 16170
rect 11560 16010 11570 16030
rect 11590 16010 11600 16030
rect 11560 15870 11600 16010
rect 11560 15850 11570 15870
rect 11590 15850 11600 15870
rect 11560 15710 11600 15850
rect 11560 15690 11570 15710
rect 11590 15690 11600 15710
rect 11560 15550 11600 15690
rect 11560 15530 11570 15550
rect 11590 15530 11600 15550
rect 11560 15390 11600 15530
rect 11560 15370 11570 15390
rect 11590 15370 11600 15390
rect 11560 15230 11600 15370
rect 11560 15210 11570 15230
rect 11590 15210 11600 15230
rect 11560 15200 11600 15210
rect 11640 16190 11680 16200
rect 11640 16170 11650 16190
rect 11670 16170 11680 16190
rect 11640 16030 11680 16170
rect 11640 16010 11650 16030
rect 11670 16010 11680 16030
rect 11640 15870 11680 16010
rect 11640 15850 11650 15870
rect 11670 15850 11680 15870
rect 11640 15710 11680 15850
rect 11640 15690 11650 15710
rect 11670 15690 11680 15710
rect 11640 15550 11680 15690
rect 11640 15530 11650 15550
rect 11670 15530 11680 15550
rect 11640 15390 11680 15530
rect 11640 15370 11650 15390
rect 11670 15370 11680 15390
rect 11640 15230 11680 15370
rect 11640 15210 11650 15230
rect 11670 15210 11680 15230
rect 11640 15200 11680 15210
rect 11720 16190 11760 16200
rect 11720 16170 11730 16190
rect 11750 16170 11760 16190
rect 11720 16030 11760 16170
rect 11720 16010 11730 16030
rect 11750 16010 11760 16030
rect 11720 15870 11760 16010
rect 11720 15850 11730 15870
rect 11750 15850 11760 15870
rect 11720 15710 11760 15850
rect 11720 15690 11730 15710
rect 11750 15690 11760 15710
rect 11720 15550 11760 15690
rect 11720 15530 11730 15550
rect 11750 15530 11760 15550
rect 11720 15390 11760 15530
rect 11720 15370 11730 15390
rect 11750 15370 11760 15390
rect 11720 15230 11760 15370
rect 11720 15210 11730 15230
rect 11750 15210 11760 15230
rect 11720 15200 11760 15210
rect 11800 16190 11840 16200
rect 11800 16170 11810 16190
rect 11830 16170 11840 16190
rect 11800 16030 11840 16170
rect 11800 16010 11810 16030
rect 11830 16010 11840 16030
rect 11800 15870 11840 16010
rect 11800 15850 11810 15870
rect 11830 15850 11840 15870
rect 11800 15710 11840 15850
rect 11800 15690 11810 15710
rect 11830 15690 11840 15710
rect 11800 15550 11840 15690
rect 11800 15530 11810 15550
rect 11830 15530 11840 15550
rect 11800 15390 11840 15530
rect 11800 15370 11810 15390
rect 11830 15370 11840 15390
rect 11800 15230 11840 15370
rect 11800 15210 11810 15230
rect 11830 15210 11840 15230
rect 11800 15200 11840 15210
rect 11880 16190 11920 16200
rect 11880 16170 11890 16190
rect 11910 16170 11920 16190
rect 11880 16030 11920 16170
rect 11880 16010 11890 16030
rect 11910 16010 11920 16030
rect 11880 15870 11920 16010
rect 11880 15850 11890 15870
rect 11910 15850 11920 15870
rect 11880 15710 11920 15850
rect 11880 15690 11890 15710
rect 11910 15690 11920 15710
rect 11880 15550 11920 15690
rect 11880 15530 11890 15550
rect 11910 15530 11920 15550
rect 11880 15390 11920 15530
rect 11880 15370 11890 15390
rect 11910 15370 11920 15390
rect 11880 15230 11920 15370
rect 11880 15210 11890 15230
rect 11910 15210 11920 15230
rect 11880 15200 11920 15210
rect 11960 16190 12000 16200
rect 11960 16170 11970 16190
rect 11990 16170 12000 16190
rect 11960 16030 12000 16170
rect 11960 16010 11970 16030
rect 11990 16010 12000 16030
rect 11960 15870 12000 16010
rect 11960 15850 11970 15870
rect 11990 15850 12000 15870
rect 11960 15710 12000 15850
rect 11960 15690 11970 15710
rect 11990 15690 12000 15710
rect 11960 15550 12000 15690
rect 11960 15530 11970 15550
rect 11990 15530 12000 15550
rect 11960 15390 12000 15530
rect 11960 15370 11970 15390
rect 11990 15370 12000 15390
rect 11960 15230 12000 15370
rect 11960 15210 11970 15230
rect 11990 15210 12000 15230
rect 11960 15200 12000 15210
rect 12040 16190 12080 16200
rect 12040 16170 12050 16190
rect 12070 16170 12080 16190
rect 12040 16030 12080 16170
rect 12040 16010 12050 16030
rect 12070 16010 12080 16030
rect 12040 15870 12080 16010
rect 12040 15850 12050 15870
rect 12070 15850 12080 15870
rect 12040 15710 12080 15850
rect 12040 15690 12050 15710
rect 12070 15690 12080 15710
rect 12040 15550 12080 15690
rect 12040 15530 12050 15550
rect 12070 15530 12080 15550
rect 12040 15390 12080 15530
rect 12040 15370 12050 15390
rect 12070 15370 12080 15390
rect 12040 15230 12080 15370
rect 12040 15210 12050 15230
rect 12070 15210 12080 15230
rect 12040 15200 12080 15210
rect 12120 16190 12160 16200
rect 12120 16170 12130 16190
rect 12150 16170 12160 16190
rect 12120 16030 12160 16170
rect 12120 16010 12130 16030
rect 12150 16010 12160 16030
rect 12120 15870 12160 16010
rect 12120 15850 12130 15870
rect 12150 15850 12160 15870
rect 12120 15710 12160 15850
rect 12120 15690 12130 15710
rect 12150 15690 12160 15710
rect 12120 15550 12160 15690
rect 12120 15530 12130 15550
rect 12150 15530 12160 15550
rect 12120 15390 12160 15530
rect 12120 15370 12130 15390
rect 12150 15370 12160 15390
rect 12120 15230 12160 15370
rect 12120 15210 12130 15230
rect 12150 15210 12160 15230
rect 12120 15200 12160 15210
rect 12200 16190 12240 16200
rect 12200 16170 12210 16190
rect 12230 16170 12240 16190
rect 12200 16030 12240 16170
rect 12200 16010 12210 16030
rect 12230 16010 12240 16030
rect 12200 15870 12240 16010
rect 12200 15850 12210 15870
rect 12230 15850 12240 15870
rect 12200 15710 12240 15850
rect 12200 15690 12210 15710
rect 12230 15690 12240 15710
rect 12200 15550 12240 15690
rect 12200 15530 12210 15550
rect 12230 15530 12240 15550
rect 12200 15390 12240 15530
rect 12200 15370 12210 15390
rect 12230 15370 12240 15390
rect 12200 15230 12240 15370
rect 12200 15210 12210 15230
rect 12230 15210 12240 15230
rect 12200 15200 12240 15210
rect 12280 16190 12320 16200
rect 12280 16170 12290 16190
rect 12310 16170 12320 16190
rect 12280 16030 12320 16170
rect 12280 16010 12290 16030
rect 12310 16010 12320 16030
rect 12280 15870 12320 16010
rect 12280 15850 12290 15870
rect 12310 15850 12320 15870
rect 12280 15710 12320 15850
rect 12280 15690 12290 15710
rect 12310 15690 12320 15710
rect 12280 15550 12320 15690
rect 12280 15530 12290 15550
rect 12310 15530 12320 15550
rect 12280 15390 12320 15530
rect 12280 15370 12290 15390
rect 12310 15370 12320 15390
rect 12280 15230 12320 15370
rect 12280 15210 12290 15230
rect 12310 15210 12320 15230
rect 12280 15200 12320 15210
rect 12360 16190 12400 16200
rect 12360 16170 12370 16190
rect 12390 16170 12400 16190
rect 12360 16030 12400 16170
rect 12360 16010 12370 16030
rect 12390 16010 12400 16030
rect 12360 15870 12400 16010
rect 12360 15850 12370 15870
rect 12390 15850 12400 15870
rect 12360 15710 12400 15850
rect 12360 15690 12370 15710
rect 12390 15690 12400 15710
rect 12360 15550 12400 15690
rect 12360 15530 12370 15550
rect 12390 15530 12400 15550
rect 12360 15390 12400 15530
rect 12360 15370 12370 15390
rect 12390 15370 12400 15390
rect 12360 15230 12400 15370
rect 12360 15210 12370 15230
rect 12390 15210 12400 15230
rect 12360 15200 12400 15210
rect 12440 16190 12480 16200
rect 12440 16170 12450 16190
rect 12470 16170 12480 16190
rect 12440 16030 12480 16170
rect 12440 16010 12450 16030
rect 12470 16010 12480 16030
rect 12440 15870 12480 16010
rect 12440 15850 12450 15870
rect 12470 15850 12480 15870
rect 12440 15710 12480 15850
rect 12440 15690 12450 15710
rect 12470 15690 12480 15710
rect 12440 15550 12480 15690
rect 12440 15530 12450 15550
rect 12470 15530 12480 15550
rect 12440 15390 12480 15530
rect 12440 15370 12450 15390
rect 12470 15370 12480 15390
rect 12440 15230 12480 15370
rect 12440 15210 12450 15230
rect 12470 15210 12480 15230
rect 12440 15200 12480 15210
rect 12520 16190 12560 16200
rect 12520 16170 12530 16190
rect 12550 16170 12560 16190
rect 12520 16030 12560 16170
rect 12520 16010 12530 16030
rect 12550 16010 12560 16030
rect 12520 15870 12560 16010
rect 12520 15850 12530 15870
rect 12550 15850 12560 15870
rect 12520 15710 12560 15850
rect 12520 15690 12530 15710
rect 12550 15690 12560 15710
rect 12520 15550 12560 15690
rect 12520 15530 12530 15550
rect 12550 15530 12560 15550
rect 12520 15390 12560 15530
rect 12520 15370 12530 15390
rect 12550 15370 12560 15390
rect 12520 15230 12560 15370
rect 12520 15210 12530 15230
rect 12550 15210 12560 15230
rect 12520 15200 12560 15210
rect 12600 16190 12640 16200
rect 12600 16170 12610 16190
rect 12630 16170 12640 16190
rect 12600 16030 12640 16170
rect 12600 16010 12610 16030
rect 12630 16010 12640 16030
rect 12600 15870 12640 16010
rect 12600 15850 12610 15870
rect 12630 15850 12640 15870
rect 12600 15710 12640 15850
rect 12600 15690 12610 15710
rect 12630 15690 12640 15710
rect 12600 15550 12640 15690
rect 12600 15530 12610 15550
rect 12630 15530 12640 15550
rect 12600 15390 12640 15530
rect 12600 15370 12610 15390
rect 12630 15370 12640 15390
rect 12600 15230 12640 15370
rect 12600 15210 12610 15230
rect 12630 15210 12640 15230
rect 12600 15200 12640 15210
rect 12680 16190 12720 16200
rect 12680 16170 12690 16190
rect 12710 16170 12720 16190
rect 12680 16030 12720 16170
rect 12680 16010 12690 16030
rect 12710 16010 12720 16030
rect 12680 15870 12720 16010
rect 12680 15850 12690 15870
rect 12710 15850 12720 15870
rect 12680 15710 12720 15850
rect 12680 15690 12690 15710
rect 12710 15690 12720 15710
rect 12680 15550 12720 15690
rect 12680 15530 12690 15550
rect 12710 15530 12720 15550
rect 12680 15390 12720 15530
rect 12680 15370 12690 15390
rect 12710 15370 12720 15390
rect 12680 15230 12720 15370
rect 12680 15210 12690 15230
rect 12710 15210 12720 15230
rect 12680 15200 12720 15210
rect 12760 16190 12800 16200
rect 12760 16170 12770 16190
rect 12790 16170 12800 16190
rect 12760 16030 12800 16170
rect 12760 16010 12770 16030
rect 12790 16010 12800 16030
rect 12760 15870 12800 16010
rect 12760 15850 12770 15870
rect 12790 15850 12800 15870
rect 12760 15710 12800 15850
rect 12760 15690 12770 15710
rect 12790 15690 12800 15710
rect 12760 15550 12800 15690
rect 12760 15530 12770 15550
rect 12790 15530 12800 15550
rect 12760 15390 12800 15530
rect 12760 15370 12770 15390
rect 12790 15370 12800 15390
rect 12760 15230 12800 15370
rect 12760 15210 12770 15230
rect 12790 15210 12800 15230
rect 12760 15200 12800 15210
rect 12840 16190 12880 16200
rect 12840 16170 12850 16190
rect 12870 16170 12880 16190
rect 12840 16030 12880 16170
rect 12840 16010 12850 16030
rect 12870 16010 12880 16030
rect 12840 15870 12880 16010
rect 12840 15850 12850 15870
rect 12870 15850 12880 15870
rect 12840 15710 12880 15850
rect 12840 15690 12850 15710
rect 12870 15690 12880 15710
rect 12840 15550 12880 15690
rect 12840 15530 12850 15550
rect 12870 15530 12880 15550
rect 12840 15390 12880 15530
rect 12840 15370 12850 15390
rect 12870 15370 12880 15390
rect 12840 15230 12880 15370
rect 12840 15210 12850 15230
rect 12870 15210 12880 15230
rect 12840 15200 12880 15210
rect 12920 16190 12960 16200
rect 12920 16170 12930 16190
rect 12950 16170 12960 16190
rect 12920 16030 12960 16170
rect 12920 16010 12930 16030
rect 12950 16010 12960 16030
rect 12920 15870 12960 16010
rect 12920 15850 12930 15870
rect 12950 15850 12960 15870
rect 12920 15710 12960 15850
rect 12920 15690 12930 15710
rect 12950 15690 12960 15710
rect 12920 15550 12960 15690
rect 12920 15530 12930 15550
rect 12950 15530 12960 15550
rect 12920 15390 12960 15530
rect 12920 15370 12930 15390
rect 12950 15370 12960 15390
rect 12920 15230 12960 15370
rect 12920 15210 12930 15230
rect 12950 15210 12960 15230
rect 12920 15200 12960 15210
rect 13000 16190 13040 16200
rect 13000 16170 13010 16190
rect 13030 16170 13040 16190
rect 13000 16030 13040 16170
rect 13000 16010 13010 16030
rect 13030 16010 13040 16030
rect 13000 15870 13040 16010
rect 13000 15850 13010 15870
rect 13030 15850 13040 15870
rect 13000 15710 13040 15850
rect 13000 15690 13010 15710
rect 13030 15690 13040 15710
rect 13000 15550 13040 15690
rect 13000 15530 13010 15550
rect 13030 15530 13040 15550
rect 13000 15390 13040 15530
rect 13000 15370 13010 15390
rect 13030 15370 13040 15390
rect 13000 15230 13040 15370
rect 13000 15210 13010 15230
rect 13030 15210 13040 15230
rect 13000 15200 13040 15210
rect 13080 16190 13120 16200
rect 13080 16170 13090 16190
rect 13110 16170 13120 16190
rect 13080 16030 13120 16170
rect 13080 16010 13090 16030
rect 13110 16010 13120 16030
rect 13080 15870 13120 16010
rect 13080 15850 13090 15870
rect 13110 15850 13120 15870
rect 13080 15710 13120 15850
rect 13080 15690 13090 15710
rect 13110 15690 13120 15710
rect 13080 15550 13120 15690
rect 13080 15530 13090 15550
rect 13110 15530 13120 15550
rect 13080 15390 13120 15530
rect 13080 15370 13090 15390
rect 13110 15370 13120 15390
rect 13080 15230 13120 15370
rect 13080 15210 13090 15230
rect 13110 15210 13120 15230
rect 13080 15200 13120 15210
rect 13160 16190 13200 16200
rect 13160 16170 13170 16190
rect 13190 16170 13200 16190
rect 13160 16030 13200 16170
rect 13160 16010 13170 16030
rect 13190 16010 13200 16030
rect 13160 15870 13200 16010
rect 13160 15850 13170 15870
rect 13190 15850 13200 15870
rect 13160 15710 13200 15850
rect 13160 15690 13170 15710
rect 13190 15690 13200 15710
rect 13160 15550 13200 15690
rect 13160 15530 13170 15550
rect 13190 15530 13200 15550
rect 13160 15390 13200 15530
rect 13160 15370 13170 15390
rect 13190 15370 13200 15390
rect 13160 15230 13200 15370
rect 13160 15210 13170 15230
rect 13190 15210 13200 15230
rect 13160 15200 13200 15210
rect 13240 16190 13280 16200
rect 13240 16170 13250 16190
rect 13270 16170 13280 16190
rect 13240 16030 13280 16170
rect 13240 16010 13250 16030
rect 13270 16010 13280 16030
rect 13240 15870 13280 16010
rect 13240 15850 13250 15870
rect 13270 15850 13280 15870
rect 13240 15710 13280 15850
rect 13240 15690 13250 15710
rect 13270 15690 13280 15710
rect 13240 15550 13280 15690
rect 13240 15530 13250 15550
rect 13270 15530 13280 15550
rect 13240 15390 13280 15530
rect 13240 15370 13250 15390
rect 13270 15370 13280 15390
rect 13240 15230 13280 15370
rect 13240 15210 13250 15230
rect 13270 15210 13280 15230
rect 13240 15200 13280 15210
rect 13320 16190 13360 16200
rect 13320 16170 13330 16190
rect 13350 16170 13360 16190
rect 13320 16030 13360 16170
rect 13320 16010 13330 16030
rect 13350 16010 13360 16030
rect 13320 15870 13360 16010
rect 13320 15850 13330 15870
rect 13350 15850 13360 15870
rect 13320 15710 13360 15850
rect 13320 15690 13330 15710
rect 13350 15690 13360 15710
rect 13320 15550 13360 15690
rect 13320 15530 13330 15550
rect 13350 15530 13360 15550
rect 13320 15390 13360 15530
rect 13320 15370 13330 15390
rect 13350 15370 13360 15390
rect 13320 15230 13360 15370
rect 13320 15210 13330 15230
rect 13350 15210 13360 15230
rect 13320 15200 13360 15210
rect 13400 16190 13440 16200
rect 13400 16170 13410 16190
rect 13430 16170 13440 16190
rect 13400 16030 13440 16170
rect 13400 16010 13410 16030
rect 13430 16010 13440 16030
rect 13400 15870 13440 16010
rect 13400 15850 13410 15870
rect 13430 15850 13440 15870
rect 13400 15710 13440 15850
rect 13400 15690 13410 15710
rect 13430 15690 13440 15710
rect 13400 15550 13440 15690
rect 13400 15530 13410 15550
rect 13430 15530 13440 15550
rect 13400 15390 13440 15530
rect 13400 15370 13410 15390
rect 13430 15370 13440 15390
rect 13400 15230 13440 15370
rect 13400 15210 13410 15230
rect 13430 15210 13440 15230
rect 13400 15200 13440 15210
rect 13480 16190 13520 16200
rect 13480 16170 13490 16190
rect 13510 16170 13520 16190
rect 13480 16030 13520 16170
rect 13480 16010 13490 16030
rect 13510 16010 13520 16030
rect 13480 15870 13520 16010
rect 13480 15850 13490 15870
rect 13510 15850 13520 15870
rect 13480 15710 13520 15850
rect 13480 15690 13490 15710
rect 13510 15690 13520 15710
rect 13480 15550 13520 15690
rect 13480 15530 13490 15550
rect 13510 15530 13520 15550
rect 13480 15390 13520 15530
rect 13480 15370 13490 15390
rect 13510 15370 13520 15390
rect 13480 15230 13520 15370
rect 13480 15210 13490 15230
rect 13510 15210 13520 15230
rect 13480 15200 13520 15210
rect 13560 16190 13600 16200
rect 13560 16170 13570 16190
rect 13590 16170 13600 16190
rect 13560 16030 13600 16170
rect 13560 16010 13570 16030
rect 13590 16010 13600 16030
rect 13560 15870 13600 16010
rect 13560 15850 13570 15870
rect 13590 15850 13600 15870
rect 13560 15710 13600 15850
rect 13560 15690 13570 15710
rect 13590 15690 13600 15710
rect 13560 15550 13600 15690
rect 13560 15530 13570 15550
rect 13590 15530 13600 15550
rect 13560 15390 13600 15530
rect 13560 15370 13570 15390
rect 13590 15370 13600 15390
rect 13560 15230 13600 15370
rect 13560 15210 13570 15230
rect 13590 15210 13600 15230
rect 13560 15200 13600 15210
rect 13640 16190 13680 16200
rect 13640 16170 13650 16190
rect 13670 16170 13680 16190
rect 13640 16030 13680 16170
rect 13640 16010 13650 16030
rect 13670 16010 13680 16030
rect 13640 15870 13680 16010
rect 13640 15850 13650 15870
rect 13670 15850 13680 15870
rect 13640 15710 13680 15850
rect 13640 15690 13650 15710
rect 13670 15690 13680 15710
rect 13640 15550 13680 15690
rect 13640 15530 13650 15550
rect 13670 15530 13680 15550
rect 13640 15390 13680 15530
rect 13640 15370 13650 15390
rect 13670 15370 13680 15390
rect 13640 15230 13680 15370
rect 13640 15210 13650 15230
rect 13670 15210 13680 15230
rect 13640 15200 13680 15210
rect 13720 16190 13760 16200
rect 13720 16170 13730 16190
rect 13750 16170 13760 16190
rect 13720 16030 13760 16170
rect 13720 16010 13730 16030
rect 13750 16010 13760 16030
rect 13720 15870 13760 16010
rect 13720 15850 13730 15870
rect 13750 15850 13760 15870
rect 13720 15710 13760 15850
rect 13720 15690 13730 15710
rect 13750 15690 13760 15710
rect 13720 15550 13760 15690
rect 13720 15530 13730 15550
rect 13750 15530 13760 15550
rect 13720 15390 13760 15530
rect 13720 15370 13730 15390
rect 13750 15370 13760 15390
rect 13720 15230 13760 15370
rect 13720 15210 13730 15230
rect 13750 15210 13760 15230
rect 13720 15200 13760 15210
rect 13800 16190 13840 16200
rect 13800 16170 13810 16190
rect 13830 16170 13840 16190
rect 13800 16030 13840 16170
rect 13800 16010 13810 16030
rect 13830 16010 13840 16030
rect 13800 15870 13840 16010
rect 13800 15850 13810 15870
rect 13830 15850 13840 15870
rect 13800 15710 13840 15850
rect 13800 15690 13810 15710
rect 13830 15690 13840 15710
rect 13800 15550 13840 15690
rect 13800 15530 13810 15550
rect 13830 15530 13840 15550
rect 13800 15390 13840 15530
rect 13800 15370 13810 15390
rect 13830 15370 13840 15390
rect 13800 15230 13840 15370
rect 13800 15210 13810 15230
rect 13830 15210 13840 15230
rect 13800 15200 13840 15210
rect 13880 16190 13920 16200
rect 13880 16170 13890 16190
rect 13910 16170 13920 16190
rect 13880 16030 13920 16170
rect 13880 16010 13890 16030
rect 13910 16010 13920 16030
rect 13880 15870 13920 16010
rect 13880 15850 13890 15870
rect 13910 15850 13920 15870
rect 13880 15710 13920 15850
rect 13880 15690 13890 15710
rect 13910 15690 13920 15710
rect 13880 15550 13920 15690
rect 13880 15530 13890 15550
rect 13910 15530 13920 15550
rect 13880 15390 13920 15530
rect 13880 15370 13890 15390
rect 13910 15370 13920 15390
rect 13880 15230 13920 15370
rect 13880 15210 13890 15230
rect 13910 15210 13920 15230
rect 13880 15200 13920 15210
rect 13960 16190 14000 16200
rect 13960 16170 13970 16190
rect 13990 16170 14000 16190
rect 13960 16030 14000 16170
rect 13960 16010 13970 16030
rect 13990 16010 14000 16030
rect 13960 15870 14000 16010
rect 13960 15850 13970 15870
rect 13990 15850 14000 15870
rect 13960 15710 14000 15850
rect 13960 15690 13970 15710
rect 13990 15690 14000 15710
rect 13960 15550 14000 15690
rect 13960 15530 13970 15550
rect 13990 15530 14000 15550
rect 13960 15390 14000 15530
rect 13960 15370 13970 15390
rect 13990 15370 14000 15390
rect 13960 15230 14000 15370
rect 13960 15210 13970 15230
rect 13990 15210 14000 15230
rect 13960 15200 14000 15210
rect 14040 16190 14080 16200
rect 14040 16170 14050 16190
rect 14070 16170 14080 16190
rect 14040 16030 14080 16170
rect 14040 16010 14050 16030
rect 14070 16010 14080 16030
rect 14040 15870 14080 16010
rect 14040 15850 14050 15870
rect 14070 15850 14080 15870
rect 14040 15710 14080 15850
rect 14040 15690 14050 15710
rect 14070 15690 14080 15710
rect 14040 15550 14080 15690
rect 14040 15530 14050 15550
rect 14070 15530 14080 15550
rect 14040 15390 14080 15530
rect 14040 15370 14050 15390
rect 14070 15370 14080 15390
rect 14040 15230 14080 15370
rect 14040 15210 14050 15230
rect 14070 15210 14080 15230
rect 14040 15200 14080 15210
rect 14120 16190 14160 16200
rect 14120 16170 14130 16190
rect 14150 16170 14160 16190
rect 14120 16030 14160 16170
rect 14120 16010 14130 16030
rect 14150 16010 14160 16030
rect 14120 15870 14160 16010
rect 14120 15850 14130 15870
rect 14150 15850 14160 15870
rect 14120 15710 14160 15850
rect 14120 15690 14130 15710
rect 14150 15690 14160 15710
rect 14120 15550 14160 15690
rect 14120 15530 14130 15550
rect 14150 15530 14160 15550
rect 14120 15390 14160 15530
rect 14120 15370 14130 15390
rect 14150 15370 14160 15390
rect 14120 15230 14160 15370
rect 14120 15210 14130 15230
rect 14150 15210 14160 15230
rect 14120 15200 14160 15210
rect 14200 16190 14240 16200
rect 14200 16170 14210 16190
rect 14230 16170 14240 16190
rect 14200 16030 14240 16170
rect 14200 16010 14210 16030
rect 14230 16010 14240 16030
rect 14200 15870 14240 16010
rect 14200 15850 14210 15870
rect 14230 15850 14240 15870
rect 14200 15710 14240 15850
rect 14200 15690 14210 15710
rect 14230 15690 14240 15710
rect 14200 15550 14240 15690
rect 14200 15530 14210 15550
rect 14230 15530 14240 15550
rect 14200 15390 14240 15530
rect 14200 15370 14210 15390
rect 14230 15370 14240 15390
rect 14200 15230 14240 15370
rect 14200 15210 14210 15230
rect 14230 15210 14240 15230
rect 14200 15200 14240 15210
rect 14280 16190 14320 16200
rect 14280 16170 14290 16190
rect 14310 16170 14320 16190
rect 14280 16030 14320 16170
rect 14280 16010 14290 16030
rect 14310 16010 14320 16030
rect 14280 15870 14320 16010
rect 14280 15850 14290 15870
rect 14310 15850 14320 15870
rect 14280 15710 14320 15850
rect 14280 15690 14290 15710
rect 14310 15690 14320 15710
rect 14280 15550 14320 15690
rect 14280 15530 14290 15550
rect 14310 15530 14320 15550
rect 14280 15390 14320 15530
rect 14280 15370 14290 15390
rect 14310 15370 14320 15390
rect 14280 15230 14320 15370
rect 14280 15210 14290 15230
rect 14310 15210 14320 15230
rect 14280 15200 14320 15210
rect 14360 16190 14400 16200
rect 14360 16170 14370 16190
rect 14390 16170 14400 16190
rect 14360 16030 14400 16170
rect 14360 16010 14370 16030
rect 14390 16010 14400 16030
rect 14360 15870 14400 16010
rect 14360 15850 14370 15870
rect 14390 15850 14400 15870
rect 14360 15710 14400 15850
rect 14360 15690 14370 15710
rect 14390 15690 14400 15710
rect 14360 15550 14400 15690
rect 14360 15530 14370 15550
rect 14390 15530 14400 15550
rect 14360 15390 14400 15530
rect 14360 15370 14370 15390
rect 14390 15370 14400 15390
rect 14360 15230 14400 15370
rect 14360 15210 14370 15230
rect 14390 15210 14400 15230
rect 14360 15200 14400 15210
rect 14440 16190 14480 16200
rect 14440 16170 14450 16190
rect 14470 16170 14480 16190
rect 14440 16030 14480 16170
rect 14440 16010 14450 16030
rect 14470 16010 14480 16030
rect 14440 15870 14480 16010
rect 14440 15850 14450 15870
rect 14470 15850 14480 15870
rect 14440 15710 14480 15850
rect 14440 15690 14450 15710
rect 14470 15690 14480 15710
rect 14440 15550 14480 15690
rect 14440 15530 14450 15550
rect 14470 15530 14480 15550
rect 14440 15390 14480 15530
rect 14440 15370 14450 15390
rect 14470 15370 14480 15390
rect 14440 15230 14480 15370
rect 14440 15210 14450 15230
rect 14470 15210 14480 15230
rect 14440 15200 14480 15210
rect 14520 16190 14560 16200
rect 14520 16170 14530 16190
rect 14550 16170 14560 16190
rect 14520 16030 14560 16170
rect 14520 16010 14530 16030
rect 14550 16010 14560 16030
rect 14520 15870 14560 16010
rect 14520 15850 14530 15870
rect 14550 15850 14560 15870
rect 14520 15710 14560 15850
rect 14520 15690 14530 15710
rect 14550 15690 14560 15710
rect 14520 15550 14560 15690
rect 14520 15530 14530 15550
rect 14550 15530 14560 15550
rect 14520 15390 14560 15530
rect 14520 15370 14530 15390
rect 14550 15370 14560 15390
rect 14520 15230 14560 15370
rect 14520 15210 14530 15230
rect 14550 15210 14560 15230
rect 14520 15200 14560 15210
rect 14600 16190 14640 16200
rect 14600 16170 14610 16190
rect 14630 16170 14640 16190
rect 14600 16030 14640 16170
rect 14600 16010 14610 16030
rect 14630 16010 14640 16030
rect 14600 15870 14640 16010
rect 14600 15850 14610 15870
rect 14630 15850 14640 15870
rect 14600 15710 14640 15850
rect 14600 15690 14610 15710
rect 14630 15690 14640 15710
rect 14600 15550 14640 15690
rect 14600 15530 14610 15550
rect 14630 15530 14640 15550
rect 14600 15390 14640 15530
rect 14600 15370 14610 15390
rect 14630 15370 14640 15390
rect 14600 15230 14640 15370
rect 14600 15210 14610 15230
rect 14630 15210 14640 15230
rect 14600 15200 14640 15210
rect 14680 16190 14720 16200
rect 14680 16170 14690 16190
rect 14710 16170 14720 16190
rect 14680 16030 14720 16170
rect 14680 16010 14690 16030
rect 14710 16010 14720 16030
rect 14680 15870 14720 16010
rect 14680 15850 14690 15870
rect 14710 15850 14720 15870
rect 14680 15710 14720 15850
rect 14680 15690 14690 15710
rect 14710 15690 14720 15710
rect 14680 15550 14720 15690
rect 14680 15530 14690 15550
rect 14710 15530 14720 15550
rect 14680 15390 14720 15530
rect 14680 15370 14690 15390
rect 14710 15370 14720 15390
rect 14680 15230 14720 15370
rect 14680 15210 14690 15230
rect 14710 15210 14720 15230
rect 14680 15200 14720 15210
rect 14760 15200 14800 16200
rect 14840 15200 14880 16200
rect 14920 15200 14960 16200
rect 15000 15200 15040 16200
rect 15080 15200 15120 16200
rect 15160 15200 15200 16200
rect 15240 15200 15280 16200
rect 15320 15200 15360 16200
rect 15400 15200 15440 16200
rect 15480 15200 15520 16200
rect 15560 15200 15600 16200
rect 15640 15200 15680 16200
rect 15720 15200 15760 16200
rect 15800 15200 15840 16200
rect 15880 15200 15920 16200
rect 15960 15200 16000 16200
rect 16040 15200 16080 16200
rect 16120 15200 16160 16200
rect 16200 15200 16240 16200
rect 16280 15200 16320 16200
rect 16360 15200 16400 16200
rect 16440 15200 16480 16200
rect 16520 15200 16560 16200
rect 16600 15200 16640 16200
rect 16680 15200 16720 16200
rect 16760 16190 16800 16200
rect 16760 16170 16770 16190
rect 16790 16170 16800 16190
rect 16760 16030 16800 16170
rect 16760 16010 16770 16030
rect 16790 16010 16800 16030
rect 16760 15870 16800 16010
rect 16760 15850 16770 15870
rect 16790 15850 16800 15870
rect 16760 15710 16800 15850
rect 16760 15690 16770 15710
rect 16790 15690 16800 15710
rect 16760 15550 16800 15690
rect 16760 15530 16770 15550
rect 16790 15530 16800 15550
rect 16760 15390 16800 15530
rect 16760 15370 16770 15390
rect 16790 15370 16800 15390
rect 16760 15230 16800 15370
rect 16760 15210 16770 15230
rect 16790 15210 16800 15230
rect 16760 15200 16800 15210
rect 16840 16190 16880 16200
rect 16840 16170 16850 16190
rect 16870 16170 16880 16190
rect 16840 16030 16880 16170
rect 16840 16010 16850 16030
rect 16870 16010 16880 16030
rect 16840 15870 16880 16010
rect 16840 15850 16850 15870
rect 16870 15850 16880 15870
rect 16840 15710 16880 15850
rect 16840 15690 16850 15710
rect 16870 15690 16880 15710
rect 16840 15550 16880 15690
rect 16840 15530 16850 15550
rect 16870 15530 16880 15550
rect 16840 15390 16880 15530
rect 16840 15370 16850 15390
rect 16870 15370 16880 15390
rect 16840 15230 16880 15370
rect 16840 15210 16850 15230
rect 16870 15210 16880 15230
rect 16840 15200 16880 15210
rect 16920 16190 16960 16200
rect 16920 16170 16930 16190
rect 16950 16170 16960 16190
rect 16920 16030 16960 16170
rect 16920 16010 16930 16030
rect 16950 16010 16960 16030
rect 16920 15870 16960 16010
rect 16920 15850 16930 15870
rect 16950 15850 16960 15870
rect 16920 15710 16960 15850
rect 16920 15690 16930 15710
rect 16950 15690 16960 15710
rect 16920 15550 16960 15690
rect 16920 15530 16930 15550
rect 16950 15530 16960 15550
rect 16920 15390 16960 15530
rect 16920 15370 16930 15390
rect 16950 15370 16960 15390
rect 16920 15230 16960 15370
rect 16920 15210 16930 15230
rect 16950 15210 16960 15230
rect 16920 15200 16960 15210
rect 17000 16190 17040 16200
rect 17000 16170 17010 16190
rect 17030 16170 17040 16190
rect 17000 16030 17040 16170
rect 17000 16010 17010 16030
rect 17030 16010 17040 16030
rect 17000 15870 17040 16010
rect 17000 15850 17010 15870
rect 17030 15850 17040 15870
rect 17000 15710 17040 15850
rect 17000 15690 17010 15710
rect 17030 15690 17040 15710
rect 17000 15550 17040 15690
rect 17000 15530 17010 15550
rect 17030 15530 17040 15550
rect 17000 15390 17040 15530
rect 17000 15370 17010 15390
rect 17030 15370 17040 15390
rect 17000 15230 17040 15370
rect 17000 15210 17010 15230
rect 17030 15210 17040 15230
rect 17000 15200 17040 15210
rect 17080 16190 17120 16200
rect 17080 16170 17090 16190
rect 17110 16170 17120 16190
rect 17080 16030 17120 16170
rect 17080 16010 17090 16030
rect 17110 16010 17120 16030
rect 17080 15870 17120 16010
rect 17080 15850 17090 15870
rect 17110 15850 17120 15870
rect 17080 15710 17120 15850
rect 17080 15690 17090 15710
rect 17110 15690 17120 15710
rect 17080 15550 17120 15690
rect 17080 15530 17090 15550
rect 17110 15530 17120 15550
rect 17080 15390 17120 15530
rect 17080 15370 17090 15390
rect 17110 15370 17120 15390
rect 17080 15230 17120 15370
rect 17080 15210 17090 15230
rect 17110 15210 17120 15230
rect 17080 15200 17120 15210
rect 17160 16190 17200 16200
rect 17160 16170 17170 16190
rect 17190 16170 17200 16190
rect 17160 16030 17200 16170
rect 17160 16010 17170 16030
rect 17190 16010 17200 16030
rect 17160 15870 17200 16010
rect 17160 15850 17170 15870
rect 17190 15850 17200 15870
rect 17160 15710 17200 15850
rect 17160 15690 17170 15710
rect 17190 15690 17200 15710
rect 17160 15550 17200 15690
rect 17160 15530 17170 15550
rect 17190 15530 17200 15550
rect 17160 15390 17200 15530
rect 17160 15370 17170 15390
rect 17190 15370 17200 15390
rect 17160 15230 17200 15370
rect 17160 15210 17170 15230
rect 17190 15210 17200 15230
rect 17160 15200 17200 15210
rect 17240 16190 17280 16200
rect 17240 16170 17250 16190
rect 17270 16170 17280 16190
rect 17240 16030 17280 16170
rect 17240 16010 17250 16030
rect 17270 16010 17280 16030
rect 17240 15870 17280 16010
rect 17240 15850 17250 15870
rect 17270 15850 17280 15870
rect 17240 15710 17280 15850
rect 17240 15690 17250 15710
rect 17270 15690 17280 15710
rect 17240 15550 17280 15690
rect 17240 15530 17250 15550
rect 17270 15530 17280 15550
rect 17240 15390 17280 15530
rect 17240 15370 17250 15390
rect 17270 15370 17280 15390
rect 17240 15230 17280 15370
rect 17240 15210 17250 15230
rect 17270 15210 17280 15230
rect 17240 15200 17280 15210
rect 17320 16190 17360 16200
rect 17320 16170 17330 16190
rect 17350 16170 17360 16190
rect 17320 16030 17360 16170
rect 17320 16010 17330 16030
rect 17350 16010 17360 16030
rect 17320 15870 17360 16010
rect 17320 15850 17330 15870
rect 17350 15850 17360 15870
rect 17320 15710 17360 15850
rect 17320 15690 17330 15710
rect 17350 15690 17360 15710
rect 17320 15550 17360 15690
rect 17320 15530 17330 15550
rect 17350 15530 17360 15550
rect 17320 15390 17360 15530
rect 17320 15370 17330 15390
rect 17350 15370 17360 15390
rect 17320 15230 17360 15370
rect 17320 15210 17330 15230
rect 17350 15210 17360 15230
rect 17320 15200 17360 15210
rect 17400 16190 17440 16200
rect 17400 16170 17410 16190
rect 17430 16170 17440 16190
rect 17400 16030 17440 16170
rect 17400 16010 17410 16030
rect 17430 16010 17440 16030
rect 17400 15870 17440 16010
rect 17400 15850 17410 15870
rect 17430 15850 17440 15870
rect 17400 15710 17440 15850
rect 17400 15690 17410 15710
rect 17430 15690 17440 15710
rect 17400 15550 17440 15690
rect 17400 15530 17410 15550
rect 17430 15530 17440 15550
rect 17400 15390 17440 15530
rect 17400 15370 17410 15390
rect 17430 15370 17440 15390
rect 17400 15230 17440 15370
rect 17400 15210 17410 15230
rect 17430 15210 17440 15230
rect 17400 15200 17440 15210
rect 17480 16190 17520 16200
rect 17480 16170 17490 16190
rect 17510 16170 17520 16190
rect 17480 16030 17520 16170
rect 17480 16010 17490 16030
rect 17510 16010 17520 16030
rect 17480 15870 17520 16010
rect 17480 15850 17490 15870
rect 17510 15850 17520 15870
rect 17480 15710 17520 15850
rect 17480 15690 17490 15710
rect 17510 15690 17520 15710
rect 17480 15550 17520 15690
rect 17480 15530 17490 15550
rect 17510 15530 17520 15550
rect 17480 15390 17520 15530
rect 17480 15370 17490 15390
rect 17510 15370 17520 15390
rect 17480 15230 17520 15370
rect 17480 15210 17490 15230
rect 17510 15210 17520 15230
rect 17480 15200 17520 15210
rect 17560 16190 17600 16200
rect 17560 16170 17570 16190
rect 17590 16170 17600 16190
rect 17560 16030 17600 16170
rect 17560 16010 17570 16030
rect 17590 16010 17600 16030
rect 17560 15870 17600 16010
rect 17560 15850 17570 15870
rect 17590 15850 17600 15870
rect 17560 15710 17600 15850
rect 17560 15690 17570 15710
rect 17590 15690 17600 15710
rect 17560 15550 17600 15690
rect 17560 15530 17570 15550
rect 17590 15530 17600 15550
rect 17560 15390 17600 15530
rect 17560 15370 17570 15390
rect 17590 15370 17600 15390
rect 17560 15230 17600 15370
rect 17560 15210 17570 15230
rect 17590 15210 17600 15230
rect 17560 15200 17600 15210
rect 17640 16190 17680 16200
rect 17640 16170 17650 16190
rect 17670 16170 17680 16190
rect 17640 16030 17680 16170
rect 17640 16010 17650 16030
rect 17670 16010 17680 16030
rect 17640 15870 17680 16010
rect 17640 15850 17650 15870
rect 17670 15850 17680 15870
rect 17640 15710 17680 15850
rect 17640 15690 17650 15710
rect 17670 15690 17680 15710
rect 17640 15550 17680 15690
rect 17640 15530 17650 15550
rect 17670 15530 17680 15550
rect 17640 15390 17680 15530
rect 17640 15370 17650 15390
rect 17670 15370 17680 15390
rect 17640 15230 17680 15370
rect 17640 15210 17650 15230
rect 17670 15210 17680 15230
rect 17640 15200 17680 15210
rect 17720 16190 17760 16200
rect 17720 16170 17730 16190
rect 17750 16170 17760 16190
rect 17720 16030 17760 16170
rect 17720 16010 17730 16030
rect 17750 16010 17760 16030
rect 17720 15870 17760 16010
rect 17720 15850 17730 15870
rect 17750 15850 17760 15870
rect 17720 15710 17760 15850
rect 17720 15690 17730 15710
rect 17750 15690 17760 15710
rect 17720 15550 17760 15690
rect 17720 15530 17730 15550
rect 17750 15530 17760 15550
rect 17720 15390 17760 15530
rect 17720 15370 17730 15390
rect 17750 15370 17760 15390
rect 17720 15230 17760 15370
rect 17720 15210 17730 15230
rect 17750 15210 17760 15230
rect 17720 15200 17760 15210
rect 17800 16190 17840 16200
rect 17800 16170 17810 16190
rect 17830 16170 17840 16190
rect 17800 16030 17840 16170
rect 17800 16010 17810 16030
rect 17830 16010 17840 16030
rect 17800 15870 17840 16010
rect 17800 15850 17810 15870
rect 17830 15850 17840 15870
rect 17800 15710 17840 15850
rect 17800 15690 17810 15710
rect 17830 15690 17840 15710
rect 17800 15550 17840 15690
rect 17800 15530 17810 15550
rect 17830 15530 17840 15550
rect 17800 15390 17840 15530
rect 17800 15370 17810 15390
rect 17830 15370 17840 15390
rect 17800 15230 17840 15370
rect 17800 15210 17810 15230
rect 17830 15210 17840 15230
rect 17800 15200 17840 15210
rect 17880 16190 17920 16200
rect 17880 16170 17890 16190
rect 17910 16170 17920 16190
rect 17880 16030 17920 16170
rect 17880 16010 17890 16030
rect 17910 16010 17920 16030
rect 17880 15870 17920 16010
rect 17880 15850 17890 15870
rect 17910 15850 17920 15870
rect 17880 15710 17920 15850
rect 17880 15690 17890 15710
rect 17910 15690 17920 15710
rect 17880 15550 17920 15690
rect 17880 15530 17890 15550
rect 17910 15530 17920 15550
rect 17880 15390 17920 15530
rect 17880 15370 17890 15390
rect 17910 15370 17920 15390
rect 17880 15230 17920 15370
rect 17880 15210 17890 15230
rect 17910 15210 17920 15230
rect 17880 15200 17920 15210
rect 17960 16190 18000 16200
rect 17960 16170 17970 16190
rect 17990 16170 18000 16190
rect 17960 16030 18000 16170
rect 17960 16010 17970 16030
rect 17990 16010 18000 16030
rect 17960 15870 18000 16010
rect 17960 15850 17970 15870
rect 17990 15850 18000 15870
rect 17960 15710 18000 15850
rect 17960 15690 17970 15710
rect 17990 15690 18000 15710
rect 17960 15550 18000 15690
rect 17960 15530 17970 15550
rect 17990 15530 18000 15550
rect 17960 15390 18000 15530
rect 17960 15370 17970 15390
rect 17990 15370 18000 15390
rect 17960 15230 18000 15370
rect 17960 15210 17970 15230
rect 17990 15210 18000 15230
rect 17960 15200 18000 15210
rect 18040 16190 18080 16200
rect 18040 16170 18050 16190
rect 18070 16170 18080 16190
rect 18040 16030 18080 16170
rect 18040 16010 18050 16030
rect 18070 16010 18080 16030
rect 18040 15870 18080 16010
rect 18040 15850 18050 15870
rect 18070 15850 18080 15870
rect 18040 15710 18080 15850
rect 18040 15690 18050 15710
rect 18070 15690 18080 15710
rect 18040 15550 18080 15690
rect 18040 15530 18050 15550
rect 18070 15530 18080 15550
rect 18040 15390 18080 15530
rect 18040 15370 18050 15390
rect 18070 15370 18080 15390
rect 18040 15230 18080 15370
rect 18040 15210 18050 15230
rect 18070 15210 18080 15230
rect 18040 15200 18080 15210
rect 18120 16190 18160 16200
rect 18120 16170 18130 16190
rect 18150 16170 18160 16190
rect 18120 16030 18160 16170
rect 18120 16010 18130 16030
rect 18150 16010 18160 16030
rect 18120 15870 18160 16010
rect 18120 15850 18130 15870
rect 18150 15850 18160 15870
rect 18120 15710 18160 15850
rect 18120 15690 18130 15710
rect 18150 15690 18160 15710
rect 18120 15550 18160 15690
rect 18120 15530 18130 15550
rect 18150 15530 18160 15550
rect 18120 15390 18160 15530
rect 18120 15370 18130 15390
rect 18150 15370 18160 15390
rect 18120 15230 18160 15370
rect 18120 15210 18130 15230
rect 18150 15210 18160 15230
rect 18120 15200 18160 15210
rect 18200 16190 18240 16200
rect 18200 16170 18210 16190
rect 18230 16170 18240 16190
rect 18200 16030 18240 16170
rect 18200 16010 18210 16030
rect 18230 16010 18240 16030
rect 18200 15870 18240 16010
rect 18200 15850 18210 15870
rect 18230 15850 18240 15870
rect 18200 15710 18240 15850
rect 18200 15690 18210 15710
rect 18230 15690 18240 15710
rect 18200 15550 18240 15690
rect 18200 15530 18210 15550
rect 18230 15530 18240 15550
rect 18200 15390 18240 15530
rect 18200 15370 18210 15390
rect 18230 15370 18240 15390
rect 18200 15230 18240 15370
rect 18200 15210 18210 15230
rect 18230 15210 18240 15230
rect 18200 15200 18240 15210
rect 18280 16190 18320 16200
rect 18280 16170 18290 16190
rect 18310 16170 18320 16190
rect 18280 16030 18320 16170
rect 18280 16010 18290 16030
rect 18310 16010 18320 16030
rect 18280 15870 18320 16010
rect 18280 15850 18290 15870
rect 18310 15850 18320 15870
rect 18280 15710 18320 15850
rect 18280 15690 18290 15710
rect 18310 15690 18320 15710
rect 18280 15550 18320 15690
rect 18280 15530 18290 15550
rect 18310 15530 18320 15550
rect 18280 15390 18320 15530
rect 18280 15370 18290 15390
rect 18310 15370 18320 15390
rect 18280 15230 18320 15370
rect 18280 15210 18290 15230
rect 18310 15210 18320 15230
rect 18280 15200 18320 15210
rect 18360 16190 18400 16200
rect 18360 16170 18370 16190
rect 18390 16170 18400 16190
rect 18360 16030 18400 16170
rect 18360 16010 18370 16030
rect 18390 16010 18400 16030
rect 18360 15870 18400 16010
rect 18360 15850 18370 15870
rect 18390 15850 18400 15870
rect 18360 15710 18400 15850
rect 18360 15690 18370 15710
rect 18390 15690 18400 15710
rect 18360 15550 18400 15690
rect 18360 15530 18370 15550
rect 18390 15530 18400 15550
rect 18360 15390 18400 15530
rect 18360 15370 18370 15390
rect 18390 15370 18400 15390
rect 18360 15230 18400 15370
rect 18360 15210 18370 15230
rect 18390 15210 18400 15230
rect 18360 15200 18400 15210
rect 18440 16190 18480 16200
rect 18440 16170 18450 16190
rect 18470 16170 18480 16190
rect 18440 16030 18480 16170
rect 18440 16010 18450 16030
rect 18470 16010 18480 16030
rect 18440 15870 18480 16010
rect 18440 15850 18450 15870
rect 18470 15850 18480 15870
rect 18440 15710 18480 15850
rect 18440 15690 18450 15710
rect 18470 15690 18480 15710
rect 18440 15550 18480 15690
rect 18440 15530 18450 15550
rect 18470 15530 18480 15550
rect 18440 15390 18480 15530
rect 18440 15370 18450 15390
rect 18470 15370 18480 15390
rect 18440 15230 18480 15370
rect 18440 15210 18450 15230
rect 18470 15210 18480 15230
rect 18440 15200 18480 15210
rect 18520 16190 18560 16200
rect 18520 16170 18530 16190
rect 18550 16170 18560 16190
rect 18520 16030 18560 16170
rect 18520 16010 18530 16030
rect 18550 16010 18560 16030
rect 18520 15870 18560 16010
rect 18520 15850 18530 15870
rect 18550 15850 18560 15870
rect 18520 15710 18560 15850
rect 18520 15690 18530 15710
rect 18550 15690 18560 15710
rect 18520 15550 18560 15690
rect 18520 15530 18530 15550
rect 18550 15530 18560 15550
rect 18520 15390 18560 15530
rect 18520 15370 18530 15390
rect 18550 15370 18560 15390
rect 18520 15230 18560 15370
rect 18520 15210 18530 15230
rect 18550 15210 18560 15230
rect 18520 15200 18560 15210
rect 18600 16190 18640 16200
rect 18600 16170 18610 16190
rect 18630 16170 18640 16190
rect 18600 16030 18640 16170
rect 18600 16010 18610 16030
rect 18630 16010 18640 16030
rect 18600 15870 18640 16010
rect 18600 15850 18610 15870
rect 18630 15850 18640 15870
rect 18600 15710 18640 15850
rect 18600 15690 18610 15710
rect 18630 15690 18640 15710
rect 18600 15550 18640 15690
rect 18600 15530 18610 15550
rect 18630 15530 18640 15550
rect 18600 15390 18640 15530
rect 18600 15370 18610 15390
rect 18630 15370 18640 15390
rect 18600 15230 18640 15370
rect 18600 15210 18610 15230
rect 18630 15210 18640 15230
rect 18600 15200 18640 15210
rect 18680 16190 18720 16200
rect 18680 16170 18690 16190
rect 18710 16170 18720 16190
rect 18680 16030 18720 16170
rect 18680 16010 18690 16030
rect 18710 16010 18720 16030
rect 18680 15870 18720 16010
rect 18680 15850 18690 15870
rect 18710 15850 18720 15870
rect 18680 15710 18720 15850
rect 18680 15690 18690 15710
rect 18710 15690 18720 15710
rect 18680 15550 18720 15690
rect 18680 15530 18690 15550
rect 18710 15530 18720 15550
rect 18680 15390 18720 15530
rect 18680 15370 18690 15390
rect 18710 15370 18720 15390
rect 18680 15230 18720 15370
rect 18680 15210 18690 15230
rect 18710 15210 18720 15230
rect 18680 15200 18720 15210
rect 18760 16190 18800 16200
rect 18760 16170 18770 16190
rect 18790 16170 18800 16190
rect 18760 16030 18800 16170
rect 18760 16010 18770 16030
rect 18790 16010 18800 16030
rect 18760 15870 18800 16010
rect 18760 15850 18770 15870
rect 18790 15850 18800 15870
rect 18760 15710 18800 15850
rect 18760 15690 18770 15710
rect 18790 15690 18800 15710
rect 18760 15550 18800 15690
rect 18760 15530 18770 15550
rect 18790 15530 18800 15550
rect 18760 15390 18800 15530
rect 18760 15370 18770 15390
rect 18790 15370 18800 15390
rect 18760 15230 18800 15370
rect 18760 15210 18770 15230
rect 18790 15210 18800 15230
rect 18760 15200 18800 15210
rect 18840 16190 18880 16200
rect 18840 16170 18850 16190
rect 18870 16170 18880 16190
rect 18840 16030 18880 16170
rect 18840 16010 18850 16030
rect 18870 16010 18880 16030
rect 18840 15870 18880 16010
rect 18840 15850 18850 15870
rect 18870 15850 18880 15870
rect 18840 15710 18880 15850
rect 18840 15690 18850 15710
rect 18870 15690 18880 15710
rect 18840 15550 18880 15690
rect 18840 15530 18850 15550
rect 18870 15530 18880 15550
rect 18840 15390 18880 15530
rect 18840 15370 18850 15390
rect 18870 15370 18880 15390
rect 18840 15230 18880 15370
rect 18840 15210 18850 15230
rect 18870 15210 18880 15230
rect 18840 15200 18880 15210
rect 18920 16190 18960 16200
rect 18920 16170 18930 16190
rect 18950 16170 18960 16190
rect 18920 16030 18960 16170
rect 18920 16010 18930 16030
rect 18950 16010 18960 16030
rect 18920 15870 18960 16010
rect 18920 15850 18930 15870
rect 18950 15850 18960 15870
rect 18920 15710 18960 15850
rect 18920 15690 18930 15710
rect 18950 15690 18960 15710
rect 18920 15550 18960 15690
rect 18920 15530 18930 15550
rect 18950 15530 18960 15550
rect 18920 15390 18960 15530
rect 18920 15370 18930 15390
rect 18950 15370 18960 15390
rect 18920 15230 18960 15370
rect 18920 15210 18930 15230
rect 18950 15210 18960 15230
rect 18920 15200 18960 15210
rect 19000 16190 19040 16200
rect 19000 16170 19010 16190
rect 19030 16170 19040 16190
rect 19000 16030 19040 16170
rect 19000 16010 19010 16030
rect 19030 16010 19040 16030
rect 19000 15870 19040 16010
rect 19000 15850 19010 15870
rect 19030 15850 19040 15870
rect 19000 15710 19040 15850
rect 19000 15690 19010 15710
rect 19030 15690 19040 15710
rect 19000 15550 19040 15690
rect 19000 15530 19010 15550
rect 19030 15530 19040 15550
rect 19000 15390 19040 15530
rect 19000 15370 19010 15390
rect 19030 15370 19040 15390
rect 19000 15230 19040 15370
rect 19000 15210 19010 15230
rect 19030 15210 19040 15230
rect 19000 15200 19040 15210
rect 19080 16190 19120 16200
rect 19080 16170 19090 16190
rect 19110 16170 19120 16190
rect 19080 16030 19120 16170
rect 19080 16010 19090 16030
rect 19110 16010 19120 16030
rect 19080 15870 19120 16010
rect 19080 15850 19090 15870
rect 19110 15850 19120 15870
rect 19080 15710 19120 15850
rect 19080 15690 19090 15710
rect 19110 15690 19120 15710
rect 19080 15550 19120 15690
rect 19080 15530 19090 15550
rect 19110 15530 19120 15550
rect 19080 15390 19120 15530
rect 19080 15370 19090 15390
rect 19110 15370 19120 15390
rect 19080 15230 19120 15370
rect 19080 15210 19090 15230
rect 19110 15210 19120 15230
rect 19080 15200 19120 15210
rect 19160 16190 19200 16200
rect 19160 16170 19170 16190
rect 19190 16170 19200 16190
rect 19160 16030 19200 16170
rect 19160 16010 19170 16030
rect 19190 16010 19200 16030
rect 19160 15870 19200 16010
rect 19160 15850 19170 15870
rect 19190 15850 19200 15870
rect 19160 15710 19200 15850
rect 19160 15690 19170 15710
rect 19190 15690 19200 15710
rect 19160 15550 19200 15690
rect 19160 15530 19170 15550
rect 19190 15530 19200 15550
rect 19160 15390 19200 15530
rect 19160 15370 19170 15390
rect 19190 15370 19200 15390
rect 19160 15230 19200 15370
rect 19160 15210 19170 15230
rect 19190 15210 19200 15230
rect 19160 15200 19200 15210
rect 19240 16190 19280 16200
rect 19240 16170 19250 16190
rect 19270 16170 19280 16190
rect 19240 16030 19280 16170
rect 19240 16010 19250 16030
rect 19270 16010 19280 16030
rect 19240 15870 19280 16010
rect 19240 15850 19250 15870
rect 19270 15850 19280 15870
rect 19240 15710 19280 15850
rect 19240 15690 19250 15710
rect 19270 15690 19280 15710
rect 19240 15550 19280 15690
rect 19240 15530 19250 15550
rect 19270 15530 19280 15550
rect 19240 15390 19280 15530
rect 19240 15370 19250 15390
rect 19270 15370 19280 15390
rect 19240 15230 19280 15370
rect 19240 15210 19250 15230
rect 19270 15210 19280 15230
rect 19240 15200 19280 15210
rect 19320 16190 19360 16200
rect 19320 16170 19330 16190
rect 19350 16170 19360 16190
rect 19320 16030 19360 16170
rect 19320 16010 19330 16030
rect 19350 16010 19360 16030
rect 19320 15870 19360 16010
rect 19320 15850 19330 15870
rect 19350 15850 19360 15870
rect 19320 15710 19360 15850
rect 19320 15690 19330 15710
rect 19350 15690 19360 15710
rect 19320 15550 19360 15690
rect 19320 15530 19330 15550
rect 19350 15530 19360 15550
rect 19320 15390 19360 15530
rect 19320 15370 19330 15390
rect 19350 15370 19360 15390
rect 19320 15230 19360 15370
rect 19320 15210 19330 15230
rect 19350 15210 19360 15230
rect 19320 15200 19360 15210
rect 19400 16190 19440 16200
rect 19400 16170 19410 16190
rect 19430 16170 19440 16190
rect 19400 16030 19440 16170
rect 19400 16010 19410 16030
rect 19430 16010 19440 16030
rect 19400 15870 19440 16010
rect 19400 15850 19410 15870
rect 19430 15850 19440 15870
rect 19400 15710 19440 15850
rect 19400 15690 19410 15710
rect 19430 15690 19440 15710
rect 19400 15550 19440 15690
rect 19400 15530 19410 15550
rect 19430 15530 19440 15550
rect 19400 15390 19440 15530
rect 19400 15370 19410 15390
rect 19430 15370 19440 15390
rect 19400 15230 19440 15370
rect 19400 15210 19410 15230
rect 19430 15210 19440 15230
rect 19400 15200 19440 15210
rect 19480 16190 19520 16200
rect 19480 16170 19490 16190
rect 19510 16170 19520 16190
rect 19480 16030 19520 16170
rect 19480 16010 19490 16030
rect 19510 16010 19520 16030
rect 19480 15870 19520 16010
rect 19480 15850 19490 15870
rect 19510 15850 19520 15870
rect 19480 15710 19520 15850
rect 19480 15690 19490 15710
rect 19510 15690 19520 15710
rect 19480 15550 19520 15690
rect 19480 15530 19490 15550
rect 19510 15530 19520 15550
rect 19480 15390 19520 15530
rect 19480 15370 19490 15390
rect 19510 15370 19520 15390
rect 19480 15230 19520 15370
rect 19480 15210 19490 15230
rect 19510 15210 19520 15230
rect 19480 15200 19520 15210
rect 19560 16190 19600 16200
rect 19560 16170 19570 16190
rect 19590 16170 19600 16190
rect 19560 16030 19600 16170
rect 19560 16010 19570 16030
rect 19590 16010 19600 16030
rect 19560 15870 19600 16010
rect 19560 15850 19570 15870
rect 19590 15850 19600 15870
rect 19560 15710 19600 15850
rect 19560 15690 19570 15710
rect 19590 15690 19600 15710
rect 19560 15550 19600 15690
rect 19560 15530 19570 15550
rect 19590 15530 19600 15550
rect 19560 15390 19600 15530
rect 19560 15370 19570 15390
rect 19590 15370 19600 15390
rect 19560 15230 19600 15370
rect 19560 15210 19570 15230
rect 19590 15210 19600 15230
rect 19560 15200 19600 15210
rect 19640 16190 19680 16200
rect 19640 16170 19650 16190
rect 19670 16170 19680 16190
rect 19640 16030 19680 16170
rect 19640 16010 19650 16030
rect 19670 16010 19680 16030
rect 19640 15870 19680 16010
rect 19640 15850 19650 15870
rect 19670 15850 19680 15870
rect 19640 15710 19680 15850
rect 19640 15690 19650 15710
rect 19670 15690 19680 15710
rect 19640 15550 19680 15690
rect 19640 15530 19650 15550
rect 19670 15530 19680 15550
rect 19640 15390 19680 15530
rect 19640 15370 19650 15390
rect 19670 15370 19680 15390
rect 19640 15230 19680 15370
rect 19640 15210 19650 15230
rect 19670 15210 19680 15230
rect 19640 15200 19680 15210
rect 19720 16190 19760 16200
rect 19720 16170 19730 16190
rect 19750 16170 19760 16190
rect 19720 16030 19760 16170
rect 19720 16010 19730 16030
rect 19750 16010 19760 16030
rect 19720 15870 19760 16010
rect 19720 15850 19730 15870
rect 19750 15850 19760 15870
rect 19720 15710 19760 15850
rect 19720 15690 19730 15710
rect 19750 15690 19760 15710
rect 19720 15550 19760 15690
rect 19720 15530 19730 15550
rect 19750 15530 19760 15550
rect 19720 15390 19760 15530
rect 19720 15370 19730 15390
rect 19750 15370 19760 15390
rect 19720 15230 19760 15370
rect 19720 15210 19730 15230
rect 19750 15210 19760 15230
rect 19720 15200 19760 15210
rect 19800 16190 19840 16200
rect 19800 16170 19810 16190
rect 19830 16170 19840 16190
rect 19800 16030 19840 16170
rect 19800 16010 19810 16030
rect 19830 16010 19840 16030
rect 19800 15870 19840 16010
rect 19800 15850 19810 15870
rect 19830 15850 19840 15870
rect 19800 15710 19840 15850
rect 19800 15690 19810 15710
rect 19830 15690 19840 15710
rect 19800 15550 19840 15690
rect 19800 15530 19810 15550
rect 19830 15530 19840 15550
rect 19800 15390 19840 15530
rect 19800 15370 19810 15390
rect 19830 15370 19840 15390
rect 19800 15230 19840 15370
rect 19800 15210 19810 15230
rect 19830 15210 19840 15230
rect 19800 15200 19840 15210
rect 19880 16190 19920 16200
rect 19880 16170 19890 16190
rect 19910 16170 19920 16190
rect 19880 16030 19920 16170
rect 19880 16010 19890 16030
rect 19910 16010 19920 16030
rect 19880 15870 19920 16010
rect 19880 15850 19890 15870
rect 19910 15850 19920 15870
rect 19880 15710 19920 15850
rect 19880 15690 19890 15710
rect 19910 15690 19920 15710
rect 19880 15550 19920 15690
rect 19880 15530 19890 15550
rect 19910 15530 19920 15550
rect 19880 15390 19920 15530
rect 19880 15370 19890 15390
rect 19910 15370 19920 15390
rect 19880 15230 19920 15370
rect 19880 15210 19890 15230
rect 19910 15210 19920 15230
rect 19880 15200 19920 15210
rect 19960 16190 20000 16200
rect 19960 16170 19970 16190
rect 19990 16170 20000 16190
rect 19960 16030 20000 16170
rect 19960 16010 19970 16030
rect 19990 16010 20000 16030
rect 19960 15870 20000 16010
rect 19960 15850 19970 15870
rect 19990 15850 20000 15870
rect 19960 15710 20000 15850
rect 19960 15690 19970 15710
rect 19990 15690 20000 15710
rect 19960 15550 20000 15690
rect 19960 15530 19970 15550
rect 19990 15530 20000 15550
rect 19960 15390 20000 15530
rect 19960 15370 19970 15390
rect 19990 15370 20000 15390
rect 19960 15230 20000 15370
rect 19960 15210 19970 15230
rect 19990 15210 20000 15230
rect 19960 15200 20000 15210
rect 20040 16190 20080 16200
rect 20040 16170 20050 16190
rect 20070 16170 20080 16190
rect 20040 16030 20080 16170
rect 20040 16010 20050 16030
rect 20070 16010 20080 16030
rect 20040 15870 20080 16010
rect 20040 15850 20050 15870
rect 20070 15850 20080 15870
rect 20040 15710 20080 15850
rect 20040 15690 20050 15710
rect 20070 15690 20080 15710
rect 20040 15550 20080 15690
rect 20040 15530 20050 15550
rect 20070 15530 20080 15550
rect 20040 15390 20080 15530
rect 20040 15370 20050 15390
rect 20070 15370 20080 15390
rect 20040 15230 20080 15370
rect 20040 15210 20050 15230
rect 20070 15210 20080 15230
rect 20040 15200 20080 15210
rect 20120 16190 20160 16200
rect 20120 16170 20130 16190
rect 20150 16170 20160 16190
rect 20120 16030 20160 16170
rect 20120 16010 20130 16030
rect 20150 16010 20160 16030
rect 20120 15870 20160 16010
rect 20120 15850 20130 15870
rect 20150 15850 20160 15870
rect 20120 15710 20160 15850
rect 20120 15690 20130 15710
rect 20150 15690 20160 15710
rect 20120 15550 20160 15690
rect 20120 15530 20130 15550
rect 20150 15530 20160 15550
rect 20120 15390 20160 15530
rect 20120 15370 20130 15390
rect 20150 15370 20160 15390
rect 20120 15230 20160 15370
rect 20120 15210 20130 15230
rect 20150 15210 20160 15230
rect 20120 15200 20160 15210
rect 20200 16190 20240 16200
rect 20200 16170 20210 16190
rect 20230 16170 20240 16190
rect 20200 16030 20240 16170
rect 20200 16010 20210 16030
rect 20230 16010 20240 16030
rect 20200 15870 20240 16010
rect 20200 15850 20210 15870
rect 20230 15850 20240 15870
rect 20200 15710 20240 15850
rect 20200 15690 20210 15710
rect 20230 15690 20240 15710
rect 20200 15550 20240 15690
rect 20200 15530 20210 15550
rect 20230 15530 20240 15550
rect 20200 15390 20240 15530
rect 20200 15370 20210 15390
rect 20230 15370 20240 15390
rect 20200 15230 20240 15370
rect 20200 15210 20210 15230
rect 20230 15210 20240 15230
rect 20200 15200 20240 15210
rect 20280 16190 20320 16200
rect 20280 16170 20290 16190
rect 20310 16170 20320 16190
rect 20280 16030 20320 16170
rect 20280 16010 20290 16030
rect 20310 16010 20320 16030
rect 20280 15870 20320 16010
rect 20280 15850 20290 15870
rect 20310 15850 20320 15870
rect 20280 15710 20320 15850
rect 20280 15690 20290 15710
rect 20310 15690 20320 15710
rect 20280 15550 20320 15690
rect 20280 15530 20290 15550
rect 20310 15530 20320 15550
rect 20280 15390 20320 15530
rect 20280 15370 20290 15390
rect 20310 15370 20320 15390
rect 20280 15230 20320 15370
rect 20280 15210 20290 15230
rect 20310 15210 20320 15230
rect 20280 15200 20320 15210
rect 20360 16190 20400 16200
rect 20360 16170 20370 16190
rect 20390 16170 20400 16190
rect 20360 16030 20400 16170
rect 20360 16010 20370 16030
rect 20390 16010 20400 16030
rect 20360 15870 20400 16010
rect 20360 15850 20370 15870
rect 20390 15850 20400 15870
rect 20360 15710 20400 15850
rect 20360 15690 20370 15710
rect 20390 15690 20400 15710
rect 20360 15550 20400 15690
rect 20360 15530 20370 15550
rect 20390 15530 20400 15550
rect 20360 15390 20400 15530
rect 20360 15370 20370 15390
rect 20390 15370 20400 15390
rect 20360 15230 20400 15370
rect 20360 15210 20370 15230
rect 20390 15210 20400 15230
rect 20360 15200 20400 15210
rect 20440 16190 20480 16200
rect 20440 16170 20450 16190
rect 20470 16170 20480 16190
rect 20440 16030 20480 16170
rect 20440 16010 20450 16030
rect 20470 16010 20480 16030
rect 20440 15870 20480 16010
rect 20440 15850 20450 15870
rect 20470 15850 20480 15870
rect 20440 15710 20480 15850
rect 20440 15690 20450 15710
rect 20470 15690 20480 15710
rect 20440 15550 20480 15690
rect 20440 15530 20450 15550
rect 20470 15530 20480 15550
rect 20440 15390 20480 15530
rect 20440 15370 20450 15390
rect 20470 15370 20480 15390
rect 20440 15230 20480 15370
rect 20440 15210 20450 15230
rect 20470 15210 20480 15230
rect 20440 15200 20480 15210
rect 20520 16190 20560 16200
rect 20520 16170 20530 16190
rect 20550 16170 20560 16190
rect 20520 16030 20560 16170
rect 20520 16010 20530 16030
rect 20550 16010 20560 16030
rect 20520 15870 20560 16010
rect 20520 15850 20530 15870
rect 20550 15850 20560 15870
rect 20520 15710 20560 15850
rect 20520 15690 20530 15710
rect 20550 15690 20560 15710
rect 20520 15550 20560 15690
rect 20520 15530 20530 15550
rect 20550 15530 20560 15550
rect 20520 15390 20560 15530
rect 20520 15370 20530 15390
rect 20550 15370 20560 15390
rect 20520 15230 20560 15370
rect 20520 15210 20530 15230
rect 20550 15210 20560 15230
rect 20520 15200 20560 15210
rect 20600 16190 20640 16200
rect 20600 16170 20610 16190
rect 20630 16170 20640 16190
rect 20600 16030 20640 16170
rect 20600 16010 20610 16030
rect 20630 16010 20640 16030
rect 20600 15870 20640 16010
rect 20600 15850 20610 15870
rect 20630 15850 20640 15870
rect 20600 15710 20640 15850
rect 20600 15690 20610 15710
rect 20630 15690 20640 15710
rect 20600 15550 20640 15690
rect 20600 15530 20610 15550
rect 20630 15530 20640 15550
rect 20600 15390 20640 15530
rect 20600 15370 20610 15390
rect 20630 15370 20640 15390
rect 20600 15230 20640 15370
rect 20600 15210 20610 15230
rect 20630 15210 20640 15230
rect 20600 15200 20640 15210
rect 20680 16190 20720 16200
rect 20680 16170 20690 16190
rect 20710 16170 20720 16190
rect 20680 16030 20720 16170
rect 20680 16010 20690 16030
rect 20710 16010 20720 16030
rect 20680 15870 20720 16010
rect 20680 15850 20690 15870
rect 20710 15850 20720 15870
rect 20680 15710 20720 15850
rect 20680 15690 20690 15710
rect 20710 15690 20720 15710
rect 20680 15550 20720 15690
rect 20680 15530 20690 15550
rect 20710 15530 20720 15550
rect 20680 15390 20720 15530
rect 20680 15370 20690 15390
rect 20710 15370 20720 15390
rect 20680 15230 20720 15370
rect 20680 15210 20690 15230
rect 20710 15210 20720 15230
rect 20680 15200 20720 15210
rect 20760 16190 20800 16200
rect 20760 16170 20770 16190
rect 20790 16170 20800 16190
rect 20760 16030 20800 16170
rect 20760 16010 20770 16030
rect 20790 16010 20800 16030
rect 20760 15870 20800 16010
rect 20760 15850 20770 15870
rect 20790 15850 20800 15870
rect 20760 15710 20800 15850
rect 20760 15690 20770 15710
rect 20790 15690 20800 15710
rect 20760 15550 20800 15690
rect 20760 15530 20770 15550
rect 20790 15530 20800 15550
rect 20760 15390 20800 15530
rect 20760 15370 20770 15390
rect 20790 15370 20800 15390
rect 20760 15230 20800 15370
rect 20760 15210 20770 15230
rect 20790 15210 20800 15230
rect 20760 15200 20800 15210
rect 20840 16190 20880 16200
rect 20840 16170 20850 16190
rect 20870 16170 20880 16190
rect 20840 16030 20880 16170
rect 20840 16010 20850 16030
rect 20870 16010 20880 16030
rect 20840 15870 20880 16010
rect 20840 15850 20850 15870
rect 20870 15850 20880 15870
rect 20840 15710 20880 15850
rect 20840 15690 20850 15710
rect 20870 15690 20880 15710
rect 20840 15550 20880 15690
rect 20840 15530 20850 15550
rect 20870 15530 20880 15550
rect 20840 15390 20880 15530
rect 20840 15370 20850 15390
rect 20870 15370 20880 15390
rect 20840 15230 20880 15370
rect 20840 15210 20850 15230
rect 20870 15210 20880 15230
rect 20840 15200 20880 15210
rect 20920 16190 20960 16200
rect 20920 16170 20930 16190
rect 20950 16170 20960 16190
rect 20920 16030 20960 16170
rect 20920 16010 20930 16030
rect 20950 16010 20960 16030
rect 20920 15870 20960 16010
rect 20920 15850 20930 15870
rect 20950 15850 20960 15870
rect 20920 15710 20960 15850
rect 20920 15690 20930 15710
rect 20950 15690 20960 15710
rect 20920 15550 20960 15690
rect 20920 15530 20930 15550
rect 20950 15530 20960 15550
rect 20920 15390 20960 15530
rect 20920 15370 20930 15390
rect 20950 15370 20960 15390
rect 20920 15230 20960 15370
rect 20920 15210 20930 15230
rect 20950 15210 20960 15230
rect 20920 15200 20960 15210
rect 0 15150 40 15160
rect 0 15130 10 15150
rect 30 15130 40 15150
rect 0 14990 40 15130
rect 0 14970 10 14990
rect 30 14970 40 14990
rect 0 14960 40 14970
rect 80 15150 120 15160
rect 80 15130 90 15150
rect 110 15130 120 15150
rect 80 14990 120 15130
rect 80 14970 90 14990
rect 110 14970 120 14990
rect 80 14960 120 14970
rect 160 15150 200 15160
rect 160 15130 170 15150
rect 190 15130 200 15150
rect 160 14990 200 15130
rect 160 14970 170 14990
rect 190 14970 200 14990
rect 160 14960 200 14970
rect 240 15150 280 15160
rect 240 15130 250 15150
rect 270 15130 280 15150
rect 240 14990 280 15130
rect 240 14970 250 14990
rect 270 14970 280 14990
rect 240 14960 280 14970
rect 320 15150 360 15160
rect 320 15130 330 15150
rect 350 15130 360 15150
rect 320 14990 360 15130
rect 320 14970 330 14990
rect 350 14970 360 14990
rect 320 14960 360 14970
rect 400 15150 440 15160
rect 400 15130 410 15150
rect 430 15130 440 15150
rect 400 14990 440 15130
rect 400 14970 410 14990
rect 430 14970 440 14990
rect 400 14960 440 14970
rect 480 15150 520 15160
rect 480 15130 490 15150
rect 510 15130 520 15150
rect 480 14990 520 15130
rect 480 14970 490 14990
rect 510 14970 520 14990
rect 480 14960 520 14970
rect 560 15150 600 15160
rect 560 15130 570 15150
rect 590 15130 600 15150
rect 560 14990 600 15130
rect 560 14970 570 14990
rect 590 14970 600 14990
rect 560 14960 600 14970
rect 640 15150 680 15160
rect 640 15130 650 15150
rect 670 15130 680 15150
rect 640 14990 680 15130
rect 640 14970 650 14990
rect 670 14970 680 14990
rect 640 14960 680 14970
rect 720 15150 760 15160
rect 720 15130 730 15150
rect 750 15130 760 15150
rect 720 14990 760 15130
rect 720 14970 730 14990
rect 750 14970 760 14990
rect 720 14960 760 14970
rect 800 15150 840 15160
rect 800 15130 810 15150
rect 830 15130 840 15150
rect 800 14990 840 15130
rect 800 14970 810 14990
rect 830 14970 840 14990
rect 800 14960 840 14970
rect 880 15150 920 15160
rect 880 15130 890 15150
rect 910 15130 920 15150
rect 880 14990 920 15130
rect 880 14970 890 14990
rect 910 14970 920 14990
rect 880 14960 920 14970
rect 960 15150 1000 15160
rect 960 15130 970 15150
rect 990 15130 1000 15150
rect 960 14990 1000 15130
rect 960 14970 970 14990
rect 990 14970 1000 14990
rect 960 14960 1000 14970
rect 1040 15150 1080 15160
rect 1040 15130 1050 15150
rect 1070 15130 1080 15150
rect 1040 14990 1080 15130
rect 1040 14970 1050 14990
rect 1070 14970 1080 14990
rect 1040 14960 1080 14970
rect 1120 15150 1160 15160
rect 1120 15130 1130 15150
rect 1150 15130 1160 15150
rect 1120 14990 1160 15130
rect 1120 14970 1130 14990
rect 1150 14970 1160 14990
rect 1120 14960 1160 14970
rect 1200 15150 1240 15160
rect 1200 15130 1210 15150
rect 1230 15130 1240 15150
rect 1200 14990 1240 15130
rect 1200 14970 1210 14990
rect 1230 14970 1240 14990
rect 1200 14960 1240 14970
rect 1280 15150 1320 15160
rect 1280 15130 1290 15150
rect 1310 15130 1320 15150
rect 1280 14990 1320 15130
rect 1280 14970 1290 14990
rect 1310 14970 1320 14990
rect 1280 14960 1320 14970
rect 1360 15150 1400 15160
rect 1360 15130 1370 15150
rect 1390 15130 1400 15150
rect 1360 14990 1400 15130
rect 1360 14970 1370 14990
rect 1390 14970 1400 14990
rect 1360 14960 1400 14970
rect 1440 15150 1480 15160
rect 1440 15130 1450 15150
rect 1470 15130 1480 15150
rect 1440 14990 1480 15130
rect 1440 14970 1450 14990
rect 1470 14970 1480 14990
rect 1440 14960 1480 14970
rect 1520 15150 1560 15160
rect 1520 15130 1530 15150
rect 1550 15130 1560 15150
rect 1520 14990 1560 15130
rect 1520 14970 1530 14990
rect 1550 14970 1560 14990
rect 1520 14960 1560 14970
rect 1600 15150 1640 15160
rect 1600 15130 1610 15150
rect 1630 15130 1640 15150
rect 1600 14990 1640 15130
rect 1600 14970 1610 14990
rect 1630 14970 1640 14990
rect 1600 14960 1640 14970
rect 1680 15150 1720 15160
rect 1680 15130 1690 15150
rect 1710 15130 1720 15150
rect 1680 14990 1720 15130
rect 1680 14970 1690 14990
rect 1710 14970 1720 14990
rect 1680 14960 1720 14970
rect 1760 15150 1800 15160
rect 1760 15130 1770 15150
rect 1790 15130 1800 15150
rect 1760 14990 1800 15130
rect 1760 14970 1770 14990
rect 1790 14970 1800 14990
rect 1760 14960 1800 14970
rect 1840 15150 1880 15160
rect 1840 15130 1850 15150
rect 1870 15130 1880 15150
rect 1840 14990 1880 15130
rect 1840 14970 1850 14990
rect 1870 14970 1880 14990
rect 1840 14960 1880 14970
rect 1920 15150 1960 15160
rect 1920 15130 1930 15150
rect 1950 15130 1960 15150
rect 1920 14990 1960 15130
rect 1920 14970 1930 14990
rect 1950 14970 1960 14990
rect 1920 14960 1960 14970
rect 2000 15150 2040 15160
rect 2000 15130 2010 15150
rect 2030 15130 2040 15150
rect 2000 14990 2040 15130
rect 2000 14970 2010 14990
rect 2030 14970 2040 14990
rect 2000 14960 2040 14970
rect 2080 15150 2120 15160
rect 2080 15130 2090 15150
rect 2110 15130 2120 15150
rect 2080 14990 2120 15130
rect 2080 14970 2090 14990
rect 2110 14970 2120 14990
rect 2080 14960 2120 14970
rect 2160 15150 2200 15160
rect 2160 15130 2170 15150
rect 2190 15130 2200 15150
rect 2160 14990 2200 15130
rect 2160 14970 2170 14990
rect 2190 14970 2200 14990
rect 2160 14960 2200 14970
rect 2240 15150 2280 15160
rect 2240 15130 2250 15150
rect 2270 15130 2280 15150
rect 2240 14990 2280 15130
rect 2240 14970 2250 14990
rect 2270 14970 2280 14990
rect 2240 14960 2280 14970
rect 2320 15150 2360 15160
rect 2320 15130 2330 15150
rect 2350 15130 2360 15150
rect 2320 14990 2360 15130
rect 2320 14970 2330 14990
rect 2350 14970 2360 14990
rect 2320 14960 2360 14970
rect 2400 15150 2440 15160
rect 2400 15130 2410 15150
rect 2430 15130 2440 15150
rect 2400 14990 2440 15130
rect 2400 14970 2410 14990
rect 2430 14970 2440 14990
rect 2400 14960 2440 14970
rect 2480 15150 2520 15160
rect 2480 15130 2490 15150
rect 2510 15130 2520 15150
rect 2480 14990 2520 15130
rect 2480 14970 2490 14990
rect 2510 14970 2520 14990
rect 2480 14960 2520 14970
rect 2560 15150 2600 15160
rect 2560 15130 2570 15150
rect 2590 15130 2600 15150
rect 2560 14990 2600 15130
rect 2560 14970 2570 14990
rect 2590 14970 2600 14990
rect 2560 14960 2600 14970
rect 2640 15150 2680 15160
rect 2640 15130 2650 15150
rect 2670 15130 2680 15150
rect 2640 14990 2680 15130
rect 2640 14970 2650 14990
rect 2670 14970 2680 14990
rect 2640 14960 2680 14970
rect 2720 15150 2760 15160
rect 2720 15130 2730 15150
rect 2750 15130 2760 15150
rect 2720 14990 2760 15130
rect 2720 14970 2730 14990
rect 2750 14970 2760 14990
rect 2720 14960 2760 14970
rect 2800 15150 2840 15160
rect 2800 15130 2810 15150
rect 2830 15130 2840 15150
rect 2800 14990 2840 15130
rect 2800 14970 2810 14990
rect 2830 14970 2840 14990
rect 2800 14960 2840 14970
rect 2880 15150 2920 15160
rect 2880 15130 2890 15150
rect 2910 15130 2920 15150
rect 2880 14990 2920 15130
rect 2880 14970 2890 14990
rect 2910 14970 2920 14990
rect 2880 14960 2920 14970
rect 2960 15150 3000 15160
rect 2960 15130 2970 15150
rect 2990 15130 3000 15150
rect 2960 14990 3000 15130
rect 2960 14970 2970 14990
rect 2990 14970 3000 14990
rect 2960 14960 3000 14970
rect 3040 15150 3080 15160
rect 3040 15130 3050 15150
rect 3070 15130 3080 15150
rect 3040 14990 3080 15130
rect 3040 14970 3050 14990
rect 3070 14970 3080 14990
rect 3040 14960 3080 14970
rect 3120 15150 3160 15160
rect 3120 15130 3130 15150
rect 3150 15130 3160 15150
rect 3120 14990 3160 15130
rect 3120 14970 3130 14990
rect 3150 14970 3160 14990
rect 3120 14960 3160 14970
rect 3200 15150 3240 15160
rect 3200 15130 3210 15150
rect 3230 15130 3240 15150
rect 3200 14990 3240 15130
rect 3200 14970 3210 14990
rect 3230 14970 3240 14990
rect 3200 14960 3240 14970
rect 3280 15150 3320 15160
rect 3280 15130 3290 15150
rect 3310 15130 3320 15150
rect 3280 14990 3320 15130
rect 3280 14970 3290 14990
rect 3310 14970 3320 14990
rect 3280 14960 3320 14970
rect 3360 15150 3400 15160
rect 3360 15130 3370 15150
rect 3390 15130 3400 15150
rect 3360 14990 3400 15130
rect 3360 14970 3370 14990
rect 3390 14970 3400 14990
rect 3360 14960 3400 14970
rect 3440 15150 3480 15160
rect 3440 15130 3450 15150
rect 3470 15130 3480 15150
rect 3440 14990 3480 15130
rect 3440 14970 3450 14990
rect 3470 14970 3480 14990
rect 3440 14960 3480 14970
rect 3520 15150 3560 15160
rect 3520 15130 3530 15150
rect 3550 15130 3560 15150
rect 3520 14990 3560 15130
rect 3520 14970 3530 14990
rect 3550 14970 3560 14990
rect 3520 14960 3560 14970
rect 3600 15150 3640 15160
rect 3600 15130 3610 15150
rect 3630 15130 3640 15150
rect 3600 14990 3640 15130
rect 3600 14970 3610 14990
rect 3630 14970 3640 14990
rect 3600 14960 3640 14970
rect 3680 15150 3720 15160
rect 3680 15130 3690 15150
rect 3710 15130 3720 15150
rect 3680 14990 3720 15130
rect 3680 14970 3690 14990
rect 3710 14970 3720 14990
rect 3680 14960 3720 14970
rect 3760 15150 3800 15160
rect 3760 15130 3770 15150
rect 3790 15130 3800 15150
rect 3760 14990 3800 15130
rect 3760 14970 3770 14990
rect 3790 14970 3800 14990
rect 3760 14960 3800 14970
rect 3840 15150 3880 15160
rect 3840 15130 3850 15150
rect 3870 15130 3880 15150
rect 3840 14990 3880 15130
rect 3840 14970 3850 14990
rect 3870 14970 3880 14990
rect 3840 14960 3880 14970
rect 3920 15150 3960 15160
rect 3920 15130 3930 15150
rect 3950 15130 3960 15150
rect 3920 14990 3960 15130
rect 3920 14970 3930 14990
rect 3950 14970 3960 14990
rect 3920 14960 3960 14970
rect 4000 15150 4040 15160
rect 4000 15130 4010 15150
rect 4030 15130 4040 15150
rect 4000 14990 4040 15130
rect 4000 14970 4010 14990
rect 4030 14970 4040 14990
rect 4000 14960 4040 14970
rect 4080 15150 4120 15160
rect 4080 15130 4090 15150
rect 4110 15130 4120 15150
rect 4080 14990 4120 15130
rect 4080 14970 4090 14990
rect 4110 14970 4120 14990
rect 4080 14960 4120 14970
rect 4160 15150 4200 15160
rect 4160 15130 4170 15150
rect 4190 15130 4200 15150
rect 4160 14990 4200 15130
rect 4160 14970 4170 14990
rect 4190 14970 4200 14990
rect 4160 14960 4200 14970
rect 4240 14960 4280 15160
rect 4320 14960 4360 15160
rect 4400 14960 4440 15160
rect 4480 14960 4520 15160
rect 4560 14960 4600 15160
rect 4640 14960 4680 15160
rect 4720 14960 4760 15160
rect 4800 14960 4840 15160
rect 4880 14960 4920 15160
rect 4960 14960 5000 15160
rect 5040 14960 5080 15160
rect 5120 14960 5160 15160
rect 5200 14960 5240 15160
rect 5280 14960 5320 15160
rect 5360 14960 5400 15160
rect 5440 14960 5480 15160
rect 5520 14960 5560 15160
rect 5600 14960 5640 15160
rect 5680 14960 5720 15160
rect 5760 14960 5800 15160
rect 5840 14960 5880 15160
rect 5920 14960 5960 15160
rect 6000 14960 6040 15160
rect 6080 14960 6120 15160
rect 6160 14960 6200 15160
rect 6240 15150 6280 15160
rect 6240 15130 6250 15150
rect 6270 15130 6280 15150
rect 6240 14990 6280 15130
rect 6240 14970 6250 14990
rect 6270 14970 6280 14990
rect 6240 14960 6280 14970
rect 6320 15150 6360 15160
rect 6320 15130 6330 15150
rect 6350 15130 6360 15150
rect 6320 14990 6360 15130
rect 6320 14970 6330 14990
rect 6350 14970 6360 14990
rect 6320 14960 6360 14970
rect 6400 15150 6440 15160
rect 6400 15130 6410 15150
rect 6430 15130 6440 15150
rect 6400 14990 6440 15130
rect 6400 14970 6410 14990
rect 6430 14970 6440 14990
rect 6400 14960 6440 14970
rect 6480 15150 6520 15160
rect 6480 15130 6490 15150
rect 6510 15130 6520 15150
rect 6480 14990 6520 15130
rect 6480 14970 6490 14990
rect 6510 14970 6520 14990
rect 6480 14960 6520 14970
rect 6560 15150 6600 15160
rect 6560 15130 6570 15150
rect 6590 15130 6600 15150
rect 6560 14990 6600 15130
rect 6560 14970 6570 14990
rect 6590 14970 6600 14990
rect 6560 14960 6600 14970
rect 6640 15150 6680 15160
rect 6640 15130 6650 15150
rect 6670 15130 6680 15150
rect 6640 14990 6680 15130
rect 6640 14970 6650 14990
rect 6670 14970 6680 14990
rect 6640 14960 6680 14970
rect 6720 15150 6760 15160
rect 6720 15130 6730 15150
rect 6750 15130 6760 15150
rect 6720 14990 6760 15130
rect 6720 14970 6730 14990
rect 6750 14970 6760 14990
rect 6720 14960 6760 14970
rect 6800 15150 6840 15160
rect 6800 15130 6810 15150
rect 6830 15130 6840 15150
rect 6800 14990 6840 15130
rect 6800 14970 6810 14990
rect 6830 14970 6840 14990
rect 6800 14960 6840 14970
rect 6880 15150 6920 15160
rect 6880 15130 6890 15150
rect 6910 15130 6920 15150
rect 6880 14990 6920 15130
rect 6880 14970 6890 14990
rect 6910 14970 6920 14990
rect 6880 14960 6920 14970
rect 6960 15150 7000 15160
rect 6960 15130 6970 15150
rect 6990 15130 7000 15150
rect 6960 14990 7000 15130
rect 6960 14970 6970 14990
rect 6990 14970 7000 14990
rect 6960 14960 7000 14970
rect 7040 15150 7080 15160
rect 7040 15130 7050 15150
rect 7070 15130 7080 15150
rect 7040 14990 7080 15130
rect 7040 14970 7050 14990
rect 7070 14970 7080 14990
rect 7040 14960 7080 14970
rect 7120 15150 7160 15160
rect 7120 15130 7130 15150
rect 7150 15130 7160 15150
rect 7120 14990 7160 15130
rect 7120 14970 7130 14990
rect 7150 14970 7160 14990
rect 7120 14960 7160 14970
rect 7200 15150 7240 15160
rect 7200 15130 7210 15150
rect 7230 15130 7240 15150
rect 7200 14990 7240 15130
rect 7200 14970 7210 14990
rect 7230 14970 7240 14990
rect 7200 14960 7240 14970
rect 7280 15150 7320 15160
rect 7280 15130 7290 15150
rect 7310 15130 7320 15150
rect 7280 14990 7320 15130
rect 7280 14970 7290 14990
rect 7310 14970 7320 14990
rect 7280 14960 7320 14970
rect 7360 15150 7400 15160
rect 7360 15130 7370 15150
rect 7390 15130 7400 15150
rect 7360 14990 7400 15130
rect 7360 14970 7370 14990
rect 7390 14970 7400 14990
rect 7360 14960 7400 14970
rect 7440 15150 7480 15160
rect 7440 15130 7450 15150
rect 7470 15130 7480 15150
rect 7440 14990 7480 15130
rect 7440 14970 7450 14990
rect 7470 14970 7480 14990
rect 7440 14960 7480 14970
rect 7520 15150 7560 15160
rect 7520 15130 7530 15150
rect 7550 15130 7560 15150
rect 7520 14990 7560 15130
rect 7520 14970 7530 14990
rect 7550 14970 7560 14990
rect 7520 14960 7560 14970
rect 7600 15150 7640 15160
rect 7600 15130 7610 15150
rect 7630 15130 7640 15150
rect 7600 14990 7640 15130
rect 7600 14970 7610 14990
rect 7630 14970 7640 14990
rect 7600 14960 7640 14970
rect 7680 15150 7720 15160
rect 7680 15130 7690 15150
rect 7710 15130 7720 15150
rect 7680 14990 7720 15130
rect 7680 14970 7690 14990
rect 7710 14970 7720 14990
rect 7680 14960 7720 14970
rect 7760 15150 7800 15160
rect 7760 15130 7770 15150
rect 7790 15130 7800 15150
rect 7760 14990 7800 15130
rect 7760 14970 7770 14990
rect 7790 14970 7800 14990
rect 7760 14960 7800 14970
rect 7840 15150 7880 15160
rect 7840 15130 7850 15150
rect 7870 15130 7880 15150
rect 7840 14990 7880 15130
rect 7840 14970 7850 14990
rect 7870 14970 7880 14990
rect 7840 14960 7880 14970
rect 7920 15150 7960 15160
rect 7920 15130 7930 15150
rect 7950 15130 7960 15150
rect 7920 14990 7960 15130
rect 7920 14970 7930 14990
rect 7950 14970 7960 14990
rect 7920 14960 7960 14970
rect 8000 15150 8040 15160
rect 8000 15130 8010 15150
rect 8030 15130 8040 15150
rect 8000 14990 8040 15130
rect 8000 14970 8010 14990
rect 8030 14970 8040 14990
rect 8000 14960 8040 14970
rect 8080 15150 8120 15160
rect 8080 15130 8090 15150
rect 8110 15130 8120 15150
rect 8080 14990 8120 15130
rect 8080 14970 8090 14990
rect 8110 14970 8120 14990
rect 8080 14960 8120 14970
rect 8160 15150 8200 15160
rect 8160 15130 8170 15150
rect 8190 15130 8200 15150
rect 8160 14990 8200 15130
rect 8160 14970 8170 14990
rect 8190 14970 8200 14990
rect 8160 14960 8200 14970
rect 8240 15150 8280 15160
rect 8240 15130 8250 15150
rect 8270 15130 8280 15150
rect 8240 14990 8280 15130
rect 8240 14970 8250 14990
rect 8270 14970 8280 14990
rect 8240 14960 8280 14970
rect 8320 15150 8360 15160
rect 8320 15130 8330 15150
rect 8350 15130 8360 15150
rect 8320 14990 8360 15130
rect 8320 14970 8330 14990
rect 8350 14970 8360 14990
rect 8320 14960 8360 14970
rect 8400 15150 8440 15160
rect 8400 15130 8410 15150
rect 8430 15130 8440 15150
rect 8400 14990 8440 15130
rect 8400 14970 8410 14990
rect 8430 14970 8440 14990
rect 8400 14960 8440 14970
rect 8480 15150 8520 15160
rect 8480 15130 8490 15150
rect 8510 15130 8520 15150
rect 8480 14990 8520 15130
rect 8480 14970 8490 14990
rect 8510 14970 8520 14990
rect 8480 14960 8520 14970
rect 8560 15150 8600 15160
rect 8560 15130 8570 15150
rect 8590 15130 8600 15150
rect 8560 14990 8600 15130
rect 8560 14970 8570 14990
rect 8590 14970 8600 14990
rect 8560 14960 8600 14970
rect 8640 15150 8680 15160
rect 8640 15130 8650 15150
rect 8670 15130 8680 15150
rect 8640 14990 8680 15130
rect 8640 14970 8650 14990
rect 8670 14970 8680 14990
rect 8640 14960 8680 14970
rect 8720 15150 8760 15160
rect 8720 15130 8730 15150
rect 8750 15130 8760 15150
rect 8720 14990 8760 15130
rect 8720 14970 8730 14990
rect 8750 14970 8760 14990
rect 8720 14960 8760 14970
rect 8800 15150 8840 15160
rect 8800 15130 8810 15150
rect 8830 15130 8840 15150
rect 8800 14990 8840 15130
rect 8800 14970 8810 14990
rect 8830 14970 8840 14990
rect 8800 14960 8840 14970
rect 8880 15150 8920 15160
rect 8880 15130 8890 15150
rect 8910 15130 8920 15150
rect 8880 14990 8920 15130
rect 8880 14970 8890 14990
rect 8910 14970 8920 14990
rect 8880 14960 8920 14970
rect 8960 15150 9000 15160
rect 8960 15130 8970 15150
rect 8990 15130 9000 15150
rect 8960 14990 9000 15130
rect 8960 14970 8970 14990
rect 8990 14970 9000 14990
rect 8960 14960 9000 14970
rect 9040 15150 9080 15160
rect 9040 15130 9050 15150
rect 9070 15130 9080 15150
rect 9040 14990 9080 15130
rect 9040 14970 9050 14990
rect 9070 14970 9080 14990
rect 9040 14960 9080 14970
rect 9120 15150 9160 15160
rect 9120 15130 9130 15150
rect 9150 15130 9160 15150
rect 9120 14990 9160 15130
rect 9120 14970 9130 14990
rect 9150 14970 9160 14990
rect 9120 14960 9160 14970
rect 9200 15150 9240 15160
rect 9200 15130 9210 15150
rect 9230 15130 9240 15150
rect 9200 14990 9240 15130
rect 9200 14970 9210 14990
rect 9230 14970 9240 14990
rect 9200 14960 9240 14970
rect 9280 15150 9320 15160
rect 9280 15130 9290 15150
rect 9310 15130 9320 15150
rect 9280 14990 9320 15130
rect 9280 14970 9290 14990
rect 9310 14970 9320 14990
rect 9280 14960 9320 14970
rect 9360 15150 9400 15160
rect 9360 15130 9370 15150
rect 9390 15130 9400 15150
rect 9360 14990 9400 15130
rect 9360 14970 9370 14990
rect 9390 14970 9400 14990
rect 9360 14960 9400 14970
rect 9440 15150 9480 15160
rect 9440 15130 9450 15150
rect 9470 15130 9480 15150
rect 9440 14990 9480 15130
rect 9440 14970 9450 14990
rect 9470 14970 9480 14990
rect 9440 14960 9480 14970
rect 9520 14960 9560 15160
rect 9600 14960 9640 15160
rect 9680 14960 9720 15160
rect 9760 14960 9800 15160
rect 9840 14960 9880 15160
rect 9920 14960 9960 15160
rect 10000 14960 10040 15160
rect 10080 14960 10120 15160
rect 10160 14960 10200 15160
rect 10240 14960 10280 15160
rect 10320 14960 10360 15160
rect 10400 14960 10440 15160
rect 10480 14960 10520 15160
rect 10560 14960 10600 15160
rect 10640 14960 10680 15160
rect 10720 14960 10760 15160
rect 10800 14960 10840 15160
rect 10880 14960 10920 15160
rect 10960 14960 11000 15160
rect 11040 14960 11080 15160
rect 11120 14960 11160 15160
rect 11200 14960 11240 15160
rect 11280 14960 11320 15160
rect 11360 14960 11400 15160
rect 11440 14960 11480 15160
rect 11560 15150 11600 15160
rect 11560 15130 11570 15150
rect 11590 15130 11600 15150
rect 11560 14990 11600 15130
rect 11560 14970 11570 14990
rect 11590 14970 11600 14990
rect 11560 14960 11600 14970
rect 11640 15150 11680 15160
rect 11640 15130 11650 15150
rect 11670 15130 11680 15150
rect 11640 14990 11680 15130
rect 11640 14970 11650 14990
rect 11670 14970 11680 14990
rect 11640 14960 11680 14970
rect 11720 15150 11760 15160
rect 11720 15130 11730 15150
rect 11750 15130 11760 15150
rect 11720 14990 11760 15130
rect 11720 14970 11730 14990
rect 11750 14970 11760 14990
rect 11720 14960 11760 14970
rect 11800 15150 11840 15160
rect 11800 15130 11810 15150
rect 11830 15130 11840 15150
rect 11800 14990 11840 15130
rect 11800 14970 11810 14990
rect 11830 14970 11840 14990
rect 11800 14960 11840 14970
rect 11880 15150 11920 15160
rect 11880 15130 11890 15150
rect 11910 15130 11920 15150
rect 11880 14990 11920 15130
rect 11880 14970 11890 14990
rect 11910 14970 11920 14990
rect 11880 14960 11920 14970
rect 11960 15150 12000 15160
rect 11960 15130 11970 15150
rect 11990 15130 12000 15150
rect 11960 14990 12000 15130
rect 11960 14970 11970 14990
rect 11990 14970 12000 14990
rect 11960 14960 12000 14970
rect 12040 15150 12080 15160
rect 12040 15130 12050 15150
rect 12070 15130 12080 15150
rect 12040 14990 12080 15130
rect 12040 14970 12050 14990
rect 12070 14970 12080 14990
rect 12040 14960 12080 14970
rect 12120 15150 12160 15160
rect 12120 15130 12130 15150
rect 12150 15130 12160 15150
rect 12120 14990 12160 15130
rect 12120 14970 12130 14990
rect 12150 14970 12160 14990
rect 12120 14960 12160 14970
rect 12200 15150 12240 15160
rect 12200 15130 12210 15150
rect 12230 15130 12240 15150
rect 12200 14990 12240 15130
rect 12200 14970 12210 14990
rect 12230 14970 12240 14990
rect 12200 14960 12240 14970
rect 12280 15150 12320 15160
rect 12280 15130 12290 15150
rect 12310 15130 12320 15150
rect 12280 14990 12320 15130
rect 12280 14970 12290 14990
rect 12310 14970 12320 14990
rect 12280 14960 12320 14970
rect 12360 15150 12400 15160
rect 12360 15130 12370 15150
rect 12390 15130 12400 15150
rect 12360 14990 12400 15130
rect 12360 14970 12370 14990
rect 12390 14970 12400 14990
rect 12360 14960 12400 14970
rect 12440 15150 12480 15160
rect 12440 15130 12450 15150
rect 12470 15130 12480 15150
rect 12440 14990 12480 15130
rect 12440 14970 12450 14990
rect 12470 14970 12480 14990
rect 12440 14960 12480 14970
rect 12520 15150 12560 15160
rect 12520 15130 12530 15150
rect 12550 15130 12560 15150
rect 12520 14990 12560 15130
rect 12520 14970 12530 14990
rect 12550 14970 12560 14990
rect 12520 14960 12560 14970
rect 12600 15150 12640 15160
rect 12600 15130 12610 15150
rect 12630 15130 12640 15150
rect 12600 14990 12640 15130
rect 12600 14970 12610 14990
rect 12630 14970 12640 14990
rect 12600 14960 12640 14970
rect 12680 15150 12720 15160
rect 12680 15130 12690 15150
rect 12710 15130 12720 15150
rect 12680 14990 12720 15130
rect 12680 14970 12690 14990
rect 12710 14970 12720 14990
rect 12680 14960 12720 14970
rect 12760 15150 12800 15160
rect 12760 15130 12770 15150
rect 12790 15130 12800 15150
rect 12760 14990 12800 15130
rect 12760 14970 12770 14990
rect 12790 14970 12800 14990
rect 12760 14960 12800 14970
rect 12840 15150 12880 15160
rect 12840 15130 12850 15150
rect 12870 15130 12880 15150
rect 12840 14990 12880 15130
rect 12840 14970 12850 14990
rect 12870 14970 12880 14990
rect 12840 14960 12880 14970
rect 12920 15150 12960 15160
rect 12920 15130 12930 15150
rect 12950 15130 12960 15150
rect 12920 14990 12960 15130
rect 12920 14970 12930 14990
rect 12950 14970 12960 14990
rect 12920 14960 12960 14970
rect 13000 15150 13040 15160
rect 13000 15130 13010 15150
rect 13030 15130 13040 15150
rect 13000 14990 13040 15130
rect 13000 14970 13010 14990
rect 13030 14970 13040 14990
rect 13000 14960 13040 14970
rect 13080 15150 13120 15160
rect 13080 15130 13090 15150
rect 13110 15130 13120 15150
rect 13080 14990 13120 15130
rect 13080 14970 13090 14990
rect 13110 14970 13120 14990
rect 13080 14960 13120 14970
rect 13160 15150 13200 15160
rect 13160 15130 13170 15150
rect 13190 15130 13200 15150
rect 13160 14990 13200 15130
rect 13160 14970 13170 14990
rect 13190 14970 13200 14990
rect 13160 14960 13200 14970
rect 13240 15150 13280 15160
rect 13240 15130 13250 15150
rect 13270 15130 13280 15150
rect 13240 14990 13280 15130
rect 13240 14970 13250 14990
rect 13270 14970 13280 14990
rect 13240 14960 13280 14970
rect 13320 15150 13360 15160
rect 13320 15130 13330 15150
rect 13350 15130 13360 15150
rect 13320 14990 13360 15130
rect 13320 14970 13330 14990
rect 13350 14970 13360 14990
rect 13320 14960 13360 14970
rect 13400 15150 13440 15160
rect 13400 15130 13410 15150
rect 13430 15130 13440 15150
rect 13400 14990 13440 15130
rect 13400 14970 13410 14990
rect 13430 14970 13440 14990
rect 13400 14960 13440 14970
rect 13480 15150 13520 15160
rect 13480 15130 13490 15150
rect 13510 15130 13520 15150
rect 13480 14990 13520 15130
rect 13480 14970 13490 14990
rect 13510 14970 13520 14990
rect 13480 14960 13520 14970
rect 13560 15150 13600 15160
rect 13560 15130 13570 15150
rect 13590 15130 13600 15150
rect 13560 14990 13600 15130
rect 13560 14970 13570 14990
rect 13590 14970 13600 14990
rect 13560 14960 13600 14970
rect 13640 15150 13680 15160
rect 13640 15130 13650 15150
rect 13670 15130 13680 15150
rect 13640 14990 13680 15130
rect 13640 14970 13650 14990
rect 13670 14970 13680 14990
rect 13640 14960 13680 14970
rect 13720 15150 13760 15160
rect 13720 15130 13730 15150
rect 13750 15130 13760 15150
rect 13720 14990 13760 15130
rect 13720 14970 13730 14990
rect 13750 14970 13760 14990
rect 13720 14960 13760 14970
rect 13800 15150 13840 15160
rect 13800 15130 13810 15150
rect 13830 15130 13840 15150
rect 13800 14990 13840 15130
rect 13800 14970 13810 14990
rect 13830 14970 13840 14990
rect 13800 14960 13840 14970
rect 13880 15150 13920 15160
rect 13880 15130 13890 15150
rect 13910 15130 13920 15150
rect 13880 14990 13920 15130
rect 13880 14970 13890 14990
rect 13910 14970 13920 14990
rect 13880 14960 13920 14970
rect 13960 15150 14000 15160
rect 13960 15130 13970 15150
rect 13990 15130 14000 15150
rect 13960 14990 14000 15130
rect 13960 14970 13970 14990
rect 13990 14970 14000 14990
rect 13960 14960 14000 14970
rect 14040 15150 14080 15160
rect 14040 15130 14050 15150
rect 14070 15130 14080 15150
rect 14040 14990 14080 15130
rect 14040 14970 14050 14990
rect 14070 14970 14080 14990
rect 14040 14960 14080 14970
rect 14120 15150 14160 15160
rect 14120 15130 14130 15150
rect 14150 15130 14160 15150
rect 14120 14990 14160 15130
rect 14120 14970 14130 14990
rect 14150 14970 14160 14990
rect 14120 14960 14160 14970
rect 14200 15150 14240 15160
rect 14200 15130 14210 15150
rect 14230 15130 14240 15150
rect 14200 14990 14240 15130
rect 14200 14970 14210 14990
rect 14230 14970 14240 14990
rect 14200 14960 14240 14970
rect 14280 15150 14320 15160
rect 14280 15130 14290 15150
rect 14310 15130 14320 15150
rect 14280 14990 14320 15130
rect 14280 14970 14290 14990
rect 14310 14970 14320 14990
rect 14280 14960 14320 14970
rect 14360 15150 14400 15160
rect 14360 15130 14370 15150
rect 14390 15130 14400 15150
rect 14360 14990 14400 15130
rect 14360 14970 14370 14990
rect 14390 14970 14400 14990
rect 14360 14960 14400 14970
rect 14440 15150 14480 15160
rect 14440 15130 14450 15150
rect 14470 15130 14480 15150
rect 14440 14990 14480 15130
rect 14440 14970 14450 14990
rect 14470 14970 14480 14990
rect 14440 14960 14480 14970
rect 14520 15150 14560 15160
rect 14520 15130 14530 15150
rect 14550 15130 14560 15150
rect 14520 14990 14560 15130
rect 14520 14970 14530 14990
rect 14550 14970 14560 14990
rect 14520 14960 14560 14970
rect 14600 15150 14640 15160
rect 14600 15130 14610 15150
rect 14630 15130 14640 15150
rect 14600 14990 14640 15130
rect 14600 14970 14610 14990
rect 14630 14970 14640 14990
rect 14600 14960 14640 14970
rect 14680 15150 14720 15160
rect 14680 15130 14690 15150
rect 14710 15130 14720 15150
rect 14680 14990 14720 15130
rect 14680 14970 14690 14990
rect 14710 14970 14720 14990
rect 14680 14960 14720 14970
rect 14760 14960 14800 15160
rect 14840 14960 14880 15160
rect 14920 14960 14960 15160
rect 15000 14960 15040 15160
rect 15080 14960 15120 15160
rect 15160 14960 15200 15160
rect 15240 14960 15280 15160
rect 15320 14960 15360 15160
rect 15400 14960 15440 15160
rect 15480 14960 15520 15160
rect 15560 14960 15600 15160
rect 15640 14960 15680 15160
rect 15720 14960 15760 15160
rect 15800 14960 15840 15160
rect 15880 14960 15920 15160
rect 15960 14960 16000 15160
rect 16040 14960 16080 15160
rect 16120 14960 16160 15160
rect 16200 14960 16240 15160
rect 16280 14960 16320 15160
rect 16360 14960 16400 15160
rect 16440 14960 16480 15160
rect 16520 14960 16560 15160
rect 16600 14960 16640 15160
rect 16680 14960 16720 15160
rect 16760 15150 16800 15160
rect 16760 15130 16770 15150
rect 16790 15130 16800 15150
rect 16760 14990 16800 15130
rect 16760 14970 16770 14990
rect 16790 14970 16800 14990
rect 16760 14960 16800 14970
rect 16840 15150 16880 15160
rect 16840 15130 16850 15150
rect 16870 15130 16880 15150
rect 16840 14990 16880 15130
rect 16840 14970 16850 14990
rect 16870 14970 16880 14990
rect 16840 14960 16880 14970
rect 16920 15150 16960 15160
rect 16920 15130 16930 15150
rect 16950 15130 16960 15150
rect 16920 14990 16960 15130
rect 16920 14970 16930 14990
rect 16950 14970 16960 14990
rect 16920 14960 16960 14970
rect 17000 15150 17040 15160
rect 17000 15130 17010 15150
rect 17030 15130 17040 15150
rect 17000 14990 17040 15130
rect 17000 14970 17010 14990
rect 17030 14970 17040 14990
rect 17000 14960 17040 14970
rect 17080 15150 17120 15160
rect 17080 15130 17090 15150
rect 17110 15130 17120 15150
rect 17080 14990 17120 15130
rect 17080 14970 17090 14990
rect 17110 14970 17120 14990
rect 17080 14960 17120 14970
rect 17160 15150 17200 15160
rect 17160 15130 17170 15150
rect 17190 15130 17200 15150
rect 17160 14990 17200 15130
rect 17160 14970 17170 14990
rect 17190 14970 17200 14990
rect 17160 14960 17200 14970
rect 17240 15150 17280 15160
rect 17240 15130 17250 15150
rect 17270 15130 17280 15150
rect 17240 14990 17280 15130
rect 17240 14970 17250 14990
rect 17270 14970 17280 14990
rect 17240 14960 17280 14970
rect 17320 15150 17360 15160
rect 17320 15130 17330 15150
rect 17350 15130 17360 15150
rect 17320 14990 17360 15130
rect 17320 14970 17330 14990
rect 17350 14970 17360 14990
rect 17320 14960 17360 14970
rect 17400 15150 17440 15160
rect 17400 15130 17410 15150
rect 17430 15130 17440 15150
rect 17400 14990 17440 15130
rect 17400 14970 17410 14990
rect 17430 14970 17440 14990
rect 17400 14960 17440 14970
rect 17480 15150 17520 15160
rect 17480 15130 17490 15150
rect 17510 15130 17520 15150
rect 17480 14990 17520 15130
rect 17480 14970 17490 14990
rect 17510 14970 17520 14990
rect 17480 14960 17520 14970
rect 17560 15150 17600 15160
rect 17560 15130 17570 15150
rect 17590 15130 17600 15150
rect 17560 14990 17600 15130
rect 17560 14970 17570 14990
rect 17590 14970 17600 14990
rect 17560 14960 17600 14970
rect 17640 15150 17680 15160
rect 17640 15130 17650 15150
rect 17670 15130 17680 15150
rect 17640 14990 17680 15130
rect 17640 14970 17650 14990
rect 17670 14970 17680 14990
rect 17640 14960 17680 14970
rect 17720 15150 17760 15160
rect 17720 15130 17730 15150
rect 17750 15130 17760 15150
rect 17720 14990 17760 15130
rect 17720 14970 17730 14990
rect 17750 14970 17760 14990
rect 17720 14960 17760 14970
rect 17800 15150 17840 15160
rect 17800 15130 17810 15150
rect 17830 15130 17840 15150
rect 17800 14990 17840 15130
rect 17800 14970 17810 14990
rect 17830 14970 17840 14990
rect 17800 14960 17840 14970
rect 17880 15150 17920 15160
rect 17880 15130 17890 15150
rect 17910 15130 17920 15150
rect 17880 14990 17920 15130
rect 17880 14970 17890 14990
rect 17910 14970 17920 14990
rect 17880 14960 17920 14970
rect 17960 15150 18000 15160
rect 17960 15130 17970 15150
rect 17990 15130 18000 15150
rect 17960 14990 18000 15130
rect 17960 14970 17970 14990
rect 17990 14970 18000 14990
rect 17960 14960 18000 14970
rect 18040 15150 18080 15160
rect 18040 15130 18050 15150
rect 18070 15130 18080 15150
rect 18040 14990 18080 15130
rect 18040 14970 18050 14990
rect 18070 14970 18080 14990
rect 18040 14960 18080 14970
rect 18120 15150 18160 15160
rect 18120 15130 18130 15150
rect 18150 15130 18160 15150
rect 18120 14990 18160 15130
rect 18120 14970 18130 14990
rect 18150 14970 18160 14990
rect 18120 14960 18160 14970
rect 18200 15150 18240 15160
rect 18200 15130 18210 15150
rect 18230 15130 18240 15150
rect 18200 14990 18240 15130
rect 18200 14970 18210 14990
rect 18230 14970 18240 14990
rect 18200 14960 18240 14970
rect 18280 15150 18320 15160
rect 18280 15130 18290 15150
rect 18310 15130 18320 15150
rect 18280 14990 18320 15130
rect 18280 14970 18290 14990
rect 18310 14970 18320 14990
rect 18280 14960 18320 14970
rect 18360 15150 18400 15160
rect 18360 15130 18370 15150
rect 18390 15130 18400 15150
rect 18360 14990 18400 15130
rect 18360 14970 18370 14990
rect 18390 14970 18400 14990
rect 18360 14960 18400 14970
rect 18440 15150 18480 15160
rect 18440 15130 18450 15150
rect 18470 15130 18480 15150
rect 18440 14990 18480 15130
rect 18440 14970 18450 14990
rect 18470 14970 18480 14990
rect 18440 14960 18480 14970
rect 18520 15150 18560 15160
rect 18520 15130 18530 15150
rect 18550 15130 18560 15150
rect 18520 14990 18560 15130
rect 18520 14970 18530 14990
rect 18550 14970 18560 14990
rect 18520 14960 18560 14970
rect 18600 15150 18640 15160
rect 18600 15130 18610 15150
rect 18630 15130 18640 15150
rect 18600 14990 18640 15130
rect 18600 14970 18610 14990
rect 18630 14970 18640 14990
rect 18600 14960 18640 14970
rect 18680 15150 18720 15160
rect 18680 15130 18690 15150
rect 18710 15130 18720 15150
rect 18680 14990 18720 15130
rect 18680 14970 18690 14990
rect 18710 14970 18720 14990
rect 18680 14960 18720 14970
rect 18760 15150 18800 15160
rect 18760 15130 18770 15150
rect 18790 15130 18800 15150
rect 18760 14990 18800 15130
rect 18760 14970 18770 14990
rect 18790 14970 18800 14990
rect 18760 14960 18800 14970
rect 18840 15150 18880 15160
rect 18840 15130 18850 15150
rect 18870 15130 18880 15150
rect 18840 14990 18880 15130
rect 18840 14970 18850 14990
rect 18870 14970 18880 14990
rect 18840 14960 18880 14970
rect 18920 15150 18960 15160
rect 18920 15130 18930 15150
rect 18950 15130 18960 15150
rect 18920 14990 18960 15130
rect 18920 14970 18930 14990
rect 18950 14970 18960 14990
rect 18920 14960 18960 14970
rect 19000 15150 19040 15160
rect 19000 15130 19010 15150
rect 19030 15130 19040 15150
rect 19000 14990 19040 15130
rect 19000 14970 19010 14990
rect 19030 14970 19040 14990
rect 19000 14960 19040 14970
rect 19080 15150 19120 15160
rect 19080 15130 19090 15150
rect 19110 15130 19120 15150
rect 19080 14990 19120 15130
rect 19080 14970 19090 14990
rect 19110 14970 19120 14990
rect 19080 14960 19120 14970
rect 19160 15150 19200 15160
rect 19160 15130 19170 15150
rect 19190 15130 19200 15150
rect 19160 14990 19200 15130
rect 19160 14970 19170 14990
rect 19190 14970 19200 14990
rect 19160 14960 19200 14970
rect 19240 15150 19280 15160
rect 19240 15130 19250 15150
rect 19270 15130 19280 15150
rect 19240 14990 19280 15130
rect 19240 14970 19250 14990
rect 19270 14970 19280 14990
rect 19240 14960 19280 14970
rect 19320 15150 19360 15160
rect 19320 15130 19330 15150
rect 19350 15130 19360 15150
rect 19320 14990 19360 15130
rect 19320 14970 19330 14990
rect 19350 14970 19360 14990
rect 19320 14960 19360 14970
rect 19400 15150 19440 15160
rect 19400 15130 19410 15150
rect 19430 15130 19440 15150
rect 19400 14990 19440 15130
rect 19400 14970 19410 14990
rect 19430 14970 19440 14990
rect 19400 14960 19440 14970
rect 19480 15150 19520 15160
rect 19480 15130 19490 15150
rect 19510 15130 19520 15150
rect 19480 14990 19520 15130
rect 19480 14970 19490 14990
rect 19510 14970 19520 14990
rect 19480 14960 19520 14970
rect 19560 15150 19600 15160
rect 19560 15130 19570 15150
rect 19590 15130 19600 15150
rect 19560 14990 19600 15130
rect 19560 14970 19570 14990
rect 19590 14970 19600 14990
rect 19560 14960 19600 14970
rect 19640 15150 19680 15160
rect 19640 15130 19650 15150
rect 19670 15130 19680 15150
rect 19640 14990 19680 15130
rect 19640 14970 19650 14990
rect 19670 14970 19680 14990
rect 19640 14960 19680 14970
rect 19720 15150 19760 15160
rect 19720 15130 19730 15150
rect 19750 15130 19760 15150
rect 19720 14990 19760 15130
rect 19720 14970 19730 14990
rect 19750 14970 19760 14990
rect 19720 14960 19760 14970
rect 19800 15150 19840 15160
rect 19800 15130 19810 15150
rect 19830 15130 19840 15150
rect 19800 14990 19840 15130
rect 19800 14970 19810 14990
rect 19830 14970 19840 14990
rect 19800 14960 19840 14970
rect 19880 15150 19920 15160
rect 19880 15130 19890 15150
rect 19910 15130 19920 15150
rect 19880 14990 19920 15130
rect 19880 14970 19890 14990
rect 19910 14970 19920 14990
rect 19880 14960 19920 14970
rect 19960 15150 20000 15160
rect 19960 15130 19970 15150
rect 19990 15130 20000 15150
rect 19960 14990 20000 15130
rect 19960 14970 19970 14990
rect 19990 14970 20000 14990
rect 19960 14960 20000 14970
rect 20040 15150 20080 15160
rect 20040 15130 20050 15150
rect 20070 15130 20080 15150
rect 20040 14990 20080 15130
rect 20040 14970 20050 14990
rect 20070 14970 20080 14990
rect 20040 14960 20080 14970
rect 20120 15150 20160 15160
rect 20120 15130 20130 15150
rect 20150 15130 20160 15150
rect 20120 14990 20160 15130
rect 20120 14970 20130 14990
rect 20150 14970 20160 14990
rect 20120 14960 20160 14970
rect 20200 15150 20240 15160
rect 20200 15130 20210 15150
rect 20230 15130 20240 15150
rect 20200 14990 20240 15130
rect 20200 14970 20210 14990
rect 20230 14970 20240 14990
rect 20200 14960 20240 14970
rect 20280 15150 20320 15160
rect 20280 15130 20290 15150
rect 20310 15130 20320 15150
rect 20280 14990 20320 15130
rect 20280 14970 20290 14990
rect 20310 14970 20320 14990
rect 20280 14960 20320 14970
rect 20360 15150 20400 15160
rect 20360 15130 20370 15150
rect 20390 15130 20400 15150
rect 20360 14990 20400 15130
rect 20360 14970 20370 14990
rect 20390 14970 20400 14990
rect 20360 14960 20400 14970
rect 20440 15150 20480 15160
rect 20440 15130 20450 15150
rect 20470 15130 20480 15150
rect 20440 14990 20480 15130
rect 20440 14970 20450 14990
rect 20470 14970 20480 14990
rect 20440 14960 20480 14970
rect 20520 15150 20560 15160
rect 20520 15130 20530 15150
rect 20550 15130 20560 15150
rect 20520 14990 20560 15130
rect 20520 14970 20530 14990
rect 20550 14970 20560 14990
rect 20520 14960 20560 14970
rect 20600 15150 20640 15160
rect 20600 15130 20610 15150
rect 20630 15130 20640 15150
rect 20600 14990 20640 15130
rect 20600 14970 20610 14990
rect 20630 14970 20640 14990
rect 20600 14960 20640 14970
rect 20680 15150 20720 15160
rect 20680 15130 20690 15150
rect 20710 15130 20720 15150
rect 20680 14990 20720 15130
rect 20680 14970 20690 14990
rect 20710 14970 20720 14990
rect 20680 14960 20720 14970
rect 20760 15150 20800 15160
rect 20760 15130 20770 15150
rect 20790 15130 20800 15150
rect 20760 14990 20800 15130
rect 20760 14970 20770 14990
rect 20790 14970 20800 14990
rect 20760 14960 20800 14970
rect 20840 15150 20880 15160
rect 20840 15130 20850 15150
rect 20870 15130 20880 15150
rect 20840 14990 20880 15130
rect 20840 14970 20850 14990
rect 20870 14970 20880 14990
rect 20840 14960 20880 14970
rect 20920 15150 20960 15160
rect 20920 15130 20930 15150
rect 20950 15130 20960 15150
rect 20920 14990 20960 15130
rect 20920 14970 20930 14990
rect 20950 14970 20960 14990
rect 20920 14960 20960 14970
rect 0 14910 40 14920
rect 0 14890 10 14910
rect 30 14890 40 14910
rect 0 14750 40 14890
rect 0 14730 10 14750
rect 30 14730 40 14750
rect 0 14720 40 14730
rect 80 14910 120 14920
rect 80 14890 90 14910
rect 110 14890 120 14910
rect 80 14750 120 14890
rect 80 14730 90 14750
rect 110 14730 120 14750
rect 80 14720 120 14730
rect 160 14910 200 14920
rect 160 14890 170 14910
rect 190 14890 200 14910
rect 160 14750 200 14890
rect 160 14730 170 14750
rect 190 14730 200 14750
rect 160 14720 200 14730
rect 240 14910 280 14920
rect 240 14890 250 14910
rect 270 14890 280 14910
rect 240 14750 280 14890
rect 240 14730 250 14750
rect 270 14730 280 14750
rect 240 14720 280 14730
rect 320 14910 360 14920
rect 320 14890 330 14910
rect 350 14890 360 14910
rect 320 14750 360 14890
rect 320 14730 330 14750
rect 350 14730 360 14750
rect 320 14720 360 14730
rect 400 14910 440 14920
rect 400 14890 410 14910
rect 430 14890 440 14910
rect 400 14750 440 14890
rect 400 14730 410 14750
rect 430 14730 440 14750
rect 400 14720 440 14730
rect 480 14910 520 14920
rect 480 14890 490 14910
rect 510 14890 520 14910
rect 480 14750 520 14890
rect 480 14730 490 14750
rect 510 14730 520 14750
rect 480 14720 520 14730
rect 560 14910 600 14920
rect 560 14890 570 14910
rect 590 14890 600 14910
rect 560 14750 600 14890
rect 560 14730 570 14750
rect 590 14730 600 14750
rect 560 14720 600 14730
rect 640 14910 680 14920
rect 640 14890 650 14910
rect 670 14890 680 14910
rect 640 14750 680 14890
rect 640 14730 650 14750
rect 670 14730 680 14750
rect 640 14720 680 14730
rect 720 14910 760 14920
rect 720 14890 730 14910
rect 750 14890 760 14910
rect 720 14750 760 14890
rect 720 14730 730 14750
rect 750 14730 760 14750
rect 720 14720 760 14730
rect 800 14910 840 14920
rect 800 14890 810 14910
rect 830 14890 840 14910
rect 800 14750 840 14890
rect 800 14730 810 14750
rect 830 14730 840 14750
rect 800 14720 840 14730
rect 880 14910 920 14920
rect 880 14890 890 14910
rect 910 14890 920 14910
rect 880 14750 920 14890
rect 880 14730 890 14750
rect 910 14730 920 14750
rect 880 14720 920 14730
rect 960 14910 1000 14920
rect 960 14890 970 14910
rect 990 14890 1000 14910
rect 960 14750 1000 14890
rect 960 14730 970 14750
rect 990 14730 1000 14750
rect 960 14720 1000 14730
rect 1040 14910 1080 14920
rect 1040 14890 1050 14910
rect 1070 14890 1080 14910
rect 1040 14750 1080 14890
rect 1040 14730 1050 14750
rect 1070 14730 1080 14750
rect 1040 14720 1080 14730
rect 1120 14910 1160 14920
rect 1120 14890 1130 14910
rect 1150 14890 1160 14910
rect 1120 14750 1160 14890
rect 1120 14730 1130 14750
rect 1150 14730 1160 14750
rect 1120 14720 1160 14730
rect 1200 14910 1240 14920
rect 1200 14890 1210 14910
rect 1230 14890 1240 14910
rect 1200 14750 1240 14890
rect 1200 14730 1210 14750
rect 1230 14730 1240 14750
rect 1200 14720 1240 14730
rect 1280 14910 1320 14920
rect 1280 14890 1290 14910
rect 1310 14890 1320 14910
rect 1280 14750 1320 14890
rect 1280 14730 1290 14750
rect 1310 14730 1320 14750
rect 1280 14720 1320 14730
rect 1360 14910 1400 14920
rect 1360 14890 1370 14910
rect 1390 14890 1400 14910
rect 1360 14750 1400 14890
rect 1360 14730 1370 14750
rect 1390 14730 1400 14750
rect 1360 14720 1400 14730
rect 1440 14910 1480 14920
rect 1440 14890 1450 14910
rect 1470 14890 1480 14910
rect 1440 14750 1480 14890
rect 1440 14730 1450 14750
rect 1470 14730 1480 14750
rect 1440 14720 1480 14730
rect 1520 14910 1560 14920
rect 1520 14890 1530 14910
rect 1550 14890 1560 14910
rect 1520 14750 1560 14890
rect 1520 14730 1530 14750
rect 1550 14730 1560 14750
rect 1520 14720 1560 14730
rect 1600 14910 1640 14920
rect 1600 14890 1610 14910
rect 1630 14890 1640 14910
rect 1600 14750 1640 14890
rect 1600 14730 1610 14750
rect 1630 14730 1640 14750
rect 1600 14720 1640 14730
rect 1680 14910 1720 14920
rect 1680 14890 1690 14910
rect 1710 14890 1720 14910
rect 1680 14750 1720 14890
rect 1680 14730 1690 14750
rect 1710 14730 1720 14750
rect 1680 14720 1720 14730
rect 1760 14910 1800 14920
rect 1760 14890 1770 14910
rect 1790 14890 1800 14910
rect 1760 14750 1800 14890
rect 1760 14730 1770 14750
rect 1790 14730 1800 14750
rect 1760 14720 1800 14730
rect 1840 14910 1880 14920
rect 1840 14890 1850 14910
rect 1870 14890 1880 14910
rect 1840 14750 1880 14890
rect 1840 14730 1850 14750
rect 1870 14730 1880 14750
rect 1840 14720 1880 14730
rect 1920 14910 1960 14920
rect 1920 14890 1930 14910
rect 1950 14890 1960 14910
rect 1920 14750 1960 14890
rect 1920 14730 1930 14750
rect 1950 14730 1960 14750
rect 1920 14720 1960 14730
rect 2000 14910 2040 14920
rect 2000 14890 2010 14910
rect 2030 14890 2040 14910
rect 2000 14750 2040 14890
rect 2000 14730 2010 14750
rect 2030 14730 2040 14750
rect 2000 14720 2040 14730
rect 2080 14910 2120 14920
rect 2080 14890 2090 14910
rect 2110 14890 2120 14910
rect 2080 14750 2120 14890
rect 2080 14730 2090 14750
rect 2110 14730 2120 14750
rect 2080 14720 2120 14730
rect 2160 14910 2200 14920
rect 2160 14890 2170 14910
rect 2190 14890 2200 14910
rect 2160 14750 2200 14890
rect 2160 14730 2170 14750
rect 2190 14730 2200 14750
rect 2160 14720 2200 14730
rect 2240 14910 2280 14920
rect 2240 14890 2250 14910
rect 2270 14890 2280 14910
rect 2240 14750 2280 14890
rect 2240 14730 2250 14750
rect 2270 14730 2280 14750
rect 2240 14720 2280 14730
rect 2320 14910 2360 14920
rect 2320 14890 2330 14910
rect 2350 14890 2360 14910
rect 2320 14750 2360 14890
rect 2320 14730 2330 14750
rect 2350 14730 2360 14750
rect 2320 14720 2360 14730
rect 2400 14910 2440 14920
rect 2400 14890 2410 14910
rect 2430 14890 2440 14910
rect 2400 14750 2440 14890
rect 2400 14730 2410 14750
rect 2430 14730 2440 14750
rect 2400 14720 2440 14730
rect 2480 14910 2520 14920
rect 2480 14890 2490 14910
rect 2510 14890 2520 14910
rect 2480 14750 2520 14890
rect 2480 14730 2490 14750
rect 2510 14730 2520 14750
rect 2480 14720 2520 14730
rect 2560 14910 2600 14920
rect 2560 14890 2570 14910
rect 2590 14890 2600 14910
rect 2560 14750 2600 14890
rect 2560 14730 2570 14750
rect 2590 14730 2600 14750
rect 2560 14720 2600 14730
rect 2640 14910 2680 14920
rect 2640 14890 2650 14910
rect 2670 14890 2680 14910
rect 2640 14750 2680 14890
rect 2640 14730 2650 14750
rect 2670 14730 2680 14750
rect 2640 14720 2680 14730
rect 2720 14910 2760 14920
rect 2720 14890 2730 14910
rect 2750 14890 2760 14910
rect 2720 14750 2760 14890
rect 2720 14730 2730 14750
rect 2750 14730 2760 14750
rect 2720 14720 2760 14730
rect 2800 14910 2840 14920
rect 2800 14890 2810 14910
rect 2830 14890 2840 14910
rect 2800 14750 2840 14890
rect 2800 14730 2810 14750
rect 2830 14730 2840 14750
rect 2800 14720 2840 14730
rect 2880 14910 2920 14920
rect 2880 14890 2890 14910
rect 2910 14890 2920 14910
rect 2880 14750 2920 14890
rect 2880 14730 2890 14750
rect 2910 14730 2920 14750
rect 2880 14720 2920 14730
rect 2960 14910 3000 14920
rect 2960 14890 2970 14910
rect 2990 14890 3000 14910
rect 2960 14750 3000 14890
rect 2960 14730 2970 14750
rect 2990 14730 3000 14750
rect 2960 14720 3000 14730
rect 3040 14910 3080 14920
rect 3040 14890 3050 14910
rect 3070 14890 3080 14910
rect 3040 14750 3080 14890
rect 3040 14730 3050 14750
rect 3070 14730 3080 14750
rect 3040 14720 3080 14730
rect 3120 14910 3160 14920
rect 3120 14890 3130 14910
rect 3150 14890 3160 14910
rect 3120 14750 3160 14890
rect 3120 14730 3130 14750
rect 3150 14730 3160 14750
rect 3120 14720 3160 14730
rect 3200 14910 3240 14920
rect 3200 14890 3210 14910
rect 3230 14890 3240 14910
rect 3200 14750 3240 14890
rect 3200 14730 3210 14750
rect 3230 14730 3240 14750
rect 3200 14720 3240 14730
rect 3280 14910 3320 14920
rect 3280 14890 3290 14910
rect 3310 14890 3320 14910
rect 3280 14750 3320 14890
rect 3280 14730 3290 14750
rect 3310 14730 3320 14750
rect 3280 14720 3320 14730
rect 3360 14910 3400 14920
rect 3360 14890 3370 14910
rect 3390 14890 3400 14910
rect 3360 14750 3400 14890
rect 3360 14730 3370 14750
rect 3390 14730 3400 14750
rect 3360 14720 3400 14730
rect 3440 14910 3480 14920
rect 3440 14890 3450 14910
rect 3470 14890 3480 14910
rect 3440 14750 3480 14890
rect 3440 14730 3450 14750
rect 3470 14730 3480 14750
rect 3440 14720 3480 14730
rect 3520 14910 3560 14920
rect 3520 14890 3530 14910
rect 3550 14890 3560 14910
rect 3520 14750 3560 14890
rect 3520 14730 3530 14750
rect 3550 14730 3560 14750
rect 3520 14720 3560 14730
rect 3600 14910 3640 14920
rect 3600 14890 3610 14910
rect 3630 14890 3640 14910
rect 3600 14750 3640 14890
rect 3600 14730 3610 14750
rect 3630 14730 3640 14750
rect 3600 14720 3640 14730
rect 3680 14910 3720 14920
rect 3680 14890 3690 14910
rect 3710 14890 3720 14910
rect 3680 14750 3720 14890
rect 3680 14730 3690 14750
rect 3710 14730 3720 14750
rect 3680 14720 3720 14730
rect 3760 14910 3800 14920
rect 3760 14890 3770 14910
rect 3790 14890 3800 14910
rect 3760 14750 3800 14890
rect 3760 14730 3770 14750
rect 3790 14730 3800 14750
rect 3760 14720 3800 14730
rect 3840 14910 3880 14920
rect 3840 14890 3850 14910
rect 3870 14890 3880 14910
rect 3840 14750 3880 14890
rect 3840 14730 3850 14750
rect 3870 14730 3880 14750
rect 3840 14720 3880 14730
rect 3920 14910 3960 14920
rect 3920 14890 3930 14910
rect 3950 14890 3960 14910
rect 3920 14750 3960 14890
rect 3920 14730 3930 14750
rect 3950 14730 3960 14750
rect 3920 14720 3960 14730
rect 4000 14910 4040 14920
rect 4000 14890 4010 14910
rect 4030 14890 4040 14910
rect 4000 14750 4040 14890
rect 4000 14730 4010 14750
rect 4030 14730 4040 14750
rect 4000 14720 4040 14730
rect 4080 14910 4120 14920
rect 4080 14890 4090 14910
rect 4110 14890 4120 14910
rect 4080 14750 4120 14890
rect 4080 14730 4090 14750
rect 4110 14730 4120 14750
rect 4080 14720 4120 14730
rect 4160 14910 4200 14920
rect 4160 14890 4170 14910
rect 4190 14890 4200 14910
rect 4160 14750 4200 14890
rect 4160 14730 4170 14750
rect 4190 14730 4200 14750
rect 4160 14720 4200 14730
rect 4240 14720 4280 14920
rect 4320 14720 4360 14920
rect 4400 14720 4440 14920
rect 4480 14720 4520 14920
rect 4560 14720 4600 14920
rect 4640 14720 4680 14920
rect 4720 14720 4760 14920
rect 4800 14720 4840 14920
rect 4880 14720 4920 14920
rect 4960 14720 5000 14920
rect 5040 14720 5080 14920
rect 5120 14720 5160 14920
rect 5200 14720 5240 14920
rect 5280 14720 5320 14920
rect 5360 14720 5400 14920
rect 5440 14720 5480 14920
rect 5520 14720 5560 14920
rect 5600 14720 5640 14920
rect 5680 14720 5720 14920
rect 5760 14720 5800 14920
rect 5840 14720 5880 14920
rect 5920 14720 5960 14920
rect 6000 14720 6040 14920
rect 6080 14720 6120 14920
rect 6160 14720 6200 14920
rect 6240 14910 6280 14920
rect 6240 14890 6250 14910
rect 6270 14890 6280 14910
rect 6240 14750 6280 14890
rect 6240 14730 6250 14750
rect 6270 14730 6280 14750
rect 6240 14720 6280 14730
rect 6320 14910 6360 14920
rect 6320 14890 6330 14910
rect 6350 14890 6360 14910
rect 6320 14750 6360 14890
rect 6320 14730 6330 14750
rect 6350 14730 6360 14750
rect 6320 14720 6360 14730
rect 6400 14910 6440 14920
rect 6400 14890 6410 14910
rect 6430 14890 6440 14910
rect 6400 14750 6440 14890
rect 6400 14730 6410 14750
rect 6430 14730 6440 14750
rect 6400 14720 6440 14730
rect 6480 14910 6520 14920
rect 6480 14890 6490 14910
rect 6510 14890 6520 14910
rect 6480 14750 6520 14890
rect 6480 14730 6490 14750
rect 6510 14730 6520 14750
rect 6480 14720 6520 14730
rect 6560 14910 6600 14920
rect 6560 14890 6570 14910
rect 6590 14890 6600 14910
rect 6560 14750 6600 14890
rect 6560 14730 6570 14750
rect 6590 14730 6600 14750
rect 6560 14720 6600 14730
rect 6640 14910 6680 14920
rect 6640 14890 6650 14910
rect 6670 14890 6680 14910
rect 6640 14750 6680 14890
rect 6640 14730 6650 14750
rect 6670 14730 6680 14750
rect 6640 14720 6680 14730
rect 6720 14910 6760 14920
rect 6720 14890 6730 14910
rect 6750 14890 6760 14910
rect 6720 14750 6760 14890
rect 6720 14730 6730 14750
rect 6750 14730 6760 14750
rect 6720 14720 6760 14730
rect 6800 14910 6840 14920
rect 6800 14890 6810 14910
rect 6830 14890 6840 14910
rect 6800 14750 6840 14890
rect 6800 14730 6810 14750
rect 6830 14730 6840 14750
rect 6800 14720 6840 14730
rect 6880 14910 6920 14920
rect 6880 14890 6890 14910
rect 6910 14890 6920 14910
rect 6880 14750 6920 14890
rect 6880 14730 6890 14750
rect 6910 14730 6920 14750
rect 6880 14720 6920 14730
rect 6960 14910 7000 14920
rect 6960 14890 6970 14910
rect 6990 14890 7000 14910
rect 6960 14750 7000 14890
rect 6960 14730 6970 14750
rect 6990 14730 7000 14750
rect 6960 14720 7000 14730
rect 7040 14910 7080 14920
rect 7040 14890 7050 14910
rect 7070 14890 7080 14910
rect 7040 14750 7080 14890
rect 7040 14730 7050 14750
rect 7070 14730 7080 14750
rect 7040 14720 7080 14730
rect 7120 14910 7160 14920
rect 7120 14890 7130 14910
rect 7150 14890 7160 14910
rect 7120 14750 7160 14890
rect 7120 14730 7130 14750
rect 7150 14730 7160 14750
rect 7120 14720 7160 14730
rect 7200 14910 7240 14920
rect 7200 14890 7210 14910
rect 7230 14890 7240 14910
rect 7200 14750 7240 14890
rect 7200 14730 7210 14750
rect 7230 14730 7240 14750
rect 7200 14720 7240 14730
rect 7280 14910 7320 14920
rect 7280 14890 7290 14910
rect 7310 14890 7320 14910
rect 7280 14750 7320 14890
rect 7280 14730 7290 14750
rect 7310 14730 7320 14750
rect 7280 14720 7320 14730
rect 7360 14910 7400 14920
rect 7360 14890 7370 14910
rect 7390 14890 7400 14910
rect 7360 14750 7400 14890
rect 7360 14730 7370 14750
rect 7390 14730 7400 14750
rect 7360 14720 7400 14730
rect 7440 14910 7480 14920
rect 7440 14890 7450 14910
rect 7470 14890 7480 14910
rect 7440 14750 7480 14890
rect 7440 14730 7450 14750
rect 7470 14730 7480 14750
rect 7440 14720 7480 14730
rect 7520 14910 7560 14920
rect 7520 14890 7530 14910
rect 7550 14890 7560 14910
rect 7520 14750 7560 14890
rect 7520 14730 7530 14750
rect 7550 14730 7560 14750
rect 7520 14720 7560 14730
rect 7600 14910 7640 14920
rect 7600 14890 7610 14910
rect 7630 14890 7640 14910
rect 7600 14750 7640 14890
rect 7600 14730 7610 14750
rect 7630 14730 7640 14750
rect 7600 14720 7640 14730
rect 7680 14910 7720 14920
rect 7680 14890 7690 14910
rect 7710 14890 7720 14910
rect 7680 14750 7720 14890
rect 7680 14730 7690 14750
rect 7710 14730 7720 14750
rect 7680 14720 7720 14730
rect 7760 14910 7800 14920
rect 7760 14890 7770 14910
rect 7790 14890 7800 14910
rect 7760 14750 7800 14890
rect 7760 14730 7770 14750
rect 7790 14730 7800 14750
rect 7760 14720 7800 14730
rect 7840 14910 7880 14920
rect 7840 14890 7850 14910
rect 7870 14890 7880 14910
rect 7840 14750 7880 14890
rect 7840 14730 7850 14750
rect 7870 14730 7880 14750
rect 7840 14720 7880 14730
rect 7920 14910 7960 14920
rect 7920 14890 7930 14910
rect 7950 14890 7960 14910
rect 7920 14750 7960 14890
rect 7920 14730 7930 14750
rect 7950 14730 7960 14750
rect 7920 14720 7960 14730
rect 8000 14910 8040 14920
rect 8000 14890 8010 14910
rect 8030 14890 8040 14910
rect 8000 14750 8040 14890
rect 8000 14730 8010 14750
rect 8030 14730 8040 14750
rect 8000 14720 8040 14730
rect 8080 14910 8120 14920
rect 8080 14890 8090 14910
rect 8110 14890 8120 14910
rect 8080 14750 8120 14890
rect 8080 14730 8090 14750
rect 8110 14730 8120 14750
rect 8080 14720 8120 14730
rect 8160 14910 8200 14920
rect 8160 14890 8170 14910
rect 8190 14890 8200 14910
rect 8160 14750 8200 14890
rect 8160 14730 8170 14750
rect 8190 14730 8200 14750
rect 8160 14720 8200 14730
rect 8240 14910 8280 14920
rect 8240 14890 8250 14910
rect 8270 14890 8280 14910
rect 8240 14750 8280 14890
rect 8240 14730 8250 14750
rect 8270 14730 8280 14750
rect 8240 14720 8280 14730
rect 8320 14910 8360 14920
rect 8320 14890 8330 14910
rect 8350 14890 8360 14910
rect 8320 14750 8360 14890
rect 8320 14730 8330 14750
rect 8350 14730 8360 14750
rect 8320 14720 8360 14730
rect 8400 14910 8440 14920
rect 8400 14890 8410 14910
rect 8430 14890 8440 14910
rect 8400 14750 8440 14890
rect 8400 14730 8410 14750
rect 8430 14730 8440 14750
rect 8400 14720 8440 14730
rect 8480 14910 8520 14920
rect 8480 14890 8490 14910
rect 8510 14890 8520 14910
rect 8480 14750 8520 14890
rect 8480 14730 8490 14750
rect 8510 14730 8520 14750
rect 8480 14720 8520 14730
rect 8560 14910 8600 14920
rect 8560 14890 8570 14910
rect 8590 14890 8600 14910
rect 8560 14750 8600 14890
rect 8560 14730 8570 14750
rect 8590 14730 8600 14750
rect 8560 14720 8600 14730
rect 8640 14910 8680 14920
rect 8640 14890 8650 14910
rect 8670 14890 8680 14910
rect 8640 14750 8680 14890
rect 8640 14730 8650 14750
rect 8670 14730 8680 14750
rect 8640 14720 8680 14730
rect 8720 14910 8760 14920
rect 8720 14890 8730 14910
rect 8750 14890 8760 14910
rect 8720 14750 8760 14890
rect 8720 14730 8730 14750
rect 8750 14730 8760 14750
rect 8720 14720 8760 14730
rect 8800 14910 8840 14920
rect 8800 14890 8810 14910
rect 8830 14890 8840 14910
rect 8800 14750 8840 14890
rect 8800 14730 8810 14750
rect 8830 14730 8840 14750
rect 8800 14720 8840 14730
rect 8880 14910 8920 14920
rect 8880 14890 8890 14910
rect 8910 14890 8920 14910
rect 8880 14750 8920 14890
rect 8880 14730 8890 14750
rect 8910 14730 8920 14750
rect 8880 14720 8920 14730
rect 8960 14910 9000 14920
rect 8960 14890 8970 14910
rect 8990 14890 9000 14910
rect 8960 14750 9000 14890
rect 8960 14730 8970 14750
rect 8990 14730 9000 14750
rect 8960 14720 9000 14730
rect 9040 14910 9080 14920
rect 9040 14890 9050 14910
rect 9070 14890 9080 14910
rect 9040 14750 9080 14890
rect 9040 14730 9050 14750
rect 9070 14730 9080 14750
rect 9040 14720 9080 14730
rect 9120 14910 9160 14920
rect 9120 14890 9130 14910
rect 9150 14890 9160 14910
rect 9120 14750 9160 14890
rect 9120 14730 9130 14750
rect 9150 14730 9160 14750
rect 9120 14720 9160 14730
rect 9200 14910 9240 14920
rect 9200 14890 9210 14910
rect 9230 14890 9240 14910
rect 9200 14750 9240 14890
rect 9200 14730 9210 14750
rect 9230 14730 9240 14750
rect 9200 14720 9240 14730
rect 9280 14910 9320 14920
rect 9280 14890 9290 14910
rect 9310 14890 9320 14910
rect 9280 14750 9320 14890
rect 9280 14730 9290 14750
rect 9310 14730 9320 14750
rect 9280 14720 9320 14730
rect 9360 14910 9400 14920
rect 9360 14890 9370 14910
rect 9390 14890 9400 14910
rect 9360 14750 9400 14890
rect 9360 14730 9370 14750
rect 9390 14730 9400 14750
rect 9360 14720 9400 14730
rect 9440 14910 9480 14920
rect 9440 14890 9450 14910
rect 9470 14890 9480 14910
rect 9440 14750 9480 14890
rect 9440 14730 9450 14750
rect 9470 14730 9480 14750
rect 9440 14720 9480 14730
rect 9520 14720 9560 14920
rect 9600 14720 9640 14920
rect 9680 14720 9720 14920
rect 9760 14720 9800 14920
rect 9840 14720 9880 14920
rect 9920 14720 9960 14920
rect 10000 14720 10040 14920
rect 10080 14720 10120 14920
rect 10160 14720 10200 14920
rect 10240 14720 10280 14920
rect 10320 14720 10360 14920
rect 10400 14720 10440 14920
rect 10480 14720 10520 14920
rect 10560 14720 10600 14920
rect 10640 14720 10680 14920
rect 10720 14720 10760 14920
rect 10800 14720 10840 14920
rect 10880 14720 10920 14920
rect 10960 14720 11000 14920
rect 11040 14720 11080 14920
rect 11120 14720 11160 14920
rect 11200 14720 11240 14920
rect 11280 14720 11320 14920
rect 11360 14720 11400 14920
rect 11440 14720 11480 14920
rect 11560 14910 11600 14920
rect 11560 14890 11570 14910
rect 11590 14890 11600 14910
rect 11560 14750 11600 14890
rect 11560 14730 11570 14750
rect 11590 14730 11600 14750
rect 11560 14720 11600 14730
rect 11640 14910 11680 14920
rect 11640 14890 11650 14910
rect 11670 14890 11680 14910
rect 11640 14750 11680 14890
rect 11640 14730 11650 14750
rect 11670 14730 11680 14750
rect 11640 14720 11680 14730
rect 11720 14910 11760 14920
rect 11720 14890 11730 14910
rect 11750 14890 11760 14910
rect 11720 14750 11760 14890
rect 11720 14730 11730 14750
rect 11750 14730 11760 14750
rect 11720 14720 11760 14730
rect 11800 14910 11840 14920
rect 11800 14890 11810 14910
rect 11830 14890 11840 14910
rect 11800 14750 11840 14890
rect 11800 14730 11810 14750
rect 11830 14730 11840 14750
rect 11800 14720 11840 14730
rect 11880 14910 11920 14920
rect 11880 14890 11890 14910
rect 11910 14890 11920 14910
rect 11880 14750 11920 14890
rect 11880 14730 11890 14750
rect 11910 14730 11920 14750
rect 11880 14720 11920 14730
rect 11960 14910 12000 14920
rect 11960 14890 11970 14910
rect 11990 14890 12000 14910
rect 11960 14750 12000 14890
rect 11960 14730 11970 14750
rect 11990 14730 12000 14750
rect 11960 14720 12000 14730
rect 12040 14910 12080 14920
rect 12040 14890 12050 14910
rect 12070 14890 12080 14910
rect 12040 14750 12080 14890
rect 12040 14730 12050 14750
rect 12070 14730 12080 14750
rect 12040 14720 12080 14730
rect 12120 14910 12160 14920
rect 12120 14890 12130 14910
rect 12150 14890 12160 14910
rect 12120 14750 12160 14890
rect 12120 14730 12130 14750
rect 12150 14730 12160 14750
rect 12120 14720 12160 14730
rect 12200 14910 12240 14920
rect 12200 14890 12210 14910
rect 12230 14890 12240 14910
rect 12200 14750 12240 14890
rect 12200 14730 12210 14750
rect 12230 14730 12240 14750
rect 12200 14720 12240 14730
rect 12280 14910 12320 14920
rect 12280 14890 12290 14910
rect 12310 14890 12320 14910
rect 12280 14750 12320 14890
rect 12280 14730 12290 14750
rect 12310 14730 12320 14750
rect 12280 14720 12320 14730
rect 12360 14910 12400 14920
rect 12360 14890 12370 14910
rect 12390 14890 12400 14910
rect 12360 14750 12400 14890
rect 12360 14730 12370 14750
rect 12390 14730 12400 14750
rect 12360 14720 12400 14730
rect 12440 14910 12480 14920
rect 12440 14890 12450 14910
rect 12470 14890 12480 14910
rect 12440 14750 12480 14890
rect 12440 14730 12450 14750
rect 12470 14730 12480 14750
rect 12440 14720 12480 14730
rect 12520 14910 12560 14920
rect 12520 14890 12530 14910
rect 12550 14890 12560 14910
rect 12520 14750 12560 14890
rect 12520 14730 12530 14750
rect 12550 14730 12560 14750
rect 12520 14720 12560 14730
rect 12600 14910 12640 14920
rect 12600 14890 12610 14910
rect 12630 14890 12640 14910
rect 12600 14750 12640 14890
rect 12600 14730 12610 14750
rect 12630 14730 12640 14750
rect 12600 14720 12640 14730
rect 12680 14910 12720 14920
rect 12680 14890 12690 14910
rect 12710 14890 12720 14910
rect 12680 14750 12720 14890
rect 12680 14730 12690 14750
rect 12710 14730 12720 14750
rect 12680 14720 12720 14730
rect 12760 14910 12800 14920
rect 12760 14890 12770 14910
rect 12790 14890 12800 14910
rect 12760 14750 12800 14890
rect 12760 14730 12770 14750
rect 12790 14730 12800 14750
rect 12760 14720 12800 14730
rect 12840 14910 12880 14920
rect 12840 14890 12850 14910
rect 12870 14890 12880 14910
rect 12840 14750 12880 14890
rect 12840 14730 12850 14750
rect 12870 14730 12880 14750
rect 12840 14720 12880 14730
rect 12920 14910 12960 14920
rect 12920 14890 12930 14910
rect 12950 14890 12960 14910
rect 12920 14750 12960 14890
rect 12920 14730 12930 14750
rect 12950 14730 12960 14750
rect 12920 14720 12960 14730
rect 13000 14910 13040 14920
rect 13000 14890 13010 14910
rect 13030 14890 13040 14910
rect 13000 14750 13040 14890
rect 13000 14730 13010 14750
rect 13030 14730 13040 14750
rect 13000 14720 13040 14730
rect 13080 14910 13120 14920
rect 13080 14890 13090 14910
rect 13110 14890 13120 14910
rect 13080 14750 13120 14890
rect 13080 14730 13090 14750
rect 13110 14730 13120 14750
rect 13080 14720 13120 14730
rect 13160 14910 13200 14920
rect 13160 14890 13170 14910
rect 13190 14890 13200 14910
rect 13160 14750 13200 14890
rect 13160 14730 13170 14750
rect 13190 14730 13200 14750
rect 13160 14720 13200 14730
rect 13240 14910 13280 14920
rect 13240 14890 13250 14910
rect 13270 14890 13280 14910
rect 13240 14750 13280 14890
rect 13240 14730 13250 14750
rect 13270 14730 13280 14750
rect 13240 14720 13280 14730
rect 13320 14910 13360 14920
rect 13320 14890 13330 14910
rect 13350 14890 13360 14910
rect 13320 14750 13360 14890
rect 13320 14730 13330 14750
rect 13350 14730 13360 14750
rect 13320 14720 13360 14730
rect 13400 14910 13440 14920
rect 13400 14890 13410 14910
rect 13430 14890 13440 14910
rect 13400 14750 13440 14890
rect 13400 14730 13410 14750
rect 13430 14730 13440 14750
rect 13400 14720 13440 14730
rect 13480 14910 13520 14920
rect 13480 14890 13490 14910
rect 13510 14890 13520 14910
rect 13480 14750 13520 14890
rect 13480 14730 13490 14750
rect 13510 14730 13520 14750
rect 13480 14720 13520 14730
rect 13560 14910 13600 14920
rect 13560 14890 13570 14910
rect 13590 14890 13600 14910
rect 13560 14750 13600 14890
rect 13560 14730 13570 14750
rect 13590 14730 13600 14750
rect 13560 14720 13600 14730
rect 13640 14910 13680 14920
rect 13640 14890 13650 14910
rect 13670 14890 13680 14910
rect 13640 14750 13680 14890
rect 13640 14730 13650 14750
rect 13670 14730 13680 14750
rect 13640 14720 13680 14730
rect 13720 14910 13760 14920
rect 13720 14890 13730 14910
rect 13750 14890 13760 14910
rect 13720 14750 13760 14890
rect 13720 14730 13730 14750
rect 13750 14730 13760 14750
rect 13720 14720 13760 14730
rect 13800 14910 13840 14920
rect 13800 14890 13810 14910
rect 13830 14890 13840 14910
rect 13800 14750 13840 14890
rect 13800 14730 13810 14750
rect 13830 14730 13840 14750
rect 13800 14720 13840 14730
rect 13880 14910 13920 14920
rect 13880 14890 13890 14910
rect 13910 14890 13920 14910
rect 13880 14750 13920 14890
rect 13880 14730 13890 14750
rect 13910 14730 13920 14750
rect 13880 14720 13920 14730
rect 13960 14910 14000 14920
rect 13960 14890 13970 14910
rect 13990 14890 14000 14910
rect 13960 14750 14000 14890
rect 13960 14730 13970 14750
rect 13990 14730 14000 14750
rect 13960 14720 14000 14730
rect 14040 14910 14080 14920
rect 14040 14890 14050 14910
rect 14070 14890 14080 14910
rect 14040 14750 14080 14890
rect 14040 14730 14050 14750
rect 14070 14730 14080 14750
rect 14040 14720 14080 14730
rect 14120 14910 14160 14920
rect 14120 14890 14130 14910
rect 14150 14890 14160 14910
rect 14120 14750 14160 14890
rect 14120 14730 14130 14750
rect 14150 14730 14160 14750
rect 14120 14720 14160 14730
rect 14200 14910 14240 14920
rect 14200 14890 14210 14910
rect 14230 14890 14240 14910
rect 14200 14750 14240 14890
rect 14200 14730 14210 14750
rect 14230 14730 14240 14750
rect 14200 14720 14240 14730
rect 14280 14910 14320 14920
rect 14280 14890 14290 14910
rect 14310 14890 14320 14910
rect 14280 14750 14320 14890
rect 14280 14730 14290 14750
rect 14310 14730 14320 14750
rect 14280 14720 14320 14730
rect 14360 14910 14400 14920
rect 14360 14890 14370 14910
rect 14390 14890 14400 14910
rect 14360 14750 14400 14890
rect 14360 14730 14370 14750
rect 14390 14730 14400 14750
rect 14360 14720 14400 14730
rect 14440 14910 14480 14920
rect 14440 14890 14450 14910
rect 14470 14890 14480 14910
rect 14440 14750 14480 14890
rect 14440 14730 14450 14750
rect 14470 14730 14480 14750
rect 14440 14720 14480 14730
rect 14520 14910 14560 14920
rect 14520 14890 14530 14910
rect 14550 14890 14560 14910
rect 14520 14750 14560 14890
rect 14520 14730 14530 14750
rect 14550 14730 14560 14750
rect 14520 14720 14560 14730
rect 14600 14910 14640 14920
rect 14600 14890 14610 14910
rect 14630 14890 14640 14910
rect 14600 14750 14640 14890
rect 14600 14730 14610 14750
rect 14630 14730 14640 14750
rect 14600 14720 14640 14730
rect 14680 14910 14720 14920
rect 14680 14890 14690 14910
rect 14710 14890 14720 14910
rect 14680 14750 14720 14890
rect 14680 14730 14690 14750
rect 14710 14730 14720 14750
rect 14680 14720 14720 14730
rect 14760 14720 14800 14920
rect 14840 14720 14880 14920
rect 14920 14720 14960 14920
rect 15000 14720 15040 14920
rect 15080 14720 15120 14920
rect 15160 14720 15200 14920
rect 15240 14720 15280 14920
rect 15320 14720 15360 14920
rect 15400 14720 15440 14920
rect 15480 14720 15520 14920
rect 15560 14720 15600 14920
rect 15640 14720 15680 14920
rect 15720 14720 15760 14920
rect 15800 14720 15840 14920
rect 15880 14720 15920 14920
rect 15960 14720 16000 14920
rect 16040 14720 16080 14920
rect 16120 14720 16160 14920
rect 16200 14720 16240 14920
rect 16280 14720 16320 14920
rect 16360 14720 16400 14920
rect 16440 14720 16480 14920
rect 16520 14720 16560 14920
rect 16600 14720 16640 14920
rect 16680 14720 16720 14920
rect 16760 14910 16800 14920
rect 16760 14890 16770 14910
rect 16790 14890 16800 14910
rect 16760 14750 16800 14890
rect 16760 14730 16770 14750
rect 16790 14730 16800 14750
rect 16760 14720 16800 14730
rect 16840 14910 16880 14920
rect 16840 14890 16850 14910
rect 16870 14890 16880 14910
rect 16840 14750 16880 14890
rect 16840 14730 16850 14750
rect 16870 14730 16880 14750
rect 16840 14720 16880 14730
rect 16920 14910 16960 14920
rect 16920 14890 16930 14910
rect 16950 14890 16960 14910
rect 16920 14750 16960 14890
rect 16920 14730 16930 14750
rect 16950 14730 16960 14750
rect 16920 14720 16960 14730
rect 17000 14910 17040 14920
rect 17000 14890 17010 14910
rect 17030 14890 17040 14910
rect 17000 14750 17040 14890
rect 17000 14730 17010 14750
rect 17030 14730 17040 14750
rect 17000 14720 17040 14730
rect 17080 14910 17120 14920
rect 17080 14890 17090 14910
rect 17110 14890 17120 14910
rect 17080 14750 17120 14890
rect 17080 14730 17090 14750
rect 17110 14730 17120 14750
rect 17080 14720 17120 14730
rect 17160 14910 17200 14920
rect 17160 14890 17170 14910
rect 17190 14890 17200 14910
rect 17160 14750 17200 14890
rect 17160 14730 17170 14750
rect 17190 14730 17200 14750
rect 17160 14720 17200 14730
rect 17240 14910 17280 14920
rect 17240 14890 17250 14910
rect 17270 14890 17280 14910
rect 17240 14750 17280 14890
rect 17240 14730 17250 14750
rect 17270 14730 17280 14750
rect 17240 14720 17280 14730
rect 17320 14910 17360 14920
rect 17320 14890 17330 14910
rect 17350 14890 17360 14910
rect 17320 14750 17360 14890
rect 17320 14730 17330 14750
rect 17350 14730 17360 14750
rect 17320 14720 17360 14730
rect 17400 14910 17440 14920
rect 17400 14890 17410 14910
rect 17430 14890 17440 14910
rect 17400 14750 17440 14890
rect 17400 14730 17410 14750
rect 17430 14730 17440 14750
rect 17400 14720 17440 14730
rect 17480 14910 17520 14920
rect 17480 14890 17490 14910
rect 17510 14890 17520 14910
rect 17480 14750 17520 14890
rect 17480 14730 17490 14750
rect 17510 14730 17520 14750
rect 17480 14720 17520 14730
rect 17560 14910 17600 14920
rect 17560 14890 17570 14910
rect 17590 14890 17600 14910
rect 17560 14750 17600 14890
rect 17560 14730 17570 14750
rect 17590 14730 17600 14750
rect 17560 14720 17600 14730
rect 17640 14910 17680 14920
rect 17640 14890 17650 14910
rect 17670 14890 17680 14910
rect 17640 14750 17680 14890
rect 17640 14730 17650 14750
rect 17670 14730 17680 14750
rect 17640 14720 17680 14730
rect 17720 14910 17760 14920
rect 17720 14890 17730 14910
rect 17750 14890 17760 14910
rect 17720 14750 17760 14890
rect 17720 14730 17730 14750
rect 17750 14730 17760 14750
rect 17720 14720 17760 14730
rect 17800 14910 17840 14920
rect 17800 14890 17810 14910
rect 17830 14890 17840 14910
rect 17800 14750 17840 14890
rect 17800 14730 17810 14750
rect 17830 14730 17840 14750
rect 17800 14720 17840 14730
rect 17880 14910 17920 14920
rect 17880 14890 17890 14910
rect 17910 14890 17920 14910
rect 17880 14750 17920 14890
rect 17880 14730 17890 14750
rect 17910 14730 17920 14750
rect 17880 14720 17920 14730
rect 17960 14910 18000 14920
rect 17960 14890 17970 14910
rect 17990 14890 18000 14910
rect 17960 14750 18000 14890
rect 17960 14730 17970 14750
rect 17990 14730 18000 14750
rect 17960 14720 18000 14730
rect 18040 14910 18080 14920
rect 18040 14890 18050 14910
rect 18070 14890 18080 14910
rect 18040 14750 18080 14890
rect 18040 14730 18050 14750
rect 18070 14730 18080 14750
rect 18040 14720 18080 14730
rect 18120 14910 18160 14920
rect 18120 14890 18130 14910
rect 18150 14890 18160 14910
rect 18120 14750 18160 14890
rect 18120 14730 18130 14750
rect 18150 14730 18160 14750
rect 18120 14720 18160 14730
rect 18200 14910 18240 14920
rect 18200 14890 18210 14910
rect 18230 14890 18240 14910
rect 18200 14750 18240 14890
rect 18200 14730 18210 14750
rect 18230 14730 18240 14750
rect 18200 14720 18240 14730
rect 18280 14910 18320 14920
rect 18280 14890 18290 14910
rect 18310 14890 18320 14910
rect 18280 14750 18320 14890
rect 18280 14730 18290 14750
rect 18310 14730 18320 14750
rect 18280 14720 18320 14730
rect 18360 14910 18400 14920
rect 18360 14890 18370 14910
rect 18390 14890 18400 14910
rect 18360 14750 18400 14890
rect 18360 14730 18370 14750
rect 18390 14730 18400 14750
rect 18360 14720 18400 14730
rect 18440 14910 18480 14920
rect 18440 14890 18450 14910
rect 18470 14890 18480 14910
rect 18440 14750 18480 14890
rect 18440 14730 18450 14750
rect 18470 14730 18480 14750
rect 18440 14720 18480 14730
rect 18520 14910 18560 14920
rect 18520 14890 18530 14910
rect 18550 14890 18560 14910
rect 18520 14750 18560 14890
rect 18520 14730 18530 14750
rect 18550 14730 18560 14750
rect 18520 14720 18560 14730
rect 18600 14910 18640 14920
rect 18600 14890 18610 14910
rect 18630 14890 18640 14910
rect 18600 14750 18640 14890
rect 18600 14730 18610 14750
rect 18630 14730 18640 14750
rect 18600 14720 18640 14730
rect 18680 14910 18720 14920
rect 18680 14890 18690 14910
rect 18710 14890 18720 14910
rect 18680 14750 18720 14890
rect 18680 14730 18690 14750
rect 18710 14730 18720 14750
rect 18680 14720 18720 14730
rect 18760 14910 18800 14920
rect 18760 14890 18770 14910
rect 18790 14890 18800 14910
rect 18760 14750 18800 14890
rect 18760 14730 18770 14750
rect 18790 14730 18800 14750
rect 18760 14720 18800 14730
rect 18840 14910 18880 14920
rect 18840 14890 18850 14910
rect 18870 14890 18880 14910
rect 18840 14750 18880 14890
rect 18840 14730 18850 14750
rect 18870 14730 18880 14750
rect 18840 14720 18880 14730
rect 18920 14910 18960 14920
rect 18920 14890 18930 14910
rect 18950 14890 18960 14910
rect 18920 14750 18960 14890
rect 18920 14730 18930 14750
rect 18950 14730 18960 14750
rect 18920 14720 18960 14730
rect 19000 14910 19040 14920
rect 19000 14890 19010 14910
rect 19030 14890 19040 14910
rect 19000 14750 19040 14890
rect 19000 14730 19010 14750
rect 19030 14730 19040 14750
rect 19000 14720 19040 14730
rect 19080 14910 19120 14920
rect 19080 14890 19090 14910
rect 19110 14890 19120 14910
rect 19080 14750 19120 14890
rect 19080 14730 19090 14750
rect 19110 14730 19120 14750
rect 19080 14720 19120 14730
rect 19160 14910 19200 14920
rect 19160 14890 19170 14910
rect 19190 14890 19200 14910
rect 19160 14750 19200 14890
rect 19160 14730 19170 14750
rect 19190 14730 19200 14750
rect 19160 14720 19200 14730
rect 19240 14910 19280 14920
rect 19240 14890 19250 14910
rect 19270 14890 19280 14910
rect 19240 14750 19280 14890
rect 19240 14730 19250 14750
rect 19270 14730 19280 14750
rect 19240 14720 19280 14730
rect 19320 14910 19360 14920
rect 19320 14890 19330 14910
rect 19350 14890 19360 14910
rect 19320 14750 19360 14890
rect 19320 14730 19330 14750
rect 19350 14730 19360 14750
rect 19320 14720 19360 14730
rect 19400 14910 19440 14920
rect 19400 14890 19410 14910
rect 19430 14890 19440 14910
rect 19400 14750 19440 14890
rect 19400 14730 19410 14750
rect 19430 14730 19440 14750
rect 19400 14720 19440 14730
rect 19480 14910 19520 14920
rect 19480 14890 19490 14910
rect 19510 14890 19520 14910
rect 19480 14750 19520 14890
rect 19480 14730 19490 14750
rect 19510 14730 19520 14750
rect 19480 14720 19520 14730
rect 19560 14910 19600 14920
rect 19560 14890 19570 14910
rect 19590 14890 19600 14910
rect 19560 14750 19600 14890
rect 19560 14730 19570 14750
rect 19590 14730 19600 14750
rect 19560 14720 19600 14730
rect 19640 14910 19680 14920
rect 19640 14890 19650 14910
rect 19670 14890 19680 14910
rect 19640 14750 19680 14890
rect 19640 14730 19650 14750
rect 19670 14730 19680 14750
rect 19640 14720 19680 14730
rect 19720 14910 19760 14920
rect 19720 14890 19730 14910
rect 19750 14890 19760 14910
rect 19720 14750 19760 14890
rect 19720 14730 19730 14750
rect 19750 14730 19760 14750
rect 19720 14720 19760 14730
rect 19800 14910 19840 14920
rect 19800 14890 19810 14910
rect 19830 14890 19840 14910
rect 19800 14750 19840 14890
rect 19800 14730 19810 14750
rect 19830 14730 19840 14750
rect 19800 14720 19840 14730
rect 19880 14910 19920 14920
rect 19880 14890 19890 14910
rect 19910 14890 19920 14910
rect 19880 14750 19920 14890
rect 19880 14730 19890 14750
rect 19910 14730 19920 14750
rect 19880 14720 19920 14730
rect 19960 14910 20000 14920
rect 19960 14890 19970 14910
rect 19990 14890 20000 14910
rect 19960 14750 20000 14890
rect 19960 14730 19970 14750
rect 19990 14730 20000 14750
rect 19960 14720 20000 14730
rect 20040 14910 20080 14920
rect 20040 14890 20050 14910
rect 20070 14890 20080 14910
rect 20040 14750 20080 14890
rect 20040 14730 20050 14750
rect 20070 14730 20080 14750
rect 20040 14720 20080 14730
rect 20120 14910 20160 14920
rect 20120 14890 20130 14910
rect 20150 14890 20160 14910
rect 20120 14750 20160 14890
rect 20120 14730 20130 14750
rect 20150 14730 20160 14750
rect 20120 14720 20160 14730
rect 20200 14910 20240 14920
rect 20200 14890 20210 14910
rect 20230 14890 20240 14910
rect 20200 14750 20240 14890
rect 20200 14730 20210 14750
rect 20230 14730 20240 14750
rect 20200 14720 20240 14730
rect 20280 14910 20320 14920
rect 20280 14890 20290 14910
rect 20310 14890 20320 14910
rect 20280 14750 20320 14890
rect 20280 14730 20290 14750
rect 20310 14730 20320 14750
rect 20280 14720 20320 14730
rect 20360 14910 20400 14920
rect 20360 14890 20370 14910
rect 20390 14890 20400 14910
rect 20360 14750 20400 14890
rect 20360 14730 20370 14750
rect 20390 14730 20400 14750
rect 20360 14720 20400 14730
rect 20440 14910 20480 14920
rect 20440 14890 20450 14910
rect 20470 14890 20480 14910
rect 20440 14750 20480 14890
rect 20440 14730 20450 14750
rect 20470 14730 20480 14750
rect 20440 14720 20480 14730
rect 20520 14910 20560 14920
rect 20520 14890 20530 14910
rect 20550 14890 20560 14910
rect 20520 14750 20560 14890
rect 20520 14730 20530 14750
rect 20550 14730 20560 14750
rect 20520 14720 20560 14730
rect 20600 14910 20640 14920
rect 20600 14890 20610 14910
rect 20630 14890 20640 14910
rect 20600 14750 20640 14890
rect 20600 14730 20610 14750
rect 20630 14730 20640 14750
rect 20600 14720 20640 14730
rect 20680 14910 20720 14920
rect 20680 14890 20690 14910
rect 20710 14890 20720 14910
rect 20680 14750 20720 14890
rect 20680 14730 20690 14750
rect 20710 14730 20720 14750
rect 20680 14720 20720 14730
rect 20760 14910 20800 14920
rect 20760 14890 20770 14910
rect 20790 14890 20800 14910
rect 20760 14750 20800 14890
rect 20760 14730 20770 14750
rect 20790 14730 20800 14750
rect 20760 14720 20800 14730
rect 20840 14910 20880 14920
rect 20840 14890 20850 14910
rect 20870 14890 20880 14910
rect 20840 14750 20880 14890
rect 20840 14730 20850 14750
rect 20870 14730 20880 14750
rect 20840 14720 20880 14730
rect 20920 14910 20960 14920
rect 20920 14890 20930 14910
rect 20950 14890 20960 14910
rect 20920 14750 20960 14890
rect 20920 14730 20930 14750
rect 20950 14730 20960 14750
rect 20920 14720 20960 14730
<< viali >>
rect 10 18650 30 18670
rect 10 18490 30 18510
rect 90 18650 110 18670
rect 90 18490 110 18510
rect 170 18650 190 18670
rect 170 18490 190 18510
rect 250 18650 270 18670
rect 250 18490 270 18510
rect 330 18650 350 18670
rect 330 18490 350 18510
rect 410 18650 430 18670
rect 410 18490 430 18510
rect 490 18650 510 18670
rect 490 18490 510 18510
rect 570 18650 590 18670
rect 570 18490 590 18510
rect 650 18650 670 18670
rect 650 18490 670 18510
rect 730 18650 750 18670
rect 730 18490 750 18510
rect 810 18650 830 18670
rect 810 18490 830 18510
rect 890 18650 910 18670
rect 890 18490 910 18510
rect 970 18650 990 18670
rect 970 18490 990 18510
rect 1050 18650 1070 18670
rect 1050 18490 1070 18510
rect 1130 18650 1150 18670
rect 1130 18490 1150 18510
rect 1210 18650 1230 18670
rect 1210 18490 1230 18510
rect 1290 18650 1310 18670
rect 1290 18490 1310 18510
rect 1370 18650 1390 18670
rect 1370 18490 1390 18510
rect 1450 18650 1470 18670
rect 1450 18490 1470 18510
rect 1530 18650 1550 18670
rect 1530 18490 1550 18510
rect 1610 18650 1630 18670
rect 1610 18490 1630 18510
rect 1690 18650 1710 18670
rect 1690 18490 1710 18510
rect 1770 18650 1790 18670
rect 1770 18490 1790 18510
rect 1850 18650 1870 18670
rect 1850 18490 1870 18510
rect 1930 18650 1950 18670
rect 1930 18490 1950 18510
rect 2010 18650 2030 18670
rect 2010 18490 2030 18510
rect 2090 18650 2110 18670
rect 2090 18490 2110 18510
rect 2170 18650 2190 18670
rect 2170 18490 2190 18510
rect 2250 18650 2270 18670
rect 2250 18490 2270 18510
rect 2330 18650 2350 18670
rect 2330 18490 2350 18510
rect 2410 18650 2430 18670
rect 2410 18490 2430 18510
rect 2490 18650 2510 18670
rect 2490 18490 2510 18510
rect 2570 18650 2590 18670
rect 2570 18490 2590 18510
rect 2650 18650 2670 18670
rect 2650 18490 2670 18510
rect 2730 18650 2750 18670
rect 2730 18490 2750 18510
rect 2810 18650 2830 18670
rect 2810 18490 2830 18510
rect 2890 18650 2910 18670
rect 2890 18490 2910 18510
rect 2970 18650 2990 18670
rect 2970 18490 2990 18510
rect 3050 18650 3070 18670
rect 3050 18490 3070 18510
rect 3130 18650 3150 18670
rect 3130 18490 3150 18510
rect 3210 18650 3230 18670
rect 3210 18490 3230 18510
rect 3290 18650 3310 18670
rect 3290 18490 3310 18510
rect 3370 18650 3390 18670
rect 3370 18490 3390 18510
rect 3450 18650 3470 18670
rect 3450 18490 3470 18510
rect 3530 18650 3550 18670
rect 3530 18490 3550 18510
rect 3610 18650 3630 18670
rect 3610 18490 3630 18510
rect 3690 18650 3710 18670
rect 3690 18490 3710 18510
rect 3770 18650 3790 18670
rect 3770 18490 3790 18510
rect 3850 18650 3870 18670
rect 3850 18490 3870 18510
rect 3930 18650 3950 18670
rect 3930 18490 3950 18510
rect 4010 18650 4030 18670
rect 4010 18490 4030 18510
rect 4090 18650 4110 18670
rect 4090 18490 4110 18510
rect 4170 18650 4190 18670
rect 4170 18490 4190 18510
rect 6250 18650 6270 18670
rect 6250 18490 6270 18510
rect 6330 18650 6350 18670
rect 6330 18490 6350 18510
rect 6410 18650 6430 18670
rect 6410 18490 6430 18510
rect 6490 18650 6510 18670
rect 6490 18490 6510 18510
rect 6570 18650 6590 18670
rect 6570 18490 6590 18510
rect 6650 18650 6670 18670
rect 6650 18490 6670 18510
rect 6730 18650 6750 18670
rect 6730 18490 6750 18510
rect 6810 18650 6830 18670
rect 6810 18490 6830 18510
rect 6890 18650 6910 18670
rect 6890 18490 6910 18510
rect 6970 18650 6990 18670
rect 6970 18490 6990 18510
rect 7050 18650 7070 18670
rect 7050 18490 7070 18510
rect 7130 18650 7150 18670
rect 7130 18490 7150 18510
rect 7210 18650 7230 18670
rect 7210 18490 7230 18510
rect 7290 18650 7310 18670
rect 7290 18490 7310 18510
rect 7370 18650 7390 18670
rect 7370 18490 7390 18510
rect 7450 18650 7470 18670
rect 7450 18490 7470 18510
rect 7530 18650 7550 18670
rect 7530 18490 7550 18510
rect 7610 18650 7630 18670
rect 7610 18490 7630 18510
rect 7690 18650 7710 18670
rect 7690 18490 7710 18510
rect 7770 18650 7790 18670
rect 7770 18490 7790 18510
rect 7850 18650 7870 18670
rect 7850 18490 7870 18510
rect 7930 18650 7950 18670
rect 7930 18490 7950 18510
rect 8010 18650 8030 18670
rect 8010 18490 8030 18510
rect 8090 18650 8110 18670
rect 8090 18490 8110 18510
rect 8170 18650 8190 18670
rect 8170 18490 8190 18510
rect 8250 18650 8270 18670
rect 8250 18490 8270 18510
rect 8330 18650 8350 18670
rect 8330 18490 8350 18510
rect 8410 18650 8430 18670
rect 8410 18490 8430 18510
rect 8490 18650 8510 18670
rect 8490 18490 8510 18510
rect 8570 18650 8590 18670
rect 8570 18490 8590 18510
rect 8650 18650 8670 18670
rect 8650 18490 8670 18510
rect 8730 18650 8750 18670
rect 8730 18490 8750 18510
rect 8810 18650 8830 18670
rect 8810 18490 8830 18510
rect 8890 18650 8910 18670
rect 8890 18490 8910 18510
rect 8970 18650 8990 18670
rect 8970 18490 8990 18510
rect 9050 18650 9070 18670
rect 9050 18490 9070 18510
rect 9130 18650 9150 18670
rect 9130 18490 9150 18510
rect 9210 18650 9230 18670
rect 9210 18490 9230 18510
rect 9290 18650 9310 18670
rect 9290 18490 9310 18510
rect 9370 18650 9390 18670
rect 9370 18490 9390 18510
rect 9450 18650 9470 18670
rect 9450 18490 9470 18510
rect 11570 18650 11590 18670
rect 11570 18490 11590 18510
rect 11650 18650 11670 18670
rect 11650 18490 11670 18510
rect 11730 18650 11750 18670
rect 11730 18490 11750 18510
rect 11810 18650 11830 18670
rect 11810 18490 11830 18510
rect 11890 18650 11910 18670
rect 11890 18490 11910 18510
rect 11970 18650 11990 18670
rect 11970 18490 11990 18510
rect 12050 18650 12070 18670
rect 12050 18490 12070 18510
rect 12130 18650 12150 18670
rect 12130 18490 12150 18510
rect 12210 18650 12230 18670
rect 12210 18490 12230 18510
rect 12290 18650 12310 18670
rect 12290 18490 12310 18510
rect 12370 18650 12390 18670
rect 12370 18490 12390 18510
rect 12450 18650 12470 18670
rect 12450 18490 12470 18510
rect 12530 18650 12550 18670
rect 12530 18490 12550 18510
rect 12610 18650 12630 18670
rect 12610 18490 12630 18510
rect 12690 18650 12710 18670
rect 12690 18490 12710 18510
rect 12770 18650 12790 18670
rect 12770 18490 12790 18510
rect 12850 18650 12870 18670
rect 12850 18490 12870 18510
rect 12930 18650 12950 18670
rect 12930 18490 12950 18510
rect 13010 18650 13030 18670
rect 13010 18490 13030 18510
rect 13090 18650 13110 18670
rect 13090 18490 13110 18510
rect 13170 18650 13190 18670
rect 13170 18490 13190 18510
rect 13250 18650 13270 18670
rect 13250 18490 13270 18510
rect 13330 18650 13350 18670
rect 13330 18490 13350 18510
rect 13410 18650 13430 18670
rect 13410 18490 13430 18510
rect 13490 18650 13510 18670
rect 13490 18490 13510 18510
rect 13570 18650 13590 18670
rect 13570 18490 13590 18510
rect 13650 18650 13670 18670
rect 13650 18490 13670 18510
rect 13730 18650 13750 18670
rect 13730 18490 13750 18510
rect 13810 18650 13830 18670
rect 13810 18490 13830 18510
rect 13890 18650 13910 18670
rect 13890 18490 13910 18510
rect 13970 18650 13990 18670
rect 13970 18490 13990 18510
rect 14050 18650 14070 18670
rect 14050 18490 14070 18510
rect 14130 18650 14150 18670
rect 14130 18490 14150 18510
rect 14210 18650 14230 18670
rect 14210 18490 14230 18510
rect 14290 18650 14310 18670
rect 14290 18490 14310 18510
rect 14370 18650 14390 18670
rect 14370 18490 14390 18510
rect 14450 18650 14470 18670
rect 14450 18490 14470 18510
rect 14530 18650 14550 18670
rect 14530 18490 14550 18510
rect 14610 18650 14630 18670
rect 14610 18490 14630 18510
rect 14690 18650 14710 18670
rect 14690 18490 14710 18510
rect 16770 18650 16790 18670
rect 16770 18490 16790 18510
rect 16850 18650 16870 18670
rect 16850 18490 16870 18510
rect 16930 18650 16950 18670
rect 16930 18490 16950 18510
rect 17010 18650 17030 18670
rect 17010 18490 17030 18510
rect 17090 18650 17110 18670
rect 17090 18490 17110 18510
rect 17170 18650 17190 18670
rect 17170 18490 17190 18510
rect 17250 18650 17270 18670
rect 17250 18490 17270 18510
rect 17330 18650 17350 18670
rect 17330 18490 17350 18510
rect 17410 18650 17430 18670
rect 17410 18490 17430 18510
rect 17490 18650 17510 18670
rect 17490 18490 17510 18510
rect 17570 18650 17590 18670
rect 17570 18490 17590 18510
rect 17650 18650 17670 18670
rect 17650 18490 17670 18510
rect 17730 18650 17750 18670
rect 17730 18490 17750 18510
rect 17810 18650 17830 18670
rect 17810 18490 17830 18510
rect 17890 18650 17910 18670
rect 17890 18490 17910 18510
rect 17970 18650 17990 18670
rect 17970 18490 17990 18510
rect 18050 18650 18070 18670
rect 18050 18490 18070 18510
rect 18130 18650 18150 18670
rect 18130 18490 18150 18510
rect 18210 18650 18230 18670
rect 18210 18490 18230 18510
rect 18290 18650 18310 18670
rect 18290 18490 18310 18510
rect 18370 18650 18390 18670
rect 18370 18490 18390 18510
rect 18450 18650 18470 18670
rect 18450 18490 18470 18510
rect 18530 18650 18550 18670
rect 18530 18490 18550 18510
rect 18610 18650 18630 18670
rect 18610 18490 18630 18510
rect 18690 18650 18710 18670
rect 18690 18490 18710 18510
rect 18770 18650 18790 18670
rect 18770 18490 18790 18510
rect 18850 18650 18870 18670
rect 18850 18490 18870 18510
rect 18930 18650 18950 18670
rect 18930 18490 18950 18510
rect 19010 18650 19030 18670
rect 19010 18490 19030 18510
rect 19090 18650 19110 18670
rect 19090 18490 19110 18510
rect 19170 18650 19190 18670
rect 19170 18490 19190 18510
rect 19250 18650 19270 18670
rect 19250 18490 19270 18510
rect 19330 18650 19350 18670
rect 19330 18490 19350 18510
rect 19410 18650 19430 18670
rect 19410 18490 19430 18510
rect 19490 18650 19510 18670
rect 19490 18490 19510 18510
rect 19570 18650 19590 18670
rect 19570 18490 19590 18510
rect 19650 18650 19670 18670
rect 19650 18490 19670 18510
rect 19730 18650 19750 18670
rect 19730 18490 19750 18510
rect 19810 18650 19830 18670
rect 19810 18490 19830 18510
rect 19890 18650 19910 18670
rect 19890 18490 19910 18510
rect 19970 18650 19990 18670
rect 19970 18490 19990 18510
rect 20050 18650 20070 18670
rect 20050 18490 20070 18510
rect 20130 18650 20150 18670
rect 20130 18490 20150 18510
rect 20210 18650 20230 18670
rect 20210 18490 20230 18510
rect 20290 18650 20310 18670
rect 20290 18490 20310 18510
rect 20370 18650 20390 18670
rect 20370 18490 20390 18510
rect 20450 18650 20470 18670
rect 20450 18490 20470 18510
rect 20530 18650 20550 18670
rect 20530 18490 20550 18510
rect 20610 18650 20630 18670
rect 20610 18490 20630 18510
rect 20690 18650 20710 18670
rect 20690 18490 20710 18510
rect 20770 18650 20790 18670
rect 20770 18490 20790 18510
rect 20850 18650 20870 18670
rect 20850 18490 20870 18510
rect 20930 18650 20950 18670
rect 20930 18490 20950 18510
rect 10 18410 30 18430
rect 10 18250 30 18270
rect 90 18410 110 18430
rect 90 18250 110 18270
rect 170 18410 190 18430
rect 170 18250 190 18270
rect 250 18410 270 18430
rect 250 18250 270 18270
rect 330 18410 350 18430
rect 330 18250 350 18270
rect 410 18410 430 18430
rect 410 18250 430 18270
rect 490 18410 510 18430
rect 490 18250 510 18270
rect 570 18410 590 18430
rect 570 18250 590 18270
rect 650 18410 670 18430
rect 650 18250 670 18270
rect 730 18410 750 18430
rect 730 18250 750 18270
rect 810 18410 830 18430
rect 810 18250 830 18270
rect 890 18410 910 18430
rect 890 18250 910 18270
rect 970 18410 990 18430
rect 970 18250 990 18270
rect 1050 18410 1070 18430
rect 1050 18250 1070 18270
rect 1130 18410 1150 18430
rect 1130 18250 1150 18270
rect 1210 18410 1230 18430
rect 1210 18250 1230 18270
rect 1290 18410 1310 18430
rect 1290 18250 1310 18270
rect 1370 18410 1390 18430
rect 1370 18250 1390 18270
rect 1450 18410 1470 18430
rect 1450 18250 1470 18270
rect 1530 18410 1550 18430
rect 1530 18250 1550 18270
rect 1610 18410 1630 18430
rect 1610 18250 1630 18270
rect 1690 18410 1710 18430
rect 1690 18250 1710 18270
rect 1770 18410 1790 18430
rect 1770 18250 1790 18270
rect 1850 18410 1870 18430
rect 1850 18250 1870 18270
rect 1930 18410 1950 18430
rect 1930 18250 1950 18270
rect 2010 18410 2030 18430
rect 2010 18250 2030 18270
rect 2090 18410 2110 18430
rect 2090 18250 2110 18270
rect 2170 18410 2190 18430
rect 2170 18250 2190 18270
rect 2250 18410 2270 18430
rect 2250 18250 2270 18270
rect 2330 18410 2350 18430
rect 2330 18250 2350 18270
rect 2410 18410 2430 18430
rect 2410 18250 2430 18270
rect 2490 18410 2510 18430
rect 2490 18250 2510 18270
rect 2570 18410 2590 18430
rect 2570 18250 2590 18270
rect 2650 18410 2670 18430
rect 2650 18250 2670 18270
rect 2730 18410 2750 18430
rect 2730 18250 2750 18270
rect 2810 18410 2830 18430
rect 2810 18250 2830 18270
rect 2890 18410 2910 18430
rect 2890 18250 2910 18270
rect 2970 18410 2990 18430
rect 2970 18250 2990 18270
rect 3050 18410 3070 18430
rect 3050 18250 3070 18270
rect 3130 18410 3150 18430
rect 3130 18250 3150 18270
rect 3210 18410 3230 18430
rect 3210 18250 3230 18270
rect 3290 18410 3310 18430
rect 3290 18250 3310 18270
rect 3370 18410 3390 18430
rect 3370 18250 3390 18270
rect 3450 18410 3470 18430
rect 3450 18250 3470 18270
rect 3530 18410 3550 18430
rect 3530 18250 3550 18270
rect 3610 18410 3630 18430
rect 3610 18250 3630 18270
rect 3690 18410 3710 18430
rect 3690 18250 3710 18270
rect 3770 18410 3790 18430
rect 3770 18250 3790 18270
rect 3850 18410 3870 18430
rect 3850 18250 3870 18270
rect 3930 18410 3950 18430
rect 3930 18250 3950 18270
rect 4010 18410 4030 18430
rect 4010 18250 4030 18270
rect 4090 18410 4110 18430
rect 4090 18250 4110 18270
rect 4170 18410 4190 18430
rect 4170 18250 4190 18270
rect 6250 18410 6270 18430
rect 6250 18250 6270 18270
rect 6330 18410 6350 18430
rect 6330 18250 6350 18270
rect 6410 18410 6430 18430
rect 6410 18250 6430 18270
rect 6490 18410 6510 18430
rect 6490 18250 6510 18270
rect 6570 18410 6590 18430
rect 6570 18250 6590 18270
rect 6650 18410 6670 18430
rect 6650 18250 6670 18270
rect 6730 18410 6750 18430
rect 6730 18250 6750 18270
rect 6810 18410 6830 18430
rect 6810 18250 6830 18270
rect 6890 18410 6910 18430
rect 6890 18250 6910 18270
rect 6970 18410 6990 18430
rect 6970 18250 6990 18270
rect 7050 18410 7070 18430
rect 7050 18250 7070 18270
rect 7130 18410 7150 18430
rect 7130 18250 7150 18270
rect 7210 18410 7230 18430
rect 7210 18250 7230 18270
rect 7290 18410 7310 18430
rect 7290 18250 7310 18270
rect 7370 18410 7390 18430
rect 7370 18250 7390 18270
rect 7450 18410 7470 18430
rect 7450 18250 7470 18270
rect 7530 18410 7550 18430
rect 7530 18250 7550 18270
rect 7610 18410 7630 18430
rect 7610 18250 7630 18270
rect 7690 18410 7710 18430
rect 7690 18250 7710 18270
rect 7770 18410 7790 18430
rect 7770 18250 7790 18270
rect 7850 18410 7870 18430
rect 7850 18250 7870 18270
rect 7930 18410 7950 18430
rect 7930 18250 7950 18270
rect 8010 18410 8030 18430
rect 8010 18250 8030 18270
rect 8090 18410 8110 18430
rect 8090 18250 8110 18270
rect 8170 18410 8190 18430
rect 8170 18250 8190 18270
rect 8250 18410 8270 18430
rect 8250 18250 8270 18270
rect 8330 18410 8350 18430
rect 8330 18250 8350 18270
rect 8410 18410 8430 18430
rect 8410 18250 8430 18270
rect 8490 18410 8510 18430
rect 8490 18250 8510 18270
rect 8570 18410 8590 18430
rect 8570 18250 8590 18270
rect 8650 18410 8670 18430
rect 8650 18250 8670 18270
rect 8730 18410 8750 18430
rect 8730 18250 8750 18270
rect 8810 18410 8830 18430
rect 8810 18250 8830 18270
rect 8890 18410 8910 18430
rect 8890 18250 8910 18270
rect 8970 18410 8990 18430
rect 8970 18250 8990 18270
rect 9050 18410 9070 18430
rect 9050 18250 9070 18270
rect 9130 18410 9150 18430
rect 9130 18250 9150 18270
rect 9210 18410 9230 18430
rect 9210 18250 9230 18270
rect 9290 18410 9310 18430
rect 9290 18250 9310 18270
rect 9370 18410 9390 18430
rect 9370 18250 9390 18270
rect 9450 18410 9470 18430
rect 9450 18250 9470 18270
rect 11570 18410 11590 18430
rect 11570 18250 11590 18270
rect 11650 18410 11670 18430
rect 11650 18250 11670 18270
rect 11730 18410 11750 18430
rect 11730 18250 11750 18270
rect 11810 18410 11830 18430
rect 11810 18250 11830 18270
rect 11890 18410 11910 18430
rect 11890 18250 11910 18270
rect 11970 18410 11990 18430
rect 11970 18250 11990 18270
rect 12050 18410 12070 18430
rect 12050 18250 12070 18270
rect 12130 18410 12150 18430
rect 12130 18250 12150 18270
rect 12210 18410 12230 18430
rect 12210 18250 12230 18270
rect 12290 18410 12310 18430
rect 12290 18250 12310 18270
rect 12370 18410 12390 18430
rect 12370 18250 12390 18270
rect 12450 18410 12470 18430
rect 12450 18250 12470 18270
rect 12530 18410 12550 18430
rect 12530 18250 12550 18270
rect 12610 18410 12630 18430
rect 12610 18250 12630 18270
rect 12690 18410 12710 18430
rect 12690 18250 12710 18270
rect 12770 18410 12790 18430
rect 12770 18250 12790 18270
rect 12850 18410 12870 18430
rect 12850 18250 12870 18270
rect 12930 18410 12950 18430
rect 12930 18250 12950 18270
rect 13010 18410 13030 18430
rect 13010 18250 13030 18270
rect 13090 18410 13110 18430
rect 13090 18250 13110 18270
rect 13170 18410 13190 18430
rect 13170 18250 13190 18270
rect 13250 18410 13270 18430
rect 13250 18250 13270 18270
rect 13330 18410 13350 18430
rect 13330 18250 13350 18270
rect 13410 18410 13430 18430
rect 13410 18250 13430 18270
rect 13490 18410 13510 18430
rect 13490 18250 13510 18270
rect 13570 18410 13590 18430
rect 13570 18250 13590 18270
rect 13650 18410 13670 18430
rect 13650 18250 13670 18270
rect 13730 18410 13750 18430
rect 13730 18250 13750 18270
rect 13810 18410 13830 18430
rect 13810 18250 13830 18270
rect 13890 18410 13910 18430
rect 13890 18250 13910 18270
rect 13970 18410 13990 18430
rect 13970 18250 13990 18270
rect 14050 18410 14070 18430
rect 14050 18250 14070 18270
rect 14130 18410 14150 18430
rect 14130 18250 14150 18270
rect 14210 18410 14230 18430
rect 14210 18250 14230 18270
rect 14290 18410 14310 18430
rect 14290 18250 14310 18270
rect 14370 18410 14390 18430
rect 14370 18250 14390 18270
rect 14450 18410 14470 18430
rect 14450 18250 14470 18270
rect 14530 18410 14550 18430
rect 14530 18250 14550 18270
rect 14610 18410 14630 18430
rect 14610 18250 14630 18270
rect 14690 18410 14710 18430
rect 14690 18250 14710 18270
rect 16770 18410 16790 18430
rect 16770 18250 16790 18270
rect 16850 18410 16870 18430
rect 16850 18250 16870 18270
rect 16930 18410 16950 18430
rect 16930 18250 16950 18270
rect 17010 18410 17030 18430
rect 17010 18250 17030 18270
rect 17090 18410 17110 18430
rect 17090 18250 17110 18270
rect 17170 18410 17190 18430
rect 17170 18250 17190 18270
rect 17250 18410 17270 18430
rect 17250 18250 17270 18270
rect 17330 18410 17350 18430
rect 17330 18250 17350 18270
rect 17410 18410 17430 18430
rect 17410 18250 17430 18270
rect 17490 18410 17510 18430
rect 17490 18250 17510 18270
rect 17570 18410 17590 18430
rect 17570 18250 17590 18270
rect 17650 18410 17670 18430
rect 17650 18250 17670 18270
rect 17730 18410 17750 18430
rect 17730 18250 17750 18270
rect 17810 18410 17830 18430
rect 17810 18250 17830 18270
rect 17890 18410 17910 18430
rect 17890 18250 17910 18270
rect 17970 18410 17990 18430
rect 17970 18250 17990 18270
rect 18050 18410 18070 18430
rect 18050 18250 18070 18270
rect 18130 18410 18150 18430
rect 18130 18250 18150 18270
rect 18210 18410 18230 18430
rect 18210 18250 18230 18270
rect 18290 18410 18310 18430
rect 18290 18250 18310 18270
rect 18370 18410 18390 18430
rect 18370 18250 18390 18270
rect 18450 18410 18470 18430
rect 18450 18250 18470 18270
rect 18530 18410 18550 18430
rect 18530 18250 18550 18270
rect 18610 18410 18630 18430
rect 18610 18250 18630 18270
rect 18690 18410 18710 18430
rect 18690 18250 18710 18270
rect 18770 18410 18790 18430
rect 18770 18250 18790 18270
rect 18850 18410 18870 18430
rect 18850 18250 18870 18270
rect 18930 18410 18950 18430
rect 18930 18250 18950 18270
rect 19010 18410 19030 18430
rect 19010 18250 19030 18270
rect 19090 18410 19110 18430
rect 19090 18250 19110 18270
rect 19170 18410 19190 18430
rect 19170 18250 19190 18270
rect 19250 18410 19270 18430
rect 19250 18250 19270 18270
rect 19330 18410 19350 18430
rect 19330 18250 19350 18270
rect 19410 18410 19430 18430
rect 19410 18250 19430 18270
rect 19490 18410 19510 18430
rect 19490 18250 19510 18270
rect 19570 18410 19590 18430
rect 19570 18250 19590 18270
rect 19650 18410 19670 18430
rect 19650 18250 19670 18270
rect 19730 18410 19750 18430
rect 19730 18250 19750 18270
rect 19810 18410 19830 18430
rect 19810 18250 19830 18270
rect 19890 18410 19910 18430
rect 19890 18250 19910 18270
rect 19970 18410 19990 18430
rect 19970 18250 19990 18270
rect 20050 18410 20070 18430
rect 20050 18250 20070 18270
rect 20130 18410 20150 18430
rect 20130 18250 20150 18270
rect 20210 18410 20230 18430
rect 20210 18250 20230 18270
rect 20290 18410 20310 18430
rect 20290 18250 20310 18270
rect 20370 18410 20390 18430
rect 20370 18250 20390 18270
rect 20450 18410 20470 18430
rect 20450 18250 20470 18270
rect 20530 18410 20550 18430
rect 20530 18250 20550 18270
rect 20610 18410 20630 18430
rect 20610 18250 20630 18270
rect 20690 18410 20710 18430
rect 20690 18250 20710 18270
rect 20770 18410 20790 18430
rect 20770 18250 20790 18270
rect 20850 18410 20870 18430
rect 20850 18250 20870 18270
rect 20930 18410 20950 18430
rect 20930 18250 20950 18270
rect 10 18170 30 18190
rect 10 18010 30 18030
rect 10 17850 30 17870
rect 10 17690 30 17710
rect 10 17530 30 17550
rect 10 17370 30 17390
rect 10 17210 30 17230
rect 90 18170 110 18190
rect 90 18010 110 18030
rect 90 17850 110 17870
rect 90 17690 110 17710
rect 90 17530 110 17550
rect 90 17370 110 17390
rect 90 17210 110 17230
rect 170 18170 190 18190
rect 170 18010 190 18030
rect 170 17850 190 17870
rect 170 17690 190 17710
rect 170 17530 190 17550
rect 170 17370 190 17390
rect 170 17210 190 17230
rect 250 18170 270 18190
rect 250 18010 270 18030
rect 250 17850 270 17870
rect 250 17690 270 17710
rect 250 17530 270 17550
rect 250 17370 270 17390
rect 250 17210 270 17230
rect 330 18170 350 18190
rect 330 18010 350 18030
rect 330 17850 350 17870
rect 330 17690 350 17710
rect 330 17530 350 17550
rect 330 17370 350 17390
rect 330 17210 350 17230
rect 410 18170 430 18190
rect 410 18010 430 18030
rect 410 17850 430 17870
rect 410 17690 430 17710
rect 410 17530 430 17550
rect 410 17370 430 17390
rect 410 17210 430 17230
rect 490 18170 510 18190
rect 490 18010 510 18030
rect 490 17850 510 17870
rect 490 17690 510 17710
rect 490 17530 510 17550
rect 490 17370 510 17390
rect 490 17210 510 17230
rect 570 18170 590 18190
rect 570 18010 590 18030
rect 570 17850 590 17870
rect 570 17690 590 17710
rect 570 17530 590 17550
rect 570 17370 590 17390
rect 570 17210 590 17230
rect 650 18170 670 18190
rect 650 18010 670 18030
rect 650 17850 670 17870
rect 650 17690 670 17710
rect 650 17530 670 17550
rect 650 17370 670 17390
rect 650 17210 670 17230
rect 730 18170 750 18190
rect 730 18010 750 18030
rect 730 17850 750 17870
rect 730 17690 750 17710
rect 730 17530 750 17550
rect 730 17370 750 17390
rect 730 17210 750 17230
rect 810 18170 830 18190
rect 810 18010 830 18030
rect 810 17850 830 17870
rect 810 17690 830 17710
rect 810 17530 830 17550
rect 810 17370 830 17390
rect 810 17210 830 17230
rect 890 18170 910 18190
rect 890 18010 910 18030
rect 890 17850 910 17870
rect 890 17690 910 17710
rect 890 17530 910 17550
rect 890 17370 910 17390
rect 890 17210 910 17230
rect 970 18170 990 18190
rect 970 18010 990 18030
rect 970 17850 990 17870
rect 970 17690 990 17710
rect 970 17530 990 17550
rect 970 17370 990 17390
rect 970 17210 990 17230
rect 1050 18170 1070 18190
rect 1050 18010 1070 18030
rect 1050 17850 1070 17870
rect 1050 17690 1070 17710
rect 1050 17530 1070 17550
rect 1050 17370 1070 17390
rect 1050 17210 1070 17230
rect 1130 18170 1150 18190
rect 1130 18010 1150 18030
rect 1130 17850 1150 17870
rect 1130 17690 1150 17710
rect 1130 17530 1150 17550
rect 1130 17370 1150 17390
rect 1130 17210 1150 17230
rect 1210 18170 1230 18190
rect 1210 18010 1230 18030
rect 1210 17850 1230 17870
rect 1210 17690 1230 17710
rect 1210 17530 1230 17550
rect 1210 17370 1230 17390
rect 1210 17210 1230 17230
rect 1290 18170 1310 18190
rect 1290 18010 1310 18030
rect 1290 17850 1310 17870
rect 1290 17690 1310 17710
rect 1290 17530 1310 17550
rect 1290 17370 1310 17390
rect 1290 17210 1310 17230
rect 1370 18170 1390 18190
rect 1370 18010 1390 18030
rect 1370 17850 1390 17870
rect 1370 17690 1390 17710
rect 1370 17530 1390 17550
rect 1370 17370 1390 17390
rect 1370 17210 1390 17230
rect 1450 18170 1470 18190
rect 1450 18010 1470 18030
rect 1450 17850 1470 17870
rect 1450 17690 1470 17710
rect 1450 17530 1470 17550
rect 1450 17370 1470 17390
rect 1450 17210 1470 17230
rect 1530 18170 1550 18190
rect 1530 18010 1550 18030
rect 1530 17850 1550 17870
rect 1530 17690 1550 17710
rect 1530 17530 1550 17550
rect 1530 17370 1550 17390
rect 1530 17210 1550 17230
rect 1610 18170 1630 18190
rect 1610 18010 1630 18030
rect 1610 17850 1630 17870
rect 1610 17690 1630 17710
rect 1610 17530 1630 17550
rect 1610 17370 1630 17390
rect 1610 17210 1630 17230
rect 1690 18170 1710 18190
rect 1690 18010 1710 18030
rect 1690 17850 1710 17870
rect 1690 17690 1710 17710
rect 1690 17530 1710 17550
rect 1690 17370 1710 17390
rect 1690 17210 1710 17230
rect 1770 18170 1790 18190
rect 1770 18010 1790 18030
rect 1770 17850 1790 17870
rect 1770 17690 1790 17710
rect 1770 17530 1790 17550
rect 1770 17370 1790 17390
rect 1770 17210 1790 17230
rect 1850 18170 1870 18190
rect 1850 18010 1870 18030
rect 1850 17850 1870 17870
rect 1850 17690 1870 17710
rect 1850 17530 1870 17550
rect 1850 17370 1870 17390
rect 1850 17210 1870 17230
rect 1930 18170 1950 18190
rect 1930 18010 1950 18030
rect 1930 17850 1950 17870
rect 1930 17690 1950 17710
rect 1930 17530 1950 17550
rect 1930 17370 1950 17390
rect 1930 17210 1950 17230
rect 2010 18170 2030 18190
rect 2010 18010 2030 18030
rect 2010 17850 2030 17870
rect 2010 17690 2030 17710
rect 2010 17530 2030 17550
rect 2010 17370 2030 17390
rect 2010 17210 2030 17230
rect 2090 18170 2110 18190
rect 2090 18010 2110 18030
rect 2090 17850 2110 17870
rect 2090 17690 2110 17710
rect 2090 17530 2110 17550
rect 2090 17370 2110 17390
rect 2090 17210 2110 17230
rect 2170 18170 2190 18190
rect 2170 18010 2190 18030
rect 2170 17850 2190 17870
rect 2170 17690 2190 17710
rect 2170 17530 2190 17550
rect 2170 17370 2190 17390
rect 2170 17210 2190 17230
rect 2250 18170 2270 18190
rect 2250 18010 2270 18030
rect 2250 17850 2270 17870
rect 2250 17690 2270 17710
rect 2250 17530 2270 17550
rect 2250 17370 2270 17390
rect 2250 17210 2270 17230
rect 2330 18170 2350 18190
rect 2330 18010 2350 18030
rect 2330 17850 2350 17870
rect 2330 17690 2350 17710
rect 2330 17530 2350 17550
rect 2330 17370 2350 17390
rect 2330 17210 2350 17230
rect 2410 18170 2430 18190
rect 2410 18010 2430 18030
rect 2410 17850 2430 17870
rect 2410 17690 2430 17710
rect 2410 17530 2430 17550
rect 2410 17370 2430 17390
rect 2410 17210 2430 17230
rect 2490 18170 2510 18190
rect 2490 18010 2510 18030
rect 2490 17850 2510 17870
rect 2490 17690 2510 17710
rect 2490 17530 2510 17550
rect 2490 17370 2510 17390
rect 2490 17210 2510 17230
rect 2570 18170 2590 18190
rect 2570 18010 2590 18030
rect 2570 17850 2590 17870
rect 2570 17690 2590 17710
rect 2570 17530 2590 17550
rect 2570 17370 2590 17390
rect 2570 17210 2590 17230
rect 2650 18170 2670 18190
rect 2650 18010 2670 18030
rect 2650 17850 2670 17870
rect 2650 17690 2670 17710
rect 2650 17530 2670 17550
rect 2650 17370 2670 17390
rect 2650 17210 2670 17230
rect 2730 18170 2750 18190
rect 2730 18010 2750 18030
rect 2730 17850 2750 17870
rect 2730 17690 2750 17710
rect 2730 17530 2750 17550
rect 2730 17370 2750 17390
rect 2730 17210 2750 17230
rect 2810 18170 2830 18190
rect 2810 18010 2830 18030
rect 2810 17850 2830 17870
rect 2810 17690 2830 17710
rect 2810 17530 2830 17550
rect 2810 17370 2830 17390
rect 2810 17210 2830 17230
rect 2890 18170 2910 18190
rect 2890 18010 2910 18030
rect 2890 17850 2910 17870
rect 2890 17690 2910 17710
rect 2890 17530 2910 17550
rect 2890 17370 2910 17390
rect 2890 17210 2910 17230
rect 2970 18170 2990 18190
rect 2970 18010 2990 18030
rect 2970 17850 2990 17870
rect 2970 17690 2990 17710
rect 2970 17530 2990 17550
rect 2970 17370 2990 17390
rect 2970 17210 2990 17230
rect 3050 18170 3070 18190
rect 3050 18010 3070 18030
rect 3050 17850 3070 17870
rect 3050 17690 3070 17710
rect 3050 17530 3070 17550
rect 3050 17370 3070 17390
rect 3050 17210 3070 17230
rect 3130 18170 3150 18190
rect 3130 18010 3150 18030
rect 3130 17850 3150 17870
rect 3130 17690 3150 17710
rect 3130 17530 3150 17550
rect 3130 17370 3150 17390
rect 3130 17210 3150 17230
rect 3210 18170 3230 18190
rect 3210 18010 3230 18030
rect 3210 17850 3230 17870
rect 3210 17690 3230 17710
rect 3210 17530 3230 17550
rect 3210 17370 3230 17390
rect 3210 17210 3230 17230
rect 3290 18170 3310 18190
rect 3290 18010 3310 18030
rect 3290 17850 3310 17870
rect 3290 17690 3310 17710
rect 3290 17530 3310 17550
rect 3290 17370 3310 17390
rect 3290 17210 3310 17230
rect 3370 18170 3390 18190
rect 3370 18010 3390 18030
rect 3370 17850 3390 17870
rect 3370 17690 3390 17710
rect 3370 17530 3390 17550
rect 3370 17370 3390 17390
rect 3370 17210 3390 17230
rect 3450 18170 3470 18190
rect 3450 18010 3470 18030
rect 3450 17850 3470 17870
rect 3450 17690 3470 17710
rect 3450 17530 3470 17550
rect 3450 17370 3470 17390
rect 3450 17210 3470 17230
rect 3530 18170 3550 18190
rect 3530 18010 3550 18030
rect 3530 17850 3550 17870
rect 3530 17690 3550 17710
rect 3530 17530 3550 17550
rect 3530 17370 3550 17390
rect 3530 17210 3550 17230
rect 3610 18170 3630 18190
rect 3610 18010 3630 18030
rect 3610 17850 3630 17870
rect 3610 17690 3630 17710
rect 3610 17530 3630 17550
rect 3610 17370 3630 17390
rect 3610 17210 3630 17230
rect 3690 18170 3710 18190
rect 3690 18010 3710 18030
rect 3690 17850 3710 17870
rect 3690 17690 3710 17710
rect 3690 17530 3710 17550
rect 3690 17370 3710 17390
rect 3690 17210 3710 17230
rect 3770 18170 3790 18190
rect 3770 18010 3790 18030
rect 3770 17850 3790 17870
rect 3770 17690 3790 17710
rect 3770 17530 3790 17550
rect 3770 17370 3790 17390
rect 3770 17210 3790 17230
rect 3850 18170 3870 18190
rect 3850 18010 3870 18030
rect 3850 17850 3870 17870
rect 3850 17690 3870 17710
rect 3850 17530 3870 17550
rect 3850 17370 3870 17390
rect 3850 17210 3870 17230
rect 3930 18170 3950 18190
rect 3930 18010 3950 18030
rect 3930 17850 3950 17870
rect 3930 17690 3950 17710
rect 3930 17530 3950 17550
rect 3930 17370 3950 17390
rect 3930 17210 3950 17230
rect 4010 18170 4030 18190
rect 4010 18010 4030 18030
rect 4010 17850 4030 17870
rect 4010 17690 4030 17710
rect 4010 17530 4030 17550
rect 4010 17370 4030 17390
rect 4010 17210 4030 17230
rect 4090 18170 4110 18190
rect 4090 18010 4110 18030
rect 4090 17850 4110 17870
rect 4090 17690 4110 17710
rect 4090 17530 4110 17550
rect 4090 17370 4110 17390
rect 4090 17210 4110 17230
rect 4170 18170 4190 18190
rect 4170 18010 4190 18030
rect 4170 17850 4190 17870
rect 4170 17690 4190 17710
rect 4170 17530 4190 17550
rect 4170 17370 4190 17390
rect 4170 17210 4190 17230
rect 6250 18170 6270 18190
rect 6250 18010 6270 18030
rect 6250 17850 6270 17870
rect 6250 17690 6270 17710
rect 6250 17530 6270 17550
rect 6250 17370 6270 17390
rect 6250 17210 6270 17230
rect 6330 18170 6350 18190
rect 6330 18010 6350 18030
rect 6330 17850 6350 17870
rect 6330 17690 6350 17710
rect 6330 17530 6350 17550
rect 6330 17370 6350 17390
rect 6330 17210 6350 17230
rect 6410 18170 6430 18190
rect 6410 18010 6430 18030
rect 6410 17850 6430 17870
rect 6410 17690 6430 17710
rect 6410 17530 6430 17550
rect 6410 17370 6430 17390
rect 6410 17210 6430 17230
rect 6490 18170 6510 18190
rect 6490 18010 6510 18030
rect 6490 17850 6510 17870
rect 6490 17690 6510 17710
rect 6490 17530 6510 17550
rect 6490 17370 6510 17390
rect 6490 17210 6510 17230
rect 6570 18170 6590 18190
rect 6570 18010 6590 18030
rect 6570 17850 6590 17870
rect 6570 17690 6590 17710
rect 6570 17530 6590 17550
rect 6570 17370 6590 17390
rect 6570 17210 6590 17230
rect 6650 18170 6670 18190
rect 6650 18010 6670 18030
rect 6650 17850 6670 17870
rect 6650 17690 6670 17710
rect 6650 17530 6670 17550
rect 6650 17370 6670 17390
rect 6650 17210 6670 17230
rect 6730 18170 6750 18190
rect 6730 18010 6750 18030
rect 6730 17850 6750 17870
rect 6730 17690 6750 17710
rect 6730 17530 6750 17550
rect 6730 17370 6750 17390
rect 6730 17210 6750 17230
rect 6810 18170 6830 18190
rect 6810 18010 6830 18030
rect 6810 17850 6830 17870
rect 6810 17690 6830 17710
rect 6810 17530 6830 17550
rect 6810 17370 6830 17390
rect 6810 17210 6830 17230
rect 6890 18170 6910 18190
rect 6890 18010 6910 18030
rect 6890 17850 6910 17870
rect 6890 17690 6910 17710
rect 6890 17530 6910 17550
rect 6890 17370 6910 17390
rect 6890 17210 6910 17230
rect 6970 18170 6990 18190
rect 6970 18010 6990 18030
rect 6970 17850 6990 17870
rect 6970 17690 6990 17710
rect 6970 17530 6990 17550
rect 6970 17370 6990 17390
rect 6970 17210 6990 17230
rect 7050 18170 7070 18190
rect 7050 18010 7070 18030
rect 7050 17850 7070 17870
rect 7050 17690 7070 17710
rect 7050 17530 7070 17550
rect 7050 17370 7070 17390
rect 7050 17210 7070 17230
rect 7130 18170 7150 18190
rect 7130 18010 7150 18030
rect 7130 17850 7150 17870
rect 7130 17690 7150 17710
rect 7130 17530 7150 17550
rect 7130 17370 7150 17390
rect 7130 17210 7150 17230
rect 7210 18170 7230 18190
rect 7210 18010 7230 18030
rect 7210 17850 7230 17870
rect 7210 17690 7230 17710
rect 7210 17530 7230 17550
rect 7210 17370 7230 17390
rect 7210 17210 7230 17230
rect 7290 18170 7310 18190
rect 7290 18010 7310 18030
rect 7290 17850 7310 17870
rect 7290 17690 7310 17710
rect 7290 17530 7310 17550
rect 7290 17370 7310 17390
rect 7290 17210 7310 17230
rect 7370 18170 7390 18190
rect 7370 18010 7390 18030
rect 7370 17850 7390 17870
rect 7370 17690 7390 17710
rect 7370 17530 7390 17550
rect 7370 17370 7390 17390
rect 7370 17210 7390 17230
rect 7450 18170 7470 18190
rect 7450 18010 7470 18030
rect 7450 17850 7470 17870
rect 7450 17690 7470 17710
rect 7450 17530 7470 17550
rect 7450 17370 7470 17390
rect 7450 17210 7470 17230
rect 7530 18170 7550 18190
rect 7530 18010 7550 18030
rect 7530 17850 7550 17870
rect 7530 17690 7550 17710
rect 7530 17530 7550 17550
rect 7530 17370 7550 17390
rect 7530 17210 7550 17230
rect 7610 18170 7630 18190
rect 7610 18010 7630 18030
rect 7610 17850 7630 17870
rect 7610 17690 7630 17710
rect 7610 17530 7630 17550
rect 7610 17370 7630 17390
rect 7610 17210 7630 17230
rect 7690 18170 7710 18190
rect 7690 18010 7710 18030
rect 7690 17850 7710 17870
rect 7690 17690 7710 17710
rect 7690 17530 7710 17550
rect 7690 17370 7710 17390
rect 7690 17210 7710 17230
rect 7770 18170 7790 18190
rect 7770 18010 7790 18030
rect 7770 17850 7790 17870
rect 7770 17690 7790 17710
rect 7770 17530 7790 17550
rect 7770 17370 7790 17390
rect 7770 17210 7790 17230
rect 7850 18170 7870 18190
rect 7850 18010 7870 18030
rect 7850 17850 7870 17870
rect 7850 17690 7870 17710
rect 7850 17530 7870 17550
rect 7850 17370 7870 17390
rect 7850 17210 7870 17230
rect 7930 18170 7950 18190
rect 7930 18010 7950 18030
rect 7930 17850 7950 17870
rect 7930 17690 7950 17710
rect 7930 17530 7950 17550
rect 7930 17370 7950 17390
rect 7930 17210 7950 17230
rect 8010 18170 8030 18190
rect 8010 18010 8030 18030
rect 8010 17850 8030 17870
rect 8010 17690 8030 17710
rect 8010 17530 8030 17550
rect 8010 17370 8030 17390
rect 8010 17210 8030 17230
rect 8090 18170 8110 18190
rect 8090 18010 8110 18030
rect 8090 17850 8110 17870
rect 8090 17690 8110 17710
rect 8090 17530 8110 17550
rect 8090 17370 8110 17390
rect 8090 17210 8110 17230
rect 8170 18170 8190 18190
rect 8170 18010 8190 18030
rect 8170 17850 8190 17870
rect 8170 17690 8190 17710
rect 8170 17530 8190 17550
rect 8170 17370 8190 17390
rect 8170 17210 8190 17230
rect 8250 18170 8270 18190
rect 8250 18010 8270 18030
rect 8250 17850 8270 17870
rect 8250 17690 8270 17710
rect 8250 17530 8270 17550
rect 8250 17370 8270 17390
rect 8250 17210 8270 17230
rect 8330 18170 8350 18190
rect 8330 18010 8350 18030
rect 8330 17850 8350 17870
rect 8330 17690 8350 17710
rect 8330 17530 8350 17550
rect 8330 17370 8350 17390
rect 8330 17210 8350 17230
rect 8410 18170 8430 18190
rect 8410 18010 8430 18030
rect 8410 17850 8430 17870
rect 8410 17690 8430 17710
rect 8410 17530 8430 17550
rect 8410 17370 8430 17390
rect 8410 17210 8430 17230
rect 8490 18170 8510 18190
rect 8490 18010 8510 18030
rect 8490 17850 8510 17870
rect 8490 17690 8510 17710
rect 8490 17530 8510 17550
rect 8490 17370 8510 17390
rect 8490 17210 8510 17230
rect 8570 18170 8590 18190
rect 8570 18010 8590 18030
rect 8570 17850 8590 17870
rect 8570 17690 8590 17710
rect 8570 17530 8590 17550
rect 8570 17370 8590 17390
rect 8570 17210 8590 17230
rect 8650 18170 8670 18190
rect 8650 18010 8670 18030
rect 8650 17850 8670 17870
rect 8650 17690 8670 17710
rect 8650 17530 8670 17550
rect 8650 17370 8670 17390
rect 8650 17210 8670 17230
rect 8730 18170 8750 18190
rect 8730 18010 8750 18030
rect 8730 17850 8750 17870
rect 8730 17690 8750 17710
rect 8730 17530 8750 17550
rect 8730 17370 8750 17390
rect 8730 17210 8750 17230
rect 8810 18170 8830 18190
rect 8810 18010 8830 18030
rect 8810 17850 8830 17870
rect 8810 17690 8830 17710
rect 8810 17530 8830 17550
rect 8810 17370 8830 17390
rect 8810 17210 8830 17230
rect 8890 18170 8910 18190
rect 8890 18010 8910 18030
rect 8890 17850 8910 17870
rect 8890 17690 8910 17710
rect 8890 17530 8910 17550
rect 8890 17370 8910 17390
rect 8890 17210 8910 17230
rect 8970 18170 8990 18190
rect 8970 18010 8990 18030
rect 8970 17850 8990 17870
rect 8970 17690 8990 17710
rect 8970 17530 8990 17550
rect 8970 17370 8990 17390
rect 8970 17210 8990 17230
rect 9050 18170 9070 18190
rect 9050 18010 9070 18030
rect 9050 17850 9070 17870
rect 9050 17690 9070 17710
rect 9050 17530 9070 17550
rect 9050 17370 9070 17390
rect 9050 17210 9070 17230
rect 9130 18170 9150 18190
rect 9130 18010 9150 18030
rect 9130 17850 9150 17870
rect 9130 17690 9150 17710
rect 9130 17530 9150 17550
rect 9130 17370 9150 17390
rect 9130 17210 9150 17230
rect 9210 18170 9230 18190
rect 9210 18010 9230 18030
rect 9210 17850 9230 17870
rect 9210 17690 9230 17710
rect 9210 17530 9230 17550
rect 9210 17370 9230 17390
rect 9210 17210 9230 17230
rect 9290 18170 9310 18190
rect 9290 18010 9310 18030
rect 9290 17850 9310 17870
rect 9290 17690 9310 17710
rect 9290 17530 9310 17550
rect 9290 17370 9310 17390
rect 9290 17210 9310 17230
rect 9370 18170 9390 18190
rect 9370 18010 9390 18030
rect 9370 17850 9390 17870
rect 9370 17690 9390 17710
rect 9370 17530 9390 17550
rect 9370 17370 9390 17390
rect 9370 17210 9390 17230
rect 9450 18170 9470 18190
rect 9450 18010 9470 18030
rect 9450 17850 9470 17870
rect 9450 17690 9470 17710
rect 9450 17530 9470 17550
rect 9450 17370 9470 17390
rect 9450 17210 9470 17230
rect 11570 18170 11590 18190
rect 11570 18010 11590 18030
rect 11570 17850 11590 17870
rect 11570 17690 11590 17710
rect 11570 17530 11590 17550
rect 11570 17370 11590 17390
rect 11570 17210 11590 17230
rect 11650 18170 11670 18190
rect 11650 18010 11670 18030
rect 11650 17850 11670 17870
rect 11650 17690 11670 17710
rect 11650 17530 11670 17550
rect 11650 17370 11670 17390
rect 11650 17210 11670 17230
rect 11730 18170 11750 18190
rect 11730 18010 11750 18030
rect 11730 17850 11750 17870
rect 11730 17690 11750 17710
rect 11730 17530 11750 17550
rect 11730 17370 11750 17390
rect 11730 17210 11750 17230
rect 11810 18170 11830 18190
rect 11810 18010 11830 18030
rect 11810 17850 11830 17870
rect 11810 17690 11830 17710
rect 11810 17530 11830 17550
rect 11810 17370 11830 17390
rect 11810 17210 11830 17230
rect 11890 18170 11910 18190
rect 11890 18010 11910 18030
rect 11890 17850 11910 17870
rect 11890 17690 11910 17710
rect 11890 17530 11910 17550
rect 11890 17370 11910 17390
rect 11890 17210 11910 17230
rect 11970 18170 11990 18190
rect 11970 18010 11990 18030
rect 11970 17850 11990 17870
rect 11970 17690 11990 17710
rect 11970 17530 11990 17550
rect 11970 17370 11990 17390
rect 11970 17210 11990 17230
rect 12050 18170 12070 18190
rect 12050 18010 12070 18030
rect 12050 17850 12070 17870
rect 12050 17690 12070 17710
rect 12050 17530 12070 17550
rect 12050 17370 12070 17390
rect 12050 17210 12070 17230
rect 12130 18170 12150 18190
rect 12130 18010 12150 18030
rect 12130 17850 12150 17870
rect 12130 17690 12150 17710
rect 12130 17530 12150 17550
rect 12130 17370 12150 17390
rect 12130 17210 12150 17230
rect 12210 18170 12230 18190
rect 12210 18010 12230 18030
rect 12210 17850 12230 17870
rect 12210 17690 12230 17710
rect 12210 17530 12230 17550
rect 12210 17370 12230 17390
rect 12210 17210 12230 17230
rect 12290 18170 12310 18190
rect 12290 18010 12310 18030
rect 12290 17850 12310 17870
rect 12290 17690 12310 17710
rect 12290 17530 12310 17550
rect 12290 17370 12310 17390
rect 12290 17210 12310 17230
rect 12370 18170 12390 18190
rect 12370 18010 12390 18030
rect 12370 17850 12390 17870
rect 12370 17690 12390 17710
rect 12370 17530 12390 17550
rect 12370 17370 12390 17390
rect 12370 17210 12390 17230
rect 12450 18170 12470 18190
rect 12450 18010 12470 18030
rect 12450 17850 12470 17870
rect 12450 17690 12470 17710
rect 12450 17530 12470 17550
rect 12450 17370 12470 17390
rect 12450 17210 12470 17230
rect 12530 18170 12550 18190
rect 12530 18010 12550 18030
rect 12530 17850 12550 17870
rect 12530 17690 12550 17710
rect 12530 17530 12550 17550
rect 12530 17370 12550 17390
rect 12530 17210 12550 17230
rect 12610 18170 12630 18190
rect 12610 18010 12630 18030
rect 12610 17850 12630 17870
rect 12610 17690 12630 17710
rect 12610 17530 12630 17550
rect 12610 17370 12630 17390
rect 12610 17210 12630 17230
rect 12690 18170 12710 18190
rect 12690 18010 12710 18030
rect 12690 17850 12710 17870
rect 12690 17690 12710 17710
rect 12690 17530 12710 17550
rect 12690 17370 12710 17390
rect 12690 17210 12710 17230
rect 12770 18170 12790 18190
rect 12770 18010 12790 18030
rect 12770 17850 12790 17870
rect 12770 17690 12790 17710
rect 12770 17530 12790 17550
rect 12770 17370 12790 17390
rect 12770 17210 12790 17230
rect 12850 18170 12870 18190
rect 12850 18010 12870 18030
rect 12850 17850 12870 17870
rect 12850 17690 12870 17710
rect 12850 17530 12870 17550
rect 12850 17370 12870 17390
rect 12850 17210 12870 17230
rect 12930 18170 12950 18190
rect 12930 18010 12950 18030
rect 12930 17850 12950 17870
rect 12930 17690 12950 17710
rect 12930 17530 12950 17550
rect 12930 17370 12950 17390
rect 12930 17210 12950 17230
rect 13010 18170 13030 18190
rect 13010 18010 13030 18030
rect 13010 17850 13030 17870
rect 13010 17690 13030 17710
rect 13010 17530 13030 17550
rect 13010 17370 13030 17390
rect 13010 17210 13030 17230
rect 13090 18170 13110 18190
rect 13090 18010 13110 18030
rect 13090 17850 13110 17870
rect 13090 17690 13110 17710
rect 13090 17530 13110 17550
rect 13090 17370 13110 17390
rect 13090 17210 13110 17230
rect 13170 18170 13190 18190
rect 13170 18010 13190 18030
rect 13170 17850 13190 17870
rect 13170 17690 13190 17710
rect 13170 17530 13190 17550
rect 13170 17370 13190 17390
rect 13170 17210 13190 17230
rect 13250 18170 13270 18190
rect 13250 18010 13270 18030
rect 13250 17850 13270 17870
rect 13250 17690 13270 17710
rect 13250 17530 13270 17550
rect 13250 17370 13270 17390
rect 13250 17210 13270 17230
rect 13330 18170 13350 18190
rect 13330 18010 13350 18030
rect 13330 17850 13350 17870
rect 13330 17690 13350 17710
rect 13330 17530 13350 17550
rect 13330 17370 13350 17390
rect 13330 17210 13350 17230
rect 13410 18170 13430 18190
rect 13410 18010 13430 18030
rect 13410 17850 13430 17870
rect 13410 17690 13430 17710
rect 13410 17530 13430 17550
rect 13410 17370 13430 17390
rect 13410 17210 13430 17230
rect 13490 18170 13510 18190
rect 13490 18010 13510 18030
rect 13490 17850 13510 17870
rect 13490 17690 13510 17710
rect 13490 17530 13510 17550
rect 13490 17370 13510 17390
rect 13490 17210 13510 17230
rect 13570 18170 13590 18190
rect 13570 18010 13590 18030
rect 13570 17850 13590 17870
rect 13570 17690 13590 17710
rect 13570 17530 13590 17550
rect 13570 17370 13590 17390
rect 13570 17210 13590 17230
rect 13650 18170 13670 18190
rect 13650 18010 13670 18030
rect 13650 17850 13670 17870
rect 13650 17690 13670 17710
rect 13650 17530 13670 17550
rect 13650 17370 13670 17390
rect 13650 17210 13670 17230
rect 13730 18170 13750 18190
rect 13730 18010 13750 18030
rect 13730 17850 13750 17870
rect 13730 17690 13750 17710
rect 13730 17530 13750 17550
rect 13730 17370 13750 17390
rect 13730 17210 13750 17230
rect 13810 18170 13830 18190
rect 13810 18010 13830 18030
rect 13810 17850 13830 17870
rect 13810 17690 13830 17710
rect 13810 17530 13830 17550
rect 13810 17370 13830 17390
rect 13810 17210 13830 17230
rect 13890 18170 13910 18190
rect 13890 18010 13910 18030
rect 13890 17850 13910 17870
rect 13890 17690 13910 17710
rect 13890 17530 13910 17550
rect 13890 17370 13910 17390
rect 13890 17210 13910 17230
rect 13970 18170 13990 18190
rect 13970 18010 13990 18030
rect 13970 17850 13990 17870
rect 13970 17690 13990 17710
rect 13970 17530 13990 17550
rect 13970 17370 13990 17390
rect 13970 17210 13990 17230
rect 14050 18170 14070 18190
rect 14050 18010 14070 18030
rect 14050 17850 14070 17870
rect 14050 17690 14070 17710
rect 14050 17530 14070 17550
rect 14050 17370 14070 17390
rect 14050 17210 14070 17230
rect 14130 18170 14150 18190
rect 14130 18010 14150 18030
rect 14130 17850 14150 17870
rect 14130 17690 14150 17710
rect 14130 17530 14150 17550
rect 14130 17370 14150 17390
rect 14130 17210 14150 17230
rect 14210 18170 14230 18190
rect 14210 18010 14230 18030
rect 14210 17850 14230 17870
rect 14210 17690 14230 17710
rect 14210 17530 14230 17550
rect 14210 17370 14230 17390
rect 14210 17210 14230 17230
rect 14290 18170 14310 18190
rect 14290 18010 14310 18030
rect 14290 17850 14310 17870
rect 14290 17690 14310 17710
rect 14290 17530 14310 17550
rect 14290 17370 14310 17390
rect 14290 17210 14310 17230
rect 14370 18170 14390 18190
rect 14370 18010 14390 18030
rect 14370 17850 14390 17870
rect 14370 17690 14390 17710
rect 14370 17530 14390 17550
rect 14370 17370 14390 17390
rect 14370 17210 14390 17230
rect 14450 18170 14470 18190
rect 14450 18010 14470 18030
rect 14450 17850 14470 17870
rect 14450 17690 14470 17710
rect 14450 17530 14470 17550
rect 14450 17370 14470 17390
rect 14450 17210 14470 17230
rect 14530 18170 14550 18190
rect 14530 18010 14550 18030
rect 14530 17850 14550 17870
rect 14530 17690 14550 17710
rect 14530 17530 14550 17550
rect 14530 17370 14550 17390
rect 14530 17210 14550 17230
rect 14610 18170 14630 18190
rect 14610 18010 14630 18030
rect 14610 17850 14630 17870
rect 14610 17690 14630 17710
rect 14610 17530 14630 17550
rect 14610 17370 14630 17390
rect 14610 17210 14630 17230
rect 14690 18170 14710 18190
rect 14690 18010 14710 18030
rect 14690 17850 14710 17870
rect 14690 17690 14710 17710
rect 14690 17530 14710 17550
rect 14690 17370 14710 17390
rect 14690 17210 14710 17230
rect 16770 18170 16790 18190
rect 16770 18010 16790 18030
rect 16770 17850 16790 17870
rect 16770 17690 16790 17710
rect 16770 17530 16790 17550
rect 16770 17370 16790 17390
rect 16770 17210 16790 17230
rect 16850 18170 16870 18190
rect 16850 18010 16870 18030
rect 16850 17850 16870 17870
rect 16850 17690 16870 17710
rect 16850 17530 16870 17550
rect 16850 17370 16870 17390
rect 16850 17210 16870 17230
rect 16930 18170 16950 18190
rect 16930 18010 16950 18030
rect 16930 17850 16950 17870
rect 16930 17690 16950 17710
rect 16930 17530 16950 17550
rect 16930 17370 16950 17390
rect 16930 17210 16950 17230
rect 17010 18170 17030 18190
rect 17010 18010 17030 18030
rect 17010 17850 17030 17870
rect 17010 17690 17030 17710
rect 17010 17530 17030 17550
rect 17010 17370 17030 17390
rect 17010 17210 17030 17230
rect 17090 18170 17110 18190
rect 17090 18010 17110 18030
rect 17090 17850 17110 17870
rect 17090 17690 17110 17710
rect 17090 17530 17110 17550
rect 17090 17370 17110 17390
rect 17090 17210 17110 17230
rect 17170 18170 17190 18190
rect 17170 18010 17190 18030
rect 17170 17850 17190 17870
rect 17170 17690 17190 17710
rect 17170 17530 17190 17550
rect 17170 17370 17190 17390
rect 17170 17210 17190 17230
rect 17250 18170 17270 18190
rect 17250 18010 17270 18030
rect 17250 17850 17270 17870
rect 17250 17690 17270 17710
rect 17250 17530 17270 17550
rect 17250 17370 17270 17390
rect 17250 17210 17270 17230
rect 17330 18170 17350 18190
rect 17330 18010 17350 18030
rect 17330 17850 17350 17870
rect 17330 17690 17350 17710
rect 17330 17530 17350 17550
rect 17330 17370 17350 17390
rect 17330 17210 17350 17230
rect 17410 18170 17430 18190
rect 17410 18010 17430 18030
rect 17410 17850 17430 17870
rect 17410 17690 17430 17710
rect 17410 17530 17430 17550
rect 17410 17370 17430 17390
rect 17410 17210 17430 17230
rect 17490 18170 17510 18190
rect 17490 18010 17510 18030
rect 17490 17850 17510 17870
rect 17490 17690 17510 17710
rect 17490 17530 17510 17550
rect 17490 17370 17510 17390
rect 17490 17210 17510 17230
rect 17570 18170 17590 18190
rect 17570 18010 17590 18030
rect 17570 17850 17590 17870
rect 17570 17690 17590 17710
rect 17570 17530 17590 17550
rect 17570 17370 17590 17390
rect 17570 17210 17590 17230
rect 17650 18170 17670 18190
rect 17650 18010 17670 18030
rect 17650 17850 17670 17870
rect 17650 17690 17670 17710
rect 17650 17530 17670 17550
rect 17650 17370 17670 17390
rect 17650 17210 17670 17230
rect 17730 18170 17750 18190
rect 17730 18010 17750 18030
rect 17730 17850 17750 17870
rect 17730 17690 17750 17710
rect 17730 17530 17750 17550
rect 17730 17370 17750 17390
rect 17730 17210 17750 17230
rect 17810 18170 17830 18190
rect 17810 18010 17830 18030
rect 17810 17850 17830 17870
rect 17810 17690 17830 17710
rect 17810 17530 17830 17550
rect 17810 17370 17830 17390
rect 17810 17210 17830 17230
rect 17890 18170 17910 18190
rect 17890 18010 17910 18030
rect 17890 17850 17910 17870
rect 17890 17690 17910 17710
rect 17890 17530 17910 17550
rect 17890 17370 17910 17390
rect 17890 17210 17910 17230
rect 17970 18170 17990 18190
rect 17970 18010 17990 18030
rect 17970 17850 17990 17870
rect 17970 17690 17990 17710
rect 17970 17530 17990 17550
rect 17970 17370 17990 17390
rect 17970 17210 17990 17230
rect 18050 18170 18070 18190
rect 18050 18010 18070 18030
rect 18050 17850 18070 17870
rect 18050 17690 18070 17710
rect 18050 17530 18070 17550
rect 18050 17370 18070 17390
rect 18050 17210 18070 17230
rect 18130 18170 18150 18190
rect 18130 18010 18150 18030
rect 18130 17850 18150 17870
rect 18130 17690 18150 17710
rect 18130 17530 18150 17550
rect 18130 17370 18150 17390
rect 18130 17210 18150 17230
rect 18210 18170 18230 18190
rect 18210 18010 18230 18030
rect 18210 17850 18230 17870
rect 18210 17690 18230 17710
rect 18210 17530 18230 17550
rect 18210 17370 18230 17390
rect 18210 17210 18230 17230
rect 18290 18170 18310 18190
rect 18290 18010 18310 18030
rect 18290 17850 18310 17870
rect 18290 17690 18310 17710
rect 18290 17530 18310 17550
rect 18290 17370 18310 17390
rect 18290 17210 18310 17230
rect 18370 18170 18390 18190
rect 18370 18010 18390 18030
rect 18370 17850 18390 17870
rect 18370 17690 18390 17710
rect 18370 17530 18390 17550
rect 18370 17370 18390 17390
rect 18370 17210 18390 17230
rect 18450 18170 18470 18190
rect 18450 18010 18470 18030
rect 18450 17850 18470 17870
rect 18450 17690 18470 17710
rect 18450 17530 18470 17550
rect 18450 17370 18470 17390
rect 18450 17210 18470 17230
rect 18530 18170 18550 18190
rect 18530 18010 18550 18030
rect 18530 17850 18550 17870
rect 18530 17690 18550 17710
rect 18530 17530 18550 17550
rect 18530 17370 18550 17390
rect 18530 17210 18550 17230
rect 18610 18170 18630 18190
rect 18610 18010 18630 18030
rect 18610 17850 18630 17870
rect 18610 17690 18630 17710
rect 18610 17530 18630 17550
rect 18610 17370 18630 17390
rect 18610 17210 18630 17230
rect 18690 18170 18710 18190
rect 18690 18010 18710 18030
rect 18690 17850 18710 17870
rect 18690 17690 18710 17710
rect 18690 17530 18710 17550
rect 18690 17370 18710 17390
rect 18690 17210 18710 17230
rect 18770 18170 18790 18190
rect 18770 18010 18790 18030
rect 18770 17850 18790 17870
rect 18770 17690 18790 17710
rect 18770 17530 18790 17550
rect 18770 17370 18790 17390
rect 18770 17210 18790 17230
rect 18850 18170 18870 18190
rect 18850 18010 18870 18030
rect 18850 17850 18870 17870
rect 18850 17690 18870 17710
rect 18850 17530 18870 17550
rect 18850 17370 18870 17390
rect 18850 17210 18870 17230
rect 18930 18170 18950 18190
rect 18930 18010 18950 18030
rect 18930 17850 18950 17870
rect 18930 17690 18950 17710
rect 18930 17530 18950 17550
rect 18930 17370 18950 17390
rect 18930 17210 18950 17230
rect 19010 18170 19030 18190
rect 19010 18010 19030 18030
rect 19010 17850 19030 17870
rect 19010 17690 19030 17710
rect 19010 17530 19030 17550
rect 19010 17370 19030 17390
rect 19010 17210 19030 17230
rect 19090 18170 19110 18190
rect 19090 18010 19110 18030
rect 19090 17850 19110 17870
rect 19090 17690 19110 17710
rect 19090 17530 19110 17550
rect 19090 17370 19110 17390
rect 19090 17210 19110 17230
rect 19170 18170 19190 18190
rect 19170 18010 19190 18030
rect 19170 17850 19190 17870
rect 19170 17690 19190 17710
rect 19170 17530 19190 17550
rect 19170 17370 19190 17390
rect 19170 17210 19190 17230
rect 19250 18170 19270 18190
rect 19250 18010 19270 18030
rect 19250 17850 19270 17870
rect 19250 17690 19270 17710
rect 19250 17530 19270 17550
rect 19250 17370 19270 17390
rect 19250 17210 19270 17230
rect 19330 18170 19350 18190
rect 19330 18010 19350 18030
rect 19330 17850 19350 17870
rect 19330 17690 19350 17710
rect 19330 17530 19350 17550
rect 19330 17370 19350 17390
rect 19330 17210 19350 17230
rect 19410 18170 19430 18190
rect 19410 18010 19430 18030
rect 19410 17850 19430 17870
rect 19410 17690 19430 17710
rect 19410 17530 19430 17550
rect 19410 17370 19430 17390
rect 19410 17210 19430 17230
rect 19490 18170 19510 18190
rect 19490 18010 19510 18030
rect 19490 17850 19510 17870
rect 19490 17690 19510 17710
rect 19490 17530 19510 17550
rect 19490 17370 19510 17390
rect 19490 17210 19510 17230
rect 19570 18170 19590 18190
rect 19570 18010 19590 18030
rect 19570 17850 19590 17870
rect 19570 17690 19590 17710
rect 19570 17530 19590 17550
rect 19570 17370 19590 17390
rect 19570 17210 19590 17230
rect 19650 18170 19670 18190
rect 19650 18010 19670 18030
rect 19650 17850 19670 17870
rect 19650 17690 19670 17710
rect 19650 17530 19670 17550
rect 19650 17370 19670 17390
rect 19650 17210 19670 17230
rect 19730 18170 19750 18190
rect 19730 18010 19750 18030
rect 19730 17850 19750 17870
rect 19730 17690 19750 17710
rect 19730 17530 19750 17550
rect 19730 17370 19750 17390
rect 19730 17210 19750 17230
rect 19810 18170 19830 18190
rect 19810 18010 19830 18030
rect 19810 17850 19830 17870
rect 19810 17690 19830 17710
rect 19810 17530 19830 17550
rect 19810 17370 19830 17390
rect 19810 17210 19830 17230
rect 19890 18170 19910 18190
rect 19890 18010 19910 18030
rect 19890 17850 19910 17870
rect 19890 17690 19910 17710
rect 19890 17530 19910 17550
rect 19890 17370 19910 17390
rect 19890 17210 19910 17230
rect 19970 18170 19990 18190
rect 19970 18010 19990 18030
rect 19970 17850 19990 17870
rect 19970 17690 19990 17710
rect 19970 17530 19990 17550
rect 19970 17370 19990 17390
rect 19970 17210 19990 17230
rect 20050 18170 20070 18190
rect 20050 18010 20070 18030
rect 20050 17850 20070 17870
rect 20050 17690 20070 17710
rect 20050 17530 20070 17550
rect 20050 17370 20070 17390
rect 20050 17210 20070 17230
rect 20130 18170 20150 18190
rect 20130 18010 20150 18030
rect 20130 17850 20150 17870
rect 20130 17690 20150 17710
rect 20130 17530 20150 17550
rect 20130 17370 20150 17390
rect 20130 17210 20150 17230
rect 20210 18170 20230 18190
rect 20210 18010 20230 18030
rect 20210 17850 20230 17870
rect 20210 17690 20230 17710
rect 20210 17530 20230 17550
rect 20210 17370 20230 17390
rect 20210 17210 20230 17230
rect 20290 18170 20310 18190
rect 20290 18010 20310 18030
rect 20290 17850 20310 17870
rect 20290 17690 20310 17710
rect 20290 17530 20310 17550
rect 20290 17370 20310 17390
rect 20290 17210 20310 17230
rect 20370 18170 20390 18190
rect 20370 18010 20390 18030
rect 20370 17850 20390 17870
rect 20370 17690 20390 17710
rect 20370 17530 20390 17550
rect 20370 17370 20390 17390
rect 20370 17210 20390 17230
rect 20450 18170 20470 18190
rect 20450 18010 20470 18030
rect 20450 17850 20470 17870
rect 20450 17690 20470 17710
rect 20450 17530 20470 17550
rect 20450 17370 20470 17390
rect 20450 17210 20470 17230
rect 20530 18170 20550 18190
rect 20530 18010 20550 18030
rect 20530 17850 20550 17870
rect 20530 17690 20550 17710
rect 20530 17530 20550 17550
rect 20530 17370 20550 17390
rect 20530 17210 20550 17230
rect 20610 18170 20630 18190
rect 20610 18010 20630 18030
rect 20610 17850 20630 17870
rect 20610 17690 20630 17710
rect 20610 17530 20630 17550
rect 20610 17370 20630 17390
rect 20610 17210 20630 17230
rect 20690 18170 20710 18190
rect 20690 18010 20710 18030
rect 20690 17850 20710 17870
rect 20690 17690 20710 17710
rect 20690 17530 20710 17550
rect 20690 17370 20710 17390
rect 20690 17210 20710 17230
rect 20770 18170 20790 18190
rect 20770 18010 20790 18030
rect 20770 17850 20790 17870
rect 20770 17690 20790 17710
rect 20770 17530 20790 17550
rect 20770 17370 20790 17390
rect 20770 17210 20790 17230
rect 20850 18170 20870 18190
rect 20850 18010 20870 18030
rect 20850 17850 20870 17870
rect 20850 17690 20870 17710
rect 20850 17530 20870 17550
rect 20850 17370 20870 17390
rect 20850 17210 20870 17230
rect 20930 18170 20950 18190
rect 20930 18010 20950 18030
rect 20930 17850 20950 17870
rect 20930 17690 20950 17710
rect 20930 17530 20950 17550
rect 20930 17370 20950 17390
rect 20930 17210 20950 17230
rect 10 17130 30 17150
rect 10 16970 30 16990
rect 90 17130 110 17150
rect 90 16970 110 16990
rect 170 17130 190 17150
rect 170 16970 190 16990
rect 250 17130 270 17150
rect 250 16970 270 16990
rect 330 17130 350 17150
rect 330 16970 350 16990
rect 410 17130 430 17150
rect 410 16970 430 16990
rect 490 17130 510 17150
rect 490 16970 510 16990
rect 570 17130 590 17150
rect 570 16970 590 16990
rect 650 17130 670 17150
rect 650 16970 670 16990
rect 730 17130 750 17150
rect 730 16970 750 16990
rect 810 17130 830 17150
rect 810 16970 830 16990
rect 890 17130 910 17150
rect 890 16970 910 16990
rect 970 17130 990 17150
rect 970 16970 990 16990
rect 1050 17130 1070 17150
rect 1050 16970 1070 16990
rect 1130 17130 1150 17150
rect 1130 16970 1150 16990
rect 1210 17130 1230 17150
rect 1210 16970 1230 16990
rect 1290 17130 1310 17150
rect 1290 16970 1310 16990
rect 1370 17130 1390 17150
rect 1370 16970 1390 16990
rect 1450 17130 1470 17150
rect 1450 16970 1470 16990
rect 1530 17130 1550 17150
rect 1530 16970 1550 16990
rect 1610 17130 1630 17150
rect 1610 16970 1630 16990
rect 1690 17130 1710 17150
rect 1690 16970 1710 16990
rect 1770 17130 1790 17150
rect 1770 16970 1790 16990
rect 1850 17130 1870 17150
rect 1850 16970 1870 16990
rect 1930 17130 1950 17150
rect 1930 16970 1950 16990
rect 2010 17130 2030 17150
rect 2010 16970 2030 16990
rect 2090 17130 2110 17150
rect 2090 16970 2110 16990
rect 2170 17130 2190 17150
rect 2170 16970 2190 16990
rect 2250 17130 2270 17150
rect 2250 16970 2270 16990
rect 2330 17130 2350 17150
rect 2330 16970 2350 16990
rect 2410 17130 2430 17150
rect 2410 16970 2430 16990
rect 2490 17130 2510 17150
rect 2490 16970 2510 16990
rect 2570 17130 2590 17150
rect 2570 16970 2590 16990
rect 2650 17130 2670 17150
rect 2650 16970 2670 16990
rect 2730 17130 2750 17150
rect 2730 16970 2750 16990
rect 2810 17130 2830 17150
rect 2810 16970 2830 16990
rect 2890 17130 2910 17150
rect 2890 16970 2910 16990
rect 2970 17130 2990 17150
rect 2970 16970 2990 16990
rect 3050 17130 3070 17150
rect 3050 16970 3070 16990
rect 3130 17130 3150 17150
rect 3130 16970 3150 16990
rect 3210 17130 3230 17150
rect 3210 16970 3230 16990
rect 3290 17130 3310 17150
rect 3290 16970 3310 16990
rect 3370 17130 3390 17150
rect 3370 16970 3390 16990
rect 3450 17130 3470 17150
rect 3450 16970 3470 16990
rect 3530 17130 3550 17150
rect 3530 16970 3550 16990
rect 3610 17130 3630 17150
rect 3610 16970 3630 16990
rect 3690 17130 3710 17150
rect 3690 16970 3710 16990
rect 3770 17130 3790 17150
rect 3770 16970 3790 16990
rect 3850 17130 3870 17150
rect 3850 16970 3870 16990
rect 3930 17130 3950 17150
rect 3930 16970 3950 16990
rect 4010 17130 4030 17150
rect 4010 16970 4030 16990
rect 4090 17130 4110 17150
rect 4090 16970 4110 16990
rect 4170 17130 4190 17150
rect 4170 16970 4190 16990
rect 6250 17130 6270 17150
rect 6250 16970 6270 16990
rect 6330 17130 6350 17150
rect 6330 16970 6350 16990
rect 6410 17130 6430 17150
rect 6410 16970 6430 16990
rect 6490 17130 6510 17150
rect 6490 16970 6510 16990
rect 6570 17130 6590 17150
rect 6570 16970 6590 16990
rect 6650 17130 6670 17150
rect 6650 16970 6670 16990
rect 6730 17130 6750 17150
rect 6730 16970 6750 16990
rect 6810 17130 6830 17150
rect 6810 16970 6830 16990
rect 6890 17130 6910 17150
rect 6890 16970 6910 16990
rect 6970 17130 6990 17150
rect 6970 16970 6990 16990
rect 7050 17130 7070 17150
rect 7050 16970 7070 16990
rect 7130 17130 7150 17150
rect 7130 16970 7150 16990
rect 7210 17130 7230 17150
rect 7210 16970 7230 16990
rect 7290 17130 7310 17150
rect 7290 16970 7310 16990
rect 7370 17130 7390 17150
rect 7370 16970 7390 16990
rect 7450 17130 7470 17150
rect 7450 16970 7470 16990
rect 7530 17130 7550 17150
rect 7530 16970 7550 16990
rect 7610 17130 7630 17150
rect 7610 16970 7630 16990
rect 7690 17130 7710 17150
rect 7690 16970 7710 16990
rect 7770 17130 7790 17150
rect 7770 16970 7790 16990
rect 7850 17130 7870 17150
rect 7850 16970 7870 16990
rect 7930 17130 7950 17150
rect 7930 16970 7950 16990
rect 8010 17130 8030 17150
rect 8010 16970 8030 16990
rect 8090 17130 8110 17150
rect 8090 16970 8110 16990
rect 8170 17130 8190 17150
rect 8170 16970 8190 16990
rect 8250 17130 8270 17150
rect 8250 16970 8270 16990
rect 8330 17130 8350 17150
rect 8330 16970 8350 16990
rect 8410 17130 8430 17150
rect 8410 16970 8430 16990
rect 8490 17130 8510 17150
rect 8490 16970 8510 16990
rect 8570 17130 8590 17150
rect 8570 16970 8590 16990
rect 8650 17130 8670 17150
rect 8650 16970 8670 16990
rect 8730 17130 8750 17150
rect 8730 16970 8750 16990
rect 8810 17130 8830 17150
rect 8810 16970 8830 16990
rect 8890 17130 8910 17150
rect 8890 16970 8910 16990
rect 8970 17130 8990 17150
rect 8970 16970 8990 16990
rect 9050 17130 9070 17150
rect 9050 16970 9070 16990
rect 9130 17130 9150 17150
rect 9130 16970 9150 16990
rect 9210 17130 9230 17150
rect 9210 16970 9230 16990
rect 9290 17130 9310 17150
rect 9290 16970 9310 16990
rect 9370 17130 9390 17150
rect 9370 16970 9390 16990
rect 9450 17130 9470 17150
rect 9450 16970 9470 16990
rect 11570 17130 11590 17150
rect 11570 16970 11590 16990
rect 11650 17130 11670 17150
rect 11650 16970 11670 16990
rect 11730 17130 11750 17150
rect 11730 16970 11750 16990
rect 11810 17130 11830 17150
rect 11810 16970 11830 16990
rect 11890 17130 11910 17150
rect 11890 16970 11910 16990
rect 11970 17130 11990 17150
rect 11970 16970 11990 16990
rect 12050 17130 12070 17150
rect 12050 16970 12070 16990
rect 12130 17130 12150 17150
rect 12130 16970 12150 16990
rect 12210 17130 12230 17150
rect 12210 16970 12230 16990
rect 12290 17130 12310 17150
rect 12290 16970 12310 16990
rect 12370 17130 12390 17150
rect 12370 16970 12390 16990
rect 12450 17130 12470 17150
rect 12450 16970 12470 16990
rect 12530 17130 12550 17150
rect 12530 16970 12550 16990
rect 12610 17130 12630 17150
rect 12610 16970 12630 16990
rect 12690 17130 12710 17150
rect 12690 16970 12710 16990
rect 12770 17130 12790 17150
rect 12770 16970 12790 16990
rect 12850 17130 12870 17150
rect 12850 16970 12870 16990
rect 12930 17130 12950 17150
rect 12930 16970 12950 16990
rect 13010 17130 13030 17150
rect 13010 16970 13030 16990
rect 13090 17130 13110 17150
rect 13090 16970 13110 16990
rect 13170 17130 13190 17150
rect 13170 16970 13190 16990
rect 13250 17130 13270 17150
rect 13250 16970 13270 16990
rect 13330 17130 13350 17150
rect 13330 16970 13350 16990
rect 13410 17130 13430 17150
rect 13410 16970 13430 16990
rect 13490 17130 13510 17150
rect 13490 16970 13510 16990
rect 13570 17130 13590 17150
rect 13570 16970 13590 16990
rect 13650 17130 13670 17150
rect 13650 16970 13670 16990
rect 13730 17130 13750 17150
rect 13730 16970 13750 16990
rect 13810 17130 13830 17150
rect 13810 16970 13830 16990
rect 13890 17130 13910 17150
rect 13890 16970 13910 16990
rect 13970 17130 13990 17150
rect 13970 16970 13990 16990
rect 14050 17130 14070 17150
rect 14050 16970 14070 16990
rect 14130 17130 14150 17150
rect 14130 16970 14150 16990
rect 14210 17130 14230 17150
rect 14210 16970 14230 16990
rect 14290 17130 14310 17150
rect 14290 16970 14310 16990
rect 14370 17130 14390 17150
rect 14370 16970 14390 16990
rect 14450 17130 14470 17150
rect 14450 16970 14470 16990
rect 14530 17130 14550 17150
rect 14530 16970 14550 16990
rect 14610 17130 14630 17150
rect 14610 16970 14630 16990
rect 14690 17130 14710 17150
rect 14690 16970 14710 16990
rect 16770 17130 16790 17150
rect 16770 16970 16790 16990
rect 16850 17130 16870 17150
rect 16850 16970 16870 16990
rect 16930 17130 16950 17150
rect 16930 16970 16950 16990
rect 17010 17130 17030 17150
rect 17010 16970 17030 16990
rect 17090 17130 17110 17150
rect 17090 16970 17110 16990
rect 17170 17130 17190 17150
rect 17170 16970 17190 16990
rect 17250 17130 17270 17150
rect 17250 16970 17270 16990
rect 17330 17130 17350 17150
rect 17330 16970 17350 16990
rect 17410 17130 17430 17150
rect 17410 16970 17430 16990
rect 17490 17130 17510 17150
rect 17490 16970 17510 16990
rect 17570 17130 17590 17150
rect 17570 16970 17590 16990
rect 17650 17130 17670 17150
rect 17650 16970 17670 16990
rect 17730 17130 17750 17150
rect 17730 16970 17750 16990
rect 17810 17130 17830 17150
rect 17810 16970 17830 16990
rect 17890 17130 17910 17150
rect 17890 16970 17910 16990
rect 17970 17130 17990 17150
rect 17970 16970 17990 16990
rect 18050 17130 18070 17150
rect 18050 16970 18070 16990
rect 18130 17130 18150 17150
rect 18130 16970 18150 16990
rect 18210 17130 18230 17150
rect 18210 16970 18230 16990
rect 18290 17130 18310 17150
rect 18290 16970 18310 16990
rect 18370 17130 18390 17150
rect 18370 16970 18390 16990
rect 18450 17130 18470 17150
rect 18450 16970 18470 16990
rect 18530 17130 18550 17150
rect 18530 16970 18550 16990
rect 18610 17130 18630 17150
rect 18610 16970 18630 16990
rect 18690 17130 18710 17150
rect 18690 16970 18710 16990
rect 18770 17130 18790 17150
rect 18770 16970 18790 16990
rect 18850 17130 18870 17150
rect 18850 16970 18870 16990
rect 18930 17130 18950 17150
rect 18930 16970 18950 16990
rect 19010 17130 19030 17150
rect 19010 16970 19030 16990
rect 19090 17130 19110 17150
rect 19090 16970 19110 16990
rect 19170 17130 19190 17150
rect 19170 16970 19190 16990
rect 19250 17130 19270 17150
rect 19250 16970 19270 16990
rect 19330 17130 19350 17150
rect 19330 16970 19350 16990
rect 19410 17130 19430 17150
rect 19410 16970 19430 16990
rect 19490 17130 19510 17150
rect 19490 16970 19510 16990
rect 19570 17130 19590 17150
rect 19570 16970 19590 16990
rect 19650 17130 19670 17150
rect 19650 16970 19670 16990
rect 19730 17130 19750 17150
rect 19730 16970 19750 16990
rect 19810 17130 19830 17150
rect 19810 16970 19830 16990
rect 19890 17130 19910 17150
rect 19890 16970 19910 16990
rect 19970 17130 19990 17150
rect 19970 16970 19990 16990
rect 20050 17130 20070 17150
rect 20050 16970 20070 16990
rect 20130 17130 20150 17150
rect 20130 16970 20150 16990
rect 20210 17130 20230 17150
rect 20210 16970 20230 16990
rect 20290 17130 20310 17150
rect 20290 16970 20310 16990
rect 20370 17130 20390 17150
rect 20370 16970 20390 16990
rect 20450 17130 20470 17150
rect 20450 16970 20470 16990
rect 20530 17130 20550 17150
rect 20530 16970 20550 16990
rect 20610 17130 20630 17150
rect 20610 16970 20630 16990
rect 20690 17130 20710 17150
rect 20690 16970 20710 16990
rect 20770 17130 20790 17150
rect 20770 16970 20790 16990
rect 20850 17130 20870 17150
rect 20850 16970 20870 16990
rect 20930 17130 20950 17150
rect 20930 16970 20950 16990
rect 10 16890 30 16910
rect 10 16730 30 16750
rect 90 16890 110 16910
rect 90 16730 110 16750
rect 170 16890 190 16910
rect 170 16730 190 16750
rect 250 16890 270 16910
rect 250 16730 270 16750
rect 330 16890 350 16910
rect 330 16730 350 16750
rect 410 16890 430 16910
rect 410 16730 430 16750
rect 490 16890 510 16910
rect 490 16730 510 16750
rect 570 16890 590 16910
rect 570 16730 590 16750
rect 650 16890 670 16910
rect 650 16730 670 16750
rect 730 16890 750 16910
rect 730 16730 750 16750
rect 810 16890 830 16910
rect 810 16730 830 16750
rect 890 16890 910 16910
rect 890 16730 910 16750
rect 970 16890 990 16910
rect 970 16730 990 16750
rect 1050 16890 1070 16910
rect 1050 16730 1070 16750
rect 1130 16890 1150 16910
rect 1130 16730 1150 16750
rect 1210 16890 1230 16910
rect 1210 16730 1230 16750
rect 1290 16890 1310 16910
rect 1290 16730 1310 16750
rect 1370 16890 1390 16910
rect 1370 16730 1390 16750
rect 1450 16890 1470 16910
rect 1450 16730 1470 16750
rect 1530 16890 1550 16910
rect 1530 16730 1550 16750
rect 1610 16890 1630 16910
rect 1610 16730 1630 16750
rect 1690 16890 1710 16910
rect 1690 16730 1710 16750
rect 1770 16890 1790 16910
rect 1770 16730 1790 16750
rect 1850 16890 1870 16910
rect 1850 16730 1870 16750
rect 1930 16890 1950 16910
rect 1930 16730 1950 16750
rect 2010 16890 2030 16910
rect 2010 16730 2030 16750
rect 2090 16890 2110 16910
rect 2090 16730 2110 16750
rect 2170 16890 2190 16910
rect 2170 16730 2190 16750
rect 2250 16890 2270 16910
rect 2250 16730 2270 16750
rect 2330 16890 2350 16910
rect 2330 16730 2350 16750
rect 2410 16890 2430 16910
rect 2410 16730 2430 16750
rect 2490 16890 2510 16910
rect 2490 16730 2510 16750
rect 2570 16890 2590 16910
rect 2570 16730 2590 16750
rect 2650 16890 2670 16910
rect 2650 16730 2670 16750
rect 2730 16890 2750 16910
rect 2730 16730 2750 16750
rect 2810 16890 2830 16910
rect 2810 16730 2830 16750
rect 2890 16890 2910 16910
rect 2890 16730 2910 16750
rect 2970 16890 2990 16910
rect 2970 16730 2990 16750
rect 3050 16890 3070 16910
rect 3050 16730 3070 16750
rect 3130 16890 3150 16910
rect 3130 16730 3150 16750
rect 3210 16890 3230 16910
rect 3210 16730 3230 16750
rect 3290 16890 3310 16910
rect 3290 16730 3310 16750
rect 3370 16890 3390 16910
rect 3370 16730 3390 16750
rect 3450 16890 3470 16910
rect 3450 16730 3470 16750
rect 3530 16890 3550 16910
rect 3530 16730 3550 16750
rect 3610 16890 3630 16910
rect 3610 16730 3630 16750
rect 3690 16890 3710 16910
rect 3690 16730 3710 16750
rect 3770 16890 3790 16910
rect 3770 16730 3790 16750
rect 3850 16890 3870 16910
rect 3850 16730 3870 16750
rect 3930 16890 3950 16910
rect 3930 16730 3950 16750
rect 4010 16890 4030 16910
rect 4010 16730 4030 16750
rect 4090 16890 4110 16910
rect 4090 16730 4110 16750
rect 4170 16890 4190 16910
rect 4170 16730 4190 16750
rect 6250 16890 6270 16910
rect 6250 16730 6270 16750
rect 6330 16890 6350 16910
rect 6330 16730 6350 16750
rect 6410 16890 6430 16910
rect 6410 16730 6430 16750
rect 6490 16890 6510 16910
rect 6490 16730 6510 16750
rect 6570 16890 6590 16910
rect 6570 16730 6590 16750
rect 6650 16890 6670 16910
rect 6650 16730 6670 16750
rect 6730 16890 6750 16910
rect 6730 16730 6750 16750
rect 6810 16890 6830 16910
rect 6810 16730 6830 16750
rect 6890 16890 6910 16910
rect 6890 16730 6910 16750
rect 6970 16890 6990 16910
rect 6970 16730 6990 16750
rect 7050 16890 7070 16910
rect 7050 16730 7070 16750
rect 7130 16890 7150 16910
rect 7130 16730 7150 16750
rect 7210 16890 7230 16910
rect 7210 16730 7230 16750
rect 7290 16890 7310 16910
rect 7290 16730 7310 16750
rect 7370 16890 7390 16910
rect 7370 16730 7390 16750
rect 7450 16890 7470 16910
rect 7450 16730 7470 16750
rect 7530 16890 7550 16910
rect 7530 16730 7550 16750
rect 7610 16890 7630 16910
rect 7610 16730 7630 16750
rect 7690 16890 7710 16910
rect 7690 16730 7710 16750
rect 7770 16890 7790 16910
rect 7770 16730 7790 16750
rect 7850 16890 7870 16910
rect 7850 16730 7870 16750
rect 7930 16890 7950 16910
rect 7930 16730 7950 16750
rect 8010 16890 8030 16910
rect 8010 16730 8030 16750
rect 8090 16890 8110 16910
rect 8090 16730 8110 16750
rect 8170 16890 8190 16910
rect 8170 16730 8190 16750
rect 8250 16890 8270 16910
rect 8250 16730 8270 16750
rect 8330 16890 8350 16910
rect 8330 16730 8350 16750
rect 8410 16890 8430 16910
rect 8410 16730 8430 16750
rect 8490 16890 8510 16910
rect 8490 16730 8510 16750
rect 8570 16890 8590 16910
rect 8570 16730 8590 16750
rect 8650 16890 8670 16910
rect 8650 16730 8670 16750
rect 8730 16890 8750 16910
rect 8730 16730 8750 16750
rect 8810 16890 8830 16910
rect 8810 16730 8830 16750
rect 8890 16890 8910 16910
rect 8890 16730 8910 16750
rect 8970 16890 8990 16910
rect 8970 16730 8990 16750
rect 9050 16890 9070 16910
rect 9050 16730 9070 16750
rect 9130 16890 9150 16910
rect 9130 16730 9150 16750
rect 9210 16890 9230 16910
rect 9210 16730 9230 16750
rect 9290 16890 9310 16910
rect 9290 16730 9310 16750
rect 9370 16890 9390 16910
rect 9370 16730 9390 16750
rect 9450 16890 9470 16910
rect 9450 16730 9470 16750
rect 11570 16890 11590 16910
rect 11570 16730 11590 16750
rect 11650 16890 11670 16910
rect 11650 16730 11670 16750
rect 11730 16890 11750 16910
rect 11730 16730 11750 16750
rect 11810 16890 11830 16910
rect 11810 16730 11830 16750
rect 11890 16890 11910 16910
rect 11890 16730 11910 16750
rect 11970 16890 11990 16910
rect 11970 16730 11990 16750
rect 12050 16890 12070 16910
rect 12050 16730 12070 16750
rect 12130 16890 12150 16910
rect 12130 16730 12150 16750
rect 12210 16890 12230 16910
rect 12210 16730 12230 16750
rect 12290 16890 12310 16910
rect 12290 16730 12310 16750
rect 12370 16890 12390 16910
rect 12370 16730 12390 16750
rect 12450 16890 12470 16910
rect 12450 16730 12470 16750
rect 12530 16890 12550 16910
rect 12530 16730 12550 16750
rect 12610 16890 12630 16910
rect 12610 16730 12630 16750
rect 12690 16890 12710 16910
rect 12690 16730 12710 16750
rect 12770 16890 12790 16910
rect 12770 16730 12790 16750
rect 12850 16890 12870 16910
rect 12850 16730 12870 16750
rect 12930 16890 12950 16910
rect 12930 16730 12950 16750
rect 13010 16890 13030 16910
rect 13010 16730 13030 16750
rect 13090 16890 13110 16910
rect 13090 16730 13110 16750
rect 13170 16890 13190 16910
rect 13170 16730 13190 16750
rect 13250 16890 13270 16910
rect 13250 16730 13270 16750
rect 13330 16890 13350 16910
rect 13330 16730 13350 16750
rect 13410 16890 13430 16910
rect 13410 16730 13430 16750
rect 13490 16890 13510 16910
rect 13490 16730 13510 16750
rect 13570 16890 13590 16910
rect 13570 16730 13590 16750
rect 13650 16890 13670 16910
rect 13650 16730 13670 16750
rect 13730 16890 13750 16910
rect 13730 16730 13750 16750
rect 13810 16890 13830 16910
rect 13810 16730 13830 16750
rect 13890 16890 13910 16910
rect 13890 16730 13910 16750
rect 13970 16890 13990 16910
rect 13970 16730 13990 16750
rect 14050 16890 14070 16910
rect 14050 16730 14070 16750
rect 14130 16890 14150 16910
rect 14130 16730 14150 16750
rect 14210 16890 14230 16910
rect 14210 16730 14230 16750
rect 14290 16890 14310 16910
rect 14290 16730 14310 16750
rect 14370 16890 14390 16910
rect 14370 16730 14390 16750
rect 14450 16890 14470 16910
rect 14450 16730 14470 16750
rect 14530 16890 14550 16910
rect 14530 16730 14550 16750
rect 14610 16890 14630 16910
rect 14610 16730 14630 16750
rect 14690 16890 14710 16910
rect 14690 16730 14710 16750
rect 16770 16890 16790 16910
rect 16770 16730 16790 16750
rect 16850 16890 16870 16910
rect 16850 16730 16870 16750
rect 16930 16890 16950 16910
rect 16930 16730 16950 16750
rect 17010 16890 17030 16910
rect 17010 16730 17030 16750
rect 17090 16890 17110 16910
rect 17090 16730 17110 16750
rect 17170 16890 17190 16910
rect 17170 16730 17190 16750
rect 17250 16890 17270 16910
rect 17250 16730 17270 16750
rect 17330 16890 17350 16910
rect 17330 16730 17350 16750
rect 17410 16890 17430 16910
rect 17410 16730 17430 16750
rect 17490 16890 17510 16910
rect 17490 16730 17510 16750
rect 17570 16890 17590 16910
rect 17570 16730 17590 16750
rect 17650 16890 17670 16910
rect 17650 16730 17670 16750
rect 17730 16890 17750 16910
rect 17730 16730 17750 16750
rect 17810 16890 17830 16910
rect 17810 16730 17830 16750
rect 17890 16890 17910 16910
rect 17890 16730 17910 16750
rect 17970 16890 17990 16910
rect 17970 16730 17990 16750
rect 18050 16890 18070 16910
rect 18050 16730 18070 16750
rect 18130 16890 18150 16910
rect 18130 16730 18150 16750
rect 18210 16890 18230 16910
rect 18210 16730 18230 16750
rect 18290 16890 18310 16910
rect 18290 16730 18310 16750
rect 18370 16890 18390 16910
rect 18370 16730 18390 16750
rect 18450 16890 18470 16910
rect 18450 16730 18470 16750
rect 18530 16890 18550 16910
rect 18530 16730 18550 16750
rect 18610 16890 18630 16910
rect 18610 16730 18630 16750
rect 18690 16890 18710 16910
rect 18690 16730 18710 16750
rect 18770 16890 18790 16910
rect 18770 16730 18790 16750
rect 18850 16890 18870 16910
rect 18850 16730 18870 16750
rect 18930 16890 18950 16910
rect 18930 16730 18950 16750
rect 19010 16890 19030 16910
rect 19010 16730 19030 16750
rect 19090 16890 19110 16910
rect 19090 16730 19110 16750
rect 19170 16890 19190 16910
rect 19170 16730 19190 16750
rect 19250 16890 19270 16910
rect 19250 16730 19270 16750
rect 19330 16890 19350 16910
rect 19330 16730 19350 16750
rect 19410 16890 19430 16910
rect 19410 16730 19430 16750
rect 19490 16890 19510 16910
rect 19490 16730 19510 16750
rect 19570 16890 19590 16910
rect 19570 16730 19590 16750
rect 19650 16890 19670 16910
rect 19650 16730 19670 16750
rect 19730 16890 19750 16910
rect 19730 16730 19750 16750
rect 19810 16890 19830 16910
rect 19810 16730 19830 16750
rect 19890 16890 19910 16910
rect 19890 16730 19910 16750
rect 19970 16890 19990 16910
rect 19970 16730 19990 16750
rect 20050 16890 20070 16910
rect 20050 16730 20070 16750
rect 20130 16890 20150 16910
rect 20130 16730 20150 16750
rect 20210 16890 20230 16910
rect 20210 16730 20230 16750
rect 20290 16890 20310 16910
rect 20290 16730 20310 16750
rect 20370 16890 20390 16910
rect 20370 16730 20390 16750
rect 20450 16890 20470 16910
rect 20450 16730 20470 16750
rect 20530 16890 20550 16910
rect 20530 16730 20550 16750
rect 20610 16890 20630 16910
rect 20610 16730 20630 16750
rect 20690 16890 20710 16910
rect 20690 16730 20710 16750
rect 20770 16890 20790 16910
rect 20770 16730 20790 16750
rect 20850 16890 20870 16910
rect 20850 16730 20870 16750
rect 20930 16890 20950 16910
rect 20930 16730 20950 16750
rect 10 16650 30 16670
rect 10 16490 30 16510
rect 90 16650 110 16670
rect 90 16490 110 16510
rect 170 16650 190 16670
rect 170 16490 190 16510
rect 250 16650 270 16670
rect 250 16490 270 16510
rect 330 16650 350 16670
rect 330 16490 350 16510
rect 410 16650 430 16670
rect 410 16490 430 16510
rect 490 16650 510 16670
rect 490 16490 510 16510
rect 570 16650 590 16670
rect 570 16490 590 16510
rect 650 16650 670 16670
rect 650 16490 670 16510
rect 730 16650 750 16670
rect 730 16490 750 16510
rect 810 16650 830 16670
rect 810 16490 830 16510
rect 890 16650 910 16670
rect 890 16490 910 16510
rect 970 16650 990 16670
rect 970 16490 990 16510
rect 1050 16650 1070 16670
rect 1050 16490 1070 16510
rect 1130 16650 1150 16670
rect 1130 16490 1150 16510
rect 1210 16650 1230 16670
rect 1210 16490 1230 16510
rect 1290 16650 1310 16670
rect 1290 16490 1310 16510
rect 1370 16650 1390 16670
rect 1370 16490 1390 16510
rect 1450 16650 1470 16670
rect 1450 16490 1470 16510
rect 1530 16650 1550 16670
rect 1530 16490 1550 16510
rect 1610 16650 1630 16670
rect 1610 16490 1630 16510
rect 1690 16650 1710 16670
rect 1690 16490 1710 16510
rect 1770 16650 1790 16670
rect 1770 16490 1790 16510
rect 1850 16650 1870 16670
rect 1850 16490 1870 16510
rect 1930 16650 1950 16670
rect 1930 16490 1950 16510
rect 2010 16650 2030 16670
rect 2010 16490 2030 16510
rect 2090 16650 2110 16670
rect 2090 16490 2110 16510
rect 2170 16650 2190 16670
rect 2170 16490 2190 16510
rect 2250 16650 2270 16670
rect 2250 16490 2270 16510
rect 2330 16650 2350 16670
rect 2330 16490 2350 16510
rect 2410 16650 2430 16670
rect 2410 16490 2430 16510
rect 2490 16650 2510 16670
rect 2490 16490 2510 16510
rect 2570 16650 2590 16670
rect 2570 16490 2590 16510
rect 2650 16650 2670 16670
rect 2650 16490 2670 16510
rect 2730 16650 2750 16670
rect 2730 16490 2750 16510
rect 2810 16650 2830 16670
rect 2810 16490 2830 16510
rect 2890 16650 2910 16670
rect 2890 16490 2910 16510
rect 2970 16650 2990 16670
rect 2970 16490 2990 16510
rect 3050 16650 3070 16670
rect 3050 16490 3070 16510
rect 3130 16650 3150 16670
rect 3130 16490 3150 16510
rect 3210 16650 3230 16670
rect 3210 16490 3230 16510
rect 3290 16650 3310 16670
rect 3290 16490 3310 16510
rect 3370 16650 3390 16670
rect 3370 16490 3390 16510
rect 3450 16650 3470 16670
rect 3450 16490 3470 16510
rect 3530 16650 3550 16670
rect 3530 16490 3550 16510
rect 3610 16650 3630 16670
rect 3610 16490 3630 16510
rect 3690 16650 3710 16670
rect 3690 16490 3710 16510
rect 3770 16650 3790 16670
rect 3770 16490 3790 16510
rect 3850 16650 3870 16670
rect 3850 16490 3870 16510
rect 3930 16650 3950 16670
rect 3930 16490 3950 16510
rect 4010 16650 4030 16670
rect 4010 16490 4030 16510
rect 4090 16650 4110 16670
rect 4090 16490 4110 16510
rect 4170 16650 4190 16670
rect 4170 16490 4190 16510
rect 6250 16650 6270 16670
rect 6250 16490 6270 16510
rect 6330 16650 6350 16670
rect 6330 16490 6350 16510
rect 6410 16650 6430 16670
rect 6410 16490 6430 16510
rect 6490 16650 6510 16670
rect 6490 16490 6510 16510
rect 6570 16650 6590 16670
rect 6570 16490 6590 16510
rect 6650 16650 6670 16670
rect 6650 16490 6670 16510
rect 6730 16650 6750 16670
rect 6730 16490 6750 16510
rect 6810 16650 6830 16670
rect 6810 16490 6830 16510
rect 6890 16650 6910 16670
rect 6890 16490 6910 16510
rect 6970 16650 6990 16670
rect 6970 16490 6990 16510
rect 7050 16650 7070 16670
rect 7050 16490 7070 16510
rect 7130 16650 7150 16670
rect 7130 16490 7150 16510
rect 7210 16650 7230 16670
rect 7210 16490 7230 16510
rect 7290 16650 7310 16670
rect 7290 16490 7310 16510
rect 7370 16650 7390 16670
rect 7370 16490 7390 16510
rect 7450 16650 7470 16670
rect 7450 16490 7470 16510
rect 7530 16650 7550 16670
rect 7530 16490 7550 16510
rect 7610 16650 7630 16670
rect 7610 16490 7630 16510
rect 7690 16650 7710 16670
rect 7690 16490 7710 16510
rect 7770 16650 7790 16670
rect 7770 16490 7790 16510
rect 7850 16650 7870 16670
rect 7850 16490 7870 16510
rect 7930 16650 7950 16670
rect 7930 16490 7950 16510
rect 8010 16650 8030 16670
rect 8010 16490 8030 16510
rect 8090 16650 8110 16670
rect 8090 16490 8110 16510
rect 8170 16650 8190 16670
rect 8170 16490 8190 16510
rect 8250 16650 8270 16670
rect 8250 16490 8270 16510
rect 8330 16650 8350 16670
rect 8330 16490 8350 16510
rect 8410 16650 8430 16670
rect 8410 16490 8430 16510
rect 8490 16650 8510 16670
rect 8490 16490 8510 16510
rect 8570 16650 8590 16670
rect 8570 16490 8590 16510
rect 8650 16650 8670 16670
rect 8650 16490 8670 16510
rect 8730 16650 8750 16670
rect 8730 16490 8750 16510
rect 8810 16650 8830 16670
rect 8810 16490 8830 16510
rect 8890 16650 8910 16670
rect 8890 16490 8910 16510
rect 8970 16650 8990 16670
rect 8970 16490 8990 16510
rect 9050 16650 9070 16670
rect 9050 16490 9070 16510
rect 9130 16650 9150 16670
rect 9130 16490 9150 16510
rect 9210 16650 9230 16670
rect 9210 16490 9230 16510
rect 9290 16650 9310 16670
rect 9290 16490 9310 16510
rect 9370 16650 9390 16670
rect 9370 16490 9390 16510
rect 9450 16650 9470 16670
rect 9450 16490 9470 16510
rect 11570 16650 11590 16670
rect 11570 16490 11590 16510
rect 11650 16650 11670 16670
rect 11650 16490 11670 16510
rect 11730 16650 11750 16670
rect 11730 16490 11750 16510
rect 11810 16650 11830 16670
rect 11810 16490 11830 16510
rect 11890 16650 11910 16670
rect 11890 16490 11910 16510
rect 11970 16650 11990 16670
rect 11970 16490 11990 16510
rect 12050 16650 12070 16670
rect 12050 16490 12070 16510
rect 12130 16650 12150 16670
rect 12130 16490 12150 16510
rect 12210 16650 12230 16670
rect 12210 16490 12230 16510
rect 12290 16650 12310 16670
rect 12290 16490 12310 16510
rect 12370 16650 12390 16670
rect 12370 16490 12390 16510
rect 12450 16650 12470 16670
rect 12450 16490 12470 16510
rect 12530 16650 12550 16670
rect 12530 16490 12550 16510
rect 12610 16650 12630 16670
rect 12610 16490 12630 16510
rect 12690 16650 12710 16670
rect 12690 16490 12710 16510
rect 12770 16650 12790 16670
rect 12770 16490 12790 16510
rect 12850 16650 12870 16670
rect 12850 16490 12870 16510
rect 12930 16650 12950 16670
rect 12930 16490 12950 16510
rect 13010 16650 13030 16670
rect 13010 16490 13030 16510
rect 13090 16650 13110 16670
rect 13090 16490 13110 16510
rect 13170 16650 13190 16670
rect 13170 16490 13190 16510
rect 13250 16650 13270 16670
rect 13250 16490 13270 16510
rect 13330 16650 13350 16670
rect 13330 16490 13350 16510
rect 13410 16650 13430 16670
rect 13410 16490 13430 16510
rect 13490 16650 13510 16670
rect 13490 16490 13510 16510
rect 13570 16650 13590 16670
rect 13570 16490 13590 16510
rect 13650 16650 13670 16670
rect 13650 16490 13670 16510
rect 13730 16650 13750 16670
rect 13730 16490 13750 16510
rect 13810 16650 13830 16670
rect 13810 16490 13830 16510
rect 13890 16650 13910 16670
rect 13890 16490 13910 16510
rect 13970 16650 13990 16670
rect 13970 16490 13990 16510
rect 14050 16650 14070 16670
rect 14050 16490 14070 16510
rect 14130 16650 14150 16670
rect 14130 16490 14150 16510
rect 14210 16650 14230 16670
rect 14210 16490 14230 16510
rect 14290 16650 14310 16670
rect 14290 16490 14310 16510
rect 14370 16650 14390 16670
rect 14370 16490 14390 16510
rect 14450 16650 14470 16670
rect 14450 16490 14470 16510
rect 14530 16650 14550 16670
rect 14530 16490 14550 16510
rect 14610 16650 14630 16670
rect 14610 16490 14630 16510
rect 14690 16650 14710 16670
rect 14690 16490 14710 16510
rect 16770 16650 16790 16670
rect 16770 16490 16790 16510
rect 16850 16650 16870 16670
rect 16850 16490 16870 16510
rect 16930 16650 16950 16670
rect 16930 16490 16950 16510
rect 17010 16650 17030 16670
rect 17010 16490 17030 16510
rect 17090 16650 17110 16670
rect 17090 16490 17110 16510
rect 17170 16650 17190 16670
rect 17170 16490 17190 16510
rect 17250 16650 17270 16670
rect 17250 16490 17270 16510
rect 17330 16650 17350 16670
rect 17330 16490 17350 16510
rect 17410 16650 17430 16670
rect 17410 16490 17430 16510
rect 17490 16650 17510 16670
rect 17490 16490 17510 16510
rect 17570 16650 17590 16670
rect 17570 16490 17590 16510
rect 17650 16650 17670 16670
rect 17650 16490 17670 16510
rect 17730 16650 17750 16670
rect 17730 16490 17750 16510
rect 17810 16650 17830 16670
rect 17810 16490 17830 16510
rect 17890 16650 17910 16670
rect 17890 16490 17910 16510
rect 17970 16650 17990 16670
rect 17970 16490 17990 16510
rect 18050 16650 18070 16670
rect 18050 16490 18070 16510
rect 18130 16650 18150 16670
rect 18130 16490 18150 16510
rect 18210 16650 18230 16670
rect 18210 16490 18230 16510
rect 18290 16650 18310 16670
rect 18290 16490 18310 16510
rect 18370 16650 18390 16670
rect 18370 16490 18390 16510
rect 18450 16650 18470 16670
rect 18450 16490 18470 16510
rect 18530 16650 18550 16670
rect 18530 16490 18550 16510
rect 18610 16650 18630 16670
rect 18610 16490 18630 16510
rect 18690 16650 18710 16670
rect 18690 16490 18710 16510
rect 18770 16650 18790 16670
rect 18770 16490 18790 16510
rect 18850 16650 18870 16670
rect 18850 16490 18870 16510
rect 18930 16650 18950 16670
rect 18930 16490 18950 16510
rect 19010 16650 19030 16670
rect 19010 16490 19030 16510
rect 19090 16650 19110 16670
rect 19090 16490 19110 16510
rect 19170 16650 19190 16670
rect 19170 16490 19190 16510
rect 19250 16650 19270 16670
rect 19250 16490 19270 16510
rect 19330 16650 19350 16670
rect 19330 16490 19350 16510
rect 19410 16650 19430 16670
rect 19410 16490 19430 16510
rect 19490 16650 19510 16670
rect 19490 16490 19510 16510
rect 19570 16650 19590 16670
rect 19570 16490 19590 16510
rect 19650 16650 19670 16670
rect 19650 16490 19670 16510
rect 19730 16650 19750 16670
rect 19730 16490 19750 16510
rect 19810 16650 19830 16670
rect 19810 16490 19830 16510
rect 19890 16650 19910 16670
rect 19890 16490 19910 16510
rect 19970 16650 19990 16670
rect 19970 16490 19990 16510
rect 20050 16650 20070 16670
rect 20050 16490 20070 16510
rect 20130 16650 20150 16670
rect 20130 16490 20150 16510
rect 20210 16650 20230 16670
rect 20210 16490 20230 16510
rect 20290 16650 20310 16670
rect 20290 16490 20310 16510
rect 20370 16650 20390 16670
rect 20370 16490 20390 16510
rect 20450 16650 20470 16670
rect 20450 16490 20470 16510
rect 20530 16650 20550 16670
rect 20530 16490 20550 16510
rect 20610 16650 20630 16670
rect 20610 16490 20630 16510
rect 20690 16650 20710 16670
rect 20690 16490 20710 16510
rect 20770 16650 20790 16670
rect 20770 16490 20790 16510
rect 20850 16650 20870 16670
rect 20850 16490 20870 16510
rect 20930 16650 20950 16670
rect 20930 16490 20950 16510
rect 10 16410 30 16430
rect 10 16250 30 16270
rect 90 16410 110 16430
rect 90 16250 110 16270
rect 170 16410 190 16430
rect 170 16250 190 16270
rect 250 16410 270 16430
rect 250 16250 270 16270
rect 330 16410 350 16430
rect 330 16250 350 16270
rect 410 16410 430 16430
rect 410 16250 430 16270
rect 490 16410 510 16430
rect 490 16250 510 16270
rect 570 16410 590 16430
rect 570 16250 590 16270
rect 650 16410 670 16430
rect 650 16250 670 16270
rect 730 16410 750 16430
rect 730 16250 750 16270
rect 810 16410 830 16430
rect 810 16250 830 16270
rect 890 16410 910 16430
rect 890 16250 910 16270
rect 970 16410 990 16430
rect 970 16250 990 16270
rect 1050 16410 1070 16430
rect 1050 16250 1070 16270
rect 1130 16410 1150 16430
rect 1130 16250 1150 16270
rect 1210 16410 1230 16430
rect 1210 16250 1230 16270
rect 1290 16410 1310 16430
rect 1290 16250 1310 16270
rect 1370 16410 1390 16430
rect 1370 16250 1390 16270
rect 1450 16410 1470 16430
rect 1450 16250 1470 16270
rect 1530 16410 1550 16430
rect 1530 16250 1550 16270
rect 1610 16410 1630 16430
rect 1610 16250 1630 16270
rect 1690 16410 1710 16430
rect 1690 16250 1710 16270
rect 1770 16410 1790 16430
rect 1770 16250 1790 16270
rect 1850 16410 1870 16430
rect 1850 16250 1870 16270
rect 1930 16410 1950 16430
rect 1930 16250 1950 16270
rect 2010 16410 2030 16430
rect 2010 16250 2030 16270
rect 2090 16410 2110 16430
rect 2090 16250 2110 16270
rect 2170 16410 2190 16430
rect 2170 16250 2190 16270
rect 2250 16410 2270 16430
rect 2250 16250 2270 16270
rect 2330 16410 2350 16430
rect 2330 16250 2350 16270
rect 2410 16410 2430 16430
rect 2410 16250 2430 16270
rect 2490 16410 2510 16430
rect 2490 16250 2510 16270
rect 2570 16410 2590 16430
rect 2570 16250 2590 16270
rect 2650 16410 2670 16430
rect 2650 16250 2670 16270
rect 2730 16410 2750 16430
rect 2730 16250 2750 16270
rect 2810 16410 2830 16430
rect 2810 16250 2830 16270
rect 2890 16410 2910 16430
rect 2890 16250 2910 16270
rect 2970 16410 2990 16430
rect 2970 16250 2990 16270
rect 3050 16410 3070 16430
rect 3050 16250 3070 16270
rect 3130 16410 3150 16430
rect 3130 16250 3150 16270
rect 3210 16410 3230 16430
rect 3210 16250 3230 16270
rect 3290 16410 3310 16430
rect 3290 16250 3310 16270
rect 3370 16410 3390 16430
rect 3370 16250 3390 16270
rect 3450 16410 3470 16430
rect 3450 16250 3470 16270
rect 3530 16410 3550 16430
rect 3530 16250 3550 16270
rect 3610 16410 3630 16430
rect 3610 16250 3630 16270
rect 3690 16410 3710 16430
rect 3690 16250 3710 16270
rect 3770 16410 3790 16430
rect 3770 16250 3790 16270
rect 3850 16410 3870 16430
rect 3850 16250 3870 16270
rect 3930 16410 3950 16430
rect 3930 16250 3950 16270
rect 4010 16410 4030 16430
rect 4010 16250 4030 16270
rect 4090 16410 4110 16430
rect 4090 16250 4110 16270
rect 4170 16410 4190 16430
rect 4170 16250 4190 16270
rect 6250 16410 6270 16430
rect 6250 16250 6270 16270
rect 6330 16410 6350 16430
rect 6330 16250 6350 16270
rect 6410 16410 6430 16430
rect 6410 16250 6430 16270
rect 6490 16410 6510 16430
rect 6490 16250 6510 16270
rect 6570 16410 6590 16430
rect 6570 16250 6590 16270
rect 6650 16410 6670 16430
rect 6650 16250 6670 16270
rect 6730 16410 6750 16430
rect 6730 16250 6750 16270
rect 6810 16410 6830 16430
rect 6810 16250 6830 16270
rect 6890 16410 6910 16430
rect 6890 16250 6910 16270
rect 6970 16410 6990 16430
rect 6970 16250 6990 16270
rect 7050 16410 7070 16430
rect 7050 16250 7070 16270
rect 7130 16410 7150 16430
rect 7130 16250 7150 16270
rect 7210 16410 7230 16430
rect 7210 16250 7230 16270
rect 7290 16410 7310 16430
rect 7290 16250 7310 16270
rect 7370 16410 7390 16430
rect 7370 16250 7390 16270
rect 7450 16410 7470 16430
rect 7450 16250 7470 16270
rect 7530 16410 7550 16430
rect 7530 16250 7550 16270
rect 7610 16410 7630 16430
rect 7610 16250 7630 16270
rect 7690 16410 7710 16430
rect 7690 16250 7710 16270
rect 7770 16410 7790 16430
rect 7770 16250 7790 16270
rect 7850 16410 7870 16430
rect 7850 16250 7870 16270
rect 7930 16410 7950 16430
rect 7930 16250 7950 16270
rect 8010 16410 8030 16430
rect 8010 16250 8030 16270
rect 8090 16410 8110 16430
rect 8090 16250 8110 16270
rect 8170 16410 8190 16430
rect 8170 16250 8190 16270
rect 8250 16410 8270 16430
rect 8250 16250 8270 16270
rect 8330 16410 8350 16430
rect 8330 16250 8350 16270
rect 8410 16410 8430 16430
rect 8410 16250 8430 16270
rect 8490 16410 8510 16430
rect 8490 16250 8510 16270
rect 8570 16410 8590 16430
rect 8570 16250 8590 16270
rect 8650 16410 8670 16430
rect 8650 16250 8670 16270
rect 8730 16410 8750 16430
rect 8730 16250 8750 16270
rect 8810 16410 8830 16430
rect 8810 16250 8830 16270
rect 8890 16410 8910 16430
rect 8890 16250 8910 16270
rect 8970 16410 8990 16430
rect 8970 16250 8990 16270
rect 9050 16410 9070 16430
rect 9050 16250 9070 16270
rect 9130 16410 9150 16430
rect 9130 16250 9150 16270
rect 9210 16410 9230 16430
rect 9210 16250 9230 16270
rect 9290 16410 9310 16430
rect 9290 16250 9310 16270
rect 9370 16410 9390 16430
rect 9370 16250 9390 16270
rect 9450 16410 9470 16430
rect 9450 16250 9470 16270
rect 11570 16410 11590 16430
rect 11570 16250 11590 16270
rect 11650 16410 11670 16430
rect 11650 16250 11670 16270
rect 11730 16410 11750 16430
rect 11730 16250 11750 16270
rect 11810 16410 11830 16430
rect 11810 16250 11830 16270
rect 11890 16410 11910 16430
rect 11890 16250 11910 16270
rect 11970 16410 11990 16430
rect 11970 16250 11990 16270
rect 12050 16410 12070 16430
rect 12050 16250 12070 16270
rect 12130 16410 12150 16430
rect 12130 16250 12150 16270
rect 12210 16410 12230 16430
rect 12210 16250 12230 16270
rect 12290 16410 12310 16430
rect 12290 16250 12310 16270
rect 12370 16410 12390 16430
rect 12370 16250 12390 16270
rect 12450 16410 12470 16430
rect 12450 16250 12470 16270
rect 12530 16410 12550 16430
rect 12530 16250 12550 16270
rect 12610 16410 12630 16430
rect 12610 16250 12630 16270
rect 12690 16410 12710 16430
rect 12690 16250 12710 16270
rect 12770 16410 12790 16430
rect 12770 16250 12790 16270
rect 12850 16410 12870 16430
rect 12850 16250 12870 16270
rect 12930 16410 12950 16430
rect 12930 16250 12950 16270
rect 13010 16410 13030 16430
rect 13010 16250 13030 16270
rect 13090 16410 13110 16430
rect 13090 16250 13110 16270
rect 13170 16410 13190 16430
rect 13170 16250 13190 16270
rect 13250 16410 13270 16430
rect 13250 16250 13270 16270
rect 13330 16410 13350 16430
rect 13330 16250 13350 16270
rect 13410 16410 13430 16430
rect 13410 16250 13430 16270
rect 13490 16410 13510 16430
rect 13490 16250 13510 16270
rect 13570 16410 13590 16430
rect 13570 16250 13590 16270
rect 13650 16410 13670 16430
rect 13650 16250 13670 16270
rect 13730 16410 13750 16430
rect 13730 16250 13750 16270
rect 13810 16410 13830 16430
rect 13810 16250 13830 16270
rect 13890 16410 13910 16430
rect 13890 16250 13910 16270
rect 13970 16410 13990 16430
rect 13970 16250 13990 16270
rect 14050 16410 14070 16430
rect 14050 16250 14070 16270
rect 14130 16410 14150 16430
rect 14130 16250 14150 16270
rect 14210 16410 14230 16430
rect 14210 16250 14230 16270
rect 14290 16410 14310 16430
rect 14290 16250 14310 16270
rect 14370 16410 14390 16430
rect 14370 16250 14390 16270
rect 14450 16410 14470 16430
rect 14450 16250 14470 16270
rect 14530 16410 14550 16430
rect 14530 16250 14550 16270
rect 14610 16410 14630 16430
rect 14610 16250 14630 16270
rect 14690 16410 14710 16430
rect 14690 16250 14710 16270
rect 16770 16410 16790 16430
rect 16770 16250 16790 16270
rect 16850 16410 16870 16430
rect 16850 16250 16870 16270
rect 16930 16410 16950 16430
rect 16930 16250 16950 16270
rect 17010 16410 17030 16430
rect 17010 16250 17030 16270
rect 17090 16410 17110 16430
rect 17090 16250 17110 16270
rect 17170 16410 17190 16430
rect 17170 16250 17190 16270
rect 17250 16410 17270 16430
rect 17250 16250 17270 16270
rect 17330 16410 17350 16430
rect 17330 16250 17350 16270
rect 17410 16410 17430 16430
rect 17410 16250 17430 16270
rect 17490 16410 17510 16430
rect 17490 16250 17510 16270
rect 17570 16410 17590 16430
rect 17570 16250 17590 16270
rect 17650 16410 17670 16430
rect 17650 16250 17670 16270
rect 17730 16410 17750 16430
rect 17730 16250 17750 16270
rect 17810 16410 17830 16430
rect 17810 16250 17830 16270
rect 17890 16410 17910 16430
rect 17890 16250 17910 16270
rect 17970 16410 17990 16430
rect 17970 16250 17990 16270
rect 18050 16410 18070 16430
rect 18050 16250 18070 16270
rect 18130 16410 18150 16430
rect 18130 16250 18150 16270
rect 18210 16410 18230 16430
rect 18210 16250 18230 16270
rect 18290 16410 18310 16430
rect 18290 16250 18310 16270
rect 18370 16410 18390 16430
rect 18370 16250 18390 16270
rect 18450 16410 18470 16430
rect 18450 16250 18470 16270
rect 18530 16410 18550 16430
rect 18530 16250 18550 16270
rect 18610 16410 18630 16430
rect 18610 16250 18630 16270
rect 18690 16410 18710 16430
rect 18690 16250 18710 16270
rect 18770 16410 18790 16430
rect 18770 16250 18790 16270
rect 18850 16410 18870 16430
rect 18850 16250 18870 16270
rect 18930 16410 18950 16430
rect 18930 16250 18950 16270
rect 19010 16410 19030 16430
rect 19010 16250 19030 16270
rect 19090 16410 19110 16430
rect 19090 16250 19110 16270
rect 19170 16410 19190 16430
rect 19170 16250 19190 16270
rect 19250 16410 19270 16430
rect 19250 16250 19270 16270
rect 19330 16410 19350 16430
rect 19330 16250 19350 16270
rect 19410 16410 19430 16430
rect 19410 16250 19430 16270
rect 19490 16410 19510 16430
rect 19490 16250 19510 16270
rect 19570 16410 19590 16430
rect 19570 16250 19590 16270
rect 19650 16410 19670 16430
rect 19650 16250 19670 16270
rect 19730 16410 19750 16430
rect 19730 16250 19750 16270
rect 19810 16410 19830 16430
rect 19810 16250 19830 16270
rect 19890 16410 19910 16430
rect 19890 16250 19910 16270
rect 19970 16410 19990 16430
rect 19970 16250 19990 16270
rect 20050 16410 20070 16430
rect 20050 16250 20070 16270
rect 20130 16410 20150 16430
rect 20130 16250 20150 16270
rect 20210 16410 20230 16430
rect 20210 16250 20230 16270
rect 20290 16410 20310 16430
rect 20290 16250 20310 16270
rect 20370 16410 20390 16430
rect 20370 16250 20390 16270
rect 20450 16410 20470 16430
rect 20450 16250 20470 16270
rect 20530 16410 20550 16430
rect 20530 16250 20550 16270
rect 20610 16410 20630 16430
rect 20610 16250 20630 16270
rect 20690 16410 20710 16430
rect 20690 16250 20710 16270
rect 20770 16410 20790 16430
rect 20770 16250 20790 16270
rect 20850 16410 20870 16430
rect 20850 16250 20870 16270
rect 20930 16410 20950 16430
rect 20930 16250 20950 16270
rect 10 16170 30 16190
rect 10 16010 30 16030
rect 10 15850 30 15870
rect 10 15690 30 15710
rect 10 15530 30 15550
rect 10 15370 30 15390
rect 10 15210 30 15230
rect 90 16170 110 16190
rect 90 16010 110 16030
rect 90 15850 110 15870
rect 90 15690 110 15710
rect 90 15530 110 15550
rect 90 15370 110 15390
rect 90 15210 110 15230
rect 170 16170 190 16190
rect 170 16010 190 16030
rect 170 15850 190 15870
rect 170 15690 190 15710
rect 170 15530 190 15550
rect 170 15370 190 15390
rect 170 15210 190 15230
rect 250 16170 270 16190
rect 250 16010 270 16030
rect 250 15850 270 15870
rect 250 15690 270 15710
rect 250 15530 270 15550
rect 250 15370 270 15390
rect 250 15210 270 15230
rect 330 16170 350 16190
rect 330 16010 350 16030
rect 330 15850 350 15870
rect 330 15690 350 15710
rect 330 15530 350 15550
rect 330 15370 350 15390
rect 330 15210 350 15230
rect 410 16170 430 16190
rect 410 16010 430 16030
rect 410 15850 430 15870
rect 410 15690 430 15710
rect 410 15530 430 15550
rect 410 15370 430 15390
rect 410 15210 430 15230
rect 490 16170 510 16190
rect 490 16010 510 16030
rect 490 15850 510 15870
rect 490 15690 510 15710
rect 490 15530 510 15550
rect 490 15370 510 15390
rect 490 15210 510 15230
rect 570 16170 590 16190
rect 570 16010 590 16030
rect 570 15850 590 15870
rect 570 15690 590 15710
rect 570 15530 590 15550
rect 570 15370 590 15390
rect 570 15210 590 15230
rect 650 16170 670 16190
rect 650 16010 670 16030
rect 650 15850 670 15870
rect 650 15690 670 15710
rect 650 15530 670 15550
rect 650 15370 670 15390
rect 650 15210 670 15230
rect 730 16170 750 16190
rect 730 16010 750 16030
rect 730 15850 750 15870
rect 730 15690 750 15710
rect 730 15530 750 15550
rect 730 15370 750 15390
rect 730 15210 750 15230
rect 810 16170 830 16190
rect 810 16010 830 16030
rect 810 15850 830 15870
rect 810 15690 830 15710
rect 810 15530 830 15550
rect 810 15370 830 15390
rect 810 15210 830 15230
rect 890 16170 910 16190
rect 890 16010 910 16030
rect 890 15850 910 15870
rect 890 15690 910 15710
rect 890 15530 910 15550
rect 890 15370 910 15390
rect 890 15210 910 15230
rect 970 16170 990 16190
rect 970 16010 990 16030
rect 970 15850 990 15870
rect 970 15690 990 15710
rect 970 15530 990 15550
rect 970 15370 990 15390
rect 970 15210 990 15230
rect 1050 16170 1070 16190
rect 1050 16010 1070 16030
rect 1050 15850 1070 15870
rect 1050 15690 1070 15710
rect 1050 15530 1070 15550
rect 1050 15370 1070 15390
rect 1050 15210 1070 15230
rect 1130 16170 1150 16190
rect 1130 16010 1150 16030
rect 1130 15850 1150 15870
rect 1130 15690 1150 15710
rect 1130 15530 1150 15550
rect 1130 15370 1150 15390
rect 1130 15210 1150 15230
rect 1210 16170 1230 16190
rect 1210 16010 1230 16030
rect 1210 15850 1230 15870
rect 1210 15690 1230 15710
rect 1210 15530 1230 15550
rect 1210 15370 1230 15390
rect 1210 15210 1230 15230
rect 1290 16170 1310 16190
rect 1290 16010 1310 16030
rect 1290 15850 1310 15870
rect 1290 15690 1310 15710
rect 1290 15530 1310 15550
rect 1290 15370 1310 15390
rect 1290 15210 1310 15230
rect 1370 16170 1390 16190
rect 1370 16010 1390 16030
rect 1370 15850 1390 15870
rect 1370 15690 1390 15710
rect 1370 15530 1390 15550
rect 1370 15370 1390 15390
rect 1370 15210 1390 15230
rect 1450 16170 1470 16190
rect 1450 16010 1470 16030
rect 1450 15850 1470 15870
rect 1450 15690 1470 15710
rect 1450 15530 1470 15550
rect 1450 15370 1470 15390
rect 1450 15210 1470 15230
rect 1530 16170 1550 16190
rect 1530 16010 1550 16030
rect 1530 15850 1550 15870
rect 1530 15690 1550 15710
rect 1530 15530 1550 15550
rect 1530 15370 1550 15390
rect 1530 15210 1550 15230
rect 1610 16170 1630 16190
rect 1610 16010 1630 16030
rect 1610 15850 1630 15870
rect 1610 15690 1630 15710
rect 1610 15530 1630 15550
rect 1610 15370 1630 15390
rect 1610 15210 1630 15230
rect 1690 16170 1710 16190
rect 1690 16010 1710 16030
rect 1690 15850 1710 15870
rect 1690 15690 1710 15710
rect 1690 15530 1710 15550
rect 1690 15370 1710 15390
rect 1690 15210 1710 15230
rect 1770 16170 1790 16190
rect 1770 16010 1790 16030
rect 1770 15850 1790 15870
rect 1770 15690 1790 15710
rect 1770 15530 1790 15550
rect 1770 15370 1790 15390
rect 1770 15210 1790 15230
rect 1850 16170 1870 16190
rect 1850 16010 1870 16030
rect 1850 15850 1870 15870
rect 1850 15690 1870 15710
rect 1850 15530 1870 15550
rect 1850 15370 1870 15390
rect 1850 15210 1870 15230
rect 1930 16170 1950 16190
rect 1930 16010 1950 16030
rect 1930 15850 1950 15870
rect 1930 15690 1950 15710
rect 1930 15530 1950 15550
rect 1930 15370 1950 15390
rect 1930 15210 1950 15230
rect 2010 16170 2030 16190
rect 2010 16010 2030 16030
rect 2010 15850 2030 15870
rect 2010 15690 2030 15710
rect 2010 15530 2030 15550
rect 2010 15370 2030 15390
rect 2010 15210 2030 15230
rect 2090 16170 2110 16190
rect 2090 16010 2110 16030
rect 2090 15850 2110 15870
rect 2090 15690 2110 15710
rect 2090 15530 2110 15550
rect 2090 15370 2110 15390
rect 2090 15210 2110 15230
rect 2170 16170 2190 16190
rect 2170 16010 2190 16030
rect 2170 15850 2190 15870
rect 2170 15690 2190 15710
rect 2170 15530 2190 15550
rect 2170 15370 2190 15390
rect 2170 15210 2190 15230
rect 2250 16170 2270 16190
rect 2250 16010 2270 16030
rect 2250 15850 2270 15870
rect 2250 15690 2270 15710
rect 2250 15530 2270 15550
rect 2250 15370 2270 15390
rect 2250 15210 2270 15230
rect 2330 16170 2350 16190
rect 2330 16010 2350 16030
rect 2330 15850 2350 15870
rect 2330 15690 2350 15710
rect 2330 15530 2350 15550
rect 2330 15370 2350 15390
rect 2330 15210 2350 15230
rect 2410 16170 2430 16190
rect 2410 16010 2430 16030
rect 2410 15850 2430 15870
rect 2410 15690 2430 15710
rect 2410 15530 2430 15550
rect 2410 15370 2430 15390
rect 2410 15210 2430 15230
rect 2490 16170 2510 16190
rect 2490 16010 2510 16030
rect 2490 15850 2510 15870
rect 2490 15690 2510 15710
rect 2490 15530 2510 15550
rect 2490 15370 2510 15390
rect 2490 15210 2510 15230
rect 2570 16170 2590 16190
rect 2570 16010 2590 16030
rect 2570 15850 2590 15870
rect 2570 15690 2590 15710
rect 2570 15530 2590 15550
rect 2570 15370 2590 15390
rect 2570 15210 2590 15230
rect 2650 16170 2670 16190
rect 2650 16010 2670 16030
rect 2650 15850 2670 15870
rect 2650 15690 2670 15710
rect 2650 15530 2670 15550
rect 2650 15370 2670 15390
rect 2650 15210 2670 15230
rect 2730 16170 2750 16190
rect 2730 16010 2750 16030
rect 2730 15850 2750 15870
rect 2730 15690 2750 15710
rect 2730 15530 2750 15550
rect 2730 15370 2750 15390
rect 2730 15210 2750 15230
rect 2810 16170 2830 16190
rect 2810 16010 2830 16030
rect 2810 15850 2830 15870
rect 2810 15690 2830 15710
rect 2810 15530 2830 15550
rect 2810 15370 2830 15390
rect 2810 15210 2830 15230
rect 2890 16170 2910 16190
rect 2890 16010 2910 16030
rect 2890 15850 2910 15870
rect 2890 15690 2910 15710
rect 2890 15530 2910 15550
rect 2890 15370 2910 15390
rect 2890 15210 2910 15230
rect 2970 16170 2990 16190
rect 2970 16010 2990 16030
rect 2970 15850 2990 15870
rect 2970 15690 2990 15710
rect 2970 15530 2990 15550
rect 2970 15370 2990 15390
rect 2970 15210 2990 15230
rect 3050 16170 3070 16190
rect 3050 16010 3070 16030
rect 3050 15850 3070 15870
rect 3050 15690 3070 15710
rect 3050 15530 3070 15550
rect 3050 15370 3070 15390
rect 3050 15210 3070 15230
rect 3130 16170 3150 16190
rect 3130 16010 3150 16030
rect 3130 15850 3150 15870
rect 3130 15690 3150 15710
rect 3130 15530 3150 15550
rect 3130 15370 3150 15390
rect 3130 15210 3150 15230
rect 3210 16170 3230 16190
rect 3210 16010 3230 16030
rect 3210 15850 3230 15870
rect 3210 15690 3230 15710
rect 3210 15530 3230 15550
rect 3210 15370 3230 15390
rect 3210 15210 3230 15230
rect 3290 16170 3310 16190
rect 3290 16010 3310 16030
rect 3290 15850 3310 15870
rect 3290 15690 3310 15710
rect 3290 15530 3310 15550
rect 3290 15370 3310 15390
rect 3290 15210 3310 15230
rect 3370 16170 3390 16190
rect 3370 16010 3390 16030
rect 3370 15850 3390 15870
rect 3370 15690 3390 15710
rect 3370 15530 3390 15550
rect 3370 15370 3390 15390
rect 3370 15210 3390 15230
rect 3450 16170 3470 16190
rect 3450 16010 3470 16030
rect 3450 15850 3470 15870
rect 3450 15690 3470 15710
rect 3450 15530 3470 15550
rect 3450 15370 3470 15390
rect 3450 15210 3470 15230
rect 3530 16170 3550 16190
rect 3530 16010 3550 16030
rect 3530 15850 3550 15870
rect 3530 15690 3550 15710
rect 3530 15530 3550 15550
rect 3530 15370 3550 15390
rect 3530 15210 3550 15230
rect 3610 16170 3630 16190
rect 3610 16010 3630 16030
rect 3610 15850 3630 15870
rect 3610 15690 3630 15710
rect 3610 15530 3630 15550
rect 3610 15370 3630 15390
rect 3610 15210 3630 15230
rect 3690 16170 3710 16190
rect 3690 16010 3710 16030
rect 3690 15850 3710 15870
rect 3690 15690 3710 15710
rect 3690 15530 3710 15550
rect 3690 15370 3710 15390
rect 3690 15210 3710 15230
rect 3770 16170 3790 16190
rect 3770 16010 3790 16030
rect 3770 15850 3790 15870
rect 3770 15690 3790 15710
rect 3770 15530 3790 15550
rect 3770 15370 3790 15390
rect 3770 15210 3790 15230
rect 3850 16170 3870 16190
rect 3850 16010 3870 16030
rect 3850 15850 3870 15870
rect 3850 15690 3870 15710
rect 3850 15530 3870 15550
rect 3850 15370 3870 15390
rect 3850 15210 3870 15230
rect 3930 16170 3950 16190
rect 3930 16010 3950 16030
rect 3930 15850 3950 15870
rect 3930 15690 3950 15710
rect 3930 15530 3950 15550
rect 3930 15370 3950 15390
rect 3930 15210 3950 15230
rect 4010 16170 4030 16190
rect 4010 16010 4030 16030
rect 4010 15850 4030 15870
rect 4010 15690 4030 15710
rect 4010 15530 4030 15550
rect 4010 15370 4030 15390
rect 4010 15210 4030 15230
rect 4090 16170 4110 16190
rect 4090 16010 4110 16030
rect 4090 15850 4110 15870
rect 4090 15690 4110 15710
rect 4090 15530 4110 15550
rect 4090 15370 4110 15390
rect 4090 15210 4110 15230
rect 4170 16170 4190 16190
rect 4170 16010 4190 16030
rect 4170 15850 4190 15870
rect 4170 15690 4190 15710
rect 4170 15530 4190 15550
rect 4170 15370 4190 15390
rect 4170 15210 4190 15230
rect 6250 16170 6270 16190
rect 6250 16010 6270 16030
rect 6250 15850 6270 15870
rect 6250 15690 6270 15710
rect 6250 15530 6270 15550
rect 6250 15370 6270 15390
rect 6250 15210 6270 15230
rect 6330 16170 6350 16190
rect 6330 16010 6350 16030
rect 6330 15850 6350 15870
rect 6330 15690 6350 15710
rect 6330 15530 6350 15550
rect 6330 15370 6350 15390
rect 6330 15210 6350 15230
rect 6410 16170 6430 16190
rect 6410 16010 6430 16030
rect 6410 15850 6430 15870
rect 6410 15690 6430 15710
rect 6410 15530 6430 15550
rect 6410 15370 6430 15390
rect 6410 15210 6430 15230
rect 6490 16170 6510 16190
rect 6490 16010 6510 16030
rect 6490 15850 6510 15870
rect 6490 15690 6510 15710
rect 6490 15530 6510 15550
rect 6490 15370 6510 15390
rect 6490 15210 6510 15230
rect 6570 16170 6590 16190
rect 6570 16010 6590 16030
rect 6570 15850 6590 15870
rect 6570 15690 6590 15710
rect 6570 15530 6590 15550
rect 6570 15370 6590 15390
rect 6570 15210 6590 15230
rect 6650 16170 6670 16190
rect 6650 16010 6670 16030
rect 6650 15850 6670 15870
rect 6650 15690 6670 15710
rect 6650 15530 6670 15550
rect 6650 15370 6670 15390
rect 6650 15210 6670 15230
rect 6730 16170 6750 16190
rect 6730 16010 6750 16030
rect 6730 15850 6750 15870
rect 6730 15690 6750 15710
rect 6730 15530 6750 15550
rect 6730 15370 6750 15390
rect 6730 15210 6750 15230
rect 6810 16170 6830 16190
rect 6810 16010 6830 16030
rect 6810 15850 6830 15870
rect 6810 15690 6830 15710
rect 6810 15530 6830 15550
rect 6810 15370 6830 15390
rect 6810 15210 6830 15230
rect 6890 16170 6910 16190
rect 6890 16010 6910 16030
rect 6890 15850 6910 15870
rect 6890 15690 6910 15710
rect 6890 15530 6910 15550
rect 6890 15370 6910 15390
rect 6890 15210 6910 15230
rect 6970 16170 6990 16190
rect 6970 16010 6990 16030
rect 6970 15850 6990 15870
rect 6970 15690 6990 15710
rect 6970 15530 6990 15550
rect 6970 15370 6990 15390
rect 6970 15210 6990 15230
rect 7050 16170 7070 16190
rect 7050 16010 7070 16030
rect 7050 15850 7070 15870
rect 7050 15690 7070 15710
rect 7050 15530 7070 15550
rect 7050 15370 7070 15390
rect 7050 15210 7070 15230
rect 7130 16170 7150 16190
rect 7130 16010 7150 16030
rect 7130 15850 7150 15870
rect 7130 15690 7150 15710
rect 7130 15530 7150 15550
rect 7130 15370 7150 15390
rect 7130 15210 7150 15230
rect 7210 16170 7230 16190
rect 7210 16010 7230 16030
rect 7210 15850 7230 15870
rect 7210 15690 7230 15710
rect 7210 15530 7230 15550
rect 7210 15370 7230 15390
rect 7210 15210 7230 15230
rect 7290 16170 7310 16190
rect 7290 16010 7310 16030
rect 7290 15850 7310 15870
rect 7290 15690 7310 15710
rect 7290 15530 7310 15550
rect 7290 15370 7310 15390
rect 7290 15210 7310 15230
rect 7370 16170 7390 16190
rect 7370 16010 7390 16030
rect 7370 15850 7390 15870
rect 7370 15690 7390 15710
rect 7370 15530 7390 15550
rect 7370 15370 7390 15390
rect 7370 15210 7390 15230
rect 7450 16170 7470 16190
rect 7450 16010 7470 16030
rect 7450 15850 7470 15870
rect 7450 15690 7470 15710
rect 7450 15530 7470 15550
rect 7450 15370 7470 15390
rect 7450 15210 7470 15230
rect 7530 16170 7550 16190
rect 7530 16010 7550 16030
rect 7530 15850 7550 15870
rect 7530 15690 7550 15710
rect 7530 15530 7550 15550
rect 7530 15370 7550 15390
rect 7530 15210 7550 15230
rect 7610 16170 7630 16190
rect 7610 16010 7630 16030
rect 7610 15850 7630 15870
rect 7610 15690 7630 15710
rect 7610 15530 7630 15550
rect 7610 15370 7630 15390
rect 7610 15210 7630 15230
rect 7690 16170 7710 16190
rect 7690 16010 7710 16030
rect 7690 15850 7710 15870
rect 7690 15690 7710 15710
rect 7690 15530 7710 15550
rect 7690 15370 7710 15390
rect 7690 15210 7710 15230
rect 7770 16170 7790 16190
rect 7770 16010 7790 16030
rect 7770 15850 7790 15870
rect 7770 15690 7790 15710
rect 7770 15530 7790 15550
rect 7770 15370 7790 15390
rect 7770 15210 7790 15230
rect 7850 16170 7870 16190
rect 7850 16010 7870 16030
rect 7850 15850 7870 15870
rect 7850 15690 7870 15710
rect 7850 15530 7870 15550
rect 7850 15370 7870 15390
rect 7850 15210 7870 15230
rect 7930 16170 7950 16190
rect 7930 16010 7950 16030
rect 7930 15850 7950 15870
rect 7930 15690 7950 15710
rect 7930 15530 7950 15550
rect 7930 15370 7950 15390
rect 7930 15210 7950 15230
rect 8010 16170 8030 16190
rect 8010 16010 8030 16030
rect 8010 15850 8030 15870
rect 8010 15690 8030 15710
rect 8010 15530 8030 15550
rect 8010 15370 8030 15390
rect 8010 15210 8030 15230
rect 8090 16170 8110 16190
rect 8090 16010 8110 16030
rect 8090 15850 8110 15870
rect 8090 15690 8110 15710
rect 8090 15530 8110 15550
rect 8090 15370 8110 15390
rect 8090 15210 8110 15230
rect 8170 16170 8190 16190
rect 8170 16010 8190 16030
rect 8170 15850 8190 15870
rect 8170 15690 8190 15710
rect 8170 15530 8190 15550
rect 8170 15370 8190 15390
rect 8170 15210 8190 15230
rect 8250 16170 8270 16190
rect 8250 16010 8270 16030
rect 8250 15850 8270 15870
rect 8250 15690 8270 15710
rect 8250 15530 8270 15550
rect 8250 15370 8270 15390
rect 8250 15210 8270 15230
rect 8330 16170 8350 16190
rect 8330 16010 8350 16030
rect 8330 15850 8350 15870
rect 8330 15690 8350 15710
rect 8330 15530 8350 15550
rect 8330 15370 8350 15390
rect 8330 15210 8350 15230
rect 8410 16170 8430 16190
rect 8410 16010 8430 16030
rect 8410 15850 8430 15870
rect 8410 15690 8430 15710
rect 8410 15530 8430 15550
rect 8410 15370 8430 15390
rect 8410 15210 8430 15230
rect 8490 16170 8510 16190
rect 8490 16010 8510 16030
rect 8490 15850 8510 15870
rect 8490 15690 8510 15710
rect 8490 15530 8510 15550
rect 8490 15370 8510 15390
rect 8490 15210 8510 15230
rect 8570 16170 8590 16190
rect 8570 16010 8590 16030
rect 8570 15850 8590 15870
rect 8570 15690 8590 15710
rect 8570 15530 8590 15550
rect 8570 15370 8590 15390
rect 8570 15210 8590 15230
rect 8650 16170 8670 16190
rect 8650 16010 8670 16030
rect 8650 15850 8670 15870
rect 8650 15690 8670 15710
rect 8650 15530 8670 15550
rect 8650 15370 8670 15390
rect 8650 15210 8670 15230
rect 8730 16170 8750 16190
rect 8730 16010 8750 16030
rect 8730 15850 8750 15870
rect 8730 15690 8750 15710
rect 8730 15530 8750 15550
rect 8730 15370 8750 15390
rect 8730 15210 8750 15230
rect 8810 16170 8830 16190
rect 8810 16010 8830 16030
rect 8810 15850 8830 15870
rect 8810 15690 8830 15710
rect 8810 15530 8830 15550
rect 8810 15370 8830 15390
rect 8810 15210 8830 15230
rect 8890 16170 8910 16190
rect 8890 16010 8910 16030
rect 8890 15850 8910 15870
rect 8890 15690 8910 15710
rect 8890 15530 8910 15550
rect 8890 15370 8910 15390
rect 8890 15210 8910 15230
rect 8970 16170 8990 16190
rect 8970 16010 8990 16030
rect 8970 15850 8990 15870
rect 8970 15690 8990 15710
rect 8970 15530 8990 15550
rect 8970 15370 8990 15390
rect 8970 15210 8990 15230
rect 9050 16170 9070 16190
rect 9050 16010 9070 16030
rect 9050 15850 9070 15870
rect 9050 15690 9070 15710
rect 9050 15530 9070 15550
rect 9050 15370 9070 15390
rect 9050 15210 9070 15230
rect 9130 16170 9150 16190
rect 9130 16010 9150 16030
rect 9130 15850 9150 15870
rect 9130 15690 9150 15710
rect 9130 15530 9150 15550
rect 9130 15370 9150 15390
rect 9130 15210 9150 15230
rect 9210 16170 9230 16190
rect 9210 16010 9230 16030
rect 9210 15850 9230 15870
rect 9210 15690 9230 15710
rect 9210 15530 9230 15550
rect 9210 15370 9230 15390
rect 9210 15210 9230 15230
rect 9290 16170 9310 16190
rect 9290 16010 9310 16030
rect 9290 15850 9310 15870
rect 9290 15690 9310 15710
rect 9290 15530 9310 15550
rect 9290 15370 9310 15390
rect 9290 15210 9310 15230
rect 9370 16170 9390 16190
rect 9370 16010 9390 16030
rect 9370 15850 9390 15870
rect 9370 15690 9390 15710
rect 9370 15530 9390 15550
rect 9370 15370 9390 15390
rect 9370 15210 9390 15230
rect 9450 16170 9470 16190
rect 9450 16010 9470 16030
rect 9450 15850 9470 15870
rect 9450 15690 9470 15710
rect 9450 15530 9470 15550
rect 9450 15370 9470 15390
rect 9450 15210 9470 15230
rect 11570 16170 11590 16190
rect 11570 16010 11590 16030
rect 11570 15850 11590 15870
rect 11570 15690 11590 15710
rect 11570 15530 11590 15550
rect 11570 15370 11590 15390
rect 11570 15210 11590 15230
rect 11650 16170 11670 16190
rect 11650 16010 11670 16030
rect 11650 15850 11670 15870
rect 11650 15690 11670 15710
rect 11650 15530 11670 15550
rect 11650 15370 11670 15390
rect 11650 15210 11670 15230
rect 11730 16170 11750 16190
rect 11730 16010 11750 16030
rect 11730 15850 11750 15870
rect 11730 15690 11750 15710
rect 11730 15530 11750 15550
rect 11730 15370 11750 15390
rect 11730 15210 11750 15230
rect 11810 16170 11830 16190
rect 11810 16010 11830 16030
rect 11810 15850 11830 15870
rect 11810 15690 11830 15710
rect 11810 15530 11830 15550
rect 11810 15370 11830 15390
rect 11810 15210 11830 15230
rect 11890 16170 11910 16190
rect 11890 16010 11910 16030
rect 11890 15850 11910 15870
rect 11890 15690 11910 15710
rect 11890 15530 11910 15550
rect 11890 15370 11910 15390
rect 11890 15210 11910 15230
rect 11970 16170 11990 16190
rect 11970 16010 11990 16030
rect 11970 15850 11990 15870
rect 11970 15690 11990 15710
rect 11970 15530 11990 15550
rect 11970 15370 11990 15390
rect 11970 15210 11990 15230
rect 12050 16170 12070 16190
rect 12050 16010 12070 16030
rect 12050 15850 12070 15870
rect 12050 15690 12070 15710
rect 12050 15530 12070 15550
rect 12050 15370 12070 15390
rect 12050 15210 12070 15230
rect 12130 16170 12150 16190
rect 12130 16010 12150 16030
rect 12130 15850 12150 15870
rect 12130 15690 12150 15710
rect 12130 15530 12150 15550
rect 12130 15370 12150 15390
rect 12130 15210 12150 15230
rect 12210 16170 12230 16190
rect 12210 16010 12230 16030
rect 12210 15850 12230 15870
rect 12210 15690 12230 15710
rect 12210 15530 12230 15550
rect 12210 15370 12230 15390
rect 12210 15210 12230 15230
rect 12290 16170 12310 16190
rect 12290 16010 12310 16030
rect 12290 15850 12310 15870
rect 12290 15690 12310 15710
rect 12290 15530 12310 15550
rect 12290 15370 12310 15390
rect 12290 15210 12310 15230
rect 12370 16170 12390 16190
rect 12370 16010 12390 16030
rect 12370 15850 12390 15870
rect 12370 15690 12390 15710
rect 12370 15530 12390 15550
rect 12370 15370 12390 15390
rect 12370 15210 12390 15230
rect 12450 16170 12470 16190
rect 12450 16010 12470 16030
rect 12450 15850 12470 15870
rect 12450 15690 12470 15710
rect 12450 15530 12470 15550
rect 12450 15370 12470 15390
rect 12450 15210 12470 15230
rect 12530 16170 12550 16190
rect 12530 16010 12550 16030
rect 12530 15850 12550 15870
rect 12530 15690 12550 15710
rect 12530 15530 12550 15550
rect 12530 15370 12550 15390
rect 12530 15210 12550 15230
rect 12610 16170 12630 16190
rect 12610 16010 12630 16030
rect 12610 15850 12630 15870
rect 12610 15690 12630 15710
rect 12610 15530 12630 15550
rect 12610 15370 12630 15390
rect 12610 15210 12630 15230
rect 12690 16170 12710 16190
rect 12690 16010 12710 16030
rect 12690 15850 12710 15870
rect 12690 15690 12710 15710
rect 12690 15530 12710 15550
rect 12690 15370 12710 15390
rect 12690 15210 12710 15230
rect 12770 16170 12790 16190
rect 12770 16010 12790 16030
rect 12770 15850 12790 15870
rect 12770 15690 12790 15710
rect 12770 15530 12790 15550
rect 12770 15370 12790 15390
rect 12770 15210 12790 15230
rect 12850 16170 12870 16190
rect 12850 16010 12870 16030
rect 12850 15850 12870 15870
rect 12850 15690 12870 15710
rect 12850 15530 12870 15550
rect 12850 15370 12870 15390
rect 12850 15210 12870 15230
rect 12930 16170 12950 16190
rect 12930 16010 12950 16030
rect 12930 15850 12950 15870
rect 12930 15690 12950 15710
rect 12930 15530 12950 15550
rect 12930 15370 12950 15390
rect 12930 15210 12950 15230
rect 13010 16170 13030 16190
rect 13010 16010 13030 16030
rect 13010 15850 13030 15870
rect 13010 15690 13030 15710
rect 13010 15530 13030 15550
rect 13010 15370 13030 15390
rect 13010 15210 13030 15230
rect 13090 16170 13110 16190
rect 13090 16010 13110 16030
rect 13090 15850 13110 15870
rect 13090 15690 13110 15710
rect 13090 15530 13110 15550
rect 13090 15370 13110 15390
rect 13090 15210 13110 15230
rect 13170 16170 13190 16190
rect 13170 16010 13190 16030
rect 13170 15850 13190 15870
rect 13170 15690 13190 15710
rect 13170 15530 13190 15550
rect 13170 15370 13190 15390
rect 13170 15210 13190 15230
rect 13250 16170 13270 16190
rect 13250 16010 13270 16030
rect 13250 15850 13270 15870
rect 13250 15690 13270 15710
rect 13250 15530 13270 15550
rect 13250 15370 13270 15390
rect 13250 15210 13270 15230
rect 13330 16170 13350 16190
rect 13330 16010 13350 16030
rect 13330 15850 13350 15870
rect 13330 15690 13350 15710
rect 13330 15530 13350 15550
rect 13330 15370 13350 15390
rect 13330 15210 13350 15230
rect 13410 16170 13430 16190
rect 13410 16010 13430 16030
rect 13410 15850 13430 15870
rect 13410 15690 13430 15710
rect 13410 15530 13430 15550
rect 13410 15370 13430 15390
rect 13410 15210 13430 15230
rect 13490 16170 13510 16190
rect 13490 16010 13510 16030
rect 13490 15850 13510 15870
rect 13490 15690 13510 15710
rect 13490 15530 13510 15550
rect 13490 15370 13510 15390
rect 13490 15210 13510 15230
rect 13570 16170 13590 16190
rect 13570 16010 13590 16030
rect 13570 15850 13590 15870
rect 13570 15690 13590 15710
rect 13570 15530 13590 15550
rect 13570 15370 13590 15390
rect 13570 15210 13590 15230
rect 13650 16170 13670 16190
rect 13650 16010 13670 16030
rect 13650 15850 13670 15870
rect 13650 15690 13670 15710
rect 13650 15530 13670 15550
rect 13650 15370 13670 15390
rect 13650 15210 13670 15230
rect 13730 16170 13750 16190
rect 13730 16010 13750 16030
rect 13730 15850 13750 15870
rect 13730 15690 13750 15710
rect 13730 15530 13750 15550
rect 13730 15370 13750 15390
rect 13730 15210 13750 15230
rect 13810 16170 13830 16190
rect 13810 16010 13830 16030
rect 13810 15850 13830 15870
rect 13810 15690 13830 15710
rect 13810 15530 13830 15550
rect 13810 15370 13830 15390
rect 13810 15210 13830 15230
rect 13890 16170 13910 16190
rect 13890 16010 13910 16030
rect 13890 15850 13910 15870
rect 13890 15690 13910 15710
rect 13890 15530 13910 15550
rect 13890 15370 13910 15390
rect 13890 15210 13910 15230
rect 13970 16170 13990 16190
rect 13970 16010 13990 16030
rect 13970 15850 13990 15870
rect 13970 15690 13990 15710
rect 13970 15530 13990 15550
rect 13970 15370 13990 15390
rect 13970 15210 13990 15230
rect 14050 16170 14070 16190
rect 14050 16010 14070 16030
rect 14050 15850 14070 15870
rect 14050 15690 14070 15710
rect 14050 15530 14070 15550
rect 14050 15370 14070 15390
rect 14050 15210 14070 15230
rect 14130 16170 14150 16190
rect 14130 16010 14150 16030
rect 14130 15850 14150 15870
rect 14130 15690 14150 15710
rect 14130 15530 14150 15550
rect 14130 15370 14150 15390
rect 14130 15210 14150 15230
rect 14210 16170 14230 16190
rect 14210 16010 14230 16030
rect 14210 15850 14230 15870
rect 14210 15690 14230 15710
rect 14210 15530 14230 15550
rect 14210 15370 14230 15390
rect 14210 15210 14230 15230
rect 14290 16170 14310 16190
rect 14290 16010 14310 16030
rect 14290 15850 14310 15870
rect 14290 15690 14310 15710
rect 14290 15530 14310 15550
rect 14290 15370 14310 15390
rect 14290 15210 14310 15230
rect 14370 16170 14390 16190
rect 14370 16010 14390 16030
rect 14370 15850 14390 15870
rect 14370 15690 14390 15710
rect 14370 15530 14390 15550
rect 14370 15370 14390 15390
rect 14370 15210 14390 15230
rect 14450 16170 14470 16190
rect 14450 16010 14470 16030
rect 14450 15850 14470 15870
rect 14450 15690 14470 15710
rect 14450 15530 14470 15550
rect 14450 15370 14470 15390
rect 14450 15210 14470 15230
rect 14530 16170 14550 16190
rect 14530 16010 14550 16030
rect 14530 15850 14550 15870
rect 14530 15690 14550 15710
rect 14530 15530 14550 15550
rect 14530 15370 14550 15390
rect 14530 15210 14550 15230
rect 14610 16170 14630 16190
rect 14610 16010 14630 16030
rect 14610 15850 14630 15870
rect 14610 15690 14630 15710
rect 14610 15530 14630 15550
rect 14610 15370 14630 15390
rect 14610 15210 14630 15230
rect 14690 16170 14710 16190
rect 14690 16010 14710 16030
rect 14690 15850 14710 15870
rect 14690 15690 14710 15710
rect 14690 15530 14710 15550
rect 14690 15370 14710 15390
rect 14690 15210 14710 15230
rect 16770 16170 16790 16190
rect 16770 16010 16790 16030
rect 16770 15850 16790 15870
rect 16770 15690 16790 15710
rect 16770 15530 16790 15550
rect 16770 15370 16790 15390
rect 16770 15210 16790 15230
rect 16850 16170 16870 16190
rect 16850 16010 16870 16030
rect 16850 15850 16870 15870
rect 16850 15690 16870 15710
rect 16850 15530 16870 15550
rect 16850 15370 16870 15390
rect 16850 15210 16870 15230
rect 16930 16170 16950 16190
rect 16930 16010 16950 16030
rect 16930 15850 16950 15870
rect 16930 15690 16950 15710
rect 16930 15530 16950 15550
rect 16930 15370 16950 15390
rect 16930 15210 16950 15230
rect 17010 16170 17030 16190
rect 17010 16010 17030 16030
rect 17010 15850 17030 15870
rect 17010 15690 17030 15710
rect 17010 15530 17030 15550
rect 17010 15370 17030 15390
rect 17010 15210 17030 15230
rect 17090 16170 17110 16190
rect 17090 16010 17110 16030
rect 17090 15850 17110 15870
rect 17090 15690 17110 15710
rect 17090 15530 17110 15550
rect 17090 15370 17110 15390
rect 17090 15210 17110 15230
rect 17170 16170 17190 16190
rect 17170 16010 17190 16030
rect 17170 15850 17190 15870
rect 17170 15690 17190 15710
rect 17170 15530 17190 15550
rect 17170 15370 17190 15390
rect 17170 15210 17190 15230
rect 17250 16170 17270 16190
rect 17250 16010 17270 16030
rect 17250 15850 17270 15870
rect 17250 15690 17270 15710
rect 17250 15530 17270 15550
rect 17250 15370 17270 15390
rect 17250 15210 17270 15230
rect 17330 16170 17350 16190
rect 17330 16010 17350 16030
rect 17330 15850 17350 15870
rect 17330 15690 17350 15710
rect 17330 15530 17350 15550
rect 17330 15370 17350 15390
rect 17330 15210 17350 15230
rect 17410 16170 17430 16190
rect 17410 16010 17430 16030
rect 17410 15850 17430 15870
rect 17410 15690 17430 15710
rect 17410 15530 17430 15550
rect 17410 15370 17430 15390
rect 17410 15210 17430 15230
rect 17490 16170 17510 16190
rect 17490 16010 17510 16030
rect 17490 15850 17510 15870
rect 17490 15690 17510 15710
rect 17490 15530 17510 15550
rect 17490 15370 17510 15390
rect 17490 15210 17510 15230
rect 17570 16170 17590 16190
rect 17570 16010 17590 16030
rect 17570 15850 17590 15870
rect 17570 15690 17590 15710
rect 17570 15530 17590 15550
rect 17570 15370 17590 15390
rect 17570 15210 17590 15230
rect 17650 16170 17670 16190
rect 17650 16010 17670 16030
rect 17650 15850 17670 15870
rect 17650 15690 17670 15710
rect 17650 15530 17670 15550
rect 17650 15370 17670 15390
rect 17650 15210 17670 15230
rect 17730 16170 17750 16190
rect 17730 16010 17750 16030
rect 17730 15850 17750 15870
rect 17730 15690 17750 15710
rect 17730 15530 17750 15550
rect 17730 15370 17750 15390
rect 17730 15210 17750 15230
rect 17810 16170 17830 16190
rect 17810 16010 17830 16030
rect 17810 15850 17830 15870
rect 17810 15690 17830 15710
rect 17810 15530 17830 15550
rect 17810 15370 17830 15390
rect 17810 15210 17830 15230
rect 17890 16170 17910 16190
rect 17890 16010 17910 16030
rect 17890 15850 17910 15870
rect 17890 15690 17910 15710
rect 17890 15530 17910 15550
rect 17890 15370 17910 15390
rect 17890 15210 17910 15230
rect 17970 16170 17990 16190
rect 17970 16010 17990 16030
rect 17970 15850 17990 15870
rect 17970 15690 17990 15710
rect 17970 15530 17990 15550
rect 17970 15370 17990 15390
rect 17970 15210 17990 15230
rect 18050 16170 18070 16190
rect 18050 16010 18070 16030
rect 18050 15850 18070 15870
rect 18050 15690 18070 15710
rect 18050 15530 18070 15550
rect 18050 15370 18070 15390
rect 18050 15210 18070 15230
rect 18130 16170 18150 16190
rect 18130 16010 18150 16030
rect 18130 15850 18150 15870
rect 18130 15690 18150 15710
rect 18130 15530 18150 15550
rect 18130 15370 18150 15390
rect 18130 15210 18150 15230
rect 18210 16170 18230 16190
rect 18210 16010 18230 16030
rect 18210 15850 18230 15870
rect 18210 15690 18230 15710
rect 18210 15530 18230 15550
rect 18210 15370 18230 15390
rect 18210 15210 18230 15230
rect 18290 16170 18310 16190
rect 18290 16010 18310 16030
rect 18290 15850 18310 15870
rect 18290 15690 18310 15710
rect 18290 15530 18310 15550
rect 18290 15370 18310 15390
rect 18290 15210 18310 15230
rect 18370 16170 18390 16190
rect 18370 16010 18390 16030
rect 18370 15850 18390 15870
rect 18370 15690 18390 15710
rect 18370 15530 18390 15550
rect 18370 15370 18390 15390
rect 18370 15210 18390 15230
rect 18450 16170 18470 16190
rect 18450 16010 18470 16030
rect 18450 15850 18470 15870
rect 18450 15690 18470 15710
rect 18450 15530 18470 15550
rect 18450 15370 18470 15390
rect 18450 15210 18470 15230
rect 18530 16170 18550 16190
rect 18530 16010 18550 16030
rect 18530 15850 18550 15870
rect 18530 15690 18550 15710
rect 18530 15530 18550 15550
rect 18530 15370 18550 15390
rect 18530 15210 18550 15230
rect 18610 16170 18630 16190
rect 18610 16010 18630 16030
rect 18610 15850 18630 15870
rect 18610 15690 18630 15710
rect 18610 15530 18630 15550
rect 18610 15370 18630 15390
rect 18610 15210 18630 15230
rect 18690 16170 18710 16190
rect 18690 16010 18710 16030
rect 18690 15850 18710 15870
rect 18690 15690 18710 15710
rect 18690 15530 18710 15550
rect 18690 15370 18710 15390
rect 18690 15210 18710 15230
rect 18770 16170 18790 16190
rect 18770 16010 18790 16030
rect 18770 15850 18790 15870
rect 18770 15690 18790 15710
rect 18770 15530 18790 15550
rect 18770 15370 18790 15390
rect 18770 15210 18790 15230
rect 18850 16170 18870 16190
rect 18850 16010 18870 16030
rect 18850 15850 18870 15870
rect 18850 15690 18870 15710
rect 18850 15530 18870 15550
rect 18850 15370 18870 15390
rect 18850 15210 18870 15230
rect 18930 16170 18950 16190
rect 18930 16010 18950 16030
rect 18930 15850 18950 15870
rect 18930 15690 18950 15710
rect 18930 15530 18950 15550
rect 18930 15370 18950 15390
rect 18930 15210 18950 15230
rect 19010 16170 19030 16190
rect 19010 16010 19030 16030
rect 19010 15850 19030 15870
rect 19010 15690 19030 15710
rect 19010 15530 19030 15550
rect 19010 15370 19030 15390
rect 19010 15210 19030 15230
rect 19090 16170 19110 16190
rect 19090 16010 19110 16030
rect 19090 15850 19110 15870
rect 19090 15690 19110 15710
rect 19090 15530 19110 15550
rect 19090 15370 19110 15390
rect 19090 15210 19110 15230
rect 19170 16170 19190 16190
rect 19170 16010 19190 16030
rect 19170 15850 19190 15870
rect 19170 15690 19190 15710
rect 19170 15530 19190 15550
rect 19170 15370 19190 15390
rect 19170 15210 19190 15230
rect 19250 16170 19270 16190
rect 19250 16010 19270 16030
rect 19250 15850 19270 15870
rect 19250 15690 19270 15710
rect 19250 15530 19270 15550
rect 19250 15370 19270 15390
rect 19250 15210 19270 15230
rect 19330 16170 19350 16190
rect 19330 16010 19350 16030
rect 19330 15850 19350 15870
rect 19330 15690 19350 15710
rect 19330 15530 19350 15550
rect 19330 15370 19350 15390
rect 19330 15210 19350 15230
rect 19410 16170 19430 16190
rect 19410 16010 19430 16030
rect 19410 15850 19430 15870
rect 19410 15690 19430 15710
rect 19410 15530 19430 15550
rect 19410 15370 19430 15390
rect 19410 15210 19430 15230
rect 19490 16170 19510 16190
rect 19490 16010 19510 16030
rect 19490 15850 19510 15870
rect 19490 15690 19510 15710
rect 19490 15530 19510 15550
rect 19490 15370 19510 15390
rect 19490 15210 19510 15230
rect 19570 16170 19590 16190
rect 19570 16010 19590 16030
rect 19570 15850 19590 15870
rect 19570 15690 19590 15710
rect 19570 15530 19590 15550
rect 19570 15370 19590 15390
rect 19570 15210 19590 15230
rect 19650 16170 19670 16190
rect 19650 16010 19670 16030
rect 19650 15850 19670 15870
rect 19650 15690 19670 15710
rect 19650 15530 19670 15550
rect 19650 15370 19670 15390
rect 19650 15210 19670 15230
rect 19730 16170 19750 16190
rect 19730 16010 19750 16030
rect 19730 15850 19750 15870
rect 19730 15690 19750 15710
rect 19730 15530 19750 15550
rect 19730 15370 19750 15390
rect 19730 15210 19750 15230
rect 19810 16170 19830 16190
rect 19810 16010 19830 16030
rect 19810 15850 19830 15870
rect 19810 15690 19830 15710
rect 19810 15530 19830 15550
rect 19810 15370 19830 15390
rect 19810 15210 19830 15230
rect 19890 16170 19910 16190
rect 19890 16010 19910 16030
rect 19890 15850 19910 15870
rect 19890 15690 19910 15710
rect 19890 15530 19910 15550
rect 19890 15370 19910 15390
rect 19890 15210 19910 15230
rect 19970 16170 19990 16190
rect 19970 16010 19990 16030
rect 19970 15850 19990 15870
rect 19970 15690 19990 15710
rect 19970 15530 19990 15550
rect 19970 15370 19990 15390
rect 19970 15210 19990 15230
rect 20050 16170 20070 16190
rect 20050 16010 20070 16030
rect 20050 15850 20070 15870
rect 20050 15690 20070 15710
rect 20050 15530 20070 15550
rect 20050 15370 20070 15390
rect 20050 15210 20070 15230
rect 20130 16170 20150 16190
rect 20130 16010 20150 16030
rect 20130 15850 20150 15870
rect 20130 15690 20150 15710
rect 20130 15530 20150 15550
rect 20130 15370 20150 15390
rect 20130 15210 20150 15230
rect 20210 16170 20230 16190
rect 20210 16010 20230 16030
rect 20210 15850 20230 15870
rect 20210 15690 20230 15710
rect 20210 15530 20230 15550
rect 20210 15370 20230 15390
rect 20210 15210 20230 15230
rect 20290 16170 20310 16190
rect 20290 16010 20310 16030
rect 20290 15850 20310 15870
rect 20290 15690 20310 15710
rect 20290 15530 20310 15550
rect 20290 15370 20310 15390
rect 20290 15210 20310 15230
rect 20370 16170 20390 16190
rect 20370 16010 20390 16030
rect 20370 15850 20390 15870
rect 20370 15690 20390 15710
rect 20370 15530 20390 15550
rect 20370 15370 20390 15390
rect 20370 15210 20390 15230
rect 20450 16170 20470 16190
rect 20450 16010 20470 16030
rect 20450 15850 20470 15870
rect 20450 15690 20470 15710
rect 20450 15530 20470 15550
rect 20450 15370 20470 15390
rect 20450 15210 20470 15230
rect 20530 16170 20550 16190
rect 20530 16010 20550 16030
rect 20530 15850 20550 15870
rect 20530 15690 20550 15710
rect 20530 15530 20550 15550
rect 20530 15370 20550 15390
rect 20530 15210 20550 15230
rect 20610 16170 20630 16190
rect 20610 16010 20630 16030
rect 20610 15850 20630 15870
rect 20610 15690 20630 15710
rect 20610 15530 20630 15550
rect 20610 15370 20630 15390
rect 20610 15210 20630 15230
rect 20690 16170 20710 16190
rect 20690 16010 20710 16030
rect 20690 15850 20710 15870
rect 20690 15690 20710 15710
rect 20690 15530 20710 15550
rect 20690 15370 20710 15390
rect 20690 15210 20710 15230
rect 20770 16170 20790 16190
rect 20770 16010 20790 16030
rect 20770 15850 20790 15870
rect 20770 15690 20790 15710
rect 20770 15530 20790 15550
rect 20770 15370 20790 15390
rect 20770 15210 20790 15230
rect 20850 16170 20870 16190
rect 20850 16010 20870 16030
rect 20850 15850 20870 15870
rect 20850 15690 20870 15710
rect 20850 15530 20870 15550
rect 20850 15370 20870 15390
rect 20850 15210 20870 15230
rect 20930 16170 20950 16190
rect 20930 16010 20950 16030
rect 20930 15850 20950 15870
rect 20930 15690 20950 15710
rect 20930 15530 20950 15550
rect 20930 15370 20950 15390
rect 20930 15210 20950 15230
rect 10 15130 30 15150
rect 10 14970 30 14990
rect 90 15130 110 15150
rect 90 14970 110 14990
rect 170 15130 190 15150
rect 170 14970 190 14990
rect 250 15130 270 15150
rect 250 14970 270 14990
rect 330 15130 350 15150
rect 330 14970 350 14990
rect 410 15130 430 15150
rect 410 14970 430 14990
rect 490 15130 510 15150
rect 490 14970 510 14990
rect 570 15130 590 15150
rect 570 14970 590 14990
rect 650 15130 670 15150
rect 650 14970 670 14990
rect 730 15130 750 15150
rect 730 14970 750 14990
rect 810 15130 830 15150
rect 810 14970 830 14990
rect 890 15130 910 15150
rect 890 14970 910 14990
rect 970 15130 990 15150
rect 970 14970 990 14990
rect 1050 15130 1070 15150
rect 1050 14970 1070 14990
rect 1130 15130 1150 15150
rect 1130 14970 1150 14990
rect 1210 15130 1230 15150
rect 1210 14970 1230 14990
rect 1290 15130 1310 15150
rect 1290 14970 1310 14990
rect 1370 15130 1390 15150
rect 1370 14970 1390 14990
rect 1450 15130 1470 15150
rect 1450 14970 1470 14990
rect 1530 15130 1550 15150
rect 1530 14970 1550 14990
rect 1610 15130 1630 15150
rect 1610 14970 1630 14990
rect 1690 15130 1710 15150
rect 1690 14970 1710 14990
rect 1770 15130 1790 15150
rect 1770 14970 1790 14990
rect 1850 15130 1870 15150
rect 1850 14970 1870 14990
rect 1930 15130 1950 15150
rect 1930 14970 1950 14990
rect 2010 15130 2030 15150
rect 2010 14970 2030 14990
rect 2090 15130 2110 15150
rect 2090 14970 2110 14990
rect 2170 15130 2190 15150
rect 2170 14970 2190 14990
rect 2250 15130 2270 15150
rect 2250 14970 2270 14990
rect 2330 15130 2350 15150
rect 2330 14970 2350 14990
rect 2410 15130 2430 15150
rect 2410 14970 2430 14990
rect 2490 15130 2510 15150
rect 2490 14970 2510 14990
rect 2570 15130 2590 15150
rect 2570 14970 2590 14990
rect 2650 15130 2670 15150
rect 2650 14970 2670 14990
rect 2730 15130 2750 15150
rect 2730 14970 2750 14990
rect 2810 15130 2830 15150
rect 2810 14970 2830 14990
rect 2890 15130 2910 15150
rect 2890 14970 2910 14990
rect 2970 15130 2990 15150
rect 2970 14970 2990 14990
rect 3050 15130 3070 15150
rect 3050 14970 3070 14990
rect 3130 15130 3150 15150
rect 3130 14970 3150 14990
rect 3210 15130 3230 15150
rect 3210 14970 3230 14990
rect 3290 15130 3310 15150
rect 3290 14970 3310 14990
rect 3370 15130 3390 15150
rect 3370 14970 3390 14990
rect 3450 15130 3470 15150
rect 3450 14970 3470 14990
rect 3530 15130 3550 15150
rect 3530 14970 3550 14990
rect 3610 15130 3630 15150
rect 3610 14970 3630 14990
rect 3690 15130 3710 15150
rect 3690 14970 3710 14990
rect 3770 15130 3790 15150
rect 3770 14970 3790 14990
rect 3850 15130 3870 15150
rect 3850 14970 3870 14990
rect 3930 15130 3950 15150
rect 3930 14970 3950 14990
rect 4010 15130 4030 15150
rect 4010 14970 4030 14990
rect 4090 15130 4110 15150
rect 4090 14970 4110 14990
rect 4170 15130 4190 15150
rect 4170 14970 4190 14990
rect 6250 15130 6270 15150
rect 6250 14970 6270 14990
rect 6330 15130 6350 15150
rect 6330 14970 6350 14990
rect 6410 15130 6430 15150
rect 6410 14970 6430 14990
rect 6490 15130 6510 15150
rect 6490 14970 6510 14990
rect 6570 15130 6590 15150
rect 6570 14970 6590 14990
rect 6650 15130 6670 15150
rect 6650 14970 6670 14990
rect 6730 15130 6750 15150
rect 6730 14970 6750 14990
rect 6810 15130 6830 15150
rect 6810 14970 6830 14990
rect 6890 15130 6910 15150
rect 6890 14970 6910 14990
rect 6970 15130 6990 15150
rect 6970 14970 6990 14990
rect 7050 15130 7070 15150
rect 7050 14970 7070 14990
rect 7130 15130 7150 15150
rect 7130 14970 7150 14990
rect 7210 15130 7230 15150
rect 7210 14970 7230 14990
rect 7290 15130 7310 15150
rect 7290 14970 7310 14990
rect 7370 15130 7390 15150
rect 7370 14970 7390 14990
rect 7450 15130 7470 15150
rect 7450 14970 7470 14990
rect 7530 15130 7550 15150
rect 7530 14970 7550 14990
rect 7610 15130 7630 15150
rect 7610 14970 7630 14990
rect 7690 15130 7710 15150
rect 7690 14970 7710 14990
rect 7770 15130 7790 15150
rect 7770 14970 7790 14990
rect 7850 15130 7870 15150
rect 7850 14970 7870 14990
rect 7930 15130 7950 15150
rect 7930 14970 7950 14990
rect 8010 15130 8030 15150
rect 8010 14970 8030 14990
rect 8090 15130 8110 15150
rect 8090 14970 8110 14990
rect 8170 15130 8190 15150
rect 8170 14970 8190 14990
rect 8250 15130 8270 15150
rect 8250 14970 8270 14990
rect 8330 15130 8350 15150
rect 8330 14970 8350 14990
rect 8410 15130 8430 15150
rect 8410 14970 8430 14990
rect 8490 15130 8510 15150
rect 8490 14970 8510 14990
rect 8570 15130 8590 15150
rect 8570 14970 8590 14990
rect 8650 15130 8670 15150
rect 8650 14970 8670 14990
rect 8730 15130 8750 15150
rect 8730 14970 8750 14990
rect 8810 15130 8830 15150
rect 8810 14970 8830 14990
rect 8890 15130 8910 15150
rect 8890 14970 8910 14990
rect 8970 15130 8990 15150
rect 8970 14970 8990 14990
rect 9050 15130 9070 15150
rect 9050 14970 9070 14990
rect 9130 15130 9150 15150
rect 9130 14970 9150 14990
rect 9210 15130 9230 15150
rect 9210 14970 9230 14990
rect 9290 15130 9310 15150
rect 9290 14970 9310 14990
rect 9370 15130 9390 15150
rect 9370 14970 9390 14990
rect 9450 15130 9470 15150
rect 9450 14970 9470 14990
rect 11570 15130 11590 15150
rect 11570 14970 11590 14990
rect 11650 15130 11670 15150
rect 11650 14970 11670 14990
rect 11730 15130 11750 15150
rect 11730 14970 11750 14990
rect 11810 15130 11830 15150
rect 11810 14970 11830 14990
rect 11890 15130 11910 15150
rect 11890 14970 11910 14990
rect 11970 15130 11990 15150
rect 11970 14970 11990 14990
rect 12050 15130 12070 15150
rect 12050 14970 12070 14990
rect 12130 15130 12150 15150
rect 12130 14970 12150 14990
rect 12210 15130 12230 15150
rect 12210 14970 12230 14990
rect 12290 15130 12310 15150
rect 12290 14970 12310 14990
rect 12370 15130 12390 15150
rect 12370 14970 12390 14990
rect 12450 15130 12470 15150
rect 12450 14970 12470 14990
rect 12530 15130 12550 15150
rect 12530 14970 12550 14990
rect 12610 15130 12630 15150
rect 12610 14970 12630 14990
rect 12690 15130 12710 15150
rect 12690 14970 12710 14990
rect 12770 15130 12790 15150
rect 12770 14970 12790 14990
rect 12850 15130 12870 15150
rect 12850 14970 12870 14990
rect 12930 15130 12950 15150
rect 12930 14970 12950 14990
rect 13010 15130 13030 15150
rect 13010 14970 13030 14990
rect 13090 15130 13110 15150
rect 13090 14970 13110 14990
rect 13170 15130 13190 15150
rect 13170 14970 13190 14990
rect 13250 15130 13270 15150
rect 13250 14970 13270 14990
rect 13330 15130 13350 15150
rect 13330 14970 13350 14990
rect 13410 15130 13430 15150
rect 13410 14970 13430 14990
rect 13490 15130 13510 15150
rect 13490 14970 13510 14990
rect 13570 15130 13590 15150
rect 13570 14970 13590 14990
rect 13650 15130 13670 15150
rect 13650 14970 13670 14990
rect 13730 15130 13750 15150
rect 13730 14970 13750 14990
rect 13810 15130 13830 15150
rect 13810 14970 13830 14990
rect 13890 15130 13910 15150
rect 13890 14970 13910 14990
rect 13970 15130 13990 15150
rect 13970 14970 13990 14990
rect 14050 15130 14070 15150
rect 14050 14970 14070 14990
rect 14130 15130 14150 15150
rect 14130 14970 14150 14990
rect 14210 15130 14230 15150
rect 14210 14970 14230 14990
rect 14290 15130 14310 15150
rect 14290 14970 14310 14990
rect 14370 15130 14390 15150
rect 14370 14970 14390 14990
rect 14450 15130 14470 15150
rect 14450 14970 14470 14990
rect 14530 15130 14550 15150
rect 14530 14970 14550 14990
rect 14610 15130 14630 15150
rect 14610 14970 14630 14990
rect 14690 15130 14710 15150
rect 14690 14970 14710 14990
rect 16770 15130 16790 15150
rect 16770 14970 16790 14990
rect 16850 15130 16870 15150
rect 16850 14970 16870 14990
rect 16930 15130 16950 15150
rect 16930 14970 16950 14990
rect 17010 15130 17030 15150
rect 17010 14970 17030 14990
rect 17090 15130 17110 15150
rect 17090 14970 17110 14990
rect 17170 15130 17190 15150
rect 17170 14970 17190 14990
rect 17250 15130 17270 15150
rect 17250 14970 17270 14990
rect 17330 15130 17350 15150
rect 17330 14970 17350 14990
rect 17410 15130 17430 15150
rect 17410 14970 17430 14990
rect 17490 15130 17510 15150
rect 17490 14970 17510 14990
rect 17570 15130 17590 15150
rect 17570 14970 17590 14990
rect 17650 15130 17670 15150
rect 17650 14970 17670 14990
rect 17730 15130 17750 15150
rect 17730 14970 17750 14990
rect 17810 15130 17830 15150
rect 17810 14970 17830 14990
rect 17890 15130 17910 15150
rect 17890 14970 17910 14990
rect 17970 15130 17990 15150
rect 17970 14970 17990 14990
rect 18050 15130 18070 15150
rect 18050 14970 18070 14990
rect 18130 15130 18150 15150
rect 18130 14970 18150 14990
rect 18210 15130 18230 15150
rect 18210 14970 18230 14990
rect 18290 15130 18310 15150
rect 18290 14970 18310 14990
rect 18370 15130 18390 15150
rect 18370 14970 18390 14990
rect 18450 15130 18470 15150
rect 18450 14970 18470 14990
rect 18530 15130 18550 15150
rect 18530 14970 18550 14990
rect 18610 15130 18630 15150
rect 18610 14970 18630 14990
rect 18690 15130 18710 15150
rect 18690 14970 18710 14990
rect 18770 15130 18790 15150
rect 18770 14970 18790 14990
rect 18850 15130 18870 15150
rect 18850 14970 18870 14990
rect 18930 15130 18950 15150
rect 18930 14970 18950 14990
rect 19010 15130 19030 15150
rect 19010 14970 19030 14990
rect 19090 15130 19110 15150
rect 19090 14970 19110 14990
rect 19170 15130 19190 15150
rect 19170 14970 19190 14990
rect 19250 15130 19270 15150
rect 19250 14970 19270 14990
rect 19330 15130 19350 15150
rect 19330 14970 19350 14990
rect 19410 15130 19430 15150
rect 19410 14970 19430 14990
rect 19490 15130 19510 15150
rect 19490 14970 19510 14990
rect 19570 15130 19590 15150
rect 19570 14970 19590 14990
rect 19650 15130 19670 15150
rect 19650 14970 19670 14990
rect 19730 15130 19750 15150
rect 19730 14970 19750 14990
rect 19810 15130 19830 15150
rect 19810 14970 19830 14990
rect 19890 15130 19910 15150
rect 19890 14970 19910 14990
rect 19970 15130 19990 15150
rect 19970 14970 19990 14990
rect 20050 15130 20070 15150
rect 20050 14970 20070 14990
rect 20130 15130 20150 15150
rect 20130 14970 20150 14990
rect 20210 15130 20230 15150
rect 20210 14970 20230 14990
rect 20290 15130 20310 15150
rect 20290 14970 20310 14990
rect 20370 15130 20390 15150
rect 20370 14970 20390 14990
rect 20450 15130 20470 15150
rect 20450 14970 20470 14990
rect 20530 15130 20550 15150
rect 20530 14970 20550 14990
rect 20610 15130 20630 15150
rect 20610 14970 20630 14990
rect 20690 15130 20710 15150
rect 20690 14970 20710 14990
rect 20770 15130 20790 15150
rect 20770 14970 20790 14990
rect 20850 15130 20870 15150
rect 20850 14970 20870 14990
rect 20930 15130 20950 15150
rect 20930 14970 20950 14990
rect 10 14890 30 14910
rect 10 14730 30 14750
rect 90 14890 110 14910
rect 90 14730 110 14750
rect 170 14890 190 14910
rect 170 14730 190 14750
rect 250 14890 270 14910
rect 250 14730 270 14750
rect 330 14890 350 14910
rect 330 14730 350 14750
rect 410 14890 430 14910
rect 410 14730 430 14750
rect 490 14890 510 14910
rect 490 14730 510 14750
rect 570 14890 590 14910
rect 570 14730 590 14750
rect 650 14890 670 14910
rect 650 14730 670 14750
rect 730 14890 750 14910
rect 730 14730 750 14750
rect 810 14890 830 14910
rect 810 14730 830 14750
rect 890 14890 910 14910
rect 890 14730 910 14750
rect 970 14890 990 14910
rect 970 14730 990 14750
rect 1050 14890 1070 14910
rect 1050 14730 1070 14750
rect 1130 14890 1150 14910
rect 1130 14730 1150 14750
rect 1210 14890 1230 14910
rect 1210 14730 1230 14750
rect 1290 14890 1310 14910
rect 1290 14730 1310 14750
rect 1370 14890 1390 14910
rect 1370 14730 1390 14750
rect 1450 14890 1470 14910
rect 1450 14730 1470 14750
rect 1530 14890 1550 14910
rect 1530 14730 1550 14750
rect 1610 14890 1630 14910
rect 1610 14730 1630 14750
rect 1690 14890 1710 14910
rect 1690 14730 1710 14750
rect 1770 14890 1790 14910
rect 1770 14730 1790 14750
rect 1850 14890 1870 14910
rect 1850 14730 1870 14750
rect 1930 14890 1950 14910
rect 1930 14730 1950 14750
rect 2010 14890 2030 14910
rect 2010 14730 2030 14750
rect 2090 14890 2110 14910
rect 2090 14730 2110 14750
rect 2170 14890 2190 14910
rect 2170 14730 2190 14750
rect 2250 14890 2270 14910
rect 2250 14730 2270 14750
rect 2330 14890 2350 14910
rect 2330 14730 2350 14750
rect 2410 14890 2430 14910
rect 2410 14730 2430 14750
rect 2490 14890 2510 14910
rect 2490 14730 2510 14750
rect 2570 14890 2590 14910
rect 2570 14730 2590 14750
rect 2650 14890 2670 14910
rect 2650 14730 2670 14750
rect 2730 14890 2750 14910
rect 2730 14730 2750 14750
rect 2810 14890 2830 14910
rect 2810 14730 2830 14750
rect 2890 14890 2910 14910
rect 2890 14730 2910 14750
rect 2970 14890 2990 14910
rect 2970 14730 2990 14750
rect 3050 14890 3070 14910
rect 3050 14730 3070 14750
rect 3130 14890 3150 14910
rect 3130 14730 3150 14750
rect 3210 14890 3230 14910
rect 3210 14730 3230 14750
rect 3290 14890 3310 14910
rect 3290 14730 3310 14750
rect 3370 14890 3390 14910
rect 3370 14730 3390 14750
rect 3450 14890 3470 14910
rect 3450 14730 3470 14750
rect 3530 14890 3550 14910
rect 3530 14730 3550 14750
rect 3610 14890 3630 14910
rect 3610 14730 3630 14750
rect 3690 14890 3710 14910
rect 3690 14730 3710 14750
rect 3770 14890 3790 14910
rect 3770 14730 3790 14750
rect 3850 14890 3870 14910
rect 3850 14730 3870 14750
rect 3930 14890 3950 14910
rect 3930 14730 3950 14750
rect 4010 14890 4030 14910
rect 4010 14730 4030 14750
rect 4090 14890 4110 14910
rect 4090 14730 4110 14750
rect 4170 14890 4190 14910
rect 4170 14730 4190 14750
rect 6250 14890 6270 14910
rect 6250 14730 6270 14750
rect 6330 14890 6350 14910
rect 6330 14730 6350 14750
rect 6410 14890 6430 14910
rect 6410 14730 6430 14750
rect 6490 14890 6510 14910
rect 6490 14730 6510 14750
rect 6570 14890 6590 14910
rect 6570 14730 6590 14750
rect 6650 14890 6670 14910
rect 6650 14730 6670 14750
rect 6730 14890 6750 14910
rect 6730 14730 6750 14750
rect 6810 14890 6830 14910
rect 6810 14730 6830 14750
rect 6890 14890 6910 14910
rect 6890 14730 6910 14750
rect 6970 14890 6990 14910
rect 6970 14730 6990 14750
rect 7050 14890 7070 14910
rect 7050 14730 7070 14750
rect 7130 14890 7150 14910
rect 7130 14730 7150 14750
rect 7210 14890 7230 14910
rect 7210 14730 7230 14750
rect 7290 14890 7310 14910
rect 7290 14730 7310 14750
rect 7370 14890 7390 14910
rect 7370 14730 7390 14750
rect 7450 14890 7470 14910
rect 7450 14730 7470 14750
rect 7530 14890 7550 14910
rect 7530 14730 7550 14750
rect 7610 14890 7630 14910
rect 7610 14730 7630 14750
rect 7690 14890 7710 14910
rect 7690 14730 7710 14750
rect 7770 14890 7790 14910
rect 7770 14730 7790 14750
rect 7850 14890 7870 14910
rect 7850 14730 7870 14750
rect 7930 14890 7950 14910
rect 7930 14730 7950 14750
rect 8010 14890 8030 14910
rect 8010 14730 8030 14750
rect 8090 14890 8110 14910
rect 8090 14730 8110 14750
rect 8170 14890 8190 14910
rect 8170 14730 8190 14750
rect 8250 14890 8270 14910
rect 8250 14730 8270 14750
rect 8330 14890 8350 14910
rect 8330 14730 8350 14750
rect 8410 14890 8430 14910
rect 8410 14730 8430 14750
rect 8490 14890 8510 14910
rect 8490 14730 8510 14750
rect 8570 14890 8590 14910
rect 8570 14730 8590 14750
rect 8650 14890 8670 14910
rect 8650 14730 8670 14750
rect 8730 14890 8750 14910
rect 8730 14730 8750 14750
rect 8810 14890 8830 14910
rect 8810 14730 8830 14750
rect 8890 14890 8910 14910
rect 8890 14730 8910 14750
rect 8970 14890 8990 14910
rect 8970 14730 8990 14750
rect 9050 14890 9070 14910
rect 9050 14730 9070 14750
rect 9130 14890 9150 14910
rect 9130 14730 9150 14750
rect 9210 14890 9230 14910
rect 9210 14730 9230 14750
rect 9290 14890 9310 14910
rect 9290 14730 9310 14750
rect 9370 14890 9390 14910
rect 9370 14730 9390 14750
rect 9450 14890 9470 14910
rect 9450 14730 9470 14750
rect 11570 14890 11590 14910
rect 11570 14730 11590 14750
rect 11650 14890 11670 14910
rect 11650 14730 11670 14750
rect 11730 14890 11750 14910
rect 11730 14730 11750 14750
rect 11810 14890 11830 14910
rect 11810 14730 11830 14750
rect 11890 14890 11910 14910
rect 11890 14730 11910 14750
rect 11970 14890 11990 14910
rect 11970 14730 11990 14750
rect 12050 14890 12070 14910
rect 12050 14730 12070 14750
rect 12130 14890 12150 14910
rect 12130 14730 12150 14750
rect 12210 14890 12230 14910
rect 12210 14730 12230 14750
rect 12290 14890 12310 14910
rect 12290 14730 12310 14750
rect 12370 14890 12390 14910
rect 12370 14730 12390 14750
rect 12450 14890 12470 14910
rect 12450 14730 12470 14750
rect 12530 14890 12550 14910
rect 12530 14730 12550 14750
rect 12610 14890 12630 14910
rect 12610 14730 12630 14750
rect 12690 14890 12710 14910
rect 12690 14730 12710 14750
rect 12770 14890 12790 14910
rect 12770 14730 12790 14750
rect 12850 14890 12870 14910
rect 12850 14730 12870 14750
rect 12930 14890 12950 14910
rect 12930 14730 12950 14750
rect 13010 14890 13030 14910
rect 13010 14730 13030 14750
rect 13090 14890 13110 14910
rect 13090 14730 13110 14750
rect 13170 14890 13190 14910
rect 13170 14730 13190 14750
rect 13250 14890 13270 14910
rect 13250 14730 13270 14750
rect 13330 14890 13350 14910
rect 13330 14730 13350 14750
rect 13410 14890 13430 14910
rect 13410 14730 13430 14750
rect 13490 14890 13510 14910
rect 13490 14730 13510 14750
rect 13570 14890 13590 14910
rect 13570 14730 13590 14750
rect 13650 14890 13670 14910
rect 13650 14730 13670 14750
rect 13730 14890 13750 14910
rect 13730 14730 13750 14750
rect 13810 14890 13830 14910
rect 13810 14730 13830 14750
rect 13890 14890 13910 14910
rect 13890 14730 13910 14750
rect 13970 14890 13990 14910
rect 13970 14730 13990 14750
rect 14050 14890 14070 14910
rect 14050 14730 14070 14750
rect 14130 14890 14150 14910
rect 14130 14730 14150 14750
rect 14210 14890 14230 14910
rect 14210 14730 14230 14750
rect 14290 14890 14310 14910
rect 14290 14730 14310 14750
rect 14370 14890 14390 14910
rect 14370 14730 14390 14750
rect 14450 14890 14470 14910
rect 14450 14730 14470 14750
rect 14530 14890 14550 14910
rect 14530 14730 14550 14750
rect 14610 14890 14630 14910
rect 14610 14730 14630 14750
rect 14690 14890 14710 14910
rect 14690 14730 14710 14750
rect 16770 14890 16790 14910
rect 16770 14730 16790 14750
rect 16850 14890 16870 14910
rect 16850 14730 16870 14750
rect 16930 14890 16950 14910
rect 16930 14730 16950 14750
rect 17010 14890 17030 14910
rect 17010 14730 17030 14750
rect 17090 14890 17110 14910
rect 17090 14730 17110 14750
rect 17170 14890 17190 14910
rect 17170 14730 17190 14750
rect 17250 14890 17270 14910
rect 17250 14730 17270 14750
rect 17330 14890 17350 14910
rect 17330 14730 17350 14750
rect 17410 14890 17430 14910
rect 17410 14730 17430 14750
rect 17490 14890 17510 14910
rect 17490 14730 17510 14750
rect 17570 14890 17590 14910
rect 17570 14730 17590 14750
rect 17650 14890 17670 14910
rect 17650 14730 17670 14750
rect 17730 14890 17750 14910
rect 17730 14730 17750 14750
rect 17810 14890 17830 14910
rect 17810 14730 17830 14750
rect 17890 14890 17910 14910
rect 17890 14730 17910 14750
rect 17970 14890 17990 14910
rect 17970 14730 17990 14750
rect 18050 14890 18070 14910
rect 18050 14730 18070 14750
rect 18130 14890 18150 14910
rect 18130 14730 18150 14750
rect 18210 14890 18230 14910
rect 18210 14730 18230 14750
rect 18290 14890 18310 14910
rect 18290 14730 18310 14750
rect 18370 14890 18390 14910
rect 18370 14730 18390 14750
rect 18450 14890 18470 14910
rect 18450 14730 18470 14750
rect 18530 14890 18550 14910
rect 18530 14730 18550 14750
rect 18610 14890 18630 14910
rect 18610 14730 18630 14750
rect 18690 14890 18710 14910
rect 18690 14730 18710 14750
rect 18770 14890 18790 14910
rect 18770 14730 18790 14750
rect 18850 14890 18870 14910
rect 18850 14730 18870 14750
rect 18930 14890 18950 14910
rect 18930 14730 18950 14750
rect 19010 14890 19030 14910
rect 19010 14730 19030 14750
rect 19090 14890 19110 14910
rect 19090 14730 19110 14750
rect 19170 14890 19190 14910
rect 19170 14730 19190 14750
rect 19250 14890 19270 14910
rect 19250 14730 19270 14750
rect 19330 14890 19350 14910
rect 19330 14730 19350 14750
rect 19410 14890 19430 14910
rect 19410 14730 19430 14750
rect 19490 14890 19510 14910
rect 19490 14730 19510 14750
rect 19570 14890 19590 14910
rect 19570 14730 19590 14750
rect 19650 14890 19670 14910
rect 19650 14730 19670 14750
rect 19730 14890 19750 14910
rect 19730 14730 19750 14750
rect 19810 14890 19830 14910
rect 19810 14730 19830 14750
rect 19890 14890 19910 14910
rect 19890 14730 19910 14750
rect 19970 14890 19990 14910
rect 19970 14730 19990 14750
rect 20050 14890 20070 14910
rect 20050 14730 20070 14750
rect 20130 14890 20150 14910
rect 20130 14730 20150 14750
rect 20210 14890 20230 14910
rect 20210 14730 20230 14750
rect 20290 14890 20310 14910
rect 20290 14730 20310 14750
rect 20370 14890 20390 14910
rect 20370 14730 20390 14750
rect 20450 14890 20470 14910
rect 20450 14730 20470 14750
rect 20530 14890 20550 14910
rect 20530 14730 20550 14750
rect 20610 14890 20630 14910
rect 20610 14730 20630 14750
rect 20690 14890 20710 14910
rect 20690 14730 20710 14750
rect 20770 14890 20790 14910
rect 20770 14730 20790 14750
rect 20850 14890 20870 14910
rect 20850 14730 20870 14750
rect 20930 14890 20950 14910
rect 20930 14730 20950 14750
<< metal1 >>
rect 0 18675 40 18680
rect 0 18645 5 18675
rect 35 18645 40 18675
rect 0 18640 40 18645
rect 80 18675 120 18680
rect 80 18645 85 18675
rect 115 18645 120 18675
rect 80 18640 120 18645
rect 160 18675 200 18680
rect 160 18645 165 18675
rect 195 18645 200 18675
rect 160 18640 200 18645
rect 240 18675 280 18680
rect 240 18645 245 18675
rect 275 18645 280 18675
rect 240 18640 280 18645
rect 320 18675 360 18680
rect 320 18645 325 18675
rect 355 18645 360 18675
rect 320 18640 360 18645
rect 400 18675 440 18680
rect 400 18645 405 18675
rect 435 18645 440 18675
rect 400 18640 440 18645
rect 480 18675 520 18680
rect 480 18645 485 18675
rect 515 18645 520 18675
rect 480 18640 520 18645
rect 560 18675 600 18680
rect 560 18645 565 18675
rect 595 18645 600 18675
rect 560 18640 600 18645
rect 640 18675 680 18680
rect 640 18645 645 18675
rect 675 18645 680 18675
rect 640 18640 680 18645
rect 720 18675 760 18680
rect 720 18645 725 18675
rect 755 18645 760 18675
rect 720 18640 760 18645
rect 800 18675 840 18680
rect 800 18645 805 18675
rect 835 18645 840 18675
rect 800 18640 840 18645
rect 880 18675 920 18680
rect 880 18645 885 18675
rect 915 18645 920 18675
rect 880 18640 920 18645
rect 960 18675 1000 18680
rect 960 18645 965 18675
rect 995 18645 1000 18675
rect 960 18640 1000 18645
rect 1040 18675 1080 18680
rect 1040 18645 1045 18675
rect 1075 18645 1080 18675
rect 1040 18640 1080 18645
rect 1120 18675 1160 18680
rect 1120 18645 1125 18675
rect 1155 18645 1160 18675
rect 1120 18640 1160 18645
rect 1200 18675 1240 18680
rect 1200 18645 1205 18675
rect 1235 18645 1240 18675
rect 1200 18640 1240 18645
rect 1280 18675 1320 18680
rect 1280 18645 1285 18675
rect 1315 18645 1320 18675
rect 1280 18640 1320 18645
rect 1360 18675 1400 18680
rect 1360 18645 1365 18675
rect 1395 18645 1400 18675
rect 1360 18640 1400 18645
rect 1440 18675 1480 18680
rect 1440 18645 1445 18675
rect 1475 18645 1480 18675
rect 1440 18640 1480 18645
rect 1520 18675 1560 18680
rect 1520 18645 1525 18675
rect 1555 18645 1560 18675
rect 1520 18640 1560 18645
rect 1600 18675 1640 18680
rect 1600 18645 1605 18675
rect 1635 18645 1640 18675
rect 1600 18640 1640 18645
rect 1680 18675 1720 18680
rect 1680 18645 1685 18675
rect 1715 18645 1720 18675
rect 1680 18640 1720 18645
rect 1760 18675 1800 18680
rect 1760 18645 1765 18675
rect 1795 18645 1800 18675
rect 1760 18640 1800 18645
rect 1840 18675 1880 18680
rect 1840 18645 1845 18675
rect 1875 18645 1880 18675
rect 1840 18640 1880 18645
rect 1920 18675 1960 18680
rect 1920 18645 1925 18675
rect 1955 18645 1960 18675
rect 1920 18640 1960 18645
rect 2000 18675 2040 18680
rect 2000 18645 2005 18675
rect 2035 18645 2040 18675
rect 2000 18640 2040 18645
rect 2080 18675 2120 18680
rect 2080 18645 2085 18675
rect 2115 18645 2120 18675
rect 2080 18640 2120 18645
rect 2160 18675 2200 18680
rect 2160 18645 2165 18675
rect 2195 18645 2200 18675
rect 2160 18640 2200 18645
rect 2240 18675 2280 18680
rect 2240 18645 2245 18675
rect 2275 18645 2280 18675
rect 2240 18640 2280 18645
rect 2320 18675 2360 18680
rect 2320 18645 2325 18675
rect 2355 18645 2360 18675
rect 2320 18640 2360 18645
rect 2400 18675 2440 18680
rect 2400 18645 2405 18675
rect 2435 18645 2440 18675
rect 2400 18640 2440 18645
rect 2480 18675 2520 18680
rect 2480 18645 2485 18675
rect 2515 18645 2520 18675
rect 2480 18640 2520 18645
rect 2560 18675 2600 18680
rect 2560 18645 2565 18675
rect 2595 18645 2600 18675
rect 2560 18640 2600 18645
rect 2640 18675 2680 18680
rect 2640 18645 2645 18675
rect 2675 18645 2680 18675
rect 2640 18640 2680 18645
rect 2720 18675 2760 18680
rect 2720 18645 2725 18675
rect 2755 18645 2760 18675
rect 2720 18640 2760 18645
rect 2800 18675 2840 18680
rect 2800 18645 2805 18675
rect 2835 18645 2840 18675
rect 2800 18640 2840 18645
rect 2880 18675 2920 18680
rect 2880 18645 2885 18675
rect 2915 18645 2920 18675
rect 2880 18640 2920 18645
rect 2960 18675 3000 18680
rect 2960 18645 2965 18675
rect 2995 18645 3000 18675
rect 2960 18640 3000 18645
rect 3040 18675 3080 18680
rect 3040 18645 3045 18675
rect 3075 18645 3080 18675
rect 3040 18640 3080 18645
rect 3120 18675 3160 18680
rect 3120 18645 3125 18675
rect 3155 18645 3160 18675
rect 3120 18640 3160 18645
rect 3200 18675 3240 18680
rect 3200 18645 3205 18675
rect 3235 18645 3240 18675
rect 3200 18640 3240 18645
rect 3280 18675 3320 18680
rect 3280 18645 3285 18675
rect 3315 18645 3320 18675
rect 3280 18640 3320 18645
rect 3360 18675 3400 18680
rect 3360 18645 3365 18675
rect 3395 18645 3400 18675
rect 3360 18640 3400 18645
rect 3440 18675 3480 18680
rect 3440 18645 3445 18675
rect 3475 18645 3480 18675
rect 3440 18640 3480 18645
rect 3520 18675 3560 18680
rect 3520 18645 3525 18675
rect 3555 18645 3560 18675
rect 3520 18640 3560 18645
rect 3600 18675 3640 18680
rect 3600 18645 3605 18675
rect 3635 18645 3640 18675
rect 3600 18640 3640 18645
rect 3680 18675 3720 18680
rect 3680 18645 3685 18675
rect 3715 18645 3720 18675
rect 3680 18640 3720 18645
rect 3760 18675 3800 18680
rect 3760 18645 3765 18675
rect 3795 18645 3800 18675
rect 3760 18640 3800 18645
rect 3840 18675 3880 18680
rect 3840 18645 3845 18675
rect 3875 18645 3880 18675
rect 3840 18640 3880 18645
rect 3920 18675 3960 18680
rect 3920 18645 3925 18675
rect 3955 18645 3960 18675
rect 3920 18640 3960 18645
rect 4000 18675 4040 18680
rect 4000 18645 4005 18675
rect 4035 18645 4040 18675
rect 4000 18640 4040 18645
rect 4080 18675 4120 18680
rect 4080 18645 4085 18675
rect 4115 18645 4120 18675
rect 4080 18640 4120 18645
rect 4160 18675 4200 18680
rect 4160 18645 4165 18675
rect 4195 18645 4200 18675
rect 4160 18640 4200 18645
rect 6240 18675 6280 18680
rect 6240 18645 6245 18675
rect 6275 18645 6280 18675
rect 6240 18640 6280 18645
rect 6320 18675 6360 18680
rect 6320 18645 6325 18675
rect 6355 18645 6360 18675
rect 6320 18640 6360 18645
rect 6400 18675 6440 18680
rect 6400 18645 6405 18675
rect 6435 18645 6440 18675
rect 6400 18640 6440 18645
rect 6480 18675 6520 18680
rect 6480 18645 6485 18675
rect 6515 18645 6520 18675
rect 6480 18640 6520 18645
rect 6560 18675 6600 18680
rect 6560 18645 6565 18675
rect 6595 18645 6600 18675
rect 6560 18640 6600 18645
rect 6640 18675 6680 18680
rect 6640 18645 6645 18675
rect 6675 18645 6680 18675
rect 6640 18640 6680 18645
rect 6720 18675 6760 18680
rect 6720 18645 6725 18675
rect 6755 18645 6760 18675
rect 6720 18640 6760 18645
rect 6800 18675 6840 18680
rect 6800 18645 6805 18675
rect 6835 18645 6840 18675
rect 6800 18640 6840 18645
rect 6880 18675 6920 18680
rect 6880 18645 6885 18675
rect 6915 18645 6920 18675
rect 6880 18640 6920 18645
rect 6960 18675 7000 18680
rect 6960 18645 6965 18675
rect 6995 18645 7000 18675
rect 6960 18640 7000 18645
rect 7040 18675 7080 18680
rect 7040 18645 7045 18675
rect 7075 18645 7080 18675
rect 7040 18640 7080 18645
rect 7120 18675 7160 18680
rect 7120 18645 7125 18675
rect 7155 18645 7160 18675
rect 7120 18640 7160 18645
rect 7200 18675 7240 18680
rect 7200 18645 7205 18675
rect 7235 18645 7240 18675
rect 7200 18640 7240 18645
rect 7280 18675 7320 18680
rect 7280 18645 7285 18675
rect 7315 18645 7320 18675
rect 7280 18640 7320 18645
rect 7360 18675 7400 18680
rect 7360 18645 7365 18675
rect 7395 18645 7400 18675
rect 7360 18640 7400 18645
rect 7440 18675 7480 18680
rect 7440 18645 7445 18675
rect 7475 18645 7480 18675
rect 7440 18640 7480 18645
rect 7520 18675 7560 18680
rect 7520 18645 7525 18675
rect 7555 18645 7560 18675
rect 7520 18640 7560 18645
rect 7600 18675 7640 18680
rect 7600 18645 7605 18675
rect 7635 18645 7640 18675
rect 7600 18640 7640 18645
rect 7680 18675 7720 18680
rect 7680 18645 7685 18675
rect 7715 18645 7720 18675
rect 7680 18640 7720 18645
rect 7760 18675 7800 18680
rect 7760 18645 7765 18675
rect 7795 18645 7800 18675
rect 7760 18640 7800 18645
rect 7840 18675 7880 18680
rect 7840 18645 7845 18675
rect 7875 18645 7880 18675
rect 7840 18640 7880 18645
rect 7920 18675 7960 18680
rect 7920 18645 7925 18675
rect 7955 18645 7960 18675
rect 7920 18640 7960 18645
rect 8000 18675 8040 18680
rect 8000 18645 8005 18675
rect 8035 18645 8040 18675
rect 8000 18640 8040 18645
rect 8080 18675 8120 18680
rect 8080 18645 8085 18675
rect 8115 18645 8120 18675
rect 8080 18640 8120 18645
rect 8160 18675 8200 18680
rect 8160 18645 8165 18675
rect 8195 18645 8200 18675
rect 8160 18640 8200 18645
rect 8240 18675 8280 18680
rect 8240 18645 8245 18675
rect 8275 18645 8280 18675
rect 8240 18640 8280 18645
rect 8320 18675 8360 18680
rect 8320 18645 8325 18675
rect 8355 18645 8360 18675
rect 8320 18640 8360 18645
rect 8400 18675 8440 18680
rect 8400 18645 8405 18675
rect 8435 18645 8440 18675
rect 8400 18640 8440 18645
rect 8480 18675 8520 18680
rect 8480 18645 8485 18675
rect 8515 18645 8520 18675
rect 8480 18640 8520 18645
rect 8560 18675 8600 18680
rect 8560 18645 8565 18675
rect 8595 18645 8600 18675
rect 8560 18640 8600 18645
rect 8640 18675 8680 18680
rect 8640 18645 8645 18675
rect 8675 18645 8680 18675
rect 8640 18640 8680 18645
rect 8720 18675 8760 18680
rect 8720 18645 8725 18675
rect 8755 18645 8760 18675
rect 8720 18640 8760 18645
rect 8800 18675 8840 18680
rect 8800 18645 8805 18675
rect 8835 18645 8840 18675
rect 8800 18640 8840 18645
rect 8880 18675 8920 18680
rect 8880 18645 8885 18675
rect 8915 18645 8920 18675
rect 8880 18640 8920 18645
rect 8960 18675 9000 18680
rect 8960 18645 8965 18675
rect 8995 18645 9000 18675
rect 8960 18640 9000 18645
rect 9040 18675 9080 18680
rect 9040 18645 9045 18675
rect 9075 18645 9080 18675
rect 9040 18640 9080 18645
rect 9120 18675 9160 18680
rect 9120 18645 9125 18675
rect 9155 18645 9160 18675
rect 9120 18640 9160 18645
rect 9200 18675 9240 18680
rect 9200 18645 9205 18675
rect 9235 18645 9240 18675
rect 9200 18640 9240 18645
rect 9280 18675 9320 18680
rect 9280 18645 9285 18675
rect 9315 18645 9320 18675
rect 9280 18640 9320 18645
rect 9360 18675 9400 18680
rect 9360 18645 9365 18675
rect 9395 18645 9400 18675
rect 9360 18640 9400 18645
rect 9440 18675 9480 18680
rect 9440 18645 9445 18675
rect 9475 18645 9480 18675
rect 9440 18640 9480 18645
rect 11560 18675 11600 18680
rect 11560 18645 11565 18675
rect 11595 18645 11600 18675
rect 11560 18640 11600 18645
rect 11640 18675 11680 18680
rect 11640 18645 11645 18675
rect 11675 18645 11680 18675
rect 11640 18640 11680 18645
rect 11720 18675 11760 18680
rect 11720 18645 11725 18675
rect 11755 18645 11760 18675
rect 11720 18640 11760 18645
rect 11800 18675 11840 18680
rect 11800 18645 11805 18675
rect 11835 18645 11840 18675
rect 11800 18640 11840 18645
rect 11880 18675 11920 18680
rect 11880 18645 11885 18675
rect 11915 18645 11920 18675
rect 11880 18640 11920 18645
rect 11960 18675 12000 18680
rect 11960 18645 11965 18675
rect 11995 18645 12000 18675
rect 11960 18640 12000 18645
rect 12040 18675 12080 18680
rect 12040 18645 12045 18675
rect 12075 18645 12080 18675
rect 12040 18640 12080 18645
rect 12120 18675 12160 18680
rect 12120 18645 12125 18675
rect 12155 18645 12160 18675
rect 12120 18640 12160 18645
rect 12200 18675 12240 18680
rect 12200 18645 12205 18675
rect 12235 18645 12240 18675
rect 12200 18640 12240 18645
rect 12280 18675 12320 18680
rect 12280 18645 12285 18675
rect 12315 18645 12320 18675
rect 12280 18640 12320 18645
rect 12360 18675 12400 18680
rect 12360 18645 12365 18675
rect 12395 18645 12400 18675
rect 12360 18640 12400 18645
rect 12440 18675 12480 18680
rect 12440 18645 12445 18675
rect 12475 18645 12480 18675
rect 12440 18640 12480 18645
rect 12520 18675 12560 18680
rect 12520 18645 12525 18675
rect 12555 18645 12560 18675
rect 12520 18640 12560 18645
rect 12600 18675 12640 18680
rect 12600 18645 12605 18675
rect 12635 18645 12640 18675
rect 12600 18640 12640 18645
rect 12680 18675 12720 18680
rect 12680 18645 12685 18675
rect 12715 18645 12720 18675
rect 12680 18640 12720 18645
rect 12760 18675 12800 18680
rect 12760 18645 12765 18675
rect 12795 18645 12800 18675
rect 12760 18640 12800 18645
rect 12840 18675 12880 18680
rect 12840 18645 12845 18675
rect 12875 18645 12880 18675
rect 12840 18640 12880 18645
rect 12920 18675 12960 18680
rect 12920 18645 12925 18675
rect 12955 18645 12960 18675
rect 12920 18640 12960 18645
rect 13000 18675 13040 18680
rect 13000 18645 13005 18675
rect 13035 18645 13040 18675
rect 13000 18640 13040 18645
rect 13080 18675 13120 18680
rect 13080 18645 13085 18675
rect 13115 18645 13120 18675
rect 13080 18640 13120 18645
rect 13160 18675 13200 18680
rect 13160 18645 13165 18675
rect 13195 18645 13200 18675
rect 13160 18640 13200 18645
rect 13240 18675 13280 18680
rect 13240 18645 13245 18675
rect 13275 18645 13280 18675
rect 13240 18640 13280 18645
rect 13320 18675 13360 18680
rect 13320 18645 13325 18675
rect 13355 18645 13360 18675
rect 13320 18640 13360 18645
rect 13400 18675 13440 18680
rect 13400 18645 13405 18675
rect 13435 18645 13440 18675
rect 13400 18640 13440 18645
rect 13480 18675 13520 18680
rect 13480 18645 13485 18675
rect 13515 18645 13520 18675
rect 13480 18640 13520 18645
rect 13560 18675 13600 18680
rect 13560 18645 13565 18675
rect 13595 18645 13600 18675
rect 13560 18640 13600 18645
rect 13640 18675 13680 18680
rect 13640 18645 13645 18675
rect 13675 18645 13680 18675
rect 13640 18640 13680 18645
rect 13720 18675 13760 18680
rect 13720 18645 13725 18675
rect 13755 18645 13760 18675
rect 13720 18640 13760 18645
rect 13800 18675 13840 18680
rect 13800 18645 13805 18675
rect 13835 18645 13840 18675
rect 13800 18640 13840 18645
rect 13880 18675 13920 18680
rect 13880 18645 13885 18675
rect 13915 18645 13920 18675
rect 13880 18640 13920 18645
rect 13960 18675 14000 18680
rect 13960 18645 13965 18675
rect 13995 18645 14000 18675
rect 13960 18640 14000 18645
rect 14040 18675 14080 18680
rect 14040 18645 14045 18675
rect 14075 18645 14080 18675
rect 14040 18640 14080 18645
rect 14120 18675 14160 18680
rect 14120 18645 14125 18675
rect 14155 18645 14160 18675
rect 14120 18640 14160 18645
rect 14200 18675 14240 18680
rect 14200 18645 14205 18675
rect 14235 18645 14240 18675
rect 14200 18640 14240 18645
rect 14280 18675 14320 18680
rect 14280 18645 14285 18675
rect 14315 18645 14320 18675
rect 14280 18640 14320 18645
rect 14360 18675 14400 18680
rect 14360 18645 14365 18675
rect 14395 18645 14400 18675
rect 14360 18640 14400 18645
rect 14440 18675 14480 18680
rect 14440 18645 14445 18675
rect 14475 18645 14480 18675
rect 14440 18640 14480 18645
rect 14520 18675 14560 18680
rect 14520 18645 14525 18675
rect 14555 18645 14560 18675
rect 14520 18640 14560 18645
rect 14600 18675 14640 18680
rect 14600 18645 14605 18675
rect 14635 18645 14640 18675
rect 14600 18640 14640 18645
rect 14680 18675 14720 18680
rect 14680 18645 14685 18675
rect 14715 18645 14720 18675
rect 14680 18640 14720 18645
rect 16760 18675 16800 18680
rect 16760 18645 16765 18675
rect 16795 18645 16800 18675
rect 16760 18640 16800 18645
rect 16840 18675 16880 18680
rect 16840 18645 16845 18675
rect 16875 18645 16880 18675
rect 16840 18640 16880 18645
rect 16920 18675 16960 18680
rect 16920 18645 16925 18675
rect 16955 18645 16960 18675
rect 16920 18640 16960 18645
rect 17000 18675 17040 18680
rect 17000 18645 17005 18675
rect 17035 18645 17040 18675
rect 17000 18640 17040 18645
rect 17080 18675 17120 18680
rect 17080 18645 17085 18675
rect 17115 18645 17120 18675
rect 17080 18640 17120 18645
rect 17160 18675 17200 18680
rect 17160 18645 17165 18675
rect 17195 18645 17200 18675
rect 17160 18640 17200 18645
rect 17240 18675 17280 18680
rect 17240 18645 17245 18675
rect 17275 18645 17280 18675
rect 17240 18640 17280 18645
rect 17320 18675 17360 18680
rect 17320 18645 17325 18675
rect 17355 18645 17360 18675
rect 17320 18640 17360 18645
rect 17400 18675 17440 18680
rect 17400 18645 17405 18675
rect 17435 18645 17440 18675
rect 17400 18640 17440 18645
rect 17480 18675 17520 18680
rect 17480 18645 17485 18675
rect 17515 18645 17520 18675
rect 17480 18640 17520 18645
rect 17560 18675 17600 18680
rect 17560 18645 17565 18675
rect 17595 18645 17600 18675
rect 17560 18640 17600 18645
rect 17640 18675 17680 18680
rect 17640 18645 17645 18675
rect 17675 18645 17680 18675
rect 17640 18640 17680 18645
rect 17720 18675 17760 18680
rect 17720 18645 17725 18675
rect 17755 18645 17760 18675
rect 17720 18640 17760 18645
rect 17800 18675 17840 18680
rect 17800 18645 17805 18675
rect 17835 18645 17840 18675
rect 17800 18640 17840 18645
rect 17880 18675 17920 18680
rect 17880 18645 17885 18675
rect 17915 18645 17920 18675
rect 17880 18640 17920 18645
rect 17960 18675 18000 18680
rect 17960 18645 17965 18675
rect 17995 18645 18000 18675
rect 17960 18640 18000 18645
rect 18040 18675 18080 18680
rect 18040 18645 18045 18675
rect 18075 18645 18080 18675
rect 18040 18640 18080 18645
rect 18120 18675 18160 18680
rect 18120 18645 18125 18675
rect 18155 18645 18160 18675
rect 18120 18640 18160 18645
rect 18200 18675 18240 18680
rect 18200 18645 18205 18675
rect 18235 18645 18240 18675
rect 18200 18640 18240 18645
rect 18280 18675 18320 18680
rect 18280 18645 18285 18675
rect 18315 18645 18320 18675
rect 18280 18640 18320 18645
rect 18360 18675 18400 18680
rect 18360 18645 18365 18675
rect 18395 18645 18400 18675
rect 18360 18640 18400 18645
rect 18440 18675 18480 18680
rect 18440 18645 18445 18675
rect 18475 18645 18480 18675
rect 18440 18640 18480 18645
rect 18520 18675 18560 18680
rect 18520 18645 18525 18675
rect 18555 18645 18560 18675
rect 18520 18640 18560 18645
rect 18600 18675 18640 18680
rect 18600 18645 18605 18675
rect 18635 18645 18640 18675
rect 18600 18640 18640 18645
rect 18680 18675 18720 18680
rect 18680 18645 18685 18675
rect 18715 18645 18720 18675
rect 18680 18640 18720 18645
rect 18760 18675 18800 18680
rect 18760 18645 18765 18675
rect 18795 18645 18800 18675
rect 18760 18640 18800 18645
rect 18840 18675 18880 18680
rect 18840 18645 18845 18675
rect 18875 18645 18880 18675
rect 18840 18640 18880 18645
rect 18920 18675 18960 18680
rect 18920 18645 18925 18675
rect 18955 18645 18960 18675
rect 18920 18640 18960 18645
rect 19000 18675 19040 18680
rect 19000 18645 19005 18675
rect 19035 18645 19040 18675
rect 19000 18640 19040 18645
rect 19080 18675 19120 18680
rect 19080 18645 19085 18675
rect 19115 18645 19120 18675
rect 19080 18640 19120 18645
rect 19160 18675 19200 18680
rect 19160 18645 19165 18675
rect 19195 18645 19200 18675
rect 19160 18640 19200 18645
rect 19240 18675 19280 18680
rect 19240 18645 19245 18675
rect 19275 18645 19280 18675
rect 19240 18640 19280 18645
rect 19320 18675 19360 18680
rect 19320 18645 19325 18675
rect 19355 18645 19360 18675
rect 19320 18640 19360 18645
rect 19400 18675 19440 18680
rect 19400 18645 19405 18675
rect 19435 18645 19440 18675
rect 19400 18640 19440 18645
rect 19480 18675 19520 18680
rect 19480 18645 19485 18675
rect 19515 18645 19520 18675
rect 19480 18640 19520 18645
rect 19560 18675 19600 18680
rect 19560 18645 19565 18675
rect 19595 18645 19600 18675
rect 19560 18640 19600 18645
rect 19640 18675 19680 18680
rect 19640 18645 19645 18675
rect 19675 18645 19680 18675
rect 19640 18640 19680 18645
rect 19720 18675 19760 18680
rect 19720 18645 19725 18675
rect 19755 18645 19760 18675
rect 19720 18640 19760 18645
rect 19800 18675 19840 18680
rect 19800 18645 19805 18675
rect 19835 18645 19840 18675
rect 19800 18640 19840 18645
rect 19880 18675 19920 18680
rect 19880 18645 19885 18675
rect 19915 18645 19920 18675
rect 19880 18640 19920 18645
rect 19960 18675 20000 18680
rect 19960 18645 19965 18675
rect 19995 18645 20000 18675
rect 19960 18640 20000 18645
rect 20040 18675 20080 18680
rect 20040 18645 20045 18675
rect 20075 18645 20080 18675
rect 20040 18640 20080 18645
rect 20120 18675 20160 18680
rect 20120 18645 20125 18675
rect 20155 18645 20160 18675
rect 20120 18640 20160 18645
rect 20200 18675 20240 18680
rect 20200 18645 20205 18675
rect 20235 18645 20240 18675
rect 20200 18640 20240 18645
rect 20280 18675 20320 18680
rect 20280 18645 20285 18675
rect 20315 18645 20320 18675
rect 20280 18640 20320 18645
rect 20360 18675 20400 18680
rect 20360 18645 20365 18675
rect 20395 18645 20400 18675
rect 20360 18640 20400 18645
rect 20440 18675 20480 18680
rect 20440 18645 20445 18675
rect 20475 18645 20480 18675
rect 20440 18640 20480 18645
rect 20520 18675 20560 18680
rect 20520 18645 20525 18675
rect 20555 18645 20560 18675
rect 20520 18640 20560 18645
rect 20600 18675 20640 18680
rect 20600 18645 20605 18675
rect 20635 18645 20640 18675
rect 20600 18640 20640 18645
rect 20680 18675 20720 18680
rect 20680 18645 20685 18675
rect 20715 18645 20720 18675
rect 20680 18640 20720 18645
rect 20760 18675 20800 18680
rect 20760 18645 20765 18675
rect 20795 18645 20800 18675
rect 20760 18640 20800 18645
rect 20840 18675 20880 18680
rect 20840 18645 20845 18675
rect 20875 18645 20880 18675
rect 20840 18640 20880 18645
rect 20920 18675 20960 18680
rect 20920 18645 20925 18675
rect 20955 18645 20960 18675
rect 20920 18640 20960 18645
rect 0 18515 40 18520
rect 0 18485 5 18515
rect 35 18485 40 18515
rect 0 18480 40 18485
rect 80 18515 120 18520
rect 80 18485 85 18515
rect 115 18485 120 18515
rect 80 18480 120 18485
rect 160 18515 200 18520
rect 160 18485 165 18515
rect 195 18485 200 18515
rect 160 18480 200 18485
rect 240 18515 280 18520
rect 240 18485 245 18515
rect 275 18485 280 18515
rect 240 18480 280 18485
rect 320 18515 360 18520
rect 320 18485 325 18515
rect 355 18485 360 18515
rect 320 18480 360 18485
rect 400 18515 440 18520
rect 400 18485 405 18515
rect 435 18485 440 18515
rect 400 18480 440 18485
rect 480 18515 520 18520
rect 480 18485 485 18515
rect 515 18485 520 18515
rect 480 18480 520 18485
rect 560 18515 600 18520
rect 560 18485 565 18515
rect 595 18485 600 18515
rect 560 18480 600 18485
rect 640 18515 680 18520
rect 640 18485 645 18515
rect 675 18485 680 18515
rect 640 18480 680 18485
rect 720 18515 760 18520
rect 720 18485 725 18515
rect 755 18485 760 18515
rect 720 18480 760 18485
rect 800 18515 840 18520
rect 800 18485 805 18515
rect 835 18485 840 18515
rect 800 18480 840 18485
rect 880 18515 920 18520
rect 880 18485 885 18515
rect 915 18485 920 18515
rect 880 18480 920 18485
rect 960 18515 1000 18520
rect 960 18485 965 18515
rect 995 18485 1000 18515
rect 960 18480 1000 18485
rect 1040 18515 1080 18520
rect 1040 18485 1045 18515
rect 1075 18485 1080 18515
rect 1040 18480 1080 18485
rect 1120 18515 1160 18520
rect 1120 18485 1125 18515
rect 1155 18485 1160 18515
rect 1120 18480 1160 18485
rect 1200 18515 1240 18520
rect 1200 18485 1205 18515
rect 1235 18485 1240 18515
rect 1200 18480 1240 18485
rect 1280 18515 1320 18520
rect 1280 18485 1285 18515
rect 1315 18485 1320 18515
rect 1280 18480 1320 18485
rect 1360 18515 1400 18520
rect 1360 18485 1365 18515
rect 1395 18485 1400 18515
rect 1360 18480 1400 18485
rect 1440 18515 1480 18520
rect 1440 18485 1445 18515
rect 1475 18485 1480 18515
rect 1440 18480 1480 18485
rect 1520 18515 1560 18520
rect 1520 18485 1525 18515
rect 1555 18485 1560 18515
rect 1520 18480 1560 18485
rect 1600 18515 1640 18520
rect 1600 18485 1605 18515
rect 1635 18485 1640 18515
rect 1600 18480 1640 18485
rect 1680 18515 1720 18520
rect 1680 18485 1685 18515
rect 1715 18485 1720 18515
rect 1680 18480 1720 18485
rect 1760 18515 1800 18520
rect 1760 18485 1765 18515
rect 1795 18485 1800 18515
rect 1760 18480 1800 18485
rect 1840 18515 1880 18520
rect 1840 18485 1845 18515
rect 1875 18485 1880 18515
rect 1840 18480 1880 18485
rect 1920 18515 1960 18520
rect 1920 18485 1925 18515
rect 1955 18485 1960 18515
rect 1920 18480 1960 18485
rect 2000 18515 2040 18520
rect 2000 18485 2005 18515
rect 2035 18485 2040 18515
rect 2000 18480 2040 18485
rect 2080 18515 2120 18520
rect 2080 18485 2085 18515
rect 2115 18485 2120 18515
rect 2080 18480 2120 18485
rect 2160 18515 2200 18520
rect 2160 18485 2165 18515
rect 2195 18485 2200 18515
rect 2160 18480 2200 18485
rect 2240 18515 2280 18520
rect 2240 18485 2245 18515
rect 2275 18485 2280 18515
rect 2240 18480 2280 18485
rect 2320 18515 2360 18520
rect 2320 18485 2325 18515
rect 2355 18485 2360 18515
rect 2320 18480 2360 18485
rect 2400 18515 2440 18520
rect 2400 18485 2405 18515
rect 2435 18485 2440 18515
rect 2400 18480 2440 18485
rect 2480 18515 2520 18520
rect 2480 18485 2485 18515
rect 2515 18485 2520 18515
rect 2480 18480 2520 18485
rect 2560 18515 2600 18520
rect 2560 18485 2565 18515
rect 2595 18485 2600 18515
rect 2560 18480 2600 18485
rect 2640 18515 2680 18520
rect 2640 18485 2645 18515
rect 2675 18485 2680 18515
rect 2640 18480 2680 18485
rect 2720 18515 2760 18520
rect 2720 18485 2725 18515
rect 2755 18485 2760 18515
rect 2720 18480 2760 18485
rect 2800 18515 2840 18520
rect 2800 18485 2805 18515
rect 2835 18485 2840 18515
rect 2800 18480 2840 18485
rect 2880 18515 2920 18520
rect 2880 18485 2885 18515
rect 2915 18485 2920 18515
rect 2880 18480 2920 18485
rect 2960 18515 3000 18520
rect 2960 18485 2965 18515
rect 2995 18485 3000 18515
rect 2960 18480 3000 18485
rect 3040 18515 3080 18520
rect 3040 18485 3045 18515
rect 3075 18485 3080 18515
rect 3040 18480 3080 18485
rect 3120 18515 3160 18520
rect 3120 18485 3125 18515
rect 3155 18485 3160 18515
rect 3120 18480 3160 18485
rect 3200 18515 3240 18520
rect 3200 18485 3205 18515
rect 3235 18485 3240 18515
rect 3200 18480 3240 18485
rect 3280 18515 3320 18520
rect 3280 18485 3285 18515
rect 3315 18485 3320 18515
rect 3280 18480 3320 18485
rect 3360 18515 3400 18520
rect 3360 18485 3365 18515
rect 3395 18485 3400 18515
rect 3360 18480 3400 18485
rect 3440 18515 3480 18520
rect 3440 18485 3445 18515
rect 3475 18485 3480 18515
rect 3440 18480 3480 18485
rect 3520 18515 3560 18520
rect 3520 18485 3525 18515
rect 3555 18485 3560 18515
rect 3520 18480 3560 18485
rect 3600 18515 3640 18520
rect 3600 18485 3605 18515
rect 3635 18485 3640 18515
rect 3600 18480 3640 18485
rect 3680 18515 3720 18520
rect 3680 18485 3685 18515
rect 3715 18485 3720 18515
rect 3680 18480 3720 18485
rect 3760 18515 3800 18520
rect 3760 18485 3765 18515
rect 3795 18485 3800 18515
rect 3760 18480 3800 18485
rect 3840 18515 3880 18520
rect 3840 18485 3845 18515
rect 3875 18485 3880 18515
rect 3840 18480 3880 18485
rect 3920 18515 3960 18520
rect 3920 18485 3925 18515
rect 3955 18485 3960 18515
rect 3920 18480 3960 18485
rect 4000 18515 4040 18520
rect 4000 18485 4005 18515
rect 4035 18485 4040 18515
rect 4000 18480 4040 18485
rect 4080 18515 4120 18520
rect 4080 18485 4085 18515
rect 4115 18485 4120 18515
rect 4080 18480 4120 18485
rect 4160 18515 4200 18520
rect 4160 18485 4165 18515
rect 4195 18485 4200 18515
rect 4160 18480 4200 18485
rect 6240 18515 6280 18520
rect 6240 18485 6245 18515
rect 6275 18485 6280 18515
rect 6240 18480 6280 18485
rect 6320 18515 6360 18520
rect 6320 18485 6325 18515
rect 6355 18485 6360 18515
rect 6320 18480 6360 18485
rect 6400 18515 6440 18520
rect 6400 18485 6405 18515
rect 6435 18485 6440 18515
rect 6400 18480 6440 18485
rect 6480 18515 6520 18520
rect 6480 18485 6485 18515
rect 6515 18485 6520 18515
rect 6480 18480 6520 18485
rect 6560 18515 6600 18520
rect 6560 18485 6565 18515
rect 6595 18485 6600 18515
rect 6560 18480 6600 18485
rect 6640 18515 6680 18520
rect 6640 18485 6645 18515
rect 6675 18485 6680 18515
rect 6640 18480 6680 18485
rect 6720 18515 6760 18520
rect 6720 18485 6725 18515
rect 6755 18485 6760 18515
rect 6720 18480 6760 18485
rect 6800 18515 6840 18520
rect 6800 18485 6805 18515
rect 6835 18485 6840 18515
rect 6800 18480 6840 18485
rect 6880 18515 6920 18520
rect 6880 18485 6885 18515
rect 6915 18485 6920 18515
rect 6880 18480 6920 18485
rect 6960 18515 7000 18520
rect 6960 18485 6965 18515
rect 6995 18485 7000 18515
rect 6960 18480 7000 18485
rect 7040 18515 7080 18520
rect 7040 18485 7045 18515
rect 7075 18485 7080 18515
rect 7040 18480 7080 18485
rect 7120 18515 7160 18520
rect 7120 18485 7125 18515
rect 7155 18485 7160 18515
rect 7120 18480 7160 18485
rect 7200 18515 7240 18520
rect 7200 18485 7205 18515
rect 7235 18485 7240 18515
rect 7200 18480 7240 18485
rect 7280 18515 7320 18520
rect 7280 18485 7285 18515
rect 7315 18485 7320 18515
rect 7280 18480 7320 18485
rect 7360 18515 7400 18520
rect 7360 18485 7365 18515
rect 7395 18485 7400 18515
rect 7360 18480 7400 18485
rect 7440 18515 7480 18520
rect 7440 18485 7445 18515
rect 7475 18485 7480 18515
rect 7440 18480 7480 18485
rect 7520 18515 7560 18520
rect 7520 18485 7525 18515
rect 7555 18485 7560 18515
rect 7520 18480 7560 18485
rect 7600 18515 7640 18520
rect 7600 18485 7605 18515
rect 7635 18485 7640 18515
rect 7600 18480 7640 18485
rect 7680 18515 7720 18520
rect 7680 18485 7685 18515
rect 7715 18485 7720 18515
rect 7680 18480 7720 18485
rect 7760 18515 7800 18520
rect 7760 18485 7765 18515
rect 7795 18485 7800 18515
rect 7760 18480 7800 18485
rect 7840 18515 7880 18520
rect 7840 18485 7845 18515
rect 7875 18485 7880 18515
rect 7840 18480 7880 18485
rect 7920 18515 7960 18520
rect 7920 18485 7925 18515
rect 7955 18485 7960 18515
rect 7920 18480 7960 18485
rect 8000 18515 8040 18520
rect 8000 18485 8005 18515
rect 8035 18485 8040 18515
rect 8000 18480 8040 18485
rect 8080 18515 8120 18520
rect 8080 18485 8085 18515
rect 8115 18485 8120 18515
rect 8080 18480 8120 18485
rect 8160 18515 8200 18520
rect 8160 18485 8165 18515
rect 8195 18485 8200 18515
rect 8160 18480 8200 18485
rect 8240 18515 8280 18520
rect 8240 18485 8245 18515
rect 8275 18485 8280 18515
rect 8240 18480 8280 18485
rect 8320 18515 8360 18520
rect 8320 18485 8325 18515
rect 8355 18485 8360 18515
rect 8320 18480 8360 18485
rect 8400 18515 8440 18520
rect 8400 18485 8405 18515
rect 8435 18485 8440 18515
rect 8400 18480 8440 18485
rect 8480 18515 8520 18520
rect 8480 18485 8485 18515
rect 8515 18485 8520 18515
rect 8480 18480 8520 18485
rect 8560 18515 8600 18520
rect 8560 18485 8565 18515
rect 8595 18485 8600 18515
rect 8560 18480 8600 18485
rect 8640 18515 8680 18520
rect 8640 18485 8645 18515
rect 8675 18485 8680 18515
rect 8640 18480 8680 18485
rect 8720 18515 8760 18520
rect 8720 18485 8725 18515
rect 8755 18485 8760 18515
rect 8720 18480 8760 18485
rect 8800 18515 8840 18520
rect 8800 18485 8805 18515
rect 8835 18485 8840 18515
rect 8800 18480 8840 18485
rect 8880 18515 8920 18520
rect 8880 18485 8885 18515
rect 8915 18485 8920 18515
rect 8880 18480 8920 18485
rect 8960 18515 9000 18520
rect 8960 18485 8965 18515
rect 8995 18485 9000 18515
rect 8960 18480 9000 18485
rect 9040 18515 9080 18520
rect 9040 18485 9045 18515
rect 9075 18485 9080 18515
rect 9040 18480 9080 18485
rect 9120 18515 9160 18520
rect 9120 18485 9125 18515
rect 9155 18485 9160 18515
rect 9120 18480 9160 18485
rect 9200 18515 9240 18520
rect 9200 18485 9205 18515
rect 9235 18485 9240 18515
rect 9200 18480 9240 18485
rect 9280 18515 9320 18520
rect 9280 18485 9285 18515
rect 9315 18485 9320 18515
rect 9280 18480 9320 18485
rect 9360 18515 9400 18520
rect 9360 18485 9365 18515
rect 9395 18485 9400 18515
rect 9360 18480 9400 18485
rect 9440 18515 9480 18520
rect 9440 18485 9445 18515
rect 9475 18485 9480 18515
rect 9440 18480 9480 18485
rect 11560 18515 11600 18520
rect 11560 18485 11565 18515
rect 11595 18485 11600 18515
rect 11560 18480 11600 18485
rect 11640 18515 11680 18520
rect 11640 18485 11645 18515
rect 11675 18485 11680 18515
rect 11640 18480 11680 18485
rect 11720 18515 11760 18520
rect 11720 18485 11725 18515
rect 11755 18485 11760 18515
rect 11720 18480 11760 18485
rect 11800 18515 11840 18520
rect 11800 18485 11805 18515
rect 11835 18485 11840 18515
rect 11800 18480 11840 18485
rect 11880 18515 11920 18520
rect 11880 18485 11885 18515
rect 11915 18485 11920 18515
rect 11880 18480 11920 18485
rect 11960 18515 12000 18520
rect 11960 18485 11965 18515
rect 11995 18485 12000 18515
rect 11960 18480 12000 18485
rect 12040 18515 12080 18520
rect 12040 18485 12045 18515
rect 12075 18485 12080 18515
rect 12040 18480 12080 18485
rect 12120 18515 12160 18520
rect 12120 18485 12125 18515
rect 12155 18485 12160 18515
rect 12120 18480 12160 18485
rect 12200 18515 12240 18520
rect 12200 18485 12205 18515
rect 12235 18485 12240 18515
rect 12200 18480 12240 18485
rect 12280 18515 12320 18520
rect 12280 18485 12285 18515
rect 12315 18485 12320 18515
rect 12280 18480 12320 18485
rect 12360 18515 12400 18520
rect 12360 18485 12365 18515
rect 12395 18485 12400 18515
rect 12360 18480 12400 18485
rect 12440 18515 12480 18520
rect 12440 18485 12445 18515
rect 12475 18485 12480 18515
rect 12440 18480 12480 18485
rect 12520 18515 12560 18520
rect 12520 18485 12525 18515
rect 12555 18485 12560 18515
rect 12520 18480 12560 18485
rect 12600 18515 12640 18520
rect 12600 18485 12605 18515
rect 12635 18485 12640 18515
rect 12600 18480 12640 18485
rect 12680 18515 12720 18520
rect 12680 18485 12685 18515
rect 12715 18485 12720 18515
rect 12680 18480 12720 18485
rect 12760 18515 12800 18520
rect 12760 18485 12765 18515
rect 12795 18485 12800 18515
rect 12760 18480 12800 18485
rect 12840 18515 12880 18520
rect 12840 18485 12845 18515
rect 12875 18485 12880 18515
rect 12840 18480 12880 18485
rect 12920 18515 12960 18520
rect 12920 18485 12925 18515
rect 12955 18485 12960 18515
rect 12920 18480 12960 18485
rect 13000 18515 13040 18520
rect 13000 18485 13005 18515
rect 13035 18485 13040 18515
rect 13000 18480 13040 18485
rect 13080 18515 13120 18520
rect 13080 18485 13085 18515
rect 13115 18485 13120 18515
rect 13080 18480 13120 18485
rect 13160 18515 13200 18520
rect 13160 18485 13165 18515
rect 13195 18485 13200 18515
rect 13160 18480 13200 18485
rect 13240 18515 13280 18520
rect 13240 18485 13245 18515
rect 13275 18485 13280 18515
rect 13240 18480 13280 18485
rect 13320 18515 13360 18520
rect 13320 18485 13325 18515
rect 13355 18485 13360 18515
rect 13320 18480 13360 18485
rect 13400 18515 13440 18520
rect 13400 18485 13405 18515
rect 13435 18485 13440 18515
rect 13400 18480 13440 18485
rect 13480 18515 13520 18520
rect 13480 18485 13485 18515
rect 13515 18485 13520 18515
rect 13480 18480 13520 18485
rect 13560 18515 13600 18520
rect 13560 18485 13565 18515
rect 13595 18485 13600 18515
rect 13560 18480 13600 18485
rect 13640 18515 13680 18520
rect 13640 18485 13645 18515
rect 13675 18485 13680 18515
rect 13640 18480 13680 18485
rect 13720 18515 13760 18520
rect 13720 18485 13725 18515
rect 13755 18485 13760 18515
rect 13720 18480 13760 18485
rect 13800 18515 13840 18520
rect 13800 18485 13805 18515
rect 13835 18485 13840 18515
rect 13800 18480 13840 18485
rect 13880 18515 13920 18520
rect 13880 18485 13885 18515
rect 13915 18485 13920 18515
rect 13880 18480 13920 18485
rect 13960 18515 14000 18520
rect 13960 18485 13965 18515
rect 13995 18485 14000 18515
rect 13960 18480 14000 18485
rect 14040 18515 14080 18520
rect 14040 18485 14045 18515
rect 14075 18485 14080 18515
rect 14040 18480 14080 18485
rect 14120 18515 14160 18520
rect 14120 18485 14125 18515
rect 14155 18485 14160 18515
rect 14120 18480 14160 18485
rect 14200 18515 14240 18520
rect 14200 18485 14205 18515
rect 14235 18485 14240 18515
rect 14200 18480 14240 18485
rect 14280 18515 14320 18520
rect 14280 18485 14285 18515
rect 14315 18485 14320 18515
rect 14280 18480 14320 18485
rect 14360 18515 14400 18520
rect 14360 18485 14365 18515
rect 14395 18485 14400 18515
rect 14360 18480 14400 18485
rect 14440 18515 14480 18520
rect 14440 18485 14445 18515
rect 14475 18485 14480 18515
rect 14440 18480 14480 18485
rect 14520 18515 14560 18520
rect 14520 18485 14525 18515
rect 14555 18485 14560 18515
rect 14520 18480 14560 18485
rect 14600 18515 14640 18520
rect 14600 18485 14605 18515
rect 14635 18485 14640 18515
rect 14600 18480 14640 18485
rect 14680 18515 14720 18520
rect 14680 18485 14685 18515
rect 14715 18485 14720 18515
rect 14680 18480 14720 18485
rect 16760 18515 16800 18520
rect 16760 18485 16765 18515
rect 16795 18485 16800 18515
rect 16760 18480 16800 18485
rect 16840 18515 16880 18520
rect 16840 18485 16845 18515
rect 16875 18485 16880 18515
rect 16840 18480 16880 18485
rect 16920 18515 16960 18520
rect 16920 18485 16925 18515
rect 16955 18485 16960 18515
rect 16920 18480 16960 18485
rect 17000 18515 17040 18520
rect 17000 18485 17005 18515
rect 17035 18485 17040 18515
rect 17000 18480 17040 18485
rect 17080 18515 17120 18520
rect 17080 18485 17085 18515
rect 17115 18485 17120 18515
rect 17080 18480 17120 18485
rect 17160 18515 17200 18520
rect 17160 18485 17165 18515
rect 17195 18485 17200 18515
rect 17160 18480 17200 18485
rect 17240 18515 17280 18520
rect 17240 18485 17245 18515
rect 17275 18485 17280 18515
rect 17240 18480 17280 18485
rect 17320 18515 17360 18520
rect 17320 18485 17325 18515
rect 17355 18485 17360 18515
rect 17320 18480 17360 18485
rect 17400 18515 17440 18520
rect 17400 18485 17405 18515
rect 17435 18485 17440 18515
rect 17400 18480 17440 18485
rect 17480 18515 17520 18520
rect 17480 18485 17485 18515
rect 17515 18485 17520 18515
rect 17480 18480 17520 18485
rect 17560 18515 17600 18520
rect 17560 18485 17565 18515
rect 17595 18485 17600 18515
rect 17560 18480 17600 18485
rect 17640 18515 17680 18520
rect 17640 18485 17645 18515
rect 17675 18485 17680 18515
rect 17640 18480 17680 18485
rect 17720 18515 17760 18520
rect 17720 18485 17725 18515
rect 17755 18485 17760 18515
rect 17720 18480 17760 18485
rect 17800 18515 17840 18520
rect 17800 18485 17805 18515
rect 17835 18485 17840 18515
rect 17800 18480 17840 18485
rect 17880 18515 17920 18520
rect 17880 18485 17885 18515
rect 17915 18485 17920 18515
rect 17880 18480 17920 18485
rect 17960 18515 18000 18520
rect 17960 18485 17965 18515
rect 17995 18485 18000 18515
rect 17960 18480 18000 18485
rect 18040 18515 18080 18520
rect 18040 18485 18045 18515
rect 18075 18485 18080 18515
rect 18040 18480 18080 18485
rect 18120 18515 18160 18520
rect 18120 18485 18125 18515
rect 18155 18485 18160 18515
rect 18120 18480 18160 18485
rect 18200 18515 18240 18520
rect 18200 18485 18205 18515
rect 18235 18485 18240 18515
rect 18200 18480 18240 18485
rect 18280 18515 18320 18520
rect 18280 18485 18285 18515
rect 18315 18485 18320 18515
rect 18280 18480 18320 18485
rect 18360 18515 18400 18520
rect 18360 18485 18365 18515
rect 18395 18485 18400 18515
rect 18360 18480 18400 18485
rect 18440 18515 18480 18520
rect 18440 18485 18445 18515
rect 18475 18485 18480 18515
rect 18440 18480 18480 18485
rect 18520 18515 18560 18520
rect 18520 18485 18525 18515
rect 18555 18485 18560 18515
rect 18520 18480 18560 18485
rect 18600 18515 18640 18520
rect 18600 18485 18605 18515
rect 18635 18485 18640 18515
rect 18600 18480 18640 18485
rect 18680 18515 18720 18520
rect 18680 18485 18685 18515
rect 18715 18485 18720 18515
rect 18680 18480 18720 18485
rect 18760 18515 18800 18520
rect 18760 18485 18765 18515
rect 18795 18485 18800 18515
rect 18760 18480 18800 18485
rect 18840 18515 18880 18520
rect 18840 18485 18845 18515
rect 18875 18485 18880 18515
rect 18840 18480 18880 18485
rect 18920 18515 18960 18520
rect 18920 18485 18925 18515
rect 18955 18485 18960 18515
rect 18920 18480 18960 18485
rect 19000 18515 19040 18520
rect 19000 18485 19005 18515
rect 19035 18485 19040 18515
rect 19000 18480 19040 18485
rect 19080 18515 19120 18520
rect 19080 18485 19085 18515
rect 19115 18485 19120 18515
rect 19080 18480 19120 18485
rect 19160 18515 19200 18520
rect 19160 18485 19165 18515
rect 19195 18485 19200 18515
rect 19160 18480 19200 18485
rect 19240 18515 19280 18520
rect 19240 18485 19245 18515
rect 19275 18485 19280 18515
rect 19240 18480 19280 18485
rect 19320 18515 19360 18520
rect 19320 18485 19325 18515
rect 19355 18485 19360 18515
rect 19320 18480 19360 18485
rect 19400 18515 19440 18520
rect 19400 18485 19405 18515
rect 19435 18485 19440 18515
rect 19400 18480 19440 18485
rect 19480 18515 19520 18520
rect 19480 18485 19485 18515
rect 19515 18485 19520 18515
rect 19480 18480 19520 18485
rect 19560 18515 19600 18520
rect 19560 18485 19565 18515
rect 19595 18485 19600 18515
rect 19560 18480 19600 18485
rect 19640 18515 19680 18520
rect 19640 18485 19645 18515
rect 19675 18485 19680 18515
rect 19640 18480 19680 18485
rect 19720 18515 19760 18520
rect 19720 18485 19725 18515
rect 19755 18485 19760 18515
rect 19720 18480 19760 18485
rect 19800 18515 19840 18520
rect 19800 18485 19805 18515
rect 19835 18485 19840 18515
rect 19800 18480 19840 18485
rect 19880 18515 19920 18520
rect 19880 18485 19885 18515
rect 19915 18485 19920 18515
rect 19880 18480 19920 18485
rect 19960 18515 20000 18520
rect 19960 18485 19965 18515
rect 19995 18485 20000 18515
rect 19960 18480 20000 18485
rect 20040 18515 20080 18520
rect 20040 18485 20045 18515
rect 20075 18485 20080 18515
rect 20040 18480 20080 18485
rect 20120 18515 20160 18520
rect 20120 18485 20125 18515
rect 20155 18485 20160 18515
rect 20120 18480 20160 18485
rect 20200 18515 20240 18520
rect 20200 18485 20205 18515
rect 20235 18485 20240 18515
rect 20200 18480 20240 18485
rect 20280 18515 20320 18520
rect 20280 18485 20285 18515
rect 20315 18485 20320 18515
rect 20280 18480 20320 18485
rect 20360 18515 20400 18520
rect 20360 18485 20365 18515
rect 20395 18485 20400 18515
rect 20360 18480 20400 18485
rect 20440 18515 20480 18520
rect 20440 18485 20445 18515
rect 20475 18485 20480 18515
rect 20440 18480 20480 18485
rect 20520 18515 20560 18520
rect 20520 18485 20525 18515
rect 20555 18485 20560 18515
rect 20520 18480 20560 18485
rect 20600 18515 20640 18520
rect 20600 18485 20605 18515
rect 20635 18485 20640 18515
rect 20600 18480 20640 18485
rect 20680 18515 20720 18520
rect 20680 18485 20685 18515
rect 20715 18485 20720 18515
rect 20680 18480 20720 18485
rect 20760 18515 20800 18520
rect 20760 18485 20765 18515
rect 20795 18485 20800 18515
rect 20760 18480 20800 18485
rect 20840 18515 20880 18520
rect 20840 18485 20845 18515
rect 20875 18485 20880 18515
rect 20840 18480 20880 18485
rect 20920 18515 20960 18520
rect 20920 18485 20925 18515
rect 20955 18485 20960 18515
rect 20920 18480 20960 18485
rect 0 18435 40 18440
rect 0 18405 5 18435
rect 35 18405 40 18435
rect 0 18400 40 18405
rect 80 18435 120 18440
rect 80 18405 85 18435
rect 115 18405 120 18435
rect 80 18400 120 18405
rect 160 18435 200 18440
rect 160 18405 165 18435
rect 195 18405 200 18435
rect 160 18400 200 18405
rect 240 18435 280 18440
rect 240 18405 245 18435
rect 275 18405 280 18435
rect 240 18400 280 18405
rect 320 18435 360 18440
rect 320 18405 325 18435
rect 355 18405 360 18435
rect 320 18400 360 18405
rect 400 18435 440 18440
rect 400 18405 405 18435
rect 435 18405 440 18435
rect 400 18400 440 18405
rect 480 18435 520 18440
rect 480 18405 485 18435
rect 515 18405 520 18435
rect 480 18400 520 18405
rect 560 18435 600 18440
rect 560 18405 565 18435
rect 595 18405 600 18435
rect 560 18400 600 18405
rect 640 18435 680 18440
rect 640 18405 645 18435
rect 675 18405 680 18435
rect 640 18400 680 18405
rect 720 18435 760 18440
rect 720 18405 725 18435
rect 755 18405 760 18435
rect 720 18400 760 18405
rect 800 18435 840 18440
rect 800 18405 805 18435
rect 835 18405 840 18435
rect 800 18400 840 18405
rect 880 18435 920 18440
rect 880 18405 885 18435
rect 915 18405 920 18435
rect 880 18400 920 18405
rect 960 18435 1000 18440
rect 960 18405 965 18435
rect 995 18405 1000 18435
rect 960 18400 1000 18405
rect 1040 18435 1080 18440
rect 1040 18405 1045 18435
rect 1075 18405 1080 18435
rect 1040 18400 1080 18405
rect 1120 18435 1160 18440
rect 1120 18405 1125 18435
rect 1155 18405 1160 18435
rect 1120 18400 1160 18405
rect 1200 18435 1240 18440
rect 1200 18405 1205 18435
rect 1235 18405 1240 18435
rect 1200 18400 1240 18405
rect 1280 18435 1320 18440
rect 1280 18405 1285 18435
rect 1315 18405 1320 18435
rect 1280 18400 1320 18405
rect 1360 18435 1400 18440
rect 1360 18405 1365 18435
rect 1395 18405 1400 18435
rect 1360 18400 1400 18405
rect 1440 18435 1480 18440
rect 1440 18405 1445 18435
rect 1475 18405 1480 18435
rect 1440 18400 1480 18405
rect 1520 18435 1560 18440
rect 1520 18405 1525 18435
rect 1555 18405 1560 18435
rect 1520 18400 1560 18405
rect 1600 18435 1640 18440
rect 1600 18405 1605 18435
rect 1635 18405 1640 18435
rect 1600 18400 1640 18405
rect 1680 18435 1720 18440
rect 1680 18405 1685 18435
rect 1715 18405 1720 18435
rect 1680 18400 1720 18405
rect 1760 18435 1800 18440
rect 1760 18405 1765 18435
rect 1795 18405 1800 18435
rect 1760 18400 1800 18405
rect 1840 18435 1880 18440
rect 1840 18405 1845 18435
rect 1875 18405 1880 18435
rect 1840 18400 1880 18405
rect 1920 18435 1960 18440
rect 1920 18405 1925 18435
rect 1955 18405 1960 18435
rect 1920 18400 1960 18405
rect 2000 18435 2040 18440
rect 2000 18405 2005 18435
rect 2035 18405 2040 18435
rect 2000 18400 2040 18405
rect 2080 18435 2120 18440
rect 2080 18405 2085 18435
rect 2115 18405 2120 18435
rect 2080 18400 2120 18405
rect 2160 18435 2200 18440
rect 2160 18405 2165 18435
rect 2195 18405 2200 18435
rect 2160 18400 2200 18405
rect 2240 18435 2280 18440
rect 2240 18405 2245 18435
rect 2275 18405 2280 18435
rect 2240 18400 2280 18405
rect 2320 18435 2360 18440
rect 2320 18405 2325 18435
rect 2355 18405 2360 18435
rect 2320 18400 2360 18405
rect 2400 18435 2440 18440
rect 2400 18405 2405 18435
rect 2435 18405 2440 18435
rect 2400 18400 2440 18405
rect 2480 18435 2520 18440
rect 2480 18405 2485 18435
rect 2515 18405 2520 18435
rect 2480 18400 2520 18405
rect 2560 18435 2600 18440
rect 2560 18405 2565 18435
rect 2595 18405 2600 18435
rect 2560 18400 2600 18405
rect 2640 18435 2680 18440
rect 2640 18405 2645 18435
rect 2675 18405 2680 18435
rect 2640 18400 2680 18405
rect 2720 18435 2760 18440
rect 2720 18405 2725 18435
rect 2755 18405 2760 18435
rect 2720 18400 2760 18405
rect 2800 18435 2840 18440
rect 2800 18405 2805 18435
rect 2835 18405 2840 18435
rect 2800 18400 2840 18405
rect 2880 18435 2920 18440
rect 2880 18405 2885 18435
rect 2915 18405 2920 18435
rect 2880 18400 2920 18405
rect 2960 18435 3000 18440
rect 2960 18405 2965 18435
rect 2995 18405 3000 18435
rect 2960 18400 3000 18405
rect 3040 18435 3080 18440
rect 3040 18405 3045 18435
rect 3075 18405 3080 18435
rect 3040 18400 3080 18405
rect 3120 18435 3160 18440
rect 3120 18405 3125 18435
rect 3155 18405 3160 18435
rect 3120 18400 3160 18405
rect 3200 18435 3240 18440
rect 3200 18405 3205 18435
rect 3235 18405 3240 18435
rect 3200 18400 3240 18405
rect 3280 18435 3320 18440
rect 3280 18405 3285 18435
rect 3315 18405 3320 18435
rect 3280 18400 3320 18405
rect 3360 18435 3400 18440
rect 3360 18405 3365 18435
rect 3395 18405 3400 18435
rect 3360 18400 3400 18405
rect 3440 18435 3480 18440
rect 3440 18405 3445 18435
rect 3475 18405 3480 18435
rect 3440 18400 3480 18405
rect 3520 18435 3560 18440
rect 3520 18405 3525 18435
rect 3555 18405 3560 18435
rect 3520 18400 3560 18405
rect 3600 18435 3640 18440
rect 3600 18405 3605 18435
rect 3635 18405 3640 18435
rect 3600 18400 3640 18405
rect 3680 18435 3720 18440
rect 3680 18405 3685 18435
rect 3715 18405 3720 18435
rect 3680 18400 3720 18405
rect 3760 18435 3800 18440
rect 3760 18405 3765 18435
rect 3795 18405 3800 18435
rect 3760 18400 3800 18405
rect 3840 18435 3880 18440
rect 3840 18405 3845 18435
rect 3875 18405 3880 18435
rect 3840 18400 3880 18405
rect 3920 18435 3960 18440
rect 3920 18405 3925 18435
rect 3955 18405 3960 18435
rect 3920 18400 3960 18405
rect 4000 18435 4040 18440
rect 4000 18405 4005 18435
rect 4035 18405 4040 18435
rect 4000 18400 4040 18405
rect 4080 18435 4120 18440
rect 4080 18405 4085 18435
rect 4115 18405 4120 18435
rect 4080 18400 4120 18405
rect 4160 18435 4200 18440
rect 4160 18405 4165 18435
rect 4195 18405 4200 18435
rect 4160 18400 4200 18405
rect 6240 18435 6280 18440
rect 6240 18405 6245 18435
rect 6275 18405 6280 18435
rect 6240 18400 6280 18405
rect 6320 18435 6360 18440
rect 6320 18405 6325 18435
rect 6355 18405 6360 18435
rect 6320 18400 6360 18405
rect 6400 18435 6440 18440
rect 6400 18405 6405 18435
rect 6435 18405 6440 18435
rect 6400 18400 6440 18405
rect 6480 18435 6520 18440
rect 6480 18405 6485 18435
rect 6515 18405 6520 18435
rect 6480 18400 6520 18405
rect 6560 18435 6600 18440
rect 6560 18405 6565 18435
rect 6595 18405 6600 18435
rect 6560 18400 6600 18405
rect 6640 18435 6680 18440
rect 6640 18405 6645 18435
rect 6675 18405 6680 18435
rect 6640 18400 6680 18405
rect 6720 18435 6760 18440
rect 6720 18405 6725 18435
rect 6755 18405 6760 18435
rect 6720 18400 6760 18405
rect 6800 18435 6840 18440
rect 6800 18405 6805 18435
rect 6835 18405 6840 18435
rect 6800 18400 6840 18405
rect 6880 18435 6920 18440
rect 6880 18405 6885 18435
rect 6915 18405 6920 18435
rect 6880 18400 6920 18405
rect 6960 18435 7000 18440
rect 6960 18405 6965 18435
rect 6995 18405 7000 18435
rect 6960 18400 7000 18405
rect 7040 18435 7080 18440
rect 7040 18405 7045 18435
rect 7075 18405 7080 18435
rect 7040 18400 7080 18405
rect 7120 18435 7160 18440
rect 7120 18405 7125 18435
rect 7155 18405 7160 18435
rect 7120 18400 7160 18405
rect 7200 18435 7240 18440
rect 7200 18405 7205 18435
rect 7235 18405 7240 18435
rect 7200 18400 7240 18405
rect 7280 18435 7320 18440
rect 7280 18405 7285 18435
rect 7315 18405 7320 18435
rect 7280 18400 7320 18405
rect 7360 18435 7400 18440
rect 7360 18405 7365 18435
rect 7395 18405 7400 18435
rect 7360 18400 7400 18405
rect 7440 18435 7480 18440
rect 7440 18405 7445 18435
rect 7475 18405 7480 18435
rect 7440 18400 7480 18405
rect 7520 18435 7560 18440
rect 7520 18405 7525 18435
rect 7555 18405 7560 18435
rect 7520 18400 7560 18405
rect 7600 18435 7640 18440
rect 7600 18405 7605 18435
rect 7635 18405 7640 18435
rect 7600 18400 7640 18405
rect 7680 18435 7720 18440
rect 7680 18405 7685 18435
rect 7715 18405 7720 18435
rect 7680 18400 7720 18405
rect 7760 18435 7800 18440
rect 7760 18405 7765 18435
rect 7795 18405 7800 18435
rect 7760 18400 7800 18405
rect 7840 18435 7880 18440
rect 7840 18405 7845 18435
rect 7875 18405 7880 18435
rect 7840 18400 7880 18405
rect 7920 18435 7960 18440
rect 7920 18405 7925 18435
rect 7955 18405 7960 18435
rect 7920 18400 7960 18405
rect 8000 18435 8040 18440
rect 8000 18405 8005 18435
rect 8035 18405 8040 18435
rect 8000 18400 8040 18405
rect 8080 18435 8120 18440
rect 8080 18405 8085 18435
rect 8115 18405 8120 18435
rect 8080 18400 8120 18405
rect 8160 18435 8200 18440
rect 8160 18405 8165 18435
rect 8195 18405 8200 18435
rect 8160 18400 8200 18405
rect 8240 18435 8280 18440
rect 8240 18405 8245 18435
rect 8275 18405 8280 18435
rect 8240 18400 8280 18405
rect 8320 18435 8360 18440
rect 8320 18405 8325 18435
rect 8355 18405 8360 18435
rect 8320 18400 8360 18405
rect 8400 18435 8440 18440
rect 8400 18405 8405 18435
rect 8435 18405 8440 18435
rect 8400 18400 8440 18405
rect 8480 18435 8520 18440
rect 8480 18405 8485 18435
rect 8515 18405 8520 18435
rect 8480 18400 8520 18405
rect 8560 18435 8600 18440
rect 8560 18405 8565 18435
rect 8595 18405 8600 18435
rect 8560 18400 8600 18405
rect 8640 18435 8680 18440
rect 8640 18405 8645 18435
rect 8675 18405 8680 18435
rect 8640 18400 8680 18405
rect 8720 18435 8760 18440
rect 8720 18405 8725 18435
rect 8755 18405 8760 18435
rect 8720 18400 8760 18405
rect 8800 18435 8840 18440
rect 8800 18405 8805 18435
rect 8835 18405 8840 18435
rect 8800 18400 8840 18405
rect 8880 18435 8920 18440
rect 8880 18405 8885 18435
rect 8915 18405 8920 18435
rect 8880 18400 8920 18405
rect 8960 18435 9000 18440
rect 8960 18405 8965 18435
rect 8995 18405 9000 18435
rect 8960 18400 9000 18405
rect 9040 18435 9080 18440
rect 9040 18405 9045 18435
rect 9075 18405 9080 18435
rect 9040 18400 9080 18405
rect 9120 18435 9160 18440
rect 9120 18405 9125 18435
rect 9155 18405 9160 18435
rect 9120 18400 9160 18405
rect 9200 18435 9240 18440
rect 9200 18405 9205 18435
rect 9235 18405 9240 18435
rect 9200 18400 9240 18405
rect 9280 18435 9320 18440
rect 9280 18405 9285 18435
rect 9315 18405 9320 18435
rect 9280 18400 9320 18405
rect 9360 18435 9400 18440
rect 9360 18405 9365 18435
rect 9395 18405 9400 18435
rect 9360 18400 9400 18405
rect 9440 18435 9480 18440
rect 9440 18405 9445 18435
rect 9475 18405 9480 18435
rect 9440 18400 9480 18405
rect 11560 18435 11600 18440
rect 11560 18405 11565 18435
rect 11595 18405 11600 18435
rect 11560 18400 11600 18405
rect 11640 18435 11680 18440
rect 11640 18405 11645 18435
rect 11675 18405 11680 18435
rect 11640 18400 11680 18405
rect 11720 18435 11760 18440
rect 11720 18405 11725 18435
rect 11755 18405 11760 18435
rect 11720 18400 11760 18405
rect 11800 18435 11840 18440
rect 11800 18405 11805 18435
rect 11835 18405 11840 18435
rect 11800 18400 11840 18405
rect 11880 18435 11920 18440
rect 11880 18405 11885 18435
rect 11915 18405 11920 18435
rect 11880 18400 11920 18405
rect 11960 18435 12000 18440
rect 11960 18405 11965 18435
rect 11995 18405 12000 18435
rect 11960 18400 12000 18405
rect 12040 18435 12080 18440
rect 12040 18405 12045 18435
rect 12075 18405 12080 18435
rect 12040 18400 12080 18405
rect 12120 18435 12160 18440
rect 12120 18405 12125 18435
rect 12155 18405 12160 18435
rect 12120 18400 12160 18405
rect 12200 18435 12240 18440
rect 12200 18405 12205 18435
rect 12235 18405 12240 18435
rect 12200 18400 12240 18405
rect 12280 18435 12320 18440
rect 12280 18405 12285 18435
rect 12315 18405 12320 18435
rect 12280 18400 12320 18405
rect 12360 18435 12400 18440
rect 12360 18405 12365 18435
rect 12395 18405 12400 18435
rect 12360 18400 12400 18405
rect 12440 18435 12480 18440
rect 12440 18405 12445 18435
rect 12475 18405 12480 18435
rect 12440 18400 12480 18405
rect 12520 18435 12560 18440
rect 12520 18405 12525 18435
rect 12555 18405 12560 18435
rect 12520 18400 12560 18405
rect 12600 18435 12640 18440
rect 12600 18405 12605 18435
rect 12635 18405 12640 18435
rect 12600 18400 12640 18405
rect 12680 18435 12720 18440
rect 12680 18405 12685 18435
rect 12715 18405 12720 18435
rect 12680 18400 12720 18405
rect 12760 18435 12800 18440
rect 12760 18405 12765 18435
rect 12795 18405 12800 18435
rect 12760 18400 12800 18405
rect 12840 18435 12880 18440
rect 12840 18405 12845 18435
rect 12875 18405 12880 18435
rect 12840 18400 12880 18405
rect 12920 18435 12960 18440
rect 12920 18405 12925 18435
rect 12955 18405 12960 18435
rect 12920 18400 12960 18405
rect 13000 18435 13040 18440
rect 13000 18405 13005 18435
rect 13035 18405 13040 18435
rect 13000 18400 13040 18405
rect 13080 18435 13120 18440
rect 13080 18405 13085 18435
rect 13115 18405 13120 18435
rect 13080 18400 13120 18405
rect 13160 18435 13200 18440
rect 13160 18405 13165 18435
rect 13195 18405 13200 18435
rect 13160 18400 13200 18405
rect 13240 18435 13280 18440
rect 13240 18405 13245 18435
rect 13275 18405 13280 18435
rect 13240 18400 13280 18405
rect 13320 18435 13360 18440
rect 13320 18405 13325 18435
rect 13355 18405 13360 18435
rect 13320 18400 13360 18405
rect 13400 18435 13440 18440
rect 13400 18405 13405 18435
rect 13435 18405 13440 18435
rect 13400 18400 13440 18405
rect 13480 18435 13520 18440
rect 13480 18405 13485 18435
rect 13515 18405 13520 18435
rect 13480 18400 13520 18405
rect 13560 18435 13600 18440
rect 13560 18405 13565 18435
rect 13595 18405 13600 18435
rect 13560 18400 13600 18405
rect 13640 18435 13680 18440
rect 13640 18405 13645 18435
rect 13675 18405 13680 18435
rect 13640 18400 13680 18405
rect 13720 18435 13760 18440
rect 13720 18405 13725 18435
rect 13755 18405 13760 18435
rect 13720 18400 13760 18405
rect 13800 18435 13840 18440
rect 13800 18405 13805 18435
rect 13835 18405 13840 18435
rect 13800 18400 13840 18405
rect 13880 18435 13920 18440
rect 13880 18405 13885 18435
rect 13915 18405 13920 18435
rect 13880 18400 13920 18405
rect 13960 18435 14000 18440
rect 13960 18405 13965 18435
rect 13995 18405 14000 18435
rect 13960 18400 14000 18405
rect 14040 18435 14080 18440
rect 14040 18405 14045 18435
rect 14075 18405 14080 18435
rect 14040 18400 14080 18405
rect 14120 18435 14160 18440
rect 14120 18405 14125 18435
rect 14155 18405 14160 18435
rect 14120 18400 14160 18405
rect 14200 18435 14240 18440
rect 14200 18405 14205 18435
rect 14235 18405 14240 18435
rect 14200 18400 14240 18405
rect 14280 18435 14320 18440
rect 14280 18405 14285 18435
rect 14315 18405 14320 18435
rect 14280 18400 14320 18405
rect 14360 18435 14400 18440
rect 14360 18405 14365 18435
rect 14395 18405 14400 18435
rect 14360 18400 14400 18405
rect 14440 18435 14480 18440
rect 14440 18405 14445 18435
rect 14475 18405 14480 18435
rect 14440 18400 14480 18405
rect 14520 18435 14560 18440
rect 14520 18405 14525 18435
rect 14555 18405 14560 18435
rect 14520 18400 14560 18405
rect 14600 18435 14640 18440
rect 14600 18405 14605 18435
rect 14635 18405 14640 18435
rect 14600 18400 14640 18405
rect 14680 18435 14720 18440
rect 14680 18405 14685 18435
rect 14715 18405 14720 18435
rect 14680 18400 14720 18405
rect 16760 18435 16800 18440
rect 16760 18405 16765 18435
rect 16795 18405 16800 18435
rect 16760 18400 16800 18405
rect 16840 18435 16880 18440
rect 16840 18405 16845 18435
rect 16875 18405 16880 18435
rect 16840 18400 16880 18405
rect 16920 18435 16960 18440
rect 16920 18405 16925 18435
rect 16955 18405 16960 18435
rect 16920 18400 16960 18405
rect 17000 18435 17040 18440
rect 17000 18405 17005 18435
rect 17035 18405 17040 18435
rect 17000 18400 17040 18405
rect 17080 18435 17120 18440
rect 17080 18405 17085 18435
rect 17115 18405 17120 18435
rect 17080 18400 17120 18405
rect 17160 18435 17200 18440
rect 17160 18405 17165 18435
rect 17195 18405 17200 18435
rect 17160 18400 17200 18405
rect 17240 18435 17280 18440
rect 17240 18405 17245 18435
rect 17275 18405 17280 18435
rect 17240 18400 17280 18405
rect 17320 18435 17360 18440
rect 17320 18405 17325 18435
rect 17355 18405 17360 18435
rect 17320 18400 17360 18405
rect 17400 18435 17440 18440
rect 17400 18405 17405 18435
rect 17435 18405 17440 18435
rect 17400 18400 17440 18405
rect 17480 18435 17520 18440
rect 17480 18405 17485 18435
rect 17515 18405 17520 18435
rect 17480 18400 17520 18405
rect 17560 18435 17600 18440
rect 17560 18405 17565 18435
rect 17595 18405 17600 18435
rect 17560 18400 17600 18405
rect 17640 18435 17680 18440
rect 17640 18405 17645 18435
rect 17675 18405 17680 18435
rect 17640 18400 17680 18405
rect 17720 18435 17760 18440
rect 17720 18405 17725 18435
rect 17755 18405 17760 18435
rect 17720 18400 17760 18405
rect 17800 18435 17840 18440
rect 17800 18405 17805 18435
rect 17835 18405 17840 18435
rect 17800 18400 17840 18405
rect 17880 18435 17920 18440
rect 17880 18405 17885 18435
rect 17915 18405 17920 18435
rect 17880 18400 17920 18405
rect 17960 18435 18000 18440
rect 17960 18405 17965 18435
rect 17995 18405 18000 18435
rect 17960 18400 18000 18405
rect 18040 18435 18080 18440
rect 18040 18405 18045 18435
rect 18075 18405 18080 18435
rect 18040 18400 18080 18405
rect 18120 18435 18160 18440
rect 18120 18405 18125 18435
rect 18155 18405 18160 18435
rect 18120 18400 18160 18405
rect 18200 18435 18240 18440
rect 18200 18405 18205 18435
rect 18235 18405 18240 18435
rect 18200 18400 18240 18405
rect 18280 18435 18320 18440
rect 18280 18405 18285 18435
rect 18315 18405 18320 18435
rect 18280 18400 18320 18405
rect 18360 18435 18400 18440
rect 18360 18405 18365 18435
rect 18395 18405 18400 18435
rect 18360 18400 18400 18405
rect 18440 18435 18480 18440
rect 18440 18405 18445 18435
rect 18475 18405 18480 18435
rect 18440 18400 18480 18405
rect 18520 18435 18560 18440
rect 18520 18405 18525 18435
rect 18555 18405 18560 18435
rect 18520 18400 18560 18405
rect 18600 18435 18640 18440
rect 18600 18405 18605 18435
rect 18635 18405 18640 18435
rect 18600 18400 18640 18405
rect 18680 18435 18720 18440
rect 18680 18405 18685 18435
rect 18715 18405 18720 18435
rect 18680 18400 18720 18405
rect 18760 18435 18800 18440
rect 18760 18405 18765 18435
rect 18795 18405 18800 18435
rect 18760 18400 18800 18405
rect 18840 18435 18880 18440
rect 18840 18405 18845 18435
rect 18875 18405 18880 18435
rect 18840 18400 18880 18405
rect 18920 18435 18960 18440
rect 18920 18405 18925 18435
rect 18955 18405 18960 18435
rect 18920 18400 18960 18405
rect 19000 18435 19040 18440
rect 19000 18405 19005 18435
rect 19035 18405 19040 18435
rect 19000 18400 19040 18405
rect 19080 18435 19120 18440
rect 19080 18405 19085 18435
rect 19115 18405 19120 18435
rect 19080 18400 19120 18405
rect 19160 18435 19200 18440
rect 19160 18405 19165 18435
rect 19195 18405 19200 18435
rect 19160 18400 19200 18405
rect 19240 18435 19280 18440
rect 19240 18405 19245 18435
rect 19275 18405 19280 18435
rect 19240 18400 19280 18405
rect 19320 18435 19360 18440
rect 19320 18405 19325 18435
rect 19355 18405 19360 18435
rect 19320 18400 19360 18405
rect 19400 18435 19440 18440
rect 19400 18405 19405 18435
rect 19435 18405 19440 18435
rect 19400 18400 19440 18405
rect 19480 18435 19520 18440
rect 19480 18405 19485 18435
rect 19515 18405 19520 18435
rect 19480 18400 19520 18405
rect 19560 18435 19600 18440
rect 19560 18405 19565 18435
rect 19595 18405 19600 18435
rect 19560 18400 19600 18405
rect 19640 18435 19680 18440
rect 19640 18405 19645 18435
rect 19675 18405 19680 18435
rect 19640 18400 19680 18405
rect 19720 18435 19760 18440
rect 19720 18405 19725 18435
rect 19755 18405 19760 18435
rect 19720 18400 19760 18405
rect 19800 18435 19840 18440
rect 19800 18405 19805 18435
rect 19835 18405 19840 18435
rect 19800 18400 19840 18405
rect 19880 18435 19920 18440
rect 19880 18405 19885 18435
rect 19915 18405 19920 18435
rect 19880 18400 19920 18405
rect 19960 18435 20000 18440
rect 19960 18405 19965 18435
rect 19995 18405 20000 18435
rect 19960 18400 20000 18405
rect 20040 18435 20080 18440
rect 20040 18405 20045 18435
rect 20075 18405 20080 18435
rect 20040 18400 20080 18405
rect 20120 18435 20160 18440
rect 20120 18405 20125 18435
rect 20155 18405 20160 18435
rect 20120 18400 20160 18405
rect 20200 18435 20240 18440
rect 20200 18405 20205 18435
rect 20235 18405 20240 18435
rect 20200 18400 20240 18405
rect 20280 18435 20320 18440
rect 20280 18405 20285 18435
rect 20315 18405 20320 18435
rect 20280 18400 20320 18405
rect 20360 18435 20400 18440
rect 20360 18405 20365 18435
rect 20395 18405 20400 18435
rect 20360 18400 20400 18405
rect 20440 18435 20480 18440
rect 20440 18405 20445 18435
rect 20475 18405 20480 18435
rect 20440 18400 20480 18405
rect 20520 18435 20560 18440
rect 20520 18405 20525 18435
rect 20555 18405 20560 18435
rect 20520 18400 20560 18405
rect 20600 18435 20640 18440
rect 20600 18405 20605 18435
rect 20635 18405 20640 18435
rect 20600 18400 20640 18405
rect 20680 18435 20720 18440
rect 20680 18405 20685 18435
rect 20715 18405 20720 18435
rect 20680 18400 20720 18405
rect 20760 18435 20800 18440
rect 20760 18405 20765 18435
rect 20795 18405 20800 18435
rect 20760 18400 20800 18405
rect 20840 18435 20880 18440
rect 20840 18405 20845 18435
rect 20875 18405 20880 18435
rect 20840 18400 20880 18405
rect 20920 18435 20960 18440
rect 20920 18405 20925 18435
rect 20955 18405 20960 18435
rect 20920 18400 20960 18405
rect 0 18275 40 18280
rect 0 18245 5 18275
rect 35 18245 40 18275
rect 0 18240 40 18245
rect 80 18275 120 18280
rect 80 18245 85 18275
rect 115 18245 120 18275
rect 80 18240 120 18245
rect 160 18275 200 18280
rect 160 18245 165 18275
rect 195 18245 200 18275
rect 160 18240 200 18245
rect 240 18275 280 18280
rect 240 18245 245 18275
rect 275 18245 280 18275
rect 240 18240 280 18245
rect 320 18275 360 18280
rect 320 18245 325 18275
rect 355 18245 360 18275
rect 320 18240 360 18245
rect 400 18275 440 18280
rect 400 18245 405 18275
rect 435 18245 440 18275
rect 400 18240 440 18245
rect 480 18275 520 18280
rect 480 18245 485 18275
rect 515 18245 520 18275
rect 480 18240 520 18245
rect 560 18275 600 18280
rect 560 18245 565 18275
rect 595 18245 600 18275
rect 560 18240 600 18245
rect 640 18275 680 18280
rect 640 18245 645 18275
rect 675 18245 680 18275
rect 640 18240 680 18245
rect 720 18275 760 18280
rect 720 18245 725 18275
rect 755 18245 760 18275
rect 720 18240 760 18245
rect 800 18275 840 18280
rect 800 18245 805 18275
rect 835 18245 840 18275
rect 800 18240 840 18245
rect 880 18275 920 18280
rect 880 18245 885 18275
rect 915 18245 920 18275
rect 880 18240 920 18245
rect 960 18275 1000 18280
rect 960 18245 965 18275
rect 995 18245 1000 18275
rect 960 18240 1000 18245
rect 1040 18275 1080 18280
rect 1040 18245 1045 18275
rect 1075 18245 1080 18275
rect 1040 18240 1080 18245
rect 1120 18275 1160 18280
rect 1120 18245 1125 18275
rect 1155 18245 1160 18275
rect 1120 18240 1160 18245
rect 1200 18275 1240 18280
rect 1200 18245 1205 18275
rect 1235 18245 1240 18275
rect 1200 18240 1240 18245
rect 1280 18275 1320 18280
rect 1280 18245 1285 18275
rect 1315 18245 1320 18275
rect 1280 18240 1320 18245
rect 1360 18275 1400 18280
rect 1360 18245 1365 18275
rect 1395 18245 1400 18275
rect 1360 18240 1400 18245
rect 1440 18275 1480 18280
rect 1440 18245 1445 18275
rect 1475 18245 1480 18275
rect 1440 18240 1480 18245
rect 1520 18275 1560 18280
rect 1520 18245 1525 18275
rect 1555 18245 1560 18275
rect 1520 18240 1560 18245
rect 1600 18275 1640 18280
rect 1600 18245 1605 18275
rect 1635 18245 1640 18275
rect 1600 18240 1640 18245
rect 1680 18275 1720 18280
rect 1680 18245 1685 18275
rect 1715 18245 1720 18275
rect 1680 18240 1720 18245
rect 1760 18275 1800 18280
rect 1760 18245 1765 18275
rect 1795 18245 1800 18275
rect 1760 18240 1800 18245
rect 1840 18275 1880 18280
rect 1840 18245 1845 18275
rect 1875 18245 1880 18275
rect 1840 18240 1880 18245
rect 1920 18275 1960 18280
rect 1920 18245 1925 18275
rect 1955 18245 1960 18275
rect 1920 18240 1960 18245
rect 2000 18275 2040 18280
rect 2000 18245 2005 18275
rect 2035 18245 2040 18275
rect 2000 18240 2040 18245
rect 2080 18275 2120 18280
rect 2080 18245 2085 18275
rect 2115 18245 2120 18275
rect 2080 18240 2120 18245
rect 2160 18275 2200 18280
rect 2160 18245 2165 18275
rect 2195 18245 2200 18275
rect 2160 18240 2200 18245
rect 2240 18275 2280 18280
rect 2240 18245 2245 18275
rect 2275 18245 2280 18275
rect 2240 18240 2280 18245
rect 2320 18275 2360 18280
rect 2320 18245 2325 18275
rect 2355 18245 2360 18275
rect 2320 18240 2360 18245
rect 2400 18275 2440 18280
rect 2400 18245 2405 18275
rect 2435 18245 2440 18275
rect 2400 18240 2440 18245
rect 2480 18275 2520 18280
rect 2480 18245 2485 18275
rect 2515 18245 2520 18275
rect 2480 18240 2520 18245
rect 2560 18275 2600 18280
rect 2560 18245 2565 18275
rect 2595 18245 2600 18275
rect 2560 18240 2600 18245
rect 2640 18275 2680 18280
rect 2640 18245 2645 18275
rect 2675 18245 2680 18275
rect 2640 18240 2680 18245
rect 2720 18275 2760 18280
rect 2720 18245 2725 18275
rect 2755 18245 2760 18275
rect 2720 18240 2760 18245
rect 2800 18275 2840 18280
rect 2800 18245 2805 18275
rect 2835 18245 2840 18275
rect 2800 18240 2840 18245
rect 2880 18275 2920 18280
rect 2880 18245 2885 18275
rect 2915 18245 2920 18275
rect 2880 18240 2920 18245
rect 2960 18275 3000 18280
rect 2960 18245 2965 18275
rect 2995 18245 3000 18275
rect 2960 18240 3000 18245
rect 3040 18275 3080 18280
rect 3040 18245 3045 18275
rect 3075 18245 3080 18275
rect 3040 18240 3080 18245
rect 3120 18275 3160 18280
rect 3120 18245 3125 18275
rect 3155 18245 3160 18275
rect 3120 18240 3160 18245
rect 3200 18275 3240 18280
rect 3200 18245 3205 18275
rect 3235 18245 3240 18275
rect 3200 18240 3240 18245
rect 3280 18275 3320 18280
rect 3280 18245 3285 18275
rect 3315 18245 3320 18275
rect 3280 18240 3320 18245
rect 3360 18275 3400 18280
rect 3360 18245 3365 18275
rect 3395 18245 3400 18275
rect 3360 18240 3400 18245
rect 3440 18275 3480 18280
rect 3440 18245 3445 18275
rect 3475 18245 3480 18275
rect 3440 18240 3480 18245
rect 3520 18275 3560 18280
rect 3520 18245 3525 18275
rect 3555 18245 3560 18275
rect 3520 18240 3560 18245
rect 3600 18275 3640 18280
rect 3600 18245 3605 18275
rect 3635 18245 3640 18275
rect 3600 18240 3640 18245
rect 3680 18275 3720 18280
rect 3680 18245 3685 18275
rect 3715 18245 3720 18275
rect 3680 18240 3720 18245
rect 3760 18275 3800 18280
rect 3760 18245 3765 18275
rect 3795 18245 3800 18275
rect 3760 18240 3800 18245
rect 3840 18275 3880 18280
rect 3840 18245 3845 18275
rect 3875 18245 3880 18275
rect 3840 18240 3880 18245
rect 3920 18275 3960 18280
rect 3920 18245 3925 18275
rect 3955 18245 3960 18275
rect 3920 18240 3960 18245
rect 4000 18275 4040 18280
rect 4000 18245 4005 18275
rect 4035 18245 4040 18275
rect 4000 18240 4040 18245
rect 4080 18275 4120 18280
rect 4080 18245 4085 18275
rect 4115 18245 4120 18275
rect 4080 18240 4120 18245
rect 4160 18275 4200 18280
rect 4160 18245 4165 18275
rect 4195 18245 4200 18275
rect 4160 18240 4200 18245
rect 6240 18275 6280 18280
rect 6240 18245 6245 18275
rect 6275 18245 6280 18275
rect 6240 18240 6280 18245
rect 6320 18275 6360 18280
rect 6320 18245 6325 18275
rect 6355 18245 6360 18275
rect 6320 18240 6360 18245
rect 6400 18275 6440 18280
rect 6400 18245 6405 18275
rect 6435 18245 6440 18275
rect 6400 18240 6440 18245
rect 6480 18275 6520 18280
rect 6480 18245 6485 18275
rect 6515 18245 6520 18275
rect 6480 18240 6520 18245
rect 6560 18275 6600 18280
rect 6560 18245 6565 18275
rect 6595 18245 6600 18275
rect 6560 18240 6600 18245
rect 6640 18275 6680 18280
rect 6640 18245 6645 18275
rect 6675 18245 6680 18275
rect 6640 18240 6680 18245
rect 6720 18275 6760 18280
rect 6720 18245 6725 18275
rect 6755 18245 6760 18275
rect 6720 18240 6760 18245
rect 6800 18275 6840 18280
rect 6800 18245 6805 18275
rect 6835 18245 6840 18275
rect 6800 18240 6840 18245
rect 6880 18275 6920 18280
rect 6880 18245 6885 18275
rect 6915 18245 6920 18275
rect 6880 18240 6920 18245
rect 6960 18275 7000 18280
rect 6960 18245 6965 18275
rect 6995 18245 7000 18275
rect 6960 18240 7000 18245
rect 7040 18275 7080 18280
rect 7040 18245 7045 18275
rect 7075 18245 7080 18275
rect 7040 18240 7080 18245
rect 7120 18275 7160 18280
rect 7120 18245 7125 18275
rect 7155 18245 7160 18275
rect 7120 18240 7160 18245
rect 7200 18275 7240 18280
rect 7200 18245 7205 18275
rect 7235 18245 7240 18275
rect 7200 18240 7240 18245
rect 7280 18275 7320 18280
rect 7280 18245 7285 18275
rect 7315 18245 7320 18275
rect 7280 18240 7320 18245
rect 7360 18275 7400 18280
rect 7360 18245 7365 18275
rect 7395 18245 7400 18275
rect 7360 18240 7400 18245
rect 7440 18275 7480 18280
rect 7440 18245 7445 18275
rect 7475 18245 7480 18275
rect 7440 18240 7480 18245
rect 7520 18275 7560 18280
rect 7520 18245 7525 18275
rect 7555 18245 7560 18275
rect 7520 18240 7560 18245
rect 7600 18275 7640 18280
rect 7600 18245 7605 18275
rect 7635 18245 7640 18275
rect 7600 18240 7640 18245
rect 7680 18275 7720 18280
rect 7680 18245 7685 18275
rect 7715 18245 7720 18275
rect 7680 18240 7720 18245
rect 7760 18275 7800 18280
rect 7760 18245 7765 18275
rect 7795 18245 7800 18275
rect 7760 18240 7800 18245
rect 7840 18275 7880 18280
rect 7840 18245 7845 18275
rect 7875 18245 7880 18275
rect 7840 18240 7880 18245
rect 7920 18275 7960 18280
rect 7920 18245 7925 18275
rect 7955 18245 7960 18275
rect 7920 18240 7960 18245
rect 8000 18275 8040 18280
rect 8000 18245 8005 18275
rect 8035 18245 8040 18275
rect 8000 18240 8040 18245
rect 8080 18275 8120 18280
rect 8080 18245 8085 18275
rect 8115 18245 8120 18275
rect 8080 18240 8120 18245
rect 8160 18275 8200 18280
rect 8160 18245 8165 18275
rect 8195 18245 8200 18275
rect 8160 18240 8200 18245
rect 8240 18275 8280 18280
rect 8240 18245 8245 18275
rect 8275 18245 8280 18275
rect 8240 18240 8280 18245
rect 8320 18275 8360 18280
rect 8320 18245 8325 18275
rect 8355 18245 8360 18275
rect 8320 18240 8360 18245
rect 8400 18275 8440 18280
rect 8400 18245 8405 18275
rect 8435 18245 8440 18275
rect 8400 18240 8440 18245
rect 8480 18275 8520 18280
rect 8480 18245 8485 18275
rect 8515 18245 8520 18275
rect 8480 18240 8520 18245
rect 8560 18275 8600 18280
rect 8560 18245 8565 18275
rect 8595 18245 8600 18275
rect 8560 18240 8600 18245
rect 8640 18275 8680 18280
rect 8640 18245 8645 18275
rect 8675 18245 8680 18275
rect 8640 18240 8680 18245
rect 8720 18275 8760 18280
rect 8720 18245 8725 18275
rect 8755 18245 8760 18275
rect 8720 18240 8760 18245
rect 8800 18275 8840 18280
rect 8800 18245 8805 18275
rect 8835 18245 8840 18275
rect 8800 18240 8840 18245
rect 8880 18275 8920 18280
rect 8880 18245 8885 18275
rect 8915 18245 8920 18275
rect 8880 18240 8920 18245
rect 8960 18275 9000 18280
rect 8960 18245 8965 18275
rect 8995 18245 9000 18275
rect 8960 18240 9000 18245
rect 9040 18275 9080 18280
rect 9040 18245 9045 18275
rect 9075 18245 9080 18275
rect 9040 18240 9080 18245
rect 9120 18275 9160 18280
rect 9120 18245 9125 18275
rect 9155 18245 9160 18275
rect 9120 18240 9160 18245
rect 9200 18275 9240 18280
rect 9200 18245 9205 18275
rect 9235 18245 9240 18275
rect 9200 18240 9240 18245
rect 9280 18275 9320 18280
rect 9280 18245 9285 18275
rect 9315 18245 9320 18275
rect 9280 18240 9320 18245
rect 9360 18275 9400 18280
rect 9360 18245 9365 18275
rect 9395 18245 9400 18275
rect 9360 18240 9400 18245
rect 9440 18275 9480 18280
rect 9440 18245 9445 18275
rect 9475 18245 9480 18275
rect 9440 18240 9480 18245
rect 11560 18275 11600 18280
rect 11560 18245 11565 18275
rect 11595 18245 11600 18275
rect 11560 18240 11600 18245
rect 11640 18275 11680 18280
rect 11640 18245 11645 18275
rect 11675 18245 11680 18275
rect 11640 18240 11680 18245
rect 11720 18275 11760 18280
rect 11720 18245 11725 18275
rect 11755 18245 11760 18275
rect 11720 18240 11760 18245
rect 11800 18275 11840 18280
rect 11800 18245 11805 18275
rect 11835 18245 11840 18275
rect 11800 18240 11840 18245
rect 11880 18275 11920 18280
rect 11880 18245 11885 18275
rect 11915 18245 11920 18275
rect 11880 18240 11920 18245
rect 11960 18275 12000 18280
rect 11960 18245 11965 18275
rect 11995 18245 12000 18275
rect 11960 18240 12000 18245
rect 12040 18275 12080 18280
rect 12040 18245 12045 18275
rect 12075 18245 12080 18275
rect 12040 18240 12080 18245
rect 12120 18275 12160 18280
rect 12120 18245 12125 18275
rect 12155 18245 12160 18275
rect 12120 18240 12160 18245
rect 12200 18275 12240 18280
rect 12200 18245 12205 18275
rect 12235 18245 12240 18275
rect 12200 18240 12240 18245
rect 12280 18275 12320 18280
rect 12280 18245 12285 18275
rect 12315 18245 12320 18275
rect 12280 18240 12320 18245
rect 12360 18275 12400 18280
rect 12360 18245 12365 18275
rect 12395 18245 12400 18275
rect 12360 18240 12400 18245
rect 12440 18275 12480 18280
rect 12440 18245 12445 18275
rect 12475 18245 12480 18275
rect 12440 18240 12480 18245
rect 12520 18275 12560 18280
rect 12520 18245 12525 18275
rect 12555 18245 12560 18275
rect 12520 18240 12560 18245
rect 12600 18275 12640 18280
rect 12600 18245 12605 18275
rect 12635 18245 12640 18275
rect 12600 18240 12640 18245
rect 12680 18275 12720 18280
rect 12680 18245 12685 18275
rect 12715 18245 12720 18275
rect 12680 18240 12720 18245
rect 12760 18275 12800 18280
rect 12760 18245 12765 18275
rect 12795 18245 12800 18275
rect 12760 18240 12800 18245
rect 12840 18275 12880 18280
rect 12840 18245 12845 18275
rect 12875 18245 12880 18275
rect 12840 18240 12880 18245
rect 12920 18275 12960 18280
rect 12920 18245 12925 18275
rect 12955 18245 12960 18275
rect 12920 18240 12960 18245
rect 13000 18275 13040 18280
rect 13000 18245 13005 18275
rect 13035 18245 13040 18275
rect 13000 18240 13040 18245
rect 13080 18275 13120 18280
rect 13080 18245 13085 18275
rect 13115 18245 13120 18275
rect 13080 18240 13120 18245
rect 13160 18275 13200 18280
rect 13160 18245 13165 18275
rect 13195 18245 13200 18275
rect 13160 18240 13200 18245
rect 13240 18275 13280 18280
rect 13240 18245 13245 18275
rect 13275 18245 13280 18275
rect 13240 18240 13280 18245
rect 13320 18275 13360 18280
rect 13320 18245 13325 18275
rect 13355 18245 13360 18275
rect 13320 18240 13360 18245
rect 13400 18275 13440 18280
rect 13400 18245 13405 18275
rect 13435 18245 13440 18275
rect 13400 18240 13440 18245
rect 13480 18275 13520 18280
rect 13480 18245 13485 18275
rect 13515 18245 13520 18275
rect 13480 18240 13520 18245
rect 13560 18275 13600 18280
rect 13560 18245 13565 18275
rect 13595 18245 13600 18275
rect 13560 18240 13600 18245
rect 13640 18275 13680 18280
rect 13640 18245 13645 18275
rect 13675 18245 13680 18275
rect 13640 18240 13680 18245
rect 13720 18275 13760 18280
rect 13720 18245 13725 18275
rect 13755 18245 13760 18275
rect 13720 18240 13760 18245
rect 13800 18275 13840 18280
rect 13800 18245 13805 18275
rect 13835 18245 13840 18275
rect 13800 18240 13840 18245
rect 13880 18275 13920 18280
rect 13880 18245 13885 18275
rect 13915 18245 13920 18275
rect 13880 18240 13920 18245
rect 13960 18275 14000 18280
rect 13960 18245 13965 18275
rect 13995 18245 14000 18275
rect 13960 18240 14000 18245
rect 14040 18275 14080 18280
rect 14040 18245 14045 18275
rect 14075 18245 14080 18275
rect 14040 18240 14080 18245
rect 14120 18275 14160 18280
rect 14120 18245 14125 18275
rect 14155 18245 14160 18275
rect 14120 18240 14160 18245
rect 14200 18275 14240 18280
rect 14200 18245 14205 18275
rect 14235 18245 14240 18275
rect 14200 18240 14240 18245
rect 14280 18275 14320 18280
rect 14280 18245 14285 18275
rect 14315 18245 14320 18275
rect 14280 18240 14320 18245
rect 14360 18275 14400 18280
rect 14360 18245 14365 18275
rect 14395 18245 14400 18275
rect 14360 18240 14400 18245
rect 14440 18275 14480 18280
rect 14440 18245 14445 18275
rect 14475 18245 14480 18275
rect 14440 18240 14480 18245
rect 14520 18275 14560 18280
rect 14520 18245 14525 18275
rect 14555 18245 14560 18275
rect 14520 18240 14560 18245
rect 14600 18275 14640 18280
rect 14600 18245 14605 18275
rect 14635 18245 14640 18275
rect 14600 18240 14640 18245
rect 14680 18275 14720 18280
rect 14680 18245 14685 18275
rect 14715 18245 14720 18275
rect 14680 18240 14720 18245
rect 16760 18275 16800 18280
rect 16760 18245 16765 18275
rect 16795 18245 16800 18275
rect 16760 18240 16800 18245
rect 16840 18275 16880 18280
rect 16840 18245 16845 18275
rect 16875 18245 16880 18275
rect 16840 18240 16880 18245
rect 16920 18275 16960 18280
rect 16920 18245 16925 18275
rect 16955 18245 16960 18275
rect 16920 18240 16960 18245
rect 17000 18275 17040 18280
rect 17000 18245 17005 18275
rect 17035 18245 17040 18275
rect 17000 18240 17040 18245
rect 17080 18275 17120 18280
rect 17080 18245 17085 18275
rect 17115 18245 17120 18275
rect 17080 18240 17120 18245
rect 17160 18275 17200 18280
rect 17160 18245 17165 18275
rect 17195 18245 17200 18275
rect 17160 18240 17200 18245
rect 17240 18275 17280 18280
rect 17240 18245 17245 18275
rect 17275 18245 17280 18275
rect 17240 18240 17280 18245
rect 17320 18275 17360 18280
rect 17320 18245 17325 18275
rect 17355 18245 17360 18275
rect 17320 18240 17360 18245
rect 17400 18275 17440 18280
rect 17400 18245 17405 18275
rect 17435 18245 17440 18275
rect 17400 18240 17440 18245
rect 17480 18275 17520 18280
rect 17480 18245 17485 18275
rect 17515 18245 17520 18275
rect 17480 18240 17520 18245
rect 17560 18275 17600 18280
rect 17560 18245 17565 18275
rect 17595 18245 17600 18275
rect 17560 18240 17600 18245
rect 17640 18275 17680 18280
rect 17640 18245 17645 18275
rect 17675 18245 17680 18275
rect 17640 18240 17680 18245
rect 17720 18275 17760 18280
rect 17720 18245 17725 18275
rect 17755 18245 17760 18275
rect 17720 18240 17760 18245
rect 17800 18275 17840 18280
rect 17800 18245 17805 18275
rect 17835 18245 17840 18275
rect 17800 18240 17840 18245
rect 17880 18275 17920 18280
rect 17880 18245 17885 18275
rect 17915 18245 17920 18275
rect 17880 18240 17920 18245
rect 17960 18275 18000 18280
rect 17960 18245 17965 18275
rect 17995 18245 18000 18275
rect 17960 18240 18000 18245
rect 18040 18275 18080 18280
rect 18040 18245 18045 18275
rect 18075 18245 18080 18275
rect 18040 18240 18080 18245
rect 18120 18275 18160 18280
rect 18120 18245 18125 18275
rect 18155 18245 18160 18275
rect 18120 18240 18160 18245
rect 18200 18275 18240 18280
rect 18200 18245 18205 18275
rect 18235 18245 18240 18275
rect 18200 18240 18240 18245
rect 18280 18275 18320 18280
rect 18280 18245 18285 18275
rect 18315 18245 18320 18275
rect 18280 18240 18320 18245
rect 18360 18275 18400 18280
rect 18360 18245 18365 18275
rect 18395 18245 18400 18275
rect 18360 18240 18400 18245
rect 18440 18275 18480 18280
rect 18440 18245 18445 18275
rect 18475 18245 18480 18275
rect 18440 18240 18480 18245
rect 18520 18275 18560 18280
rect 18520 18245 18525 18275
rect 18555 18245 18560 18275
rect 18520 18240 18560 18245
rect 18600 18275 18640 18280
rect 18600 18245 18605 18275
rect 18635 18245 18640 18275
rect 18600 18240 18640 18245
rect 18680 18275 18720 18280
rect 18680 18245 18685 18275
rect 18715 18245 18720 18275
rect 18680 18240 18720 18245
rect 18760 18275 18800 18280
rect 18760 18245 18765 18275
rect 18795 18245 18800 18275
rect 18760 18240 18800 18245
rect 18840 18275 18880 18280
rect 18840 18245 18845 18275
rect 18875 18245 18880 18275
rect 18840 18240 18880 18245
rect 18920 18275 18960 18280
rect 18920 18245 18925 18275
rect 18955 18245 18960 18275
rect 18920 18240 18960 18245
rect 19000 18275 19040 18280
rect 19000 18245 19005 18275
rect 19035 18245 19040 18275
rect 19000 18240 19040 18245
rect 19080 18275 19120 18280
rect 19080 18245 19085 18275
rect 19115 18245 19120 18275
rect 19080 18240 19120 18245
rect 19160 18275 19200 18280
rect 19160 18245 19165 18275
rect 19195 18245 19200 18275
rect 19160 18240 19200 18245
rect 19240 18275 19280 18280
rect 19240 18245 19245 18275
rect 19275 18245 19280 18275
rect 19240 18240 19280 18245
rect 19320 18275 19360 18280
rect 19320 18245 19325 18275
rect 19355 18245 19360 18275
rect 19320 18240 19360 18245
rect 19400 18275 19440 18280
rect 19400 18245 19405 18275
rect 19435 18245 19440 18275
rect 19400 18240 19440 18245
rect 19480 18275 19520 18280
rect 19480 18245 19485 18275
rect 19515 18245 19520 18275
rect 19480 18240 19520 18245
rect 19560 18275 19600 18280
rect 19560 18245 19565 18275
rect 19595 18245 19600 18275
rect 19560 18240 19600 18245
rect 19640 18275 19680 18280
rect 19640 18245 19645 18275
rect 19675 18245 19680 18275
rect 19640 18240 19680 18245
rect 19720 18275 19760 18280
rect 19720 18245 19725 18275
rect 19755 18245 19760 18275
rect 19720 18240 19760 18245
rect 19800 18275 19840 18280
rect 19800 18245 19805 18275
rect 19835 18245 19840 18275
rect 19800 18240 19840 18245
rect 19880 18275 19920 18280
rect 19880 18245 19885 18275
rect 19915 18245 19920 18275
rect 19880 18240 19920 18245
rect 19960 18275 20000 18280
rect 19960 18245 19965 18275
rect 19995 18245 20000 18275
rect 19960 18240 20000 18245
rect 20040 18275 20080 18280
rect 20040 18245 20045 18275
rect 20075 18245 20080 18275
rect 20040 18240 20080 18245
rect 20120 18275 20160 18280
rect 20120 18245 20125 18275
rect 20155 18245 20160 18275
rect 20120 18240 20160 18245
rect 20200 18275 20240 18280
rect 20200 18245 20205 18275
rect 20235 18245 20240 18275
rect 20200 18240 20240 18245
rect 20280 18275 20320 18280
rect 20280 18245 20285 18275
rect 20315 18245 20320 18275
rect 20280 18240 20320 18245
rect 20360 18275 20400 18280
rect 20360 18245 20365 18275
rect 20395 18245 20400 18275
rect 20360 18240 20400 18245
rect 20440 18275 20480 18280
rect 20440 18245 20445 18275
rect 20475 18245 20480 18275
rect 20440 18240 20480 18245
rect 20520 18275 20560 18280
rect 20520 18245 20525 18275
rect 20555 18245 20560 18275
rect 20520 18240 20560 18245
rect 20600 18275 20640 18280
rect 20600 18245 20605 18275
rect 20635 18245 20640 18275
rect 20600 18240 20640 18245
rect 20680 18275 20720 18280
rect 20680 18245 20685 18275
rect 20715 18245 20720 18275
rect 20680 18240 20720 18245
rect 20760 18275 20800 18280
rect 20760 18245 20765 18275
rect 20795 18245 20800 18275
rect 20760 18240 20800 18245
rect 20840 18275 20880 18280
rect 20840 18245 20845 18275
rect 20875 18245 20880 18275
rect 20840 18240 20880 18245
rect 20920 18275 20960 18280
rect 20920 18245 20925 18275
rect 20955 18245 20960 18275
rect 20920 18240 20960 18245
rect 0 18195 40 18200
rect 0 18165 5 18195
rect 35 18165 40 18195
rect 0 18160 40 18165
rect 80 18195 120 18200
rect 80 18165 85 18195
rect 115 18165 120 18195
rect 80 18160 120 18165
rect 160 18195 200 18200
rect 160 18165 165 18195
rect 195 18165 200 18195
rect 160 18160 200 18165
rect 240 18195 280 18200
rect 240 18165 245 18195
rect 275 18165 280 18195
rect 240 18160 280 18165
rect 320 18195 360 18200
rect 320 18165 325 18195
rect 355 18165 360 18195
rect 320 18160 360 18165
rect 400 18195 440 18200
rect 400 18165 405 18195
rect 435 18165 440 18195
rect 400 18160 440 18165
rect 480 18195 520 18200
rect 480 18165 485 18195
rect 515 18165 520 18195
rect 480 18160 520 18165
rect 560 18195 600 18200
rect 560 18165 565 18195
rect 595 18165 600 18195
rect 560 18160 600 18165
rect 640 18195 680 18200
rect 640 18165 645 18195
rect 675 18165 680 18195
rect 640 18160 680 18165
rect 720 18195 760 18200
rect 720 18165 725 18195
rect 755 18165 760 18195
rect 720 18160 760 18165
rect 800 18195 840 18200
rect 800 18165 805 18195
rect 835 18165 840 18195
rect 800 18160 840 18165
rect 880 18195 920 18200
rect 880 18165 885 18195
rect 915 18165 920 18195
rect 880 18160 920 18165
rect 960 18195 1000 18200
rect 960 18165 965 18195
rect 995 18165 1000 18195
rect 960 18160 1000 18165
rect 1040 18195 1080 18200
rect 1040 18165 1045 18195
rect 1075 18165 1080 18195
rect 1040 18160 1080 18165
rect 1120 18195 1160 18200
rect 1120 18165 1125 18195
rect 1155 18165 1160 18195
rect 1120 18160 1160 18165
rect 1200 18195 1240 18200
rect 1200 18165 1205 18195
rect 1235 18165 1240 18195
rect 1200 18160 1240 18165
rect 1280 18195 1320 18200
rect 1280 18165 1285 18195
rect 1315 18165 1320 18195
rect 1280 18160 1320 18165
rect 1360 18195 1400 18200
rect 1360 18165 1365 18195
rect 1395 18165 1400 18195
rect 1360 18160 1400 18165
rect 1440 18195 1480 18200
rect 1440 18165 1445 18195
rect 1475 18165 1480 18195
rect 1440 18160 1480 18165
rect 1520 18195 1560 18200
rect 1520 18165 1525 18195
rect 1555 18165 1560 18195
rect 1520 18160 1560 18165
rect 1600 18195 1640 18200
rect 1600 18165 1605 18195
rect 1635 18165 1640 18195
rect 1600 18160 1640 18165
rect 1680 18195 1720 18200
rect 1680 18165 1685 18195
rect 1715 18165 1720 18195
rect 1680 18160 1720 18165
rect 1760 18195 1800 18200
rect 1760 18165 1765 18195
rect 1795 18165 1800 18195
rect 1760 18160 1800 18165
rect 1840 18195 1880 18200
rect 1840 18165 1845 18195
rect 1875 18165 1880 18195
rect 1840 18160 1880 18165
rect 1920 18195 1960 18200
rect 1920 18165 1925 18195
rect 1955 18165 1960 18195
rect 1920 18160 1960 18165
rect 2000 18195 2040 18200
rect 2000 18165 2005 18195
rect 2035 18165 2040 18195
rect 2000 18160 2040 18165
rect 2080 18195 2120 18200
rect 2080 18165 2085 18195
rect 2115 18165 2120 18195
rect 2080 18160 2120 18165
rect 2160 18195 2200 18200
rect 2160 18165 2165 18195
rect 2195 18165 2200 18195
rect 2160 18160 2200 18165
rect 2240 18195 2280 18200
rect 2240 18165 2245 18195
rect 2275 18165 2280 18195
rect 2240 18160 2280 18165
rect 2320 18195 2360 18200
rect 2320 18165 2325 18195
rect 2355 18165 2360 18195
rect 2320 18160 2360 18165
rect 2400 18195 2440 18200
rect 2400 18165 2405 18195
rect 2435 18165 2440 18195
rect 2400 18160 2440 18165
rect 2480 18195 2520 18200
rect 2480 18165 2485 18195
rect 2515 18165 2520 18195
rect 2480 18160 2520 18165
rect 2560 18195 2600 18200
rect 2560 18165 2565 18195
rect 2595 18165 2600 18195
rect 2560 18160 2600 18165
rect 2640 18195 2680 18200
rect 2640 18165 2645 18195
rect 2675 18165 2680 18195
rect 2640 18160 2680 18165
rect 2720 18195 2760 18200
rect 2720 18165 2725 18195
rect 2755 18165 2760 18195
rect 2720 18160 2760 18165
rect 2800 18195 2840 18200
rect 2800 18165 2805 18195
rect 2835 18165 2840 18195
rect 2800 18160 2840 18165
rect 2880 18195 2920 18200
rect 2880 18165 2885 18195
rect 2915 18165 2920 18195
rect 2880 18160 2920 18165
rect 2960 18195 3000 18200
rect 2960 18165 2965 18195
rect 2995 18165 3000 18195
rect 2960 18160 3000 18165
rect 3040 18195 3080 18200
rect 3040 18165 3045 18195
rect 3075 18165 3080 18195
rect 3040 18160 3080 18165
rect 3120 18195 3160 18200
rect 3120 18165 3125 18195
rect 3155 18165 3160 18195
rect 3120 18160 3160 18165
rect 3200 18195 3240 18200
rect 3200 18165 3205 18195
rect 3235 18165 3240 18195
rect 3200 18160 3240 18165
rect 3280 18195 3320 18200
rect 3280 18165 3285 18195
rect 3315 18165 3320 18195
rect 3280 18160 3320 18165
rect 3360 18195 3400 18200
rect 3360 18165 3365 18195
rect 3395 18165 3400 18195
rect 3360 18160 3400 18165
rect 3440 18195 3480 18200
rect 3440 18165 3445 18195
rect 3475 18165 3480 18195
rect 3440 18160 3480 18165
rect 3520 18195 3560 18200
rect 3520 18165 3525 18195
rect 3555 18165 3560 18195
rect 3520 18160 3560 18165
rect 3600 18195 3640 18200
rect 3600 18165 3605 18195
rect 3635 18165 3640 18195
rect 3600 18160 3640 18165
rect 3680 18195 3720 18200
rect 3680 18165 3685 18195
rect 3715 18165 3720 18195
rect 3680 18160 3720 18165
rect 3760 18195 3800 18200
rect 3760 18165 3765 18195
rect 3795 18165 3800 18195
rect 3760 18160 3800 18165
rect 3840 18195 3880 18200
rect 3840 18165 3845 18195
rect 3875 18165 3880 18195
rect 3840 18160 3880 18165
rect 3920 18195 3960 18200
rect 3920 18165 3925 18195
rect 3955 18165 3960 18195
rect 3920 18160 3960 18165
rect 4000 18195 4040 18200
rect 4000 18165 4005 18195
rect 4035 18165 4040 18195
rect 4000 18160 4040 18165
rect 4080 18195 4120 18200
rect 4080 18165 4085 18195
rect 4115 18165 4120 18195
rect 4080 18160 4120 18165
rect 4160 18195 4200 18200
rect 4160 18165 4165 18195
rect 4195 18165 4200 18195
rect 4160 18160 4200 18165
rect 6240 18195 6280 18200
rect 6240 18165 6245 18195
rect 6275 18165 6280 18195
rect 6240 18160 6280 18165
rect 6320 18195 6360 18200
rect 6320 18165 6325 18195
rect 6355 18165 6360 18195
rect 6320 18160 6360 18165
rect 6400 18195 6440 18200
rect 6400 18165 6405 18195
rect 6435 18165 6440 18195
rect 6400 18160 6440 18165
rect 6480 18195 6520 18200
rect 6480 18165 6485 18195
rect 6515 18165 6520 18195
rect 6480 18160 6520 18165
rect 6560 18195 6600 18200
rect 6560 18165 6565 18195
rect 6595 18165 6600 18195
rect 6560 18160 6600 18165
rect 6640 18195 6680 18200
rect 6640 18165 6645 18195
rect 6675 18165 6680 18195
rect 6640 18160 6680 18165
rect 6720 18195 6760 18200
rect 6720 18165 6725 18195
rect 6755 18165 6760 18195
rect 6720 18160 6760 18165
rect 6800 18195 6840 18200
rect 6800 18165 6805 18195
rect 6835 18165 6840 18195
rect 6800 18160 6840 18165
rect 6880 18195 6920 18200
rect 6880 18165 6885 18195
rect 6915 18165 6920 18195
rect 6880 18160 6920 18165
rect 6960 18195 7000 18200
rect 6960 18165 6965 18195
rect 6995 18165 7000 18195
rect 6960 18160 7000 18165
rect 7040 18195 7080 18200
rect 7040 18165 7045 18195
rect 7075 18165 7080 18195
rect 7040 18160 7080 18165
rect 7120 18195 7160 18200
rect 7120 18165 7125 18195
rect 7155 18165 7160 18195
rect 7120 18160 7160 18165
rect 7200 18195 7240 18200
rect 7200 18165 7205 18195
rect 7235 18165 7240 18195
rect 7200 18160 7240 18165
rect 7280 18195 7320 18200
rect 7280 18165 7285 18195
rect 7315 18165 7320 18195
rect 7280 18160 7320 18165
rect 7360 18195 7400 18200
rect 7360 18165 7365 18195
rect 7395 18165 7400 18195
rect 7360 18160 7400 18165
rect 7440 18195 7480 18200
rect 7440 18165 7445 18195
rect 7475 18165 7480 18195
rect 7440 18160 7480 18165
rect 7520 18195 7560 18200
rect 7520 18165 7525 18195
rect 7555 18165 7560 18195
rect 7520 18160 7560 18165
rect 7600 18195 7640 18200
rect 7600 18165 7605 18195
rect 7635 18165 7640 18195
rect 7600 18160 7640 18165
rect 7680 18195 7720 18200
rect 7680 18165 7685 18195
rect 7715 18165 7720 18195
rect 7680 18160 7720 18165
rect 7760 18195 7800 18200
rect 7760 18165 7765 18195
rect 7795 18165 7800 18195
rect 7760 18160 7800 18165
rect 7840 18195 7880 18200
rect 7840 18165 7845 18195
rect 7875 18165 7880 18195
rect 7840 18160 7880 18165
rect 7920 18195 7960 18200
rect 7920 18165 7925 18195
rect 7955 18165 7960 18195
rect 7920 18160 7960 18165
rect 8000 18195 8040 18200
rect 8000 18165 8005 18195
rect 8035 18165 8040 18195
rect 8000 18160 8040 18165
rect 8080 18195 8120 18200
rect 8080 18165 8085 18195
rect 8115 18165 8120 18195
rect 8080 18160 8120 18165
rect 8160 18195 8200 18200
rect 8160 18165 8165 18195
rect 8195 18165 8200 18195
rect 8160 18160 8200 18165
rect 8240 18195 8280 18200
rect 8240 18165 8245 18195
rect 8275 18165 8280 18195
rect 8240 18160 8280 18165
rect 8320 18195 8360 18200
rect 8320 18165 8325 18195
rect 8355 18165 8360 18195
rect 8320 18160 8360 18165
rect 8400 18195 8440 18200
rect 8400 18165 8405 18195
rect 8435 18165 8440 18195
rect 8400 18160 8440 18165
rect 8480 18195 8520 18200
rect 8480 18165 8485 18195
rect 8515 18165 8520 18195
rect 8480 18160 8520 18165
rect 8560 18195 8600 18200
rect 8560 18165 8565 18195
rect 8595 18165 8600 18195
rect 8560 18160 8600 18165
rect 8640 18195 8680 18200
rect 8640 18165 8645 18195
rect 8675 18165 8680 18195
rect 8640 18160 8680 18165
rect 8720 18195 8760 18200
rect 8720 18165 8725 18195
rect 8755 18165 8760 18195
rect 8720 18160 8760 18165
rect 8800 18195 8840 18200
rect 8800 18165 8805 18195
rect 8835 18165 8840 18195
rect 8800 18160 8840 18165
rect 8880 18195 8920 18200
rect 8880 18165 8885 18195
rect 8915 18165 8920 18195
rect 8880 18160 8920 18165
rect 8960 18195 9000 18200
rect 8960 18165 8965 18195
rect 8995 18165 9000 18195
rect 8960 18160 9000 18165
rect 9040 18195 9080 18200
rect 9040 18165 9045 18195
rect 9075 18165 9080 18195
rect 9040 18160 9080 18165
rect 9120 18195 9160 18200
rect 9120 18165 9125 18195
rect 9155 18165 9160 18195
rect 9120 18160 9160 18165
rect 9200 18195 9240 18200
rect 9200 18165 9205 18195
rect 9235 18165 9240 18195
rect 9200 18160 9240 18165
rect 9280 18195 9320 18200
rect 9280 18165 9285 18195
rect 9315 18165 9320 18195
rect 9280 18160 9320 18165
rect 9360 18195 9400 18200
rect 9360 18165 9365 18195
rect 9395 18165 9400 18195
rect 9360 18160 9400 18165
rect 9440 18195 9480 18200
rect 9440 18165 9445 18195
rect 9475 18165 9480 18195
rect 9440 18160 9480 18165
rect 11560 18195 11600 18200
rect 11560 18165 11565 18195
rect 11595 18165 11600 18195
rect 11560 18160 11600 18165
rect 11640 18195 11680 18200
rect 11640 18165 11645 18195
rect 11675 18165 11680 18195
rect 11640 18160 11680 18165
rect 11720 18195 11760 18200
rect 11720 18165 11725 18195
rect 11755 18165 11760 18195
rect 11720 18160 11760 18165
rect 11800 18195 11840 18200
rect 11800 18165 11805 18195
rect 11835 18165 11840 18195
rect 11800 18160 11840 18165
rect 11880 18195 11920 18200
rect 11880 18165 11885 18195
rect 11915 18165 11920 18195
rect 11880 18160 11920 18165
rect 11960 18195 12000 18200
rect 11960 18165 11965 18195
rect 11995 18165 12000 18195
rect 11960 18160 12000 18165
rect 12040 18195 12080 18200
rect 12040 18165 12045 18195
rect 12075 18165 12080 18195
rect 12040 18160 12080 18165
rect 12120 18195 12160 18200
rect 12120 18165 12125 18195
rect 12155 18165 12160 18195
rect 12120 18160 12160 18165
rect 12200 18195 12240 18200
rect 12200 18165 12205 18195
rect 12235 18165 12240 18195
rect 12200 18160 12240 18165
rect 12280 18195 12320 18200
rect 12280 18165 12285 18195
rect 12315 18165 12320 18195
rect 12280 18160 12320 18165
rect 12360 18195 12400 18200
rect 12360 18165 12365 18195
rect 12395 18165 12400 18195
rect 12360 18160 12400 18165
rect 12440 18195 12480 18200
rect 12440 18165 12445 18195
rect 12475 18165 12480 18195
rect 12440 18160 12480 18165
rect 12520 18195 12560 18200
rect 12520 18165 12525 18195
rect 12555 18165 12560 18195
rect 12520 18160 12560 18165
rect 12600 18195 12640 18200
rect 12600 18165 12605 18195
rect 12635 18165 12640 18195
rect 12600 18160 12640 18165
rect 12680 18195 12720 18200
rect 12680 18165 12685 18195
rect 12715 18165 12720 18195
rect 12680 18160 12720 18165
rect 12760 18195 12800 18200
rect 12760 18165 12765 18195
rect 12795 18165 12800 18195
rect 12760 18160 12800 18165
rect 12840 18195 12880 18200
rect 12840 18165 12845 18195
rect 12875 18165 12880 18195
rect 12840 18160 12880 18165
rect 12920 18195 12960 18200
rect 12920 18165 12925 18195
rect 12955 18165 12960 18195
rect 12920 18160 12960 18165
rect 13000 18195 13040 18200
rect 13000 18165 13005 18195
rect 13035 18165 13040 18195
rect 13000 18160 13040 18165
rect 13080 18195 13120 18200
rect 13080 18165 13085 18195
rect 13115 18165 13120 18195
rect 13080 18160 13120 18165
rect 13160 18195 13200 18200
rect 13160 18165 13165 18195
rect 13195 18165 13200 18195
rect 13160 18160 13200 18165
rect 13240 18195 13280 18200
rect 13240 18165 13245 18195
rect 13275 18165 13280 18195
rect 13240 18160 13280 18165
rect 13320 18195 13360 18200
rect 13320 18165 13325 18195
rect 13355 18165 13360 18195
rect 13320 18160 13360 18165
rect 13400 18195 13440 18200
rect 13400 18165 13405 18195
rect 13435 18165 13440 18195
rect 13400 18160 13440 18165
rect 13480 18195 13520 18200
rect 13480 18165 13485 18195
rect 13515 18165 13520 18195
rect 13480 18160 13520 18165
rect 13560 18195 13600 18200
rect 13560 18165 13565 18195
rect 13595 18165 13600 18195
rect 13560 18160 13600 18165
rect 13640 18195 13680 18200
rect 13640 18165 13645 18195
rect 13675 18165 13680 18195
rect 13640 18160 13680 18165
rect 13720 18195 13760 18200
rect 13720 18165 13725 18195
rect 13755 18165 13760 18195
rect 13720 18160 13760 18165
rect 13800 18195 13840 18200
rect 13800 18165 13805 18195
rect 13835 18165 13840 18195
rect 13800 18160 13840 18165
rect 13880 18195 13920 18200
rect 13880 18165 13885 18195
rect 13915 18165 13920 18195
rect 13880 18160 13920 18165
rect 13960 18195 14000 18200
rect 13960 18165 13965 18195
rect 13995 18165 14000 18195
rect 13960 18160 14000 18165
rect 14040 18195 14080 18200
rect 14040 18165 14045 18195
rect 14075 18165 14080 18195
rect 14040 18160 14080 18165
rect 14120 18195 14160 18200
rect 14120 18165 14125 18195
rect 14155 18165 14160 18195
rect 14120 18160 14160 18165
rect 14200 18195 14240 18200
rect 14200 18165 14205 18195
rect 14235 18165 14240 18195
rect 14200 18160 14240 18165
rect 14280 18195 14320 18200
rect 14280 18165 14285 18195
rect 14315 18165 14320 18195
rect 14280 18160 14320 18165
rect 14360 18195 14400 18200
rect 14360 18165 14365 18195
rect 14395 18165 14400 18195
rect 14360 18160 14400 18165
rect 14440 18195 14480 18200
rect 14440 18165 14445 18195
rect 14475 18165 14480 18195
rect 14440 18160 14480 18165
rect 14520 18195 14560 18200
rect 14520 18165 14525 18195
rect 14555 18165 14560 18195
rect 14520 18160 14560 18165
rect 14600 18195 14640 18200
rect 14600 18165 14605 18195
rect 14635 18165 14640 18195
rect 14600 18160 14640 18165
rect 14680 18195 14720 18200
rect 14680 18165 14685 18195
rect 14715 18165 14720 18195
rect 14680 18160 14720 18165
rect 16760 18195 16800 18200
rect 16760 18165 16765 18195
rect 16795 18165 16800 18195
rect 16760 18160 16800 18165
rect 16840 18195 16880 18200
rect 16840 18165 16845 18195
rect 16875 18165 16880 18195
rect 16840 18160 16880 18165
rect 16920 18195 16960 18200
rect 16920 18165 16925 18195
rect 16955 18165 16960 18195
rect 16920 18160 16960 18165
rect 17000 18195 17040 18200
rect 17000 18165 17005 18195
rect 17035 18165 17040 18195
rect 17000 18160 17040 18165
rect 17080 18195 17120 18200
rect 17080 18165 17085 18195
rect 17115 18165 17120 18195
rect 17080 18160 17120 18165
rect 17160 18195 17200 18200
rect 17160 18165 17165 18195
rect 17195 18165 17200 18195
rect 17160 18160 17200 18165
rect 17240 18195 17280 18200
rect 17240 18165 17245 18195
rect 17275 18165 17280 18195
rect 17240 18160 17280 18165
rect 17320 18195 17360 18200
rect 17320 18165 17325 18195
rect 17355 18165 17360 18195
rect 17320 18160 17360 18165
rect 17400 18195 17440 18200
rect 17400 18165 17405 18195
rect 17435 18165 17440 18195
rect 17400 18160 17440 18165
rect 17480 18195 17520 18200
rect 17480 18165 17485 18195
rect 17515 18165 17520 18195
rect 17480 18160 17520 18165
rect 17560 18195 17600 18200
rect 17560 18165 17565 18195
rect 17595 18165 17600 18195
rect 17560 18160 17600 18165
rect 17640 18195 17680 18200
rect 17640 18165 17645 18195
rect 17675 18165 17680 18195
rect 17640 18160 17680 18165
rect 17720 18195 17760 18200
rect 17720 18165 17725 18195
rect 17755 18165 17760 18195
rect 17720 18160 17760 18165
rect 17800 18195 17840 18200
rect 17800 18165 17805 18195
rect 17835 18165 17840 18195
rect 17800 18160 17840 18165
rect 17880 18195 17920 18200
rect 17880 18165 17885 18195
rect 17915 18165 17920 18195
rect 17880 18160 17920 18165
rect 17960 18195 18000 18200
rect 17960 18165 17965 18195
rect 17995 18165 18000 18195
rect 17960 18160 18000 18165
rect 18040 18195 18080 18200
rect 18040 18165 18045 18195
rect 18075 18165 18080 18195
rect 18040 18160 18080 18165
rect 18120 18195 18160 18200
rect 18120 18165 18125 18195
rect 18155 18165 18160 18195
rect 18120 18160 18160 18165
rect 18200 18195 18240 18200
rect 18200 18165 18205 18195
rect 18235 18165 18240 18195
rect 18200 18160 18240 18165
rect 18280 18195 18320 18200
rect 18280 18165 18285 18195
rect 18315 18165 18320 18195
rect 18280 18160 18320 18165
rect 18360 18195 18400 18200
rect 18360 18165 18365 18195
rect 18395 18165 18400 18195
rect 18360 18160 18400 18165
rect 18440 18195 18480 18200
rect 18440 18165 18445 18195
rect 18475 18165 18480 18195
rect 18440 18160 18480 18165
rect 18520 18195 18560 18200
rect 18520 18165 18525 18195
rect 18555 18165 18560 18195
rect 18520 18160 18560 18165
rect 18600 18195 18640 18200
rect 18600 18165 18605 18195
rect 18635 18165 18640 18195
rect 18600 18160 18640 18165
rect 18680 18195 18720 18200
rect 18680 18165 18685 18195
rect 18715 18165 18720 18195
rect 18680 18160 18720 18165
rect 18760 18195 18800 18200
rect 18760 18165 18765 18195
rect 18795 18165 18800 18195
rect 18760 18160 18800 18165
rect 18840 18195 18880 18200
rect 18840 18165 18845 18195
rect 18875 18165 18880 18195
rect 18840 18160 18880 18165
rect 18920 18195 18960 18200
rect 18920 18165 18925 18195
rect 18955 18165 18960 18195
rect 18920 18160 18960 18165
rect 19000 18195 19040 18200
rect 19000 18165 19005 18195
rect 19035 18165 19040 18195
rect 19000 18160 19040 18165
rect 19080 18195 19120 18200
rect 19080 18165 19085 18195
rect 19115 18165 19120 18195
rect 19080 18160 19120 18165
rect 19160 18195 19200 18200
rect 19160 18165 19165 18195
rect 19195 18165 19200 18195
rect 19160 18160 19200 18165
rect 19240 18195 19280 18200
rect 19240 18165 19245 18195
rect 19275 18165 19280 18195
rect 19240 18160 19280 18165
rect 19320 18195 19360 18200
rect 19320 18165 19325 18195
rect 19355 18165 19360 18195
rect 19320 18160 19360 18165
rect 19400 18195 19440 18200
rect 19400 18165 19405 18195
rect 19435 18165 19440 18195
rect 19400 18160 19440 18165
rect 19480 18195 19520 18200
rect 19480 18165 19485 18195
rect 19515 18165 19520 18195
rect 19480 18160 19520 18165
rect 19560 18195 19600 18200
rect 19560 18165 19565 18195
rect 19595 18165 19600 18195
rect 19560 18160 19600 18165
rect 19640 18195 19680 18200
rect 19640 18165 19645 18195
rect 19675 18165 19680 18195
rect 19640 18160 19680 18165
rect 19720 18195 19760 18200
rect 19720 18165 19725 18195
rect 19755 18165 19760 18195
rect 19720 18160 19760 18165
rect 19800 18195 19840 18200
rect 19800 18165 19805 18195
rect 19835 18165 19840 18195
rect 19800 18160 19840 18165
rect 19880 18195 19920 18200
rect 19880 18165 19885 18195
rect 19915 18165 19920 18195
rect 19880 18160 19920 18165
rect 19960 18195 20000 18200
rect 19960 18165 19965 18195
rect 19995 18165 20000 18195
rect 19960 18160 20000 18165
rect 20040 18195 20080 18200
rect 20040 18165 20045 18195
rect 20075 18165 20080 18195
rect 20040 18160 20080 18165
rect 20120 18195 20160 18200
rect 20120 18165 20125 18195
rect 20155 18165 20160 18195
rect 20120 18160 20160 18165
rect 20200 18195 20240 18200
rect 20200 18165 20205 18195
rect 20235 18165 20240 18195
rect 20200 18160 20240 18165
rect 20280 18195 20320 18200
rect 20280 18165 20285 18195
rect 20315 18165 20320 18195
rect 20280 18160 20320 18165
rect 20360 18195 20400 18200
rect 20360 18165 20365 18195
rect 20395 18165 20400 18195
rect 20360 18160 20400 18165
rect 20440 18195 20480 18200
rect 20440 18165 20445 18195
rect 20475 18165 20480 18195
rect 20440 18160 20480 18165
rect 20520 18195 20560 18200
rect 20520 18165 20525 18195
rect 20555 18165 20560 18195
rect 20520 18160 20560 18165
rect 20600 18195 20640 18200
rect 20600 18165 20605 18195
rect 20635 18165 20640 18195
rect 20600 18160 20640 18165
rect 20680 18195 20720 18200
rect 20680 18165 20685 18195
rect 20715 18165 20720 18195
rect 20680 18160 20720 18165
rect 20760 18195 20800 18200
rect 20760 18165 20765 18195
rect 20795 18165 20800 18195
rect 20760 18160 20800 18165
rect 20840 18195 20880 18200
rect 20840 18165 20845 18195
rect 20875 18165 20880 18195
rect 20840 18160 20880 18165
rect 20920 18195 20960 18200
rect 20920 18165 20925 18195
rect 20955 18165 20960 18195
rect 20920 18160 20960 18165
rect 0 18035 40 18040
rect 0 18005 5 18035
rect 35 18005 40 18035
rect 0 18000 40 18005
rect 80 18035 120 18040
rect 80 18005 85 18035
rect 115 18005 120 18035
rect 80 18000 120 18005
rect 160 18035 200 18040
rect 160 18005 165 18035
rect 195 18005 200 18035
rect 160 18000 200 18005
rect 240 18035 280 18040
rect 240 18005 245 18035
rect 275 18005 280 18035
rect 240 18000 280 18005
rect 320 18035 360 18040
rect 320 18005 325 18035
rect 355 18005 360 18035
rect 320 18000 360 18005
rect 400 18035 440 18040
rect 400 18005 405 18035
rect 435 18005 440 18035
rect 400 18000 440 18005
rect 480 18035 520 18040
rect 480 18005 485 18035
rect 515 18005 520 18035
rect 480 18000 520 18005
rect 560 18035 600 18040
rect 560 18005 565 18035
rect 595 18005 600 18035
rect 560 18000 600 18005
rect 640 18035 680 18040
rect 640 18005 645 18035
rect 675 18005 680 18035
rect 640 18000 680 18005
rect 720 18035 760 18040
rect 720 18005 725 18035
rect 755 18005 760 18035
rect 720 18000 760 18005
rect 800 18035 840 18040
rect 800 18005 805 18035
rect 835 18005 840 18035
rect 800 18000 840 18005
rect 880 18035 920 18040
rect 880 18005 885 18035
rect 915 18005 920 18035
rect 880 18000 920 18005
rect 960 18035 1000 18040
rect 960 18005 965 18035
rect 995 18005 1000 18035
rect 960 18000 1000 18005
rect 1040 18035 1080 18040
rect 1040 18005 1045 18035
rect 1075 18005 1080 18035
rect 1040 18000 1080 18005
rect 1120 18035 1160 18040
rect 1120 18005 1125 18035
rect 1155 18005 1160 18035
rect 1120 18000 1160 18005
rect 1200 18035 1240 18040
rect 1200 18005 1205 18035
rect 1235 18005 1240 18035
rect 1200 18000 1240 18005
rect 1280 18035 1320 18040
rect 1280 18005 1285 18035
rect 1315 18005 1320 18035
rect 1280 18000 1320 18005
rect 1360 18035 1400 18040
rect 1360 18005 1365 18035
rect 1395 18005 1400 18035
rect 1360 18000 1400 18005
rect 1440 18035 1480 18040
rect 1440 18005 1445 18035
rect 1475 18005 1480 18035
rect 1440 18000 1480 18005
rect 1520 18035 1560 18040
rect 1520 18005 1525 18035
rect 1555 18005 1560 18035
rect 1520 18000 1560 18005
rect 1600 18035 1640 18040
rect 1600 18005 1605 18035
rect 1635 18005 1640 18035
rect 1600 18000 1640 18005
rect 1680 18035 1720 18040
rect 1680 18005 1685 18035
rect 1715 18005 1720 18035
rect 1680 18000 1720 18005
rect 1760 18035 1800 18040
rect 1760 18005 1765 18035
rect 1795 18005 1800 18035
rect 1760 18000 1800 18005
rect 1840 18035 1880 18040
rect 1840 18005 1845 18035
rect 1875 18005 1880 18035
rect 1840 18000 1880 18005
rect 1920 18035 1960 18040
rect 1920 18005 1925 18035
rect 1955 18005 1960 18035
rect 1920 18000 1960 18005
rect 2000 18035 2040 18040
rect 2000 18005 2005 18035
rect 2035 18005 2040 18035
rect 2000 18000 2040 18005
rect 2080 18035 2120 18040
rect 2080 18005 2085 18035
rect 2115 18005 2120 18035
rect 2080 18000 2120 18005
rect 2160 18035 2200 18040
rect 2160 18005 2165 18035
rect 2195 18005 2200 18035
rect 2160 18000 2200 18005
rect 2240 18035 2280 18040
rect 2240 18005 2245 18035
rect 2275 18005 2280 18035
rect 2240 18000 2280 18005
rect 2320 18035 2360 18040
rect 2320 18005 2325 18035
rect 2355 18005 2360 18035
rect 2320 18000 2360 18005
rect 2400 18035 2440 18040
rect 2400 18005 2405 18035
rect 2435 18005 2440 18035
rect 2400 18000 2440 18005
rect 2480 18035 2520 18040
rect 2480 18005 2485 18035
rect 2515 18005 2520 18035
rect 2480 18000 2520 18005
rect 2560 18035 2600 18040
rect 2560 18005 2565 18035
rect 2595 18005 2600 18035
rect 2560 18000 2600 18005
rect 2640 18035 2680 18040
rect 2640 18005 2645 18035
rect 2675 18005 2680 18035
rect 2640 18000 2680 18005
rect 2720 18035 2760 18040
rect 2720 18005 2725 18035
rect 2755 18005 2760 18035
rect 2720 18000 2760 18005
rect 2800 18035 2840 18040
rect 2800 18005 2805 18035
rect 2835 18005 2840 18035
rect 2800 18000 2840 18005
rect 2880 18035 2920 18040
rect 2880 18005 2885 18035
rect 2915 18005 2920 18035
rect 2880 18000 2920 18005
rect 2960 18035 3000 18040
rect 2960 18005 2965 18035
rect 2995 18005 3000 18035
rect 2960 18000 3000 18005
rect 3040 18035 3080 18040
rect 3040 18005 3045 18035
rect 3075 18005 3080 18035
rect 3040 18000 3080 18005
rect 3120 18035 3160 18040
rect 3120 18005 3125 18035
rect 3155 18005 3160 18035
rect 3120 18000 3160 18005
rect 3200 18035 3240 18040
rect 3200 18005 3205 18035
rect 3235 18005 3240 18035
rect 3200 18000 3240 18005
rect 3280 18035 3320 18040
rect 3280 18005 3285 18035
rect 3315 18005 3320 18035
rect 3280 18000 3320 18005
rect 3360 18035 3400 18040
rect 3360 18005 3365 18035
rect 3395 18005 3400 18035
rect 3360 18000 3400 18005
rect 3440 18035 3480 18040
rect 3440 18005 3445 18035
rect 3475 18005 3480 18035
rect 3440 18000 3480 18005
rect 3520 18035 3560 18040
rect 3520 18005 3525 18035
rect 3555 18005 3560 18035
rect 3520 18000 3560 18005
rect 3600 18035 3640 18040
rect 3600 18005 3605 18035
rect 3635 18005 3640 18035
rect 3600 18000 3640 18005
rect 3680 18035 3720 18040
rect 3680 18005 3685 18035
rect 3715 18005 3720 18035
rect 3680 18000 3720 18005
rect 3760 18035 3800 18040
rect 3760 18005 3765 18035
rect 3795 18005 3800 18035
rect 3760 18000 3800 18005
rect 3840 18035 3880 18040
rect 3840 18005 3845 18035
rect 3875 18005 3880 18035
rect 3840 18000 3880 18005
rect 3920 18035 3960 18040
rect 3920 18005 3925 18035
rect 3955 18005 3960 18035
rect 3920 18000 3960 18005
rect 4000 18035 4040 18040
rect 4000 18005 4005 18035
rect 4035 18005 4040 18035
rect 4000 18000 4040 18005
rect 4080 18035 4120 18040
rect 4080 18005 4085 18035
rect 4115 18005 4120 18035
rect 4080 18000 4120 18005
rect 4160 18035 4200 18040
rect 4160 18005 4165 18035
rect 4195 18005 4200 18035
rect 4160 18000 4200 18005
rect 6240 18035 6280 18040
rect 6240 18005 6245 18035
rect 6275 18005 6280 18035
rect 6240 18000 6280 18005
rect 6320 18035 6360 18040
rect 6320 18005 6325 18035
rect 6355 18005 6360 18035
rect 6320 18000 6360 18005
rect 6400 18035 6440 18040
rect 6400 18005 6405 18035
rect 6435 18005 6440 18035
rect 6400 18000 6440 18005
rect 6480 18035 6520 18040
rect 6480 18005 6485 18035
rect 6515 18005 6520 18035
rect 6480 18000 6520 18005
rect 6560 18035 6600 18040
rect 6560 18005 6565 18035
rect 6595 18005 6600 18035
rect 6560 18000 6600 18005
rect 6640 18035 6680 18040
rect 6640 18005 6645 18035
rect 6675 18005 6680 18035
rect 6640 18000 6680 18005
rect 6720 18035 6760 18040
rect 6720 18005 6725 18035
rect 6755 18005 6760 18035
rect 6720 18000 6760 18005
rect 6800 18035 6840 18040
rect 6800 18005 6805 18035
rect 6835 18005 6840 18035
rect 6800 18000 6840 18005
rect 6880 18035 6920 18040
rect 6880 18005 6885 18035
rect 6915 18005 6920 18035
rect 6880 18000 6920 18005
rect 6960 18035 7000 18040
rect 6960 18005 6965 18035
rect 6995 18005 7000 18035
rect 6960 18000 7000 18005
rect 7040 18035 7080 18040
rect 7040 18005 7045 18035
rect 7075 18005 7080 18035
rect 7040 18000 7080 18005
rect 7120 18035 7160 18040
rect 7120 18005 7125 18035
rect 7155 18005 7160 18035
rect 7120 18000 7160 18005
rect 7200 18035 7240 18040
rect 7200 18005 7205 18035
rect 7235 18005 7240 18035
rect 7200 18000 7240 18005
rect 7280 18035 7320 18040
rect 7280 18005 7285 18035
rect 7315 18005 7320 18035
rect 7280 18000 7320 18005
rect 7360 18035 7400 18040
rect 7360 18005 7365 18035
rect 7395 18005 7400 18035
rect 7360 18000 7400 18005
rect 7440 18035 7480 18040
rect 7440 18005 7445 18035
rect 7475 18005 7480 18035
rect 7440 18000 7480 18005
rect 7520 18035 7560 18040
rect 7520 18005 7525 18035
rect 7555 18005 7560 18035
rect 7520 18000 7560 18005
rect 7600 18035 7640 18040
rect 7600 18005 7605 18035
rect 7635 18005 7640 18035
rect 7600 18000 7640 18005
rect 7680 18035 7720 18040
rect 7680 18005 7685 18035
rect 7715 18005 7720 18035
rect 7680 18000 7720 18005
rect 7760 18035 7800 18040
rect 7760 18005 7765 18035
rect 7795 18005 7800 18035
rect 7760 18000 7800 18005
rect 7840 18035 7880 18040
rect 7840 18005 7845 18035
rect 7875 18005 7880 18035
rect 7840 18000 7880 18005
rect 7920 18035 7960 18040
rect 7920 18005 7925 18035
rect 7955 18005 7960 18035
rect 7920 18000 7960 18005
rect 8000 18035 8040 18040
rect 8000 18005 8005 18035
rect 8035 18005 8040 18035
rect 8000 18000 8040 18005
rect 8080 18035 8120 18040
rect 8080 18005 8085 18035
rect 8115 18005 8120 18035
rect 8080 18000 8120 18005
rect 8160 18035 8200 18040
rect 8160 18005 8165 18035
rect 8195 18005 8200 18035
rect 8160 18000 8200 18005
rect 8240 18035 8280 18040
rect 8240 18005 8245 18035
rect 8275 18005 8280 18035
rect 8240 18000 8280 18005
rect 8320 18035 8360 18040
rect 8320 18005 8325 18035
rect 8355 18005 8360 18035
rect 8320 18000 8360 18005
rect 8400 18035 8440 18040
rect 8400 18005 8405 18035
rect 8435 18005 8440 18035
rect 8400 18000 8440 18005
rect 8480 18035 8520 18040
rect 8480 18005 8485 18035
rect 8515 18005 8520 18035
rect 8480 18000 8520 18005
rect 8560 18035 8600 18040
rect 8560 18005 8565 18035
rect 8595 18005 8600 18035
rect 8560 18000 8600 18005
rect 8640 18035 8680 18040
rect 8640 18005 8645 18035
rect 8675 18005 8680 18035
rect 8640 18000 8680 18005
rect 8720 18035 8760 18040
rect 8720 18005 8725 18035
rect 8755 18005 8760 18035
rect 8720 18000 8760 18005
rect 8800 18035 8840 18040
rect 8800 18005 8805 18035
rect 8835 18005 8840 18035
rect 8800 18000 8840 18005
rect 8880 18035 8920 18040
rect 8880 18005 8885 18035
rect 8915 18005 8920 18035
rect 8880 18000 8920 18005
rect 8960 18035 9000 18040
rect 8960 18005 8965 18035
rect 8995 18005 9000 18035
rect 8960 18000 9000 18005
rect 9040 18035 9080 18040
rect 9040 18005 9045 18035
rect 9075 18005 9080 18035
rect 9040 18000 9080 18005
rect 9120 18035 9160 18040
rect 9120 18005 9125 18035
rect 9155 18005 9160 18035
rect 9120 18000 9160 18005
rect 9200 18035 9240 18040
rect 9200 18005 9205 18035
rect 9235 18005 9240 18035
rect 9200 18000 9240 18005
rect 9280 18035 9320 18040
rect 9280 18005 9285 18035
rect 9315 18005 9320 18035
rect 9280 18000 9320 18005
rect 9360 18035 9400 18040
rect 9360 18005 9365 18035
rect 9395 18005 9400 18035
rect 9360 18000 9400 18005
rect 9440 18035 9480 18040
rect 9440 18005 9445 18035
rect 9475 18005 9480 18035
rect 9440 18000 9480 18005
rect 11560 18035 11600 18040
rect 11560 18005 11565 18035
rect 11595 18005 11600 18035
rect 11560 18000 11600 18005
rect 11640 18035 11680 18040
rect 11640 18005 11645 18035
rect 11675 18005 11680 18035
rect 11640 18000 11680 18005
rect 11720 18035 11760 18040
rect 11720 18005 11725 18035
rect 11755 18005 11760 18035
rect 11720 18000 11760 18005
rect 11800 18035 11840 18040
rect 11800 18005 11805 18035
rect 11835 18005 11840 18035
rect 11800 18000 11840 18005
rect 11880 18035 11920 18040
rect 11880 18005 11885 18035
rect 11915 18005 11920 18035
rect 11880 18000 11920 18005
rect 11960 18035 12000 18040
rect 11960 18005 11965 18035
rect 11995 18005 12000 18035
rect 11960 18000 12000 18005
rect 12040 18035 12080 18040
rect 12040 18005 12045 18035
rect 12075 18005 12080 18035
rect 12040 18000 12080 18005
rect 12120 18035 12160 18040
rect 12120 18005 12125 18035
rect 12155 18005 12160 18035
rect 12120 18000 12160 18005
rect 12200 18035 12240 18040
rect 12200 18005 12205 18035
rect 12235 18005 12240 18035
rect 12200 18000 12240 18005
rect 12280 18035 12320 18040
rect 12280 18005 12285 18035
rect 12315 18005 12320 18035
rect 12280 18000 12320 18005
rect 12360 18035 12400 18040
rect 12360 18005 12365 18035
rect 12395 18005 12400 18035
rect 12360 18000 12400 18005
rect 12440 18035 12480 18040
rect 12440 18005 12445 18035
rect 12475 18005 12480 18035
rect 12440 18000 12480 18005
rect 12520 18035 12560 18040
rect 12520 18005 12525 18035
rect 12555 18005 12560 18035
rect 12520 18000 12560 18005
rect 12600 18035 12640 18040
rect 12600 18005 12605 18035
rect 12635 18005 12640 18035
rect 12600 18000 12640 18005
rect 12680 18035 12720 18040
rect 12680 18005 12685 18035
rect 12715 18005 12720 18035
rect 12680 18000 12720 18005
rect 12760 18035 12800 18040
rect 12760 18005 12765 18035
rect 12795 18005 12800 18035
rect 12760 18000 12800 18005
rect 12840 18035 12880 18040
rect 12840 18005 12845 18035
rect 12875 18005 12880 18035
rect 12840 18000 12880 18005
rect 12920 18035 12960 18040
rect 12920 18005 12925 18035
rect 12955 18005 12960 18035
rect 12920 18000 12960 18005
rect 13000 18035 13040 18040
rect 13000 18005 13005 18035
rect 13035 18005 13040 18035
rect 13000 18000 13040 18005
rect 13080 18035 13120 18040
rect 13080 18005 13085 18035
rect 13115 18005 13120 18035
rect 13080 18000 13120 18005
rect 13160 18035 13200 18040
rect 13160 18005 13165 18035
rect 13195 18005 13200 18035
rect 13160 18000 13200 18005
rect 13240 18035 13280 18040
rect 13240 18005 13245 18035
rect 13275 18005 13280 18035
rect 13240 18000 13280 18005
rect 13320 18035 13360 18040
rect 13320 18005 13325 18035
rect 13355 18005 13360 18035
rect 13320 18000 13360 18005
rect 13400 18035 13440 18040
rect 13400 18005 13405 18035
rect 13435 18005 13440 18035
rect 13400 18000 13440 18005
rect 13480 18035 13520 18040
rect 13480 18005 13485 18035
rect 13515 18005 13520 18035
rect 13480 18000 13520 18005
rect 13560 18035 13600 18040
rect 13560 18005 13565 18035
rect 13595 18005 13600 18035
rect 13560 18000 13600 18005
rect 13640 18035 13680 18040
rect 13640 18005 13645 18035
rect 13675 18005 13680 18035
rect 13640 18000 13680 18005
rect 13720 18035 13760 18040
rect 13720 18005 13725 18035
rect 13755 18005 13760 18035
rect 13720 18000 13760 18005
rect 13800 18035 13840 18040
rect 13800 18005 13805 18035
rect 13835 18005 13840 18035
rect 13800 18000 13840 18005
rect 13880 18035 13920 18040
rect 13880 18005 13885 18035
rect 13915 18005 13920 18035
rect 13880 18000 13920 18005
rect 13960 18035 14000 18040
rect 13960 18005 13965 18035
rect 13995 18005 14000 18035
rect 13960 18000 14000 18005
rect 14040 18035 14080 18040
rect 14040 18005 14045 18035
rect 14075 18005 14080 18035
rect 14040 18000 14080 18005
rect 14120 18035 14160 18040
rect 14120 18005 14125 18035
rect 14155 18005 14160 18035
rect 14120 18000 14160 18005
rect 14200 18035 14240 18040
rect 14200 18005 14205 18035
rect 14235 18005 14240 18035
rect 14200 18000 14240 18005
rect 14280 18035 14320 18040
rect 14280 18005 14285 18035
rect 14315 18005 14320 18035
rect 14280 18000 14320 18005
rect 14360 18035 14400 18040
rect 14360 18005 14365 18035
rect 14395 18005 14400 18035
rect 14360 18000 14400 18005
rect 14440 18035 14480 18040
rect 14440 18005 14445 18035
rect 14475 18005 14480 18035
rect 14440 18000 14480 18005
rect 14520 18035 14560 18040
rect 14520 18005 14525 18035
rect 14555 18005 14560 18035
rect 14520 18000 14560 18005
rect 14600 18035 14640 18040
rect 14600 18005 14605 18035
rect 14635 18005 14640 18035
rect 14600 18000 14640 18005
rect 14680 18035 14720 18040
rect 14680 18005 14685 18035
rect 14715 18005 14720 18035
rect 14680 18000 14720 18005
rect 16760 18035 16800 18040
rect 16760 18005 16765 18035
rect 16795 18005 16800 18035
rect 16760 18000 16800 18005
rect 16840 18035 16880 18040
rect 16840 18005 16845 18035
rect 16875 18005 16880 18035
rect 16840 18000 16880 18005
rect 16920 18035 16960 18040
rect 16920 18005 16925 18035
rect 16955 18005 16960 18035
rect 16920 18000 16960 18005
rect 17000 18035 17040 18040
rect 17000 18005 17005 18035
rect 17035 18005 17040 18035
rect 17000 18000 17040 18005
rect 17080 18035 17120 18040
rect 17080 18005 17085 18035
rect 17115 18005 17120 18035
rect 17080 18000 17120 18005
rect 17160 18035 17200 18040
rect 17160 18005 17165 18035
rect 17195 18005 17200 18035
rect 17160 18000 17200 18005
rect 17240 18035 17280 18040
rect 17240 18005 17245 18035
rect 17275 18005 17280 18035
rect 17240 18000 17280 18005
rect 17320 18035 17360 18040
rect 17320 18005 17325 18035
rect 17355 18005 17360 18035
rect 17320 18000 17360 18005
rect 17400 18035 17440 18040
rect 17400 18005 17405 18035
rect 17435 18005 17440 18035
rect 17400 18000 17440 18005
rect 17480 18035 17520 18040
rect 17480 18005 17485 18035
rect 17515 18005 17520 18035
rect 17480 18000 17520 18005
rect 17560 18035 17600 18040
rect 17560 18005 17565 18035
rect 17595 18005 17600 18035
rect 17560 18000 17600 18005
rect 17640 18035 17680 18040
rect 17640 18005 17645 18035
rect 17675 18005 17680 18035
rect 17640 18000 17680 18005
rect 17720 18035 17760 18040
rect 17720 18005 17725 18035
rect 17755 18005 17760 18035
rect 17720 18000 17760 18005
rect 17800 18035 17840 18040
rect 17800 18005 17805 18035
rect 17835 18005 17840 18035
rect 17800 18000 17840 18005
rect 17880 18035 17920 18040
rect 17880 18005 17885 18035
rect 17915 18005 17920 18035
rect 17880 18000 17920 18005
rect 17960 18035 18000 18040
rect 17960 18005 17965 18035
rect 17995 18005 18000 18035
rect 17960 18000 18000 18005
rect 18040 18035 18080 18040
rect 18040 18005 18045 18035
rect 18075 18005 18080 18035
rect 18040 18000 18080 18005
rect 18120 18035 18160 18040
rect 18120 18005 18125 18035
rect 18155 18005 18160 18035
rect 18120 18000 18160 18005
rect 18200 18035 18240 18040
rect 18200 18005 18205 18035
rect 18235 18005 18240 18035
rect 18200 18000 18240 18005
rect 18280 18035 18320 18040
rect 18280 18005 18285 18035
rect 18315 18005 18320 18035
rect 18280 18000 18320 18005
rect 18360 18035 18400 18040
rect 18360 18005 18365 18035
rect 18395 18005 18400 18035
rect 18360 18000 18400 18005
rect 18440 18035 18480 18040
rect 18440 18005 18445 18035
rect 18475 18005 18480 18035
rect 18440 18000 18480 18005
rect 18520 18035 18560 18040
rect 18520 18005 18525 18035
rect 18555 18005 18560 18035
rect 18520 18000 18560 18005
rect 18600 18035 18640 18040
rect 18600 18005 18605 18035
rect 18635 18005 18640 18035
rect 18600 18000 18640 18005
rect 18680 18035 18720 18040
rect 18680 18005 18685 18035
rect 18715 18005 18720 18035
rect 18680 18000 18720 18005
rect 18760 18035 18800 18040
rect 18760 18005 18765 18035
rect 18795 18005 18800 18035
rect 18760 18000 18800 18005
rect 18840 18035 18880 18040
rect 18840 18005 18845 18035
rect 18875 18005 18880 18035
rect 18840 18000 18880 18005
rect 18920 18035 18960 18040
rect 18920 18005 18925 18035
rect 18955 18005 18960 18035
rect 18920 18000 18960 18005
rect 19000 18035 19040 18040
rect 19000 18005 19005 18035
rect 19035 18005 19040 18035
rect 19000 18000 19040 18005
rect 19080 18035 19120 18040
rect 19080 18005 19085 18035
rect 19115 18005 19120 18035
rect 19080 18000 19120 18005
rect 19160 18035 19200 18040
rect 19160 18005 19165 18035
rect 19195 18005 19200 18035
rect 19160 18000 19200 18005
rect 19240 18035 19280 18040
rect 19240 18005 19245 18035
rect 19275 18005 19280 18035
rect 19240 18000 19280 18005
rect 19320 18035 19360 18040
rect 19320 18005 19325 18035
rect 19355 18005 19360 18035
rect 19320 18000 19360 18005
rect 19400 18035 19440 18040
rect 19400 18005 19405 18035
rect 19435 18005 19440 18035
rect 19400 18000 19440 18005
rect 19480 18035 19520 18040
rect 19480 18005 19485 18035
rect 19515 18005 19520 18035
rect 19480 18000 19520 18005
rect 19560 18035 19600 18040
rect 19560 18005 19565 18035
rect 19595 18005 19600 18035
rect 19560 18000 19600 18005
rect 19640 18035 19680 18040
rect 19640 18005 19645 18035
rect 19675 18005 19680 18035
rect 19640 18000 19680 18005
rect 19720 18035 19760 18040
rect 19720 18005 19725 18035
rect 19755 18005 19760 18035
rect 19720 18000 19760 18005
rect 19800 18035 19840 18040
rect 19800 18005 19805 18035
rect 19835 18005 19840 18035
rect 19800 18000 19840 18005
rect 19880 18035 19920 18040
rect 19880 18005 19885 18035
rect 19915 18005 19920 18035
rect 19880 18000 19920 18005
rect 19960 18035 20000 18040
rect 19960 18005 19965 18035
rect 19995 18005 20000 18035
rect 19960 18000 20000 18005
rect 20040 18035 20080 18040
rect 20040 18005 20045 18035
rect 20075 18005 20080 18035
rect 20040 18000 20080 18005
rect 20120 18035 20160 18040
rect 20120 18005 20125 18035
rect 20155 18005 20160 18035
rect 20120 18000 20160 18005
rect 20200 18035 20240 18040
rect 20200 18005 20205 18035
rect 20235 18005 20240 18035
rect 20200 18000 20240 18005
rect 20280 18035 20320 18040
rect 20280 18005 20285 18035
rect 20315 18005 20320 18035
rect 20280 18000 20320 18005
rect 20360 18035 20400 18040
rect 20360 18005 20365 18035
rect 20395 18005 20400 18035
rect 20360 18000 20400 18005
rect 20440 18035 20480 18040
rect 20440 18005 20445 18035
rect 20475 18005 20480 18035
rect 20440 18000 20480 18005
rect 20520 18035 20560 18040
rect 20520 18005 20525 18035
rect 20555 18005 20560 18035
rect 20520 18000 20560 18005
rect 20600 18035 20640 18040
rect 20600 18005 20605 18035
rect 20635 18005 20640 18035
rect 20600 18000 20640 18005
rect 20680 18035 20720 18040
rect 20680 18005 20685 18035
rect 20715 18005 20720 18035
rect 20680 18000 20720 18005
rect 20760 18035 20800 18040
rect 20760 18005 20765 18035
rect 20795 18005 20800 18035
rect 20760 18000 20800 18005
rect 20840 18035 20880 18040
rect 20840 18005 20845 18035
rect 20875 18005 20880 18035
rect 20840 18000 20880 18005
rect 20920 18035 20960 18040
rect 20920 18005 20925 18035
rect 20955 18005 20960 18035
rect 20920 18000 20960 18005
rect 0 17875 40 17880
rect 0 17845 5 17875
rect 35 17845 40 17875
rect 0 17840 40 17845
rect 80 17875 120 17880
rect 80 17845 85 17875
rect 115 17845 120 17875
rect 80 17840 120 17845
rect 160 17875 200 17880
rect 160 17845 165 17875
rect 195 17845 200 17875
rect 160 17840 200 17845
rect 240 17875 280 17880
rect 240 17845 245 17875
rect 275 17845 280 17875
rect 240 17840 280 17845
rect 320 17875 360 17880
rect 320 17845 325 17875
rect 355 17845 360 17875
rect 320 17840 360 17845
rect 400 17875 440 17880
rect 400 17845 405 17875
rect 435 17845 440 17875
rect 400 17840 440 17845
rect 480 17875 520 17880
rect 480 17845 485 17875
rect 515 17845 520 17875
rect 480 17840 520 17845
rect 560 17875 600 17880
rect 560 17845 565 17875
rect 595 17845 600 17875
rect 560 17840 600 17845
rect 640 17875 680 17880
rect 640 17845 645 17875
rect 675 17845 680 17875
rect 640 17840 680 17845
rect 720 17875 760 17880
rect 720 17845 725 17875
rect 755 17845 760 17875
rect 720 17840 760 17845
rect 800 17875 840 17880
rect 800 17845 805 17875
rect 835 17845 840 17875
rect 800 17840 840 17845
rect 880 17875 920 17880
rect 880 17845 885 17875
rect 915 17845 920 17875
rect 880 17840 920 17845
rect 960 17875 1000 17880
rect 960 17845 965 17875
rect 995 17845 1000 17875
rect 960 17840 1000 17845
rect 1040 17875 1080 17880
rect 1040 17845 1045 17875
rect 1075 17845 1080 17875
rect 1040 17840 1080 17845
rect 1120 17875 1160 17880
rect 1120 17845 1125 17875
rect 1155 17845 1160 17875
rect 1120 17840 1160 17845
rect 1200 17875 1240 17880
rect 1200 17845 1205 17875
rect 1235 17845 1240 17875
rect 1200 17840 1240 17845
rect 1280 17875 1320 17880
rect 1280 17845 1285 17875
rect 1315 17845 1320 17875
rect 1280 17840 1320 17845
rect 1360 17875 1400 17880
rect 1360 17845 1365 17875
rect 1395 17845 1400 17875
rect 1360 17840 1400 17845
rect 1440 17875 1480 17880
rect 1440 17845 1445 17875
rect 1475 17845 1480 17875
rect 1440 17840 1480 17845
rect 1520 17875 1560 17880
rect 1520 17845 1525 17875
rect 1555 17845 1560 17875
rect 1520 17840 1560 17845
rect 1600 17875 1640 17880
rect 1600 17845 1605 17875
rect 1635 17845 1640 17875
rect 1600 17840 1640 17845
rect 1680 17875 1720 17880
rect 1680 17845 1685 17875
rect 1715 17845 1720 17875
rect 1680 17840 1720 17845
rect 1760 17875 1800 17880
rect 1760 17845 1765 17875
rect 1795 17845 1800 17875
rect 1760 17840 1800 17845
rect 1840 17875 1880 17880
rect 1840 17845 1845 17875
rect 1875 17845 1880 17875
rect 1840 17840 1880 17845
rect 1920 17875 1960 17880
rect 1920 17845 1925 17875
rect 1955 17845 1960 17875
rect 1920 17840 1960 17845
rect 2000 17875 2040 17880
rect 2000 17845 2005 17875
rect 2035 17845 2040 17875
rect 2000 17840 2040 17845
rect 2080 17875 2120 17880
rect 2080 17845 2085 17875
rect 2115 17845 2120 17875
rect 2080 17840 2120 17845
rect 2160 17875 2200 17880
rect 2160 17845 2165 17875
rect 2195 17845 2200 17875
rect 2160 17840 2200 17845
rect 2240 17875 2280 17880
rect 2240 17845 2245 17875
rect 2275 17845 2280 17875
rect 2240 17840 2280 17845
rect 2320 17875 2360 17880
rect 2320 17845 2325 17875
rect 2355 17845 2360 17875
rect 2320 17840 2360 17845
rect 2400 17875 2440 17880
rect 2400 17845 2405 17875
rect 2435 17845 2440 17875
rect 2400 17840 2440 17845
rect 2480 17875 2520 17880
rect 2480 17845 2485 17875
rect 2515 17845 2520 17875
rect 2480 17840 2520 17845
rect 2560 17875 2600 17880
rect 2560 17845 2565 17875
rect 2595 17845 2600 17875
rect 2560 17840 2600 17845
rect 2640 17875 2680 17880
rect 2640 17845 2645 17875
rect 2675 17845 2680 17875
rect 2640 17840 2680 17845
rect 2720 17875 2760 17880
rect 2720 17845 2725 17875
rect 2755 17845 2760 17875
rect 2720 17840 2760 17845
rect 2800 17875 2840 17880
rect 2800 17845 2805 17875
rect 2835 17845 2840 17875
rect 2800 17840 2840 17845
rect 2880 17875 2920 17880
rect 2880 17845 2885 17875
rect 2915 17845 2920 17875
rect 2880 17840 2920 17845
rect 2960 17875 3000 17880
rect 2960 17845 2965 17875
rect 2995 17845 3000 17875
rect 2960 17840 3000 17845
rect 3040 17875 3080 17880
rect 3040 17845 3045 17875
rect 3075 17845 3080 17875
rect 3040 17840 3080 17845
rect 3120 17875 3160 17880
rect 3120 17845 3125 17875
rect 3155 17845 3160 17875
rect 3120 17840 3160 17845
rect 3200 17875 3240 17880
rect 3200 17845 3205 17875
rect 3235 17845 3240 17875
rect 3200 17840 3240 17845
rect 3280 17875 3320 17880
rect 3280 17845 3285 17875
rect 3315 17845 3320 17875
rect 3280 17840 3320 17845
rect 3360 17875 3400 17880
rect 3360 17845 3365 17875
rect 3395 17845 3400 17875
rect 3360 17840 3400 17845
rect 3440 17875 3480 17880
rect 3440 17845 3445 17875
rect 3475 17845 3480 17875
rect 3440 17840 3480 17845
rect 3520 17875 3560 17880
rect 3520 17845 3525 17875
rect 3555 17845 3560 17875
rect 3520 17840 3560 17845
rect 3600 17875 3640 17880
rect 3600 17845 3605 17875
rect 3635 17845 3640 17875
rect 3600 17840 3640 17845
rect 3680 17875 3720 17880
rect 3680 17845 3685 17875
rect 3715 17845 3720 17875
rect 3680 17840 3720 17845
rect 3760 17875 3800 17880
rect 3760 17845 3765 17875
rect 3795 17845 3800 17875
rect 3760 17840 3800 17845
rect 3840 17875 3880 17880
rect 3840 17845 3845 17875
rect 3875 17845 3880 17875
rect 3840 17840 3880 17845
rect 3920 17875 3960 17880
rect 3920 17845 3925 17875
rect 3955 17845 3960 17875
rect 3920 17840 3960 17845
rect 4000 17875 4040 17880
rect 4000 17845 4005 17875
rect 4035 17845 4040 17875
rect 4000 17840 4040 17845
rect 4080 17875 4120 17880
rect 4080 17845 4085 17875
rect 4115 17845 4120 17875
rect 4080 17840 4120 17845
rect 4160 17875 4200 17880
rect 4160 17845 4165 17875
rect 4195 17845 4200 17875
rect 4160 17840 4200 17845
rect 6240 17875 6280 17880
rect 6240 17845 6245 17875
rect 6275 17845 6280 17875
rect 6240 17840 6280 17845
rect 6320 17875 6360 17880
rect 6320 17845 6325 17875
rect 6355 17845 6360 17875
rect 6320 17840 6360 17845
rect 6400 17875 6440 17880
rect 6400 17845 6405 17875
rect 6435 17845 6440 17875
rect 6400 17840 6440 17845
rect 6480 17875 6520 17880
rect 6480 17845 6485 17875
rect 6515 17845 6520 17875
rect 6480 17840 6520 17845
rect 6560 17875 6600 17880
rect 6560 17845 6565 17875
rect 6595 17845 6600 17875
rect 6560 17840 6600 17845
rect 6640 17875 6680 17880
rect 6640 17845 6645 17875
rect 6675 17845 6680 17875
rect 6640 17840 6680 17845
rect 6720 17875 6760 17880
rect 6720 17845 6725 17875
rect 6755 17845 6760 17875
rect 6720 17840 6760 17845
rect 6800 17875 6840 17880
rect 6800 17845 6805 17875
rect 6835 17845 6840 17875
rect 6800 17840 6840 17845
rect 6880 17875 6920 17880
rect 6880 17845 6885 17875
rect 6915 17845 6920 17875
rect 6880 17840 6920 17845
rect 6960 17875 7000 17880
rect 6960 17845 6965 17875
rect 6995 17845 7000 17875
rect 6960 17840 7000 17845
rect 7040 17875 7080 17880
rect 7040 17845 7045 17875
rect 7075 17845 7080 17875
rect 7040 17840 7080 17845
rect 7120 17875 7160 17880
rect 7120 17845 7125 17875
rect 7155 17845 7160 17875
rect 7120 17840 7160 17845
rect 7200 17875 7240 17880
rect 7200 17845 7205 17875
rect 7235 17845 7240 17875
rect 7200 17840 7240 17845
rect 7280 17875 7320 17880
rect 7280 17845 7285 17875
rect 7315 17845 7320 17875
rect 7280 17840 7320 17845
rect 7360 17875 7400 17880
rect 7360 17845 7365 17875
rect 7395 17845 7400 17875
rect 7360 17840 7400 17845
rect 7440 17875 7480 17880
rect 7440 17845 7445 17875
rect 7475 17845 7480 17875
rect 7440 17840 7480 17845
rect 7520 17875 7560 17880
rect 7520 17845 7525 17875
rect 7555 17845 7560 17875
rect 7520 17840 7560 17845
rect 7600 17875 7640 17880
rect 7600 17845 7605 17875
rect 7635 17845 7640 17875
rect 7600 17840 7640 17845
rect 7680 17875 7720 17880
rect 7680 17845 7685 17875
rect 7715 17845 7720 17875
rect 7680 17840 7720 17845
rect 7760 17875 7800 17880
rect 7760 17845 7765 17875
rect 7795 17845 7800 17875
rect 7760 17840 7800 17845
rect 7840 17875 7880 17880
rect 7840 17845 7845 17875
rect 7875 17845 7880 17875
rect 7840 17840 7880 17845
rect 7920 17875 7960 17880
rect 7920 17845 7925 17875
rect 7955 17845 7960 17875
rect 7920 17840 7960 17845
rect 8000 17875 8040 17880
rect 8000 17845 8005 17875
rect 8035 17845 8040 17875
rect 8000 17840 8040 17845
rect 8080 17875 8120 17880
rect 8080 17845 8085 17875
rect 8115 17845 8120 17875
rect 8080 17840 8120 17845
rect 8160 17875 8200 17880
rect 8160 17845 8165 17875
rect 8195 17845 8200 17875
rect 8160 17840 8200 17845
rect 8240 17875 8280 17880
rect 8240 17845 8245 17875
rect 8275 17845 8280 17875
rect 8240 17840 8280 17845
rect 8320 17875 8360 17880
rect 8320 17845 8325 17875
rect 8355 17845 8360 17875
rect 8320 17840 8360 17845
rect 8400 17875 8440 17880
rect 8400 17845 8405 17875
rect 8435 17845 8440 17875
rect 8400 17840 8440 17845
rect 8480 17875 8520 17880
rect 8480 17845 8485 17875
rect 8515 17845 8520 17875
rect 8480 17840 8520 17845
rect 8560 17875 8600 17880
rect 8560 17845 8565 17875
rect 8595 17845 8600 17875
rect 8560 17840 8600 17845
rect 8640 17875 8680 17880
rect 8640 17845 8645 17875
rect 8675 17845 8680 17875
rect 8640 17840 8680 17845
rect 8720 17875 8760 17880
rect 8720 17845 8725 17875
rect 8755 17845 8760 17875
rect 8720 17840 8760 17845
rect 8800 17875 8840 17880
rect 8800 17845 8805 17875
rect 8835 17845 8840 17875
rect 8800 17840 8840 17845
rect 8880 17875 8920 17880
rect 8880 17845 8885 17875
rect 8915 17845 8920 17875
rect 8880 17840 8920 17845
rect 8960 17875 9000 17880
rect 8960 17845 8965 17875
rect 8995 17845 9000 17875
rect 8960 17840 9000 17845
rect 9040 17875 9080 17880
rect 9040 17845 9045 17875
rect 9075 17845 9080 17875
rect 9040 17840 9080 17845
rect 9120 17875 9160 17880
rect 9120 17845 9125 17875
rect 9155 17845 9160 17875
rect 9120 17840 9160 17845
rect 9200 17875 9240 17880
rect 9200 17845 9205 17875
rect 9235 17845 9240 17875
rect 9200 17840 9240 17845
rect 9280 17875 9320 17880
rect 9280 17845 9285 17875
rect 9315 17845 9320 17875
rect 9280 17840 9320 17845
rect 9360 17875 9400 17880
rect 9360 17845 9365 17875
rect 9395 17845 9400 17875
rect 9360 17840 9400 17845
rect 9440 17875 9480 17880
rect 9440 17845 9445 17875
rect 9475 17845 9480 17875
rect 9440 17840 9480 17845
rect 11560 17875 11600 17880
rect 11560 17845 11565 17875
rect 11595 17845 11600 17875
rect 11560 17840 11600 17845
rect 11640 17875 11680 17880
rect 11640 17845 11645 17875
rect 11675 17845 11680 17875
rect 11640 17840 11680 17845
rect 11720 17875 11760 17880
rect 11720 17845 11725 17875
rect 11755 17845 11760 17875
rect 11720 17840 11760 17845
rect 11800 17875 11840 17880
rect 11800 17845 11805 17875
rect 11835 17845 11840 17875
rect 11800 17840 11840 17845
rect 11880 17875 11920 17880
rect 11880 17845 11885 17875
rect 11915 17845 11920 17875
rect 11880 17840 11920 17845
rect 11960 17875 12000 17880
rect 11960 17845 11965 17875
rect 11995 17845 12000 17875
rect 11960 17840 12000 17845
rect 12040 17875 12080 17880
rect 12040 17845 12045 17875
rect 12075 17845 12080 17875
rect 12040 17840 12080 17845
rect 12120 17875 12160 17880
rect 12120 17845 12125 17875
rect 12155 17845 12160 17875
rect 12120 17840 12160 17845
rect 12200 17875 12240 17880
rect 12200 17845 12205 17875
rect 12235 17845 12240 17875
rect 12200 17840 12240 17845
rect 12280 17875 12320 17880
rect 12280 17845 12285 17875
rect 12315 17845 12320 17875
rect 12280 17840 12320 17845
rect 12360 17875 12400 17880
rect 12360 17845 12365 17875
rect 12395 17845 12400 17875
rect 12360 17840 12400 17845
rect 12440 17875 12480 17880
rect 12440 17845 12445 17875
rect 12475 17845 12480 17875
rect 12440 17840 12480 17845
rect 12520 17875 12560 17880
rect 12520 17845 12525 17875
rect 12555 17845 12560 17875
rect 12520 17840 12560 17845
rect 12600 17875 12640 17880
rect 12600 17845 12605 17875
rect 12635 17845 12640 17875
rect 12600 17840 12640 17845
rect 12680 17875 12720 17880
rect 12680 17845 12685 17875
rect 12715 17845 12720 17875
rect 12680 17840 12720 17845
rect 12760 17875 12800 17880
rect 12760 17845 12765 17875
rect 12795 17845 12800 17875
rect 12760 17840 12800 17845
rect 12840 17875 12880 17880
rect 12840 17845 12845 17875
rect 12875 17845 12880 17875
rect 12840 17840 12880 17845
rect 12920 17875 12960 17880
rect 12920 17845 12925 17875
rect 12955 17845 12960 17875
rect 12920 17840 12960 17845
rect 13000 17875 13040 17880
rect 13000 17845 13005 17875
rect 13035 17845 13040 17875
rect 13000 17840 13040 17845
rect 13080 17875 13120 17880
rect 13080 17845 13085 17875
rect 13115 17845 13120 17875
rect 13080 17840 13120 17845
rect 13160 17875 13200 17880
rect 13160 17845 13165 17875
rect 13195 17845 13200 17875
rect 13160 17840 13200 17845
rect 13240 17875 13280 17880
rect 13240 17845 13245 17875
rect 13275 17845 13280 17875
rect 13240 17840 13280 17845
rect 13320 17875 13360 17880
rect 13320 17845 13325 17875
rect 13355 17845 13360 17875
rect 13320 17840 13360 17845
rect 13400 17875 13440 17880
rect 13400 17845 13405 17875
rect 13435 17845 13440 17875
rect 13400 17840 13440 17845
rect 13480 17875 13520 17880
rect 13480 17845 13485 17875
rect 13515 17845 13520 17875
rect 13480 17840 13520 17845
rect 13560 17875 13600 17880
rect 13560 17845 13565 17875
rect 13595 17845 13600 17875
rect 13560 17840 13600 17845
rect 13640 17875 13680 17880
rect 13640 17845 13645 17875
rect 13675 17845 13680 17875
rect 13640 17840 13680 17845
rect 13720 17875 13760 17880
rect 13720 17845 13725 17875
rect 13755 17845 13760 17875
rect 13720 17840 13760 17845
rect 13800 17875 13840 17880
rect 13800 17845 13805 17875
rect 13835 17845 13840 17875
rect 13800 17840 13840 17845
rect 13880 17875 13920 17880
rect 13880 17845 13885 17875
rect 13915 17845 13920 17875
rect 13880 17840 13920 17845
rect 13960 17875 14000 17880
rect 13960 17845 13965 17875
rect 13995 17845 14000 17875
rect 13960 17840 14000 17845
rect 14040 17875 14080 17880
rect 14040 17845 14045 17875
rect 14075 17845 14080 17875
rect 14040 17840 14080 17845
rect 14120 17875 14160 17880
rect 14120 17845 14125 17875
rect 14155 17845 14160 17875
rect 14120 17840 14160 17845
rect 14200 17875 14240 17880
rect 14200 17845 14205 17875
rect 14235 17845 14240 17875
rect 14200 17840 14240 17845
rect 14280 17875 14320 17880
rect 14280 17845 14285 17875
rect 14315 17845 14320 17875
rect 14280 17840 14320 17845
rect 14360 17875 14400 17880
rect 14360 17845 14365 17875
rect 14395 17845 14400 17875
rect 14360 17840 14400 17845
rect 14440 17875 14480 17880
rect 14440 17845 14445 17875
rect 14475 17845 14480 17875
rect 14440 17840 14480 17845
rect 14520 17875 14560 17880
rect 14520 17845 14525 17875
rect 14555 17845 14560 17875
rect 14520 17840 14560 17845
rect 14600 17875 14640 17880
rect 14600 17845 14605 17875
rect 14635 17845 14640 17875
rect 14600 17840 14640 17845
rect 14680 17875 14720 17880
rect 14680 17845 14685 17875
rect 14715 17845 14720 17875
rect 14680 17840 14720 17845
rect 16760 17875 16800 17880
rect 16760 17845 16765 17875
rect 16795 17845 16800 17875
rect 16760 17840 16800 17845
rect 16840 17875 16880 17880
rect 16840 17845 16845 17875
rect 16875 17845 16880 17875
rect 16840 17840 16880 17845
rect 16920 17875 16960 17880
rect 16920 17845 16925 17875
rect 16955 17845 16960 17875
rect 16920 17840 16960 17845
rect 17000 17875 17040 17880
rect 17000 17845 17005 17875
rect 17035 17845 17040 17875
rect 17000 17840 17040 17845
rect 17080 17875 17120 17880
rect 17080 17845 17085 17875
rect 17115 17845 17120 17875
rect 17080 17840 17120 17845
rect 17160 17875 17200 17880
rect 17160 17845 17165 17875
rect 17195 17845 17200 17875
rect 17160 17840 17200 17845
rect 17240 17875 17280 17880
rect 17240 17845 17245 17875
rect 17275 17845 17280 17875
rect 17240 17840 17280 17845
rect 17320 17875 17360 17880
rect 17320 17845 17325 17875
rect 17355 17845 17360 17875
rect 17320 17840 17360 17845
rect 17400 17875 17440 17880
rect 17400 17845 17405 17875
rect 17435 17845 17440 17875
rect 17400 17840 17440 17845
rect 17480 17875 17520 17880
rect 17480 17845 17485 17875
rect 17515 17845 17520 17875
rect 17480 17840 17520 17845
rect 17560 17875 17600 17880
rect 17560 17845 17565 17875
rect 17595 17845 17600 17875
rect 17560 17840 17600 17845
rect 17640 17875 17680 17880
rect 17640 17845 17645 17875
rect 17675 17845 17680 17875
rect 17640 17840 17680 17845
rect 17720 17875 17760 17880
rect 17720 17845 17725 17875
rect 17755 17845 17760 17875
rect 17720 17840 17760 17845
rect 17800 17875 17840 17880
rect 17800 17845 17805 17875
rect 17835 17845 17840 17875
rect 17800 17840 17840 17845
rect 17880 17875 17920 17880
rect 17880 17845 17885 17875
rect 17915 17845 17920 17875
rect 17880 17840 17920 17845
rect 17960 17875 18000 17880
rect 17960 17845 17965 17875
rect 17995 17845 18000 17875
rect 17960 17840 18000 17845
rect 18040 17875 18080 17880
rect 18040 17845 18045 17875
rect 18075 17845 18080 17875
rect 18040 17840 18080 17845
rect 18120 17875 18160 17880
rect 18120 17845 18125 17875
rect 18155 17845 18160 17875
rect 18120 17840 18160 17845
rect 18200 17875 18240 17880
rect 18200 17845 18205 17875
rect 18235 17845 18240 17875
rect 18200 17840 18240 17845
rect 18280 17875 18320 17880
rect 18280 17845 18285 17875
rect 18315 17845 18320 17875
rect 18280 17840 18320 17845
rect 18360 17875 18400 17880
rect 18360 17845 18365 17875
rect 18395 17845 18400 17875
rect 18360 17840 18400 17845
rect 18440 17875 18480 17880
rect 18440 17845 18445 17875
rect 18475 17845 18480 17875
rect 18440 17840 18480 17845
rect 18520 17875 18560 17880
rect 18520 17845 18525 17875
rect 18555 17845 18560 17875
rect 18520 17840 18560 17845
rect 18600 17875 18640 17880
rect 18600 17845 18605 17875
rect 18635 17845 18640 17875
rect 18600 17840 18640 17845
rect 18680 17875 18720 17880
rect 18680 17845 18685 17875
rect 18715 17845 18720 17875
rect 18680 17840 18720 17845
rect 18760 17875 18800 17880
rect 18760 17845 18765 17875
rect 18795 17845 18800 17875
rect 18760 17840 18800 17845
rect 18840 17875 18880 17880
rect 18840 17845 18845 17875
rect 18875 17845 18880 17875
rect 18840 17840 18880 17845
rect 18920 17875 18960 17880
rect 18920 17845 18925 17875
rect 18955 17845 18960 17875
rect 18920 17840 18960 17845
rect 19000 17875 19040 17880
rect 19000 17845 19005 17875
rect 19035 17845 19040 17875
rect 19000 17840 19040 17845
rect 19080 17875 19120 17880
rect 19080 17845 19085 17875
rect 19115 17845 19120 17875
rect 19080 17840 19120 17845
rect 19160 17875 19200 17880
rect 19160 17845 19165 17875
rect 19195 17845 19200 17875
rect 19160 17840 19200 17845
rect 19240 17875 19280 17880
rect 19240 17845 19245 17875
rect 19275 17845 19280 17875
rect 19240 17840 19280 17845
rect 19320 17875 19360 17880
rect 19320 17845 19325 17875
rect 19355 17845 19360 17875
rect 19320 17840 19360 17845
rect 19400 17875 19440 17880
rect 19400 17845 19405 17875
rect 19435 17845 19440 17875
rect 19400 17840 19440 17845
rect 19480 17875 19520 17880
rect 19480 17845 19485 17875
rect 19515 17845 19520 17875
rect 19480 17840 19520 17845
rect 19560 17875 19600 17880
rect 19560 17845 19565 17875
rect 19595 17845 19600 17875
rect 19560 17840 19600 17845
rect 19640 17875 19680 17880
rect 19640 17845 19645 17875
rect 19675 17845 19680 17875
rect 19640 17840 19680 17845
rect 19720 17875 19760 17880
rect 19720 17845 19725 17875
rect 19755 17845 19760 17875
rect 19720 17840 19760 17845
rect 19800 17875 19840 17880
rect 19800 17845 19805 17875
rect 19835 17845 19840 17875
rect 19800 17840 19840 17845
rect 19880 17875 19920 17880
rect 19880 17845 19885 17875
rect 19915 17845 19920 17875
rect 19880 17840 19920 17845
rect 19960 17875 20000 17880
rect 19960 17845 19965 17875
rect 19995 17845 20000 17875
rect 19960 17840 20000 17845
rect 20040 17875 20080 17880
rect 20040 17845 20045 17875
rect 20075 17845 20080 17875
rect 20040 17840 20080 17845
rect 20120 17875 20160 17880
rect 20120 17845 20125 17875
rect 20155 17845 20160 17875
rect 20120 17840 20160 17845
rect 20200 17875 20240 17880
rect 20200 17845 20205 17875
rect 20235 17845 20240 17875
rect 20200 17840 20240 17845
rect 20280 17875 20320 17880
rect 20280 17845 20285 17875
rect 20315 17845 20320 17875
rect 20280 17840 20320 17845
rect 20360 17875 20400 17880
rect 20360 17845 20365 17875
rect 20395 17845 20400 17875
rect 20360 17840 20400 17845
rect 20440 17875 20480 17880
rect 20440 17845 20445 17875
rect 20475 17845 20480 17875
rect 20440 17840 20480 17845
rect 20520 17875 20560 17880
rect 20520 17845 20525 17875
rect 20555 17845 20560 17875
rect 20520 17840 20560 17845
rect 20600 17875 20640 17880
rect 20600 17845 20605 17875
rect 20635 17845 20640 17875
rect 20600 17840 20640 17845
rect 20680 17875 20720 17880
rect 20680 17845 20685 17875
rect 20715 17845 20720 17875
rect 20680 17840 20720 17845
rect 20760 17875 20800 17880
rect 20760 17845 20765 17875
rect 20795 17845 20800 17875
rect 20760 17840 20800 17845
rect 20840 17875 20880 17880
rect 20840 17845 20845 17875
rect 20875 17845 20880 17875
rect 20840 17840 20880 17845
rect 20920 17875 20960 17880
rect 20920 17845 20925 17875
rect 20955 17845 20960 17875
rect 20920 17840 20960 17845
rect 0 17715 40 17720
rect 0 17685 5 17715
rect 35 17685 40 17715
rect 0 17680 40 17685
rect 80 17715 120 17720
rect 80 17685 85 17715
rect 115 17685 120 17715
rect 80 17680 120 17685
rect 160 17715 200 17720
rect 160 17685 165 17715
rect 195 17685 200 17715
rect 160 17680 200 17685
rect 240 17715 280 17720
rect 240 17685 245 17715
rect 275 17685 280 17715
rect 240 17680 280 17685
rect 320 17715 360 17720
rect 320 17685 325 17715
rect 355 17685 360 17715
rect 320 17680 360 17685
rect 400 17715 440 17720
rect 400 17685 405 17715
rect 435 17685 440 17715
rect 400 17680 440 17685
rect 480 17715 520 17720
rect 480 17685 485 17715
rect 515 17685 520 17715
rect 480 17680 520 17685
rect 560 17715 600 17720
rect 560 17685 565 17715
rect 595 17685 600 17715
rect 560 17680 600 17685
rect 640 17715 680 17720
rect 640 17685 645 17715
rect 675 17685 680 17715
rect 640 17680 680 17685
rect 720 17715 760 17720
rect 720 17685 725 17715
rect 755 17685 760 17715
rect 720 17680 760 17685
rect 800 17715 840 17720
rect 800 17685 805 17715
rect 835 17685 840 17715
rect 800 17680 840 17685
rect 880 17715 920 17720
rect 880 17685 885 17715
rect 915 17685 920 17715
rect 880 17680 920 17685
rect 960 17715 1000 17720
rect 960 17685 965 17715
rect 995 17685 1000 17715
rect 960 17680 1000 17685
rect 1040 17715 1080 17720
rect 1040 17685 1045 17715
rect 1075 17685 1080 17715
rect 1040 17680 1080 17685
rect 1120 17715 1160 17720
rect 1120 17685 1125 17715
rect 1155 17685 1160 17715
rect 1120 17680 1160 17685
rect 1200 17715 1240 17720
rect 1200 17685 1205 17715
rect 1235 17685 1240 17715
rect 1200 17680 1240 17685
rect 1280 17715 1320 17720
rect 1280 17685 1285 17715
rect 1315 17685 1320 17715
rect 1280 17680 1320 17685
rect 1360 17715 1400 17720
rect 1360 17685 1365 17715
rect 1395 17685 1400 17715
rect 1360 17680 1400 17685
rect 1440 17715 1480 17720
rect 1440 17685 1445 17715
rect 1475 17685 1480 17715
rect 1440 17680 1480 17685
rect 1520 17715 1560 17720
rect 1520 17685 1525 17715
rect 1555 17685 1560 17715
rect 1520 17680 1560 17685
rect 1600 17715 1640 17720
rect 1600 17685 1605 17715
rect 1635 17685 1640 17715
rect 1600 17680 1640 17685
rect 1680 17715 1720 17720
rect 1680 17685 1685 17715
rect 1715 17685 1720 17715
rect 1680 17680 1720 17685
rect 1760 17715 1800 17720
rect 1760 17685 1765 17715
rect 1795 17685 1800 17715
rect 1760 17680 1800 17685
rect 1840 17715 1880 17720
rect 1840 17685 1845 17715
rect 1875 17685 1880 17715
rect 1840 17680 1880 17685
rect 1920 17715 1960 17720
rect 1920 17685 1925 17715
rect 1955 17685 1960 17715
rect 1920 17680 1960 17685
rect 2000 17715 2040 17720
rect 2000 17685 2005 17715
rect 2035 17685 2040 17715
rect 2000 17680 2040 17685
rect 2080 17715 2120 17720
rect 2080 17685 2085 17715
rect 2115 17685 2120 17715
rect 2080 17680 2120 17685
rect 2160 17715 2200 17720
rect 2160 17685 2165 17715
rect 2195 17685 2200 17715
rect 2160 17680 2200 17685
rect 2240 17715 2280 17720
rect 2240 17685 2245 17715
rect 2275 17685 2280 17715
rect 2240 17680 2280 17685
rect 2320 17715 2360 17720
rect 2320 17685 2325 17715
rect 2355 17685 2360 17715
rect 2320 17680 2360 17685
rect 2400 17715 2440 17720
rect 2400 17685 2405 17715
rect 2435 17685 2440 17715
rect 2400 17680 2440 17685
rect 2480 17715 2520 17720
rect 2480 17685 2485 17715
rect 2515 17685 2520 17715
rect 2480 17680 2520 17685
rect 2560 17715 2600 17720
rect 2560 17685 2565 17715
rect 2595 17685 2600 17715
rect 2560 17680 2600 17685
rect 2640 17715 2680 17720
rect 2640 17685 2645 17715
rect 2675 17685 2680 17715
rect 2640 17680 2680 17685
rect 2720 17715 2760 17720
rect 2720 17685 2725 17715
rect 2755 17685 2760 17715
rect 2720 17680 2760 17685
rect 2800 17715 2840 17720
rect 2800 17685 2805 17715
rect 2835 17685 2840 17715
rect 2800 17680 2840 17685
rect 2880 17715 2920 17720
rect 2880 17685 2885 17715
rect 2915 17685 2920 17715
rect 2880 17680 2920 17685
rect 2960 17715 3000 17720
rect 2960 17685 2965 17715
rect 2995 17685 3000 17715
rect 2960 17680 3000 17685
rect 3040 17715 3080 17720
rect 3040 17685 3045 17715
rect 3075 17685 3080 17715
rect 3040 17680 3080 17685
rect 3120 17715 3160 17720
rect 3120 17685 3125 17715
rect 3155 17685 3160 17715
rect 3120 17680 3160 17685
rect 3200 17715 3240 17720
rect 3200 17685 3205 17715
rect 3235 17685 3240 17715
rect 3200 17680 3240 17685
rect 3280 17715 3320 17720
rect 3280 17685 3285 17715
rect 3315 17685 3320 17715
rect 3280 17680 3320 17685
rect 3360 17715 3400 17720
rect 3360 17685 3365 17715
rect 3395 17685 3400 17715
rect 3360 17680 3400 17685
rect 3440 17715 3480 17720
rect 3440 17685 3445 17715
rect 3475 17685 3480 17715
rect 3440 17680 3480 17685
rect 3520 17715 3560 17720
rect 3520 17685 3525 17715
rect 3555 17685 3560 17715
rect 3520 17680 3560 17685
rect 3600 17715 3640 17720
rect 3600 17685 3605 17715
rect 3635 17685 3640 17715
rect 3600 17680 3640 17685
rect 3680 17715 3720 17720
rect 3680 17685 3685 17715
rect 3715 17685 3720 17715
rect 3680 17680 3720 17685
rect 3760 17715 3800 17720
rect 3760 17685 3765 17715
rect 3795 17685 3800 17715
rect 3760 17680 3800 17685
rect 3840 17715 3880 17720
rect 3840 17685 3845 17715
rect 3875 17685 3880 17715
rect 3840 17680 3880 17685
rect 3920 17715 3960 17720
rect 3920 17685 3925 17715
rect 3955 17685 3960 17715
rect 3920 17680 3960 17685
rect 4000 17715 4040 17720
rect 4000 17685 4005 17715
rect 4035 17685 4040 17715
rect 4000 17680 4040 17685
rect 4080 17715 4120 17720
rect 4080 17685 4085 17715
rect 4115 17685 4120 17715
rect 4080 17680 4120 17685
rect 4160 17715 4200 17720
rect 4160 17685 4165 17715
rect 4195 17685 4200 17715
rect 4160 17680 4200 17685
rect 6240 17715 6280 17720
rect 6240 17685 6245 17715
rect 6275 17685 6280 17715
rect 6240 17680 6280 17685
rect 6320 17715 6360 17720
rect 6320 17685 6325 17715
rect 6355 17685 6360 17715
rect 6320 17680 6360 17685
rect 6400 17715 6440 17720
rect 6400 17685 6405 17715
rect 6435 17685 6440 17715
rect 6400 17680 6440 17685
rect 6480 17715 6520 17720
rect 6480 17685 6485 17715
rect 6515 17685 6520 17715
rect 6480 17680 6520 17685
rect 6560 17715 6600 17720
rect 6560 17685 6565 17715
rect 6595 17685 6600 17715
rect 6560 17680 6600 17685
rect 6640 17715 6680 17720
rect 6640 17685 6645 17715
rect 6675 17685 6680 17715
rect 6640 17680 6680 17685
rect 6720 17715 6760 17720
rect 6720 17685 6725 17715
rect 6755 17685 6760 17715
rect 6720 17680 6760 17685
rect 6800 17715 6840 17720
rect 6800 17685 6805 17715
rect 6835 17685 6840 17715
rect 6800 17680 6840 17685
rect 6880 17715 6920 17720
rect 6880 17685 6885 17715
rect 6915 17685 6920 17715
rect 6880 17680 6920 17685
rect 6960 17715 7000 17720
rect 6960 17685 6965 17715
rect 6995 17685 7000 17715
rect 6960 17680 7000 17685
rect 7040 17715 7080 17720
rect 7040 17685 7045 17715
rect 7075 17685 7080 17715
rect 7040 17680 7080 17685
rect 7120 17715 7160 17720
rect 7120 17685 7125 17715
rect 7155 17685 7160 17715
rect 7120 17680 7160 17685
rect 7200 17715 7240 17720
rect 7200 17685 7205 17715
rect 7235 17685 7240 17715
rect 7200 17680 7240 17685
rect 7280 17715 7320 17720
rect 7280 17685 7285 17715
rect 7315 17685 7320 17715
rect 7280 17680 7320 17685
rect 7360 17715 7400 17720
rect 7360 17685 7365 17715
rect 7395 17685 7400 17715
rect 7360 17680 7400 17685
rect 7440 17715 7480 17720
rect 7440 17685 7445 17715
rect 7475 17685 7480 17715
rect 7440 17680 7480 17685
rect 7520 17715 7560 17720
rect 7520 17685 7525 17715
rect 7555 17685 7560 17715
rect 7520 17680 7560 17685
rect 7600 17715 7640 17720
rect 7600 17685 7605 17715
rect 7635 17685 7640 17715
rect 7600 17680 7640 17685
rect 7680 17715 7720 17720
rect 7680 17685 7685 17715
rect 7715 17685 7720 17715
rect 7680 17680 7720 17685
rect 7760 17715 7800 17720
rect 7760 17685 7765 17715
rect 7795 17685 7800 17715
rect 7760 17680 7800 17685
rect 7840 17715 7880 17720
rect 7840 17685 7845 17715
rect 7875 17685 7880 17715
rect 7840 17680 7880 17685
rect 7920 17715 7960 17720
rect 7920 17685 7925 17715
rect 7955 17685 7960 17715
rect 7920 17680 7960 17685
rect 8000 17715 8040 17720
rect 8000 17685 8005 17715
rect 8035 17685 8040 17715
rect 8000 17680 8040 17685
rect 8080 17715 8120 17720
rect 8080 17685 8085 17715
rect 8115 17685 8120 17715
rect 8080 17680 8120 17685
rect 8160 17715 8200 17720
rect 8160 17685 8165 17715
rect 8195 17685 8200 17715
rect 8160 17680 8200 17685
rect 8240 17715 8280 17720
rect 8240 17685 8245 17715
rect 8275 17685 8280 17715
rect 8240 17680 8280 17685
rect 8320 17715 8360 17720
rect 8320 17685 8325 17715
rect 8355 17685 8360 17715
rect 8320 17680 8360 17685
rect 8400 17715 8440 17720
rect 8400 17685 8405 17715
rect 8435 17685 8440 17715
rect 8400 17680 8440 17685
rect 8480 17715 8520 17720
rect 8480 17685 8485 17715
rect 8515 17685 8520 17715
rect 8480 17680 8520 17685
rect 8560 17715 8600 17720
rect 8560 17685 8565 17715
rect 8595 17685 8600 17715
rect 8560 17680 8600 17685
rect 8640 17715 8680 17720
rect 8640 17685 8645 17715
rect 8675 17685 8680 17715
rect 8640 17680 8680 17685
rect 8720 17715 8760 17720
rect 8720 17685 8725 17715
rect 8755 17685 8760 17715
rect 8720 17680 8760 17685
rect 8800 17715 8840 17720
rect 8800 17685 8805 17715
rect 8835 17685 8840 17715
rect 8800 17680 8840 17685
rect 8880 17715 8920 17720
rect 8880 17685 8885 17715
rect 8915 17685 8920 17715
rect 8880 17680 8920 17685
rect 8960 17715 9000 17720
rect 8960 17685 8965 17715
rect 8995 17685 9000 17715
rect 8960 17680 9000 17685
rect 9040 17715 9080 17720
rect 9040 17685 9045 17715
rect 9075 17685 9080 17715
rect 9040 17680 9080 17685
rect 9120 17715 9160 17720
rect 9120 17685 9125 17715
rect 9155 17685 9160 17715
rect 9120 17680 9160 17685
rect 9200 17715 9240 17720
rect 9200 17685 9205 17715
rect 9235 17685 9240 17715
rect 9200 17680 9240 17685
rect 9280 17715 9320 17720
rect 9280 17685 9285 17715
rect 9315 17685 9320 17715
rect 9280 17680 9320 17685
rect 9360 17715 9400 17720
rect 9360 17685 9365 17715
rect 9395 17685 9400 17715
rect 9360 17680 9400 17685
rect 9440 17715 9480 17720
rect 9440 17685 9445 17715
rect 9475 17685 9480 17715
rect 9440 17680 9480 17685
rect 11560 17715 11600 17720
rect 11560 17685 11565 17715
rect 11595 17685 11600 17715
rect 11560 17680 11600 17685
rect 11640 17715 11680 17720
rect 11640 17685 11645 17715
rect 11675 17685 11680 17715
rect 11640 17680 11680 17685
rect 11720 17715 11760 17720
rect 11720 17685 11725 17715
rect 11755 17685 11760 17715
rect 11720 17680 11760 17685
rect 11800 17715 11840 17720
rect 11800 17685 11805 17715
rect 11835 17685 11840 17715
rect 11800 17680 11840 17685
rect 11880 17715 11920 17720
rect 11880 17685 11885 17715
rect 11915 17685 11920 17715
rect 11880 17680 11920 17685
rect 11960 17715 12000 17720
rect 11960 17685 11965 17715
rect 11995 17685 12000 17715
rect 11960 17680 12000 17685
rect 12040 17715 12080 17720
rect 12040 17685 12045 17715
rect 12075 17685 12080 17715
rect 12040 17680 12080 17685
rect 12120 17715 12160 17720
rect 12120 17685 12125 17715
rect 12155 17685 12160 17715
rect 12120 17680 12160 17685
rect 12200 17715 12240 17720
rect 12200 17685 12205 17715
rect 12235 17685 12240 17715
rect 12200 17680 12240 17685
rect 12280 17715 12320 17720
rect 12280 17685 12285 17715
rect 12315 17685 12320 17715
rect 12280 17680 12320 17685
rect 12360 17715 12400 17720
rect 12360 17685 12365 17715
rect 12395 17685 12400 17715
rect 12360 17680 12400 17685
rect 12440 17715 12480 17720
rect 12440 17685 12445 17715
rect 12475 17685 12480 17715
rect 12440 17680 12480 17685
rect 12520 17715 12560 17720
rect 12520 17685 12525 17715
rect 12555 17685 12560 17715
rect 12520 17680 12560 17685
rect 12600 17715 12640 17720
rect 12600 17685 12605 17715
rect 12635 17685 12640 17715
rect 12600 17680 12640 17685
rect 12680 17715 12720 17720
rect 12680 17685 12685 17715
rect 12715 17685 12720 17715
rect 12680 17680 12720 17685
rect 12760 17715 12800 17720
rect 12760 17685 12765 17715
rect 12795 17685 12800 17715
rect 12760 17680 12800 17685
rect 12840 17715 12880 17720
rect 12840 17685 12845 17715
rect 12875 17685 12880 17715
rect 12840 17680 12880 17685
rect 12920 17715 12960 17720
rect 12920 17685 12925 17715
rect 12955 17685 12960 17715
rect 12920 17680 12960 17685
rect 13000 17715 13040 17720
rect 13000 17685 13005 17715
rect 13035 17685 13040 17715
rect 13000 17680 13040 17685
rect 13080 17715 13120 17720
rect 13080 17685 13085 17715
rect 13115 17685 13120 17715
rect 13080 17680 13120 17685
rect 13160 17715 13200 17720
rect 13160 17685 13165 17715
rect 13195 17685 13200 17715
rect 13160 17680 13200 17685
rect 13240 17715 13280 17720
rect 13240 17685 13245 17715
rect 13275 17685 13280 17715
rect 13240 17680 13280 17685
rect 13320 17715 13360 17720
rect 13320 17685 13325 17715
rect 13355 17685 13360 17715
rect 13320 17680 13360 17685
rect 13400 17715 13440 17720
rect 13400 17685 13405 17715
rect 13435 17685 13440 17715
rect 13400 17680 13440 17685
rect 13480 17715 13520 17720
rect 13480 17685 13485 17715
rect 13515 17685 13520 17715
rect 13480 17680 13520 17685
rect 13560 17715 13600 17720
rect 13560 17685 13565 17715
rect 13595 17685 13600 17715
rect 13560 17680 13600 17685
rect 13640 17715 13680 17720
rect 13640 17685 13645 17715
rect 13675 17685 13680 17715
rect 13640 17680 13680 17685
rect 13720 17715 13760 17720
rect 13720 17685 13725 17715
rect 13755 17685 13760 17715
rect 13720 17680 13760 17685
rect 13800 17715 13840 17720
rect 13800 17685 13805 17715
rect 13835 17685 13840 17715
rect 13800 17680 13840 17685
rect 13880 17715 13920 17720
rect 13880 17685 13885 17715
rect 13915 17685 13920 17715
rect 13880 17680 13920 17685
rect 13960 17715 14000 17720
rect 13960 17685 13965 17715
rect 13995 17685 14000 17715
rect 13960 17680 14000 17685
rect 14040 17715 14080 17720
rect 14040 17685 14045 17715
rect 14075 17685 14080 17715
rect 14040 17680 14080 17685
rect 14120 17715 14160 17720
rect 14120 17685 14125 17715
rect 14155 17685 14160 17715
rect 14120 17680 14160 17685
rect 14200 17715 14240 17720
rect 14200 17685 14205 17715
rect 14235 17685 14240 17715
rect 14200 17680 14240 17685
rect 14280 17715 14320 17720
rect 14280 17685 14285 17715
rect 14315 17685 14320 17715
rect 14280 17680 14320 17685
rect 14360 17715 14400 17720
rect 14360 17685 14365 17715
rect 14395 17685 14400 17715
rect 14360 17680 14400 17685
rect 14440 17715 14480 17720
rect 14440 17685 14445 17715
rect 14475 17685 14480 17715
rect 14440 17680 14480 17685
rect 14520 17715 14560 17720
rect 14520 17685 14525 17715
rect 14555 17685 14560 17715
rect 14520 17680 14560 17685
rect 14600 17715 14640 17720
rect 14600 17685 14605 17715
rect 14635 17685 14640 17715
rect 14600 17680 14640 17685
rect 14680 17715 14720 17720
rect 14680 17685 14685 17715
rect 14715 17685 14720 17715
rect 14680 17680 14720 17685
rect 16760 17715 16800 17720
rect 16760 17685 16765 17715
rect 16795 17685 16800 17715
rect 16760 17680 16800 17685
rect 16840 17715 16880 17720
rect 16840 17685 16845 17715
rect 16875 17685 16880 17715
rect 16840 17680 16880 17685
rect 16920 17715 16960 17720
rect 16920 17685 16925 17715
rect 16955 17685 16960 17715
rect 16920 17680 16960 17685
rect 17000 17715 17040 17720
rect 17000 17685 17005 17715
rect 17035 17685 17040 17715
rect 17000 17680 17040 17685
rect 17080 17715 17120 17720
rect 17080 17685 17085 17715
rect 17115 17685 17120 17715
rect 17080 17680 17120 17685
rect 17160 17715 17200 17720
rect 17160 17685 17165 17715
rect 17195 17685 17200 17715
rect 17160 17680 17200 17685
rect 17240 17715 17280 17720
rect 17240 17685 17245 17715
rect 17275 17685 17280 17715
rect 17240 17680 17280 17685
rect 17320 17715 17360 17720
rect 17320 17685 17325 17715
rect 17355 17685 17360 17715
rect 17320 17680 17360 17685
rect 17400 17715 17440 17720
rect 17400 17685 17405 17715
rect 17435 17685 17440 17715
rect 17400 17680 17440 17685
rect 17480 17715 17520 17720
rect 17480 17685 17485 17715
rect 17515 17685 17520 17715
rect 17480 17680 17520 17685
rect 17560 17715 17600 17720
rect 17560 17685 17565 17715
rect 17595 17685 17600 17715
rect 17560 17680 17600 17685
rect 17640 17715 17680 17720
rect 17640 17685 17645 17715
rect 17675 17685 17680 17715
rect 17640 17680 17680 17685
rect 17720 17715 17760 17720
rect 17720 17685 17725 17715
rect 17755 17685 17760 17715
rect 17720 17680 17760 17685
rect 17800 17715 17840 17720
rect 17800 17685 17805 17715
rect 17835 17685 17840 17715
rect 17800 17680 17840 17685
rect 17880 17715 17920 17720
rect 17880 17685 17885 17715
rect 17915 17685 17920 17715
rect 17880 17680 17920 17685
rect 17960 17715 18000 17720
rect 17960 17685 17965 17715
rect 17995 17685 18000 17715
rect 17960 17680 18000 17685
rect 18040 17715 18080 17720
rect 18040 17685 18045 17715
rect 18075 17685 18080 17715
rect 18040 17680 18080 17685
rect 18120 17715 18160 17720
rect 18120 17685 18125 17715
rect 18155 17685 18160 17715
rect 18120 17680 18160 17685
rect 18200 17715 18240 17720
rect 18200 17685 18205 17715
rect 18235 17685 18240 17715
rect 18200 17680 18240 17685
rect 18280 17715 18320 17720
rect 18280 17685 18285 17715
rect 18315 17685 18320 17715
rect 18280 17680 18320 17685
rect 18360 17715 18400 17720
rect 18360 17685 18365 17715
rect 18395 17685 18400 17715
rect 18360 17680 18400 17685
rect 18440 17715 18480 17720
rect 18440 17685 18445 17715
rect 18475 17685 18480 17715
rect 18440 17680 18480 17685
rect 18520 17715 18560 17720
rect 18520 17685 18525 17715
rect 18555 17685 18560 17715
rect 18520 17680 18560 17685
rect 18600 17715 18640 17720
rect 18600 17685 18605 17715
rect 18635 17685 18640 17715
rect 18600 17680 18640 17685
rect 18680 17715 18720 17720
rect 18680 17685 18685 17715
rect 18715 17685 18720 17715
rect 18680 17680 18720 17685
rect 18760 17715 18800 17720
rect 18760 17685 18765 17715
rect 18795 17685 18800 17715
rect 18760 17680 18800 17685
rect 18840 17715 18880 17720
rect 18840 17685 18845 17715
rect 18875 17685 18880 17715
rect 18840 17680 18880 17685
rect 18920 17715 18960 17720
rect 18920 17685 18925 17715
rect 18955 17685 18960 17715
rect 18920 17680 18960 17685
rect 19000 17715 19040 17720
rect 19000 17685 19005 17715
rect 19035 17685 19040 17715
rect 19000 17680 19040 17685
rect 19080 17715 19120 17720
rect 19080 17685 19085 17715
rect 19115 17685 19120 17715
rect 19080 17680 19120 17685
rect 19160 17715 19200 17720
rect 19160 17685 19165 17715
rect 19195 17685 19200 17715
rect 19160 17680 19200 17685
rect 19240 17715 19280 17720
rect 19240 17685 19245 17715
rect 19275 17685 19280 17715
rect 19240 17680 19280 17685
rect 19320 17715 19360 17720
rect 19320 17685 19325 17715
rect 19355 17685 19360 17715
rect 19320 17680 19360 17685
rect 19400 17715 19440 17720
rect 19400 17685 19405 17715
rect 19435 17685 19440 17715
rect 19400 17680 19440 17685
rect 19480 17715 19520 17720
rect 19480 17685 19485 17715
rect 19515 17685 19520 17715
rect 19480 17680 19520 17685
rect 19560 17715 19600 17720
rect 19560 17685 19565 17715
rect 19595 17685 19600 17715
rect 19560 17680 19600 17685
rect 19640 17715 19680 17720
rect 19640 17685 19645 17715
rect 19675 17685 19680 17715
rect 19640 17680 19680 17685
rect 19720 17715 19760 17720
rect 19720 17685 19725 17715
rect 19755 17685 19760 17715
rect 19720 17680 19760 17685
rect 19800 17715 19840 17720
rect 19800 17685 19805 17715
rect 19835 17685 19840 17715
rect 19800 17680 19840 17685
rect 19880 17715 19920 17720
rect 19880 17685 19885 17715
rect 19915 17685 19920 17715
rect 19880 17680 19920 17685
rect 19960 17715 20000 17720
rect 19960 17685 19965 17715
rect 19995 17685 20000 17715
rect 19960 17680 20000 17685
rect 20040 17715 20080 17720
rect 20040 17685 20045 17715
rect 20075 17685 20080 17715
rect 20040 17680 20080 17685
rect 20120 17715 20160 17720
rect 20120 17685 20125 17715
rect 20155 17685 20160 17715
rect 20120 17680 20160 17685
rect 20200 17715 20240 17720
rect 20200 17685 20205 17715
rect 20235 17685 20240 17715
rect 20200 17680 20240 17685
rect 20280 17715 20320 17720
rect 20280 17685 20285 17715
rect 20315 17685 20320 17715
rect 20280 17680 20320 17685
rect 20360 17715 20400 17720
rect 20360 17685 20365 17715
rect 20395 17685 20400 17715
rect 20360 17680 20400 17685
rect 20440 17715 20480 17720
rect 20440 17685 20445 17715
rect 20475 17685 20480 17715
rect 20440 17680 20480 17685
rect 20520 17715 20560 17720
rect 20520 17685 20525 17715
rect 20555 17685 20560 17715
rect 20520 17680 20560 17685
rect 20600 17715 20640 17720
rect 20600 17685 20605 17715
rect 20635 17685 20640 17715
rect 20600 17680 20640 17685
rect 20680 17715 20720 17720
rect 20680 17685 20685 17715
rect 20715 17685 20720 17715
rect 20680 17680 20720 17685
rect 20760 17715 20800 17720
rect 20760 17685 20765 17715
rect 20795 17685 20800 17715
rect 20760 17680 20800 17685
rect 20840 17715 20880 17720
rect 20840 17685 20845 17715
rect 20875 17685 20880 17715
rect 20840 17680 20880 17685
rect 20920 17715 20960 17720
rect 20920 17685 20925 17715
rect 20955 17685 20960 17715
rect 20920 17680 20960 17685
rect 0 17555 40 17560
rect 0 17525 5 17555
rect 35 17525 40 17555
rect 0 17520 40 17525
rect 80 17555 120 17560
rect 80 17525 85 17555
rect 115 17525 120 17555
rect 80 17520 120 17525
rect 160 17555 200 17560
rect 160 17525 165 17555
rect 195 17525 200 17555
rect 160 17520 200 17525
rect 240 17555 280 17560
rect 240 17525 245 17555
rect 275 17525 280 17555
rect 240 17520 280 17525
rect 320 17555 360 17560
rect 320 17525 325 17555
rect 355 17525 360 17555
rect 320 17520 360 17525
rect 400 17555 440 17560
rect 400 17525 405 17555
rect 435 17525 440 17555
rect 400 17520 440 17525
rect 480 17555 520 17560
rect 480 17525 485 17555
rect 515 17525 520 17555
rect 480 17520 520 17525
rect 560 17555 600 17560
rect 560 17525 565 17555
rect 595 17525 600 17555
rect 560 17520 600 17525
rect 640 17555 680 17560
rect 640 17525 645 17555
rect 675 17525 680 17555
rect 640 17520 680 17525
rect 720 17555 760 17560
rect 720 17525 725 17555
rect 755 17525 760 17555
rect 720 17520 760 17525
rect 800 17555 840 17560
rect 800 17525 805 17555
rect 835 17525 840 17555
rect 800 17520 840 17525
rect 880 17555 920 17560
rect 880 17525 885 17555
rect 915 17525 920 17555
rect 880 17520 920 17525
rect 960 17555 1000 17560
rect 960 17525 965 17555
rect 995 17525 1000 17555
rect 960 17520 1000 17525
rect 1040 17555 1080 17560
rect 1040 17525 1045 17555
rect 1075 17525 1080 17555
rect 1040 17520 1080 17525
rect 1120 17555 1160 17560
rect 1120 17525 1125 17555
rect 1155 17525 1160 17555
rect 1120 17520 1160 17525
rect 1200 17555 1240 17560
rect 1200 17525 1205 17555
rect 1235 17525 1240 17555
rect 1200 17520 1240 17525
rect 1280 17555 1320 17560
rect 1280 17525 1285 17555
rect 1315 17525 1320 17555
rect 1280 17520 1320 17525
rect 1360 17555 1400 17560
rect 1360 17525 1365 17555
rect 1395 17525 1400 17555
rect 1360 17520 1400 17525
rect 1440 17555 1480 17560
rect 1440 17525 1445 17555
rect 1475 17525 1480 17555
rect 1440 17520 1480 17525
rect 1520 17555 1560 17560
rect 1520 17525 1525 17555
rect 1555 17525 1560 17555
rect 1520 17520 1560 17525
rect 1600 17555 1640 17560
rect 1600 17525 1605 17555
rect 1635 17525 1640 17555
rect 1600 17520 1640 17525
rect 1680 17555 1720 17560
rect 1680 17525 1685 17555
rect 1715 17525 1720 17555
rect 1680 17520 1720 17525
rect 1760 17555 1800 17560
rect 1760 17525 1765 17555
rect 1795 17525 1800 17555
rect 1760 17520 1800 17525
rect 1840 17555 1880 17560
rect 1840 17525 1845 17555
rect 1875 17525 1880 17555
rect 1840 17520 1880 17525
rect 1920 17555 1960 17560
rect 1920 17525 1925 17555
rect 1955 17525 1960 17555
rect 1920 17520 1960 17525
rect 2000 17555 2040 17560
rect 2000 17525 2005 17555
rect 2035 17525 2040 17555
rect 2000 17520 2040 17525
rect 2080 17555 2120 17560
rect 2080 17525 2085 17555
rect 2115 17525 2120 17555
rect 2080 17520 2120 17525
rect 2160 17555 2200 17560
rect 2160 17525 2165 17555
rect 2195 17525 2200 17555
rect 2160 17520 2200 17525
rect 2240 17555 2280 17560
rect 2240 17525 2245 17555
rect 2275 17525 2280 17555
rect 2240 17520 2280 17525
rect 2320 17555 2360 17560
rect 2320 17525 2325 17555
rect 2355 17525 2360 17555
rect 2320 17520 2360 17525
rect 2400 17555 2440 17560
rect 2400 17525 2405 17555
rect 2435 17525 2440 17555
rect 2400 17520 2440 17525
rect 2480 17555 2520 17560
rect 2480 17525 2485 17555
rect 2515 17525 2520 17555
rect 2480 17520 2520 17525
rect 2560 17555 2600 17560
rect 2560 17525 2565 17555
rect 2595 17525 2600 17555
rect 2560 17520 2600 17525
rect 2640 17555 2680 17560
rect 2640 17525 2645 17555
rect 2675 17525 2680 17555
rect 2640 17520 2680 17525
rect 2720 17555 2760 17560
rect 2720 17525 2725 17555
rect 2755 17525 2760 17555
rect 2720 17520 2760 17525
rect 2800 17555 2840 17560
rect 2800 17525 2805 17555
rect 2835 17525 2840 17555
rect 2800 17520 2840 17525
rect 2880 17555 2920 17560
rect 2880 17525 2885 17555
rect 2915 17525 2920 17555
rect 2880 17520 2920 17525
rect 2960 17555 3000 17560
rect 2960 17525 2965 17555
rect 2995 17525 3000 17555
rect 2960 17520 3000 17525
rect 3040 17555 3080 17560
rect 3040 17525 3045 17555
rect 3075 17525 3080 17555
rect 3040 17520 3080 17525
rect 3120 17555 3160 17560
rect 3120 17525 3125 17555
rect 3155 17525 3160 17555
rect 3120 17520 3160 17525
rect 3200 17555 3240 17560
rect 3200 17525 3205 17555
rect 3235 17525 3240 17555
rect 3200 17520 3240 17525
rect 3280 17555 3320 17560
rect 3280 17525 3285 17555
rect 3315 17525 3320 17555
rect 3280 17520 3320 17525
rect 3360 17555 3400 17560
rect 3360 17525 3365 17555
rect 3395 17525 3400 17555
rect 3360 17520 3400 17525
rect 3440 17555 3480 17560
rect 3440 17525 3445 17555
rect 3475 17525 3480 17555
rect 3440 17520 3480 17525
rect 3520 17555 3560 17560
rect 3520 17525 3525 17555
rect 3555 17525 3560 17555
rect 3520 17520 3560 17525
rect 3600 17555 3640 17560
rect 3600 17525 3605 17555
rect 3635 17525 3640 17555
rect 3600 17520 3640 17525
rect 3680 17555 3720 17560
rect 3680 17525 3685 17555
rect 3715 17525 3720 17555
rect 3680 17520 3720 17525
rect 3760 17555 3800 17560
rect 3760 17525 3765 17555
rect 3795 17525 3800 17555
rect 3760 17520 3800 17525
rect 3840 17555 3880 17560
rect 3840 17525 3845 17555
rect 3875 17525 3880 17555
rect 3840 17520 3880 17525
rect 3920 17555 3960 17560
rect 3920 17525 3925 17555
rect 3955 17525 3960 17555
rect 3920 17520 3960 17525
rect 4000 17555 4040 17560
rect 4000 17525 4005 17555
rect 4035 17525 4040 17555
rect 4000 17520 4040 17525
rect 4080 17555 4120 17560
rect 4080 17525 4085 17555
rect 4115 17525 4120 17555
rect 4080 17520 4120 17525
rect 4160 17555 4200 17560
rect 4160 17525 4165 17555
rect 4195 17525 4200 17555
rect 4160 17520 4200 17525
rect 6240 17555 6280 17560
rect 6240 17525 6245 17555
rect 6275 17525 6280 17555
rect 6240 17520 6280 17525
rect 6320 17555 6360 17560
rect 6320 17525 6325 17555
rect 6355 17525 6360 17555
rect 6320 17520 6360 17525
rect 6400 17555 6440 17560
rect 6400 17525 6405 17555
rect 6435 17525 6440 17555
rect 6400 17520 6440 17525
rect 6480 17555 6520 17560
rect 6480 17525 6485 17555
rect 6515 17525 6520 17555
rect 6480 17520 6520 17525
rect 6560 17555 6600 17560
rect 6560 17525 6565 17555
rect 6595 17525 6600 17555
rect 6560 17520 6600 17525
rect 6640 17555 6680 17560
rect 6640 17525 6645 17555
rect 6675 17525 6680 17555
rect 6640 17520 6680 17525
rect 6720 17555 6760 17560
rect 6720 17525 6725 17555
rect 6755 17525 6760 17555
rect 6720 17520 6760 17525
rect 6800 17555 6840 17560
rect 6800 17525 6805 17555
rect 6835 17525 6840 17555
rect 6800 17520 6840 17525
rect 6880 17555 6920 17560
rect 6880 17525 6885 17555
rect 6915 17525 6920 17555
rect 6880 17520 6920 17525
rect 6960 17555 7000 17560
rect 6960 17525 6965 17555
rect 6995 17525 7000 17555
rect 6960 17520 7000 17525
rect 7040 17555 7080 17560
rect 7040 17525 7045 17555
rect 7075 17525 7080 17555
rect 7040 17520 7080 17525
rect 7120 17555 7160 17560
rect 7120 17525 7125 17555
rect 7155 17525 7160 17555
rect 7120 17520 7160 17525
rect 7200 17555 7240 17560
rect 7200 17525 7205 17555
rect 7235 17525 7240 17555
rect 7200 17520 7240 17525
rect 7280 17555 7320 17560
rect 7280 17525 7285 17555
rect 7315 17525 7320 17555
rect 7280 17520 7320 17525
rect 7360 17555 7400 17560
rect 7360 17525 7365 17555
rect 7395 17525 7400 17555
rect 7360 17520 7400 17525
rect 7440 17555 7480 17560
rect 7440 17525 7445 17555
rect 7475 17525 7480 17555
rect 7440 17520 7480 17525
rect 7520 17555 7560 17560
rect 7520 17525 7525 17555
rect 7555 17525 7560 17555
rect 7520 17520 7560 17525
rect 7600 17555 7640 17560
rect 7600 17525 7605 17555
rect 7635 17525 7640 17555
rect 7600 17520 7640 17525
rect 7680 17555 7720 17560
rect 7680 17525 7685 17555
rect 7715 17525 7720 17555
rect 7680 17520 7720 17525
rect 7760 17555 7800 17560
rect 7760 17525 7765 17555
rect 7795 17525 7800 17555
rect 7760 17520 7800 17525
rect 7840 17555 7880 17560
rect 7840 17525 7845 17555
rect 7875 17525 7880 17555
rect 7840 17520 7880 17525
rect 7920 17555 7960 17560
rect 7920 17525 7925 17555
rect 7955 17525 7960 17555
rect 7920 17520 7960 17525
rect 8000 17555 8040 17560
rect 8000 17525 8005 17555
rect 8035 17525 8040 17555
rect 8000 17520 8040 17525
rect 8080 17555 8120 17560
rect 8080 17525 8085 17555
rect 8115 17525 8120 17555
rect 8080 17520 8120 17525
rect 8160 17555 8200 17560
rect 8160 17525 8165 17555
rect 8195 17525 8200 17555
rect 8160 17520 8200 17525
rect 8240 17555 8280 17560
rect 8240 17525 8245 17555
rect 8275 17525 8280 17555
rect 8240 17520 8280 17525
rect 8320 17555 8360 17560
rect 8320 17525 8325 17555
rect 8355 17525 8360 17555
rect 8320 17520 8360 17525
rect 8400 17555 8440 17560
rect 8400 17525 8405 17555
rect 8435 17525 8440 17555
rect 8400 17520 8440 17525
rect 8480 17555 8520 17560
rect 8480 17525 8485 17555
rect 8515 17525 8520 17555
rect 8480 17520 8520 17525
rect 8560 17555 8600 17560
rect 8560 17525 8565 17555
rect 8595 17525 8600 17555
rect 8560 17520 8600 17525
rect 8640 17555 8680 17560
rect 8640 17525 8645 17555
rect 8675 17525 8680 17555
rect 8640 17520 8680 17525
rect 8720 17555 8760 17560
rect 8720 17525 8725 17555
rect 8755 17525 8760 17555
rect 8720 17520 8760 17525
rect 8800 17555 8840 17560
rect 8800 17525 8805 17555
rect 8835 17525 8840 17555
rect 8800 17520 8840 17525
rect 8880 17555 8920 17560
rect 8880 17525 8885 17555
rect 8915 17525 8920 17555
rect 8880 17520 8920 17525
rect 8960 17555 9000 17560
rect 8960 17525 8965 17555
rect 8995 17525 9000 17555
rect 8960 17520 9000 17525
rect 9040 17555 9080 17560
rect 9040 17525 9045 17555
rect 9075 17525 9080 17555
rect 9040 17520 9080 17525
rect 9120 17555 9160 17560
rect 9120 17525 9125 17555
rect 9155 17525 9160 17555
rect 9120 17520 9160 17525
rect 9200 17555 9240 17560
rect 9200 17525 9205 17555
rect 9235 17525 9240 17555
rect 9200 17520 9240 17525
rect 9280 17555 9320 17560
rect 9280 17525 9285 17555
rect 9315 17525 9320 17555
rect 9280 17520 9320 17525
rect 9360 17555 9400 17560
rect 9360 17525 9365 17555
rect 9395 17525 9400 17555
rect 9360 17520 9400 17525
rect 9440 17555 9480 17560
rect 9440 17525 9445 17555
rect 9475 17525 9480 17555
rect 9440 17520 9480 17525
rect 11560 17555 11600 17560
rect 11560 17525 11565 17555
rect 11595 17525 11600 17555
rect 11560 17520 11600 17525
rect 11640 17555 11680 17560
rect 11640 17525 11645 17555
rect 11675 17525 11680 17555
rect 11640 17520 11680 17525
rect 11720 17555 11760 17560
rect 11720 17525 11725 17555
rect 11755 17525 11760 17555
rect 11720 17520 11760 17525
rect 11800 17555 11840 17560
rect 11800 17525 11805 17555
rect 11835 17525 11840 17555
rect 11800 17520 11840 17525
rect 11880 17555 11920 17560
rect 11880 17525 11885 17555
rect 11915 17525 11920 17555
rect 11880 17520 11920 17525
rect 11960 17555 12000 17560
rect 11960 17525 11965 17555
rect 11995 17525 12000 17555
rect 11960 17520 12000 17525
rect 12040 17555 12080 17560
rect 12040 17525 12045 17555
rect 12075 17525 12080 17555
rect 12040 17520 12080 17525
rect 12120 17555 12160 17560
rect 12120 17525 12125 17555
rect 12155 17525 12160 17555
rect 12120 17520 12160 17525
rect 12200 17555 12240 17560
rect 12200 17525 12205 17555
rect 12235 17525 12240 17555
rect 12200 17520 12240 17525
rect 12280 17555 12320 17560
rect 12280 17525 12285 17555
rect 12315 17525 12320 17555
rect 12280 17520 12320 17525
rect 12360 17555 12400 17560
rect 12360 17525 12365 17555
rect 12395 17525 12400 17555
rect 12360 17520 12400 17525
rect 12440 17555 12480 17560
rect 12440 17525 12445 17555
rect 12475 17525 12480 17555
rect 12440 17520 12480 17525
rect 12520 17555 12560 17560
rect 12520 17525 12525 17555
rect 12555 17525 12560 17555
rect 12520 17520 12560 17525
rect 12600 17555 12640 17560
rect 12600 17525 12605 17555
rect 12635 17525 12640 17555
rect 12600 17520 12640 17525
rect 12680 17555 12720 17560
rect 12680 17525 12685 17555
rect 12715 17525 12720 17555
rect 12680 17520 12720 17525
rect 12760 17555 12800 17560
rect 12760 17525 12765 17555
rect 12795 17525 12800 17555
rect 12760 17520 12800 17525
rect 12840 17555 12880 17560
rect 12840 17525 12845 17555
rect 12875 17525 12880 17555
rect 12840 17520 12880 17525
rect 12920 17555 12960 17560
rect 12920 17525 12925 17555
rect 12955 17525 12960 17555
rect 12920 17520 12960 17525
rect 13000 17555 13040 17560
rect 13000 17525 13005 17555
rect 13035 17525 13040 17555
rect 13000 17520 13040 17525
rect 13080 17555 13120 17560
rect 13080 17525 13085 17555
rect 13115 17525 13120 17555
rect 13080 17520 13120 17525
rect 13160 17555 13200 17560
rect 13160 17525 13165 17555
rect 13195 17525 13200 17555
rect 13160 17520 13200 17525
rect 13240 17555 13280 17560
rect 13240 17525 13245 17555
rect 13275 17525 13280 17555
rect 13240 17520 13280 17525
rect 13320 17555 13360 17560
rect 13320 17525 13325 17555
rect 13355 17525 13360 17555
rect 13320 17520 13360 17525
rect 13400 17555 13440 17560
rect 13400 17525 13405 17555
rect 13435 17525 13440 17555
rect 13400 17520 13440 17525
rect 13480 17555 13520 17560
rect 13480 17525 13485 17555
rect 13515 17525 13520 17555
rect 13480 17520 13520 17525
rect 13560 17555 13600 17560
rect 13560 17525 13565 17555
rect 13595 17525 13600 17555
rect 13560 17520 13600 17525
rect 13640 17555 13680 17560
rect 13640 17525 13645 17555
rect 13675 17525 13680 17555
rect 13640 17520 13680 17525
rect 13720 17555 13760 17560
rect 13720 17525 13725 17555
rect 13755 17525 13760 17555
rect 13720 17520 13760 17525
rect 13800 17555 13840 17560
rect 13800 17525 13805 17555
rect 13835 17525 13840 17555
rect 13800 17520 13840 17525
rect 13880 17555 13920 17560
rect 13880 17525 13885 17555
rect 13915 17525 13920 17555
rect 13880 17520 13920 17525
rect 13960 17555 14000 17560
rect 13960 17525 13965 17555
rect 13995 17525 14000 17555
rect 13960 17520 14000 17525
rect 14040 17555 14080 17560
rect 14040 17525 14045 17555
rect 14075 17525 14080 17555
rect 14040 17520 14080 17525
rect 14120 17555 14160 17560
rect 14120 17525 14125 17555
rect 14155 17525 14160 17555
rect 14120 17520 14160 17525
rect 14200 17555 14240 17560
rect 14200 17525 14205 17555
rect 14235 17525 14240 17555
rect 14200 17520 14240 17525
rect 14280 17555 14320 17560
rect 14280 17525 14285 17555
rect 14315 17525 14320 17555
rect 14280 17520 14320 17525
rect 14360 17555 14400 17560
rect 14360 17525 14365 17555
rect 14395 17525 14400 17555
rect 14360 17520 14400 17525
rect 14440 17555 14480 17560
rect 14440 17525 14445 17555
rect 14475 17525 14480 17555
rect 14440 17520 14480 17525
rect 14520 17555 14560 17560
rect 14520 17525 14525 17555
rect 14555 17525 14560 17555
rect 14520 17520 14560 17525
rect 14600 17555 14640 17560
rect 14600 17525 14605 17555
rect 14635 17525 14640 17555
rect 14600 17520 14640 17525
rect 14680 17555 14720 17560
rect 14680 17525 14685 17555
rect 14715 17525 14720 17555
rect 14680 17520 14720 17525
rect 16760 17555 16800 17560
rect 16760 17525 16765 17555
rect 16795 17525 16800 17555
rect 16760 17520 16800 17525
rect 16840 17555 16880 17560
rect 16840 17525 16845 17555
rect 16875 17525 16880 17555
rect 16840 17520 16880 17525
rect 16920 17555 16960 17560
rect 16920 17525 16925 17555
rect 16955 17525 16960 17555
rect 16920 17520 16960 17525
rect 17000 17555 17040 17560
rect 17000 17525 17005 17555
rect 17035 17525 17040 17555
rect 17000 17520 17040 17525
rect 17080 17555 17120 17560
rect 17080 17525 17085 17555
rect 17115 17525 17120 17555
rect 17080 17520 17120 17525
rect 17160 17555 17200 17560
rect 17160 17525 17165 17555
rect 17195 17525 17200 17555
rect 17160 17520 17200 17525
rect 17240 17555 17280 17560
rect 17240 17525 17245 17555
rect 17275 17525 17280 17555
rect 17240 17520 17280 17525
rect 17320 17555 17360 17560
rect 17320 17525 17325 17555
rect 17355 17525 17360 17555
rect 17320 17520 17360 17525
rect 17400 17555 17440 17560
rect 17400 17525 17405 17555
rect 17435 17525 17440 17555
rect 17400 17520 17440 17525
rect 17480 17555 17520 17560
rect 17480 17525 17485 17555
rect 17515 17525 17520 17555
rect 17480 17520 17520 17525
rect 17560 17555 17600 17560
rect 17560 17525 17565 17555
rect 17595 17525 17600 17555
rect 17560 17520 17600 17525
rect 17640 17555 17680 17560
rect 17640 17525 17645 17555
rect 17675 17525 17680 17555
rect 17640 17520 17680 17525
rect 17720 17555 17760 17560
rect 17720 17525 17725 17555
rect 17755 17525 17760 17555
rect 17720 17520 17760 17525
rect 17800 17555 17840 17560
rect 17800 17525 17805 17555
rect 17835 17525 17840 17555
rect 17800 17520 17840 17525
rect 17880 17555 17920 17560
rect 17880 17525 17885 17555
rect 17915 17525 17920 17555
rect 17880 17520 17920 17525
rect 17960 17555 18000 17560
rect 17960 17525 17965 17555
rect 17995 17525 18000 17555
rect 17960 17520 18000 17525
rect 18040 17555 18080 17560
rect 18040 17525 18045 17555
rect 18075 17525 18080 17555
rect 18040 17520 18080 17525
rect 18120 17555 18160 17560
rect 18120 17525 18125 17555
rect 18155 17525 18160 17555
rect 18120 17520 18160 17525
rect 18200 17555 18240 17560
rect 18200 17525 18205 17555
rect 18235 17525 18240 17555
rect 18200 17520 18240 17525
rect 18280 17555 18320 17560
rect 18280 17525 18285 17555
rect 18315 17525 18320 17555
rect 18280 17520 18320 17525
rect 18360 17555 18400 17560
rect 18360 17525 18365 17555
rect 18395 17525 18400 17555
rect 18360 17520 18400 17525
rect 18440 17555 18480 17560
rect 18440 17525 18445 17555
rect 18475 17525 18480 17555
rect 18440 17520 18480 17525
rect 18520 17555 18560 17560
rect 18520 17525 18525 17555
rect 18555 17525 18560 17555
rect 18520 17520 18560 17525
rect 18600 17555 18640 17560
rect 18600 17525 18605 17555
rect 18635 17525 18640 17555
rect 18600 17520 18640 17525
rect 18680 17555 18720 17560
rect 18680 17525 18685 17555
rect 18715 17525 18720 17555
rect 18680 17520 18720 17525
rect 18760 17555 18800 17560
rect 18760 17525 18765 17555
rect 18795 17525 18800 17555
rect 18760 17520 18800 17525
rect 18840 17555 18880 17560
rect 18840 17525 18845 17555
rect 18875 17525 18880 17555
rect 18840 17520 18880 17525
rect 18920 17555 18960 17560
rect 18920 17525 18925 17555
rect 18955 17525 18960 17555
rect 18920 17520 18960 17525
rect 19000 17555 19040 17560
rect 19000 17525 19005 17555
rect 19035 17525 19040 17555
rect 19000 17520 19040 17525
rect 19080 17555 19120 17560
rect 19080 17525 19085 17555
rect 19115 17525 19120 17555
rect 19080 17520 19120 17525
rect 19160 17555 19200 17560
rect 19160 17525 19165 17555
rect 19195 17525 19200 17555
rect 19160 17520 19200 17525
rect 19240 17555 19280 17560
rect 19240 17525 19245 17555
rect 19275 17525 19280 17555
rect 19240 17520 19280 17525
rect 19320 17555 19360 17560
rect 19320 17525 19325 17555
rect 19355 17525 19360 17555
rect 19320 17520 19360 17525
rect 19400 17555 19440 17560
rect 19400 17525 19405 17555
rect 19435 17525 19440 17555
rect 19400 17520 19440 17525
rect 19480 17555 19520 17560
rect 19480 17525 19485 17555
rect 19515 17525 19520 17555
rect 19480 17520 19520 17525
rect 19560 17555 19600 17560
rect 19560 17525 19565 17555
rect 19595 17525 19600 17555
rect 19560 17520 19600 17525
rect 19640 17555 19680 17560
rect 19640 17525 19645 17555
rect 19675 17525 19680 17555
rect 19640 17520 19680 17525
rect 19720 17555 19760 17560
rect 19720 17525 19725 17555
rect 19755 17525 19760 17555
rect 19720 17520 19760 17525
rect 19800 17555 19840 17560
rect 19800 17525 19805 17555
rect 19835 17525 19840 17555
rect 19800 17520 19840 17525
rect 19880 17555 19920 17560
rect 19880 17525 19885 17555
rect 19915 17525 19920 17555
rect 19880 17520 19920 17525
rect 19960 17555 20000 17560
rect 19960 17525 19965 17555
rect 19995 17525 20000 17555
rect 19960 17520 20000 17525
rect 20040 17555 20080 17560
rect 20040 17525 20045 17555
rect 20075 17525 20080 17555
rect 20040 17520 20080 17525
rect 20120 17555 20160 17560
rect 20120 17525 20125 17555
rect 20155 17525 20160 17555
rect 20120 17520 20160 17525
rect 20200 17555 20240 17560
rect 20200 17525 20205 17555
rect 20235 17525 20240 17555
rect 20200 17520 20240 17525
rect 20280 17555 20320 17560
rect 20280 17525 20285 17555
rect 20315 17525 20320 17555
rect 20280 17520 20320 17525
rect 20360 17555 20400 17560
rect 20360 17525 20365 17555
rect 20395 17525 20400 17555
rect 20360 17520 20400 17525
rect 20440 17555 20480 17560
rect 20440 17525 20445 17555
rect 20475 17525 20480 17555
rect 20440 17520 20480 17525
rect 20520 17555 20560 17560
rect 20520 17525 20525 17555
rect 20555 17525 20560 17555
rect 20520 17520 20560 17525
rect 20600 17555 20640 17560
rect 20600 17525 20605 17555
rect 20635 17525 20640 17555
rect 20600 17520 20640 17525
rect 20680 17555 20720 17560
rect 20680 17525 20685 17555
rect 20715 17525 20720 17555
rect 20680 17520 20720 17525
rect 20760 17555 20800 17560
rect 20760 17525 20765 17555
rect 20795 17525 20800 17555
rect 20760 17520 20800 17525
rect 20840 17555 20880 17560
rect 20840 17525 20845 17555
rect 20875 17525 20880 17555
rect 20840 17520 20880 17525
rect 20920 17555 20960 17560
rect 20920 17525 20925 17555
rect 20955 17525 20960 17555
rect 20920 17520 20960 17525
rect 0 17395 40 17400
rect 0 17365 5 17395
rect 35 17365 40 17395
rect 0 17360 40 17365
rect 80 17395 120 17400
rect 80 17365 85 17395
rect 115 17365 120 17395
rect 80 17360 120 17365
rect 160 17395 200 17400
rect 160 17365 165 17395
rect 195 17365 200 17395
rect 160 17360 200 17365
rect 240 17395 280 17400
rect 240 17365 245 17395
rect 275 17365 280 17395
rect 240 17360 280 17365
rect 320 17395 360 17400
rect 320 17365 325 17395
rect 355 17365 360 17395
rect 320 17360 360 17365
rect 400 17395 440 17400
rect 400 17365 405 17395
rect 435 17365 440 17395
rect 400 17360 440 17365
rect 480 17395 520 17400
rect 480 17365 485 17395
rect 515 17365 520 17395
rect 480 17360 520 17365
rect 560 17395 600 17400
rect 560 17365 565 17395
rect 595 17365 600 17395
rect 560 17360 600 17365
rect 640 17395 680 17400
rect 640 17365 645 17395
rect 675 17365 680 17395
rect 640 17360 680 17365
rect 720 17395 760 17400
rect 720 17365 725 17395
rect 755 17365 760 17395
rect 720 17360 760 17365
rect 800 17395 840 17400
rect 800 17365 805 17395
rect 835 17365 840 17395
rect 800 17360 840 17365
rect 880 17395 920 17400
rect 880 17365 885 17395
rect 915 17365 920 17395
rect 880 17360 920 17365
rect 960 17395 1000 17400
rect 960 17365 965 17395
rect 995 17365 1000 17395
rect 960 17360 1000 17365
rect 1040 17395 1080 17400
rect 1040 17365 1045 17395
rect 1075 17365 1080 17395
rect 1040 17360 1080 17365
rect 1120 17395 1160 17400
rect 1120 17365 1125 17395
rect 1155 17365 1160 17395
rect 1120 17360 1160 17365
rect 1200 17395 1240 17400
rect 1200 17365 1205 17395
rect 1235 17365 1240 17395
rect 1200 17360 1240 17365
rect 1280 17395 1320 17400
rect 1280 17365 1285 17395
rect 1315 17365 1320 17395
rect 1280 17360 1320 17365
rect 1360 17395 1400 17400
rect 1360 17365 1365 17395
rect 1395 17365 1400 17395
rect 1360 17360 1400 17365
rect 1440 17395 1480 17400
rect 1440 17365 1445 17395
rect 1475 17365 1480 17395
rect 1440 17360 1480 17365
rect 1520 17395 1560 17400
rect 1520 17365 1525 17395
rect 1555 17365 1560 17395
rect 1520 17360 1560 17365
rect 1600 17395 1640 17400
rect 1600 17365 1605 17395
rect 1635 17365 1640 17395
rect 1600 17360 1640 17365
rect 1680 17395 1720 17400
rect 1680 17365 1685 17395
rect 1715 17365 1720 17395
rect 1680 17360 1720 17365
rect 1760 17395 1800 17400
rect 1760 17365 1765 17395
rect 1795 17365 1800 17395
rect 1760 17360 1800 17365
rect 1840 17395 1880 17400
rect 1840 17365 1845 17395
rect 1875 17365 1880 17395
rect 1840 17360 1880 17365
rect 1920 17395 1960 17400
rect 1920 17365 1925 17395
rect 1955 17365 1960 17395
rect 1920 17360 1960 17365
rect 2000 17395 2040 17400
rect 2000 17365 2005 17395
rect 2035 17365 2040 17395
rect 2000 17360 2040 17365
rect 2080 17395 2120 17400
rect 2080 17365 2085 17395
rect 2115 17365 2120 17395
rect 2080 17360 2120 17365
rect 2160 17395 2200 17400
rect 2160 17365 2165 17395
rect 2195 17365 2200 17395
rect 2160 17360 2200 17365
rect 2240 17395 2280 17400
rect 2240 17365 2245 17395
rect 2275 17365 2280 17395
rect 2240 17360 2280 17365
rect 2320 17395 2360 17400
rect 2320 17365 2325 17395
rect 2355 17365 2360 17395
rect 2320 17360 2360 17365
rect 2400 17395 2440 17400
rect 2400 17365 2405 17395
rect 2435 17365 2440 17395
rect 2400 17360 2440 17365
rect 2480 17395 2520 17400
rect 2480 17365 2485 17395
rect 2515 17365 2520 17395
rect 2480 17360 2520 17365
rect 2560 17395 2600 17400
rect 2560 17365 2565 17395
rect 2595 17365 2600 17395
rect 2560 17360 2600 17365
rect 2640 17395 2680 17400
rect 2640 17365 2645 17395
rect 2675 17365 2680 17395
rect 2640 17360 2680 17365
rect 2720 17395 2760 17400
rect 2720 17365 2725 17395
rect 2755 17365 2760 17395
rect 2720 17360 2760 17365
rect 2800 17395 2840 17400
rect 2800 17365 2805 17395
rect 2835 17365 2840 17395
rect 2800 17360 2840 17365
rect 2880 17395 2920 17400
rect 2880 17365 2885 17395
rect 2915 17365 2920 17395
rect 2880 17360 2920 17365
rect 2960 17395 3000 17400
rect 2960 17365 2965 17395
rect 2995 17365 3000 17395
rect 2960 17360 3000 17365
rect 3040 17395 3080 17400
rect 3040 17365 3045 17395
rect 3075 17365 3080 17395
rect 3040 17360 3080 17365
rect 3120 17395 3160 17400
rect 3120 17365 3125 17395
rect 3155 17365 3160 17395
rect 3120 17360 3160 17365
rect 3200 17395 3240 17400
rect 3200 17365 3205 17395
rect 3235 17365 3240 17395
rect 3200 17360 3240 17365
rect 3280 17395 3320 17400
rect 3280 17365 3285 17395
rect 3315 17365 3320 17395
rect 3280 17360 3320 17365
rect 3360 17395 3400 17400
rect 3360 17365 3365 17395
rect 3395 17365 3400 17395
rect 3360 17360 3400 17365
rect 3440 17395 3480 17400
rect 3440 17365 3445 17395
rect 3475 17365 3480 17395
rect 3440 17360 3480 17365
rect 3520 17395 3560 17400
rect 3520 17365 3525 17395
rect 3555 17365 3560 17395
rect 3520 17360 3560 17365
rect 3600 17395 3640 17400
rect 3600 17365 3605 17395
rect 3635 17365 3640 17395
rect 3600 17360 3640 17365
rect 3680 17395 3720 17400
rect 3680 17365 3685 17395
rect 3715 17365 3720 17395
rect 3680 17360 3720 17365
rect 3760 17395 3800 17400
rect 3760 17365 3765 17395
rect 3795 17365 3800 17395
rect 3760 17360 3800 17365
rect 3840 17395 3880 17400
rect 3840 17365 3845 17395
rect 3875 17365 3880 17395
rect 3840 17360 3880 17365
rect 3920 17395 3960 17400
rect 3920 17365 3925 17395
rect 3955 17365 3960 17395
rect 3920 17360 3960 17365
rect 4000 17395 4040 17400
rect 4000 17365 4005 17395
rect 4035 17365 4040 17395
rect 4000 17360 4040 17365
rect 4080 17395 4120 17400
rect 4080 17365 4085 17395
rect 4115 17365 4120 17395
rect 4080 17360 4120 17365
rect 4160 17395 4200 17400
rect 4160 17365 4165 17395
rect 4195 17365 4200 17395
rect 4160 17360 4200 17365
rect 6240 17395 6280 17400
rect 6240 17365 6245 17395
rect 6275 17365 6280 17395
rect 6240 17360 6280 17365
rect 6320 17395 6360 17400
rect 6320 17365 6325 17395
rect 6355 17365 6360 17395
rect 6320 17360 6360 17365
rect 6400 17395 6440 17400
rect 6400 17365 6405 17395
rect 6435 17365 6440 17395
rect 6400 17360 6440 17365
rect 6480 17395 6520 17400
rect 6480 17365 6485 17395
rect 6515 17365 6520 17395
rect 6480 17360 6520 17365
rect 6560 17395 6600 17400
rect 6560 17365 6565 17395
rect 6595 17365 6600 17395
rect 6560 17360 6600 17365
rect 6640 17395 6680 17400
rect 6640 17365 6645 17395
rect 6675 17365 6680 17395
rect 6640 17360 6680 17365
rect 6720 17395 6760 17400
rect 6720 17365 6725 17395
rect 6755 17365 6760 17395
rect 6720 17360 6760 17365
rect 6800 17395 6840 17400
rect 6800 17365 6805 17395
rect 6835 17365 6840 17395
rect 6800 17360 6840 17365
rect 6880 17395 6920 17400
rect 6880 17365 6885 17395
rect 6915 17365 6920 17395
rect 6880 17360 6920 17365
rect 6960 17395 7000 17400
rect 6960 17365 6965 17395
rect 6995 17365 7000 17395
rect 6960 17360 7000 17365
rect 7040 17395 7080 17400
rect 7040 17365 7045 17395
rect 7075 17365 7080 17395
rect 7040 17360 7080 17365
rect 7120 17395 7160 17400
rect 7120 17365 7125 17395
rect 7155 17365 7160 17395
rect 7120 17360 7160 17365
rect 7200 17395 7240 17400
rect 7200 17365 7205 17395
rect 7235 17365 7240 17395
rect 7200 17360 7240 17365
rect 7280 17395 7320 17400
rect 7280 17365 7285 17395
rect 7315 17365 7320 17395
rect 7280 17360 7320 17365
rect 7360 17395 7400 17400
rect 7360 17365 7365 17395
rect 7395 17365 7400 17395
rect 7360 17360 7400 17365
rect 7440 17395 7480 17400
rect 7440 17365 7445 17395
rect 7475 17365 7480 17395
rect 7440 17360 7480 17365
rect 7520 17395 7560 17400
rect 7520 17365 7525 17395
rect 7555 17365 7560 17395
rect 7520 17360 7560 17365
rect 7600 17395 7640 17400
rect 7600 17365 7605 17395
rect 7635 17365 7640 17395
rect 7600 17360 7640 17365
rect 7680 17395 7720 17400
rect 7680 17365 7685 17395
rect 7715 17365 7720 17395
rect 7680 17360 7720 17365
rect 7760 17395 7800 17400
rect 7760 17365 7765 17395
rect 7795 17365 7800 17395
rect 7760 17360 7800 17365
rect 7840 17395 7880 17400
rect 7840 17365 7845 17395
rect 7875 17365 7880 17395
rect 7840 17360 7880 17365
rect 7920 17395 7960 17400
rect 7920 17365 7925 17395
rect 7955 17365 7960 17395
rect 7920 17360 7960 17365
rect 8000 17395 8040 17400
rect 8000 17365 8005 17395
rect 8035 17365 8040 17395
rect 8000 17360 8040 17365
rect 8080 17395 8120 17400
rect 8080 17365 8085 17395
rect 8115 17365 8120 17395
rect 8080 17360 8120 17365
rect 8160 17395 8200 17400
rect 8160 17365 8165 17395
rect 8195 17365 8200 17395
rect 8160 17360 8200 17365
rect 8240 17395 8280 17400
rect 8240 17365 8245 17395
rect 8275 17365 8280 17395
rect 8240 17360 8280 17365
rect 8320 17395 8360 17400
rect 8320 17365 8325 17395
rect 8355 17365 8360 17395
rect 8320 17360 8360 17365
rect 8400 17395 8440 17400
rect 8400 17365 8405 17395
rect 8435 17365 8440 17395
rect 8400 17360 8440 17365
rect 8480 17395 8520 17400
rect 8480 17365 8485 17395
rect 8515 17365 8520 17395
rect 8480 17360 8520 17365
rect 8560 17395 8600 17400
rect 8560 17365 8565 17395
rect 8595 17365 8600 17395
rect 8560 17360 8600 17365
rect 8640 17395 8680 17400
rect 8640 17365 8645 17395
rect 8675 17365 8680 17395
rect 8640 17360 8680 17365
rect 8720 17395 8760 17400
rect 8720 17365 8725 17395
rect 8755 17365 8760 17395
rect 8720 17360 8760 17365
rect 8800 17395 8840 17400
rect 8800 17365 8805 17395
rect 8835 17365 8840 17395
rect 8800 17360 8840 17365
rect 8880 17395 8920 17400
rect 8880 17365 8885 17395
rect 8915 17365 8920 17395
rect 8880 17360 8920 17365
rect 8960 17395 9000 17400
rect 8960 17365 8965 17395
rect 8995 17365 9000 17395
rect 8960 17360 9000 17365
rect 9040 17395 9080 17400
rect 9040 17365 9045 17395
rect 9075 17365 9080 17395
rect 9040 17360 9080 17365
rect 9120 17395 9160 17400
rect 9120 17365 9125 17395
rect 9155 17365 9160 17395
rect 9120 17360 9160 17365
rect 9200 17395 9240 17400
rect 9200 17365 9205 17395
rect 9235 17365 9240 17395
rect 9200 17360 9240 17365
rect 9280 17395 9320 17400
rect 9280 17365 9285 17395
rect 9315 17365 9320 17395
rect 9280 17360 9320 17365
rect 9360 17395 9400 17400
rect 9360 17365 9365 17395
rect 9395 17365 9400 17395
rect 9360 17360 9400 17365
rect 9440 17395 9480 17400
rect 9440 17365 9445 17395
rect 9475 17365 9480 17395
rect 9440 17360 9480 17365
rect 11560 17395 11600 17400
rect 11560 17365 11565 17395
rect 11595 17365 11600 17395
rect 11560 17360 11600 17365
rect 11640 17395 11680 17400
rect 11640 17365 11645 17395
rect 11675 17365 11680 17395
rect 11640 17360 11680 17365
rect 11720 17395 11760 17400
rect 11720 17365 11725 17395
rect 11755 17365 11760 17395
rect 11720 17360 11760 17365
rect 11800 17395 11840 17400
rect 11800 17365 11805 17395
rect 11835 17365 11840 17395
rect 11800 17360 11840 17365
rect 11880 17395 11920 17400
rect 11880 17365 11885 17395
rect 11915 17365 11920 17395
rect 11880 17360 11920 17365
rect 11960 17395 12000 17400
rect 11960 17365 11965 17395
rect 11995 17365 12000 17395
rect 11960 17360 12000 17365
rect 12040 17395 12080 17400
rect 12040 17365 12045 17395
rect 12075 17365 12080 17395
rect 12040 17360 12080 17365
rect 12120 17395 12160 17400
rect 12120 17365 12125 17395
rect 12155 17365 12160 17395
rect 12120 17360 12160 17365
rect 12200 17395 12240 17400
rect 12200 17365 12205 17395
rect 12235 17365 12240 17395
rect 12200 17360 12240 17365
rect 12280 17395 12320 17400
rect 12280 17365 12285 17395
rect 12315 17365 12320 17395
rect 12280 17360 12320 17365
rect 12360 17395 12400 17400
rect 12360 17365 12365 17395
rect 12395 17365 12400 17395
rect 12360 17360 12400 17365
rect 12440 17395 12480 17400
rect 12440 17365 12445 17395
rect 12475 17365 12480 17395
rect 12440 17360 12480 17365
rect 12520 17395 12560 17400
rect 12520 17365 12525 17395
rect 12555 17365 12560 17395
rect 12520 17360 12560 17365
rect 12600 17395 12640 17400
rect 12600 17365 12605 17395
rect 12635 17365 12640 17395
rect 12600 17360 12640 17365
rect 12680 17395 12720 17400
rect 12680 17365 12685 17395
rect 12715 17365 12720 17395
rect 12680 17360 12720 17365
rect 12760 17395 12800 17400
rect 12760 17365 12765 17395
rect 12795 17365 12800 17395
rect 12760 17360 12800 17365
rect 12840 17395 12880 17400
rect 12840 17365 12845 17395
rect 12875 17365 12880 17395
rect 12840 17360 12880 17365
rect 12920 17395 12960 17400
rect 12920 17365 12925 17395
rect 12955 17365 12960 17395
rect 12920 17360 12960 17365
rect 13000 17395 13040 17400
rect 13000 17365 13005 17395
rect 13035 17365 13040 17395
rect 13000 17360 13040 17365
rect 13080 17395 13120 17400
rect 13080 17365 13085 17395
rect 13115 17365 13120 17395
rect 13080 17360 13120 17365
rect 13160 17395 13200 17400
rect 13160 17365 13165 17395
rect 13195 17365 13200 17395
rect 13160 17360 13200 17365
rect 13240 17395 13280 17400
rect 13240 17365 13245 17395
rect 13275 17365 13280 17395
rect 13240 17360 13280 17365
rect 13320 17395 13360 17400
rect 13320 17365 13325 17395
rect 13355 17365 13360 17395
rect 13320 17360 13360 17365
rect 13400 17395 13440 17400
rect 13400 17365 13405 17395
rect 13435 17365 13440 17395
rect 13400 17360 13440 17365
rect 13480 17395 13520 17400
rect 13480 17365 13485 17395
rect 13515 17365 13520 17395
rect 13480 17360 13520 17365
rect 13560 17395 13600 17400
rect 13560 17365 13565 17395
rect 13595 17365 13600 17395
rect 13560 17360 13600 17365
rect 13640 17395 13680 17400
rect 13640 17365 13645 17395
rect 13675 17365 13680 17395
rect 13640 17360 13680 17365
rect 13720 17395 13760 17400
rect 13720 17365 13725 17395
rect 13755 17365 13760 17395
rect 13720 17360 13760 17365
rect 13800 17395 13840 17400
rect 13800 17365 13805 17395
rect 13835 17365 13840 17395
rect 13800 17360 13840 17365
rect 13880 17395 13920 17400
rect 13880 17365 13885 17395
rect 13915 17365 13920 17395
rect 13880 17360 13920 17365
rect 13960 17395 14000 17400
rect 13960 17365 13965 17395
rect 13995 17365 14000 17395
rect 13960 17360 14000 17365
rect 14040 17395 14080 17400
rect 14040 17365 14045 17395
rect 14075 17365 14080 17395
rect 14040 17360 14080 17365
rect 14120 17395 14160 17400
rect 14120 17365 14125 17395
rect 14155 17365 14160 17395
rect 14120 17360 14160 17365
rect 14200 17395 14240 17400
rect 14200 17365 14205 17395
rect 14235 17365 14240 17395
rect 14200 17360 14240 17365
rect 14280 17395 14320 17400
rect 14280 17365 14285 17395
rect 14315 17365 14320 17395
rect 14280 17360 14320 17365
rect 14360 17395 14400 17400
rect 14360 17365 14365 17395
rect 14395 17365 14400 17395
rect 14360 17360 14400 17365
rect 14440 17395 14480 17400
rect 14440 17365 14445 17395
rect 14475 17365 14480 17395
rect 14440 17360 14480 17365
rect 14520 17395 14560 17400
rect 14520 17365 14525 17395
rect 14555 17365 14560 17395
rect 14520 17360 14560 17365
rect 14600 17395 14640 17400
rect 14600 17365 14605 17395
rect 14635 17365 14640 17395
rect 14600 17360 14640 17365
rect 14680 17395 14720 17400
rect 14680 17365 14685 17395
rect 14715 17365 14720 17395
rect 14680 17360 14720 17365
rect 16760 17395 16800 17400
rect 16760 17365 16765 17395
rect 16795 17365 16800 17395
rect 16760 17360 16800 17365
rect 16840 17395 16880 17400
rect 16840 17365 16845 17395
rect 16875 17365 16880 17395
rect 16840 17360 16880 17365
rect 16920 17395 16960 17400
rect 16920 17365 16925 17395
rect 16955 17365 16960 17395
rect 16920 17360 16960 17365
rect 17000 17395 17040 17400
rect 17000 17365 17005 17395
rect 17035 17365 17040 17395
rect 17000 17360 17040 17365
rect 17080 17395 17120 17400
rect 17080 17365 17085 17395
rect 17115 17365 17120 17395
rect 17080 17360 17120 17365
rect 17160 17395 17200 17400
rect 17160 17365 17165 17395
rect 17195 17365 17200 17395
rect 17160 17360 17200 17365
rect 17240 17395 17280 17400
rect 17240 17365 17245 17395
rect 17275 17365 17280 17395
rect 17240 17360 17280 17365
rect 17320 17395 17360 17400
rect 17320 17365 17325 17395
rect 17355 17365 17360 17395
rect 17320 17360 17360 17365
rect 17400 17395 17440 17400
rect 17400 17365 17405 17395
rect 17435 17365 17440 17395
rect 17400 17360 17440 17365
rect 17480 17395 17520 17400
rect 17480 17365 17485 17395
rect 17515 17365 17520 17395
rect 17480 17360 17520 17365
rect 17560 17395 17600 17400
rect 17560 17365 17565 17395
rect 17595 17365 17600 17395
rect 17560 17360 17600 17365
rect 17640 17395 17680 17400
rect 17640 17365 17645 17395
rect 17675 17365 17680 17395
rect 17640 17360 17680 17365
rect 17720 17395 17760 17400
rect 17720 17365 17725 17395
rect 17755 17365 17760 17395
rect 17720 17360 17760 17365
rect 17800 17395 17840 17400
rect 17800 17365 17805 17395
rect 17835 17365 17840 17395
rect 17800 17360 17840 17365
rect 17880 17395 17920 17400
rect 17880 17365 17885 17395
rect 17915 17365 17920 17395
rect 17880 17360 17920 17365
rect 17960 17395 18000 17400
rect 17960 17365 17965 17395
rect 17995 17365 18000 17395
rect 17960 17360 18000 17365
rect 18040 17395 18080 17400
rect 18040 17365 18045 17395
rect 18075 17365 18080 17395
rect 18040 17360 18080 17365
rect 18120 17395 18160 17400
rect 18120 17365 18125 17395
rect 18155 17365 18160 17395
rect 18120 17360 18160 17365
rect 18200 17395 18240 17400
rect 18200 17365 18205 17395
rect 18235 17365 18240 17395
rect 18200 17360 18240 17365
rect 18280 17395 18320 17400
rect 18280 17365 18285 17395
rect 18315 17365 18320 17395
rect 18280 17360 18320 17365
rect 18360 17395 18400 17400
rect 18360 17365 18365 17395
rect 18395 17365 18400 17395
rect 18360 17360 18400 17365
rect 18440 17395 18480 17400
rect 18440 17365 18445 17395
rect 18475 17365 18480 17395
rect 18440 17360 18480 17365
rect 18520 17395 18560 17400
rect 18520 17365 18525 17395
rect 18555 17365 18560 17395
rect 18520 17360 18560 17365
rect 18600 17395 18640 17400
rect 18600 17365 18605 17395
rect 18635 17365 18640 17395
rect 18600 17360 18640 17365
rect 18680 17395 18720 17400
rect 18680 17365 18685 17395
rect 18715 17365 18720 17395
rect 18680 17360 18720 17365
rect 18760 17395 18800 17400
rect 18760 17365 18765 17395
rect 18795 17365 18800 17395
rect 18760 17360 18800 17365
rect 18840 17395 18880 17400
rect 18840 17365 18845 17395
rect 18875 17365 18880 17395
rect 18840 17360 18880 17365
rect 18920 17395 18960 17400
rect 18920 17365 18925 17395
rect 18955 17365 18960 17395
rect 18920 17360 18960 17365
rect 19000 17395 19040 17400
rect 19000 17365 19005 17395
rect 19035 17365 19040 17395
rect 19000 17360 19040 17365
rect 19080 17395 19120 17400
rect 19080 17365 19085 17395
rect 19115 17365 19120 17395
rect 19080 17360 19120 17365
rect 19160 17395 19200 17400
rect 19160 17365 19165 17395
rect 19195 17365 19200 17395
rect 19160 17360 19200 17365
rect 19240 17395 19280 17400
rect 19240 17365 19245 17395
rect 19275 17365 19280 17395
rect 19240 17360 19280 17365
rect 19320 17395 19360 17400
rect 19320 17365 19325 17395
rect 19355 17365 19360 17395
rect 19320 17360 19360 17365
rect 19400 17395 19440 17400
rect 19400 17365 19405 17395
rect 19435 17365 19440 17395
rect 19400 17360 19440 17365
rect 19480 17395 19520 17400
rect 19480 17365 19485 17395
rect 19515 17365 19520 17395
rect 19480 17360 19520 17365
rect 19560 17395 19600 17400
rect 19560 17365 19565 17395
rect 19595 17365 19600 17395
rect 19560 17360 19600 17365
rect 19640 17395 19680 17400
rect 19640 17365 19645 17395
rect 19675 17365 19680 17395
rect 19640 17360 19680 17365
rect 19720 17395 19760 17400
rect 19720 17365 19725 17395
rect 19755 17365 19760 17395
rect 19720 17360 19760 17365
rect 19800 17395 19840 17400
rect 19800 17365 19805 17395
rect 19835 17365 19840 17395
rect 19800 17360 19840 17365
rect 19880 17395 19920 17400
rect 19880 17365 19885 17395
rect 19915 17365 19920 17395
rect 19880 17360 19920 17365
rect 19960 17395 20000 17400
rect 19960 17365 19965 17395
rect 19995 17365 20000 17395
rect 19960 17360 20000 17365
rect 20040 17395 20080 17400
rect 20040 17365 20045 17395
rect 20075 17365 20080 17395
rect 20040 17360 20080 17365
rect 20120 17395 20160 17400
rect 20120 17365 20125 17395
rect 20155 17365 20160 17395
rect 20120 17360 20160 17365
rect 20200 17395 20240 17400
rect 20200 17365 20205 17395
rect 20235 17365 20240 17395
rect 20200 17360 20240 17365
rect 20280 17395 20320 17400
rect 20280 17365 20285 17395
rect 20315 17365 20320 17395
rect 20280 17360 20320 17365
rect 20360 17395 20400 17400
rect 20360 17365 20365 17395
rect 20395 17365 20400 17395
rect 20360 17360 20400 17365
rect 20440 17395 20480 17400
rect 20440 17365 20445 17395
rect 20475 17365 20480 17395
rect 20440 17360 20480 17365
rect 20520 17395 20560 17400
rect 20520 17365 20525 17395
rect 20555 17365 20560 17395
rect 20520 17360 20560 17365
rect 20600 17395 20640 17400
rect 20600 17365 20605 17395
rect 20635 17365 20640 17395
rect 20600 17360 20640 17365
rect 20680 17395 20720 17400
rect 20680 17365 20685 17395
rect 20715 17365 20720 17395
rect 20680 17360 20720 17365
rect 20760 17395 20800 17400
rect 20760 17365 20765 17395
rect 20795 17365 20800 17395
rect 20760 17360 20800 17365
rect 20840 17395 20880 17400
rect 20840 17365 20845 17395
rect 20875 17365 20880 17395
rect 20840 17360 20880 17365
rect 20920 17395 20960 17400
rect 20920 17365 20925 17395
rect 20955 17365 20960 17395
rect 20920 17360 20960 17365
rect 0 17235 40 17240
rect 0 17205 5 17235
rect 35 17205 40 17235
rect 0 17200 40 17205
rect 80 17235 120 17240
rect 80 17205 85 17235
rect 115 17205 120 17235
rect 80 17200 120 17205
rect 160 17235 200 17240
rect 160 17205 165 17235
rect 195 17205 200 17235
rect 160 17200 200 17205
rect 240 17235 280 17240
rect 240 17205 245 17235
rect 275 17205 280 17235
rect 240 17200 280 17205
rect 320 17235 360 17240
rect 320 17205 325 17235
rect 355 17205 360 17235
rect 320 17200 360 17205
rect 400 17235 440 17240
rect 400 17205 405 17235
rect 435 17205 440 17235
rect 400 17200 440 17205
rect 480 17235 520 17240
rect 480 17205 485 17235
rect 515 17205 520 17235
rect 480 17200 520 17205
rect 560 17235 600 17240
rect 560 17205 565 17235
rect 595 17205 600 17235
rect 560 17200 600 17205
rect 640 17235 680 17240
rect 640 17205 645 17235
rect 675 17205 680 17235
rect 640 17200 680 17205
rect 720 17235 760 17240
rect 720 17205 725 17235
rect 755 17205 760 17235
rect 720 17200 760 17205
rect 800 17235 840 17240
rect 800 17205 805 17235
rect 835 17205 840 17235
rect 800 17200 840 17205
rect 880 17235 920 17240
rect 880 17205 885 17235
rect 915 17205 920 17235
rect 880 17200 920 17205
rect 960 17235 1000 17240
rect 960 17205 965 17235
rect 995 17205 1000 17235
rect 960 17200 1000 17205
rect 1040 17235 1080 17240
rect 1040 17205 1045 17235
rect 1075 17205 1080 17235
rect 1040 17200 1080 17205
rect 1120 17235 1160 17240
rect 1120 17205 1125 17235
rect 1155 17205 1160 17235
rect 1120 17200 1160 17205
rect 1200 17235 1240 17240
rect 1200 17205 1205 17235
rect 1235 17205 1240 17235
rect 1200 17200 1240 17205
rect 1280 17235 1320 17240
rect 1280 17205 1285 17235
rect 1315 17205 1320 17235
rect 1280 17200 1320 17205
rect 1360 17235 1400 17240
rect 1360 17205 1365 17235
rect 1395 17205 1400 17235
rect 1360 17200 1400 17205
rect 1440 17235 1480 17240
rect 1440 17205 1445 17235
rect 1475 17205 1480 17235
rect 1440 17200 1480 17205
rect 1520 17235 1560 17240
rect 1520 17205 1525 17235
rect 1555 17205 1560 17235
rect 1520 17200 1560 17205
rect 1600 17235 1640 17240
rect 1600 17205 1605 17235
rect 1635 17205 1640 17235
rect 1600 17200 1640 17205
rect 1680 17235 1720 17240
rect 1680 17205 1685 17235
rect 1715 17205 1720 17235
rect 1680 17200 1720 17205
rect 1760 17235 1800 17240
rect 1760 17205 1765 17235
rect 1795 17205 1800 17235
rect 1760 17200 1800 17205
rect 1840 17235 1880 17240
rect 1840 17205 1845 17235
rect 1875 17205 1880 17235
rect 1840 17200 1880 17205
rect 1920 17235 1960 17240
rect 1920 17205 1925 17235
rect 1955 17205 1960 17235
rect 1920 17200 1960 17205
rect 2000 17235 2040 17240
rect 2000 17205 2005 17235
rect 2035 17205 2040 17235
rect 2000 17200 2040 17205
rect 2080 17235 2120 17240
rect 2080 17205 2085 17235
rect 2115 17205 2120 17235
rect 2080 17200 2120 17205
rect 2160 17235 2200 17240
rect 2160 17205 2165 17235
rect 2195 17205 2200 17235
rect 2160 17200 2200 17205
rect 2240 17235 2280 17240
rect 2240 17205 2245 17235
rect 2275 17205 2280 17235
rect 2240 17200 2280 17205
rect 2320 17235 2360 17240
rect 2320 17205 2325 17235
rect 2355 17205 2360 17235
rect 2320 17200 2360 17205
rect 2400 17235 2440 17240
rect 2400 17205 2405 17235
rect 2435 17205 2440 17235
rect 2400 17200 2440 17205
rect 2480 17235 2520 17240
rect 2480 17205 2485 17235
rect 2515 17205 2520 17235
rect 2480 17200 2520 17205
rect 2560 17235 2600 17240
rect 2560 17205 2565 17235
rect 2595 17205 2600 17235
rect 2560 17200 2600 17205
rect 2640 17235 2680 17240
rect 2640 17205 2645 17235
rect 2675 17205 2680 17235
rect 2640 17200 2680 17205
rect 2720 17235 2760 17240
rect 2720 17205 2725 17235
rect 2755 17205 2760 17235
rect 2720 17200 2760 17205
rect 2800 17235 2840 17240
rect 2800 17205 2805 17235
rect 2835 17205 2840 17235
rect 2800 17200 2840 17205
rect 2880 17235 2920 17240
rect 2880 17205 2885 17235
rect 2915 17205 2920 17235
rect 2880 17200 2920 17205
rect 2960 17235 3000 17240
rect 2960 17205 2965 17235
rect 2995 17205 3000 17235
rect 2960 17200 3000 17205
rect 3040 17235 3080 17240
rect 3040 17205 3045 17235
rect 3075 17205 3080 17235
rect 3040 17200 3080 17205
rect 3120 17235 3160 17240
rect 3120 17205 3125 17235
rect 3155 17205 3160 17235
rect 3120 17200 3160 17205
rect 3200 17235 3240 17240
rect 3200 17205 3205 17235
rect 3235 17205 3240 17235
rect 3200 17200 3240 17205
rect 3280 17235 3320 17240
rect 3280 17205 3285 17235
rect 3315 17205 3320 17235
rect 3280 17200 3320 17205
rect 3360 17235 3400 17240
rect 3360 17205 3365 17235
rect 3395 17205 3400 17235
rect 3360 17200 3400 17205
rect 3440 17235 3480 17240
rect 3440 17205 3445 17235
rect 3475 17205 3480 17235
rect 3440 17200 3480 17205
rect 3520 17235 3560 17240
rect 3520 17205 3525 17235
rect 3555 17205 3560 17235
rect 3520 17200 3560 17205
rect 3600 17235 3640 17240
rect 3600 17205 3605 17235
rect 3635 17205 3640 17235
rect 3600 17200 3640 17205
rect 3680 17235 3720 17240
rect 3680 17205 3685 17235
rect 3715 17205 3720 17235
rect 3680 17200 3720 17205
rect 3760 17235 3800 17240
rect 3760 17205 3765 17235
rect 3795 17205 3800 17235
rect 3760 17200 3800 17205
rect 3840 17235 3880 17240
rect 3840 17205 3845 17235
rect 3875 17205 3880 17235
rect 3840 17200 3880 17205
rect 3920 17235 3960 17240
rect 3920 17205 3925 17235
rect 3955 17205 3960 17235
rect 3920 17200 3960 17205
rect 4000 17235 4040 17240
rect 4000 17205 4005 17235
rect 4035 17205 4040 17235
rect 4000 17200 4040 17205
rect 4080 17235 4120 17240
rect 4080 17205 4085 17235
rect 4115 17205 4120 17235
rect 4080 17200 4120 17205
rect 4160 17235 4200 17240
rect 4160 17205 4165 17235
rect 4195 17205 4200 17235
rect 4160 17200 4200 17205
rect 6240 17235 6280 17240
rect 6240 17205 6245 17235
rect 6275 17205 6280 17235
rect 6240 17200 6280 17205
rect 6320 17235 6360 17240
rect 6320 17205 6325 17235
rect 6355 17205 6360 17235
rect 6320 17200 6360 17205
rect 6400 17235 6440 17240
rect 6400 17205 6405 17235
rect 6435 17205 6440 17235
rect 6400 17200 6440 17205
rect 6480 17235 6520 17240
rect 6480 17205 6485 17235
rect 6515 17205 6520 17235
rect 6480 17200 6520 17205
rect 6560 17235 6600 17240
rect 6560 17205 6565 17235
rect 6595 17205 6600 17235
rect 6560 17200 6600 17205
rect 6640 17235 6680 17240
rect 6640 17205 6645 17235
rect 6675 17205 6680 17235
rect 6640 17200 6680 17205
rect 6720 17235 6760 17240
rect 6720 17205 6725 17235
rect 6755 17205 6760 17235
rect 6720 17200 6760 17205
rect 6800 17235 6840 17240
rect 6800 17205 6805 17235
rect 6835 17205 6840 17235
rect 6800 17200 6840 17205
rect 6880 17235 6920 17240
rect 6880 17205 6885 17235
rect 6915 17205 6920 17235
rect 6880 17200 6920 17205
rect 6960 17235 7000 17240
rect 6960 17205 6965 17235
rect 6995 17205 7000 17235
rect 6960 17200 7000 17205
rect 7040 17235 7080 17240
rect 7040 17205 7045 17235
rect 7075 17205 7080 17235
rect 7040 17200 7080 17205
rect 7120 17235 7160 17240
rect 7120 17205 7125 17235
rect 7155 17205 7160 17235
rect 7120 17200 7160 17205
rect 7200 17235 7240 17240
rect 7200 17205 7205 17235
rect 7235 17205 7240 17235
rect 7200 17200 7240 17205
rect 7280 17235 7320 17240
rect 7280 17205 7285 17235
rect 7315 17205 7320 17235
rect 7280 17200 7320 17205
rect 7360 17235 7400 17240
rect 7360 17205 7365 17235
rect 7395 17205 7400 17235
rect 7360 17200 7400 17205
rect 7440 17235 7480 17240
rect 7440 17205 7445 17235
rect 7475 17205 7480 17235
rect 7440 17200 7480 17205
rect 7520 17235 7560 17240
rect 7520 17205 7525 17235
rect 7555 17205 7560 17235
rect 7520 17200 7560 17205
rect 7600 17235 7640 17240
rect 7600 17205 7605 17235
rect 7635 17205 7640 17235
rect 7600 17200 7640 17205
rect 7680 17235 7720 17240
rect 7680 17205 7685 17235
rect 7715 17205 7720 17235
rect 7680 17200 7720 17205
rect 7760 17235 7800 17240
rect 7760 17205 7765 17235
rect 7795 17205 7800 17235
rect 7760 17200 7800 17205
rect 7840 17235 7880 17240
rect 7840 17205 7845 17235
rect 7875 17205 7880 17235
rect 7840 17200 7880 17205
rect 7920 17235 7960 17240
rect 7920 17205 7925 17235
rect 7955 17205 7960 17235
rect 7920 17200 7960 17205
rect 8000 17235 8040 17240
rect 8000 17205 8005 17235
rect 8035 17205 8040 17235
rect 8000 17200 8040 17205
rect 8080 17235 8120 17240
rect 8080 17205 8085 17235
rect 8115 17205 8120 17235
rect 8080 17200 8120 17205
rect 8160 17235 8200 17240
rect 8160 17205 8165 17235
rect 8195 17205 8200 17235
rect 8160 17200 8200 17205
rect 8240 17235 8280 17240
rect 8240 17205 8245 17235
rect 8275 17205 8280 17235
rect 8240 17200 8280 17205
rect 8320 17235 8360 17240
rect 8320 17205 8325 17235
rect 8355 17205 8360 17235
rect 8320 17200 8360 17205
rect 8400 17235 8440 17240
rect 8400 17205 8405 17235
rect 8435 17205 8440 17235
rect 8400 17200 8440 17205
rect 8480 17235 8520 17240
rect 8480 17205 8485 17235
rect 8515 17205 8520 17235
rect 8480 17200 8520 17205
rect 8560 17235 8600 17240
rect 8560 17205 8565 17235
rect 8595 17205 8600 17235
rect 8560 17200 8600 17205
rect 8640 17235 8680 17240
rect 8640 17205 8645 17235
rect 8675 17205 8680 17235
rect 8640 17200 8680 17205
rect 8720 17235 8760 17240
rect 8720 17205 8725 17235
rect 8755 17205 8760 17235
rect 8720 17200 8760 17205
rect 8800 17235 8840 17240
rect 8800 17205 8805 17235
rect 8835 17205 8840 17235
rect 8800 17200 8840 17205
rect 8880 17235 8920 17240
rect 8880 17205 8885 17235
rect 8915 17205 8920 17235
rect 8880 17200 8920 17205
rect 8960 17235 9000 17240
rect 8960 17205 8965 17235
rect 8995 17205 9000 17235
rect 8960 17200 9000 17205
rect 9040 17235 9080 17240
rect 9040 17205 9045 17235
rect 9075 17205 9080 17235
rect 9040 17200 9080 17205
rect 9120 17235 9160 17240
rect 9120 17205 9125 17235
rect 9155 17205 9160 17235
rect 9120 17200 9160 17205
rect 9200 17235 9240 17240
rect 9200 17205 9205 17235
rect 9235 17205 9240 17235
rect 9200 17200 9240 17205
rect 9280 17235 9320 17240
rect 9280 17205 9285 17235
rect 9315 17205 9320 17235
rect 9280 17200 9320 17205
rect 9360 17235 9400 17240
rect 9360 17205 9365 17235
rect 9395 17205 9400 17235
rect 9360 17200 9400 17205
rect 9440 17235 9480 17240
rect 9440 17205 9445 17235
rect 9475 17205 9480 17235
rect 9440 17200 9480 17205
rect 11560 17235 11600 17240
rect 11560 17205 11565 17235
rect 11595 17205 11600 17235
rect 11560 17200 11600 17205
rect 11640 17235 11680 17240
rect 11640 17205 11645 17235
rect 11675 17205 11680 17235
rect 11640 17200 11680 17205
rect 11720 17235 11760 17240
rect 11720 17205 11725 17235
rect 11755 17205 11760 17235
rect 11720 17200 11760 17205
rect 11800 17235 11840 17240
rect 11800 17205 11805 17235
rect 11835 17205 11840 17235
rect 11800 17200 11840 17205
rect 11880 17235 11920 17240
rect 11880 17205 11885 17235
rect 11915 17205 11920 17235
rect 11880 17200 11920 17205
rect 11960 17235 12000 17240
rect 11960 17205 11965 17235
rect 11995 17205 12000 17235
rect 11960 17200 12000 17205
rect 12040 17235 12080 17240
rect 12040 17205 12045 17235
rect 12075 17205 12080 17235
rect 12040 17200 12080 17205
rect 12120 17235 12160 17240
rect 12120 17205 12125 17235
rect 12155 17205 12160 17235
rect 12120 17200 12160 17205
rect 12200 17235 12240 17240
rect 12200 17205 12205 17235
rect 12235 17205 12240 17235
rect 12200 17200 12240 17205
rect 12280 17235 12320 17240
rect 12280 17205 12285 17235
rect 12315 17205 12320 17235
rect 12280 17200 12320 17205
rect 12360 17235 12400 17240
rect 12360 17205 12365 17235
rect 12395 17205 12400 17235
rect 12360 17200 12400 17205
rect 12440 17235 12480 17240
rect 12440 17205 12445 17235
rect 12475 17205 12480 17235
rect 12440 17200 12480 17205
rect 12520 17235 12560 17240
rect 12520 17205 12525 17235
rect 12555 17205 12560 17235
rect 12520 17200 12560 17205
rect 12600 17235 12640 17240
rect 12600 17205 12605 17235
rect 12635 17205 12640 17235
rect 12600 17200 12640 17205
rect 12680 17235 12720 17240
rect 12680 17205 12685 17235
rect 12715 17205 12720 17235
rect 12680 17200 12720 17205
rect 12760 17235 12800 17240
rect 12760 17205 12765 17235
rect 12795 17205 12800 17235
rect 12760 17200 12800 17205
rect 12840 17235 12880 17240
rect 12840 17205 12845 17235
rect 12875 17205 12880 17235
rect 12840 17200 12880 17205
rect 12920 17235 12960 17240
rect 12920 17205 12925 17235
rect 12955 17205 12960 17235
rect 12920 17200 12960 17205
rect 13000 17235 13040 17240
rect 13000 17205 13005 17235
rect 13035 17205 13040 17235
rect 13000 17200 13040 17205
rect 13080 17235 13120 17240
rect 13080 17205 13085 17235
rect 13115 17205 13120 17235
rect 13080 17200 13120 17205
rect 13160 17235 13200 17240
rect 13160 17205 13165 17235
rect 13195 17205 13200 17235
rect 13160 17200 13200 17205
rect 13240 17235 13280 17240
rect 13240 17205 13245 17235
rect 13275 17205 13280 17235
rect 13240 17200 13280 17205
rect 13320 17235 13360 17240
rect 13320 17205 13325 17235
rect 13355 17205 13360 17235
rect 13320 17200 13360 17205
rect 13400 17235 13440 17240
rect 13400 17205 13405 17235
rect 13435 17205 13440 17235
rect 13400 17200 13440 17205
rect 13480 17235 13520 17240
rect 13480 17205 13485 17235
rect 13515 17205 13520 17235
rect 13480 17200 13520 17205
rect 13560 17235 13600 17240
rect 13560 17205 13565 17235
rect 13595 17205 13600 17235
rect 13560 17200 13600 17205
rect 13640 17235 13680 17240
rect 13640 17205 13645 17235
rect 13675 17205 13680 17235
rect 13640 17200 13680 17205
rect 13720 17235 13760 17240
rect 13720 17205 13725 17235
rect 13755 17205 13760 17235
rect 13720 17200 13760 17205
rect 13800 17235 13840 17240
rect 13800 17205 13805 17235
rect 13835 17205 13840 17235
rect 13800 17200 13840 17205
rect 13880 17235 13920 17240
rect 13880 17205 13885 17235
rect 13915 17205 13920 17235
rect 13880 17200 13920 17205
rect 13960 17235 14000 17240
rect 13960 17205 13965 17235
rect 13995 17205 14000 17235
rect 13960 17200 14000 17205
rect 14040 17235 14080 17240
rect 14040 17205 14045 17235
rect 14075 17205 14080 17235
rect 14040 17200 14080 17205
rect 14120 17235 14160 17240
rect 14120 17205 14125 17235
rect 14155 17205 14160 17235
rect 14120 17200 14160 17205
rect 14200 17235 14240 17240
rect 14200 17205 14205 17235
rect 14235 17205 14240 17235
rect 14200 17200 14240 17205
rect 14280 17235 14320 17240
rect 14280 17205 14285 17235
rect 14315 17205 14320 17235
rect 14280 17200 14320 17205
rect 14360 17235 14400 17240
rect 14360 17205 14365 17235
rect 14395 17205 14400 17235
rect 14360 17200 14400 17205
rect 14440 17235 14480 17240
rect 14440 17205 14445 17235
rect 14475 17205 14480 17235
rect 14440 17200 14480 17205
rect 14520 17235 14560 17240
rect 14520 17205 14525 17235
rect 14555 17205 14560 17235
rect 14520 17200 14560 17205
rect 14600 17235 14640 17240
rect 14600 17205 14605 17235
rect 14635 17205 14640 17235
rect 14600 17200 14640 17205
rect 14680 17235 14720 17240
rect 14680 17205 14685 17235
rect 14715 17205 14720 17235
rect 14680 17200 14720 17205
rect 16760 17235 16800 17240
rect 16760 17205 16765 17235
rect 16795 17205 16800 17235
rect 16760 17200 16800 17205
rect 16840 17235 16880 17240
rect 16840 17205 16845 17235
rect 16875 17205 16880 17235
rect 16840 17200 16880 17205
rect 16920 17235 16960 17240
rect 16920 17205 16925 17235
rect 16955 17205 16960 17235
rect 16920 17200 16960 17205
rect 17000 17235 17040 17240
rect 17000 17205 17005 17235
rect 17035 17205 17040 17235
rect 17000 17200 17040 17205
rect 17080 17235 17120 17240
rect 17080 17205 17085 17235
rect 17115 17205 17120 17235
rect 17080 17200 17120 17205
rect 17160 17235 17200 17240
rect 17160 17205 17165 17235
rect 17195 17205 17200 17235
rect 17160 17200 17200 17205
rect 17240 17235 17280 17240
rect 17240 17205 17245 17235
rect 17275 17205 17280 17235
rect 17240 17200 17280 17205
rect 17320 17235 17360 17240
rect 17320 17205 17325 17235
rect 17355 17205 17360 17235
rect 17320 17200 17360 17205
rect 17400 17235 17440 17240
rect 17400 17205 17405 17235
rect 17435 17205 17440 17235
rect 17400 17200 17440 17205
rect 17480 17235 17520 17240
rect 17480 17205 17485 17235
rect 17515 17205 17520 17235
rect 17480 17200 17520 17205
rect 17560 17235 17600 17240
rect 17560 17205 17565 17235
rect 17595 17205 17600 17235
rect 17560 17200 17600 17205
rect 17640 17235 17680 17240
rect 17640 17205 17645 17235
rect 17675 17205 17680 17235
rect 17640 17200 17680 17205
rect 17720 17235 17760 17240
rect 17720 17205 17725 17235
rect 17755 17205 17760 17235
rect 17720 17200 17760 17205
rect 17800 17235 17840 17240
rect 17800 17205 17805 17235
rect 17835 17205 17840 17235
rect 17800 17200 17840 17205
rect 17880 17235 17920 17240
rect 17880 17205 17885 17235
rect 17915 17205 17920 17235
rect 17880 17200 17920 17205
rect 17960 17235 18000 17240
rect 17960 17205 17965 17235
rect 17995 17205 18000 17235
rect 17960 17200 18000 17205
rect 18040 17235 18080 17240
rect 18040 17205 18045 17235
rect 18075 17205 18080 17235
rect 18040 17200 18080 17205
rect 18120 17235 18160 17240
rect 18120 17205 18125 17235
rect 18155 17205 18160 17235
rect 18120 17200 18160 17205
rect 18200 17235 18240 17240
rect 18200 17205 18205 17235
rect 18235 17205 18240 17235
rect 18200 17200 18240 17205
rect 18280 17235 18320 17240
rect 18280 17205 18285 17235
rect 18315 17205 18320 17235
rect 18280 17200 18320 17205
rect 18360 17235 18400 17240
rect 18360 17205 18365 17235
rect 18395 17205 18400 17235
rect 18360 17200 18400 17205
rect 18440 17235 18480 17240
rect 18440 17205 18445 17235
rect 18475 17205 18480 17235
rect 18440 17200 18480 17205
rect 18520 17235 18560 17240
rect 18520 17205 18525 17235
rect 18555 17205 18560 17235
rect 18520 17200 18560 17205
rect 18600 17235 18640 17240
rect 18600 17205 18605 17235
rect 18635 17205 18640 17235
rect 18600 17200 18640 17205
rect 18680 17235 18720 17240
rect 18680 17205 18685 17235
rect 18715 17205 18720 17235
rect 18680 17200 18720 17205
rect 18760 17235 18800 17240
rect 18760 17205 18765 17235
rect 18795 17205 18800 17235
rect 18760 17200 18800 17205
rect 18840 17235 18880 17240
rect 18840 17205 18845 17235
rect 18875 17205 18880 17235
rect 18840 17200 18880 17205
rect 18920 17235 18960 17240
rect 18920 17205 18925 17235
rect 18955 17205 18960 17235
rect 18920 17200 18960 17205
rect 19000 17235 19040 17240
rect 19000 17205 19005 17235
rect 19035 17205 19040 17235
rect 19000 17200 19040 17205
rect 19080 17235 19120 17240
rect 19080 17205 19085 17235
rect 19115 17205 19120 17235
rect 19080 17200 19120 17205
rect 19160 17235 19200 17240
rect 19160 17205 19165 17235
rect 19195 17205 19200 17235
rect 19160 17200 19200 17205
rect 19240 17235 19280 17240
rect 19240 17205 19245 17235
rect 19275 17205 19280 17235
rect 19240 17200 19280 17205
rect 19320 17235 19360 17240
rect 19320 17205 19325 17235
rect 19355 17205 19360 17235
rect 19320 17200 19360 17205
rect 19400 17235 19440 17240
rect 19400 17205 19405 17235
rect 19435 17205 19440 17235
rect 19400 17200 19440 17205
rect 19480 17235 19520 17240
rect 19480 17205 19485 17235
rect 19515 17205 19520 17235
rect 19480 17200 19520 17205
rect 19560 17235 19600 17240
rect 19560 17205 19565 17235
rect 19595 17205 19600 17235
rect 19560 17200 19600 17205
rect 19640 17235 19680 17240
rect 19640 17205 19645 17235
rect 19675 17205 19680 17235
rect 19640 17200 19680 17205
rect 19720 17235 19760 17240
rect 19720 17205 19725 17235
rect 19755 17205 19760 17235
rect 19720 17200 19760 17205
rect 19800 17235 19840 17240
rect 19800 17205 19805 17235
rect 19835 17205 19840 17235
rect 19800 17200 19840 17205
rect 19880 17235 19920 17240
rect 19880 17205 19885 17235
rect 19915 17205 19920 17235
rect 19880 17200 19920 17205
rect 19960 17235 20000 17240
rect 19960 17205 19965 17235
rect 19995 17205 20000 17235
rect 19960 17200 20000 17205
rect 20040 17235 20080 17240
rect 20040 17205 20045 17235
rect 20075 17205 20080 17235
rect 20040 17200 20080 17205
rect 20120 17235 20160 17240
rect 20120 17205 20125 17235
rect 20155 17205 20160 17235
rect 20120 17200 20160 17205
rect 20200 17235 20240 17240
rect 20200 17205 20205 17235
rect 20235 17205 20240 17235
rect 20200 17200 20240 17205
rect 20280 17235 20320 17240
rect 20280 17205 20285 17235
rect 20315 17205 20320 17235
rect 20280 17200 20320 17205
rect 20360 17235 20400 17240
rect 20360 17205 20365 17235
rect 20395 17205 20400 17235
rect 20360 17200 20400 17205
rect 20440 17235 20480 17240
rect 20440 17205 20445 17235
rect 20475 17205 20480 17235
rect 20440 17200 20480 17205
rect 20520 17235 20560 17240
rect 20520 17205 20525 17235
rect 20555 17205 20560 17235
rect 20520 17200 20560 17205
rect 20600 17235 20640 17240
rect 20600 17205 20605 17235
rect 20635 17205 20640 17235
rect 20600 17200 20640 17205
rect 20680 17235 20720 17240
rect 20680 17205 20685 17235
rect 20715 17205 20720 17235
rect 20680 17200 20720 17205
rect 20760 17235 20800 17240
rect 20760 17205 20765 17235
rect 20795 17205 20800 17235
rect 20760 17200 20800 17205
rect 20840 17235 20880 17240
rect 20840 17205 20845 17235
rect 20875 17205 20880 17235
rect 20840 17200 20880 17205
rect 20920 17235 20960 17240
rect 20920 17205 20925 17235
rect 20955 17205 20960 17235
rect 20920 17200 20960 17205
rect 0 17155 40 17160
rect 0 17125 5 17155
rect 35 17125 40 17155
rect 0 17120 40 17125
rect 80 17155 120 17160
rect 80 17125 85 17155
rect 115 17125 120 17155
rect 80 17120 120 17125
rect 160 17155 200 17160
rect 160 17125 165 17155
rect 195 17125 200 17155
rect 160 17120 200 17125
rect 240 17155 280 17160
rect 240 17125 245 17155
rect 275 17125 280 17155
rect 240 17120 280 17125
rect 320 17155 360 17160
rect 320 17125 325 17155
rect 355 17125 360 17155
rect 320 17120 360 17125
rect 400 17155 440 17160
rect 400 17125 405 17155
rect 435 17125 440 17155
rect 400 17120 440 17125
rect 480 17155 520 17160
rect 480 17125 485 17155
rect 515 17125 520 17155
rect 480 17120 520 17125
rect 560 17155 600 17160
rect 560 17125 565 17155
rect 595 17125 600 17155
rect 560 17120 600 17125
rect 640 17155 680 17160
rect 640 17125 645 17155
rect 675 17125 680 17155
rect 640 17120 680 17125
rect 720 17155 760 17160
rect 720 17125 725 17155
rect 755 17125 760 17155
rect 720 17120 760 17125
rect 800 17155 840 17160
rect 800 17125 805 17155
rect 835 17125 840 17155
rect 800 17120 840 17125
rect 880 17155 920 17160
rect 880 17125 885 17155
rect 915 17125 920 17155
rect 880 17120 920 17125
rect 960 17155 1000 17160
rect 960 17125 965 17155
rect 995 17125 1000 17155
rect 960 17120 1000 17125
rect 1040 17155 1080 17160
rect 1040 17125 1045 17155
rect 1075 17125 1080 17155
rect 1040 17120 1080 17125
rect 1120 17155 1160 17160
rect 1120 17125 1125 17155
rect 1155 17125 1160 17155
rect 1120 17120 1160 17125
rect 1200 17155 1240 17160
rect 1200 17125 1205 17155
rect 1235 17125 1240 17155
rect 1200 17120 1240 17125
rect 1280 17155 1320 17160
rect 1280 17125 1285 17155
rect 1315 17125 1320 17155
rect 1280 17120 1320 17125
rect 1360 17155 1400 17160
rect 1360 17125 1365 17155
rect 1395 17125 1400 17155
rect 1360 17120 1400 17125
rect 1440 17155 1480 17160
rect 1440 17125 1445 17155
rect 1475 17125 1480 17155
rect 1440 17120 1480 17125
rect 1520 17155 1560 17160
rect 1520 17125 1525 17155
rect 1555 17125 1560 17155
rect 1520 17120 1560 17125
rect 1600 17155 1640 17160
rect 1600 17125 1605 17155
rect 1635 17125 1640 17155
rect 1600 17120 1640 17125
rect 1680 17155 1720 17160
rect 1680 17125 1685 17155
rect 1715 17125 1720 17155
rect 1680 17120 1720 17125
rect 1760 17155 1800 17160
rect 1760 17125 1765 17155
rect 1795 17125 1800 17155
rect 1760 17120 1800 17125
rect 1840 17155 1880 17160
rect 1840 17125 1845 17155
rect 1875 17125 1880 17155
rect 1840 17120 1880 17125
rect 1920 17155 1960 17160
rect 1920 17125 1925 17155
rect 1955 17125 1960 17155
rect 1920 17120 1960 17125
rect 2000 17155 2040 17160
rect 2000 17125 2005 17155
rect 2035 17125 2040 17155
rect 2000 17120 2040 17125
rect 2080 17155 2120 17160
rect 2080 17125 2085 17155
rect 2115 17125 2120 17155
rect 2080 17120 2120 17125
rect 2160 17155 2200 17160
rect 2160 17125 2165 17155
rect 2195 17125 2200 17155
rect 2160 17120 2200 17125
rect 2240 17155 2280 17160
rect 2240 17125 2245 17155
rect 2275 17125 2280 17155
rect 2240 17120 2280 17125
rect 2320 17155 2360 17160
rect 2320 17125 2325 17155
rect 2355 17125 2360 17155
rect 2320 17120 2360 17125
rect 2400 17155 2440 17160
rect 2400 17125 2405 17155
rect 2435 17125 2440 17155
rect 2400 17120 2440 17125
rect 2480 17155 2520 17160
rect 2480 17125 2485 17155
rect 2515 17125 2520 17155
rect 2480 17120 2520 17125
rect 2560 17155 2600 17160
rect 2560 17125 2565 17155
rect 2595 17125 2600 17155
rect 2560 17120 2600 17125
rect 2640 17155 2680 17160
rect 2640 17125 2645 17155
rect 2675 17125 2680 17155
rect 2640 17120 2680 17125
rect 2720 17155 2760 17160
rect 2720 17125 2725 17155
rect 2755 17125 2760 17155
rect 2720 17120 2760 17125
rect 2800 17155 2840 17160
rect 2800 17125 2805 17155
rect 2835 17125 2840 17155
rect 2800 17120 2840 17125
rect 2880 17155 2920 17160
rect 2880 17125 2885 17155
rect 2915 17125 2920 17155
rect 2880 17120 2920 17125
rect 2960 17155 3000 17160
rect 2960 17125 2965 17155
rect 2995 17125 3000 17155
rect 2960 17120 3000 17125
rect 3040 17155 3080 17160
rect 3040 17125 3045 17155
rect 3075 17125 3080 17155
rect 3040 17120 3080 17125
rect 3120 17155 3160 17160
rect 3120 17125 3125 17155
rect 3155 17125 3160 17155
rect 3120 17120 3160 17125
rect 3200 17155 3240 17160
rect 3200 17125 3205 17155
rect 3235 17125 3240 17155
rect 3200 17120 3240 17125
rect 3280 17155 3320 17160
rect 3280 17125 3285 17155
rect 3315 17125 3320 17155
rect 3280 17120 3320 17125
rect 3360 17155 3400 17160
rect 3360 17125 3365 17155
rect 3395 17125 3400 17155
rect 3360 17120 3400 17125
rect 3440 17155 3480 17160
rect 3440 17125 3445 17155
rect 3475 17125 3480 17155
rect 3440 17120 3480 17125
rect 3520 17155 3560 17160
rect 3520 17125 3525 17155
rect 3555 17125 3560 17155
rect 3520 17120 3560 17125
rect 3600 17155 3640 17160
rect 3600 17125 3605 17155
rect 3635 17125 3640 17155
rect 3600 17120 3640 17125
rect 3680 17155 3720 17160
rect 3680 17125 3685 17155
rect 3715 17125 3720 17155
rect 3680 17120 3720 17125
rect 3760 17155 3800 17160
rect 3760 17125 3765 17155
rect 3795 17125 3800 17155
rect 3760 17120 3800 17125
rect 3840 17155 3880 17160
rect 3840 17125 3845 17155
rect 3875 17125 3880 17155
rect 3840 17120 3880 17125
rect 3920 17155 3960 17160
rect 3920 17125 3925 17155
rect 3955 17125 3960 17155
rect 3920 17120 3960 17125
rect 4000 17155 4040 17160
rect 4000 17125 4005 17155
rect 4035 17125 4040 17155
rect 4000 17120 4040 17125
rect 4080 17155 4120 17160
rect 4080 17125 4085 17155
rect 4115 17125 4120 17155
rect 4080 17120 4120 17125
rect 4160 17155 4200 17160
rect 4160 17125 4165 17155
rect 4195 17125 4200 17155
rect 4160 17120 4200 17125
rect 6240 17155 6280 17160
rect 6240 17125 6245 17155
rect 6275 17125 6280 17155
rect 6240 17120 6280 17125
rect 6320 17155 6360 17160
rect 6320 17125 6325 17155
rect 6355 17125 6360 17155
rect 6320 17120 6360 17125
rect 6400 17155 6440 17160
rect 6400 17125 6405 17155
rect 6435 17125 6440 17155
rect 6400 17120 6440 17125
rect 6480 17155 6520 17160
rect 6480 17125 6485 17155
rect 6515 17125 6520 17155
rect 6480 17120 6520 17125
rect 6560 17155 6600 17160
rect 6560 17125 6565 17155
rect 6595 17125 6600 17155
rect 6560 17120 6600 17125
rect 6640 17155 6680 17160
rect 6640 17125 6645 17155
rect 6675 17125 6680 17155
rect 6640 17120 6680 17125
rect 6720 17155 6760 17160
rect 6720 17125 6725 17155
rect 6755 17125 6760 17155
rect 6720 17120 6760 17125
rect 6800 17155 6840 17160
rect 6800 17125 6805 17155
rect 6835 17125 6840 17155
rect 6800 17120 6840 17125
rect 6880 17155 6920 17160
rect 6880 17125 6885 17155
rect 6915 17125 6920 17155
rect 6880 17120 6920 17125
rect 6960 17155 7000 17160
rect 6960 17125 6965 17155
rect 6995 17125 7000 17155
rect 6960 17120 7000 17125
rect 7040 17155 7080 17160
rect 7040 17125 7045 17155
rect 7075 17125 7080 17155
rect 7040 17120 7080 17125
rect 7120 17155 7160 17160
rect 7120 17125 7125 17155
rect 7155 17125 7160 17155
rect 7120 17120 7160 17125
rect 7200 17155 7240 17160
rect 7200 17125 7205 17155
rect 7235 17125 7240 17155
rect 7200 17120 7240 17125
rect 7280 17155 7320 17160
rect 7280 17125 7285 17155
rect 7315 17125 7320 17155
rect 7280 17120 7320 17125
rect 7360 17155 7400 17160
rect 7360 17125 7365 17155
rect 7395 17125 7400 17155
rect 7360 17120 7400 17125
rect 7440 17155 7480 17160
rect 7440 17125 7445 17155
rect 7475 17125 7480 17155
rect 7440 17120 7480 17125
rect 7520 17155 7560 17160
rect 7520 17125 7525 17155
rect 7555 17125 7560 17155
rect 7520 17120 7560 17125
rect 7600 17155 7640 17160
rect 7600 17125 7605 17155
rect 7635 17125 7640 17155
rect 7600 17120 7640 17125
rect 7680 17155 7720 17160
rect 7680 17125 7685 17155
rect 7715 17125 7720 17155
rect 7680 17120 7720 17125
rect 7760 17155 7800 17160
rect 7760 17125 7765 17155
rect 7795 17125 7800 17155
rect 7760 17120 7800 17125
rect 7840 17155 7880 17160
rect 7840 17125 7845 17155
rect 7875 17125 7880 17155
rect 7840 17120 7880 17125
rect 7920 17155 7960 17160
rect 7920 17125 7925 17155
rect 7955 17125 7960 17155
rect 7920 17120 7960 17125
rect 8000 17155 8040 17160
rect 8000 17125 8005 17155
rect 8035 17125 8040 17155
rect 8000 17120 8040 17125
rect 8080 17155 8120 17160
rect 8080 17125 8085 17155
rect 8115 17125 8120 17155
rect 8080 17120 8120 17125
rect 8160 17155 8200 17160
rect 8160 17125 8165 17155
rect 8195 17125 8200 17155
rect 8160 17120 8200 17125
rect 8240 17155 8280 17160
rect 8240 17125 8245 17155
rect 8275 17125 8280 17155
rect 8240 17120 8280 17125
rect 8320 17155 8360 17160
rect 8320 17125 8325 17155
rect 8355 17125 8360 17155
rect 8320 17120 8360 17125
rect 8400 17155 8440 17160
rect 8400 17125 8405 17155
rect 8435 17125 8440 17155
rect 8400 17120 8440 17125
rect 8480 17155 8520 17160
rect 8480 17125 8485 17155
rect 8515 17125 8520 17155
rect 8480 17120 8520 17125
rect 8560 17155 8600 17160
rect 8560 17125 8565 17155
rect 8595 17125 8600 17155
rect 8560 17120 8600 17125
rect 8640 17155 8680 17160
rect 8640 17125 8645 17155
rect 8675 17125 8680 17155
rect 8640 17120 8680 17125
rect 8720 17155 8760 17160
rect 8720 17125 8725 17155
rect 8755 17125 8760 17155
rect 8720 17120 8760 17125
rect 8800 17155 8840 17160
rect 8800 17125 8805 17155
rect 8835 17125 8840 17155
rect 8800 17120 8840 17125
rect 8880 17155 8920 17160
rect 8880 17125 8885 17155
rect 8915 17125 8920 17155
rect 8880 17120 8920 17125
rect 8960 17155 9000 17160
rect 8960 17125 8965 17155
rect 8995 17125 9000 17155
rect 8960 17120 9000 17125
rect 9040 17155 9080 17160
rect 9040 17125 9045 17155
rect 9075 17125 9080 17155
rect 9040 17120 9080 17125
rect 9120 17155 9160 17160
rect 9120 17125 9125 17155
rect 9155 17125 9160 17155
rect 9120 17120 9160 17125
rect 9200 17155 9240 17160
rect 9200 17125 9205 17155
rect 9235 17125 9240 17155
rect 9200 17120 9240 17125
rect 9280 17155 9320 17160
rect 9280 17125 9285 17155
rect 9315 17125 9320 17155
rect 9280 17120 9320 17125
rect 9360 17155 9400 17160
rect 9360 17125 9365 17155
rect 9395 17125 9400 17155
rect 9360 17120 9400 17125
rect 9440 17155 9480 17160
rect 9440 17125 9445 17155
rect 9475 17125 9480 17155
rect 9440 17120 9480 17125
rect 11560 17155 11600 17160
rect 11560 17125 11565 17155
rect 11595 17125 11600 17155
rect 11560 17120 11600 17125
rect 11640 17155 11680 17160
rect 11640 17125 11645 17155
rect 11675 17125 11680 17155
rect 11640 17120 11680 17125
rect 11720 17155 11760 17160
rect 11720 17125 11725 17155
rect 11755 17125 11760 17155
rect 11720 17120 11760 17125
rect 11800 17155 11840 17160
rect 11800 17125 11805 17155
rect 11835 17125 11840 17155
rect 11800 17120 11840 17125
rect 11880 17155 11920 17160
rect 11880 17125 11885 17155
rect 11915 17125 11920 17155
rect 11880 17120 11920 17125
rect 11960 17155 12000 17160
rect 11960 17125 11965 17155
rect 11995 17125 12000 17155
rect 11960 17120 12000 17125
rect 12040 17155 12080 17160
rect 12040 17125 12045 17155
rect 12075 17125 12080 17155
rect 12040 17120 12080 17125
rect 12120 17155 12160 17160
rect 12120 17125 12125 17155
rect 12155 17125 12160 17155
rect 12120 17120 12160 17125
rect 12200 17155 12240 17160
rect 12200 17125 12205 17155
rect 12235 17125 12240 17155
rect 12200 17120 12240 17125
rect 12280 17155 12320 17160
rect 12280 17125 12285 17155
rect 12315 17125 12320 17155
rect 12280 17120 12320 17125
rect 12360 17155 12400 17160
rect 12360 17125 12365 17155
rect 12395 17125 12400 17155
rect 12360 17120 12400 17125
rect 12440 17155 12480 17160
rect 12440 17125 12445 17155
rect 12475 17125 12480 17155
rect 12440 17120 12480 17125
rect 12520 17155 12560 17160
rect 12520 17125 12525 17155
rect 12555 17125 12560 17155
rect 12520 17120 12560 17125
rect 12600 17155 12640 17160
rect 12600 17125 12605 17155
rect 12635 17125 12640 17155
rect 12600 17120 12640 17125
rect 12680 17155 12720 17160
rect 12680 17125 12685 17155
rect 12715 17125 12720 17155
rect 12680 17120 12720 17125
rect 12760 17155 12800 17160
rect 12760 17125 12765 17155
rect 12795 17125 12800 17155
rect 12760 17120 12800 17125
rect 12840 17155 12880 17160
rect 12840 17125 12845 17155
rect 12875 17125 12880 17155
rect 12840 17120 12880 17125
rect 12920 17155 12960 17160
rect 12920 17125 12925 17155
rect 12955 17125 12960 17155
rect 12920 17120 12960 17125
rect 13000 17155 13040 17160
rect 13000 17125 13005 17155
rect 13035 17125 13040 17155
rect 13000 17120 13040 17125
rect 13080 17155 13120 17160
rect 13080 17125 13085 17155
rect 13115 17125 13120 17155
rect 13080 17120 13120 17125
rect 13160 17155 13200 17160
rect 13160 17125 13165 17155
rect 13195 17125 13200 17155
rect 13160 17120 13200 17125
rect 13240 17155 13280 17160
rect 13240 17125 13245 17155
rect 13275 17125 13280 17155
rect 13240 17120 13280 17125
rect 13320 17155 13360 17160
rect 13320 17125 13325 17155
rect 13355 17125 13360 17155
rect 13320 17120 13360 17125
rect 13400 17155 13440 17160
rect 13400 17125 13405 17155
rect 13435 17125 13440 17155
rect 13400 17120 13440 17125
rect 13480 17155 13520 17160
rect 13480 17125 13485 17155
rect 13515 17125 13520 17155
rect 13480 17120 13520 17125
rect 13560 17155 13600 17160
rect 13560 17125 13565 17155
rect 13595 17125 13600 17155
rect 13560 17120 13600 17125
rect 13640 17155 13680 17160
rect 13640 17125 13645 17155
rect 13675 17125 13680 17155
rect 13640 17120 13680 17125
rect 13720 17155 13760 17160
rect 13720 17125 13725 17155
rect 13755 17125 13760 17155
rect 13720 17120 13760 17125
rect 13800 17155 13840 17160
rect 13800 17125 13805 17155
rect 13835 17125 13840 17155
rect 13800 17120 13840 17125
rect 13880 17155 13920 17160
rect 13880 17125 13885 17155
rect 13915 17125 13920 17155
rect 13880 17120 13920 17125
rect 13960 17155 14000 17160
rect 13960 17125 13965 17155
rect 13995 17125 14000 17155
rect 13960 17120 14000 17125
rect 14040 17155 14080 17160
rect 14040 17125 14045 17155
rect 14075 17125 14080 17155
rect 14040 17120 14080 17125
rect 14120 17155 14160 17160
rect 14120 17125 14125 17155
rect 14155 17125 14160 17155
rect 14120 17120 14160 17125
rect 14200 17155 14240 17160
rect 14200 17125 14205 17155
rect 14235 17125 14240 17155
rect 14200 17120 14240 17125
rect 14280 17155 14320 17160
rect 14280 17125 14285 17155
rect 14315 17125 14320 17155
rect 14280 17120 14320 17125
rect 14360 17155 14400 17160
rect 14360 17125 14365 17155
rect 14395 17125 14400 17155
rect 14360 17120 14400 17125
rect 14440 17155 14480 17160
rect 14440 17125 14445 17155
rect 14475 17125 14480 17155
rect 14440 17120 14480 17125
rect 14520 17155 14560 17160
rect 14520 17125 14525 17155
rect 14555 17125 14560 17155
rect 14520 17120 14560 17125
rect 14600 17155 14640 17160
rect 14600 17125 14605 17155
rect 14635 17125 14640 17155
rect 14600 17120 14640 17125
rect 14680 17155 14720 17160
rect 14680 17125 14685 17155
rect 14715 17125 14720 17155
rect 14680 17120 14720 17125
rect 16760 17155 16800 17160
rect 16760 17125 16765 17155
rect 16795 17125 16800 17155
rect 16760 17120 16800 17125
rect 16840 17155 16880 17160
rect 16840 17125 16845 17155
rect 16875 17125 16880 17155
rect 16840 17120 16880 17125
rect 16920 17155 16960 17160
rect 16920 17125 16925 17155
rect 16955 17125 16960 17155
rect 16920 17120 16960 17125
rect 17000 17155 17040 17160
rect 17000 17125 17005 17155
rect 17035 17125 17040 17155
rect 17000 17120 17040 17125
rect 17080 17155 17120 17160
rect 17080 17125 17085 17155
rect 17115 17125 17120 17155
rect 17080 17120 17120 17125
rect 17160 17155 17200 17160
rect 17160 17125 17165 17155
rect 17195 17125 17200 17155
rect 17160 17120 17200 17125
rect 17240 17155 17280 17160
rect 17240 17125 17245 17155
rect 17275 17125 17280 17155
rect 17240 17120 17280 17125
rect 17320 17155 17360 17160
rect 17320 17125 17325 17155
rect 17355 17125 17360 17155
rect 17320 17120 17360 17125
rect 17400 17155 17440 17160
rect 17400 17125 17405 17155
rect 17435 17125 17440 17155
rect 17400 17120 17440 17125
rect 17480 17155 17520 17160
rect 17480 17125 17485 17155
rect 17515 17125 17520 17155
rect 17480 17120 17520 17125
rect 17560 17155 17600 17160
rect 17560 17125 17565 17155
rect 17595 17125 17600 17155
rect 17560 17120 17600 17125
rect 17640 17155 17680 17160
rect 17640 17125 17645 17155
rect 17675 17125 17680 17155
rect 17640 17120 17680 17125
rect 17720 17155 17760 17160
rect 17720 17125 17725 17155
rect 17755 17125 17760 17155
rect 17720 17120 17760 17125
rect 17800 17155 17840 17160
rect 17800 17125 17805 17155
rect 17835 17125 17840 17155
rect 17800 17120 17840 17125
rect 17880 17155 17920 17160
rect 17880 17125 17885 17155
rect 17915 17125 17920 17155
rect 17880 17120 17920 17125
rect 17960 17155 18000 17160
rect 17960 17125 17965 17155
rect 17995 17125 18000 17155
rect 17960 17120 18000 17125
rect 18040 17155 18080 17160
rect 18040 17125 18045 17155
rect 18075 17125 18080 17155
rect 18040 17120 18080 17125
rect 18120 17155 18160 17160
rect 18120 17125 18125 17155
rect 18155 17125 18160 17155
rect 18120 17120 18160 17125
rect 18200 17155 18240 17160
rect 18200 17125 18205 17155
rect 18235 17125 18240 17155
rect 18200 17120 18240 17125
rect 18280 17155 18320 17160
rect 18280 17125 18285 17155
rect 18315 17125 18320 17155
rect 18280 17120 18320 17125
rect 18360 17155 18400 17160
rect 18360 17125 18365 17155
rect 18395 17125 18400 17155
rect 18360 17120 18400 17125
rect 18440 17155 18480 17160
rect 18440 17125 18445 17155
rect 18475 17125 18480 17155
rect 18440 17120 18480 17125
rect 18520 17155 18560 17160
rect 18520 17125 18525 17155
rect 18555 17125 18560 17155
rect 18520 17120 18560 17125
rect 18600 17155 18640 17160
rect 18600 17125 18605 17155
rect 18635 17125 18640 17155
rect 18600 17120 18640 17125
rect 18680 17155 18720 17160
rect 18680 17125 18685 17155
rect 18715 17125 18720 17155
rect 18680 17120 18720 17125
rect 18760 17155 18800 17160
rect 18760 17125 18765 17155
rect 18795 17125 18800 17155
rect 18760 17120 18800 17125
rect 18840 17155 18880 17160
rect 18840 17125 18845 17155
rect 18875 17125 18880 17155
rect 18840 17120 18880 17125
rect 18920 17155 18960 17160
rect 18920 17125 18925 17155
rect 18955 17125 18960 17155
rect 18920 17120 18960 17125
rect 19000 17155 19040 17160
rect 19000 17125 19005 17155
rect 19035 17125 19040 17155
rect 19000 17120 19040 17125
rect 19080 17155 19120 17160
rect 19080 17125 19085 17155
rect 19115 17125 19120 17155
rect 19080 17120 19120 17125
rect 19160 17155 19200 17160
rect 19160 17125 19165 17155
rect 19195 17125 19200 17155
rect 19160 17120 19200 17125
rect 19240 17155 19280 17160
rect 19240 17125 19245 17155
rect 19275 17125 19280 17155
rect 19240 17120 19280 17125
rect 19320 17155 19360 17160
rect 19320 17125 19325 17155
rect 19355 17125 19360 17155
rect 19320 17120 19360 17125
rect 19400 17155 19440 17160
rect 19400 17125 19405 17155
rect 19435 17125 19440 17155
rect 19400 17120 19440 17125
rect 19480 17155 19520 17160
rect 19480 17125 19485 17155
rect 19515 17125 19520 17155
rect 19480 17120 19520 17125
rect 19560 17155 19600 17160
rect 19560 17125 19565 17155
rect 19595 17125 19600 17155
rect 19560 17120 19600 17125
rect 19640 17155 19680 17160
rect 19640 17125 19645 17155
rect 19675 17125 19680 17155
rect 19640 17120 19680 17125
rect 19720 17155 19760 17160
rect 19720 17125 19725 17155
rect 19755 17125 19760 17155
rect 19720 17120 19760 17125
rect 19800 17155 19840 17160
rect 19800 17125 19805 17155
rect 19835 17125 19840 17155
rect 19800 17120 19840 17125
rect 19880 17155 19920 17160
rect 19880 17125 19885 17155
rect 19915 17125 19920 17155
rect 19880 17120 19920 17125
rect 19960 17155 20000 17160
rect 19960 17125 19965 17155
rect 19995 17125 20000 17155
rect 19960 17120 20000 17125
rect 20040 17155 20080 17160
rect 20040 17125 20045 17155
rect 20075 17125 20080 17155
rect 20040 17120 20080 17125
rect 20120 17155 20160 17160
rect 20120 17125 20125 17155
rect 20155 17125 20160 17155
rect 20120 17120 20160 17125
rect 20200 17155 20240 17160
rect 20200 17125 20205 17155
rect 20235 17125 20240 17155
rect 20200 17120 20240 17125
rect 20280 17155 20320 17160
rect 20280 17125 20285 17155
rect 20315 17125 20320 17155
rect 20280 17120 20320 17125
rect 20360 17155 20400 17160
rect 20360 17125 20365 17155
rect 20395 17125 20400 17155
rect 20360 17120 20400 17125
rect 20440 17155 20480 17160
rect 20440 17125 20445 17155
rect 20475 17125 20480 17155
rect 20440 17120 20480 17125
rect 20520 17155 20560 17160
rect 20520 17125 20525 17155
rect 20555 17125 20560 17155
rect 20520 17120 20560 17125
rect 20600 17155 20640 17160
rect 20600 17125 20605 17155
rect 20635 17125 20640 17155
rect 20600 17120 20640 17125
rect 20680 17155 20720 17160
rect 20680 17125 20685 17155
rect 20715 17125 20720 17155
rect 20680 17120 20720 17125
rect 20760 17155 20800 17160
rect 20760 17125 20765 17155
rect 20795 17125 20800 17155
rect 20760 17120 20800 17125
rect 20840 17155 20880 17160
rect 20840 17125 20845 17155
rect 20875 17125 20880 17155
rect 20840 17120 20880 17125
rect 20920 17155 20960 17160
rect 20920 17125 20925 17155
rect 20955 17125 20960 17155
rect 20920 17120 20960 17125
rect 0 16995 40 17000
rect 0 16965 5 16995
rect 35 16965 40 16995
rect 0 16960 40 16965
rect 80 16995 120 17000
rect 80 16965 85 16995
rect 115 16965 120 16995
rect 80 16960 120 16965
rect 160 16995 200 17000
rect 160 16965 165 16995
rect 195 16965 200 16995
rect 160 16960 200 16965
rect 240 16995 280 17000
rect 240 16965 245 16995
rect 275 16965 280 16995
rect 240 16960 280 16965
rect 320 16995 360 17000
rect 320 16965 325 16995
rect 355 16965 360 16995
rect 320 16960 360 16965
rect 400 16995 440 17000
rect 400 16965 405 16995
rect 435 16965 440 16995
rect 400 16960 440 16965
rect 480 16995 520 17000
rect 480 16965 485 16995
rect 515 16965 520 16995
rect 480 16960 520 16965
rect 560 16995 600 17000
rect 560 16965 565 16995
rect 595 16965 600 16995
rect 560 16960 600 16965
rect 640 16995 680 17000
rect 640 16965 645 16995
rect 675 16965 680 16995
rect 640 16960 680 16965
rect 720 16995 760 17000
rect 720 16965 725 16995
rect 755 16965 760 16995
rect 720 16960 760 16965
rect 800 16995 840 17000
rect 800 16965 805 16995
rect 835 16965 840 16995
rect 800 16960 840 16965
rect 880 16995 920 17000
rect 880 16965 885 16995
rect 915 16965 920 16995
rect 880 16960 920 16965
rect 960 16995 1000 17000
rect 960 16965 965 16995
rect 995 16965 1000 16995
rect 960 16960 1000 16965
rect 1040 16995 1080 17000
rect 1040 16965 1045 16995
rect 1075 16965 1080 16995
rect 1040 16960 1080 16965
rect 1120 16995 1160 17000
rect 1120 16965 1125 16995
rect 1155 16965 1160 16995
rect 1120 16960 1160 16965
rect 1200 16995 1240 17000
rect 1200 16965 1205 16995
rect 1235 16965 1240 16995
rect 1200 16960 1240 16965
rect 1280 16995 1320 17000
rect 1280 16965 1285 16995
rect 1315 16965 1320 16995
rect 1280 16960 1320 16965
rect 1360 16995 1400 17000
rect 1360 16965 1365 16995
rect 1395 16965 1400 16995
rect 1360 16960 1400 16965
rect 1440 16995 1480 17000
rect 1440 16965 1445 16995
rect 1475 16965 1480 16995
rect 1440 16960 1480 16965
rect 1520 16995 1560 17000
rect 1520 16965 1525 16995
rect 1555 16965 1560 16995
rect 1520 16960 1560 16965
rect 1600 16995 1640 17000
rect 1600 16965 1605 16995
rect 1635 16965 1640 16995
rect 1600 16960 1640 16965
rect 1680 16995 1720 17000
rect 1680 16965 1685 16995
rect 1715 16965 1720 16995
rect 1680 16960 1720 16965
rect 1760 16995 1800 17000
rect 1760 16965 1765 16995
rect 1795 16965 1800 16995
rect 1760 16960 1800 16965
rect 1840 16995 1880 17000
rect 1840 16965 1845 16995
rect 1875 16965 1880 16995
rect 1840 16960 1880 16965
rect 1920 16995 1960 17000
rect 1920 16965 1925 16995
rect 1955 16965 1960 16995
rect 1920 16960 1960 16965
rect 2000 16995 2040 17000
rect 2000 16965 2005 16995
rect 2035 16965 2040 16995
rect 2000 16960 2040 16965
rect 2080 16995 2120 17000
rect 2080 16965 2085 16995
rect 2115 16965 2120 16995
rect 2080 16960 2120 16965
rect 2160 16995 2200 17000
rect 2160 16965 2165 16995
rect 2195 16965 2200 16995
rect 2160 16960 2200 16965
rect 2240 16995 2280 17000
rect 2240 16965 2245 16995
rect 2275 16965 2280 16995
rect 2240 16960 2280 16965
rect 2320 16995 2360 17000
rect 2320 16965 2325 16995
rect 2355 16965 2360 16995
rect 2320 16960 2360 16965
rect 2400 16995 2440 17000
rect 2400 16965 2405 16995
rect 2435 16965 2440 16995
rect 2400 16960 2440 16965
rect 2480 16995 2520 17000
rect 2480 16965 2485 16995
rect 2515 16965 2520 16995
rect 2480 16960 2520 16965
rect 2560 16995 2600 17000
rect 2560 16965 2565 16995
rect 2595 16965 2600 16995
rect 2560 16960 2600 16965
rect 2640 16995 2680 17000
rect 2640 16965 2645 16995
rect 2675 16965 2680 16995
rect 2640 16960 2680 16965
rect 2720 16995 2760 17000
rect 2720 16965 2725 16995
rect 2755 16965 2760 16995
rect 2720 16960 2760 16965
rect 2800 16995 2840 17000
rect 2800 16965 2805 16995
rect 2835 16965 2840 16995
rect 2800 16960 2840 16965
rect 2880 16995 2920 17000
rect 2880 16965 2885 16995
rect 2915 16965 2920 16995
rect 2880 16960 2920 16965
rect 2960 16995 3000 17000
rect 2960 16965 2965 16995
rect 2995 16965 3000 16995
rect 2960 16960 3000 16965
rect 3040 16995 3080 17000
rect 3040 16965 3045 16995
rect 3075 16965 3080 16995
rect 3040 16960 3080 16965
rect 3120 16995 3160 17000
rect 3120 16965 3125 16995
rect 3155 16965 3160 16995
rect 3120 16960 3160 16965
rect 3200 16995 3240 17000
rect 3200 16965 3205 16995
rect 3235 16965 3240 16995
rect 3200 16960 3240 16965
rect 3280 16995 3320 17000
rect 3280 16965 3285 16995
rect 3315 16965 3320 16995
rect 3280 16960 3320 16965
rect 3360 16995 3400 17000
rect 3360 16965 3365 16995
rect 3395 16965 3400 16995
rect 3360 16960 3400 16965
rect 3440 16995 3480 17000
rect 3440 16965 3445 16995
rect 3475 16965 3480 16995
rect 3440 16960 3480 16965
rect 3520 16995 3560 17000
rect 3520 16965 3525 16995
rect 3555 16965 3560 16995
rect 3520 16960 3560 16965
rect 3600 16995 3640 17000
rect 3600 16965 3605 16995
rect 3635 16965 3640 16995
rect 3600 16960 3640 16965
rect 3680 16995 3720 17000
rect 3680 16965 3685 16995
rect 3715 16965 3720 16995
rect 3680 16960 3720 16965
rect 3760 16995 3800 17000
rect 3760 16965 3765 16995
rect 3795 16965 3800 16995
rect 3760 16960 3800 16965
rect 3840 16995 3880 17000
rect 3840 16965 3845 16995
rect 3875 16965 3880 16995
rect 3840 16960 3880 16965
rect 3920 16995 3960 17000
rect 3920 16965 3925 16995
rect 3955 16965 3960 16995
rect 3920 16960 3960 16965
rect 4000 16995 4040 17000
rect 4000 16965 4005 16995
rect 4035 16965 4040 16995
rect 4000 16960 4040 16965
rect 4080 16995 4120 17000
rect 4080 16965 4085 16995
rect 4115 16965 4120 16995
rect 4080 16960 4120 16965
rect 4160 16995 4200 17000
rect 4160 16965 4165 16995
rect 4195 16965 4200 16995
rect 4160 16960 4200 16965
rect 6240 16995 6280 17000
rect 6240 16965 6245 16995
rect 6275 16965 6280 16995
rect 6240 16960 6280 16965
rect 6320 16995 6360 17000
rect 6320 16965 6325 16995
rect 6355 16965 6360 16995
rect 6320 16960 6360 16965
rect 6400 16995 6440 17000
rect 6400 16965 6405 16995
rect 6435 16965 6440 16995
rect 6400 16960 6440 16965
rect 6480 16995 6520 17000
rect 6480 16965 6485 16995
rect 6515 16965 6520 16995
rect 6480 16960 6520 16965
rect 6560 16995 6600 17000
rect 6560 16965 6565 16995
rect 6595 16965 6600 16995
rect 6560 16960 6600 16965
rect 6640 16995 6680 17000
rect 6640 16965 6645 16995
rect 6675 16965 6680 16995
rect 6640 16960 6680 16965
rect 6720 16995 6760 17000
rect 6720 16965 6725 16995
rect 6755 16965 6760 16995
rect 6720 16960 6760 16965
rect 6800 16995 6840 17000
rect 6800 16965 6805 16995
rect 6835 16965 6840 16995
rect 6800 16960 6840 16965
rect 6880 16995 6920 17000
rect 6880 16965 6885 16995
rect 6915 16965 6920 16995
rect 6880 16960 6920 16965
rect 6960 16995 7000 17000
rect 6960 16965 6965 16995
rect 6995 16965 7000 16995
rect 6960 16960 7000 16965
rect 7040 16995 7080 17000
rect 7040 16965 7045 16995
rect 7075 16965 7080 16995
rect 7040 16960 7080 16965
rect 7120 16995 7160 17000
rect 7120 16965 7125 16995
rect 7155 16965 7160 16995
rect 7120 16960 7160 16965
rect 7200 16995 7240 17000
rect 7200 16965 7205 16995
rect 7235 16965 7240 16995
rect 7200 16960 7240 16965
rect 7280 16995 7320 17000
rect 7280 16965 7285 16995
rect 7315 16965 7320 16995
rect 7280 16960 7320 16965
rect 7360 16995 7400 17000
rect 7360 16965 7365 16995
rect 7395 16965 7400 16995
rect 7360 16960 7400 16965
rect 7440 16995 7480 17000
rect 7440 16965 7445 16995
rect 7475 16965 7480 16995
rect 7440 16960 7480 16965
rect 7520 16995 7560 17000
rect 7520 16965 7525 16995
rect 7555 16965 7560 16995
rect 7520 16960 7560 16965
rect 7600 16995 7640 17000
rect 7600 16965 7605 16995
rect 7635 16965 7640 16995
rect 7600 16960 7640 16965
rect 7680 16995 7720 17000
rect 7680 16965 7685 16995
rect 7715 16965 7720 16995
rect 7680 16960 7720 16965
rect 7760 16995 7800 17000
rect 7760 16965 7765 16995
rect 7795 16965 7800 16995
rect 7760 16960 7800 16965
rect 7840 16995 7880 17000
rect 7840 16965 7845 16995
rect 7875 16965 7880 16995
rect 7840 16960 7880 16965
rect 7920 16995 7960 17000
rect 7920 16965 7925 16995
rect 7955 16965 7960 16995
rect 7920 16960 7960 16965
rect 8000 16995 8040 17000
rect 8000 16965 8005 16995
rect 8035 16965 8040 16995
rect 8000 16960 8040 16965
rect 8080 16995 8120 17000
rect 8080 16965 8085 16995
rect 8115 16965 8120 16995
rect 8080 16960 8120 16965
rect 8160 16995 8200 17000
rect 8160 16965 8165 16995
rect 8195 16965 8200 16995
rect 8160 16960 8200 16965
rect 8240 16995 8280 17000
rect 8240 16965 8245 16995
rect 8275 16965 8280 16995
rect 8240 16960 8280 16965
rect 8320 16995 8360 17000
rect 8320 16965 8325 16995
rect 8355 16965 8360 16995
rect 8320 16960 8360 16965
rect 8400 16995 8440 17000
rect 8400 16965 8405 16995
rect 8435 16965 8440 16995
rect 8400 16960 8440 16965
rect 8480 16995 8520 17000
rect 8480 16965 8485 16995
rect 8515 16965 8520 16995
rect 8480 16960 8520 16965
rect 8560 16995 8600 17000
rect 8560 16965 8565 16995
rect 8595 16965 8600 16995
rect 8560 16960 8600 16965
rect 8640 16995 8680 17000
rect 8640 16965 8645 16995
rect 8675 16965 8680 16995
rect 8640 16960 8680 16965
rect 8720 16995 8760 17000
rect 8720 16965 8725 16995
rect 8755 16965 8760 16995
rect 8720 16960 8760 16965
rect 8800 16995 8840 17000
rect 8800 16965 8805 16995
rect 8835 16965 8840 16995
rect 8800 16960 8840 16965
rect 8880 16995 8920 17000
rect 8880 16965 8885 16995
rect 8915 16965 8920 16995
rect 8880 16960 8920 16965
rect 8960 16995 9000 17000
rect 8960 16965 8965 16995
rect 8995 16965 9000 16995
rect 8960 16960 9000 16965
rect 9040 16995 9080 17000
rect 9040 16965 9045 16995
rect 9075 16965 9080 16995
rect 9040 16960 9080 16965
rect 9120 16995 9160 17000
rect 9120 16965 9125 16995
rect 9155 16965 9160 16995
rect 9120 16960 9160 16965
rect 9200 16995 9240 17000
rect 9200 16965 9205 16995
rect 9235 16965 9240 16995
rect 9200 16960 9240 16965
rect 9280 16995 9320 17000
rect 9280 16965 9285 16995
rect 9315 16965 9320 16995
rect 9280 16960 9320 16965
rect 9360 16995 9400 17000
rect 9360 16965 9365 16995
rect 9395 16965 9400 16995
rect 9360 16960 9400 16965
rect 9440 16995 9480 17000
rect 9440 16965 9445 16995
rect 9475 16965 9480 16995
rect 9440 16960 9480 16965
rect 11560 16995 11600 17000
rect 11560 16965 11565 16995
rect 11595 16965 11600 16995
rect 11560 16960 11600 16965
rect 11640 16995 11680 17000
rect 11640 16965 11645 16995
rect 11675 16965 11680 16995
rect 11640 16960 11680 16965
rect 11720 16995 11760 17000
rect 11720 16965 11725 16995
rect 11755 16965 11760 16995
rect 11720 16960 11760 16965
rect 11800 16995 11840 17000
rect 11800 16965 11805 16995
rect 11835 16965 11840 16995
rect 11800 16960 11840 16965
rect 11880 16995 11920 17000
rect 11880 16965 11885 16995
rect 11915 16965 11920 16995
rect 11880 16960 11920 16965
rect 11960 16995 12000 17000
rect 11960 16965 11965 16995
rect 11995 16965 12000 16995
rect 11960 16960 12000 16965
rect 12040 16995 12080 17000
rect 12040 16965 12045 16995
rect 12075 16965 12080 16995
rect 12040 16960 12080 16965
rect 12120 16995 12160 17000
rect 12120 16965 12125 16995
rect 12155 16965 12160 16995
rect 12120 16960 12160 16965
rect 12200 16995 12240 17000
rect 12200 16965 12205 16995
rect 12235 16965 12240 16995
rect 12200 16960 12240 16965
rect 12280 16995 12320 17000
rect 12280 16965 12285 16995
rect 12315 16965 12320 16995
rect 12280 16960 12320 16965
rect 12360 16995 12400 17000
rect 12360 16965 12365 16995
rect 12395 16965 12400 16995
rect 12360 16960 12400 16965
rect 12440 16995 12480 17000
rect 12440 16965 12445 16995
rect 12475 16965 12480 16995
rect 12440 16960 12480 16965
rect 12520 16995 12560 17000
rect 12520 16965 12525 16995
rect 12555 16965 12560 16995
rect 12520 16960 12560 16965
rect 12600 16995 12640 17000
rect 12600 16965 12605 16995
rect 12635 16965 12640 16995
rect 12600 16960 12640 16965
rect 12680 16995 12720 17000
rect 12680 16965 12685 16995
rect 12715 16965 12720 16995
rect 12680 16960 12720 16965
rect 12760 16995 12800 17000
rect 12760 16965 12765 16995
rect 12795 16965 12800 16995
rect 12760 16960 12800 16965
rect 12840 16995 12880 17000
rect 12840 16965 12845 16995
rect 12875 16965 12880 16995
rect 12840 16960 12880 16965
rect 12920 16995 12960 17000
rect 12920 16965 12925 16995
rect 12955 16965 12960 16995
rect 12920 16960 12960 16965
rect 13000 16995 13040 17000
rect 13000 16965 13005 16995
rect 13035 16965 13040 16995
rect 13000 16960 13040 16965
rect 13080 16995 13120 17000
rect 13080 16965 13085 16995
rect 13115 16965 13120 16995
rect 13080 16960 13120 16965
rect 13160 16995 13200 17000
rect 13160 16965 13165 16995
rect 13195 16965 13200 16995
rect 13160 16960 13200 16965
rect 13240 16995 13280 17000
rect 13240 16965 13245 16995
rect 13275 16965 13280 16995
rect 13240 16960 13280 16965
rect 13320 16995 13360 17000
rect 13320 16965 13325 16995
rect 13355 16965 13360 16995
rect 13320 16960 13360 16965
rect 13400 16995 13440 17000
rect 13400 16965 13405 16995
rect 13435 16965 13440 16995
rect 13400 16960 13440 16965
rect 13480 16995 13520 17000
rect 13480 16965 13485 16995
rect 13515 16965 13520 16995
rect 13480 16960 13520 16965
rect 13560 16995 13600 17000
rect 13560 16965 13565 16995
rect 13595 16965 13600 16995
rect 13560 16960 13600 16965
rect 13640 16995 13680 17000
rect 13640 16965 13645 16995
rect 13675 16965 13680 16995
rect 13640 16960 13680 16965
rect 13720 16995 13760 17000
rect 13720 16965 13725 16995
rect 13755 16965 13760 16995
rect 13720 16960 13760 16965
rect 13800 16995 13840 17000
rect 13800 16965 13805 16995
rect 13835 16965 13840 16995
rect 13800 16960 13840 16965
rect 13880 16995 13920 17000
rect 13880 16965 13885 16995
rect 13915 16965 13920 16995
rect 13880 16960 13920 16965
rect 13960 16995 14000 17000
rect 13960 16965 13965 16995
rect 13995 16965 14000 16995
rect 13960 16960 14000 16965
rect 14040 16995 14080 17000
rect 14040 16965 14045 16995
rect 14075 16965 14080 16995
rect 14040 16960 14080 16965
rect 14120 16995 14160 17000
rect 14120 16965 14125 16995
rect 14155 16965 14160 16995
rect 14120 16960 14160 16965
rect 14200 16995 14240 17000
rect 14200 16965 14205 16995
rect 14235 16965 14240 16995
rect 14200 16960 14240 16965
rect 14280 16995 14320 17000
rect 14280 16965 14285 16995
rect 14315 16965 14320 16995
rect 14280 16960 14320 16965
rect 14360 16995 14400 17000
rect 14360 16965 14365 16995
rect 14395 16965 14400 16995
rect 14360 16960 14400 16965
rect 14440 16995 14480 17000
rect 14440 16965 14445 16995
rect 14475 16965 14480 16995
rect 14440 16960 14480 16965
rect 14520 16995 14560 17000
rect 14520 16965 14525 16995
rect 14555 16965 14560 16995
rect 14520 16960 14560 16965
rect 14600 16995 14640 17000
rect 14600 16965 14605 16995
rect 14635 16965 14640 16995
rect 14600 16960 14640 16965
rect 14680 16995 14720 17000
rect 14680 16965 14685 16995
rect 14715 16965 14720 16995
rect 14680 16960 14720 16965
rect 16760 16995 16800 17000
rect 16760 16965 16765 16995
rect 16795 16965 16800 16995
rect 16760 16960 16800 16965
rect 16840 16995 16880 17000
rect 16840 16965 16845 16995
rect 16875 16965 16880 16995
rect 16840 16960 16880 16965
rect 16920 16995 16960 17000
rect 16920 16965 16925 16995
rect 16955 16965 16960 16995
rect 16920 16960 16960 16965
rect 17000 16995 17040 17000
rect 17000 16965 17005 16995
rect 17035 16965 17040 16995
rect 17000 16960 17040 16965
rect 17080 16995 17120 17000
rect 17080 16965 17085 16995
rect 17115 16965 17120 16995
rect 17080 16960 17120 16965
rect 17160 16995 17200 17000
rect 17160 16965 17165 16995
rect 17195 16965 17200 16995
rect 17160 16960 17200 16965
rect 17240 16995 17280 17000
rect 17240 16965 17245 16995
rect 17275 16965 17280 16995
rect 17240 16960 17280 16965
rect 17320 16995 17360 17000
rect 17320 16965 17325 16995
rect 17355 16965 17360 16995
rect 17320 16960 17360 16965
rect 17400 16995 17440 17000
rect 17400 16965 17405 16995
rect 17435 16965 17440 16995
rect 17400 16960 17440 16965
rect 17480 16995 17520 17000
rect 17480 16965 17485 16995
rect 17515 16965 17520 16995
rect 17480 16960 17520 16965
rect 17560 16995 17600 17000
rect 17560 16965 17565 16995
rect 17595 16965 17600 16995
rect 17560 16960 17600 16965
rect 17640 16995 17680 17000
rect 17640 16965 17645 16995
rect 17675 16965 17680 16995
rect 17640 16960 17680 16965
rect 17720 16995 17760 17000
rect 17720 16965 17725 16995
rect 17755 16965 17760 16995
rect 17720 16960 17760 16965
rect 17800 16995 17840 17000
rect 17800 16965 17805 16995
rect 17835 16965 17840 16995
rect 17800 16960 17840 16965
rect 17880 16995 17920 17000
rect 17880 16965 17885 16995
rect 17915 16965 17920 16995
rect 17880 16960 17920 16965
rect 17960 16995 18000 17000
rect 17960 16965 17965 16995
rect 17995 16965 18000 16995
rect 17960 16960 18000 16965
rect 18040 16995 18080 17000
rect 18040 16965 18045 16995
rect 18075 16965 18080 16995
rect 18040 16960 18080 16965
rect 18120 16995 18160 17000
rect 18120 16965 18125 16995
rect 18155 16965 18160 16995
rect 18120 16960 18160 16965
rect 18200 16995 18240 17000
rect 18200 16965 18205 16995
rect 18235 16965 18240 16995
rect 18200 16960 18240 16965
rect 18280 16995 18320 17000
rect 18280 16965 18285 16995
rect 18315 16965 18320 16995
rect 18280 16960 18320 16965
rect 18360 16995 18400 17000
rect 18360 16965 18365 16995
rect 18395 16965 18400 16995
rect 18360 16960 18400 16965
rect 18440 16995 18480 17000
rect 18440 16965 18445 16995
rect 18475 16965 18480 16995
rect 18440 16960 18480 16965
rect 18520 16995 18560 17000
rect 18520 16965 18525 16995
rect 18555 16965 18560 16995
rect 18520 16960 18560 16965
rect 18600 16995 18640 17000
rect 18600 16965 18605 16995
rect 18635 16965 18640 16995
rect 18600 16960 18640 16965
rect 18680 16995 18720 17000
rect 18680 16965 18685 16995
rect 18715 16965 18720 16995
rect 18680 16960 18720 16965
rect 18760 16995 18800 17000
rect 18760 16965 18765 16995
rect 18795 16965 18800 16995
rect 18760 16960 18800 16965
rect 18840 16995 18880 17000
rect 18840 16965 18845 16995
rect 18875 16965 18880 16995
rect 18840 16960 18880 16965
rect 18920 16995 18960 17000
rect 18920 16965 18925 16995
rect 18955 16965 18960 16995
rect 18920 16960 18960 16965
rect 19000 16995 19040 17000
rect 19000 16965 19005 16995
rect 19035 16965 19040 16995
rect 19000 16960 19040 16965
rect 19080 16995 19120 17000
rect 19080 16965 19085 16995
rect 19115 16965 19120 16995
rect 19080 16960 19120 16965
rect 19160 16995 19200 17000
rect 19160 16965 19165 16995
rect 19195 16965 19200 16995
rect 19160 16960 19200 16965
rect 19240 16995 19280 17000
rect 19240 16965 19245 16995
rect 19275 16965 19280 16995
rect 19240 16960 19280 16965
rect 19320 16995 19360 17000
rect 19320 16965 19325 16995
rect 19355 16965 19360 16995
rect 19320 16960 19360 16965
rect 19400 16995 19440 17000
rect 19400 16965 19405 16995
rect 19435 16965 19440 16995
rect 19400 16960 19440 16965
rect 19480 16995 19520 17000
rect 19480 16965 19485 16995
rect 19515 16965 19520 16995
rect 19480 16960 19520 16965
rect 19560 16995 19600 17000
rect 19560 16965 19565 16995
rect 19595 16965 19600 16995
rect 19560 16960 19600 16965
rect 19640 16995 19680 17000
rect 19640 16965 19645 16995
rect 19675 16965 19680 16995
rect 19640 16960 19680 16965
rect 19720 16995 19760 17000
rect 19720 16965 19725 16995
rect 19755 16965 19760 16995
rect 19720 16960 19760 16965
rect 19800 16995 19840 17000
rect 19800 16965 19805 16995
rect 19835 16965 19840 16995
rect 19800 16960 19840 16965
rect 19880 16995 19920 17000
rect 19880 16965 19885 16995
rect 19915 16965 19920 16995
rect 19880 16960 19920 16965
rect 19960 16995 20000 17000
rect 19960 16965 19965 16995
rect 19995 16965 20000 16995
rect 19960 16960 20000 16965
rect 20040 16995 20080 17000
rect 20040 16965 20045 16995
rect 20075 16965 20080 16995
rect 20040 16960 20080 16965
rect 20120 16995 20160 17000
rect 20120 16965 20125 16995
rect 20155 16965 20160 16995
rect 20120 16960 20160 16965
rect 20200 16995 20240 17000
rect 20200 16965 20205 16995
rect 20235 16965 20240 16995
rect 20200 16960 20240 16965
rect 20280 16995 20320 17000
rect 20280 16965 20285 16995
rect 20315 16965 20320 16995
rect 20280 16960 20320 16965
rect 20360 16995 20400 17000
rect 20360 16965 20365 16995
rect 20395 16965 20400 16995
rect 20360 16960 20400 16965
rect 20440 16995 20480 17000
rect 20440 16965 20445 16995
rect 20475 16965 20480 16995
rect 20440 16960 20480 16965
rect 20520 16995 20560 17000
rect 20520 16965 20525 16995
rect 20555 16965 20560 16995
rect 20520 16960 20560 16965
rect 20600 16995 20640 17000
rect 20600 16965 20605 16995
rect 20635 16965 20640 16995
rect 20600 16960 20640 16965
rect 20680 16995 20720 17000
rect 20680 16965 20685 16995
rect 20715 16965 20720 16995
rect 20680 16960 20720 16965
rect 20760 16995 20800 17000
rect 20760 16965 20765 16995
rect 20795 16965 20800 16995
rect 20760 16960 20800 16965
rect 20840 16995 20880 17000
rect 20840 16965 20845 16995
rect 20875 16965 20880 16995
rect 20840 16960 20880 16965
rect 20920 16995 20960 17000
rect 20920 16965 20925 16995
rect 20955 16965 20960 16995
rect 20920 16960 20960 16965
rect 0 16915 40 16920
rect 0 16885 5 16915
rect 35 16885 40 16915
rect 0 16880 40 16885
rect 80 16915 120 16920
rect 80 16885 85 16915
rect 115 16885 120 16915
rect 80 16880 120 16885
rect 160 16915 200 16920
rect 160 16885 165 16915
rect 195 16885 200 16915
rect 160 16880 200 16885
rect 240 16915 280 16920
rect 240 16885 245 16915
rect 275 16885 280 16915
rect 240 16880 280 16885
rect 320 16915 360 16920
rect 320 16885 325 16915
rect 355 16885 360 16915
rect 320 16880 360 16885
rect 400 16915 440 16920
rect 400 16885 405 16915
rect 435 16885 440 16915
rect 400 16880 440 16885
rect 480 16915 520 16920
rect 480 16885 485 16915
rect 515 16885 520 16915
rect 480 16880 520 16885
rect 560 16915 600 16920
rect 560 16885 565 16915
rect 595 16885 600 16915
rect 560 16880 600 16885
rect 640 16915 680 16920
rect 640 16885 645 16915
rect 675 16885 680 16915
rect 640 16880 680 16885
rect 720 16915 760 16920
rect 720 16885 725 16915
rect 755 16885 760 16915
rect 720 16880 760 16885
rect 800 16915 840 16920
rect 800 16885 805 16915
rect 835 16885 840 16915
rect 800 16880 840 16885
rect 880 16915 920 16920
rect 880 16885 885 16915
rect 915 16885 920 16915
rect 880 16880 920 16885
rect 960 16915 1000 16920
rect 960 16885 965 16915
rect 995 16885 1000 16915
rect 960 16880 1000 16885
rect 1040 16915 1080 16920
rect 1040 16885 1045 16915
rect 1075 16885 1080 16915
rect 1040 16880 1080 16885
rect 1120 16915 1160 16920
rect 1120 16885 1125 16915
rect 1155 16885 1160 16915
rect 1120 16880 1160 16885
rect 1200 16915 1240 16920
rect 1200 16885 1205 16915
rect 1235 16885 1240 16915
rect 1200 16880 1240 16885
rect 1280 16915 1320 16920
rect 1280 16885 1285 16915
rect 1315 16885 1320 16915
rect 1280 16880 1320 16885
rect 1360 16915 1400 16920
rect 1360 16885 1365 16915
rect 1395 16885 1400 16915
rect 1360 16880 1400 16885
rect 1440 16915 1480 16920
rect 1440 16885 1445 16915
rect 1475 16885 1480 16915
rect 1440 16880 1480 16885
rect 1520 16915 1560 16920
rect 1520 16885 1525 16915
rect 1555 16885 1560 16915
rect 1520 16880 1560 16885
rect 1600 16915 1640 16920
rect 1600 16885 1605 16915
rect 1635 16885 1640 16915
rect 1600 16880 1640 16885
rect 1680 16915 1720 16920
rect 1680 16885 1685 16915
rect 1715 16885 1720 16915
rect 1680 16880 1720 16885
rect 1760 16915 1800 16920
rect 1760 16885 1765 16915
rect 1795 16885 1800 16915
rect 1760 16880 1800 16885
rect 1840 16915 1880 16920
rect 1840 16885 1845 16915
rect 1875 16885 1880 16915
rect 1840 16880 1880 16885
rect 1920 16915 1960 16920
rect 1920 16885 1925 16915
rect 1955 16885 1960 16915
rect 1920 16880 1960 16885
rect 2000 16915 2040 16920
rect 2000 16885 2005 16915
rect 2035 16885 2040 16915
rect 2000 16880 2040 16885
rect 2080 16915 2120 16920
rect 2080 16885 2085 16915
rect 2115 16885 2120 16915
rect 2080 16880 2120 16885
rect 2160 16915 2200 16920
rect 2160 16885 2165 16915
rect 2195 16885 2200 16915
rect 2160 16880 2200 16885
rect 2240 16915 2280 16920
rect 2240 16885 2245 16915
rect 2275 16885 2280 16915
rect 2240 16880 2280 16885
rect 2320 16915 2360 16920
rect 2320 16885 2325 16915
rect 2355 16885 2360 16915
rect 2320 16880 2360 16885
rect 2400 16915 2440 16920
rect 2400 16885 2405 16915
rect 2435 16885 2440 16915
rect 2400 16880 2440 16885
rect 2480 16915 2520 16920
rect 2480 16885 2485 16915
rect 2515 16885 2520 16915
rect 2480 16880 2520 16885
rect 2560 16915 2600 16920
rect 2560 16885 2565 16915
rect 2595 16885 2600 16915
rect 2560 16880 2600 16885
rect 2640 16915 2680 16920
rect 2640 16885 2645 16915
rect 2675 16885 2680 16915
rect 2640 16880 2680 16885
rect 2720 16915 2760 16920
rect 2720 16885 2725 16915
rect 2755 16885 2760 16915
rect 2720 16880 2760 16885
rect 2800 16915 2840 16920
rect 2800 16885 2805 16915
rect 2835 16885 2840 16915
rect 2800 16880 2840 16885
rect 2880 16915 2920 16920
rect 2880 16885 2885 16915
rect 2915 16885 2920 16915
rect 2880 16880 2920 16885
rect 2960 16915 3000 16920
rect 2960 16885 2965 16915
rect 2995 16885 3000 16915
rect 2960 16880 3000 16885
rect 3040 16915 3080 16920
rect 3040 16885 3045 16915
rect 3075 16885 3080 16915
rect 3040 16880 3080 16885
rect 3120 16915 3160 16920
rect 3120 16885 3125 16915
rect 3155 16885 3160 16915
rect 3120 16880 3160 16885
rect 3200 16915 3240 16920
rect 3200 16885 3205 16915
rect 3235 16885 3240 16915
rect 3200 16880 3240 16885
rect 3280 16915 3320 16920
rect 3280 16885 3285 16915
rect 3315 16885 3320 16915
rect 3280 16880 3320 16885
rect 3360 16915 3400 16920
rect 3360 16885 3365 16915
rect 3395 16885 3400 16915
rect 3360 16880 3400 16885
rect 3440 16915 3480 16920
rect 3440 16885 3445 16915
rect 3475 16885 3480 16915
rect 3440 16880 3480 16885
rect 3520 16915 3560 16920
rect 3520 16885 3525 16915
rect 3555 16885 3560 16915
rect 3520 16880 3560 16885
rect 3600 16915 3640 16920
rect 3600 16885 3605 16915
rect 3635 16885 3640 16915
rect 3600 16880 3640 16885
rect 3680 16915 3720 16920
rect 3680 16885 3685 16915
rect 3715 16885 3720 16915
rect 3680 16880 3720 16885
rect 3760 16915 3800 16920
rect 3760 16885 3765 16915
rect 3795 16885 3800 16915
rect 3760 16880 3800 16885
rect 3840 16915 3880 16920
rect 3840 16885 3845 16915
rect 3875 16885 3880 16915
rect 3840 16880 3880 16885
rect 3920 16915 3960 16920
rect 3920 16885 3925 16915
rect 3955 16885 3960 16915
rect 3920 16880 3960 16885
rect 4000 16915 4040 16920
rect 4000 16885 4005 16915
rect 4035 16885 4040 16915
rect 4000 16880 4040 16885
rect 4080 16915 4120 16920
rect 4080 16885 4085 16915
rect 4115 16885 4120 16915
rect 4080 16880 4120 16885
rect 4160 16915 4200 16920
rect 4160 16885 4165 16915
rect 4195 16885 4200 16915
rect 4160 16880 4200 16885
rect 6240 16915 6280 16920
rect 6240 16885 6245 16915
rect 6275 16885 6280 16915
rect 6240 16880 6280 16885
rect 6320 16915 6360 16920
rect 6320 16885 6325 16915
rect 6355 16885 6360 16915
rect 6320 16880 6360 16885
rect 6400 16915 6440 16920
rect 6400 16885 6405 16915
rect 6435 16885 6440 16915
rect 6400 16880 6440 16885
rect 6480 16915 6520 16920
rect 6480 16885 6485 16915
rect 6515 16885 6520 16915
rect 6480 16880 6520 16885
rect 6560 16915 6600 16920
rect 6560 16885 6565 16915
rect 6595 16885 6600 16915
rect 6560 16880 6600 16885
rect 6640 16915 6680 16920
rect 6640 16885 6645 16915
rect 6675 16885 6680 16915
rect 6640 16880 6680 16885
rect 6720 16915 6760 16920
rect 6720 16885 6725 16915
rect 6755 16885 6760 16915
rect 6720 16880 6760 16885
rect 6800 16915 6840 16920
rect 6800 16885 6805 16915
rect 6835 16885 6840 16915
rect 6800 16880 6840 16885
rect 6880 16915 6920 16920
rect 6880 16885 6885 16915
rect 6915 16885 6920 16915
rect 6880 16880 6920 16885
rect 6960 16915 7000 16920
rect 6960 16885 6965 16915
rect 6995 16885 7000 16915
rect 6960 16880 7000 16885
rect 7040 16915 7080 16920
rect 7040 16885 7045 16915
rect 7075 16885 7080 16915
rect 7040 16880 7080 16885
rect 7120 16915 7160 16920
rect 7120 16885 7125 16915
rect 7155 16885 7160 16915
rect 7120 16880 7160 16885
rect 7200 16915 7240 16920
rect 7200 16885 7205 16915
rect 7235 16885 7240 16915
rect 7200 16880 7240 16885
rect 7280 16915 7320 16920
rect 7280 16885 7285 16915
rect 7315 16885 7320 16915
rect 7280 16880 7320 16885
rect 7360 16915 7400 16920
rect 7360 16885 7365 16915
rect 7395 16885 7400 16915
rect 7360 16880 7400 16885
rect 7440 16915 7480 16920
rect 7440 16885 7445 16915
rect 7475 16885 7480 16915
rect 7440 16880 7480 16885
rect 7520 16915 7560 16920
rect 7520 16885 7525 16915
rect 7555 16885 7560 16915
rect 7520 16880 7560 16885
rect 7600 16915 7640 16920
rect 7600 16885 7605 16915
rect 7635 16885 7640 16915
rect 7600 16880 7640 16885
rect 7680 16915 7720 16920
rect 7680 16885 7685 16915
rect 7715 16885 7720 16915
rect 7680 16880 7720 16885
rect 7760 16915 7800 16920
rect 7760 16885 7765 16915
rect 7795 16885 7800 16915
rect 7760 16880 7800 16885
rect 7840 16915 7880 16920
rect 7840 16885 7845 16915
rect 7875 16885 7880 16915
rect 7840 16880 7880 16885
rect 7920 16915 7960 16920
rect 7920 16885 7925 16915
rect 7955 16885 7960 16915
rect 7920 16880 7960 16885
rect 8000 16915 8040 16920
rect 8000 16885 8005 16915
rect 8035 16885 8040 16915
rect 8000 16880 8040 16885
rect 8080 16915 8120 16920
rect 8080 16885 8085 16915
rect 8115 16885 8120 16915
rect 8080 16880 8120 16885
rect 8160 16915 8200 16920
rect 8160 16885 8165 16915
rect 8195 16885 8200 16915
rect 8160 16880 8200 16885
rect 8240 16915 8280 16920
rect 8240 16885 8245 16915
rect 8275 16885 8280 16915
rect 8240 16880 8280 16885
rect 8320 16915 8360 16920
rect 8320 16885 8325 16915
rect 8355 16885 8360 16915
rect 8320 16880 8360 16885
rect 8400 16915 8440 16920
rect 8400 16885 8405 16915
rect 8435 16885 8440 16915
rect 8400 16880 8440 16885
rect 8480 16915 8520 16920
rect 8480 16885 8485 16915
rect 8515 16885 8520 16915
rect 8480 16880 8520 16885
rect 8560 16915 8600 16920
rect 8560 16885 8565 16915
rect 8595 16885 8600 16915
rect 8560 16880 8600 16885
rect 8640 16915 8680 16920
rect 8640 16885 8645 16915
rect 8675 16885 8680 16915
rect 8640 16880 8680 16885
rect 8720 16915 8760 16920
rect 8720 16885 8725 16915
rect 8755 16885 8760 16915
rect 8720 16880 8760 16885
rect 8800 16915 8840 16920
rect 8800 16885 8805 16915
rect 8835 16885 8840 16915
rect 8800 16880 8840 16885
rect 8880 16915 8920 16920
rect 8880 16885 8885 16915
rect 8915 16885 8920 16915
rect 8880 16880 8920 16885
rect 8960 16915 9000 16920
rect 8960 16885 8965 16915
rect 8995 16885 9000 16915
rect 8960 16880 9000 16885
rect 9040 16915 9080 16920
rect 9040 16885 9045 16915
rect 9075 16885 9080 16915
rect 9040 16880 9080 16885
rect 9120 16915 9160 16920
rect 9120 16885 9125 16915
rect 9155 16885 9160 16915
rect 9120 16880 9160 16885
rect 9200 16915 9240 16920
rect 9200 16885 9205 16915
rect 9235 16885 9240 16915
rect 9200 16880 9240 16885
rect 9280 16915 9320 16920
rect 9280 16885 9285 16915
rect 9315 16885 9320 16915
rect 9280 16880 9320 16885
rect 9360 16915 9400 16920
rect 9360 16885 9365 16915
rect 9395 16885 9400 16915
rect 9360 16880 9400 16885
rect 9440 16915 9480 16920
rect 9440 16885 9445 16915
rect 9475 16885 9480 16915
rect 9440 16880 9480 16885
rect 11560 16915 11600 16920
rect 11560 16885 11565 16915
rect 11595 16885 11600 16915
rect 11560 16880 11600 16885
rect 11640 16915 11680 16920
rect 11640 16885 11645 16915
rect 11675 16885 11680 16915
rect 11640 16880 11680 16885
rect 11720 16915 11760 16920
rect 11720 16885 11725 16915
rect 11755 16885 11760 16915
rect 11720 16880 11760 16885
rect 11800 16915 11840 16920
rect 11800 16885 11805 16915
rect 11835 16885 11840 16915
rect 11800 16880 11840 16885
rect 11880 16915 11920 16920
rect 11880 16885 11885 16915
rect 11915 16885 11920 16915
rect 11880 16880 11920 16885
rect 11960 16915 12000 16920
rect 11960 16885 11965 16915
rect 11995 16885 12000 16915
rect 11960 16880 12000 16885
rect 12040 16915 12080 16920
rect 12040 16885 12045 16915
rect 12075 16885 12080 16915
rect 12040 16880 12080 16885
rect 12120 16915 12160 16920
rect 12120 16885 12125 16915
rect 12155 16885 12160 16915
rect 12120 16880 12160 16885
rect 12200 16915 12240 16920
rect 12200 16885 12205 16915
rect 12235 16885 12240 16915
rect 12200 16880 12240 16885
rect 12280 16915 12320 16920
rect 12280 16885 12285 16915
rect 12315 16885 12320 16915
rect 12280 16880 12320 16885
rect 12360 16915 12400 16920
rect 12360 16885 12365 16915
rect 12395 16885 12400 16915
rect 12360 16880 12400 16885
rect 12440 16915 12480 16920
rect 12440 16885 12445 16915
rect 12475 16885 12480 16915
rect 12440 16880 12480 16885
rect 12520 16915 12560 16920
rect 12520 16885 12525 16915
rect 12555 16885 12560 16915
rect 12520 16880 12560 16885
rect 12600 16915 12640 16920
rect 12600 16885 12605 16915
rect 12635 16885 12640 16915
rect 12600 16880 12640 16885
rect 12680 16915 12720 16920
rect 12680 16885 12685 16915
rect 12715 16885 12720 16915
rect 12680 16880 12720 16885
rect 12760 16915 12800 16920
rect 12760 16885 12765 16915
rect 12795 16885 12800 16915
rect 12760 16880 12800 16885
rect 12840 16915 12880 16920
rect 12840 16885 12845 16915
rect 12875 16885 12880 16915
rect 12840 16880 12880 16885
rect 12920 16915 12960 16920
rect 12920 16885 12925 16915
rect 12955 16885 12960 16915
rect 12920 16880 12960 16885
rect 13000 16915 13040 16920
rect 13000 16885 13005 16915
rect 13035 16885 13040 16915
rect 13000 16880 13040 16885
rect 13080 16915 13120 16920
rect 13080 16885 13085 16915
rect 13115 16885 13120 16915
rect 13080 16880 13120 16885
rect 13160 16915 13200 16920
rect 13160 16885 13165 16915
rect 13195 16885 13200 16915
rect 13160 16880 13200 16885
rect 13240 16915 13280 16920
rect 13240 16885 13245 16915
rect 13275 16885 13280 16915
rect 13240 16880 13280 16885
rect 13320 16915 13360 16920
rect 13320 16885 13325 16915
rect 13355 16885 13360 16915
rect 13320 16880 13360 16885
rect 13400 16915 13440 16920
rect 13400 16885 13405 16915
rect 13435 16885 13440 16915
rect 13400 16880 13440 16885
rect 13480 16915 13520 16920
rect 13480 16885 13485 16915
rect 13515 16885 13520 16915
rect 13480 16880 13520 16885
rect 13560 16915 13600 16920
rect 13560 16885 13565 16915
rect 13595 16885 13600 16915
rect 13560 16880 13600 16885
rect 13640 16915 13680 16920
rect 13640 16885 13645 16915
rect 13675 16885 13680 16915
rect 13640 16880 13680 16885
rect 13720 16915 13760 16920
rect 13720 16885 13725 16915
rect 13755 16885 13760 16915
rect 13720 16880 13760 16885
rect 13800 16915 13840 16920
rect 13800 16885 13805 16915
rect 13835 16885 13840 16915
rect 13800 16880 13840 16885
rect 13880 16915 13920 16920
rect 13880 16885 13885 16915
rect 13915 16885 13920 16915
rect 13880 16880 13920 16885
rect 13960 16915 14000 16920
rect 13960 16885 13965 16915
rect 13995 16885 14000 16915
rect 13960 16880 14000 16885
rect 14040 16915 14080 16920
rect 14040 16885 14045 16915
rect 14075 16885 14080 16915
rect 14040 16880 14080 16885
rect 14120 16915 14160 16920
rect 14120 16885 14125 16915
rect 14155 16885 14160 16915
rect 14120 16880 14160 16885
rect 14200 16915 14240 16920
rect 14200 16885 14205 16915
rect 14235 16885 14240 16915
rect 14200 16880 14240 16885
rect 14280 16915 14320 16920
rect 14280 16885 14285 16915
rect 14315 16885 14320 16915
rect 14280 16880 14320 16885
rect 14360 16915 14400 16920
rect 14360 16885 14365 16915
rect 14395 16885 14400 16915
rect 14360 16880 14400 16885
rect 14440 16915 14480 16920
rect 14440 16885 14445 16915
rect 14475 16885 14480 16915
rect 14440 16880 14480 16885
rect 14520 16915 14560 16920
rect 14520 16885 14525 16915
rect 14555 16885 14560 16915
rect 14520 16880 14560 16885
rect 14600 16915 14640 16920
rect 14600 16885 14605 16915
rect 14635 16885 14640 16915
rect 14600 16880 14640 16885
rect 14680 16915 14720 16920
rect 14680 16885 14685 16915
rect 14715 16885 14720 16915
rect 14680 16880 14720 16885
rect 16760 16915 16800 16920
rect 16760 16885 16765 16915
rect 16795 16885 16800 16915
rect 16760 16880 16800 16885
rect 16840 16915 16880 16920
rect 16840 16885 16845 16915
rect 16875 16885 16880 16915
rect 16840 16880 16880 16885
rect 16920 16915 16960 16920
rect 16920 16885 16925 16915
rect 16955 16885 16960 16915
rect 16920 16880 16960 16885
rect 17000 16915 17040 16920
rect 17000 16885 17005 16915
rect 17035 16885 17040 16915
rect 17000 16880 17040 16885
rect 17080 16915 17120 16920
rect 17080 16885 17085 16915
rect 17115 16885 17120 16915
rect 17080 16880 17120 16885
rect 17160 16915 17200 16920
rect 17160 16885 17165 16915
rect 17195 16885 17200 16915
rect 17160 16880 17200 16885
rect 17240 16915 17280 16920
rect 17240 16885 17245 16915
rect 17275 16885 17280 16915
rect 17240 16880 17280 16885
rect 17320 16915 17360 16920
rect 17320 16885 17325 16915
rect 17355 16885 17360 16915
rect 17320 16880 17360 16885
rect 17400 16915 17440 16920
rect 17400 16885 17405 16915
rect 17435 16885 17440 16915
rect 17400 16880 17440 16885
rect 17480 16915 17520 16920
rect 17480 16885 17485 16915
rect 17515 16885 17520 16915
rect 17480 16880 17520 16885
rect 17560 16915 17600 16920
rect 17560 16885 17565 16915
rect 17595 16885 17600 16915
rect 17560 16880 17600 16885
rect 17640 16915 17680 16920
rect 17640 16885 17645 16915
rect 17675 16885 17680 16915
rect 17640 16880 17680 16885
rect 17720 16915 17760 16920
rect 17720 16885 17725 16915
rect 17755 16885 17760 16915
rect 17720 16880 17760 16885
rect 17800 16915 17840 16920
rect 17800 16885 17805 16915
rect 17835 16885 17840 16915
rect 17800 16880 17840 16885
rect 17880 16915 17920 16920
rect 17880 16885 17885 16915
rect 17915 16885 17920 16915
rect 17880 16880 17920 16885
rect 17960 16915 18000 16920
rect 17960 16885 17965 16915
rect 17995 16885 18000 16915
rect 17960 16880 18000 16885
rect 18040 16915 18080 16920
rect 18040 16885 18045 16915
rect 18075 16885 18080 16915
rect 18040 16880 18080 16885
rect 18120 16915 18160 16920
rect 18120 16885 18125 16915
rect 18155 16885 18160 16915
rect 18120 16880 18160 16885
rect 18200 16915 18240 16920
rect 18200 16885 18205 16915
rect 18235 16885 18240 16915
rect 18200 16880 18240 16885
rect 18280 16915 18320 16920
rect 18280 16885 18285 16915
rect 18315 16885 18320 16915
rect 18280 16880 18320 16885
rect 18360 16915 18400 16920
rect 18360 16885 18365 16915
rect 18395 16885 18400 16915
rect 18360 16880 18400 16885
rect 18440 16915 18480 16920
rect 18440 16885 18445 16915
rect 18475 16885 18480 16915
rect 18440 16880 18480 16885
rect 18520 16915 18560 16920
rect 18520 16885 18525 16915
rect 18555 16885 18560 16915
rect 18520 16880 18560 16885
rect 18600 16915 18640 16920
rect 18600 16885 18605 16915
rect 18635 16885 18640 16915
rect 18600 16880 18640 16885
rect 18680 16915 18720 16920
rect 18680 16885 18685 16915
rect 18715 16885 18720 16915
rect 18680 16880 18720 16885
rect 18760 16915 18800 16920
rect 18760 16885 18765 16915
rect 18795 16885 18800 16915
rect 18760 16880 18800 16885
rect 18840 16915 18880 16920
rect 18840 16885 18845 16915
rect 18875 16885 18880 16915
rect 18840 16880 18880 16885
rect 18920 16915 18960 16920
rect 18920 16885 18925 16915
rect 18955 16885 18960 16915
rect 18920 16880 18960 16885
rect 19000 16915 19040 16920
rect 19000 16885 19005 16915
rect 19035 16885 19040 16915
rect 19000 16880 19040 16885
rect 19080 16915 19120 16920
rect 19080 16885 19085 16915
rect 19115 16885 19120 16915
rect 19080 16880 19120 16885
rect 19160 16915 19200 16920
rect 19160 16885 19165 16915
rect 19195 16885 19200 16915
rect 19160 16880 19200 16885
rect 19240 16915 19280 16920
rect 19240 16885 19245 16915
rect 19275 16885 19280 16915
rect 19240 16880 19280 16885
rect 19320 16915 19360 16920
rect 19320 16885 19325 16915
rect 19355 16885 19360 16915
rect 19320 16880 19360 16885
rect 19400 16915 19440 16920
rect 19400 16885 19405 16915
rect 19435 16885 19440 16915
rect 19400 16880 19440 16885
rect 19480 16915 19520 16920
rect 19480 16885 19485 16915
rect 19515 16885 19520 16915
rect 19480 16880 19520 16885
rect 19560 16915 19600 16920
rect 19560 16885 19565 16915
rect 19595 16885 19600 16915
rect 19560 16880 19600 16885
rect 19640 16915 19680 16920
rect 19640 16885 19645 16915
rect 19675 16885 19680 16915
rect 19640 16880 19680 16885
rect 19720 16915 19760 16920
rect 19720 16885 19725 16915
rect 19755 16885 19760 16915
rect 19720 16880 19760 16885
rect 19800 16915 19840 16920
rect 19800 16885 19805 16915
rect 19835 16885 19840 16915
rect 19800 16880 19840 16885
rect 19880 16915 19920 16920
rect 19880 16885 19885 16915
rect 19915 16885 19920 16915
rect 19880 16880 19920 16885
rect 19960 16915 20000 16920
rect 19960 16885 19965 16915
rect 19995 16885 20000 16915
rect 19960 16880 20000 16885
rect 20040 16915 20080 16920
rect 20040 16885 20045 16915
rect 20075 16885 20080 16915
rect 20040 16880 20080 16885
rect 20120 16915 20160 16920
rect 20120 16885 20125 16915
rect 20155 16885 20160 16915
rect 20120 16880 20160 16885
rect 20200 16915 20240 16920
rect 20200 16885 20205 16915
rect 20235 16885 20240 16915
rect 20200 16880 20240 16885
rect 20280 16915 20320 16920
rect 20280 16885 20285 16915
rect 20315 16885 20320 16915
rect 20280 16880 20320 16885
rect 20360 16915 20400 16920
rect 20360 16885 20365 16915
rect 20395 16885 20400 16915
rect 20360 16880 20400 16885
rect 20440 16915 20480 16920
rect 20440 16885 20445 16915
rect 20475 16885 20480 16915
rect 20440 16880 20480 16885
rect 20520 16915 20560 16920
rect 20520 16885 20525 16915
rect 20555 16885 20560 16915
rect 20520 16880 20560 16885
rect 20600 16915 20640 16920
rect 20600 16885 20605 16915
rect 20635 16885 20640 16915
rect 20600 16880 20640 16885
rect 20680 16915 20720 16920
rect 20680 16885 20685 16915
rect 20715 16885 20720 16915
rect 20680 16880 20720 16885
rect 20760 16915 20800 16920
rect 20760 16885 20765 16915
rect 20795 16885 20800 16915
rect 20760 16880 20800 16885
rect 20840 16915 20880 16920
rect 20840 16885 20845 16915
rect 20875 16885 20880 16915
rect 20840 16880 20880 16885
rect 20920 16915 20960 16920
rect 20920 16885 20925 16915
rect 20955 16885 20960 16915
rect 20920 16880 20960 16885
rect 0 16755 40 16760
rect 0 16725 5 16755
rect 35 16725 40 16755
rect 0 16720 40 16725
rect 80 16755 120 16760
rect 80 16725 85 16755
rect 115 16725 120 16755
rect 80 16720 120 16725
rect 160 16755 200 16760
rect 160 16725 165 16755
rect 195 16725 200 16755
rect 160 16720 200 16725
rect 240 16755 280 16760
rect 240 16725 245 16755
rect 275 16725 280 16755
rect 240 16720 280 16725
rect 320 16755 360 16760
rect 320 16725 325 16755
rect 355 16725 360 16755
rect 320 16720 360 16725
rect 400 16755 440 16760
rect 400 16725 405 16755
rect 435 16725 440 16755
rect 400 16720 440 16725
rect 480 16755 520 16760
rect 480 16725 485 16755
rect 515 16725 520 16755
rect 480 16720 520 16725
rect 560 16755 600 16760
rect 560 16725 565 16755
rect 595 16725 600 16755
rect 560 16720 600 16725
rect 640 16755 680 16760
rect 640 16725 645 16755
rect 675 16725 680 16755
rect 640 16720 680 16725
rect 720 16755 760 16760
rect 720 16725 725 16755
rect 755 16725 760 16755
rect 720 16720 760 16725
rect 800 16755 840 16760
rect 800 16725 805 16755
rect 835 16725 840 16755
rect 800 16720 840 16725
rect 880 16755 920 16760
rect 880 16725 885 16755
rect 915 16725 920 16755
rect 880 16720 920 16725
rect 960 16755 1000 16760
rect 960 16725 965 16755
rect 995 16725 1000 16755
rect 960 16720 1000 16725
rect 1040 16755 1080 16760
rect 1040 16725 1045 16755
rect 1075 16725 1080 16755
rect 1040 16720 1080 16725
rect 1120 16755 1160 16760
rect 1120 16725 1125 16755
rect 1155 16725 1160 16755
rect 1120 16720 1160 16725
rect 1200 16755 1240 16760
rect 1200 16725 1205 16755
rect 1235 16725 1240 16755
rect 1200 16720 1240 16725
rect 1280 16755 1320 16760
rect 1280 16725 1285 16755
rect 1315 16725 1320 16755
rect 1280 16720 1320 16725
rect 1360 16755 1400 16760
rect 1360 16725 1365 16755
rect 1395 16725 1400 16755
rect 1360 16720 1400 16725
rect 1440 16755 1480 16760
rect 1440 16725 1445 16755
rect 1475 16725 1480 16755
rect 1440 16720 1480 16725
rect 1520 16755 1560 16760
rect 1520 16725 1525 16755
rect 1555 16725 1560 16755
rect 1520 16720 1560 16725
rect 1600 16755 1640 16760
rect 1600 16725 1605 16755
rect 1635 16725 1640 16755
rect 1600 16720 1640 16725
rect 1680 16755 1720 16760
rect 1680 16725 1685 16755
rect 1715 16725 1720 16755
rect 1680 16720 1720 16725
rect 1760 16755 1800 16760
rect 1760 16725 1765 16755
rect 1795 16725 1800 16755
rect 1760 16720 1800 16725
rect 1840 16755 1880 16760
rect 1840 16725 1845 16755
rect 1875 16725 1880 16755
rect 1840 16720 1880 16725
rect 1920 16755 1960 16760
rect 1920 16725 1925 16755
rect 1955 16725 1960 16755
rect 1920 16720 1960 16725
rect 2000 16755 2040 16760
rect 2000 16725 2005 16755
rect 2035 16725 2040 16755
rect 2000 16720 2040 16725
rect 2080 16755 2120 16760
rect 2080 16725 2085 16755
rect 2115 16725 2120 16755
rect 2080 16720 2120 16725
rect 2160 16755 2200 16760
rect 2160 16725 2165 16755
rect 2195 16725 2200 16755
rect 2160 16720 2200 16725
rect 2240 16755 2280 16760
rect 2240 16725 2245 16755
rect 2275 16725 2280 16755
rect 2240 16720 2280 16725
rect 2320 16755 2360 16760
rect 2320 16725 2325 16755
rect 2355 16725 2360 16755
rect 2320 16720 2360 16725
rect 2400 16755 2440 16760
rect 2400 16725 2405 16755
rect 2435 16725 2440 16755
rect 2400 16720 2440 16725
rect 2480 16755 2520 16760
rect 2480 16725 2485 16755
rect 2515 16725 2520 16755
rect 2480 16720 2520 16725
rect 2560 16755 2600 16760
rect 2560 16725 2565 16755
rect 2595 16725 2600 16755
rect 2560 16720 2600 16725
rect 2640 16755 2680 16760
rect 2640 16725 2645 16755
rect 2675 16725 2680 16755
rect 2640 16720 2680 16725
rect 2720 16755 2760 16760
rect 2720 16725 2725 16755
rect 2755 16725 2760 16755
rect 2720 16720 2760 16725
rect 2800 16755 2840 16760
rect 2800 16725 2805 16755
rect 2835 16725 2840 16755
rect 2800 16720 2840 16725
rect 2880 16755 2920 16760
rect 2880 16725 2885 16755
rect 2915 16725 2920 16755
rect 2880 16720 2920 16725
rect 2960 16755 3000 16760
rect 2960 16725 2965 16755
rect 2995 16725 3000 16755
rect 2960 16720 3000 16725
rect 3040 16755 3080 16760
rect 3040 16725 3045 16755
rect 3075 16725 3080 16755
rect 3040 16720 3080 16725
rect 3120 16755 3160 16760
rect 3120 16725 3125 16755
rect 3155 16725 3160 16755
rect 3120 16720 3160 16725
rect 3200 16755 3240 16760
rect 3200 16725 3205 16755
rect 3235 16725 3240 16755
rect 3200 16720 3240 16725
rect 3280 16755 3320 16760
rect 3280 16725 3285 16755
rect 3315 16725 3320 16755
rect 3280 16720 3320 16725
rect 3360 16755 3400 16760
rect 3360 16725 3365 16755
rect 3395 16725 3400 16755
rect 3360 16720 3400 16725
rect 3440 16755 3480 16760
rect 3440 16725 3445 16755
rect 3475 16725 3480 16755
rect 3440 16720 3480 16725
rect 3520 16755 3560 16760
rect 3520 16725 3525 16755
rect 3555 16725 3560 16755
rect 3520 16720 3560 16725
rect 3600 16755 3640 16760
rect 3600 16725 3605 16755
rect 3635 16725 3640 16755
rect 3600 16720 3640 16725
rect 3680 16755 3720 16760
rect 3680 16725 3685 16755
rect 3715 16725 3720 16755
rect 3680 16720 3720 16725
rect 3760 16755 3800 16760
rect 3760 16725 3765 16755
rect 3795 16725 3800 16755
rect 3760 16720 3800 16725
rect 3840 16755 3880 16760
rect 3840 16725 3845 16755
rect 3875 16725 3880 16755
rect 3840 16720 3880 16725
rect 3920 16755 3960 16760
rect 3920 16725 3925 16755
rect 3955 16725 3960 16755
rect 3920 16720 3960 16725
rect 4000 16755 4040 16760
rect 4000 16725 4005 16755
rect 4035 16725 4040 16755
rect 4000 16720 4040 16725
rect 4080 16755 4120 16760
rect 4080 16725 4085 16755
rect 4115 16725 4120 16755
rect 4080 16720 4120 16725
rect 4160 16755 4200 16760
rect 4160 16725 4165 16755
rect 4195 16725 4200 16755
rect 4160 16720 4200 16725
rect 6240 16755 6280 16760
rect 6240 16725 6245 16755
rect 6275 16725 6280 16755
rect 6240 16720 6280 16725
rect 6320 16755 6360 16760
rect 6320 16725 6325 16755
rect 6355 16725 6360 16755
rect 6320 16720 6360 16725
rect 6400 16755 6440 16760
rect 6400 16725 6405 16755
rect 6435 16725 6440 16755
rect 6400 16720 6440 16725
rect 6480 16755 6520 16760
rect 6480 16725 6485 16755
rect 6515 16725 6520 16755
rect 6480 16720 6520 16725
rect 6560 16755 6600 16760
rect 6560 16725 6565 16755
rect 6595 16725 6600 16755
rect 6560 16720 6600 16725
rect 6640 16755 6680 16760
rect 6640 16725 6645 16755
rect 6675 16725 6680 16755
rect 6640 16720 6680 16725
rect 6720 16755 6760 16760
rect 6720 16725 6725 16755
rect 6755 16725 6760 16755
rect 6720 16720 6760 16725
rect 6800 16755 6840 16760
rect 6800 16725 6805 16755
rect 6835 16725 6840 16755
rect 6800 16720 6840 16725
rect 6880 16755 6920 16760
rect 6880 16725 6885 16755
rect 6915 16725 6920 16755
rect 6880 16720 6920 16725
rect 6960 16755 7000 16760
rect 6960 16725 6965 16755
rect 6995 16725 7000 16755
rect 6960 16720 7000 16725
rect 7040 16755 7080 16760
rect 7040 16725 7045 16755
rect 7075 16725 7080 16755
rect 7040 16720 7080 16725
rect 7120 16755 7160 16760
rect 7120 16725 7125 16755
rect 7155 16725 7160 16755
rect 7120 16720 7160 16725
rect 7200 16755 7240 16760
rect 7200 16725 7205 16755
rect 7235 16725 7240 16755
rect 7200 16720 7240 16725
rect 7280 16755 7320 16760
rect 7280 16725 7285 16755
rect 7315 16725 7320 16755
rect 7280 16720 7320 16725
rect 7360 16755 7400 16760
rect 7360 16725 7365 16755
rect 7395 16725 7400 16755
rect 7360 16720 7400 16725
rect 7440 16755 7480 16760
rect 7440 16725 7445 16755
rect 7475 16725 7480 16755
rect 7440 16720 7480 16725
rect 7520 16755 7560 16760
rect 7520 16725 7525 16755
rect 7555 16725 7560 16755
rect 7520 16720 7560 16725
rect 7600 16755 7640 16760
rect 7600 16725 7605 16755
rect 7635 16725 7640 16755
rect 7600 16720 7640 16725
rect 7680 16755 7720 16760
rect 7680 16725 7685 16755
rect 7715 16725 7720 16755
rect 7680 16720 7720 16725
rect 7760 16755 7800 16760
rect 7760 16725 7765 16755
rect 7795 16725 7800 16755
rect 7760 16720 7800 16725
rect 7840 16755 7880 16760
rect 7840 16725 7845 16755
rect 7875 16725 7880 16755
rect 7840 16720 7880 16725
rect 7920 16755 7960 16760
rect 7920 16725 7925 16755
rect 7955 16725 7960 16755
rect 7920 16720 7960 16725
rect 8000 16755 8040 16760
rect 8000 16725 8005 16755
rect 8035 16725 8040 16755
rect 8000 16720 8040 16725
rect 8080 16755 8120 16760
rect 8080 16725 8085 16755
rect 8115 16725 8120 16755
rect 8080 16720 8120 16725
rect 8160 16755 8200 16760
rect 8160 16725 8165 16755
rect 8195 16725 8200 16755
rect 8160 16720 8200 16725
rect 8240 16755 8280 16760
rect 8240 16725 8245 16755
rect 8275 16725 8280 16755
rect 8240 16720 8280 16725
rect 8320 16755 8360 16760
rect 8320 16725 8325 16755
rect 8355 16725 8360 16755
rect 8320 16720 8360 16725
rect 8400 16755 8440 16760
rect 8400 16725 8405 16755
rect 8435 16725 8440 16755
rect 8400 16720 8440 16725
rect 8480 16755 8520 16760
rect 8480 16725 8485 16755
rect 8515 16725 8520 16755
rect 8480 16720 8520 16725
rect 8560 16755 8600 16760
rect 8560 16725 8565 16755
rect 8595 16725 8600 16755
rect 8560 16720 8600 16725
rect 8640 16755 8680 16760
rect 8640 16725 8645 16755
rect 8675 16725 8680 16755
rect 8640 16720 8680 16725
rect 8720 16755 8760 16760
rect 8720 16725 8725 16755
rect 8755 16725 8760 16755
rect 8720 16720 8760 16725
rect 8800 16755 8840 16760
rect 8800 16725 8805 16755
rect 8835 16725 8840 16755
rect 8800 16720 8840 16725
rect 8880 16755 8920 16760
rect 8880 16725 8885 16755
rect 8915 16725 8920 16755
rect 8880 16720 8920 16725
rect 8960 16755 9000 16760
rect 8960 16725 8965 16755
rect 8995 16725 9000 16755
rect 8960 16720 9000 16725
rect 9040 16755 9080 16760
rect 9040 16725 9045 16755
rect 9075 16725 9080 16755
rect 9040 16720 9080 16725
rect 9120 16755 9160 16760
rect 9120 16725 9125 16755
rect 9155 16725 9160 16755
rect 9120 16720 9160 16725
rect 9200 16755 9240 16760
rect 9200 16725 9205 16755
rect 9235 16725 9240 16755
rect 9200 16720 9240 16725
rect 9280 16755 9320 16760
rect 9280 16725 9285 16755
rect 9315 16725 9320 16755
rect 9280 16720 9320 16725
rect 9360 16755 9400 16760
rect 9360 16725 9365 16755
rect 9395 16725 9400 16755
rect 9360 16720 9400 16725
rect 9440 16755 9480 16760
rect 9440 16725 9445 16755
rect 9475 16725 9480 16755
rect 9440 16720 9480 16725
rect 11560 16755 11600 16760
rect 11560 16725 11565 16755
rect 11595 16725 11600 16755
rect 11560 16720 11600 16725
rect 11640 16755 11680 16760
rect 11640 16725 11645 16755
rect 11675 16725 11680 16755
rect 11640 16720 11680 16725
rect 11720 16755 11760 16760
rect 11720 16725 11725 16755
rect 11755 16725 11760 16755
rect 11720 16720 11760 16725
rect 11800 16755 11840 16760
rect 11800 16725 11805 16755
rect 11835 16725 11840 16755
rect 11800 16720 11840 16725
rect 11880 16755 11920 16760
rect 11880 16725 11885 16755
rect 11915 16725 11920 16755
rect 11880 16720 11920 16725
rect 11960 16755 12000 16760
rect 11960 16725 11965 16755
rect 11995 16725 12000 16755
rect 11960 16720 12000 16725
rect 12040 16755 12080 16760
rect 12040 16725 12045 16755
rect 12075 16725 12080 16755
rect 12040 16720 12080 16725
rect 12120 16755 12160 16760
rect 12120 16725 12125 16755
rect 12155 16725 12160 16755
rect 12120 16720 12160 16725
rect 12200 16755 12240 16760
rect 12200 16725 12205 16755
rect 12235 16725 12240 16755
rect 12200 16720 12240 16725
rect 12280 16755 12320 16760
rect 12280 16725 12285 16755
rect 12315 16725 12320 16755
rect 12280 16720 12320 16725
rect 12360 16755 12400 16760
rect 12360 16725 12365 16755
rect 12395 16725 12400 16755
rect 12360 16720 12400 16725
rect 12440 16755 12480 16760
rect 12440 16725 12445 16755
rect 12475 16725 12480 16755
rect 12440 16720 12480 16725
rect 12520 16755 12560 16760
rect 12520 16725 12525 16755
rect 12555 16725 12560 16755
rect 12520 16720 12560 16725
rect 12600 16755 12640 16760
rect 12600 16725 12605 16755
rect 12635 16725 12640 16755
rect 12600 16720 12640 16725
rect 12680 16755 12720 16760
rect 12680 16725 12685 16755
rect 12715 16725 12720 16755
rect 12680 16720 12720 16725
rect 12760 16755 12800 16760
rect 12760 16725 12765 16755
rect 12795 16725 12800 16755
rect 12760 16720 12800 16725
rect 12840 16755 12880 16760
rect 12840 16725 12845 16755
rect 12875 16725 12880 16755
rect 12840 16720 12880 16725
rect 12920 16755 12960 16760
rect 12920 16725 12925 16755
rect 12955 16725 12960 16755
rect 12920 16720 12960 16725
rect 13000 16755 13040 16760
rect 13000 16725 13005 16755
rect 13035 16725 13040 16755
rect 13000 16720 13040 16725
rect 13080 16755 13120 16760
rect 13080 16725 13085 16755
rect 13115 16725 13120 16755
rect 13080 16720 13120 16725
rect 13160 16755 13200 16760
rect 13160 16725 13165 16755
rect 13195 16725 13200 16755
rect 13160 16720 13200 16725
rect 13240 16755 13280 16760
rect 13240 16725 13245 16755
rect 13275 16725 13280 16755
rect 13240 16720 13280 16725
rect 13320 16755 13360 16760
rect 13320 16725 13325 16755
rect 13355 16725 13360 16755
rect 13320 16720 13360 16725
rect 13400 16755 13440 16760
rect 13400 16725 13405 16755
rect 13435 16725 13440 16755
rect 13400 16720 13440 16725
rect 13480 16755 13520 16760
rect 13480 16725 13485 16755
rect 13515 16725 13520 16755
rect 13480 16720 13520 16725
rect 13560 16755 13600 16760
rect 13560 16725 13565 16755
rect 13595 16725 13600 16755
rect 13560 16720 13600 16725
rect 13640 16755 13680 16760
rect 13640 16725 13645 16755
rect 13675 16725 13680 16755
rect 13640 16720 13680 16725
rect 13720 16755 13760 16760
rect 13720 16725 13725 16755
rect 13755 16725 13760 16755
rect 13720 16720 13760 16725
rect 13800 16755 13840 16760
rect 13800 16725 13805 16755
rect 13835 16725 13840 16755
rect 13800 16720 13840 16725
rect 13880 16755 13920 16760
rect 13880 16725 13885 16755
rect 13915 16725 13920 16755
rect 13880 16720 13920 16725
rect 13960 16755 14000 16760
rect 13960 16725 13965 16755
rect 13995 16725 14000 16755
rect 13960 16720 14000 16725
rect 14040 16755 14080 16760
rect 14040 16725 14045 16755
rect 14075 16725 14080 16755
rect 14040 16720 14080 16725
rect 14120 16755 14160 16760
rect 14120 16725 14125 16755
rect 14155 16725 14160 16755
rect 14120 16720 14160 16725
rect 14200 16755 14240 16760
rect 14200 16725 14205 16755
rect 14235 16725 14240 16755
rect 14200 16720 14240 16725
rect 14280 16755 14320 16760
rect 14280 16725 14285 16755
rect 14315 16725 14320 16755
rect 14280 16720 14320 16725
rect 14360 16755 14400 16760
rect 14360 16725 14365 16755
rect 14395 16725 14400 16755
rect 14360 16720 14400 16725
rect 14440 16755 14480 16760
rect 14440 16725 14445 16755
rect 14475 16725 14480 16755
rect 14440 16720 14480 16725
rect 14520 16755 14560 16760
rect 14520 16725 14525 16755
rect 14555 16725 14560 16755
rect 14520 16720 14560 16725
rect 14600 16755 14640 16760
rect 14600 16725 14605 16755
rect 14635 16725 14640 16755
rect 14600 16720 14640 16725
rect 14680 16755 14720 16760
rect 14680 16725 14685 16755
rect 14715 16725 14720 16755
rect 14680 16720 14720 16725
rect 16760 16755 16800 16760
rect 16760 16725 16765 16755
rect 16795 16725 16800 16755
rect 16760 16720 16800 16725
rect 16840 16755 16880 16760
rect 16840 16725 16845 16755
rect 16875 16725 16880 16755
rect 16840 16720 16880 16725
rect 16920 16755 16960 16760
rect 16920 16725 16925 16755
rect 16955 16725 16960 16755
rect 16920 16720 16960 16725
rect 17000 16755 17040 16760
rect 17000 16725 17005 16755
rect 17035 16725 17040 16755
rect 17000 16720 17040 16725
rect 17080 16755 17120 16760
rect 17080 16725 17085 16755
rect 17115 16725 17120 16755
rect 17080 16720 17120 16725
rect 17160 16755 17200 16760
rect 17160 16725 17165 16755
rect 17195 16725 17200 16755
rect 17160 16720 17200 16725
rect 17240 16755 17280 16760
rect 17240 16725 17245 16755
rect 17275 16725 17280 16755
rect 17240 16720 17280 16725
rect 17320 16755 17360 16760
rect 17320 16725 17325 16755
rect 17355 16725 17360 16755
rect 17320 16720 17360 16725
rect 17400 16755 17440 16760
rect 17400 16725 17405 16755
rect 17435 16725 17440 16755
rect 17400 16720 17440 16725
rect 17480 16755 17520 16760
rect 17480 16725 17485 16755
rect 17515 16725 17520 16755
rect 17480 16720 17520 16725
rect 17560 16755 17600 16760
rect 17560 16725 17565 16755
rect 17595 16725 17600 16755
rect 17560 16720 17600 16725
rect 17640 16755 17680 16760
rect 17640 16725 17645 16755
rect 17675 16725 17680 16755
rect 17640 16720 17680 16725
rect 17720 16755 17760 16760
rect 17720 16725 17725 16755
rect 17755 16725 17760 16755
rect 17720 16720 17760 16725
rect 17800 16755 17840 16760
rect 17800 16725 17805 16755
rect 17835 16725 17840 16755
rect 17800 16720 17840 16725
rect 17880 16755 17920 16760
rect 17880 16725 17885 16755
rect 17915 16725 17920 16755
rect 17880 16720 17920 16725
rect 17960 16755 18000 16760
rect 17960 16725 17965 16755
rect 17995 16725 18000 16755
rect 17960 16720 18000 16725
rect 18040 16755 18080 16760
rect 18040 16725 18045 16755
rect 18075 16725 18080 16755
rect 18040 16720 18080 16725
rect 18120 16755 18160 16760
rect 18120 16725 18125 16755
rect 18155 16725 18160 16755
rect 18120 16720 18160 16725
rect 18200 16755 18240 16760
rect 18200 16725 18205 16755
rect 18235 16725 18240 16755
rect 18200 16720 18240 16725
rect 18280 16755 18320 16760
rect 18280 16725 18285 16755
rect 18315 16725 18320 16755
rect 18280 16720 18320 16725
rect 18360 16755 18400 16760
rect 18360 16725 18365 16755
rect 18395 16725 18400 16755
rect 18360 16720 18400 16725
rect 18440 16755 18480 16760
rect 18440 16725 18445 16755
rect 18475 16725 18480 16755
rect 18440 16720 18480 16725
rect 18520 16755 18560 16760
rect 18520 16725 18525 16755
rect 18555 16725 18560 16755
rect 18520 16720 18560 16725
rect 18600 16755 18640 16760
rect 18600 16725 18605 16755
rect 18635 16725 18640 16755
rect 18600 16720 18640 16725
rect 18680 16755 18720 16760
rect 18680 16725 18685 16755
rect 18715 16725 18720 16755
rect 18680 16720 18720 16725
rect 18760 16755 18800 16760
rect 18760 16725 18765 16755
rect 18795 16725 18800 16755
rect 18760 16720 18800 16725
rect 18840 16755 18880 16760
rect 18840 16725 18845 16755
rect 18875 16725 18880 16755
rect 18840 16720 18880 16725
rect 18920 16755 18960 16760
rect 18920 16725 18925 16755
rect 18955 16725 18960 16755
rect 18920 16720 18960 16725
rect 19000 16755 19040 16760
rect 19000 16725 19005 16755
rect 19035 16725 19040 16755
rect 19000 16720 19040 16725
rect 19080 16755 19120 16760
rect 19080 16725 19085 16755
rect 19115 16725 19120 16755
rect 19080 16720 19120 16725
rect 19160 16755 19200 16760
rect 19160 16725 19165 16755
rect 19195 16725 19200 16755
rect 19160 16720 19200 16725
rect 19240 16755 19280 16760
rect 19240 16725 19245 16755
rect 19275 16725 19280 16755
rect 19240 16720 19280 16725
rect 19320 16755 19360 16760
rect 19320 16725 19325 16755
rect 19355 16725 19360 16755
rect 19320 16720 19360 16725
rect 19400 16755 19440 16760
rect 19400 16725 19405 16755
rect 19435 16725 19440 16755
rect 19400 16720 19440 16725
rect 19480 16755 19520 16760
rect 19480 16725 19485 16755
rect 19515 16725 19520 16755
rect 19480 16720 19520 16725
rect 19560 16755 19600 16760
rect 19560 16725 19565 16755
rect 19595 16725 19600 16755
rect 19560 16720 19600 16725
rect 19640 16755 19680 16760
rect 19640 16725 19645 16755
rect 19675 16725 19680 16755
rect 19640 16720 19680 16725
rect 19720 16755 19760 16760
rect 19720 16725 19725 16755
rect 19755 16725 19760 16755
rect 19720 16720 19760 16725
rect 19800 16755 19840 16760
rect 19800 16725 19805 16755
rect 19835 16725 19840 16755
rect 19800 16720 19840 16725
rect 19880 16755 19920 16760
rect 19880 16725 19885 16755
rect 19915 16725 19920 16755
rect 19880 16720 19920 16725
rect 19960 16755 20000 16760
rect 19960 16725 19965 16755
rect 19995 16725 20000 16755
rect 19960 16720 20000 16725
rect 20040 16755 20080 16760
rect 20040 16725 20045 16755
rect 20075 16725 20080 16755
rect 20040 16720 20080 16725
rect 20120 16755 20160 16760
rect 20120 16725 20125 16755
rect 20155 16725 20160 16755
rect 20120 16720 20160 16725
rect 20200 16755 20240 16760
rect 20200 16725 20205 16755
rect 20235 16725 20240 16755
rect 20200 16720 20240 16725
rect 20280 16755 20320 16760
rect 20280 16725 20285 16755
rect 20315 16725 20320 16755
rect 20280 16720 20320 16725
rect 20360 16755 20400 16760
rect 20360 16725 20365 16755
rect 20395 16725 20400 16755
rect 20360 16720 20400 16725
rect 20440 16755 20480 16760
rect 20440 16725 20445 16755
rect 20475 16725 20480 16755
rect 20440 16720 20480 16725
rect 20520 16755 20560 16760
rect 20520 16725 20525 16755
rect 20555 16725 20560 16755
rect 20520 16720 20560 16725
rect 20600 16755 20640 16760
rect 20600 16725 20605 16755
rect 20635 16725 20640 16755
rect 20600 16720 20640 16725
rect 20680 16755 20720 16760
rect 20680 16725 20685 16755
rect 20715 16725 20720 16755
rect 20680 16720 20720 16725
rect 20760 16755 20800 16760
rect 20760 16725 20765 16755
rect 20795 16725 20800 16755
rect 20760 16720 20800 16725
rect 20840 16755 20880 16760
rect 20840 16725 20845 16755
rect 20875 16725 20880 16755
rect 20840 16720 20880 16725
rect 20920 16755 20960 16760
rect 20920 16725 20925 16755
rect 20955 16725 20960 16755
rect 20920 16720 20960 16725
rect 0 16675 40 16680
rect 0 16645 5 16675
rect 35 16645 40 16675
rect 0 16640 40 16645
rect 80 16675 120 16680
rect 80 16645 85 16675
rect 115 16645 120 16675
rect 80 16640 120 16645
rect 160 16675 200 16680
rect 160 16645 165 16675
rect 195 16645 200 16675
rect 160 16640 200 16645
rect 240 16675 280 16680
rect 240 16645 245 16675
rect 275 16645 280 16675
rect 240 16640 280 16645
rect 320 16675 360 16680
rect 320 16645 325 16675
rect 355 16645 360 16675
rect 320 16640 360 16645
rect 400 16675 440 16680
rect 400 16645 405 16675
rect 435 16645 440 16675
rect 400 16640 440 16645
rect 480 16675 520 16680
rect 480 16645 485 16675
rect 515 16645 520 16675
rect 480 16640 520 16645
rect 560 16675 600 16680
rect 560 16645 565 16675
rect 595 16645 600 16675
rect 560 16640 600 16645
rect 640 16675 680 16680
rect 640 16645 645 16675
rect 675 16645 680 16675
rect 640 16640 680 16645
rect 720 16675 760 16680
rect 720 16645 725 16675
rect 755 16645 760 16675
rect 720 16640 760 16645
rect 800 16675 840 16680
rect 800 16645 805 16675
rect 835 16645 840 16675
rect 800 16640 840 16645
rect 880 16675 920 16680
rect 880 16645 885 16675
rect 915 16645 920 16675
rect 880 16640 920 16645
rect 960 16675 1000 16680
rect 960 16645 965 16675
rect 995 16645 1000 16675
rect 960 16640 1000 16645
rect 1040 16675 1080 16680
rect 1040 16645 1045 16675
rect 1075 16645 1080 16675
rect 1040 16640 1080 16645
rect 1120 16675 1160 16680
rect 1120 16645 1125 16675
rect 1155 16645 1160 16675
rect 1120 16640 1160 16645
rect 1200 16675 1240 16680
rect 1200 16645 1205 16675
rect 1235 16645 1240 16675
rect 1200 16640 1240 16645
rect 1280 16675 1320 16680
rect 1280 16645 1285 16675
rect 1315 16645 1320 16675
rect 1280 16640 1320 16645
rect 1360 16675 1400 16680
rect 1360 16645 1365 16675
rect 1395 16645 1400 16675
rect 1360 16640 1400 16645
rect 1440 16675 1480 16680
rect 1440 16645 1445 16675
rect 1475 16645 1480 16675
rect 1440 16640 1480 16645
rect 1520 16675 1560 16680
rect 1520 16645 1525 16675
rect 1555 16645 1560 16675
rect 1520 16640 1560 16645
rect 1600 16675 1640 16680
rect 1600 16645 1605 16675
rect 1635 16645 1640 16675
rect 1600 16640 1640 16645
rect 1680 16675 1720 16680
rect 1680 16645 1685 16675
rect 1715 16645 1720 16675
rect 1680 16640 1720 16645
rect 1760 16675 1800 16680
rect 1760 16645 1765 16675
rect 1795 16645 1800 16675
rect 1760 16640 1800 16645
rect 1840 16675 1880 16680
rect 1840 16645 1845 16675
rect 1875 16645 1880 16675
rect 1840 16640 1880 16645
rect 1920 16675 1960 16680
rect 1920 16645 1925 16675
rect 1955 16645 1960 16675
rect 1920 16640 1960 16645
rect 2000 16675 2040 16680
rect 2000 16645 2005 16675
rect 2035 16645 2040 16675
rect 2000 16640 2040 16645
rect 2080 16675 2120 16680
rect 2080 16645 2085 16675
rect 2115 16645 2120 16675
rect 2080 16640 2120 16645
rect 2160 16675 2200 16680
rect 2160 16645 2165 16675
rect 2195 16645 2200 16675
rect 2160 16640 2200 16645
rect 2240 16675 2280 16680
rect 2240 16645 2245 16675
rect 2275 16645 2280 16675
rect 2240 16640 2280 16645
rect 2320 16675 2360 16680
rect 2320 16645 2325 16675
rect 2355 16645 2360 16675
rect 2320 16640 2360 16645
rect 2400 16675 2440 16680
rect 2400 16645 2405 16675
rect 2435 16645 2440 16675
rect 2400 16640 2440 16645
rect 2480 16675 2520 16680
rect 2480 16645 2485 16675
rect 2515 16645 2520 16675
rect 2480 16640 2520 16645
rect 2560 16675 2600 16680
rect 2560 16645 2565 16675
rect 2595 16645 2600 16675
rect 2560 16640 2600 16645
rect 2640 16675 2680 16680
rect 2640 16645 2645 16675
rect 2675 16645 2680 16675
rect 2640 16640 2680 16645
rect 2720 16675 2760 16680
rect 2720 16645 2725 16675
rect 2755 16645 2760 16675
rect 2720 16640 2760 16645
rect 2800 16675 2840 16680
rect 2800 16645 2805 16675
rect 2835 16645 2840 16675
rect 2800 16640 2840 16645
rect 2880 16675 2920 16680
rect 2880 16645 2885 16675
rect 2915 16645 2920 16675
rect 2880 16640 2920 16645
rect 2960 16675 3000 16680
rect 2960 16645 2965 16675
rect 2995 16645 3000 16675
rect 2960 16640 3000 16645
rect 3040 16675 3080 16680
rect 3040 16645 3045 16675
rect 3075 16645 3080 16675
rect 3040 16640 3080 16645
rect 3120 16675 3160 16680
rect 3120 16645 3125 16675
rect 3155 16645 3160 16675
rect 3120 16640 3160 16645
rect 3200 16675 3240 16680
rect 3200 16645 3205 16675
rect 3235 16645 3240 16675
rect 3200 16640 3240 16645
rect 3280 16675 3320 16680
rect 3280 16645 3285 16675
rect 3315 16645 3320 16675
rect 3280 16640 3320 16645
rect 3360 16675 3400 16680
rect 3360 16645 3365 16675
rect 3395 16645 3400 16675
rect 3360 16640 3400 16645
rect 3440 16675 3480 16680
rect 3440 16645 3445 16675
rect 3475 16645 3480 16675
rect 3440 16640 3480 16645
rect 3520 16675 3560 16680
rect 3520 16645 3525 16675
rect 3555 16645 3560 16675
rect 3520 16640 3560 16645
rect 3600 16675 3640 16680
rect 3600 16645 3605 16675
rect 3635 16645 3640 16675
rect 3600 16640 3640 16645
rect 3680 16675 3720 16680
rect 3680 16645 3685 16675
rect 3715 16645 3720 16675
rect 3680 16640 3720 16645
rect 3760 16675 3800 16680
rect 3760 16645 3765 16675
rect 3795 16645 3800 16675
rect 3760 16640 3800 16645
rect 3840 16675 3880 16680
rect 3840 16645 3845 16675
rect 3875 16645 3880 16675
rect 3840 16640 3880 16645
rect 3920 16675 3960 16680
rect 3920 16645 3925 16675
rect 3955 16645 3960 16675
rect 3920 16640 3960 16645
rect 4000 16675 4040 16680
rect 4000 16645 4005 16675
rect 4035 16645 4040 16675
rect 4000 16640 4040 16645
rect 4080 16675 4120 16680
rect 4080 16645 4085 16675
rect 4115 16645 4120 16675
rect 4080 16640 4120 16645
rect 4160 16675 4200 16680
rect 4160 16645 4165 16675
rect 4195 16645 4200 16675
rect 4160 16640 4200 16645
rect 6240 16675 6280 16680
rect 6240 16645 6245 16675
rect 6275 16645 6280 16675
rect 6240 16640 6280 16645
rect 6320 16675 6360 16680
rect 6320 16645 6325 16675
rect 6355 16645 6360 16675
rect 6320 16640 6360 16645
rect 6400 16675 6440 16680
rect 6400 16645 6405 16675
rect 6435 16645 6440 16675
rect 6400 16640 6440 16645
rect 6480 16675 6520 16680
rect 6480 16645 6485 16675
rect 6515 16645 6520 16675
rect 6480 16640 6520 16645
rect 6560 16675 6600 16680
rect 6560 16645 6565 16675
rect 6595 16645 6600 16675
rect 6560 16640 6600 16645
rect 6640 16675 6680 16680
rect 6640 16645 6645 16675
rect 6675 16645 6680 16675
rect 6640 16640 6680 16645
rect 6720 16675 6760 16680
rect 6720 16645 6725 16675
rect 6755 16645 6760 16675
rect 6720 16640 6760 16645
rect 6800 16675 6840 16680
rect 6800 16645 6805 16675
rect 6835 16645 6840 16675
rect 6800 16640 6840 16645
rect 6880 16675 6920 16680
rect 6880 16645 6885 16675
rect 6915 16645 6920 16675
rect 6880 16640 6920 16645
rect 6960 16675 7000 16680
rect 6960 16645 6965 16675
rect 6995 16645 7000 16675
rect 6960 16640 7000 16645
rect 7040 16675 7080 16680
rect 7040 16645 7045 16675
rect 7075 16645 7080 16675
rect 7040 16640 7080 16645
rect 7120 16675 7160 16680
rect 7120 16645 7125 16675
rect 7155 16645 7160 16675
rect 7120 16640 7160 16645
rect 7200 16675 7240 16680
rect 7200 16645 7205 16675
rect 7235 16645 7240 16675
rect 7200 16640 7240 16645
rect 7280 16675 7320 16680
rect 7280 16645 7285 16675
rect 7315 16645 7320 16675
rect 7280 16640 7320 16645
rect 7360 16675 7400 16680
rect 7360 16645 7365 16675
rect 7395 16645 7400 16675
rect 7360 16640 7400 16645
rect 7440 16675 7480 16680
rect 7440 16645 7445 16675
rect 7475 16645 7480 16675
rect 7440 16640 7480 16645
rect 7520 16675 7560 16680
rect 7520 16645 7525 16675
rect 7555 16645 7560 16675
rect 7520 16640 7560 16645
rect 7600 16675 7640 16680
rect 7600 16645 7605 16675
rect 7635 16645 7640 16675
rect 7600 16640 7640 16645
rect 7680 16675 7720 16680
rect 7680 16645 7685 16675
rect 7715 16645 7720 16675
rect 7680 16640 7720 16645
rect 7760 16675 7800 16680
rect 7760 16645 7765 16675
rect 7795 16645 7800 16675
rect 7760 16640 7800 16645
rect 7840 16675 7880 16680
rect 7840 16645 7845 16675
rect 7875 16645 7880 16675
rect 7840 16640 7880 16645
rect 7920 16675 7960 16680
rect 7920 16645 7925 16675
rect 7955 16645 7960 16675
rect 7920 16640 7960 16645
rect 8000 16675 8040 16680
rect 8000 16645 8005 16675
rect 8035 16645 8040 16675
rect 8000 16640 8040 16645
rect 8080 16675 8120 16680
rect 8080 16645 8085 16675
rect 8115 16645 8120 16675
rect 8080 16640 8120 16645
rect 8160 16675 8200 16680
rect 8160 16645 8165 16675
rect 8195 16645 8200 16675
rect 8160 16640 8200 16645
rect 8240 16675 8280 16680
rect 8240 16645 8245 16675
rect 8275 16645 8280 16675
rect 8240 16640 8280 16645
rect 8320 16675 8360 16680
rect 8320 16645 8325 16675
rect 8355 16645 8360 16675
rect 8320 16640 8360 16645
rect 8400 16675 8440 16680
rect 8400 16645 8405 16675
rect 8435 16645 8440 16675
rect 8400 16640 8440 16645
rect 8480 16675 8520 16680
rect 8480 16645 8485 16675
rect 8515 16645 8520 16675
rect 8480 16640 8520 16645
rect 8560 16675 8600 16680
rect 8560 16645 8565 16675
rect 8595 16645 8600 16675
rect 8560 16640 8600 16645
rect 8640 16675 8680 16680
rect 8640 16645 8645 16675
rect 8675 16645 8680 16675
rect 8640 16640 8680 16645
rect 8720 16675 8760 16680
rect 8720 16645 8725 16675
rect 8755 16645 8760 16675
rect 8720 16640 8760 16645
rect 8800 16675 8840 16680
rect 8800 16645 8805 16675
rect 8835 16645 8840 16675
rect 8800 16640 8840 16645
rect 8880 16675 8920 16680
rect 8880 16645 8885 16675
rect 8915 16645 8920 16675
rect 8880 16640 8920 16645
rect 8960 16675 9000 16680
rect 8960 16645 8965 16675
rect 8995 16645 9000 16675
rect 8960 16640 9000 16645
rect 9040 16675 9080 16680
rect 9040 16645 9045 16675
rect 9075 16645 9080 16675
rect 9040 16640 9080 16645
rect 9120 16675 9160 16680
rect 9120 16645 9125 16675
rect 9155 16645 9160 16675
rect 9120 16640 9160 16645
rect 9200 16675 9240 16680
rect 9200 16645 9205 16675
rect 9235 16645 9240 16675
rect 9200 16640 9240 16645
rect 9280 16675 9320 16680
rect 9280 16645 9285 16675
rect 9315 16645 9320 16675
rect 9280 16640 9320 16645
rect 9360 16675 9400 16680
rect 9360 16645 9365 16675
rect 9395 16645 9400 16675
rect 9360 16640 9400 16645
rect 9440 16675 9480 16680
rect 9440 16645 9445 16675
rect 9475 16645 9480 16675
rect 9440 16640 9480 16645
rect 11560 16675 11600 16680
rect 11560 16645 11565 16675
rect 11595 16645 11600 16675
rect 11560 16640 11600 16645
rect 11640 16675 11680 16680
rect 11640 16645 11645 16675
rect 11675 16645 11680 16675
rect 11640 16640 11680 16645
rect 11720 16675 11760 16680
rect 11720 16645 11725 16675
rect 11755 16645 11760 16675
rect 11720 16640 11760 16645
rect 11800 16675 11840 16680
rect 11800 16645 11805 16675
rect 11835 16645 11840 16675
rect 11800 16640 11840 16645
rect 11880 16675 11920 16680
rect 11880 16645 11885 16675
rect 11915 16645 11920 16675
rect 11880 16640 11920 16645
rect 11960 16675 12000 16680
rect 11960 16645 11965 16675
rect 11995 16645 12000 16675
rect 11960 16640 12000 16645
rect 12040 16675 12080 16680
rect 12040 16645 12045 16675
rect 12075 16645 12080 16675
rect 12040 16640 12080 16645
rect 12120 16675 12160 16680
rect 12120 16645 12125 16675
rect 12155 16645 12160 16675
rect 12120 16640 12160 16645
rect 12200 16675 12240 16680
rect 12200 16645 12205 16675
rect 12235 16645 12240 16675
rect 12200 16640 12240 16645
rect 12280 16675 12320 16680
rect 12280 16645 12285 16675
rect 12315 16645 12320 16675
rect 12280 16640 12320 16645
rect 12360 16675 12400 16680
rect 12360 16645 12365 16675
rect 12395 16645 12400 16675
rect 12360 16640 12400 16645
rect 12440 16675 12480 16680
rect 12440 16645 12445 16675
rect 12475 16645 12480 16675
rect 12440 16640 12480 16645
rect 12520 16675 12560 16680
rect 12520 16645 12525 16675
rect 12555 16645 12560 16675
rect 12520 16640 12560 16645
rect 12600 16675 12640 16680
rect 12600 16645 12605 16675
rect 12635 16645 12640 16675
rect 12600 16640 12640 16645
rect 12680 16675 12720 16680
rect 12680 16645 12685 16675
rect 12715 16645 12720 16675
rect 12680 16640 12720 16645
rect 12760 16675 12800 16680
rect 12760 16645 12765 16675
rect 12795 16645 12800 16675
rect 12760 16640 12800 16645
rect 12840 16675 12880 16680
rect 12840 16645 12845 16675
rect 12875 16645 12880 16675
rect 12840 16640 12880 16645
rect 12920 16675 12960 16680
rect 12920 16645 12925 16675
rect 12955 16645 12960 16675
rect 12920 16640 12960 16645
rect 13000 16675 13040 16680
rect 13000 16645 13005 16675
rect 13035 16645 13040 16675
rect 13000 16640 13040 16645
rect 13080 16675 13120 16680
rect 13080 16645 13085 16675
rect 13115 16645 13120 16675
rect 13080 16640 13120 16645
rect 13160 16675 13200 16680
rect 13160 16645 13165 16675
rect 13195 16645 13200 16675
rect 13160 16640 13200 16645
rect 13240 16675 13280 16680
rect 13240 16645 13245 16675
rect 13275 16645 13280 16675
rect 13240 16640 13280 16645
rect 13320 16675 13360 16680
rect 13320 16645 13325 16675
rect 13355 16645 13360 16675
rect 13320 16640 13360 16645
rect 13400 16675 13440 16680
rect 13400 16645 13405 16675
rect 13435 16645 13440 16675
rect 13400 16640 13440 16645
rect 13480 16675 13520 16680
rect 13480 16645 13485 16675
rect 13515 16645 13520 16675
rect 13480 16640 13520 16645
rect 13560 16675 13600 16680
rect 13560 16645 13565 16675
rect 13595 16645 13600 16675
rect 13560 16640 13600 16645
rect 13640 16675 13680 16680
rect 13640 16645 13645 16675
rect 13675 16645 13680 16675
rect 13640 16640 13680 16645
rect 13720 16675 13760 16680
rect 13720 16645 13725 16675
rect 13755 16645 13760 16675
rect 13720 16640 13760 16645
rect 13800 16675 13840 16680
rect 13800 16645 13805 16675
rect 13835 16645 13840 16675
rect 13800 16640 13840 16645
rect 13880 16675 13920 16680
rect 13880 16645 13885 16675
rect 13915 16645 13920 16675
rect 13880 16640 13920 16645
rect 13960 16675 14000 16680
rect 13960 16645 13965 16675
rect 13995 16645 14000 16675
rect 13960 16640 14000 16645
rect 14040 16675 14080 16680
rect 14040 16645 14045 16675
rect 14075 16645 14080 16675
rect 14040 16640 14080 16645
rect 14120 16675 14160 16680
rect 14120 16645 14125 16675
rect 14155 16645 14160 16675
rect 14120 16640 14160 16645
rect 14200 16675 14240 16680
rect 14200 16645 14205 16675
rect 14235 16645 14240 16675
rect 14200 16640 14240 16645
rect 14280 16675 14320 16680
rect 14280 16645 14285 16675
rect 14315 16645 14320 16675
rect 14280 16640 14320 16645
rect 14360 16675 14400 16680
rect 14360 16645 14365 16675
rect 14395 16645 14400 16675
rect 14360 16640 14400 16645
rect 14440 16675 14480 16680
rect 14440 16645 14445 16675
rect 14475 16645 14480 16675
rect 14440 16640 14480 16645
rect 14520 16675 14560 16680
rect 14520 16645 14525 16675
rect 14555 16645 14560 16675
rect 14520 16640 14560 16645
rect 14600 16675 14640 16680
rect 14600 16645 14605 16675
rect 14635 16645 14640 16675
rect 14600 16640 14640 16645
rect 14680 16675 14720 16680
rect 14680 16645 14685 16675
rect 14715 16645 14720 16675
rect 14680 16640 14720 16645
rect 16760 16675 16800 16680
rect 16760 16645 16765 16675
rect 16795 16645 16800 16675
rect 16760 16640 16800 16645
rect 16840 16675 16880 16680
rect 16840 16645 16845 16675
rect 16875 16645 16880 16675
rect 16840 16640 16880 16645
rect 16920 16675 16960 16680
rect 16920 16645 16925 16675
rect 16955 16645 16960 16675
rect 16920 16640 16960 16645
rect 17000 16675 17040 16680
rect 17000 16645 17005 16675
rect 17035 16645 17040 16675
rect 17000 16640 17040 16645
rect 17080 16675 17120 16680
rect 17080 16645 17085 16675
rect 17115 16645 17120 16675
rect 17080 16640 17120 16645
rect 17160 16675 17200 16680
rect 17160 16645 17165 16675
rect 17195 16645 17200 16675
rect 17160 16640 17200 16645
rect 17240 16675 17280 16680
rect 17240 16645 17245 16675
rect 17275 16645 17280 16675
rect 17240 16640 17280 16645
rect 17320 16675 17360 16680
rect 17320 16645 17325 16675
rect 17355 16645 17360 16675
rect 17320 16640 17360 16645
rect 17400 16675 17440 16680
rect 17400 16645 17405 16675
rect 17435 16645 17440 16675
rect 17400 16640 17440 16645
rect 17480 16675 17520 16680
rect 17480 16645 17485 16675
rect 17515 16645 17520 16675
rect 17480 16640 17520 16645
rect 17560 16675 17600 16680
rect 17560 16645 17565 16675
rect 17595 16645 17600 16675
rect 17560 16640 17600 16645
rect 17640 16675 17680 16680
rect 17640 16645 17645 16675
rect 17675 16645 17680 16675
rect 17640 16640 17680 16645
rect 17720 16675 17760 16680
rect 17720 16645 17725 16675
rect 17755 16645 17760 16675
rect 17720 16640 17760 16645
rect 17800 16675 17840 16680
rect 17800 16645 17805 16675
rect 17835 16645 17840 16675
rect 17800 16640 17840 16645
rect 17880 16675 17920 16680
rect 17880 16645 17885 16675
rect 17915 16645 17920 16675
rect 17880 16640 17920 16645
rect 17960 16675 18000 16680
rect 17960 16645 17965 16675
rect 17995 16645 18000 16675
rect 17960 16640 18000 16645
rect 18040 16675 18080 16680
rect 18040 16645 18045 16675
rect 18075 16645 18080 16675
rect 18040 16640 18080 16645
rect 18120 16675 18160 16680
rect 18120 16645 18125 16675
rect 18155 16645 18160 16675
rect 18120 16640 18160 16645
rect 18200 16675 18240 16680
rect 18200 16645 18205 16675
rect 18235 16645 18240 16675
rect 18200 16640 18240 16645
rect 18280 16675 18320 16680
rect 18280 16645 18285 16675
rect 18315 16645 18320 16675
rect 18280 16640 18320 16645
rect 18360 16675 18400 16680
rect 18360 16645 18365 16675
rect 18395 16645 18400 16675
rect 18360 16640 18400 16645
rect 18440 16675 18480 16680
rect 18440 16645 18445 16675
rect 18475 16645 18480 16675
rect 18440 16640 18480 16645
rect 18520 16675 18560 16680
rect 18520 16645 18525 16675
rect 18555 16645 18560 16675
rect 18520 16640 18560 16645
rect 18600 16675 18640 16680
rect 18600 16645 18605 16675
rect 18635 16645 18640 16675
rect 18600 16640 18640 16645
rect 18680 16675 18720 16680
rect 18680 16645 18685 16675
rect 18715 16645 18720 16675
rect 18680 16640 18720 16645
rect 18760 16675 18800 16680
rect 18760 16645 18765 16675
rect 18795 16645 18800 16675
rect 18760 16640 18800 16645
rect 18840 16675 18880 16680
rect 18840 16645 18845 16675
rect 18875 16645 18880 16675
rect 18840 16640 18880 16645
rect 18920 16675 18960 16680
rect 18920 16645 18925 16675
rect 18955 16645 18960 16675
rect 18920 16640 18960 16645
rect 19000 16675 19040 16680
rect 19000 16645 19005 16675
rect 19035 16645 19040 16675
rect 19000 16640 19040 16645
rect 19080 16675 19120 16680
rect 19080 16645 19085 16675
rect 19115 16645 19120 16675
rect 19080 16640 19120 16645
rect 19160 16675 19200 16680
rect 19160 16645 19165 16675
rect 19195 16645 19200 16675
rect 19160 16640 19200 16645
rect 19240 16675 19280 16680
rect 19240 16645 19245 16675
rect 19275 16645 19280 16675
rect 19240 16640 19280 16645
rect 19320 16675 19360 16680
rect 19320 16645 19325 16675
rect 19355 16645 19360 16675
rect 19320 16640 19360 16645
rect 19400 16675 19440 16680
rect 19400 16645 19405 16675
rect 19435 16645 19440 16675
rect 19400 16640 19440 16645
rect 19480 16675 19520 16680
rect 19480 16645 19485 16675
rect 19515 16645 19520 16675
rect 19480 16640 19520 16645
rect 19560 16675 19600 16680
rect 19560 16645 19565 16675
rect 19595 16645 19600 16675
rect 19560 16640 19600 16645
rect 19640 16675 19680 16680
rect 19640 16645 19645 16675
rect 19675 16645 19680 16675
rect 19640 16640 19680 16645
rect 19720 16675 19760 16680
rect 19720 16645 19725 16675
rect 19755 16645 19760 16675
rect 19720 16640 19760 16645
rect 19800 16675 19840 16680
rect 19800 16645 19805 16675
rect 19835 16645 19840 16675
rect 19800 16640 19840 16645
rect 19880 16675 19920 16680
rect 19880 16645 19885 16675
rect 19915 16645 19920 16675
rect 19880 16640 19920 16645
rect 19960 16675 20000 16680
rect 19960 16645 19965 16675
rect 19995 16645 20000 16675
rect 19960 16640 20000 16645
rect 20040 16675 20080 16680
rect 20040 16645 20045 16675
rect 20075 16645 20080 16675
rect 20040 16640 20080 16645
rect 20120 16675 20160 16680
rect 20120 16645 20125 16675
rect 20155 16645 20160 16675
rect 20120 16640 20160 16645
rect 20200 16675 20240 16680
rect 20200 16645 20205 16675
rect 20235 16645 20240 16675
rect 20200 16640 20240 16645
rect 20280 16675 20320 16680
rect 20280 16645 20285 16675
rect 20315 16645 20320 16675
rect 20280 16640 20320 16645
rect 20360 16675 20400 16680
rect 20360 16645 20365 16675
rect 20395 16645 20400 16675
rect 20360 16640 20400 16645
rect 20440 16675 20480 16680
rect 20440 16645 20445 16675
rect 20475 16645 20480 16675
rect 20440 16640 20480 16645
rect 20520 16675 20560 16680
rect 20520 16645 20525 16675
rect 20555 16645 20560 16675
rect 20520 16640 20560 16645
rect 20600 16675 20640 16680
rect 20600 16645 20605 16675
rect 20635 16645 20640 16675
rect 20600 16640 20640 16645
rect 20680 16675 20720 16680
rect 20680 16645 20685 16675
rect 20715 16645 20720 16675
rect 20680 16640 20720 16645
rect 20760 16675 20800 16680
rect 20760 16645 20765 16675
rect 20795 16645 20800 16675
rect 20760 16640 20800 16645
rect 20840 16675 20880 16680
rect 20840 16645 20845 16675
rect 20875 16645 20880 16675
rect 20840 16640 20880 16645
rect 20920 16675 20960 16680
rect 20920 16645 20925 16675
rect 20955 16645 20960 16675
rect 20920 16640 20960 16645
rect 0 16515 40 16520
rect 0 16485 5 16515
rect 35 16485 40 16515
rect 0 16480 40 16485
rect 80 16515 120 16520
rect 80 16485 85 16515
rect 115 16485 120 16515
rect 80 16480 120 16485
rect 160 16515 200 16520
rect 160 16485 165 16515
rect 195 16485 200 16515
rect 160 16480 200 16485
rect 240 16515 280 16520
rect 240 16485 245 16515
rect 275 16485 280 16515
rect 240 16480 280 16485
rect 320 16515 360 16520
rect 320 16485 325 16515
rect 355 16485 360 16515
rect 320 16480 360 16485
rect 400 16515 440 16520
rect 400 16485 405 16515
rect 435 16485 440 16515
rect 400 16480 440 16485
rect 480 16515 520 16520
rect 480 16485 485 16515
rect 515 16485 520 16515
rect 480 16480 520 16485
rect 560 16515 600 16520
rect 560 16485 565 16515
rect 595 16485 600 16515
rect 560 16480 600 16485
rect 640 16515 680 16520
rect 640 16485 645 16515
rect 675 16485 680 16515
rect 640 16480 680 16485
rect 720 16515 760 16520
rect 720 16485 725 16515
rect 755 16485 760 16515
rect 720 16480 760 16485
rect 800 16515 840 16520
rect 800 16485 805 16515
rect 835 16485 840 16515
rect 800 16480 840 16485
rect 880 16515 920 16520
rect 880 16485 885 16515
rect 915 16485 920 16515
rect 880 16480 920 16485
rect 960 16515 1000 16520
rect 960 16485 965 16515
rect 995 16485 1000 16515
rect 960 16480 1000 16485
rect 1040 16515 1080 16520
rect 1040 16485 1045 16515
rect 1075 16485 1080 16515
rect 1040 16480 1080 16485
rect 1120 16515 1160 16520
rect 1120 16485 1125 16515
rect 1155 16485 1160 16515
rect 1120 16480 1160 16485
rect 1200 16515 1240 16520
rect 1200 16485 1205 16515
rect 1235 16485 1240 16515
rect 1200 16480 1240 16485
rect 1280 16515 1320 16520
rect 1280 16485 1285 16515
rect 1315 16485 1320 16515
rect 1280 16480 1320 16485
rect 1360 16515 1400 16520
rect 1360 16485 1365 16515
rect 1395 16485 1400 16515
rect 1360 16480 1400 16485
rect 1440 16515 1480 16520
rect 1440 16485 1445 16515
rect 1475 16485 1480 16515
rect 1440 16480 1480 16485
rect 1520 16515 1560 16520
rect 1520 16485 1525 16515
rect 1555 16485 1560 16515
rect 1520 16480 1560 16485
rect 1600 16515 1640 16520
rect 1600 16485 1605 16515
rect 1635 16485 1640 16515
rect 1600 16480 1640 16485
rect 1680 16515 1720 16520
rect 1680 16485 1685 16515
rect 1715 16485 1720 16515
rect 1680 16480 1720 16485
rect 1760 16515 1800 16520
rect 1760 16485 1765 16515
rect 1795 16485 1800 16515
rect 1760 16480 1800 16485
rect 1840 16515 1880 16520
rect 1840 16485 1845 16515
rect 1875 16485 1880 16515
rect 1840 16480 1880 16485
rect 1920 16515 1960 16520
rect 1920 16485 1925 16515
rect 1955 16485 1960 16515
rect 1920 16480 1960 16485
rect 2000 16515 2040 16520
rect 2000 16485 2005 16515
rect 2035 16485 2040 16515
rect 2000 16480 2040 16485
rect 2080 16515 2120 16520
rect 2080 16485 2085 16515
rect 2115 16485 2120 16515
rect 2080 16480 2120 16485
rect 2160 16515 2200 16520
rect 2160 16485 2165 16515
rect 2195 16485 2200 16515
rect 2160 16480 2200 16485
rect 2240 16515 2280 16520
rect 2240 16485 2245 16515
rect 2275 16485 2280 16515
rect 2240 16480 2280 16485
rect 2320 16515 2360 16520
rect 2320 16485 2325 16515
rect 2355 16485 2360 16515
rect 2320 16480 2360 16485
rect 2400 16515 2440 16520
rect 2400 16485 2405 16515
rect 2435 16485 2440 16515
rect 2400 16480 2440 16485
rect 2480 16515 2520 16520
rect 2480 16485 2485 16515
rect 2515 16485 2520 16515
rect 2480 16480 2520 16485
rect 2560 16515 2600 16520
rect 2560 16485 2565 16515
rect 2595 16485 2600 16515
rect 2560 16480 2600 16485
rect 2640 16515 2680 16520
rect 2640 16485 2645 16515
rect 2675 16485 2680 16515
rect 2640 16480 2680 16485
rect 2720 16515 2760 16520
rect 2720 16485 2725 16515
rect 2755 16485 2760 16515
rect 2720 16480 2760 16485
rect 2800 16515 2840 16520
rect 2800 16485 2805 16515
rect 2835 16485 2840 16515
rect 2800 16480 2840 16485
rect 2880 16515 2920 16520
rect 2880 16485 2885 16515
rect 2915 16485 2920 16515
rect 2880 16480 2920 16485
rect 2960 16515 3000 16520
rect 2960 16485 2965 16515
rect 2995 16485 3000 16515
rect 2960 16480 3000 16485
rect 3040 16515 3080 16520
rect 3040 16485 3045 16515
rect 3075 16485 3080 16515
rect 3040 16480 3080 16485
rect 3120 16515 3160 16520
rect 3120 16485 3125 16515
rect 3155 16485 3160 16515
rect 3120 16480 3160 16485
rect 3200 16515 3240 16520
rect 3200 16485 3205 16515
rect 3235 16485 3240 16515
rect 3200 16480 3240 16485
rect 3280 16515 3320 16520
rect 3280 16485 3285 16515
rect 3315 16485 3320 16515
rect 3280 16480 3320 16485
rect 3360 16515 3400 16520
rect 3360 16485 3365 16515
rect 3395 16485 3400 16515
rect 3360 16480 3400 16485
rect 3440 16515 3480 16520
rect 3440 16485 3445 16515
rect 3475 16485 3480 16515
rect 3440 16480 3480 16485
rect 3520 16515 3560 16520
rect 3520 16485 3525 16515
rect 3555 16485 3560 16515
rect 3520 16480 3560 16485
rect 3600 16515 3640 16520
rect 3600 16485 3605 16515
rect 3635 16485 3640 16515
rect 3600 16480 3640 16485
rect 3680 16515 3720 16520
rect 3680 16485 3685 16515
rect 3715 16485 3720 16515
rect 3680 16480 3720 16485
rect 3760 16515 3800 16520
rect 3760 16485 3765 16515
rect 3795 16485 3800 16515
rect 3760 16480 3800 16485
rect 3840 16515 3880 16520
rect 3840 16485 3845 16515
rect 3875 16485 3880 16515
rect 3840 16480 3880 16485
rect 3920 16515 3960 16520
rect 3920 16485 3925 16515
rect 3955 16485 3960 16515
rect 3920 16480 3960 16485
rect 4000 16515 4040 16520
rect 4000 16485 4005 16515
rect 4035 16485 4040 16515
rect 4000 16480 4040 16485
rect 4080 16515 4120 16520
rect 4080 16485 4085 16515
rect 4115 16485 4120 16515
rect 4080 16480 4120 16485
rect 4160 16515 4200 16520
rect 4160 16485 4165 16515
rect 4195 16485 4200 16515
rect 4160 16480 4200 16485
rect 6240 16515 6280 16520
rect 6240 16485 6245 16515
rect 6275 16485 6280 16515
rect 6240 16480 6280 16485
rect 6320 16515 6360 16520
rect 6320 16485 6325 16515
rect 6355 16485 6360 16515
rect 6320 16480 6360 16485
rect 6400 16515 6440 16520
rect 6400 16485 6405 16515
rect 6435 16485 6440 16515
rect 6400 16480 6440 16485
rect 6480 16515 6520 16520
rect 6480 16485 6485 16515
rect 6515 16485 6520 16515
rect 6480 16480 6520 16485
rect 6560 16515 6600 16520
rect 6560 16485 6565 16515
rect 6595 16485 6600 16515
rect 6560 16480 6600 16485
rect 6640 16515 6680 16520
rect 6640 16485 6645 16515
rect 6675 16485 6680 16515
rect 6640 16480 6680 16485
rect 6720 16515 6760 16520
rect 6720 16485 6725 16515
rect 6755 16485 6760 16515
rect 6720 16480 6760 16485
rect 6800 16515 6840 16520
rect 6800 16485 6805 16515
rect 6835 16485 6840 16515
rect 6800 16480 6840 16485
rect 6880 16515 6920 16520
rect 6880 16485 6885 16515
rect 6915 16485 6920 16515
rect 6880 16480 6920 16485
rect 6960 16515 7000 16520
rect 6960 16485 6965 16515
rect 6995 16485 7000 16515
rect 6960 16480 7000 16485
rect 7040 16515 7080 16520
rect 7040 16485 7045 16515
rect 7075 16485 7080 16515
rect 7040 16480 7080 16485
rect 7120 16515 7160 16520
rect 7120 16485 7125 16515
rect 7155 16485 7160 16515
rect 7120 16480 7160 16485
rect 7200 16515 7240 16520
rect 7200 16485 7205 16515
rect 7235 16485 7240 16515
rect 7200 16480 7240 16485
rect 7280 16515 7320 16520
rect 7280 16485 7285 16515
rect 7315 16485 7320 16515
rect 7280 16480 7320 16485
rect 7360 16515 7400 16520
rect 7360 16485 7365 16515
rect 7395 16485 7400 16515
rect 7360 16480 7400 16485
rect 7440 16515 7480 16520
rect 7440 16485 7445 16515
rect 7475 16485 7480 16515
rect 7440 16480 7480 16485
rect 7520 16515 7560 16520
rect 7520 16485 7525 16515
rect 7555 16485 7560 16515
rect 7520 16480 7560 16485
rect 7600 16515 7640 16520
rect 7600 16485 7605 16515
rect 7635 16485 7640 16515
rect 7600 16480 7640 16485
rect 7680 16515 7720 16520
rect 7680 16485 7685 16515
rect 7715 16485 7720 16515
rect 7680 16480 7720 16485
rect 7760 16515 7800 16520
rect 7760 16485 7765 16515
rect 7795 16485 7800 16515
rect 7760 16480 7800 16485
rect 7840 16515 7880 16520
rect 7840 16485 7845 16515
rect 7875 16485 7880 16515
rect 7840 16480 7880 16485
rect 7920 16515 7960 16520
rect 7920 16485 7925 16515
rect 7955 16485 7960 16515
rect 7920 16480 7960 16485
rect 8000 16515 8040 16520
rect 8000 16485 8005 16515
rect 8035 16485 8040 16515
rect 8000 16480 8040 16485
rect 8080 16515 8120 16520
rect 8080 16485 8085 16515
rect 8115 16485 8120 16515
rect 8080 16480 8120 16485
rect 8160 16515 8200 16520
rect 8160 16485 8165 16515
rect 8195 16485 8200 16515
rect 8160 16480 8200 16485
rect 8240 16515 8280 16520
rect 8240 16485 8245 16515
rect 8275 16485 8280 16515
rect 8240 16480 8280 16485
rect 8320 16515 8360 16520
rect 8320 16485 8325 16515
rect 8355 16485 8360 16515
rect 8320 16480 8360 16485
rect 8400 16515 8440 16520
rect 8400 16485 8405 16515
rect 8435 16485 8440 16515
rect 8400 16480 8440 16485
rect 8480 16515 8520 16520
rect 8480 16485 8485 16515
rect 8515 16485 8520 16515
rect 8480 16480 8520 16485
rect 8560 16515 8600 16520
rect 8560 16485 8565 16515
rect 8595 16485 8600 16515
rect 8560 16480 8600 16485
rect 8640 16515 8680 16520
rect 8640 16485 8645 16515
rect 8675 16485 8680 16515
rect 8640 16480 8680 16485
rect 8720 16515 8760 16520
rect 8720 16485 8725 16515
rect 8755 16485 8760 16515
rect 8720 16480 8760 16485
rect 8800 16515 8840 16520
rect 8800 16485 8805 16515
rect 8835 16485 8840 16515
rect 8800 16480 8840 16485
rect 8880 16515 8920 16520
rect 8880 16485 8885 16515
rect 8915 16485 8920 16515
rect 8880 16480 8920 16485
rect 8960 16515 9000 16520
rect 8960 16485 8965 16515
rect 8995 16485 9000 16515
rect 8960 16480 9000 16485
rect 9040 16515 9080 16520
rect 9040 16485 9045 16515
rect 9075 16485 9080 16515
rect 9040 16480 9080 16485
rect 9120 16515 9160 16520
rect 9120 16485 9125 16515
rect 9155 16485 9160 16515
rect 9120 16480 9160 16485
rect 9200 16515 9240 16520
rect 9200 16485 9205 16515
rect 9235 16485 9240 16515
rect 9200 16480 9240 16485
rect 9280 16515 9320 16520
rect 9280 16485 9285 16515
rect 9315 16485 9320 16515
rect 9280 16480 9320 16485
rect 9360 16515 9400 16520
rect 9360 16485 9365 16515
rect 9395 16485 9400 16515
rect 9360 16480 9400 16485
rect 9440 16515 9480 16520
rect 9440 16485 9445 16515
rect 9475 16485 9480 16515
rect 9440 16480 9480 16485
rect 11560 16515 11600 16520
rect 11560 16485 11565 16515
rect 11595 16485 11600 16515
rect 11560 16480 11600 16485
rect 11640 16515 11680 16520
rect 11640 16485 11645 16515
rect 11675 16485 11680 16515
rect 11640 16480 11680 16485
rect 11720 16515 11760 16520
rect 11720 16485 11725 16515
rect 11755 16485 11760 16515
rect 11720 16480 11760 16485
rect 11800 16515 11840 16520
rect 11800 16485 11805 16515
rect 11835 16485 11840 16515
rect 11800 16480 11840 16485
rect 11880 16515 11920 16520
rect 11880 16485 11885 16515
rect 11915 16485 11920 16515
rect 11880 16480 11920 16485
rect 11960 16515 12000 16520
rect 11960 16485 11965 16515
rect 11995 16485 12000 16515
rect 11960 16480 12000 16485
rect 12040 16515 12080 16520
rect 12040 16485 12045 16515
rect 12075 16485 12080 16515
rect 12040 16480 12080 16485
rect 12120 16515 12160 16520
rect 12120 16485 12125 16515
rect 12155 16485 12160 16515
rect 12120 16480 12160 16485
rect 12200 16515 12240 16520
rect 12200 16485 12205 16515
rect 12235 16485 12240 16515
rect 12200 16480 12240 16485
rect 12280 16515 12320 16520
rect 12280 16485 12285 16515
rect 12315 16485 12320 16515
rect 12280 16480 12320 16485
rect 12360 16515 12400 16520
rect 12360 16485 12365 16515
rect 12395 16485 12400 16515
rect 12360 16480 12400 16485
rect 12440 16515 12480 16520
rect 12440 16485 12445 16515
rect 12475 16485 12480 16515
rect 12440 16480 12480 16485
rect 12520 16515 12560 16520
rect 12520 16485 12525 16515
rect 12555 16485 12560 16515
rect 12520 16480 12560 16485
rect 12600 16515 12640 16520
rect 12600 16485 12605 16515
rect 12635 16485 12640 16515
rect 12600 16480 12640 16485
rect 12680 16515 12720 16520
rect 12680 16485 12685 16515
rect 12715 16485 12720 16515
rect 12680 16480 12720 16485
rect 12760 16515 12800 16520
rect 12760 16485 12765 16515
rect 12795 16485 12800 16515
rect 12760 16480 12800 16485
rect 12840 16515 12880 16520
rect 12840 16485 12845 16515
rect 12875 16485 12880 16515
rect 12840 16480 12880 16485
rect 12920 16515 12960 16520
rect 12920 16485 12925 16515
rect 12955 16485 12960 16515
rect 12920 16480 12960 16485
rect 13000 16515 13040 16520
rect 13000 16485 13005 16515
rect 13035 16485 13040 16515
rect 13000 16480 13040 16485
rect 13080 16515 13120 16520
rect 13080 16485 13085 16515
rect 13115 16485 13120 16515
rect 13080 16480 13120 16485
rect 13160 16515 13200 16520
rect 13160 16485 13165 16515
rect 13195 16485 13200 16515
rect 13160 16480 13200 16485
rect 13240 16515 13280 16520
rect 13240 16485 13245 16515
rect 13275 16485 13280 16515
rect 13240 16480 13280 16485
rect 13320 16515 13360 16520
rect 13320 16485 13325 16515
rect 13355 16485 13360 16515
rect 13320 16480 13360 16485
rect 13400 16515 13440 16520
rect 13400 16485 13405 16515
rect 13435 16485 13440 16515
rect 13400 16480 13440 16485
rect 13480 16515 13520 16520
rect 13480 16485 13485 16515
rect 13515 16485 13520 16515
rect 13480 16480 13520 16485
rect 13560 16515 13600 16520
rect 13560 16485 13565 16515
rect 13595 16485 13600 16515
rect 13560 16480 13600 16485
rect 13640 16515 13680 16520
rect 13640 16485 13645 16515
rect 13675 16485 13680 16515
rect 13640 16480 13680 16485
rect 13720 16515 13760 16520
rect 13720 16485 13725 16515
rect 13755 16485 13760 16515
rect 13720 16480 13760 16485
rect 13800 16515 13840 16520
rect 13800 16485 13805 16515
rect 13835 16485 13840 16515
rect 13800 16480 13840 16485
rect 13880 16515 13920 16520
rect 13880 16485 13885 16515
rect 13915 16485 13920 16515
rect 13880 16480 13920 16485
rect 13960 16515 14000 16520
rect 13960 16485 13965 16515
rect 13995 16485 14000 16515
rect 13960 16480 14000 16485
rect 14040 16515 14080 16520
rect 14040 16485 14045 16515
rect 14075 16485 14080 16515
rect 14040 16480 14080 16485
rect 14120 16515 14160 16520
rect 14120 16485 14125 16515
rect 14155 16485 14160 16515
rect 14120 16480 14160 16485
rect 14200 16515 14240 16520
rect 14200 16485 14205 16515
rect 14235 16485 14240 16515
rect 14200 16480 14240 16485
rect 14280 16515 14320 16520
rect 14280 16485 14285 16515
rect 14315 16485 14320 16515
rect 14280 16480 14320 16485
rect 14360 16515 14400 16520
rect 14360 16485 14365 16515
rect 14395 16485 14400 16515
rect 14360 16480 14400 16485
rect 14440 16515 14480 16520
rect 14440 16485 14445 16515
rect 14475 16485 14480 16515
rect 14440 16480 14480 16485
rect 14520 16515 14560 16520
rect 14520 16485 14525 16515
rect 14555 16485 14560 16515
rect 14520 16480 14560 16485
rect 14600 16515 14640 16520
rect 14600 16485 14605 16515
rect 14635 16485 14640 16515
rect 14600 16480 14640 16485
rect 14680 16515 14720 16520
rect 14680 16485 14685 16515
rect 14715 16485 14720 16515
rect 14680 16480 14720 16485
rect 16760 16515 16800 16520
rect 16760 16485 16765 16515
rect 16795 16485 16800 16515
rect 16760 16480 16800 16485
rect 16840 16515 16880 16520
rect 16840 16485 16845 16515
rect 16875 16485 16880 16515
rect 16840 16480 16880 16485
rect 16920 16515 16960 16520
rect 16920 16485 16925 16515
rect 16955 16485 16960 16515
rect 16920 16480 16960 16485
rect 17000 16515 17040 16520
rect 17000 16485 17005 16515
rect 17035 16485 17040 16515
rect 17000 16480 17040 16485
rect 17080 16515 17120 16520
rect 17080 16485 17085 16515
rect 17115 16485 17120 16515
rect 17080 16480 17120 16485
rect 17160 16515 17200 16520
rect 17160 16485 17165 16515
rect 17195 16485 17200 16515
rect 17160 16480 17200 16485
rect 17240 16515 17280 16520
rect 17240 16485 17245 16515
rect 17275 16485 17280 16515
rect 17240 16480 17280 16485
rect 17320 16515 17360 16520
rect 17320 16485 17325 16515
rect 17355 16485 17360 16515
rect 17320 16480 17360 16485
rect 17400 16515 17440 16520
rect 17400 16485 17405 16515
rect 17435 16485 17440 16515
rect 17400 16480 17440 16485
rect 17480 16515 17520 16520
rect 17480 16485 17485 16515
rect 17515 16485 17520 16515
rect 17480 16480 17520 16485
rect 17560 16515 17600 16520
rect 17560 16485 17565 16515
rect 17595 16485 17600 16515
rect 17560 16480 17600 16485
rect 17640 16515 17680 16520
rect 17640 16485 17645 16515
rect 17675 16485 17680 16515
rect 17640 16480 17680 16485
rect 17720 16515 17760 16520
rect 17720 16485 17725 16515
rect 17755 16485 17760 16515
rect 17720 16480 17760 16485
rect 17800 16515 17840 16520
rect 17800 16485 17805 16515
rect 17835 16485 17840 16515
rect 17800 16480 17840 16485
rect 17880 16515 17920 16520
rect 17880 16485 17885 16515
rect 17915 16485 17920 16515
rect 17880 16480 17920 16485
rect 17960 16515 18000 16520
rect 17960 16485 17965 16515
rect 17995 16485 18000 16515
rect 17960 16480 18000 16485
rect 18040 16515 18080 16520
rect 18040 16485 18045 16515
rect 18075 16485 18080 16515
rect 18040 16480 18080 16485
rect 18120 16515 18160 16520
rect 18120 16485 18125 16515
rect 18155 16485 18160 16515
rect 18120 16480 18160 16485
rect 18200 16515 18240 16520
rect 18200 16485 18205 16515
rect 18235 16485 18240 16515
rect 18200 16480 18240 16485
rect 18280 16515 18320 16520
rect 18280 16485 18285 16515
rect 18315 16485 18320 16515
rect 18280 16480 18320 16485
rect 18360 16515 18400 16520
rect 18360 16485 18365 16515
rect 18395 16485 18400 16515
rect 18360 16480 18400 16485
rect 18440 16515 18480 16520
rect 18440 16485 18445 16515
rect 18475 16485 18480 16515
rect 18440 16480 18480 16485
rect 18520 16515 18560 16520
rect 18520 16485 18525 16515
rect 18555 16485 18560 16515
rect 18520 16480 18560 16485
rect 18600 16515 18640 16520
rect 18600 16485 18605 16515
rect 18635 16485 18640 16515
rect 18600 16480 18640 16485
rect 18680 16515 18720 16520
rect 18680 16485 18685 16515
rect 18715 16485 18720 16515
rect 18680 16480 18720 16485
rect 18760 16515 18800 16520
rect 18760 16485 18765 16515
rect 18795 16485 18800 16515
rect 18760 16480 18800 16485
rect 18840 16515 18880 16520
rect 18840 16485 18845 16515
rect 18875 16485 18880 16515
rect 18840 16480 18880 16485
rect 18920 16515 18960 16520
rect 18920 16485 18925 16515
rect 18955 16485 18960 16515
rect 18920 16480 18960 16485
rect 19000 16515 19040 16520
rect 19000 16485 19005 16515
rect 19035 16485 19040 16515
rect 19000 16480 19040 16485
rect 19080 16515 19120 16520
rect 19080 16485 19085 16515
rect 19115 16485 19120 16515
rect 19080 16480 19120 16485
rect 19160 16515 19200 16520
rect 19160 16485 19165 16515
rect 19195 16485 19200 16515
rect 19160 16480 19200 16485
rect 19240 16515 19280 16520
rect 19240 16485 19245 16515
rect 19275 16485 19280 16515
rect 19240 16480 19280 16485
rect 19320 16515 19360 16520
rect 19320 16485 19325 16515
rect 19355 16485 19360 16515
rect 19320 16480 19360 16485
rect 19400 16515 19440 16520
rect 19400 16485 19405 16515
rect 19435 16485 19440 16515
rect 19400 16480 19440 16485
rect 19480 16515 19520 16520
rect 19480 16485 19485 16515
rect 19515 16485 19520 16515
rect 19480 16480 19520 16485
rect 19560 16515 19600 16520
rect 19560 16485 19565 16515
rect 19595 16485 19600 16515
rect 19560 16480 19600 16485
rect 19640 16515 19680 16520
rect 19640 16485 19645 16515
rect 19675 16485 19680 16515
rect 19640 16480 19680 16485
rect 19720 16515 19760 16520
rect 19720 16485 19725 16515
rect 19755 16485 19760 16515
rect 19720 16480 19760 16485
rect 19800 16515 19840 16520
rect 19800 16485 19805 16515
rect 19835 16485 19840 16515
rect 19800 16480 19840 16485
rect 19880 16515 19920 16520
rect 19880 16485 19885 16515
rect 19915 16485 19920 16515
rect 19880 16480 19920 16485
rect 19960 16515 20000 16520
rect 19960 16485 19965 16515
rect 19995 16485 20000 16515
rect 19960 16480 20000 16485
rect 20040 16515 20080 16520
rect 20040 16485 20045 16515
rect 20075 16485 20080 16515
rect 20040 16480 20080 16485
rect 20120 16515 20160 16520
rect 20120 16485 20125 16515
rect 20155 16485 20160 16515
rect 20120 16480 20160 16485
rect 20200 16515 20240 16520
rect 20200 16485 20205 16515
rect 20235 16485 20240 16515
rect 20200 16480 20240 16485
rect 20280 16515 20320 16520
rect 20280 16485 20285 16515
rect 20315 16485 20320 16515
rect 20280 16480 20320 16485
rect 20360 16515 20400 16520
rect 20360 16485 20365 16515
rect 20395 16485 20400 16515
rect 20360 16480 20400 16485
rect 20440 16515 20480 16520
rect 20440 16485 20445 16515
rect 20475 16485 20480 16515
rect 20440 16480 20480 16485
rect 20520 16515 20560 16520
rect 20520 16485 20525 16515
rect 20555 16485 20560 16515
rect 20520 16480 20560 16485
rect 20600 16515 20640 16520
rect 20600 16485 20605 16515
rect 20635 16485 20640 16515
rect 20600 16480 20640 16485
rect 20680 16515 20720 16520
rect 20680 16485 20685 16515
rect 20715 16485 20720 16515
rect 20680 16480 20720 16485
rect 20760 16515 20800 16520
rect 20760 16485 20765 16515
rect 20795 16485 20800 16515
rect 20760 16480 20800 16485
rect 20840 16515 20880 16520
rect 20840 16485 20845 16515
rect 20875 16485 20880 16515
rect 20840 16480 20880 16485
rect 20920 16515 20960 16520
rect 20920 16485 20925 16515
rect 20955 16485 20960 16515
rect 20920 16480 20960 16485
rect 0 16435 40 16440
rect 0 16405 5 16435
rect 35 16405 40 16435
rect 0 16400 40 16405
rect 80 16435 120 16440
rect 80 16405 85 16435
rect 115 16405 120 16435
rect 80 16400 120 16405
rect 160 16435 200 16440
rect 160 16405 165 16435
rect 195 16405 200 16435
rect 160 16400 200 16405
rect 240 16435 280 16440
rect 240 16405 245 16435
rect 275 16405 280 16435
rect 240 16400 280 16405
rect 320 16435 360 16440
rect 320 16405 325 16435
rect 355 16405 360 16435
rect 320 16400 360 16405
rect 400 16435 440 16440
rect 400 16405 405 16435
rect 435 16405 440 16435
rect 400 16400 440 16405
rect 480 16435 520 16440
rect 480 16405 485 16435
rect 515 16405 520 16435
rect 480 16400 520 16405
rect 560 16435 600 16440
rect 560 16405 565 16435
rect 595 16405 600 16435
rect 560 16400 600 16405
rect 640 16435 680 16440
rect 640 16405 645 16435
rect 675 16405 680 16435
rect 640 16400 680 16405
rect 720 16435 760 16440
rect 720 16405 725 16435
rect 755 16405 760 16435
rect 720 16400 760 16405
rect 800 16435 840 16440
rect 800 16405 805 16435
rect 835 16405 840 16435
rect 800 16400 840 16405
rect 880 16435 920 16440
rect 880 16405 885 16435
rect 915 16405 920 16435
rect 880 16400 920 16405
rect 960 16435 1000 16440
rect 960 16405 965 16435
rect 995 16405 1000 16435
rect 960 16400 1000 16405
rect 1040 16435 1080 16440
rect 1040 16405 1045 16435
rect 1075 16405 1080 16435
rect 1040 16400 1080 16405
rect 1120 16435 1160 16440
rect 1120 16405 1125 16435
rect 1155 16405 1160 16435
rect 1120 16400 1160 16405
rect 1200 16435 1240 16440
rect 1200 16405 1205 16435
rect 1235 16405 1240 16435
rect 1200 16400 1240 16405
rect 1280 16435 1320 16440
rect 1280 16405 1285 16435
rect 1315 16405 1320 16435
rect 1280 16400 1320 16405
rect 1360 16435 1400 16440
rect 1360 16405 1365 16435
rect 1395 16405 1400 16435
rect 1360 16400 1400 16405
rect 1440 16435 1480 16440
rect 1440 16405 1445 16435
rect 1475 16405 1480 16435
rect 1440 16400 1480 16405
rect 1520 16435 1560 16440
rect 1520 16405 1525 16435
rect 1555 16405 1560 16435
rect 1520 16400 1560 16405
rect 1600 16435 1640 16440
rect 1600 16405 1605 16435
rect 1635 16405 1640 16435
rect 1600 16400 1640 16405
rect 1680 16435 1720 16440
rect 1680 16405 1685 16435
rect 1715 16405 1720 16435
rect 1680 16400 1720 16405
rect 1760 16435 1800 16440
rect 1760 16405 1765 16435
rect 1795 16405 1800 16435
rect 1760 16400 1800 16405
rect 1840 16435 1880 16440
rect 1840 16405 1845 16435
rect 1875 16405 1880 16435
rect 1840 16400 1880 16405
rect 1920 16435 1960 16440
rect 1920 16405 1925 16435
rect 1955 16405 1960 16435
rect 1920 16400 1960 16405
rect 2000 16435 2040 16440
rect 2000 16405 2005 16435
rect 2035 16405 2040 16435
rect 2000 16400 2040 16405
rect 2080 16435 2120 16440
rect 2080 16405 2085 16435
rect 2115 16405 2120 16435
rect 2080 16400 2120 16405
rect 2160 16435 2200 16440
rect 2160 16405 2165 16435
rect 2195 16405 2200 16435
rect 2160 16400 2200 16405
rect 2240 16435 2280 16440
rect 2240 16405 2245 16435
rect 2275 16405 2280 16435
rect 2240 16400 2280 16405
rect 2320 16435 2360 16440
rect 2320 16405 2325 16435
rect 2355 16405 2360 16435
rect 2320 16400 2360 16405
rect 2400 16435 2440 16440
rect 2400 16405 2405 16435
rect 2435 16405 2440 16435
rect 2400 16400 2440 16405
rect 2480 16435 2520 16440
rect 2480 16405 2485 16435
rect 2515 16405 2520 16435
rect 2480 16400 2520 16405
rect 2560 16435 2600 16440
rect 2560 16405 2565 16435
rect 2595 16405 2600 16435
rect 2560 16400 2600 16405
rect 2640 16435 2680 16440
rect 2640 16405 2645 16435
rect 2675 16405 2680 16435
rect 2640 16400 2680 16405
rect 2720 16435 2760 16440
rect 2720 16405 2725 16435
rect 2755 16405 2760 16435
rect 2720 16400 2760 16405
rect 2800 16435 2840 16440
rect 2800 16405 2805 16435
rect 2835 16405 2840 16435
rect 2800 16400 2840 16405
rect 2880 16435 2920 16440
rect 2880 16405 2885 16435
rect 2915 16405 2920 16435
rect 2880 16400 2920 16405
rect 2960 16435 3000 16440
rect 2960 16405 2965 16435
rect 2995 16405 3000 16435
rect 2960 16400 3000 16405
rect 3040 16435 3080 16440
rect 3040 16405 3045 16435
rect 3075 16405 3080 16435
rect 3040 16400 3080 16405
rect 3120 16435 3160 16440
rect 3120 16405 3125 16435
rect 3155 16405 3160 16435
rect 3120 16400 3160 16405
rect 3200 16435 3240 16440
rect 3200 16405 3205 16435
rect 3235 16405 3240 16435
rect 3200 16400 3240 16405
rect 3280 16435 3320 16440
rect 3280 16405 3285 16435
rect 3315 16405 3320 16435
rect 3280 16400 3320 16405
rect 3360 16435 3400 16440
rect 3360 16405 3365 16435
rect 3395 16405 3400 16435
rect 3360 16400 3400 16405
rect 3440 16435 3480 16440
rect 3440 16405 3445 16435
rect 3475 16405 3480 16435
rect 3440 16400 3480 16405
rect 3520 16435 3560 16440
rect 3520 16405 3525 16435
rect 3555 16405 3560 16435
rect 3520 16400 3560 16405
rect 3600 16435 3640 16440
rect 3600 16405 3605 16435
rect 3635 16405 3640 16435
rect 3600 16400 3640 16405
rect 3680 16435 3720 16440
rect 3680 16405 3685 16435
rect 3715 16405 3720 16435
rect 3680 16400 3720 16405
rect 3760 16435 3800 16440
rect 3760 16405 3765 16435
rect 3795 16405 3800 16435
rect 3760 16400 3800 16405
rect 3840 16435 3880 16440
rect 3840 16405 3845 16435
rect 3875 16405 3880 16435
rect 3840 16400 3880 16405
rect 3920 16435 3960 16440
rect 3920 16405 3925 16435
rect 3955 16405 3960 16435
rect 3920 16400 3960 16405
rect 4000 16435 4040 16440
rect 4000 16405 4005 16435
rect 4035 16405 4040 16435
rect 4000 16400 4040 16405
rect 4080 16435 4120 16440
rect 4080 16405 4085 16435
rect 4115 16405 4120 16435
rect 4080 16400 4120 16405
rect 4160 16435 4200 16440
rect 4160 16405 4165 16435
rect 4195 16405 4200 16435
rect 4160 16400 4200 16405
rect 6240 16435 6280 16440
rect 6240 16405 6245 16435
rect 6275 16405 6280 16435
rect 6240 16400 6280 16405
rect 6320 16435 6360 16440
rect 6320 16405 6325 16435
rect 6355 16405 6360 16435
rect 6320 16400 6360 16405
rect 6400 16435 6440 16440
rect 6400 16405 6405 16435
rect 6435 16405 6440 16435
rect 6400 16400 6440 16405
rect 6480 16435 6520 16440
rect 6480 16405 6485 16435
rect 6515 16405 6520 16435
rect 6480 16400 6520 16405
rect 6560 16435 6600 16440
rect 6560 16405 6565 16435
rect 6595 16405 6600 16435
rect 6560 16400 6600 16405
rect 6640 16435 6680 16440
rect 6640 16405 6645 16435
rect 6675 16405 6680 16435
rect 6640 16400 6680 16405
rect 6720 16435 6760 16440
rect 6720 16405 6725 16435
rect 6755 16405 6760 16435
rect 6720 16400 6760 16405
rect 6800 16435 6840 16440
rect 6800 16405 6805 16435
rect 6835 16405 6840 16435
rect 6800 16400 6840 16405
rect 6880 16435 6920 16440
rect 6880 16405 6885 16435
rect 6915 16405 6920 16435
rect 6880 16400 6920 16405
rect 6960 16435 7000 16440
rect 6960 16405 6965 16435
rect 6995 16405 7000 16435
rect 6960 16400 7000 16405
rect 7040 16435 7080 16440
rect 7040 16405 7045 16435
rect 7075 16405 7080 16435
rect 7040 16400 7080 16405
rect 7120 16435 7160 16440
rect 7120 16405 7125 16435
rect 7155 16405 7160 16435
rect 7120 16400 7160 16405
rect 7200 16435 7240 16440
rect 7200 16405 7205 16435
rect 7235 16405 7240 16435
rect 7200 16400 7240 16405
rect 7280 16435 7320 16440
rect 7280 16405 7285 16435
rect 7315 16405 7320 16435
rect 7280 16400 7320 16405
rect 7360 16435 7400 16440
rect 7360 16405 7365 16435
rect 7395 16405 7400 16435
rect 7360 16400 7400 16405
rect 7440 16435 7480 16440
rect 7440 16405 7445 16435
rect 7475 16405 7480 16435
rect 7440 16400 7480 16405
rect 7520 16435 7560 16440
rect 7520 16405 7525 16435
rect 7555 16405 7560 16435
rect 7520 16400 7560 16405
rect 7600 16435 7640 16440
rect 7600 16405 7605 16435
rect 7635 16405 7640 16435
rect 7600 16400 7640 16405
rect 7680 16435 7720 16440
rect 7680 16405 7685 16435
rect 7715 16405 7720 16435
rect 7680 16400 7720 16405
rect 7760 16435 7800 16440
rect 7760 16405 7765 16435
rect 7795 16405 7800 16435
rect 7760 16400 7800 16405
rect 7840 16435 7880 16440
rect 7840 16405 7845 16435
rect 7875 16405 7880 16435
rect 7840 16400 7880 16405
rect 7920 16435 7960 16440
rect 7920 16405 7925 16435
rect 7955 16405 7960 16435
rect 7920 16400 7960 16405
rect 8000 16435 8040 16440
rect 8000 16405 8005 16435
rect 8035 16405 8040 16435
rect 8000 16400 8040 16405
rect 8080 16435 8120 16440
rect 8080 16405 8085 16435
rect 8115 16405 8120 16435
rect 8080 16400 8120 16405
rect 8160 16435 8200 16440
rect 8160 16405 8165 16435
rect 8195 16405 8200 16435
rect 8160 16400 8200 16405
rect 8240 16435 8280 16440
rect 8240 16405 8245 16435
rect 8275 16405 8280 16435
rect 8240 16400 8280 16405
rect 8320 16435 8360 16440
rect 8320 16405 8325 16435
rect 8355 16405 8360 16435
rect 8320 16400 8360 16405
rect 8400 16435 8440 16440
rect 8400 16405 8405 16435
rect 8435 16405 8440 16435
rect 8400 16400 8440 16405
rect 8480 16435 8520 16440
rect 8480 16405 8485 16435
rect 8515 16405 8520 16435
rect 8480 16400 8520 16405
rect 8560 16435 8600 16440
rect 8560 16405 8565 16435
rect 8595 16405 8600 16435
rect 8560 16400 8600 16405
rect 8640 16435 8680 16440
rect 8640 16405 8645 16435
rect 8675 16405 8680 16435
rect 8640 16400 8680 16405
rect 8720 16435 8760 16440
rect 8720 16405 8725 16435
rect 8755 16405 8760 16435
rect 8720 16400 8760 16405
rect 8800 16435 8840 16440
rect 8800 16405 8805 16435
rect 8835 16405 8840 16435
rect 8800 16400 8840 16405
rect 8880 16435 8920 16440
rect 8880 16405 8885 16435
rect 8915 16405 8920 16435
rect 8880 16400 8920 16405
rect 8960 16435 9000 16440
rect 8960 16405 8965 16435
rect 8995 16405 9000 16435
rect 8960 16400 9000 16405
rect 9040 16435 9080 16440
rect 9040 16405 9045 16435
rect 9075 16405 9080 16435
rect 9040 16400 9080 16405
rect 9120 16435 9160 16440
rect 9120 16405 9125 16435
rect 9155 16405 9160 16435
rect 9120 16400 9160 16405
rect 9200 16435 9240 16440
rect 9200 16405 9205 16435
rect 9235 16405 9240 16435
rect 9200 16400 9240 16405
rect 9280 16435 9320 16440
rect 9280 16405 9285 16435
rect 9315 16405 9320 16435
rect 9280 16400 9320 16405
rect 9360 16435 9400 16440
rect 9360 16405 9365 16435
rect 9395 16405 9400 16435
rect 9360 16400 9400 16405
rect 9440 16435 9480 16440
rect 9440 16405 9445 16435
rect 9475 16405 9480 16435
rect 9440 16400 9480 16405
rect 11560 16435 11600 16440
rect 11560 16405 11565 16435
rect 11595 16405 11600 16435
rect 11560 16400 11600 16405
rect 11640 16435 11680 16440
rect 11640 16405 11645 16435
rect 11675 16405 11680 16435
rect 11640 16400 11680 16405
rect 11720 16435 11760 16440
rect 11720 16405 11725 16435
rect 11755 16405 11760 16435
rect 11720 16400 11760 16405
rect 11800 16435 11840 16440
rect 11800 16405 11805 16435
rect 11835 16405 11840 16435
rect 11800 16400 11840 16405
rect 11880 16435 11920 16440
rect 11880 16405 11885 16435
rect 11915 16405 11920 16435
rect 11880 16400 11920 16405
rect 11960 16435 12000 16440
rect 11960 16405 11965 16435
rect 11995 16405 12000 16435
rect 11960 16400 12000 16405
rect 12040 16435 12080 16440
rect 12040 16405 12045 16435
rect 12075 16405 12080 16435
rect 12040 16400 12080 16405
rect 12120 16435 12160 16440
rect 12120 16405 12125 16435
rect 12155 16405 12160 16435
rect 12120 16400 12160 16405
rect 12200 16435 12240 16440
rect 12200 16405 12205 16435
rect 12235 16405 12240 16435
rect 12200 16400 12240 16405
rect 12280 16435 12320 16440
rect 12280 16405 12285 16435
rect 12315 16405 12320 16435
rect 12280 16400 12320 16405
rect 12360 16435 12400 16440
rect 12360 16405 12365 16435
rect 12395 16405 12400 16435
rect 12360 16400 12400 16405
rect 12440 16435 12480 16440
rect 12440 16405 12445 16435
rect 12475 16405 12480 16435
rect 12440 16400 12480 16405
rect 12520 16435 12560 16440
rect 12520 16405 12525 16435
rect 12555 16405 12560 16435
rect 12520 16400 12560 16405
rect 12600 16435 12640 16440
rect 12600 16405 12605 16435
rect 12635 16405 12640 16435
rect 12600 16400 12640 16405
rect 12680 16435 12720 16440
rect 12680 16405 12685 16435
rect 12715 16405 12720 16435
rect 12680 16400 12720 16405
rect 12760 16435 12800 16440
rect 12760 16405 12765 16435
rect 12795 16405 12800 16435
rect 12760 16400 12800 16405
rect 12840 16435 12880 16440
rect 12840 16405 12845 16435
rect 12875 16405 12880 16435
rect 12840 16400 12880 16405
rect 12920 16435 12960 16440
rect 12920 16405 12925 16435
rect 12955 16405 12960 16435
rect 12920 16400 12960 16405
rect 13000 16435 13040 16440
rect 13000 16405 13005 16435
rect 13035 16405 13040 16435
rect 13000 16400 13040 16405
rect 13080 16435 13120 16440
rect 13080 16405 13085 16435
rect 13115 16405 13120 16435
rect 13080 16400 13120 16405
rect 13160 16435 13200 16440
rect 13160 16405 13165 16435
rect 13195 16405 13200 16435
rect 13160 16400 13200 16405
rect 13240 16435 13280 16440
rect 13240 16405 13245 16435
rect 13275 16405 13280 16435
rect 13240 16400 13280 16405
rect 13320 16435 13360 16440
rect 13320 16405 13325 16435
rect 13355 16405 13360 16435
rect 13320 16400 13360 16405
rect 13400 16435 13440 16440
rect 13400 16405 13405 16435
rect 13435 16405 13440 16435
rect 13400 16400 13440 16405
rect 13480 16435 13520 16440
rect 13480 16405 13485 16435
rect 13515 16405 13520 16435
rect 13480 16400 13520 16405
rect 13560 16435 13600 16440
rect 13560 16405 13565 16435
rect 13595 16405 13600 16435
rect 13560 16400 13600 16405
rect 13640 16435 13680 16440
rect 13640 16405 13645 16435
rect 13675 16405 13680 16435
rect 13640 16400 13680 16405
rect 13720 16435 13760 16440
rect 13720 16405 13725 16435
rect 13755 16405 13760 16435
rect 13720 16400 13760 16405
rect 13800 16435 13840 16440
rect 13800 16405 13805 16435
rect 13835 16405 13840 16435
rect 13800 16400 13840 16405
rect 13880 16435 13920 16440
rect 13880 16405 13885 16435
rect 13915 16405 13920 16435
rect 13880 16400 13920 16405
rect 13960 16435 14000 16440
rect 13960 16405 13965 16435
rect 13995 16405 14000 16435
rect 13960 16400 14000 16405
rect 14040 16435 14080 16440
rect 14040 16405 14045 16435
rect 14075 16405 14080 16435
rect 14040 16400 14080 16405
rect 14120 16435 14160 16440
rect 14120 16405 14125 16435
rect 14155 16405 14160 16435
rect 14120 16400 14160 16405
rect 14200 16435 14240 16440
rect 14200 16405 14205 16435
rect 14235 16405 14240 16435
rect 14200 16400 14240 16405
rect 14280 16435 14320 16440
rect 14280 16405 14285 16435
rect 14315 16405 14320 16435
rect 14280 16400 14320 16405
rect 14360 16435 14400 16440
rect 14360 16405 14365 16435
rect 14395 16405 14400 16435
rect 14360 16400 14400 16405
rect 14440 16435 14480 16440
rect 14440 16405 14445 16435
rect 14475 16405 14480 16435
rect 14440 16400 14480 16405
rect 14520 16435 14560 16440
rect 14520 16405 14525 16435
rect 14555 16405 14560 16435
rect 14520 16400 14560 16405
rect 14600 16435 14640 16440
rect 14600 16405 14605 16435
rect 14635 16405 14640 16435
rect 14600 16400 14640 16405
rect 14680 16435 14720 16440
rect 14680 16405 14685 16435
rect 14715 16405 14720 16435
rect 14680 16400 14720 16405
rect 16760 16435 16800 16440
rect 16760 16405 16765 16435
rect 16795 16405 16800 16435
rect 16760 16400 16800 16405
rect 16840 16435 16880 16440
rect 16840 16405 16845 16435
rect 16875 16405 16880 16435
rect 16840 16400 16880 16405
rect 16920 16435 16960 16440
rect 16920 16405 16925 16435
rect 16955 16405 16960 16435
rect 16920 16400 16960 16405
rect 17000 16435 17040 16440
rect 17000 16405 17005 16435
rect 17035 16405 17040 16435
rect 17000 16400 17040 16405
rect 17080 16435 17120 16440
rect 17080 16405 17085 16435
rect 17115 16405 17120 16435
rect 17080 16400 17120 16405
rect 17160 16435 17200 16440
rect 17160 16405 17165 16435
rect 17195 16405 17200 16435
rect 17160 16400 17200 16405
rect 17240 16435 17280 16440
rect 17240 16405 17245 16435
rect 17275 16405 17280 16435
rect 17240 16400 17280 16405
rect 17320 16435 17360 16440
rect 17320 16405 17325 16435
rect 17355 16405 17360 16435
rect 17320 16400 17360 16405
rect 17400 16435 17440 16440
rect 17400 16405 17405 16435
rect 17435 16405 17440 16435
rect 17400 16400 17440 16405
rect 17480 16435 17520 16440
rect 17480 16405 17485 16435
rect 17515 16405 17520 16435
rect 17480 16400 17520 16405
rect 17560 16435 17600 16440
rect 17560 16405 17565 16435
rect 17595 16405 17600 16435
rect 17560 16400 17600 16405
rect 17640 16435 17680 16440
rect 17640 16405 17645 16435
rect 17675 16405 17680 16435
rect 17640 16400 17680 16405
rect 17720 16435 17760 16440
rect 17720 16405 17725 16435
rect 17755 16405 17760 16435
rect 17720 16400 17760 16405
rect 17800 16435 17840 16440
rect 17800 16405 17805 16435
rect 17835 16405 17840 16435
rect 17800 16400 17840 16405
rect 17880 16435 17920 16440
rect 17880 16405 17885 16435
rect 17915 16405 17920 16435
rect 17880 16400 17920 16405
rect 17960 16435 18000 16440
rect 17960 16405 17965 16435
rect 17995 16405 18000 16435
rect 17960 16400 18000 16405
rect 18040 16435 18080 16440
rect 18040 16405 18045 16435
rect 18075 16405 18080 16435
rect 18040 16400 18080 16405
rect 18120 16435 18160 16440
rect 18120 16405 18125 16435
rect 18155 16405 18160 16435
rect 18120 16400 18160 16405
rect 18200 16435 18240 16440
rect 18200 16405 18205 16435
rect 18235 16405 18240 16435
rect 18200 16400 18240 16405
rect 18280 16435 18320 16440
rect 18280 16405 18285 16435
rect 18315 16405 18320 16435
rect 18280 16400 18320 16405
rect 18360 16435 18400 16440
rect 18360 16405 18365 16435
rect 18395 16405 18400 16435
rect 18360 16400 18400 16405
rect 18440 16435 18480 16440
rect 18440 16405 18445 16435
rect 18475 16405 18480 16435
rect 18440 16400 18480 16405
rect 18520 16435 18560 16440
rect 18520 16405 18525 16435
rect 18555 16405 18560 16435
rect 18520 16400 18560 16405
rect 18600 16435 18640 16440
rect 18600 16405 18605 16435
rect 18635 16405 18640 16435
rect 18600 16400 18640 16405
rect 18680 16435 18720 16440
rect 18680 16405 18685 16435
rect 18715 16405 18720 16435
rect 18680 16400 18720 16405
rect 18760 16435 18800 16440
rect 18760 16405 18765 16435
rect 18795 16405 18800 16435
rect 18760 16400 18800 16405
rect 18840 16435 18880 16440
rect 18840 16405 18845 16435
rect 18875 16405 18880 16435
rect 18840 16400 18880 16405
rect 18920 16435 18960 16440
rect 18920 16405 18925 16435
rect 18955 16405 18960 16435
rect 18920 16400 18960 16405
rect 19000 16435 19040 16440
rect 19000 16405 19005 16435
rect 19035 16405 19040 16435
rect 19000 16400 19040 16405
rect 19080 16435 19120 16440
rect 19080 16405 19085 16435
rect 19115 16405 19120 16435
rect 19080 16400 19120 16405
rect 19160 16435 19200 16440
rect 19160 16405 19165 16435
rect 19195 16405 19200 16435
rect 19160 16400 19200 16405
rect 19240 16435 19280 16440
rect 19240 16405 19245 16435
rect 19275 16405 19280 16435
rect 19240 16400 19280 16405
rect 19320 16435 19360 16440
rect 19320 16405 19325 16435
rect 19355 16405 19360 16435
rect 19320 16400 19360 16405
rect 19400 16435 19440 16440
rect 19400 16405 19405 16435
rect 19435 16405 19440 16435
rect 19400 16400 19440 16405
rect 19480 16435 19520 16440
rect 19480 16405 19485 16435
rect 19515 16405 19520 16435
rect 19480 16400 19520 16405
rect 19560 16435 19600 16440
rect 19560 16405 19565 16435
rect 19595 16405 19600 16435
rect 19560 16400 19600 16405
rect 19640 16435 19680 16440
rect 19640 16405 19645 16435
rect 19675 16405 19680 16435
rect 19640 16400 19680 16405
rect 19720 16435 19760 16440
rect 19720 16405 19725 16435
rect 19755 16405 19760 16435
rect 19720 16400 19760 16405
rect 19800 16435 19840 16440
rect 19800 16405 19805 16435
rect 19835 16405 19840 16435
rect 19800 16400 19840 16405
rect 19880 16435 19920 16440
rect 19880 16405 19885 16435
rect 19915 16405 19920 16435
rect 19880 16400 19920 16405
rect 19960 16435 20000 16440
rect 19960 16405 19965 16435
rect 19995 16405 20000 16435
rect 19960 16400 20000 16405
rect 20040 16435 20080 16440
rect 20040 16405 20045 16435
rect 20075 16405 20080 16435
rect 20040 16400 20080 16405
rect 20120 16435 20160 16440
rect 20120 16405 20125 16435
rect 20155 16405 20160 16435
rect 20120 16400 20160 16405
rect 20200 16435 20240 16440
rect 20200 16405 20205 16435
rect 20235 16405 20240 16435
rect 20200 16400 20240 16405
rect 20280 16435 20320 16440
rect 20280 16405 20285 16435
rect 20315 16405 20320 16435
rect 20280 16400 20320 16405
rect 20360 16435 20400 16440
rect 20360 16405 20365 16435
rect 20395 16405 20400 16435
rect 20360 16400 20400 16405
rect 20440 16435 20480 16440
rect 20440 16405 20445 16435
rect 20475 16405 20480 16435
rect 20440 16400 20480 16405
rect 20520 16435 20560 16440
rect 20520 16405 20525 16435
rect 20555 16405 20560 16435
rect 20520 16400 20560 16405
rect 20600 16435 20640 16440
rect 20600 16405 20605 16435
rect 20635 16405 20640 16435
rect 20600 16400 20640 16405
rect 20680 16435 20720 16440
rect 20680 16405 20685 16435
rect 20715 16405 20720 16435
rect 20680 16400 20720 16405
rect 20760 16435 20800 16440
rect 20760 16405 20765 16435
rect 20795 16405 20800 16435
rect 20760 16400 20800 16405
rect 20840 16435 20880 16440
rect 20840 16405 20845 16435
rect 20875 16405 20880 16435
rect 20840 16400 20880 16405
rect 20920 16435 20960 16440
rect 20920 16405 20925 16435
rect 20955 16405 20960 16435
rect 20920 16400 20960 16405
rect 0 16275 40 16280
rect 0 16245 5 16275
rect 35 16245 40 16275
rect 0 16240 40 16245
rect 80 16275 120 16280
rect 80 16245 85 16275
rect 115 16245 120 16275
rect 80 16240 120 16245
rect 160 16275 200 16280
rect 160 16245 165 16275
rect 195 16245 200 16275
rect 160 16240 200 16245
rect 240 16275 280 16280
rect 240 16245 245 16275
rect 275 16245 280 16275
rect 240 16240 280 16245
rect 320 16275 360 16280
rect 320 16245 325 16275
rect 355 16245 360 16275
rect 320 16240 360 16245
rect 400 16275 440 16280
rect 400 16245 405 16275
rect 435 16245 440 16275
rect 400 16240 440 16245
rect 480 16275 520 16280
rect 480 16245 485 16275
rect 515 16245 520 16275
rect 480 16240 520 16245
rect 560 16275 600 16280
rect 560 16245 565 16275
rect 595 16245 600 16275
rect 560 16240 600 16245
rect 640 16275 680 16280
rect 640 16245 645 16275
rect 675 16245 680 16275
rect 640 16240 680 16245
rect 720 16275 760 16280
rect 720 16245 725 16275
rect 755 16245 760 16275
rect 720 16240 760 16245
rect 800 16275 840 16280
rect 800 16245 805 16275
rect 835 16245 840 16275
rect 800 16240 840 16245
rect 880 16275 920 16280
rect 880 16245 885 16275
rect 915 16245 920 16275
rect 880 16240 920 16245
rect 960 16275 1000 16280
rect 960 16245 965 16275
rect 995 16245 1000 16275
rect 960 16240 1000 16245
rect 1040 16275 1080 16280
rect 1040 16245 1045 16275
rect 1075 16245 1080 16275
rect 1040 16240 1080 16245
rect 1120 16275 1160 16280
rect 1120 16245 1125 16275
rect 1155 16245 1160 16275
rect 1120 16240 1160 16245
rect 1200 16275 1240 16280
rect 1200 16245 1205 16275
rect 1235 16245 1240 16275
rect 1200 16240 1240 16245
rect 1280 16275 1320 16280
rect 1280 16245 1285 16275
rect 1315 16245 1320 16275
rect 1280 16240 1320 16245
rect 1360 16275 1400 16280
rect 1360 16245 1365 16275
rect 1395 16245 1400 16275
rect 1360 16240 1400 16245
rect 1440 16275 1480 16280
rect 1440 16245 1445 16275
rect 1475 16245 1480 16275
rect 1440 16240 1480 16245
rect 1520 16275 1560 16280
rect 1520 16245 1525 16275
rect 1555 16245 1560 16275
rect 1520 16240 1560 16245
rect 1600 16275 1640 16280
rect 1600 16245 1605 16275
rect 1635 16245 1640 16275
rect 1600 16240 1640 16245
rect 1680 16275 1720 16280
rect 1680 16245 1685 16275
rect 1715 16245 1720 16275
rect 1680 16240 1720 16245
rect 1760 16275 1800 16280
rect 1760 16245 1765 16275
rect 1795 16245 1800 16275
rect 1760 16240 1800 16245
rect 1840 16275 1880 16280
rect 1840 16245 1845 16275
rect 1875 16245 1880 16275
rect 1840 16240 1880 16245
rect 1920 16275 1960 16280
rect 1920 16245 1925 16275
rect 1955 16245 1960 16275
rect 1920 16240 1960 16245
rect 2000 16275 2040 16280
rect 2000 16245 2005 16275
rect 2035 16245 2040 16275
rect 2000 16240 2040 16245
rect 2080 16275 2120 16280
rect 2080 16245 2085 16275
rect 2115 16245 2120 16275
rect 2080 16240 2120 16245
rect 2160 16275 2200 16280
rect 2160 16245 2165 16275
rect 2195 16245 2200 16275
rect 2160 16240 2200 16245
rect 2240 16275 2280 16280
rect 2240 16245 2245 16275
rect 2275 16245 2280 16275
rect 2240 16240 2280 16245
rect 2320 16275 2360 16280
rect 2320 16245 2325 16275
rect 2355 16245 2360 16275
rect 2320 16240 2360 16245
rect 2400 16275 2440 16280
rect 2400 16245 2405 16275
rect 2435 16245 2440 16275
rect 2400 16240 2440 16245
rect 2480 16275 2520 16280
rect 2480 16245 2485 16275
rect 2515 16245 2520 16275
rect 2480 16240 2520 16245
rect 2560 16275 2600 16280
rect 2560 16245 2565 16275
rect 2595 16245 2600 16275
rect 2560 16240 2600 16245
rect 2640 16275 2680 16280
rect 2640 16245 2645 16275
rect 2675 16245 2680 16275
rect 2640 16240 2680 16245
rect 2720 16275 2760 16280
rect 2720 16245 2725 16275
rect 2755 16245 2760 16275
rect 2720 16240 2760 16245
rect 2800 16275 2840 16280
rect 2800 16245 2805 16275
rect 2835 16245 2840 16275
rect 2800 16240 2840 16245
rect 2880 16275 2920 16280
rect 2880 16245 2885 16275
rect 2915 16245 2920 16275
rect 2880 16240 2920 16245
rect 2960 16275 3000 16280
rect 2960 16245 2965 16275
rect 2995 16245 3000 16275
rect 2960 16240 3000 16245
rect 3040 16275 3080 16280
rect 3040 16245 3045 16275
rect 3075 16245 3080 16275
rect 3040 16240 3080 16245
rect 3120 16275 3160 16280
rect 3120 16245 3125 16275
rect 3155 16245 3160 16275
rect 3120 16240 3160 16245
rect 3200 16275 3240 16280
rect 3200 16245 3205 16275
rect 3235 16245 3240 16275
rect 3200 16240 3240 16245
rect 3280 16275 3320 16280
rect 3280 16245 3285 16275
rect 3315 16245 3320 16275
rect 3280 16240 3320 16245
rect 3360 16275 3400 16280
rect 3360 16245 3365 16275
rect 3395 16245 3400 16275
rect 3360 16240 3400 16245
rect 3440 16275 3480 16280
rect 3440 16245 3445 16275
rect 3475 16245 3480 16275
rect 3440 16240 3480 16245
rect 3520 16275 3560 16280
rect 3520 16245 3525 16275
rect 3555 16245 3560 16275
rect 3520 16240 3560 16245
rect 3600 16275 3640 16280
rect 3600 16245 3605 16275
rect 3635 16245 3640 16275
rect 3600 16240 3640 16245
rect 3680 16275 3720 16280
rect 3680 16245 3685 16275
rect 3715 16245 3720 16275
rect 3680 16240 3720 16245
rect 3760 16275 3800 16280
rect 3760 16245 3765 16275
rect 3795 16245 3800 16275
rect 3760 16240 3800 16245
rect 3840 16275 3880 16280
rect 3840 16245 3845 16275
rect 3875 16245 3880 16275
rect 3840 16240 3880 16245
rect 3920 16275 3960 16280
rect 3920 16245 3925 16275
rect 3955 16245 3960 16275
rect 3920 16240 3960 16245
rect 4000 16275 4040 16280
rect 4000 16245 4005 16275
rect 4035 16245 4040 16275
rect 4000 16240 4040 16245
rect 4080 16275 4120 16280
rect 4080 16245 4085 16275
rect 4115 16245 4120 16275
rect 4080 16240 4120 16245
rect 4160 16275 4200 16280
rect 4160 16245 4165 16275
rect 4195 16245 4200 16275
rect 4160 16240 4200 16245
rect 6240 16275 6280 16280
rect 6240 16245 6245 16275
rect 6275 16245 6280 16275
rect 6240 16240 6280 16245
rect 6320 16275 6360 16280
rect 6320 16245 6325 16275
rect 6355 16245 6360 16275
rect 6320 16240 6360 16245
rect 6400 16275 6440 16280
rect 6400 16245 6405 16275
rect 6435 16245 6440 16275
rect 6400 16240 6440 16245
rect 6480 16275 6520 16280
rect 6480 16245 6485 16275
rect 6515 16245 6520 16275
rect 6480 16240 6520 16245
rect 6560 16275 6600 16280
rect 6560 16245 6565 16275
rect 6595 16245 6600 16275
rect 6560 16240 6600 16245
rect 6640 16275 6680 16280
rect 6640 16245 6645 16275
rect 6675 16245 6680 16275
rect 6640 16240 6680 16245
rect 6720 16275 6760 16280
rect 6720 16245 6725 16275
rect 6755 16245 6760 16275
rect 6720 16240 6760 16245
rect 6800 16275 6840 16280
rect 6800 16245 6805 16275
rect 6835 16245 6840 16275
rect 6800 16240 6840 16245
rect 6880 16275 6920 16280
rect 6880 16245 6885 16275
rect 6915 16245 6920 16275
rect 6880 16240 6920 16245
rect 6960 16275 7000 16280
rect 6960 16245 6965 16275
rect 6995 16245 7000 16275
rect 6960 16240 7000 16245
rect 7040 16275 7080 16280
rect 7040 16245 7045 16275
rect 7075 16245 7080 16275
rect 7040 16240 7080 16245
rect 7120 16275 7160 16280
rect 7120 16245 7125 16275
rect 7155 16245 7160 16275
rect 7120 16240 7160 16245
rect 7200 16275 7240 16280
rect 7200 16245 7205 16275
rect 7235 16245 7240 16275
rect 7200 16240 7240 16245
rect 7280 16275 7320 16280
rect 7280 16245 7285 16275
rect 7315 16245 7320 16275
rect 7280 16240 7320 16245
rect 7360 16275 7400 16280
rect 7360 16245 7365 16275
rect 7395 16245 7400 16275
rect 7360 16240 7400 16245
rect 7440 16275 7480 16280
rect 7440 16245 7445 16275
rect 7475 16245 7480 16275
rect 7440 16240 7480 16245
rect 7520 16275 7560 16280
rect 7520 16245 7525 16275
rect 7555 16245 7560 16275
rect 7520 16240 7560 16245
rect 7600 16275 7640 16280
rect 7600 16245 7605 16275
rect 7635 16245 7640 16275
rect 7600 16240 7640 16245
rect 7680 16275 7720 16280
rect 7680 16245 7685 16275
rect 7715 16245 7720 16275
rect 7680 16240 7720 16245
rect 7760 16275 7800 16280
rect 7760 16245 7765 16275
rect 7795 16245 7800 16275
rect 7760 16240 7800 16245
rect 7840 16275 7880 16280
rect 7840 16245 7845 16275
rect 7875 16245 7880 16275
rect 7840 16240 7880 16245
rect 7920 16275 7960 16280
rect 7920 16245 7925 16275
rect 7955 16245 7960 16275
rect 7920 16240 7960 16245
rect 8000 16275 8040 16280
rect 8000 16245 8005 16275
rect 8035 16245 8040 16275
rect 8000 16240 8040 16245
rect 8080 16275 8120 16280
rect 8080 16245 8085 16275
rect 8115 16245 8120 16275
rect 8080 16240 8120 16245
rect 8160 16275 8200 16280
rect 8160 16245 8165 16275
rect 8195 16245 8200 16275
rect 8160 16240 8200 16245
rect 8240 16275 8280 16280
rect 8240 16245 8245 16275
rect 8275 16245 8280 16275
rect 8240 16240 8280 16245
rect 8320 16275 8360 16280
rect 8320 16245 8325 16275
rect 8355 16245 8360 16275
rect 8320 16240 8360 16245
rect 8400 16275 8440 16280
rect 8400 16245 8405 16275
rect 8435 16245 8440 16275
rect 8400 16240 8440 16245
rect 8480 16275 8520 16280
rect 8480 16245 8485 16275
rect 8515 16245 8520 16275
rect 8480 16240 8520 16245
rect 8560 16275 8600 16280
rect 8560 16245 8565 16275
rect 8595 16245 8600 16275
rect 8560 16240 8600 16245
rect 8640 16275 8680 16280
rect 8640 16245 8645 16275
rect 8675 16245 8680 16275
rect 8640 16240 8680 16245
rect 8720 16275 8760 16280
rect 8720 16245 8725 16275
rect 8755 16245 8760 16275
rect 8720 16240 8760 16245
rect 8800 16275 8840 16280
rect 8800 16245 8805 16275
rect 8835 16245 8840 16275
rect 8800 16240 8840 16245
rect 8880 16275 8920 16280
rect 8880 16245 8885 16275
rect 8915 16245 8920 16275
rect 8880 16240 8920 16245
rect 8960 16275 9000 16280
rect 8960 16245 8965 16275
rect 8995 16245 9000 16275
rect 8960 16240 9000 16245
rect 9040 16275 9080 16280
rect 9040 16245 9045 16275
rect 9075 16245 9080 16275
rect 9040 16240 9080 16245
rect 9120 16275 9160 16280
rect 9120 16245 9125 16275
rect 9155 16245 9160 16275
rect 9120 16240 9160 16245
rect 9200 16275 9240 16280
rect 9200 16245 9205 16275
rect 9235 16245 9240 16275
rect 9200 16240 9240 16245
rect 9280 16275 9320 16280
rect 9280 16245 9285 16275
rect 9315 16245 9320 16275
rect 9280 16240 9320 16245
rect 9360 16275 9400 16280
rect 9360 16245 9365 16275
rect 9395 16245 9400 16275
rect 9360 16240 9400 16245
rect 9440 16275 9480 16280
rect 9440 16245 9445 16275
rect 9475 16245 9480 16275
rect 9440 16240 9480 16245
rect 11560 16275 11600 16280
rect 11560 16245 11565 16275
rect 11595 16245 11600 16275
rect 11560 16240 11600 16245
rect 11640 16275 11680 16280
rect 11640 16245 11645 16275
rect 11675 16245 11680 16275
rect 11640 16240 11680 16245
rect 11720 16275 11760 16280
rect 11720 16245 11725 16275
rect 11755 16245 11760 16275
rect 11720 16240 11760 16245
rect 11800 16275 11840 16280
rect 11800 16245 11805 16275
rect 11835 16245 11840 16275
rect 11800 16240 11840 16245
rect 11880 16275 11920 16280
rect 11880 16245 11885 16275
rect 11915 16245 11920 16275
rect 11880 16240 11920 16245
rect 11960 16275 12000 16280
rect 11960 16245 11965 16275
rect 11995 16245 12000 16275
rect 11960 16240 12000 16245
rect 12040 16275 12080 16280
rect 12040 16245 12045 16275
rect 12075 16245 12080 16275
rect 12040 16240 12080 16245
rect 12120 16275 12160 16280
rect 12120 16245 12125 16275
rect 12155 16245 12160 16275
rect 12120 16240 12160 16245
rect 12200 16275 12240 16280
rect 12200 16245 12205 16275
rect 12235 16245 12240 16275
rect 12200 16240 12240 16245
rect 12280 16275 12320 16280
rect 12280 16245 12285 16275
rect 12315 16245 12320 16275
rect 12280 16240 12320 16245
rect 12360 16275 12400 16280
rect 12360 16245 12365 16275
rect 12395 16245 12400 16275
rect 12360 16240 12400 16245
rect 12440 16275 12480 16280
rect 12440 16245 12445 16275
rect 12475 16245 12480 16275
rect 12440 16240 12480 16245
rect 12520 16275 12560 16280
rect 12520 16245 12525 16275
rect 12555 16245 12560 16275
rect 12520 16240 12560 16245
rect 12600 16275 12640 16280
rect 12600 16245 12605 16275
rect 12635 16245 12640 16275
rect 12600 16240 12640 16245
rect 12680 16275 12720 16280
rect 12680 16245 12685 16275
rect 12715 16245 12720 16275
rect 12680 16240 12720 16245
rect 12760 16275 12800 16280
rect 12760 16245 12765 16275
rect 12795 16245 12800 16275
rect 12760 16240 12800 16245
rect 12840 16275 12880 16280
rect 12840 16245 12845 16275
rect 12875 16245 12880 16275
rect 12840 16240 12880 16245
rect 12920 16275 12960 16280
rect 12920 16245 12925 16275
rect 12955 16245 12960 16275
rect 12920 16240 12960 16245
rect 13000 16275 13040 16280
rect 13000 16245 13005 16275
rect 13035 16245 13040 16275
rect 13000 16240 13040 16245
rect 13080 16275 13120 16280
rect 13080 16245 13085 16275
rect 13115 16245 13120 16275
rect 13080 16240 13120 16245
rect 13160 16275 13200 16280
rect 13160 16245 13165 16275
rect 13195 16245 13200 16275
rect 13160 16240 13200 16245
rect 13240 16275 13280 16280
rect 13240 16245 13245 16275
rect 13275 16245 13280 16275
rect 13240 16240 13280 16245
rect 13320 16275 13360 16280
rect 13320 16245 13325 16275
rect 13355 16245 13360 16275
rect 13320 16240 13360 16245
rect 13400 16275 13440 16280
rect 13400 16245 13405 16275
rect 13435 16245 13440 16275
rect 13400 16240 13440 16245
rect 13480 16275 13520 16280
rect 13480 16245 13485 16275
rect 13515 16245 13520 16275
rect 13480 16240 13520 16245
rect 13560 16275 13600 16280
rect 13560 16245 13565 16275
rect 13595 16245 13600 16275
rect 13560 16240 13600 16245
rect 13640 16275 13680 16280
rect 13640 16245 13645 16275
rect 13675 16245 13680 16275
rect 13640 16240 13680 16245
rect 13720 16275 13760 16280
rect 13720 16245 13725 16275
rect 13755 16245 13760 16275
rect 13720 16240 13760 16245
rect 13800 16275 13840 16280
rect 13800 16245 13805 16275
rect 13835 16245 13840 16275
rect 13800 16240 13840 16245
rect 13880 16275 13920 16280
rect 13880 16245 13885 16275
rect 13915 16245 13920 16275
rect 13880 16240 13920 16245
rect 13960 16275 14000 16280
rect 13960 16245 13965 16275
rect 13995 16245 14000 16275
rect 13960 16240 14000 16245
rect 14040 16275 14080 16280
rect 14040 16245 14045 16275
rect 14075 16245 14080 16275
rect 14040 16240 14080 16245
rect 14120 16275 14160 16280
rect 14120 16245 14125 16275
rect 14155 16245 14160 16275
rect 14120 16240 14160 16245
rect 14200 16275 14240 16280
rect 14200 16245 14205 16275
rect 14235 16245 14240 16275
rect 14200 16240 14240 16245
rect 14280 16275 14320 16280
rect 14280 16245 14285 16275
rect 14315 16245 14320 16275
rect 14280 16240 14320 16245
rect 14360 16275 14400 16280
rect 14360 16245 14365 16275
rect 14395 16245 14400 16275
rect 14360 16240 14400 16245
rect 14440 16275 14480 16280
rect 14440 16245 14445 16275
rect 14475 16245 14480 16275
rect 14440 16240 14480 16245
rect 14520 16275 14560 16280
rect 14520 16245 14525 16275
rect 14555 16245 14560 16275
rect 14520 16240 14560 16245
rect 14600 16275 14640 16280
rect 14600 16245 14605 16275
rect 14635 16245 14640 16275
rect 14600 16240 14640 16245
rect 14680 16275 14720 16280
rect 14680 16245 14685 16275
rect 14715 16245 14720 16275
rect 14680 16240 14720 16245
rect 16760 16275 16800 16280
rect 16760 16245 16765 16275
rect 16795 16245 16800 16275
rect 16760 16240 16800 16245
rect 16840 16275 16880 16280
rect 16840 16245 16845 16275
rect 16875 16245 16880 16275
rect 16840 16240 16880 16245
rect 16920 16275 16960 16280
rect 16920 16245 16925 16275
rect 16955 16245 16960 16275
rect 16920 16240 16960 16245
rect 17000 16275 17040 16280
rect 17000 16245 17005 16275
rect 17035 16245 17040 16275
rect 17000 16240 17040 16245
rect 17080 16275 17120 16280
rect 17080 16245 17085 16275
rect 17115 16245 17120 16275
rect 17080 16240 17120 16245
rect 17160 16275 17200 16280
rect 17160 16245 17165 16275
rect 17195 16245 17200 16275
rect 17160 16240 17200 16245
rect 17240 16275 17280 16280
rect 17240 16245 17245 16275
rect 17275 16245 17280 16275
rect 17240 16240 17280 16245
rect 17320 16275 17360 16280
rect 17320 16245 17325 16275
rect 17355 16245 17360 16275
rect 17320 16240 17360 16245
rect 17400 16275 17440 16280
rect 17400 16245 17405 16275
rect 17435 16245 17440 16275
rect 17400 16240 17440 16245
rect 17480 16275 17520 16280
rect 17480 16245 17485 16275
rect 17515 16245 17520 16275
rect 17480 16240 17520 16245
rect 17560 16275 17600 16280
rect 17560 16245 17565 16275
rect 17595 16245 17600 16275
rect 17560 16240 17600 16245
rect 17640 16275 17680 16280
rect 17640 16245 17645 16275
rect 17675 16245 17680 16275
rect 17640 16240 17680 16245
rect 17720 16275 17760 16280
rect 17720 16245 17725 16275
rect 17755 16245 17760 16275
rect 17720 16240 17760 16245
rect 17800 16275 17840 16280
rect 17800 16245 17805 16275
rect 17835 16245 17840 16275
rect 17800 16240 17840 16245
rect 17880 16275 17920 16280
rect 17880 16245 17885 16275
rect 17915 16245 17920 16275
rect 17880 16240 17920 16245
rect 17960 16275 18000 16280
rect 17960 16245 17965 16275
rect 17995 16245 18000 16275
rect 17960 16240 18000 16245
rect 18040 16275 18080 16280
rect 18040 16245 18045 16275
rect 18075 16245 18080 16275
rect 18040 16240 18080 16245
rect 18120 16275 18160 16280
rect 18120 16245 18125 16275
rect 18155 16245 18160 16275
rect 18120 16240 18160 16245
rect 18200 16275 18240 16280
rect 18200 16245 18205 16275
rect 18235 16245 18240 16275
rect 18200 16240 18240 16245
rect 18280 16275 18320 16280
rect 18280 16245 18285 16275
rect 18315 16245 18320 16275
rect 18280 16240 18320 16245
rect 18360 16275 18400 16280
rect 18360 16245 18365 16275
rect 18395 16245 18400 16275
rect 18360 16240 18400 16245
rect 18440 16275 18480 16280
rect 18440 16245 18445 16275
rect 18475 16245 18480 16275
rect 18440 16240 18480 16245
rect 18520 16275 18560 16280
rect 18520 16245 18525 16275
rect 18555 16245 18560 16275
rect 18520 16240 18560 16245
rect 18600 16275 18640 16280
rect 18600 16245 18605 16275
rect 18635 16245 18640 16275
rect 18600 16240 18640 16245
rect 18680 16275 18720 16280
rect 18680 16245 18685 16275
rect 18715 16245 18720 16275
rect 18680 16240 18720 16245
rect 18760 16275 18800 16280
rect 18760 16245 18765 16275
rect 18795 16245 18800 16275
rect 18760 16240 18800 16245
rect 18840 16275 18880 16280
rect 18840 16245 18845 16275
rect 18875 16245 18880 16275
rect 18840 16240 18880 16245
rect 18920 16275 18960 16280
rect 18920 16245 18925 16275
rect 18955 16245 18960 16275
rect 18920 16240 18960 16245
rect 19000 16275 19040 16280
rect 19000 16245 19005 16275
rect 19035 16245 19040 16275
rect 19000 16240 19040 16245
rect 19080 16275 19120 16280
rect 19080 16245 19085 16275
rect 19115 16245 19120 16275
rect 19080 16240 19120 16245
rect 19160 16275 19200 16280
rect 19160 16245 19165 16275
rect 19195 16245 19200 16275
rect 19160 16240 19200 16245
rect 19240 16275 19280 16280
rect 19240 16245 19245 16275
rect 19275 16245 19280 16275
rect 19240 16240 19280 16245
rect 19320 16275 19360 16280
rect 19320 16245 19325 16275
rect 19355 16245 19360 16275
rect 19320 16240 19360 16245
rect 19400 16275 19440 16280
rect 19400 16245 19405 16275
rect 19435 16245 19440 16275
rect 19400 16240 19440 16245
rect 19480 16275 19520 16280
rect 19480 16245 19485 16275
rect 19515 16245 19520 16275
rect 19480 16240 19520 16245
rect 19560 16275 19600 16280
rect 19560 16245 19565 16275
rect 19595 16245 19600 16275
rect 19560 16240 19600 16245
rect 19640 16275 19680 16280
rect 19640 16245 19645 16275
rect 19675 16245 19680 16275
rect 19640 16240 19680 16245
rect 19720 16275 19760 16280
rect 19720 16245 19725 16275
rect 19755 16245 19760 16275
rect 19720 16240 19760 16245
rect 19800 16275 19840 16280
rect 19800 16245 19805 16275
rect 19835 16245 19840 16275
rect 19800 16240 19840 16245
rect 19880 16275 19920 16280
rect 19880 16245 19885 16275
rect 19915 16245 19920 16275
rect 19880 16240 19920 16245
rect 19960 16275 20000 16280
rect 19960 16245 19965 16275
rect 19995 16245 20000 16275
rect 19960 16240 20000 16245
rect 20040 16275 20080 16280
rect 20040 16245 20045 16275
rect 20075 16245 20080 16275
rect 20040 16240 20080 16245
rect 20120 16275 20160 16280
rect 20120 16245 20125 16275
rect 20155 16245 20160 16275
rect 20120 16240 20160 16245
rect 20200 16275 20240 16280
rect 20200 16245 20205 16275
rect 20235 16245 20240 16275
rect 20200 16240 20240 16245
rect 20280 16275 20320 16280
rect 20280 16245 20285 16275
rect 20315 16245 20320 16275
rect 20280 16240 20320 16245
rect 20360 16275 20400 16280
rect 20360 16245 20365 16275
rect 20395 16245 20400 16275
rect 20360 16240 20400 16245
rect 20440 16275 20480 16280
rect 20440 16245 20445 16275
rect 20475 16245 20480 16275
rect 20440 16240 20480 16245
rect 20520 16275 20560 16280
rect 20520 16245 20525 16275
rect 20555 16245 20560 16275
rect 20520 16240 20560 16245
rect 20600 16275 20640 16280
rect 20600 16245 20605 16275
rect 20635 16245 20640 16275
rect 20600 16240 20640 16245
rect 20680 16275 20720 16280
rect 20680 16245 20685 16275
rect 20715 16245 20720 16275
rect 20680 16240 20720 16245
rect 20760 16275 20800 16280
rect 20760 16245 20765 16275
rect 20795 16245 20800 16275
rect 20760 16240 20800 16245
rect 20840 16275 20880 16280
rect 20840 16245 20845 16275
rect 20875 16245 20880 16275
rect 20840 16240 20880 16245
rect 20920 16275 20960 16280
rect 20920 16245 20925 16275
rect 20955 16245 20960 16275
rect 20920 16240 20960 16245
rect 0 16195 40 16200
rect 0 16165 5 16195
rect 35 16165 40 16195
rect 0 16160 40 16165
rect 80 16195 120 16200
rect 80 16165 85 16195
rect 115 16165 120 16195
rect 80 16160 120 16165
rect 160 16195 200 16200
rect 160 16165 165 16195
rect 195 16165 200 16195
rect 160 16160 200 16165
rect 240 16195 280 16200
rect 240 16165 245 16195
rect 275 16165 280 16195
rect 240 16160 280 16165
rect 320 16195 360 16200
rect 320 16165 325 16195
rect 355 16165 360 16195
rect 320 16160 360 16165
rect 400 16195 440 16200
rect 400 16165 405 16195
rect 435 16165 440 16195
rect 400 16160 440 16165
rect 480 16195 520 16200
rect 480 16165 485 16195
rect 515 16165 520 16195
rect 480 16160 520 16165
rect 560 16195 600 16200
rect 560 16165 565 16195
rect 595 16165 600 16195
rect 560 16160 600 16165
rect 640 16195 680 16200
rect 640 16165 645 16195
rect 675 16165 680 16195
rect 640 16160 680 16165
rect 720 16195 760 16200
rect 720 16165 725 16195
rect 755 16165 760 16195
rect 720 16160 760 16165
rect 800 16195 840 16200
rect 800 16165 805 16195
rect 835 16165 840 16195
rect 800 16160 840 16165
rect 880 16195 920 16200
rect 880 16165 885 16195
rect 915 16165 920 16195
rect 880 16160 920 16165
rect 960 16195 1000 16200
rect 960 16165 965 16195
rect 995 16165 1000 16195
rect 960 16160 1000 16165
rect 1040 16195 1080 16200
rect 1040 16165 1045 16195
rect 1075 16165 1080 16195
rect 1040 16160 1080 16165
rect 1120 16195 1160 16200
rect 1120 16165 1125 16195
rect 1155 16165 1160 16195
rect 1120 16160 1160 16165
rect 1200 16195 1240 16200
rect 1200 16165 1205 16195
rect 1235 16165 1240 16195
rect 1200 16160 1240 16165
rect 1280 16195 1320 16200
rect 1280 16165 1285 16195
rect 1315 16165 1320 16195
rect 1280 16160 1320 16165
rect 1360 16195 1400 16200
rect 1360 16165 1365 16195
rect 1395 16165 1400 16195
rect 1360 16160 1400 16165
rect 1440 16195 1480 16200
rect 1440 16165 1445 16195
rect 1475 16165 1480 16195
rect 1440 16160 1480 16165
rect 1520 16195 1560 16200
rect 1520 16165 1525 16195
rect 1555 16165 1560 16195
rect 1520 16160 1560 16165
rect 1600 16195 1640 16200
rect 1600 16165 1605 16195
rect 1635 16165 1640 16195
rect 1600 16160 1640 16165
rect 1680 16195 1720 16200
rect 1680 16165 1685 16195
rect 1715 16165 1720 16195
rect 1680 16160 1720 16165
rect 1760 16195 1800 16200
rect 1760 16165 1765 16195
rect 1795 16165 1800 16195
rect 1760 16160 1800 16165
rect 1840 16195 1880 16200
rect 1840 16165 1845 16195
rect 1875 16165 1880 16195
rect 1840 16160 1880 16165
rect 1920 16195 1960 16200
rect 1920 16165 1925 16195
rect 1955 16165 1960 16195
rect 1920 16160 1960 16165
rect 2000 16195 2040 16200
rect 2000 16165 2005 16195
rect 2035 16165 2040 16195
rect 2000 16160 2040 16165
rect 2080 16195 2120 16200
rect 2080 16165 2085 16195
rect 2115 16165 2120 16195
rect 2080 16160 2120 16165
rect 2160 16195 2200 16200
rect 2160 16165 2165 16195
rect 2195 16165 2200 16195
rect 2160 16160 2200 16165
rect 2240 16195 2280 16200
rect 2240 16165 2245 16195
rect 2275 16165 2280 16195
rect 2240 16160 2280 16165
rect 2320 16195 2360 16200
rect 2320 16165 2325 16195
rect 2355 16165 2360 16195
rect 2320 16160 2360 16165
rect 2400 16195 2440 16200
rect 2400 16165 2405 16195
rect 2435 16165 2440 16195
rect 2400 16160 2440 16165
rect 2480 16195 2520 16200
rect 2480 16165 2485 16195
rect 2515 16165 2520 16195
rect 2480 16160 2520 16165
rect 2560 16195 2600 16200
rect 2560 16165 2565 16195
rect 2595 16165 2600 16195
rect 2560 16160 2600 16165
rect 2640 16195 2680 16200
rect 2640 16165 2645 16195
rect 2675 16165 2680 16195
rect 2640 16160 2680 16165
rect 2720 16195 2760 16200
rect 2720 16165 2725 16195
rect 2755 16165 2760 16195
rect 2720 16160 2760 16165
rect 2800 16195 2840 16200
rect 2800 16165 2805 16195
rect 2835 16165 2840 16195
rect 2800 16160 2840 16165
rect 2880 16195 2920 16200
rect 2880 16165 2885 16195
rect 2915 16165 2920 16195
rect 2880 16160 2920 16165
rect 2960 16195 3000 16200
rect 2960 16165 2965 16195
rect 2995 16165 3000 16195
rect 2960 16160 3000 16165
rect 3040 16195 3080 16200
rect 3040 16165 3045 16195
rect 3075 16165 3080 16195
rect 3040 16160 3080 16165
rect 3120 16195 3160 16200
rect 3120 16165 3125 16195
rect 3155 16165 3160 16195
rect 3120 16160 3160 16165
rect 3200 16195 3240 16200
rect 3200 16165 3205 16195
rect 3235 16165 3240 16195
rect 3200 16160 3240 16165
rect 3280 16195 3320 16200
rect 3280 16165 3285 16195
rect 3315 16165 3320 16195
rect 3280 16160 3320 16165
rect 3360 16195 3400 16200
rect 3360 16165 3365 16195
rect 3395 16165 3400 16195
rect 3360 16160 3400 16165
rect 3440 16195 3480 16200
rect 3440 16165 3445 16195
rect 3475 16165 3480 16195
rect 3440 16160 3480 16165
rect 3520 16195 3560 16200
rect 3520 16165 3525 16195
rect 3555 16165 3560 16195
rect 3520 16160 3560 16165
rect 3600 16195 3640 16200
rect 3600 16165 3605 16195
rect 3635 16165 3640 16195
rect 3600 16160 3640 16165
rect 3680 16195 3720 16200
rect 3680 16165 3685 16195
rect 3715 16165 3720 16195
rect 3680 16160 3720 16165
rect 3760 16195 3800 16200
rect 3760 16165 3765 16195
rect 3795 16165 3800 16195
rect 3760 16160 3800 16165
rect 3840 16195 3880 16200
rect 3840 16165 3845 16195
rect 3875 16165 3880 16195
rect 3840 16160 3880 16165
rect 3920 16195 3960 16200
rect 3920 16165 3925 16195
rect 3955 16165 3960 16195
rect 3920 16160 3960 16165
rect 4000 16195 4040 16200
rect 4000 16165 4005 16195
rect 4035 16165 4040 16195
rect 4000 16160 4040 16165
rect 4080 16195 4120 16200
rect 4080 16165 4085 16195
rect 4115 16165 4120 16195
rect 4080 16160 4120 16165
rect 4160 16195 4200 16200
rect 4160 16165 4165 16195
rect 4195 16165 4200 16195
rect 4160 16160 4200 16165
rect 6240 16195 6280 16200
rect 6240 16165 6245 16195
rect 6275 16165 6280 16195
rect 6240 16160 6280 16165
rect 6320 16195 6360 16200
rect 6320 16165 6325 16195
rect 6355 16165 6360 16195
rect 6320 16160 6360 16165
rect 6400 16195 6440 16200
rect 6400 16165 6405 16195
rect 6435 16165 6440 16195
rect 6400 16160 6440 16165
rect 6480 16195 6520 16200
rect 6480 16165 6485 16195
rect 6515 16165 6520 16195
rect 6480 16160 6520 16165
rect 6560 16195 6600 16200
rect 6560 16165 6565 16195
rect 6595 16165 6600 16195
rect 6560 16160 6600 16165
rect 6640 16195 6680 16200
rect 6640 16165 6645 16195
rect 6675 16165 6680 16195
rect 6640 16160 6680 16165
rect 6720 16195 6760 16200
rect 6720 16165 6725 16195
rect 6755 16165 6760 16195
rect 6720 16160 6760 16165
rect 6800 16195 6840 16200
rect 6800 16165 6805 16195
rect 6835 16165 6840 16195
rect 6800 16160 6840 16165
rect 6880 16195 6920 16200
rect 6880 16165 6885 16195
rect 6915 16165 6920 16195
rect 6880 16160 6920 16165
rect 6960 16195 7000 16200
rect 6960 16165 6965 16195
rect 6995 16165 7000 16195
rect 6960 16160 7000 16165
rect 7040 16195 7080 16200
rect 7040 16165 7045 16195
rect 7075 16165 7080 16195
rect 7040 16160 7080 16165
rect 7120 16195 7160 16200
rect 7120 16165 7125 16195
rect 7155 16165 7160 16195
rect 7120 16160 7160 16165
rect 7200 16195 7240 16200
rect 7200 16165 7205 16195
rect 7235 16165 7240 16195
rect 7200 16160 7240 16165
rect 7280 16195 7320 16200
rect 7280 16165 7285 16195
rect 7315 16165 7320 16195
rect 7280 16160 7320 16165
rect 7360 16195 7400 16200
rect 7360 16165 7365 16195
rect 7395 16165 7400 16195
rect 7360 16160 7400 16165
rect 7440 16195 7480 16200
rect 7440 16165 7445 16195
rect 7475 16165 7480 16195
rect 7440 16160 7480 16165
rect 7520 16195 7560 16200
rect 7520 16165 7525 16195
rect 7555 16165 7560 16195
rect 7520 16160 7560 16165
rect 7600 16195 7640 16200
rect 7600 16165 7605 16195
rect 7635 16165 7640 16195
rect 7600 16160 7640 16165
rect 7680 16195 7720 16200
rect 7680 16165 7685 16195
rect 7715 16165 7720 16195
rect 7680 16160 7720 16165
rect 7760 16195 7800 16200
rect 7760 16165 7765 16195
rect 7795 16165 7800 16195
rect 7760 16160 7800 16165
rect 7840 16195 7880 16200
rect 7840 16165 7845 16195
rect 7875 16165 7880 16195
rect 7840 16160 7880 16165
rect 7920 16195 7960 16200
rect 7920 16165 7925 16195
rect 7955 16165 7960 16195
rect 7920 16160 7960 16165
rect 8000 16195 8040 16200
rect 8000 16165 8005 16195
rect 8035 16165 8040 16195
rect 8000 16160 8040 16165
rect 8080 16195 8120 16200
rect 8080 16165 8085 16195
rect 8115 16165 8120 16195
rect 8080 16160 8120 16165
rect 8160 16195 8200 16200
rect 8160 16165 8165 16195
rect 8195 16165 8200 16195
rect 8160 16160 8200 16165
rect 8240 16195 8280 16200
rect 8240 16165 8245 16195
rect 8275 16165 8280 16195
rect 8240 16160 8280 16165
rect 8320 16195 8360 16200
rect 8320 16165 8325 16195
rect 8355 16165 8360 16195
rect 8320 16160 8360 16165
rect 8400 16195 8440 16200
rect 8400 16165 8405 16195
rect 8435 16165 8440 16195
rect 8400 16160 8440 16165
rect 8480 16195 8520 16200
rect 8480 16165 8485 16195
rect 8515 16165 8520 16195
rect 8480 16160 8520 16165
rect 8560 16195 8600 16200
rect 8560 16165 8565 16195
rect 8595 16165 8600 16195
rect 8560 16160 8600 16165
rect 8640 16195 8680 16200
rect 8640 16165 8645 16195
rect 8675 16165 8680 16195
rect 8640 16160 8680 16165
rect 8720 16195 8760 16200
rect 8720 16165 8725 16195
rect 8755 16165 8760 16195
rect 8720 16160 8760 16165
rect 8800 16195 8840 16200
rect 8800 16165 8805 16195
rect 8835 16165 8840 16195
rect 8800 16160 8840 16165
rect 8880 16195 8920 16200
rect 8880 16165 8885 16195
rect 8915 16165 8920 16195
rect 8880 16160 8920 16165
rect 8960 16195 9000 16200
rect 8960 16165 8965 16195
rect 8995 16165 9000 16195
rect 8960 16160 9000 16165
rect 9040 16195 9080 16200
rect 9040 16165 9045 16195
rect 9075 16165 9080 16195
rect 9040 16160 9080 16165
rect 9120 16195 9160 16200
rect 9120 16165 9125 16195
rect 9155 16165 9160 16195
rect 9120 16160 9160 16165
rect 9200 16195 9240 16200
rect 9200 16165 9205 16195
rect 9235 16165 9240 16195
rect 9200 16160 9240 16165
rect 9280 16195 9320 16200
rect 9280 16165 9285 16195
rect 9315 16165 9320 16195
rect 9280 16160 9320 16165
rect 9360 16195 9400 16200
rect 9360 16165 9365 16195
rect 9395 16165 9400 16195
rect 9360 16160 9400 16165
rect 9440 16195 9480 16200
rect 9440 16165 9445 16195
rect 9475 16165 9480 16195
rect 9440 16160 9480 16165
rect 11560 16195 11600 16200
rect 11560 16165 11565 16195
rect 11595 16165 11600 16195
rect 11560 16160 11600 16165
rect 11640 16195 11680 16200
rect 11640 16165 11645 16195
rect 11675 16165 11680 16195
rect 11640 16160 11680 16165
rect 11720 16195 11760 16200
rect 11720 16165 11725 16195
rect 11755 16165 11760 16195
rect 11720 16160 11760 16165
rect 11800 16195 11840 16200
rect 11800 16165 11805 16195
rect 11835 16165 11840 16195
rect 11800 16160 11840 16165
rect 11880 16195 11920 16200
rect 11880 16165 11885 16195
rect 11915 16165 11920 16195
rect 11880 16160 11920 16165
rect 11960 16195 12000 16200
rect 11960 16165 11965 16195
rect 11995 16165 12000 16195
rect 11960 16160 12000 16165
rect 12040 16195 12080 16200
rect 12040 16165 12045 16195
rect 12075 16165 12080 16195
rect 12040 16160 12080 16165
rect 12120 16195 12160 16200
rect 12120 16165 12125 16195
rect 12155 16165 12160 16195
rect 12120 16160 12160 16165
rect 12200 16195 12240 16200
rect 12200 16165 12205 16195
rect 12235 16165 12240 16195
rect 12200 16160 12240 16165
rect 12280 16195 12320 16200
rect 12280 16165 12285 16195
rect 12315 16165 12320 16195
rect 12280 16160 12320 16165
rect 12360 16195 12400 16200
rect 12360 16165 12365 16195
rect 12395 16165 12400 16195
rect 12360 16160 12400 16165
rect 12440 16195 12480 16200
rect 12440 16165 12445 16195
rect 12475 16165 12480 16195
rect 12440 16160 12480 16165
rect 12520 16195 12560 16200
rect 12520 16165 12525 16195
rect 12555 16165 12560 16195
rect 12520 16160 12560 16165
rect 12600 16195 12640 16200
rect 12600 16165 12605 16195
rect 12635 16165 12640 16195
rect 12600 16160 12640 16165
rect 12680 16195 12720 16200
rect 12680 16165 12685 16195
rect 12715 16165 12720 16195
rect 12680 16160 12720 16165
rect 12760 16195 12800 16200
rect 12760 16165 12765 16195
rect 12795 16165 12800 16195
rect 12760 16160 12800 16165
rect 12840 16195 12880 16200
rect 12840 16165 12845 16195
rect 12875 16165 12880 16195
rect 12840 16160 12880 16165
rect 12920 16195 12960 16200
rect 12920 16165 12925 16195
rect 12955 16165 12960 16195
rect 12920 16160 12960 16165
rect 13000 16195 13040 16200
rect 13000 16165 13005 16195
rect 13035 16165 13040 16195
rect 13000 16160 13040 16165
rect 13080 16195 13120 16200
rect 13080 16165 13085 16195
rect 13115 16165 13120 16195
rect 13080 16160 13120 16165
rect 13160 16195 13200 16200
rect 13160 16165 13165 16195
rect 13195 16165 13200 16195
rect 13160 16160 13200 16165
rect 13240 16195 13280 16200
rect 13240 16165 13245 16195
rect 13275 16165 13280 16195
rect 13240 16160 13280 16165
rect 13320 16195 13360 16200
rect 13320 16165 13325 16195
rect 13355 16165 13360 16195
rect 13320 16160 13360 16165
rect 13400 16195 13440 16200
rect 13400 16165 13405 16195
rect 13435 16165 13440 16195
rect 13400 16160 13440 16165
rect 13480 16195 13520 16200
rect 13480 16165 13485 16195
rect 13515 16165 13520 16195
rect 13480 16160 13520 16165
rect 13560 16195 13600 16200
rect 13560 16165 13565 16195
rect 13595 16165 13600 16195
rect 13560 16160 13600 16165
rect 13640 16195 13680 16200
rect 13640 16165 13645 16195
rect 13675 16165 13680 16195
rect 13640 16160 13680 16165
rect 13720 16195 13760 16200
rect 13720 16165 13725 16195
rect 13755 16165 13760 16195
rect 13720 16160 13760 16165
rect 13800 16195 13840 16200
rect 13800 16165 13805 16195
rect 13835 16165 13840 16195
rect 13800 16160 13840 16165
rect 13880 16195 13920 16200
rect 13880 16165 13885 16195
rect 13915 16165 13920 16195
rect 13880 16160 13920 16165
rect 13960 16195 14000 16200
rect 13960 16165 13965 16195
rect 13995 16165 14000 16195
rect 13960 16160 14000 16165
rect 14040 16195 14080 16200
rect 14040 16165 14045 16195
rect 14075 16165 14080 16195
rect 14040 16160 14080 16165
rect 14120 16195 14160 16200
rect 14120 16165 14125 16195
rect 14155 16165 14160 16195
rect 14120 16160 14160 16165
rect 14200 16195 14240 16200
rect 14200 16165 14205 16195
rect 14235 16165 14240 16195
rect 14200 16160 14240 16165
rect 14280 16195 14320 16200
rect 14280 16165 14285 16195
rect 14315 16165 14320 16195
rect 14280 16160 14320 16165
rect 14360 16195 14400 16200
rect 14360 16165 14365 16195
rect 14395 16165 14400 16195
rect 14360 16160 14400 16165
rect 14440 16195 14480 16200
rect 14440 16165 14445 16195
rect 14475 16165 14480 16195
rect 14440 16160 14480 16165
rect 14520 16195 14560 16200
rect 14520 16165 14525 16195
rect 14555 16165 14560 16195
rect 14520 16160 14560 16165
rect 14600 16195 14640 16200
rect 14600 16165 14605 16195
rect 14635 16165 14640 16195
rect 14600 16160 14640 16165
rect 14680 16195 14720 16200
rect 14680 16165 14685 16195
rect 14715 16165 14720 16195
rect 14680 16160 14720 16165
rect 16760 16195 16800 16200
rect 16760 16165 16765 16195
rect 16795 16165 16800 16195
rect 16760 16160 16800 16165
rect 16840 16195 16880 16200
rect 16840 16165 16845 16195
rect 16875 16165 16880 16195
rect 16840 16160 16880 16165
rect 16920 16195 16960 16200
rect 16920 16165 16925 16195
rect 16955 16165 16960 16195
rect 16920 16160 16960 16165
rect 17000 16195 17040 16200
rect 17000 16165 17005 16195
rect 17035 16165 17040 16195
rect 17000 16160 17040 16165
rect 17080 16195 17120 16200
rect 17080 16165 17085 16195
rect 17115 16165 17120 16195
rect 17080 16160 17120 16165
rect 17160 16195 17200 16200
rect 17160 16165 17165 16195
rect 17195 16165 17200 16195
rect 17160 16160 17200 16165
rect 17240 16195 17280 16200
rect 17240 16165 17245 16195
rect 17275 16165 17280 16195
rect 17240 16160 17280 16165
rect 17320 16195 17360 16200
rect 17320 16165 17325 16195
rect 17355 16165 17360 16195
rect 17320 16160 17360 16165
rect 17400 16195 17440 16200
rect 17400 16165 17405 16195
rect 17435 16165 17440 16195
rect 17400 16160 17440 16165
rect 17480 16195 17520 16200
rect 17480 16165 17485 16195
rect 17515 16165 17520 16195
rect 17480 16160 17520 16165
rect 17560 16195 17600 16200
rect 17560 16165 17565 16195
rect 17595 16165 17600 16195
rect 17560 16160 17600 16165
rect 17640 16195 17680 16200
rect 17640 16165 17645 16195
rect 17675 16165 17680 16195
rect 17640 16160 17680 16165
rect 17720 16195 17760 16200
rect 17720 16165 17725 16195
rect 17755 16165 17760 16195
rect 17720 16160 17760 16165
rect 17800 16195 17840 16200
rect 17800 16165 17805 16195
rect 17835 16165 17840 16195
rect 17800 16160 17840 16165
rect 17880 16195 17920 16200
rect 17880 16165 17885 16195
rect 17915 16165 17920 16195
rect 17880 16160 17920 16165
rect 17960 16195 18000 16200
rect 17960 16165 17965 16195
rect 17995 16165 18000 16195
rect 17960 16160 18000 16165
rect 18040 16195 18080 16200
rect 18040 16165 18045 16195
rect 18075 16165 18080 16195
rect 18040 16160 18080 16165
rect 18120 16195 18160 16200
rect 18120 16165 18125 16195
rect 18155 16165 18160 16195
rect 18120 16160 18160 16165
rect 18200 16195 18240 16200
rect 18200 16165 18205 16195
rect 18235 16165 18240 16195
rect 18200 16160 18240 16165
rect 18280 16195 18320 16200
rect 18280 16165 18285 16195
rect 18315 16165 18320 16195
rect 18280 16160 18320 16165
rect 18360 16195 18400 16200
rect 18360 16165 18365 16195
rect 18395 16165 18400 16195
rect 18360 16160 18400 16165
rect 18440 16195 18480 16200
rect 18440 16165 18445 16195
rect 18475 16165 18480 16195
rect 18440 16160 18480 16165
rect 18520 16195 18560 16200
rect 18520 16165 18525 16195
rect 18555 16165 18560 16195
rect 18520 16160 18560 16165
rect 18600 16195 18640 16200
rect 18600 16165 18605 16195
rect 18635 16165 18640 16195
rect 18600 16160 18640 16165
rect 18680 16195 18720 16200
rect 18680 16165 18685 16195
rect 18715 16165 18720 16195
rect 18680 16160 18720 16165
rect 18760 16195 18800 16200
rect 18760 16165 18765 16195
rect 18795 16165 18800 16195
rect 18760 16160 18800 16165
rect 18840 16195 18880 16200
rect 18840 16165 18845 16195
rect 18875 16165 18880 16195
rect 18840 16160 18880 16165
rect 18920 16195 18960 16200
rect 18920 16165 18925 16195
rect 18955 16165 18960 16195
rect 18920 16160 18960 16165
rect 19000 16195 19040 16200
rect 19000 16165 19005 16195
rect 19035 16165 19040 16195
rect 19000 16160 19040 16165
rect 19080 16195 19120 16200
rect 19080 16165 19085 16195
rect 19115 16165 19120 16195
rect 19080 16160 19120 16165
rect 19160 16195 19200 16200
rect 19160 16165 19165 16195
rect 19195 16165 19200 16195
rect 19160 16160 19200 16165
rect 19240 16195 19280 16200
rect 19240 16165 19245 16195
rect 19275 16165 19280 16195
rect 19240 16160 19280 16165
rect 19320 16195 19360 16200
rect 19320 16165 19325 16195
rect 19355 16165 19360 16195
rect 19320 16160 19360 16165
rect 19400 16195 19440 16200
rect 19400 16165 19405 16195
rect 19435 16165 19440 16195
rect 19400 16160 19440 16165
rect 19480 16195 19520 16200
rect 19480 16165 19485 16195
rect 19515 16165 19520 16195
rect 19480 16160 19520 16165
rect 19560 16195 19600 16200
rect 19560 16165 19565 16195
rect 19595 16165 19600 16195
rect 19560 16160 19600 16165
rect 19640 16195 19680 16200
rect 19640 16165 19645 16195
rect 19675 16165 19680 16195
rect 19640 16160 19680 16165
rect 19720 16195 19760 16200
rect 19720 16165 19725 16195
rect 19755 16165 19760 16195
rect 19720 16160 19760 16165
rect 19800 16195 19840 16200
rect 19800 16165 19805 16195
rect 19835 16165 19840 16195
rect 19800 16160 19840 16165
rect 19880 16195 19920 16200
rect 19880 16165 19885 16195
rect 19915 16165 19920 16195
rect 19880 16160 19920 16165
rect 19960 16195 20000 16200
rect 19960 16165 19965 16195
rect 19995 16165 20000 16195
rect 19960 16160 20000 16165
rect 20040 16195 20080 16200
rect 20040 16165 20045 16195
rect 20075 16165 20080 16195
rect 20040 16160 20080 16165
rect 20120 16195 20160 16200
rect 20120 16165 20125 16195
rect 20155 16165 20160 16195
rect 20120 16160 20160 16165
rect 20200 16195 20240 16200
rect 20200 16165 20205 16195
rect 20235 16165 20240 16195
rect 20200 16160 20240 16165
rect 20280 16195 20320 16200
rect 20280 16165 20285 16195
rect 20315 16165 20320 16195
rect 20280 16160 20320 16165
rect 20360 16195 20400 16200
rect 20360 16165 20365 16195
rect 20395 16165 20400 16195
rect 20360 16160 20400 16165
rect 20440 16195 20480 16200
rect 20440 16165 20445 16195
rect 20475 16165 20480 16195
rect 20440 16160 20480 16165
rect 20520 16195 20560 16200
rect 20520 16165 20525 16195
rect 20555 16165 20560 16195
rect 20520 16160 20560 16165
rect 20600 16195 20640 16200
rect 20600 16165 20605 16195
rect 20635 16165 20640 16195
rect 20600 16160 20640 16165
rect 20680 16195 20720 16200
rect 20680 16165 20685 16195
rect 20715 16165 20720 16195
rect 20680 16160 20720 16165
rect 20760 16195 20800 16200
rect 20760 16165 20765 16195
rect 20795 16165 20800 16195
rect 20760 16160 20800 16165
rect 20840 16195 20880 16200
rect 20840 16165 20845 16195
rect 20875 16165 20880 16195
rect 20840 16160 20880 16165
rect 20920 16195 20960 16200
rect 20920 16165 20925 16195
rect 20955 16165 20960 16195
rect 20920 16160 20960 16165
rect 0 16035 40 16040
rect 0 16005 5 16035
rect 35 16005 40 16035
rect 0 16000 40 16005
rect 80 16035 120 16040
rect 80 16005 85 16035
rect 115 16005 120 16035
rect 80 16000 120 16005
rect 160 16035 200 16040
rect 160 16005 165 16035
rect 195 16005 200 16035
rect 160 16000 200 16005
rect 240 16035 280 16040
rect 240 16005 245 16035
rect 275 16005 280 16035
rect 240 16000 280 16005
rect 320 16035 360 16040
rect 320 16005 325 16035
rect 355 16005 360 16035
rect 320 16000 360 16005
rect 400 16035 440 16040
rect 400 16005 405 16035
rect 435 16005 440 16035
rect 400 16000 440 16005
rect 480 16035 520 16040
rect 480 16005 485 16035
rect 515 16005 520 16035
rect 480 16000 520 16005
rect 560 16035 600 16040
rect 560 16005 565 16035
rect 595 16005 600 16035
rect 560 16000 600 16005
rect 640 16035 680 16040
rect 640 16005 645 16035
rect 675 16005 680 16035
rect 640 16000 680 16005
rect 720 16035 760 16040
rect 720 16005 725 16035
rect 755 16005 760 16035
rect 720 16000 760 16005
rect 800 16035 840 16040
rect 800 16005 805 16035
rect 835 16005 840 16035
rect 800 16000 840 16005
rect 880 16035 920 16040
rect 880 16005 885 16035
rect 915 16005 920 16035
rect 880 16000 920 16005
rect 960 16035 1000 16040
rect 960 16005 965 16035
rect 995 16005 1000 16035
rect 960 16000 1000 16005
rect 1040 16035 1080 16040
rect 1040 16005 1045 16035
rect 1075 16005 1080 16035
rect 1040 16000 1080 16005
rect 1120 16035 1160 16040
rect 1120 16005 1125 16035
rect 1155 16005 1160 16035
rect 1120 16000 1160 16005
rect 1200 16035 1240 16040
rect 1200 16005 1205 16035
rect 1235 16005 1240 16035
rect 1200 16000 1240 16005
rect 1280 16035 1320 16040
rect 1280 16005 1285 16035
rect 1315 16005 1320 16035
rect 1280 16000 1320 16005
rect 1360 16035 1400 16040
rect 1360 16005 1365 16035
rect 1395 16005 1400 16035
rect 1360 16000 1400 16005
rect 1440 16035 1480 16040
rect 1440 16005 1445 16035
rect 1475 16005 1480 16035
rect 1440 16000 1480 16005
rect 1520 16035 1560 16040
rect 1520 16005 1525 16035
rect 1555 16005 1560 16035
rect 1520 16000 1560 16005
rect 1600 16035 1640 16040
rect 1600 16005 1605 16035
rect 1635 16005 1640 16035
rect 1600 16000 1640 16005
rect 1680 16035 1720 16040
rect 1680 16005 1685 16035
rect 1715 16005 1720 16035
rect 1680 16000 1720 16005
rect 1760 16035 1800 16040
rect 1760 16005 1765 16035
rect 1795 16005 1800 16035
rect 1760 16000 1800 16005
rect 1840 16035 1880 16040
rect 1840 16005 1845 16035
rect 1875 16005 1880 16035
rect 1840 16000 1880 16005
rect 1920 16035 1960 16040
rect 1920 16005 1925 16035
rect 1955 16005 1960 16035
rect 1920 16000 1960 16005
rect 2000 16035 2040 16040
rect 2000 16005 2005 16035
rect 2035 16005 2040 16035
rect 2000 16000 2040 16005
rect 2080 16035 2120 16040
rect 2080 16005 2085 16035
rect 2115 16005 2120 16035
rect 2080 16000 2120 16005
rect 2160 16035 2200 16040
rect 2160 16005 2165 16035
rect 2195 16005 2200 16035
rect 2160 16000 2200 16005
rect 2240 16035 2280 16040
rect 2240 16005 2245 16035
rect 2275 16005 2280 16035
rect 2240 16000 2280 16005
rect 2320 16035 2360 16040
rect 2320 16005 2325 16035
rect 2355 16005 2360 16035
rect 2320 16000 2360 16005
rect 2400 16035 2440 16040
rect 2400 16005 2405 16035
rect 2435 16005 2440 16035
rect 2400 16000 2440 16005
rect 2480 16035 2520 16040
rect 2480 16005 2485 16035
rect 2515 16005 2520 16035
rect 2480 16000 2520 16005
rect 2560 16035 2600 16040
rect 2560 16005 2565 16035
rect 2595 16005 2600 16035
rect 2560 16000 2600 16005
rect 2640 16035 2680 16040
rect 2640 16005 2645 16035
rect 2675 16005 2680 16035
rect 2640 16000 2680 16005
rect 2720 16035 2760 16040
rect 2720 16005 2725 16035
rect 2755 16005 2760 16035
rect 2720 16000 2760 16005
rect 2800 16035 2840 16040
rect 2800 16005 2805 16035
rect 2835 16005 2840 16035
rect 2800 16000 2840 16005
rect 2880 16035 2920 16040
rect 2880 16005 2885 16035
rect 2915 16005 2920 16035
rect 2880 16000 2920 16005
rect 2960 16035 3000 16040
rect 2960 16005 2965 16035
rect 2995 16005 3000 16035
rect 2960 16000 3000 16005
rect 3040 16035 3080 16040
rect 3040 16005 3045 16035
rect 3075 16005 3080 16035
rect 3040 16000 3080 16005
rect 3120 16035 3160 16040
rect 3120 16005 3125 16035
rect 3155 16005 3160 16035
rect 3120 16000 3160 16005
rect 3200 16035 3240 16040
rect 3200 16005 3205 16035
rect 3235 16005 3240 16035
rect 3200 16000 3240 16005
rect 3280 16035 3320 16040
rect 3280 16005 3285 16035
rect 3315 16005 3320 16035
rect 3280 16000 3320 16005
rect 3360 16035 3400 16040
rect 3360 16005 3365 16035
rect 3395 16005 3400 16035
rect 3360 16000 3400 16005
rect 3440 16035 3480 16040
rect 3440 16005 3445 16035
rect 3475 16005 3480 16035
rect 3440 16000 3480 16005
rect 3520 16035 3560 16040
rect 3520 16005 3525 16035
rect 3555 16005 3560 16035
rect 3520 16000 3560 16005
rect 3600 16035 3640 16040
rect 3600 16005 3605 16035
rect 3635 16005 3640 16035
rect 3600 16000 3640 16005
rect 3680 16035 3720 16040
rect 3680 16005 3685 16035
rect 3715 16005 3720 16035
rect 3680 16000 3720 16005
rect 3760 16035 3800 16040
rect 3760 16005 3765 16035
rect 3795 16005 3800 16035
rect 3760 16000 3800 16005
rect 3840 16035 3880 16040
rect 3840 16005 3845 16035
rect 3875 16005 3880 16035
rect 3840 16000 3880 16005
rect 3920 16035 3960 16040
rect 3920 16005 3925 16035
rect 3955 16005 3960 16035
rect 3920 16000 3960 16005
rect 4000 16035 4040 16040
rect 4000 16005 4005 16035
rect 4035 16005 4040 16035
rect 4000 16000 4040 16005
rect 4080 16035 4120 16040
rect 4080 16005 4085 16035
rect 4115 16005 4120 16035
rect 4080 16000 4120 16005
rect 4160 16035 4200 16040
rect 4160 16005 4165 16035
rect 4195 16005 4200 16035
rect 4160 16000 4200 16005
rect 6240 16035 6280 16040
rect 6240 16005 6245 16035
rect 6275 16005 6280 16035
rect 6240 16000 6280 16005
rect 6320 16035 6360 16040
rect 6320 16005 6325 16035
rect 6355 16005 6360 16035
rect 6320 16000 6360 16005
rect 6400 16035 6440 16040
rect 6400 16005 6405 16035
rect 6435 16005 6440 16035
rect 6400 16000 6440 16005
rect 6480 16035 6520 16040
rect 6480 16005 6485 16035
rect 6515 16005 6520 16035
rect 6480 16000 6520 16005
rect 6560 16035 6600 16040
rect 6560 16005 6565 16035
rect 6595 16005 6600 16035
rect 6560 16000 6600 16005
rect 6640 16035 6680 16040
rect 6640 16005 6645 16035
rect 6675 16005 6680 16035
rect 6640 16000 6680 16005
rect 6720 16035 6760 16040
rect 6720 16005 6725 16035
rect 6755 16005 6760 16035
rect 6720 16000 6760 16005
rect 6800 16035 6840 16040
rect 6800 16005 6805 16035
rect 6835 16005 6840 16035
rect 6800 16000 6840 16005
rect 6880 16035 6920 16040
rect 6880 16005 6885 16035
rect 6915 16005 6920 16035
rect 6880 16000 6920 16005
rect 6960 16035 7000 16040
rect 6960 16005 6965 16035
rect 6995 16005 7000 16035
rect 6960 16000 7000 16005
rect 7040 16035 7080 16040
rect 7040 16005 7045 16035
rect 7075 16005 7080 16035
rect 7040 16000 7080 16005
rect 7120 16035 7160 16040
rect 7120 16005 7125 16035
rect 7155 16005 7160 16035
rect 7120 16000 7160 16005
rect 7200 16035 7240 16040
rect 7200 16005 7205 16035
rect 7235 16005 7240 16035
rect 7200 16000 7240 16005
rect 7280 16035 7320 16040
rect 7280 16005 7285 16035
rect 7315 16005 7320 16035
rect 7280 16000 7320 16005
rect 7360 16035 7400 16040
rect 7360 16005 7365 16035
rect 7395 16005 7400 16035
rect 7360 16000 7400 16005
rect 7440 16035 7480 16040
rect 7440 16005 7445 16035
rect 7475 16005 7480 16035
rect 7440 16000 7480 16005
rect 7520 16035 7560 16040
rect 7520 16005 7525 16035
rect 7555 16005 7560 16035
rect 7520 16000 7560 16005
rect 7600 16035 7640 16040
rect 7600 16005 7605 16035
rect 7635 16005 7640 16035
rect 7600 16000 7640 16005
rect 7680 16035 7720 16040
rect 7680 16005 7685 16035
rect 7715 16005 7720 16035
rect 7680 16000 7720 16005
rect 7760 16035 7800 16040
rect 7760 16005 7765 16035
rect 7795 16005 7800 16035
rect 7760 16000 7800 16005
rect 7840 16035 7880 16040
rect 7840 16005 7845 16035
rect 7875 16005 7880 16035
rect 7840 16000 7880 16005
rect 7920 16035 7960 16040
rect 7920 16005 7925 16035
rect 7955 16005 7960 16035
rect 7920 16000 7960 16005
rect 8000 16035 8040 16040
rect 8000 16005 8005 16035
rect 8035 16005 8040 16035
rect 8000 16000 8040 16005
rect 8080 16035 8120 16040
rect 8080 16005 8085 16035
rect 8115 16005 8120 16035
rect 8080 16000 8120 16005
rect 8160 16035 8200 16040
rect 8160 16005 8165 16035
rect 8195 16005 8200 16035
rect 8160 16000 8200 16005
rect 8240 16035 8280 16040
rect 8240 16005 8245 16035
rect 8275 16005 8280 16035
rect 8240 16000 8280 16005
rect 8320 16035 8360 16040
rect 8320 16005 8325 16035
rect 8355 16005 8360 16035
rect 8320 16000 8360 16005
rect 8400 16035 8440 16040
rect 8400 16005 8405 16035
rect 8435 16005 8440 16035
rect 8400 16000 8440 16005
rect 8480 16035 8520 16040
rect 8480 16005 8485 16035
rect 8515 16005 8520 16035
rect 8480 16000 8520 16005
rect 8560 16035 8600 16040
rect 8560 16005 8565 16035
rect 8595 16005 8600 16035
rect 8560 16000 8600 16005
rect 8640 16035 8680 16040
rect 8640 16005 8645 16035
rect 8675 16005 8680 16035
rect 8640 16000 8680 16005
rect 8720 16035 8760 16040
rect 8720 16005 8725 16035
rect 8755 16005 8760 16035
rect 8720 16000 8760 16005
rect 8800 16035 8840 16040
rect 8800 16005 8805 16035
rect 8835 16005 8840 16035
rect 8800 16000 8840 16005
rect 8880 16035 8920 16040
rect 8880 16005 8885 16035
rect 8915 16005 8920 16035
rect 8880 16000 8920 16005
rect 8960 16035 9000 16040
rect 8960 16005 8965 16035
rect 8995 16005 9000 16035
rect 8960 16000 9000 16005
rect 9040 16035 9080 16040
rect 9040 16005 9045 16035
rect 9075 16005 9080 16035
rect 9040 16000 9080 16005
rect 9120 16035 9160 16040
rect 9120 16005 9125 16035
rect 9155 16005 9160 16035
rect 9120 16000 9160 16005
rect 9200 16035 9240 16040
rect 9200 16005 9205 16035
rect 9235 16005 9240 16035
rect 9200 16000 9240 16005
rect 9280 16035 9320 16040
rect 9280 16005 9285 16035
rect 9315 16005 9320 16035
rect 9280 16000 9320 16005
rect 9360 16035 9400 16040
rect 9360 16005 9365 16035
rect 9395 16005 9400 16035
rect 9360 16000 9400 16005
rect 9440 16035 9480 16040
rect 9440 16005 9445 16035
rect 9475 16005 9480 16035
rect 9440 16000 9480 16005
rect 11560 16035 11600 16040
rect 11560 16005 11565 16035
rect 11595 16005 11600 16035
rect 11560 16000 11600 16005
rect 11640 16035 11680 16040
rect 11640 16005 11645 16035
rect 11675 16005 11680 16035
rect 11640 16000 11680 16005
rect 11720 16035 11760 16040
rect 11720 16005 11725 16035
rect 11755 16005 11760 16035
rect 11720 16000 11760 16005
rect 11800 16035 11840 16040
rect 11800 16005 11805 16035
rect 11835 16005 11840 16035
rect 11800 16000 11840 16005
rect 11880 16035 11920 16040
rect 11880 16005 11885 16035
rect 11915 16005 11920 16035
rect 11880 16000 11920 16005
rect 11960 16035 12000 16040
rect 11960 16005 11965 16035
rect 11995 16005 12000 16035
rect 11960 16000 12000 16005
rect 12040 16035 12080 16040
rect 12040 16005 12045 16035
rect 12075 16005 12080 16035
rect 12040 16000 12080 16005
rect 12120 16035 12160 16040
rect 12120 16005 12125 16035
rect 12155 16005 12160 16035
rect 12120 16000 12160 16005
rect 12200 16035 12240 16040
rect 12200 16005 12205 16035
rect 12235 16005 12240 16035
rect 12200 16000 12240 16005
rect 12280 16035 12320 16040
rect 12280 16005 12285 16035
rect 12315 16005 12320 16035
rect 12280 16000 12320 16005
rect 12360 16035 12400 16040
rect 12360 16005 12365 16035
rect 12395 16005 12400 16035
rect 12360 16000 12400 16005
rect 12440 16035 12480 16040
rect 12440 16005 12445 16035
rect 12475 16005 12480 16035
rect 12440 16000 12480 16005
rect 12520 16035 12560 16040
rect 12520 16005 12525 16035
rect 12555 16005 12560 16035
rect 12520 16000 12560 16005
rect 12600 16035 12640 16040
rect 12600 16005 12605 16035
rect 12635 16005 12640 16035
rect 12600 16000 12640 16005
rect 12680 16035 12720 16040
rect 12680 16005 12685 16035
rect 12715 16005 12720 16035
rect 12680 16000 12720 16005
rect 12760 16035 12800 16040
rect 12760 16005 12765 16035
rect 12795 16005 12800 16035
rect 12760 16000 12800 16005
rect 12840 16035 12880 16040
rect 12840 16005 12845 16035
rect 12875 16005 12880 16035
rect 12840 16000 12880 16005
rect 12920 16035 12960 16040
rect 12920 16005 12925 16035
rect 12955 16005 12960 16035
rect 12920 16000 12960 16005
rect 13000 16035 13040 16040
rect 13000 16005 13005 16035
rect 13035 16005 13040 16035
rect 13000 16000 13040 16005
rect 13080 16035 13120 16040
rect 13080 16005 13085 16035
rect 13115 16005 13120 16035
rect 13080 16000 13120 16005
rect 13160 16035 13200 16040
rect 13160 16005 13165 16035
rect 13195 16005 13200 16035
rect 13160 16000 13200 16005
rect 13240 16035 13280 16040
rect 13240 16005 13245 16035
rect 13275 16005 13280 16035
rect 13240 16000 13280 16005
rect 13320 16035 13360 16040
rect 13320 16005 13325 16035
rect 13355 16005 13360 16035
rect 13320 16000 13360 16005
rect 13400 16035 13440 16040
rect 13400 16005 13405 16035
rect 13435 16005 13440 16035
rect 13400 16000 13440 16005
rect 13480 16035 13520 16040
rect 13480 16005 13485 16035
rect 13515 16005 13520 16035
rect 13480 16000 13520 16005
rect 13560 16035 13600 16040
rect 13560 16005 13565 16035
rect 13595 16005 13600 16035
rect 13560 16000 13600 16005
rect 13640 16035 13680 16040
rect 13640 16005 13645 16035
rect 13675 16005 13680 16035
rect 13640 16000 13680 16005
rect 13720 16035 13760 16040
rect 13720 16005 13725 16035
rect 13755 16005 13760 16035
rect 13720 16000 13760 16005
rect 13800 16035 13840 16040
rect 13800 16005 13805 16035
rect 13835 16005 13840 16035
rect 13800 16000 13840 16005
rect 13880 16035 13920 16040
rect 13880 16005 13885 16035
rect 13915 16005 13920 16035
rect 13880 16000 13920 16005
rect 13960 16035 14000 16040
rect 13960 16005 13965 16035
rect 13995 16005 14000 16035
rect 13960 16000 14000 16005
rect 14040 16035 14080 16040
rect 14040 16005 14045 16035
rect 14075 16005 14080 16035
rect 14040 16000 14080 16005
rect 14120 16035 14160 16040
rect 14120 16005 14125 16035
rect 14155 16005 14160 16035
rect 14120 16000 14160 16005
rect 14200 16035 14240 16040
rect 14200 16005 14205 16035
rect 14235 16005 14240 16035
rect 14200 16000 14240 16005
rect 14280 16035 14320 16040
rect 14280 16005 14285 16035
rect 14315 16005 14320 16035
rect 14280 16000 14320 16005
rect 14360 16035 14400 16040
rect 14360 16005 14365 16035
rect 14395 16005 14400 16035
rect 14360 16000 14400 16005
rect 14440 16035 14480 16040
rect 14440 16005 14445 16035
rect 14475 16005 14480 16035
rect 14440 16000 14480 16005
rect 14520 16035 14560 16040
rect 14520 16005 14525 16035
rect 14555 16005 14560 16035
rect 14520 16000 14560 16005
rect 14600 16035 14640 16040
rect 14600 16005 14605 16035
rect 14635 16005 14640 16035
rect 14600 16000 14640 16005
rect 14680 16035 14720 16040
rect 14680 16005 14685 16035
rect 14715 16005 14720 16035
rect 14680 16000 14720 16005
rect 16760 16035 16800 16040
rect 16760 16005 16765 16035
rect 16795 16005 16800 16035
rect 16760 16000 16800 16005
rect 16840 16035 16880 16040
rect 16840 16005 16845 16035
rect 16875 16005 16880 16035
rect 16840 16000 16880 16005
rect 16920 16035 16960 16040
rect 16920 16005 16925 16035
rect 16955 16005 16960 16035
rect 16920 16000 16960 16005
rect 17000 16035 17040 16040
rect 17000 16005 17005 16035
rect 17035 16005 17040 16035
rect 17000 16000 17040 16005
rect 17080 16035 17120 16040
rect 17080 16005 17085 16035
rect 17115 16005 17120 16035
rect 17080 16000 17120 16005
rect 17160 16035 17200 16040
rect 17160 16005 17165 16035
rect 17195 16005 17200 16035
rect 17160 16000 17200 16005
rect 17240 16035 17280 16040
rect 17240 16005 17245 16035
rect 17275 16005 17280 16035
rect 17240 16000 17280 16005
rect 17320 16035 17360 16040
rect 17320 16005 17325 16035
rect 17355 16005 17360 16035
rect 17320 16000 17360 16005
rect 17400 16035 17440 16040
rect 17400 16005 17405 16035
rect 17435 16005 17440 16035
rect 17400 16000 17440 16005
rect 17480 16035 17520 16040
rect 17480 16005 17485 16035
rect 17515 16005 17520 16035
rect 17480 16000 17520 16005
rect 17560 16035 17600 16040
rect 17560 16005 17565 16035
rect 17595 16005 17600 16035
rect 17560 16000 17600 16005
rect 17640 16035 17680 16040
rect 17640 16005 17645 16035
rect 17675 16005 17680 16035
rect 17640 16000 17680 16005
rect 17720 16035 17760 16040
rect 17720 16005 17725 16035
rect 17755 16005 17760 16035
rect 17720 16000 17760 16005
rect 17800 16035 17840 16040
rect 17800 16005 17805 16035
rect 17835 16005 17840 16035
rect 17800 16000 17840 16005
rect 17880 16035 17920 16040
rect 17880 16005 17885 16035
rect 17915 16005 17920 16035
rect 17880 16000 17920 16005
rect 17960 16035 18000 16040
rect 17960 16005 17965 16035
rect 17995 16005 18000 16035
rect 17960 16000 18000 16005
rect 18040 16035 18080 16040
rect 18040 16005 18045 16035
rect 18075 16005 18080 16035
rect 18040 16000 18080 16005
rect 18120 16035 18160 16040
rect 18120 16005 18125 16035
rect 18155 16005 18160 16035
rect 18120 16000 18160 16005
rect 18200 16035 18240 16040
rect 18200 16005 18205 16035
rect 18235 16005 18240 16035
rect 18200 16000 18240 16005
rect 18280 16035 18320 16040
rect 18280 16005 18285 16035
rect 18315 16005 18320 16035
rect 18280 16000 18320 16005
rect 18360 16035 18400 16040
rect 18360 16005 18365 16035
rect 18395 16005 18400 16035
rect 18360 16000 18400 16005
rect 18440 16035 18480 16040
rect 18440 16005 18445 16035
rect 18475 16005 18480 16035
rect 18440 16000 18480 16005
rect 18520 16035 18560 16040
rect 18520 16005 18525 16035
rect 18555 16005 18560 16035
rect 18520 16000 18560 16005
rect 18600 16035 18640 16040
rect 18600 16005 18605 16035
rect 18635 16005 18640 16035
rect 18600 16000 18640 16005
rect 18680 16035 18720 16040
rect 18680 16005 18685 16035
rect 18715 16005 18720 16035
rect 18680 16000 18720 16005
rect 18760 16035 18800 16040
rect 18760 16005 18765 16035
rect 18795 16005 18800 16035
rect 18760 16000 18800 16005
rect 18840 16035 18880 16040
rect 18840 16005 18845 16035
rect 18875 16005 18880 16035
rect 18840 16000 18880 16005
rect 18920 16035 18960 16040
rect 18920 16005 18925 16035
rect 18955 16005 18960 16035
rect 18920 16000 18960 16005
rect 19000 16035 19040 16040
rect 19000 16005 19005 16035
rect 19035 16005 19040 16035
rect 19000 16000 19040 16005
rect 19080 16035 19120 16040
rect 19080 16005 19085 16035
rect 19115 16005 19120 16035
rect 19080 16000 19120 16005
rect 19160 16035 19200 16040
rect 19160 16005 19165 16035
rect 19195 16005 19200 16035
rect 19160 16000 19200 16005
rect 19240 16035 19280 16040
rect 19240 16005 19245 16035
rect 19275 16005 19280 16035
rect 19240 16000 19280 16005
rect 19320 16035 19360 16040
rect 19320 16005 19325 16035
rect 19355 16005 19360 16035
rect 19320 16000 19360 16005
rect 19400 16035 19440 16040
rect 19400 16005 19405 16035
rect 19435 16005 19440 16035
rect 19400 16000 19440 16005
rect 19480 16035 19520 16040
rect 19480 16005 19485 16035
rect 19515 16005 19520 16035
rect 19480 16000 19520 16005
rect 19560 16035 19600 16040
rect 19560 16005 19565 16035
rect 19595 16005 19600 16035
rect 19560 16000 19600 16005
rect 19640 16035 19680 16040
rect 19640 16005 19645 16035
rect 19675 16005 19680 16035
rect 19640 16000 19680 16005
rect 19720 16035 19760 16040
rect 19720 16005 19725 16035
rect 19755 16005 19760 16035
rect 19720 16000 19760 16005
rect 19800 16035 19840 16040
rect 19800 16005 19805 16035
rect 19835 16005 19840 16035
rect 19800 16000 19840 16005
rect 19880 16035 19920 16040
rect 19880 16005 19885 16035
rect 19915 16005 19920 16035
rect 19880 16000 19920 16005
rect 19960 16035 20000 16040
rect 19960 16005 19965 16035
rect 19995 16005 20000 16035
rect 19960 16000 20000 16005
rect 20040 16035 20080 16040
rect 20040 16005 20045 16035
rect 20075 16005 20080 16035
rect 20040 16000 20080 16005
rect 20120 16035 20160 16040
rect 20120 16005 20125 16035
rect 20155 16005 20160 16035
rect 20120 16000 20160 16005
rect 20200 16035 20240 16040
rect 20200 16005 20205 16035
rect 20235 16005 20240 16035
rect 20200 16000 20240 16005
rect 20280 16035 20320 16040
rect 20280 16005 20285 16035
rect 20315 16005 20320 16035
rect 20280 16000 20320 16005
rect 20360 16035 20400 16040
rect 20360 16005 20365 16035
rect 20395 16005 20400 16035
rect 20360 16000 20400 16005
rect 20440 16035 20480 16040
rect 20440 16005 20445 16035
rect 20475 16005 20480 16035
rect 20440 16000 20480 16005
rect 20520 16035 20560 16040
rect 20520 16005 20525 16035
rect 20555 16005 20560 16035
rect 20520 16000 20560 16005
rect 20600 16035 20640 16040
rect 20600 16005 20605 16035
rect 20635 16005 20640 16035
rect 20600 16000 20640 16005
rect 20680 16035 20720 16040
rect 20680 16005 20685 16035
rect 20715 16005 20720 16035
rect 20680 16000 20720 16005
rect 20760 16035 20800 16040
rect 20760 16005 20765 16035
rect 20795 16005 20800 16035
rect 20760 16000 20800 16005
rect 20840 16035 20880 16040
rect 20840 16005 20845 16035
rect 20875 16005 20880 16035
rect 20840 16000 20880 16005
rect 20920 16035 20960 16040
rect 20920 16005 20925 16035
rect 20955 16005 20960 16035
rect 20920 16000 20960 16005
rect 0 15875 40 15880
rect 0 15845 5 15875
rect 35 15845 40 15875
rect 0 15840 40 15845
rect 80 15875 120 15880
rect 80 15845 85 15875
rect 115 15845 120 15875
rect 80 15840 120 15845
rect 160 15875 200 15880
rect 160 15845 165 15875
rect 195 15845 200 15875
rect 160 15840 200 15845
rect 240 15875 280 15880
rect 240 15845 245 15875
rect 275 15845 280 15875
rect 240 15840 280 15845
rect 320 15875 360 15880
rect 320 15845 325 15875
rect 355 15845 360 15875
rect 320 15840 360 15845
rect 400 15875 440 15880
rect 400 15845 405 15875
rect 435 15845 440 15875
rect 400 15840 440 15845
rect 480 15875 520 15880
rect 480 15845 485 15875
rect 515 15845 520 15875
rect 480 15840 520 15845
rect 560 15875 600 15880
rect 560 15845 565 15875
rect 595 15845 600 15875
rect 560 15840 600 15845
rect 640 15875 680 15880
rect 640 15845 645 15875
rect 675 15845 680 15875
rect 640 15840 680 15845
rect 720 15875 760 15880
rect 720 15845 725 15875
rect 755 15845 760 15875
rect 720 15840 760 15845
rect 800 15875 840 15880
rect 800 15845 805 15875
rect 835 15845 840 15875
rect 800 15840 840 15845
rect 880 15875 920 15880
rect 880 15845 885 15875
rect 915 15845 920 15875
rect 880 15840 920 15845
rect 960 15875 1000 15880
rect 960 15845 965 15875
rect 995 15845 1000 15875
rect 960 15840 1000 15845
rect 1040 15875 1080 15880
rect 1040 15845 1045 15875
rect 1075 15845 1080 15875
rect 1040 15840 1080 15845
rect 1120 15875 1160 15880
rect 1120 15845 1125 15875
rect 1155 15845 1160 15875
rect 1120 15840 1160 15845
rect 1200 15875 1240 15880
rect 1200 15845 1205 15875
rect 1235 15845 1240 15875
rect 1200 15840 1240 15845
rect 1280 15875 1320 15880
rect 1280 15845 1285 15875
rect 1315 15845 1320 15875
rect 1280 15840 1320 15845
rect 1360 15875 1400 15880
rect 1360 15845 1365 15875
rect 1395 15845 1400 15875
rect 1360 15840 1400 15845
rect 1440 15875 1480 15880
rect 1440 15845 1445 15875
rect 1475 15845 1480 15875
rect 1440 15840 1480 15845
rect 1520 15875 1560 15880
rect 1520 15845 1525 15875
rect 1555 15845 1560 15875
rect 1520 15840 1560 15845
rect 1600 15875 1640 15880
rect 1600 15845 1605 15875
rect 1635 15845 1640 15875
rect 1600 15840 1640 15845
rect 1680 15875 1720 15880
rect 1680 15845 1685 15875
rect 1715 15845 1720 15875
rect 1680 15840 1720 15845
rect 1760 15875 1800 15880
rect 1760 15845 1765 15875
rect 1795 15845 1800 15875
rect 1760 15840 1800 15845
rect 1840 15875 1880 15880
rect 1840 15845 1845 15875
rect 1875 15845 1880 15875
rect 1840 15840 1880 15845
rect 1920 15875 1960 15880
rect 1920 15845 1925 15875
rect 1955 15845 1960 15875
rect 1920 15840 1960 15845
rect 2000 15875 2040 15880
rect 2000 15845 2005 15875
rect 2035 15845 2040 15875
rect 2000 15840 2040 15845
rect 2080 15875 2120 15880
rect 2080 15845 2085 15875
rect 2115 15845 2120 15875
rect 2080 15840 2120 15845
rect 2160 15875 2200 15880
rect 2160 15845 2165 15875
rect 2195 15845 2200 15875
rect 2160 15840 2200 15845
rect 2240 15875 2280 15880
rect 2240 15845 2245 15875
rect 2275 15845 2280 15875
rect 2240 15840 2280 15845
rect 2320 15875 2360 15880
rect 2320 15845 2325 15875
rect 2355 15845 2360 15875
rect 2320 15840 2360 15845
rect 2400 15875 2440 15880
rect 2400 15845 2405 15875
rect 2435 15845 2440 15875
rect 2400 15840 2440 15845
rect 2480 15875 2520 15880
rect 2480 15845 2485 15875
rect 2515 15845 2520 15875
rect 2480 15840 2520 15845
rect 2560 15875 2600 15880
rect 2560 15845 2565 15875
rect 2595 15845 2600 15875
rect 2560 15840 2600 15845
rect 2640 15875 2680 15880
rect 2640 15845 2645 15875
rect 2675 15845 2680 15875
rect 2640 15840 2680 15845
rect 2720 15875 2760 15880
rect 2720 15845 2725 15875
rect 2755 15845 2760 15875
rect 2720 15840 2760 15845
rect 2800 15875 2840 15880
rect 2800 15845 2805 15875
rect 2835 15845 2840 15875
rect 2800 15840 2840 15845
rect 2880 15875 2920 15880
rect 2880 15845 2885 15875
rect 2915 15845 2920 15875
rect 2880 15840 2920 15845
rect 2960 15875 3000 15880
rect 2960 15845 2965 15875
rect 2995 15845 3000 15875
rect 2960 15840 3000 15845
rect 3040 15875 3080 15880
rect 3040 15845 3045 15875
rect 3075 15845 3080 15875
rect 3040 15840 3080 15845
rect 3120 15875 3160 15880
rect 3120 15845 3125 15875
rect 3155 15845 3160 15875
rect 3120 15840 3160 15845
rect 3200 15875 3240 15880
rect 3200 15845 3205 15875
rect 3235 15845 3240 15875
rect 3200 15840 3240 15845
rect 3280 15875 3320 15880
rect 3280 15845 3285 15875
rect 3315 15845 3320 15875
rect 3280 15840 3320 15845
rect 3360 15875 3400 15880
rect 3360 15845 3365 15875
rect 3395 15845 3400 15875
rect 3360 15840 3400 15845
rect 3440 15875 3480 15880
rect 3440 15845 3445 15875
rect 3475 15845 3480 15875
rect 3440 15840 3480 15845
rect 3520 15875 3560 15880
rect 3520 15845 3525 15875
rect 3555 15845 3560 15875
rect 3520 15840 3560 15845
rect 3600 15875 3640 15880
rect 3600 15845 3605 15875
rect 3635 15845 3640 15875
rect 3600 15840 3640 15845
rect 3680 15875 3720 15880
rect 3680 15845 3685 15875
rect 3715 15845 3720 15875
rect 3680 15840 3720 15845
rect 3760 15875 3800 15880
rect 3760 15845 3765 15875
rect 3795 15845 3800 15875
rect 3760 15840 3800 15845
rect 3840 15875 3880 15880
rect 3840 15845 3845 15875
rect 3875 15845 3880 15875
rect 3840 15840 3880 15845
rect 3920 15875 3960 15880
rect 3920 15845 3925 15875
rect 3955 15845 3960 15875
rect 3920 15840 3960 15845
rect 4000 15875 4040 15880
rect 4000 15845 4005 15875
rect 4035 15845 4040 15875
rect 4000 15840 4040 15845
rect 4080 15875 4120 15880
rect 4080 15845 4085 15875
rect 4115 15845 4120 15875
rect 4080 15840 4120 15845
rect 4160 15875 4200 15880
rect 4160 15845 4165 15875
rect 4195 15845 4200 15875
rect 4160 15840 4200 15845
rect 6240 15875 6280 15880
rect 6240 15845 6245 15875
rect 6275 15845 6280 15875
rect 6240 15840 6280 15845
rect 6320 15875 6360 15880
rect 6320 15845 6325 15875
rect 6355 15845 6360 15875
rect 6320 15840 6360 15845
rect 6400 15875 6440 15880
rect 6400 15845 6405 15875
rect 6435 15845 6440 15875
rect 6400 15840 6440 15845
rect 6480 15875 6520 15880
rect 6480 15845 6485 15875
rect 6515 15845 6520 15875
rect 6480 15840 6520 15845
rect 6560 15875 6600 15880
rect 6560 15845 6565 15875
rect 6595 15845 6600 15875
rect 6560 15840 6600 15845
rect 6640 15875 6680 15880
rect 6640 15845 6645 15875
rect 6675 15845 6680 15875
rect 6640 15840 6680 15845
rect 6720 15875 6760 15880
rect 6720 15845 6725 15875
rect 6755 15845 6760 15875
rect 6720 15840 6760 15845
rect 6800 15875 6840 15880
rect 6800 15845 6805 15875
rect 6835 15845 6840 15875
rect 6800 15840 6840 15845
rect 6880 15875 6920 15880
rect 6880 15845 6885 15875
rect 6915 15845 6920 15875
rect 6880 15840 6920 15845
rect 6960 15875 7000 15880
rect 6960 15845 6965 15875
rect 6995 15845 7000 15875
rect 6960 15840 7000 15845
rect 7040 15875 7080 15880
rect 7040 15845 7045 15875
rect 7075 15845 7080 15875
rect 7040 15840 7080 15845
rect 7120 15875 7160 15880
rect 7120 15845 7125 15875
rect 7155 15845 7160 15875
rect 7120 15840 7160 15845
rect 7200 15875 7240 15880
rect 7200 15845 7205 15875
rect 7235 15845 7240 15875
rect 7200 15840 7240 15845
rect 7280 15875 7320 15880
rect 7280 15845 7285 15875
rect 7315 15845 7320 15875
rect 7280 15840 7320 15845
rect 7360 15875 7400 15880
rect 7360 15845 7365 15875
rect 7395 15845 7400 15875
rect 7360 15840 7400 15845
rect 7440 15875 7480 15880
rect 7440 15845 7445 15875
rect 7475 15845 7480 15875
rect 7440 15840 7480 15845
rect 7520 15875 7560 15880
rect 7520 15845 7525 15875
rect 7555 15845 7560 15875
rect 7520 15840 7560 15845
rect 7600 15875 7640 15880
rect 7600 15845 7605 15875
rect 7635 15845 7640 15875
rect 7600 15840 7640 15845
rect 7680 15875 7720 15880
rect 7680 15845 7685 15875
rect 7715 15845 7720 15875
rect 7680 15840 7720 15845
rect 7760 15875 7800 15880
rect 7760 15845 7765 15875
rect 7795 15845 7800 15875
rect 7760 15840 7800 15845
rect 7840 15875 7880 15880
rect 7840 15845 7845 15875
rect 7875 15845 7880 15875
rect 7840 15840 7880 15845
rect 7920 15875 7960 15880
rect 7920 15845 7925 15875
rect 7955 15845 7960 15875
rect 7920 15840 7960 15845
rect 8000 15875 8040 15880
rect 8000 15845 8005 15875
rect 8035 15845 8040 15875
rect 8000 15840 8040 15845
rect 8080 15875 8120 15880
rect 8080 15845 8085 15875
rect 8115 15845 8120 15875
rect 8080 15840 8120 15845
rect 8160 15875 8200 15880
rect 8160 15845 8165 15875
rect 8195 15845 8200 15875
rect 8160 15840 8200 15845
rect 8240 15875 8280 15880
rect 8240 15845 8245 15875
rect 8275 15845 8280 15875
rect 8240 15840 8280 15845
rect 8320 15875 8360 15880
rect 8320 15845 8325 15875
rect 8355 15845 8360 15875
rect 8320 15840 8360 15845
rect 8400 15875 8440 15880
rect 8400 15845 8405 15875
rect 8435 15845 8440 15875
rect 8400 15840 8440 15845
rect 8480 15875 8520 15880
rect 8480 15845 8485 15875
rect 8515 15845 8520 15875
rect 8480 15840 8520 15845
rect 8560 15875 8600 15880
rect 8560 15845 8565 15875
rect 8595 15845 8600 15875
rect 8560 15840 8600 15845
rect 8640 15875 8680 15880
rect 8640 15845 8645 15875
rect 8675 15845 8680 15875
rect 8640 15840 8680 15845
rect 8720 15875 8760 15880
rect 8720 15845 8725 15875
rect 8755 15845 8760 15875
rect 8720 15840 8760 15845
rect 8800 15875 8840 15880
rect 8800 15845 8805 15875
rect 8835 15845 8840 15875
rect 8800 15840 8840 15845
rect 8880 15875 8920 15880
rect 8880 15845 8885 15875
rect 8915 15845 8920 15875
rect 8880 15840 8920 15845
rect 8960 15875 9000 15880
rect 8960 15845 8965 15875
rect 8995 15845 9000 15875
rect 8960 15840 9000 15845
rect 9040 15875 9080 15880
rect 9040 15845 9045 15875
rect 9075 15845 9080 15875
rect 9040 15840 9080 15845
rect 9120 15875 9160 15880
rect 9120 15845 9125 15875
rect 9155 15845 9160 15875
rect 9120 15840 9160 15845
rect 9200 15875 9240 15880
rect 9200 15845 9205 15875
rect 9235 15845 9240 15875
rect 9200 15840 9240 15845
rect 9280 15875 9320 15880
rect 9280 15845 9285 15875
rect 9315 15845 9320 15875
rect 9280 15840 9320 15845
rect 9360 15875 9400 15880
rect 9360 15845 9365 15875
rect 9395 15845 9400 15875
rect 9360 15840 9400 15845
rect 9440 15875 9480 15880
rect 9440 15845 9445 15875
rect 9475 15845 9480 15875
rect 9440 15840 9480 15845
rect 11560 15875 11600 15880
rect 11560 15845 11565 15875
rect 11595 15845 11600 15875
rect 11560 15840 11600 15845
rect 11640 15875 11680 15880
rect 11640 15845 11645 15875
rect 11675 15845 11680 15875
rect 11640 15840 11680 15845
rect 11720 15875 11760 15880
rect 11720 15845 11725 15875
rect 11755 15845 11760 15875
rect 11720 15840 11760 15845
rect 11800 15875 11840 15880
rect 11800 15845 11805 15875
rect 11835 15845 11840 15875
rect 11800 15840 11840 15845
rect 11880 15875 11920 15880
rect 11880 15845 11885 15875
rect 11915 15845 11920 15875
rect 11880 15840 11920 15845
rect 11960 15875 12000 15880
rect 11960 15845 11965 15875
rect 11995 15845 12000 15875
rect 11960 15840 12000 15845
rect 12040 15875 12080 15880
rect 12040 15845 12045 15875
rect 12075 15845 12080 15875
rect 12040 15840 12080 15845
rect 12120 15875 12160 15880
rect 12120 15845 12125 15875
rect 12155 15845 12160 15875
rect 12120 15840 12160 15845
rect 12200 15875 12240 15880
rect 12200 15845 12205 15875
rect 12235 15845 12240 15875
rect 12200 15840 12240 15845
rect 12280 15875 12320 15880
rect 12280 15845 12285 15875
rect 12315 15845 12320 15875
rect 12280 15840 12320 15845
rect 12360 15875 12400 15880
rect 12360 15845 12365 15875
rect 12395 15845 12400 15875
rect 12360 15840 12400 15845
rect 12440 15875 12480 15880
rect 12440 15845 12445 15875
rect 12475 15845 12480 15875
rect 12440 15840 12480 15845
rect 12520 15875 12560 15880
rect 12520 15845 12525 15875
rect 12555 15845 12560 15875
rect 12520 15840 12560 15845
rect 12600 15875 12640 15880
rect 12600 15845 12605 15875
rect 12635 15845 12640 15875
rect 12600 15840 12640 15845
rect 12680 15875 12720 15880
rect 12680 15845 12685 15875
rect 12715 15845 12720 15875
rect 12680 15840 12720 15845
rect 12760 15875 12800 15880
rect 12760 15845 12765 15875
rect 12795 15845 12800 15875
rect 12760 15840 12800 15845
rect 12840 15875 12880 15880
rect 12840 15845 12845 15875
rect 12875 15845 12880 15875
rect 12840 15840 12880 15845
rect 12920 15875 12960 15880
rect 12920 15845 12925 15875
rect 12955 15845 12960 15875
rect 12920 15840 12960 15845
rect 13000 15875 13040 15880
rect 13000 15845 13005 15875
rect 13035 15845 13040 15875
rect 13000 15840 13040 15845
rect 13080 15875 13120 15880
rect 13080 15845 13085 15875
rect 13115 15845 13120 15875
rect 13080 15840 13120 15845
rect 13160 15875 13200 15880
rect 13160 15845 13165 15875
rect 13195 15845 13200 15875
rect 13160 15840 13200 15845
rect 13240 15875 13280 15880
rect 13240 15845 13245 15875
rect 13275 15845 13280 15875
rect 13240 15840 13280 15845
rect 13320 15875 13360 15880
rect 13320 15845 13325 15875
rect 13355 15845 13360 15875
rect 13320 15840 13360 15845
rect 13400 15875 13440 15880
rect 13400 15845 13405 15875
rect 13435 15845 13440 15875
rect 13400 15840 13440 15845
rect 13480 15875 13520 15880
rect 13480 15845 13485 15875
rect 13515 15845 13520 15875
rect 13480 15840 13520 15845
rect 13560 15875 13600 15880
rect 13560 15845 13565 15875
rect 13595 15845 13600 15875
rect 13560 15840 13600 15845
rect 13640 15875 13680 15880
rect 13640 15845 13645 15875
rect 13675 15845 13680 15875
rect 13640 15840 13680 15845
rect 13720 15875 13760 15880
rect 13720 15845 13725 15875
rect 13755 15845 13760 15875
rect 13720 15840 13760 15845
rect 13800 15875 13840 15880
rect 13800 15845 13805 15875
rect 13835 15845 13840 15875
rect 13800 15840 13840 15845
rect 13880 15875 13920 15880
rect 13880 15845 13885 15875
rect 13915 15845 13920 15875
rect 13880 15840 13920 15845
rect 13960 15875 14000 15880
rect 13960 15845 13965 15875
rect 13995 15845 14000 15875
rect 13960 15840 14000 15845
rect 14040 15875 14080 15880
rect 14040 15845 14045 15875
rect 14075 15845 14080 15875
rect 14040 15840 14080 15845
rect 14120 15875 14160 15880
rect 14120 15845 14125 15875
rect 14155 15845 14160 15875
rect 14120 15840 14160 15845
rect 14200 15875 14240 15880
rect 14200 15845 14205 15875
rect 14235 15845 14240 15875
rect 14200 15840 14240 15845
rect 14280 15875 14320 15880
rect 14280 15845 14285 15875
rect 14315 15845 14320 15875
rect 14280 15840 14320 15845
rect 14360 15875 14400 15880
rect 14360 15845 14365 15875
rect 14395 15845 14400 15875
rect 14360 15840 14400 15845
rect 14440 15875 14480 15880
rect 14440 15845 14445 15875
rect 14475 15845 14480 15875
rect 14440 15840 14480 15845
rect 14520 15875 14560 15880
rect 14520 15845 14525 15875
rect 14555 15845 14560 15875
rect 14520 15840 14560 15845
rect 14600 15875 14640 15880
rect 14600 15845 14605 15875
rect 14635 15845 14640 15875
rect 14600 15840 14640 15845
rect 14680 15875 14720 15880
rect 14680 15845 14685 15875
rect 14715 15845 14720 15875
rect 14680 15840 14720 15845
rect 16760 15875 16800 15880
rect 16760 15845 16765 15875
rect 16795 15845 16800 15875
rect 16760 15840 16800 15845
rect 16840 15875 16880 15880
rect 16840 15845 16845 15875
rect 16875 15845 16880 15875
rect 16840 15840 16880 15845
rect 16920 15875 16960 15880
rect 16920 15845 16925 15875
rect 16955 15845 16960 15875
rect 16920 15840 16960 15845
rect 17000 15875 17040 15880
rect 17000 15845 17005 15875
rect 17035 15845 17040 15875
rect 17000 15840 17040 15845
rect 17080 15875 17120 15880
rect 17080 15845 17085 15875
rect 17115 15845 17120 15875
rect 17080 15840 17120 15845
rect 17160 15875 17200 15880
rect 17160 15845 17165 15875
rect 17195 15845 17200 15875
rect 17160 15840 17200 15845
rect 17240 15875 17280 15880
rect 17240 15845 17245 15875
rect 17275 15845 17280 15875
rect 17240 15840 17280 15845
rect 17320 15875 17360 15880
rect 17320 15845 17325 15875
rect 17355 15845 17360 15875
rect 17320 15840 17360 15845
rect 17400 15875 17440 15880
rect 17400 15845 17405 15875
rect 17435 15845 17440 15875
rect 17400 15840 17440 15845
rect 17480 15875 17520 15880
rect 17480 15845 17485 15875
rect 17515 15845 17520 15875
rect 17480 15840 17520 15845
rect 17560 15875 17600 15880
rect 17560 15845 17565 15875
rect 17595 15845 17600 15875
rect 17560 15840 17600 15845
rect 17640 15875 17680 15880
rect 17640 15845 17645 15875
rect 17675 15845 17680 15875
rect 17640 15840 17680 15845
rect 17720 15875 17760 15880
rect 17720 15845 17725 15875
rect 17755 15845 17760 15875
rect 17720 15840 17760 15845
rect 17800 15875 17840 15880
rect 17800 15845 17805 15875
rect 17835 15845 17840 15875
rect 17800 15840 17840 15845
rect 17880 15875 17920 15880
rect 17880 15845 17885 15875
rect 17915 15845 17920 15875
rect 17880 15840 17920 15845
rect 17960 15875 18000 15880
rect 17960 15845 17965 15875
rect 17995 15845 18000 15875
rect 17960 15840 18000 15845
rect 18040 15875 18080 15880
rect 18040 15845 18045 15875
rect 18075 15845 18080 15875
rect 18040 15840 18080 15845
rect 18120 15875 18160 15880
rect 18120 15845 18125 15875
rect 18155 15845 18160 15875
rect 18120 15840 18160 15845
rect 18200 15875 18240 15880
rect 18200 15845 18205 15875
rect 18235 15845 18240 15875
rect 18200 15840 18240 15845
rect 18280 15875 18320 15880
rect 18280 15845 18285 15875
rect 18315 15845 18320 15875
rect 18280 15840 18320 15845
rect 18360 15875 18400 15880
rect 18360 15845 18365 15875
rect 18395 15845 18400 15875
rect 18360 15840 18400 15845
rect 18440 15875 18480 15880
rect 18440 15845 18445 15875
rect 18475 15845 18480 15875
rect 18440 15840 18480 15845
rect 18520 15875 18560 15880
rect 18520 15845 18525 15875
rect 18555 15845 18560 15875
rect 18520 15840 18560 15845
rect 18600 15875 18640 15880
rect 18600 15845 18605 15875
rect 18635 15845 18640 15875
rect 18600 15840 18640 15845
rect 18680 15875 18720 15880
rect 18680 15845 18685 15875
rect 18715 15845 18720 15875
rect 18680 15840 18720 15845
rect 18760 15875 18800 15880
rect 18760 15845 18765 15875
rect 18795 15845 18800 15875
rect 18760 15840 18800 15845
rect 18840 15875 18880 15880
rect 18840 15845 18845 15875
rect 18875 15845 18880 15875
rect 18840 15840 18880 15845
rect 18920 15875 18960 15880
rect 18920 15845 18925 15875
rect 18955 15845 18960 15875
rect 18920 15840 18960 15845
rect 19000 15875 19040 15880
rect 19000 15845 19005 15875
rect 19035 15845 19040 15875
rect 19000 15840 19040 15845
rect 19080 15875 19120 15880
rect 19080 15845 19085 15875
rect 19115 15845 19120 15875
rect 19080 15840 19120 15845
rect 19160 15875 19200 15880
rect 19160 15845 19165 15875
rect 19195 15845 19200 15875
rect 19160 15840 19200 15845
rect 19240 15875 19280 15880
rect 19240 15845 19245 15875
rect 19275 15845 19280 15875
rect 19240 15840 19280 15845
rect 19320 15875 19360 15880
rect 19320 15845 19325 15875
rect 19355 15845 19360 15875
rect 19320 15840 19360 15845
rect 19400 15875 19440 15880
rect 19400 15845 19405 15875
rect 19435 15845 19440 15875
rect 19400 15840 19440 15845
rect 19480 15875 19520 15880
rect 19480 15845 19485 15875
rect 19515 15845 19520 15875
rect 19480 15840 19520 15845
rect 19560 15875 19600 15880
rect 19560 15845 19565 15875
rect 19595 15845 19600 15875
rect 19560 15840 19600 15845
rect 19640 15875 19680 15880
rect 19640 15845 19645 15875
rect 19675 15845 19680 15875
rect 19640 15840 19680 15845
rect 19720 15875 19760 15880
rect 19720 15845 19725 15875
rect 19755 15845 19760 15875
rect 19720 15840 19760 15845
rect 19800 15875 19840 15880
rect 19800 15845 19805 15875
rect 19835 15845 19840 15875
rect 19800 15840 19840 15845
rect 19880 15875 19920 15880
rect 19880 15845 19885 15875
rect 19915 15845 19920 15875
rect 19880 15840 19920 15845
rect 19960 15875 20000 15880
rect 19960 15845 19965 15875
rect 19995 15845 20000 15875
rect 19960 15840 20000 15845
rect 20040 15875 20080 15880
rect 20040 15845 20045 15875
rect 20075 15845 20080 15875
rect 20040 15840 20080 15845
rect 20120 15875 20160 15880
rect 20120 15845 20125 15875
rect 20155 15845 20160 15875
rect 20120 15840 20160 15845
rect 20200 15875 20240 15880
rect 20200 15845 20205 15875
rect 20235 15845 20240 15875
rect 20200 15840 20240 15845
rect 20280 15875 20320 15880
rect 20280 15845 20285 15875
rect 20315 15845 20320 15875
rect 20280 15840 20320 15845
rect 20360 15875 20400 15880
rect 20360 15845 20365 15875
rect 20395 15845 20400 15875
rect 20360 15840 20400 15845
rect 20440 15875 20480 15880
rect 20440 15845 20445 15875
rect 20475 15845 20480 15875
rect 20440 15840 20480 15845
rect 20520 15875 20560 15880
rect 20520 15845 20525 15875
rect 20555 15845 20560 15875
rect 20520 15840 20560 15845
rect 20600 15875 20640 15880
rect 20600 15845 20605 15875
rect 20635 15845 20640 15875
rect 20600 15840 20640 15845
rect 20680 15875 20720 15880
rect 20680 15845 20685 15875
rect 20715 15845 20720 15875
rect 20680 15840 20720 15845
rect 20760 15875 20800 15880
rect 20760 15845 20765 15875
rect 20795 15845 20800 15875
rect 20760 15840 20800 15845
rect 20840 15875 20880 15880
rect 20840 15845 20845 15875
rect 20875 15845 20880 15875
rect 20840 15840 20880 15845
rect 20920 15875 20960 15880
rect 20920 15845 20925 15875
rect 20955 15845 20960 15875
rect 20920 15840 20960 15845
rect 0 15715 40 15720
rect 0 15685 5 15715
rect 35 15685 40 15715
rect 0 15680 40 15685
rect 80 15715 120 15720
rect 80 15685 85 15715
rect 115 15685 120 15715
rect 80 15680 120 15685
rect 160 15715 200 15720
rect 160 15685 165 15715
rect 195 15685 200 15715
rect 160 15680 200 15685
rect 240 15715 280 15720
rect 240 15685 245 15715
rect 275 15685 280 15715
rect 240 15680 280 15685
rect 320 15715 360 15720
rect 320 15685 325 15715
rect 355 15685 360 15715
rect 320 15680 360 15685
rect 400 15715 440 15720
rect 400 15685 405 15715
rect 435 15685 440 15715
rect 400 15680 440 15685
rect 480 15715 520 15720
rect 480 15685 485 15715
rect 515 15685 520 15715
rect 480 15680 520 15685
rect 560 15715 600 15720
rect 560 15685 565 15715
rect 595 15685 600 15715
rect 560 15680 600 15685
rect 640 15715 680 15720
rect 640 15685 645 15715
rect 675 15685 680 15715
rect 640 15680 680 15685
rect 720 15715 760 15720
rect 720 15685 725 15715
rect 755 15685 760 15715
rect 720 15680 760 15685
rect 800 15715 840 15720
rect 800 15685 805 15715
rect 835 15685 840 15715
rect 800 15680 840 15685
rect 880 15715 920 15720
rect 880 15685 885 15715
rect 915 15685 920 15715
rect 880 15680 920 15685
rect 960 15715 1000 15720
rect 960 15685 965 15715
rect 995 15685 1000 15715
rect 960 15680 1000 15685
rect 1040 15715 1080 15720
rect 1040 15685 1045 15715
rect 1075 15685 1080 15715
rect 1040 15680 1080 15685
rect 1120 15715 1160 15720
rect 1120 15685 1125 15715
rect 1155 15685 1160 15715
rect 1120 15680 1160 15685
rect 1200 15715 1240 15720
rect 1200 15685 1205 15715
rect 1235 15685 1240 15715
rect 1200 15680 1240 15685
rect 1280 15715 1320 15720
rect 1280 15685 1285 15715
rect 1315 15685 1320 15715
rect 1280 15680 1320 15685
rect 1360 15715 1400 15720
rect 1360 15685 1365 15715
rect 1395 15685 1400 15715
rect 1360 15680 1400 15685
rect 1440 15715 1480 15720
rect 1440 15685 1445 15715
rect 1475 15685 1480 15715
rect 1440 15680 1480 15685
rect 1520 15715 1560 15720
rect 1520 15685 1525 15715
rect 1555 15685 1560 15715
rect 1520 15680 1560 15685
rect 1600 15715 1640 15720
rect 1600 15685 1605 15715
rect 1635 15685 1640 15715
rect 1600 15680 1640 15685
rect 1680 15715 1720 15720
rect 1680 15685 1685 15715
rect 1715 15685 1720 15715
rect 1680 15680 1720 15685
rect 1760 15715 1800 15720
rect 1760 15685 1765 15715
rect 1795 15685 1800 15715
rect 1760 15680 1800 15685
rect 1840 15715 1880 15720
rect 1840 15685 1845 15715
rect 1875 15685 1880 15715
rect 1840 15680 1880 15685
rect 1920 15715 1960 15720
rect 1920 15685 1925 15715
rect 1955 15685 1960 15715
rect 1920 15680 1960 15685
rect 2000 15715 2040 15720
rect 2000 15685 2005 15715
rect 2035 15685 2040 15715
rect 2000 15680 2040 15685
rect 2080 15715 2120 15720
rect 2080 15685 2085 15715
rect 2115 15685 2120 15715
rect 2080 15680 2120 15685
rect 2160 15715 2200 15720
rect 2160 15685 2165 15715
rect 2195 15685 2200 15715
rect 2160 15680 2200 15685
rect 2240 15715 2280 15720
rect 2240 15685 2245 15715
rect 2275 15685 2280 15715
rect 2240 15680 2280 15685
rect 2320 15715 2360 15720
rect 2320 15685 2325 15715
rect 2355 15685 2360 15715
rect 2320 15680 2360 15685
rect 2400 15715 2440 15720
rect 2400 15685 2405 15715
rect 2435 15685 2440 15715
rect 2400 15680 2440 15685
rect 2480 15715 2520 15720
rect 2480 15685 2485 15715
rect 2515 15685 2520 15715
rect 2480 15680 2520 15685
rect 2560 15715 2600 15720
rect 2560 15685 2565 15715
rect 2595 15685 2600 15715
rect 2560 15680 2600 15685
rect 2640 15715 2680 15720
rect 2640 15685 2645 15715
rect 2675 15685 2680 15715
rect 2640 15680 2680 15685
rect 2720 15715 2760 15720
rect 2720 15685 2725 15715
rect 2755 15685 2760 15715
rect 2720 15680 2760 15685
rect 2800 15715 2840 15720
rect 2800 15685 2805 15715
rect 2835 15685 2840 15715
rect 2800 15680 2840 15685
rect 2880 15715 2920 15720
rect 2880 15685 2885 15715
rect 2915 15685 2920 15715
rect 2880 15680 2920 15685
rect 2960 15715 3000 15720
rect 2960 15685 2965 15715
rect 2995 15685 3000 15715
rect 2960 15680 3000 15685
rect 3040 15715 3080 15720
rect 3040 15685 3045 15715
rect 3075 15685 3080 15715
rect 3040 15680 3080 15685
rect 3120 15715 3160 15720
rect 3120 15685 3125 15715
rect 3155 15685 3160 15715
rect 3120 15680 3160 15685
rect 3200 15715 3240 15720
rect 3200 15685 3205 15715
rect 3235 15685 3240 15715
rect 3200 15680 3240 15685
rect 3280 15715 3320 15720
rect 3280 15685 3285 15715
rect 3315 15685 3320 15715
rect 3280 15680 3320 15685
rect 3360 15715 3400 15720
rect 3360 15685 3365 15715
rect 3395 15685 3400 15715
rect 3360 15680 3400 15685
rect 3440 15715 3480 15720
rect 3440 15685 3445 15715
rect 3475 15685 3480 15715
rect 3440 15680 3480 15685
rect 3520 15715 3560 15720
rect 3520 15685 3525 15715
rect 3555 15685 3560 15715
rect 3520 15680 3560 15685
rect 3600 15715 3640 15720
rect 3600 15685 3605 15715
rect 3635 15685 3640 15715
rect 3600 15680 3640 15685
rect 3680 15715 3720 15720
rect 3680 15685 3685 15715
rect 3715 15685 3720 15715
rect 3680 15680 3720 15685
rect 3760 15715 3800 15720
rect 3760 15685 3765 15715
rect 3795 15685 3800 15715
rect 3760 15680 3800 15685
rect 3840 15715 3880 15720
rect 3840 15685 3845 15715
rect 3875 15685 3880 15715
rect 3840 15680 3880 15685
rect 3920 15715 3960 15720
rect 3920 15685 3925 15715
rect 3955 15685 3960 15715
rect 3920 15680 3960 15685
rect 4000 15715 4040 15720
rect 4000 15685 4005 15715
rect 4035 15685 4040 15715
rect 4000 15680 4040 15685
rect 4080 15715 4120 15720
rect 4080 15685 4085 15715
rect 4115 15685 4120 15715
rect 4080 15680 4120 15685
rect 4160 15715 4200 15720
rect 4160 15685 4165 15715
rect 4195 15685 4200 15715
rect 4160 15680 4200 15685
rect 6240 15715 6280 15720
rect 6240 15685 6245 15715
rect 6275 15685 6280 15715
rect 6240 15680 6280 15685
rect 6320 15715 6360 15720
rect 6320 15685 6325 15715
rect 6355 15685 6360 15715
rect 6320 15680 6360 15685
rect 6400 15715 6440 15720
rect 6400 15685 6405 15715
rect 6435 15685 6440 15715
rect 6400 15680 6440 15685
rect 6480 15715 6520 15720
rect 6480 15685 6485 15715
rect 6515 15685 6520 15715
rect 6480 15680 6520 15685
rect 6560 15715 6600 15720
rect 6560 15685 6565 15715
rect 6595 15685 6600 15715
rect 6560 15680 6600 15685
rect 6640 15715 6680 15720
rect 6640 15685 6645 15715
rect 6675 15685 6680 15715
rect 6640 15680 6680 15685
rect 6720 15715 6760 15720
rect 6720 15685 6725 15715
rect 6755 15685 6760 15715
rect 6720 15680 6760 15685
rect 6800 15715 6840 15720
rect 6800 15685 6805 15715
rect 6835 15685 6840 15715
rect 6800 15680 6840 15685
rect 6880 15715 6920 15720
rect 6880 15685 6885 15715
rect 6915 15685 6920 15715
rect 6880 15680 6920 15685
rect 6960 15715 7000 15720
rect 6960 15685 6965 15715
rect 6995 15685 7000 15715
rect 6960 15680 7000 15685
rect 7040 15715 7080 15720
rect 7040 15685 7045 15715
rect 7075 15685 7080 15715
rect 7040 15680 7080 15685
rect 7120 15715 7160 15720
rect 7120 15685 7125 15715
rect 7155 15685 7160 15715
rect 7120 15680 7160 15685
rect 7200 15715 7240 15720
rect 7200 15685 7205 15715
rect 7235 15685 7240 15715
rect 7200 15680 7240 15685
rect 7280 15715 7320 15720
rect 7280 15685 7285 15715
rect 7315 15685 7320 15715
rect 7280 15680 7320 15685
rect 7360 15715 7400 15720
rect 7360 15685 7365 15715
rect 7395 15685 7400 15715
rect 7360 15680 7400 15685
rect 7440 15715 7480 15720
rect 7440 15685 7445 15715
rect 7475 15685 7480 15715
rect 7440 15680 7480 15685
rect 7520 15715 7560 15720
rect 7520 15685 7525 15715
rect 7555 15685 7560 15715
rect 7520 15680 7560 15685
rect 7600 15715 7640 15720
rect 7600 15685 7605 15715
rect 7635 15685 7640 15715
rect 7600 15680 7640 15685
rect 7680 15715 7720 15720
rect 7680 15685 7685 15715
rect 7715 15685 7720 15715
rect 7680 15680 7720 15685
rect 7760 15715 7800 15720
rect 7760 15685 7765 15715
rect 7795 15685 7800 15715
rect 7760 15680 7800 15685
rect 7840 15715 7880 15720
rect 7840 15685 7845 15715
rect 7875 15685 7880 15715
rect 7840 15680 7880 15685
rect 7920 15715 7960 15720
rect 7920 15685 7925 15715
rect 7955 15685 7960 15715
rect 7920 15680 7960 15685
rect 8000 15715 8040 15720
rect 8000 15685 8005 15715
rect 8035 15685 8040 15715
rect 8000 15680 8040 15685
rect 8080 15715 8120 15720
rect 8080 15685 8085 15715
rect 8115 15685 8120 15715
rect 8080 15680 8120 15685
rect 8160 15715 8200 15720
rect 8160 15685 8165 15715
rect 8195 15685 8200 15715
rect 8160 15680 8200 15685
rect 8240 15715 8280 15720
rect 8240 15685 8245 15715
rect 8275 15685 8280 15715
rect 8240 15680 8280 15685
rect 8320 15715 8360 15720
rect 8320 15685 8325 15715
rect 8355 15685 8360 15715
rect 8320 15680 8360 15685
rect 8400 15715 8440 15720
rect 8400 15685 8405 15715
rect 8435 15685 8440 15715
rect 8400 15680 8440 15685
rect 8480 15715 8520 15720
rect 8480 15685 8485 15715
rect 8515 15685 8520 15715
rect 8480 15680 8520 15685
rect 8560 15715 8600 15720
rect 8560 15685 8565 15715
rect 8595 15685 8600 15715
rect 8560 15680 8600 15685
rect 8640 15715 8680 15720
rect 8640 15685 8645 15715
rect 8675 15685 8680 15715
rect 8640 15680 8680 15685
rect 8720 15715 8760 15720
rect 8720 15685 8725 15715
rect 8755 15685 8760 15715
rect 8720 15680 8760 15685
rect 8800 15715 8840 15720
rect 8800 15685 8805 15715
rect 8835 15685 8840 15715
rect 8800 15680 8840 15685
rect 8880 15715 8920 15720
rect 8880 15685 8885 15715
rect 8915 15685 8920 15715
rect 8880 15680 8920 15685
rect 8960 15715 9000 15720
rect 8960 15685 8965 15715
rect 8995 15685 9000 15715
rect 8960 15680 9000 15685
rect 9040 15715 9080 15720
rect 9040 15685 9045 15715
rect 9075 15685 9080 15715
rect 9040 15680 9080 15685
rect 9120 15715 9160 15720
rect 9120 15685 9125 15715
rect 9155 15685 9160 15715
rect 9120 15680 9160 15685
rect 9200 15715 9240 15720
rect 9200 15685 9205 15715
rect 9235 15685 9240 15715
rect 9200 15680 9240 15685
rect 9280 15715 9320 15720
rect 9280 15685 9285 15715
rect 9315 15685 9320 15715
rect 9280 15680 9320 15685
rect 9360 15715 9400 15720
rect 9360 15685 9365 15715
rect 9395 15685 9400 15715
rect 9360 15680 9400 15685
rect 9440 15715 9480 15720
rect 9440 15685 9445 15715
rect 9475 15685 9480 15715
rect 9440 15680 9480 15685
rect 11560 15715 11600 15720
rect 11560 15685 11565 15715
rect 11595 15685 11600 15715
rect 11560 15680 11600 15685
rect 11640 15715 11680 15720
rect 11640 15685 11645 15715
rect 11675 15685 11680 15715
rect 11640 15680 11680 15685
rect 11720 15715 11760 15720
rect 11720 15685 11725 15715
rect 11755 15685 11760 15715
rect 11720 15680 11760 15685
rect 11800 15715 11840 15720
rect 11800 15685 11805 15715
rect 11835 15685 11840 15715
rect 11800 15680 11840 15685
rect 11880 15715 11920 15720
rect 11880 15685 11885 15715
rect 11915 15685 11920 15715
rect 11880 15680 11920 15685
rect 11960 15715 12000 15720
rect 11960 15685 11965 15715
rect 11995 15685 12000 15715
rect 11960 15680 12000 15685
rect 12040 15715 12080 15720
rect 12040 15685 12045 15715
rect 12075 15685 12080 15715
rect 12040 15680 12080 15685
rect 12120 15715 12160 15720
rect 12120 15685 12125 15715
rect 12155 15685 12160 15715
rect 12120 15680 12160 15685
rect 12200 15715 12240 15720
rect 12200 15685 12205 15715
rect 12235 15685 12240 15715
rect 12200 15680 12240 15685
rect 12280 15715 12320 15720
rect 12280 15685 12285 15715
rect 12315 15685 12320 15715
rect 12280 15680 12320 15685
rect 12360 15715 12400 15720
rect 12360 15685 12365 15715
rect 12395 15685 12400 15715
rect 12360 15680 12400 15685
rect 12440 15715 12480 15720
rect 12440 15685 12445 15715
rect 12475 15685 12480 15715
rect 12440 15680 12480 15685
rect 12520 15715 12560 15720
rect 12520 15685 12525 15715
rect 12555 15685 12560 15715
rect 12520 15680 12560 15685
rect 12600 15715 12640 15720
rect 12600 15685 12605 15715
rect 12635 15685 12640 15715
rect 12600 15680 12640 15685
rect 12680 15715 12720 15720
rect 12680 15685 12685 15715
rect 12715 15685 12720 15715
rect 12680 15680 12720 15685
rect 12760 15715 12800 15720
rect 12760 15685 12765 15715
rect 12795 15685 12800 15715
rect 12760 15680 12800 15685
rect 12840 15715 12880 15720
rect 12840 15685 12845 15715
rect 12875 15685 12880 15715
rect 12840 15680 12880 15685
rect 12920 15715 12960 15720
rect 12920 15685 12925 15715
rect 12955 15685 12960 15715
rect 12920 15680 12960 15685
rect 13000 15715 13040 15720
rect 13000 15685 13005 15715
rect 13035 15685 13040 15715
rect 13000 15680 13040 15685
rect 13080 15715 13120 15720
rect 13080 15685 13085 15715
rect 13115 15685 13120 15715
rect 13080 15680 13120 15685
rect 13160 15715 13200 15720
rect 13160 15685 13165 15715
rect 13195 15685 13200 15715
rect 13160 15680 13200 15685
rect 13240 15715 13280 15720
rect 13240 15685 13245 15715
rect 13275 15685 13280 15715
rect 13240 15680 13280 15685
rect 13320 15715 13360 15720
rect 13320 15685 13325 15715
rect 13355 15685 13360 15715
rect 13320 15680 13360 15685
rect 13400 15715 13440 15720
rect 13400 15685 13405 15715
rect 13435 15685 13440 15715
rect 13400 15680 13440 15685
rect 13480 15715 13520 15720
rect 13480 15685 13485 15715
rect 13515 15685 13520 15715
rect 13480 15680 13520 15685
rect 13560 15715 13600 15720
rect 13560 15685 13565 15715
rect 13595 15685 13600 15715
rect 13560 15680 13600 15685
rect 13640 15715 13680 15720
rect 13640 15685 13645 15715
rect 13675 15685 13680 15715
rect 13640 15680 13680 15685
rect 13720 15715 13760 15720
rect 13720 15685 13725 15715
rect 13755 15685 13760 15715
rect 13720 15680 13760 15685
rect 13800 15715 13840 15720
rect 13800 15685 13805 15715
rect 13835 15685 13840 15715
rect 13800 15680 13840 15685
rect 13880 15715 13920 15720
rect 13880 15685 13885 15715
rect 13915 15685 13920 15715
rect 13880 15680 13920 15685
rect 13960 15715 14000 15720
rect 13960 15685 13965 15715
rect 13995 15685 14000 15715
rect 13960 15680 14000 15685
rect 14040 15715 14080 15720
rect 14040 15685 14045 15715
rect 14075 15685 14080 15715
rect 14040 15680 14080 15685
rect 14120 15715 14160 15720
rect 14120 15685 14125 15715
rect 14155 15685 14160 15715
rect 14120 15680 14160 15685
rect 14200 15715 14240 15720
rect 14200 15685 14205 15715
rect 14235 15685 14240 15715
rect 14200 15680 14240 15685
rect 14280 15715 14320 15720
rect 14280 15685 14285 15715
rect 14315 15685 14320 15715
rect 14280 15680 14320 15685
rect 14360 15715 14400 15720
rect 14360 15685 14365 15715
rect 14395 15685 14400 15715
rect 14360 15680 14400 15685
rect 14440 15715 14480 15720
rect 14440 15685 14445 15715
rect 14475 15685 14480 15715
rect 14440 15680 14480 15685
rect 14520 15715 14560 15720
rect 14520 15685 14525 15715
rect 14555 15685 14560 15715
rect 14520 15680 14560 15685
rect 14600 15715 14640 15720
rect 14600 15685 14605 15715
rect 14635 15685 14640 15715
rect 14600 15680 14640 15685
rect 14680 15715 14720 15720
rect 14680 15685 14685 15715
rect 14715 15685 14720 15715
rect 14680 15680 14720 15685
rect 16760 15715 16800 15720
rect 16760 15685 16765 15715
rect 16795 15685 16800 15715
rect 16760 15680 16800 15685
rect 16840 15715 16880 15720
rect 16840 15685 16845 15715
rect 16875 15685 16880 15715
rect 16840 15680 16880 15685
rect 16920 15715 16960 15720
rect 16920 15685 16925 15715
rect 16955 15685 16960 15715
rect 16920 15680 16960 15685
rect 17000 15715 17040 15720
rect 17000 15685 17005 15715
rect 17035 15685 17040 15715
rect 17000 15680 17040 15685
rect 17080 15715 17120 15720
rect 17080 15685 17085 15715
rect 17115 15685 17120 15715
rect 17080 15680 17120 15685
rect 17160 15715 17200 15720
rect 17160 15685 17165 15715
rect 17195 15685 17200 15715
rect 17160 15680 17200 15685
rect 17240 15715 17280 15720
rect 17240 15685 17245 15715
rect 17275 15685 17280 15715
rect 17240 15680 17280 15685
rect 17320 15715 17360 15720
rect 17320 15685 17325 15715
rect 17355 15685 17360 15715
rect 17320 15680 17360 15685
rect 17400 15715 17440 15720
rect 17400 15685 17405 15715
rect 17435 15685 17440 15715
rect 17400 15680 17440 15685
rect 17480 15715 17520 15720
rect 17480 15685 17485 15715
rect 17515 15685 17520 15715
rect 17480 15680 17520 15685
rect 17560 15715 17600 15720
rect 17560 15685 17565 15715
rect 17595 15685 17600 15715
rect 17560 15680 17600 15685
rect 17640 15715 17680 15720
rect 17640 15685 17645 15715
rect 17675 15685 17680 15715
rect 17640 15680 17680 15685
rect 17720 15715 17760 15720
rect 17720 15685 17725 15715
rect 17755 15685 17760 15715
rect 17720 15680 17760 15685
rect 17800 15715 17840 15720
rect 17800 15685 17805 15715
rect 17835 15685 17840 15715
rect 17800 15680 17840 15685
rect 17880 15715 17920 15720
rect 17880 15685 17885 15715
rect 17915 15685 17920 15715
rect 17880 15680 17920 15685
rect 17960 15715 18000 15720
rect 17960 15685 17965 15715
rect 17995 15685 18000 15715
rect 17960 15680 18000 15685
rect 18040 15715 18080 15720
rect 18040 15685 18045 15715
rect 18075 15685 18080 15715
rect 18040 15680 18080 15685
rect 18120 15715 18160 15720
rect 18120 15685 18125 15715
rect 18155 15685 18160 15715
rect 18120 15680 18160 15685
rect 18200 15715 18240 15720
rect 18200 15685 18205 15715
rect 18235 15685 18240 15715
rect 18200 15680 18240 15685
rect 18280 15715 18320 15720
rect 18280 15685 18285 15715
rect 18315 15685 18320 15715
rect 18280 15680 18320 15685
rect 18360 15715 18400 15720
rect 18360 15685 18365 15715
rect 18395 15685 18400 15715
rect 18360 15680 18400 15685
rect 18440 15715 18480 15720
rect 18440 15685 18445 15715
rect 18475 15685 18480 15715
rect 18440 15680 18480 15685
rect 18520 15715 18560 15720
rect 18520 15685 18525 15715
rect 18555 15685 18560 15715
rect 18520 15680 18560 15685
rect 18600 15715 18640 15720
rect 18600 15685 18605 15715
rect 18635 15685 18640 15715
rect 18600 15680 18640 15685
rect 18680 15715 18720 15720
rect 18680 15685 18685 15715
rect 18715 15685 18720 15715
rect 18680 15680 18720 15685
rect 18760 15715 18800 15720
rect 18760 15685 18765 15715
rect 18795 15685 18800 15715
rect 18760 15680 18800 15685
rect 18840 15715 18880 15720
rect 18840 15685 18845 15715
rect 18875 15685 18880 15715
rect 18840 15680 18880 15685
rect 18920 15715 18960 15720
rect 18920 15685 18925 15715
rect 18955 15685 18960 15715
rect 18920 15680 18960 15685
rect 19000 15715 19040 15720
rect 19000 15685 19005 15715
rect 19035 15685 19040 15715
rect 19000 15680 19040 15685
rect 19080 15715 19120 15720
rect 19080 15685 19085 15715
rect 19115 15685 19120 15715
rect 19080 15680 19120 15685
rect 19160 15715 19200 15720
rect 19160 15685 19165 15715
rect 19195 15685 19200 15715
rect 19160 15680 19200 15685
rect 19240 15715 19280 15720
rect 19240 15685 19245 15715
rect 19275 15685 19280 15715
rect 19240 15680 19280 15685
rect 19320 15715 19360 15720
rect 19320 15685 19325 15715
rect 19355 15685 19360 15715
rect 19320 15680 19360 15685
rect 19400 15715 19440 15720
rect 19400 15685 19405 15715
rect 19435 15685 19440 15715
rect 19400 15680 19440 15685
rect 19480 15715 19520 15720
rect 19480 15685 19485 15715
rect 19515 15685 19520 15715
rect 19480 15680 19520 15685
rect 19560 15715 19600 15720
rect 19560 15685 19565 15715
rect 19595 15685 19600 15715
rect 19560 15680 19600 15685
rect 19640 15715 19680 15720
rect 19640 15685 19645 15715
rect 19675 15685 19680 15715
rect 19640 15680 19680 15685
rect 19720 15715 19760 15720
rect 19720 15685 19725 15715
rect 19755 15685 19760 15715
rect 19720 15680 19760 15685
rect 19800 15715 19840 15720
rect 19800 15685 19805 15715
rect 19835 15685 19840 15715
rect 19800 15680 19840 15685
rect 19880 15715 19920 15720
rect 19880 15685 19885 15715
rect 19915 15685 19920 15715
rect 19880 15680 19920 15685
rect 19960 15715 20000 15720
rect 19960 15685 19965 15715
rect 19995 15685 20000 15715
rect 19960 15680 20000 15685
rect 20040 15715 20080 15720
rect 20040 15685 20045 15715
rect 20075 15685 20080 15715
rect 20040 15680 20080 15685
rect 20120 15715 20160 15720
rect 20120 15685 20125 15715
rect 20155 15685 20160 15715
rect 20120 15680 20160 15685
rect 20200 15715 20240 15720
rect 20200 15685 20205 15715
rect 20235 15685 20240 15715
rect 20200 15680 20240 15685
rect 20280 15715 20320 15720
rect 20280 15685 20285 15715
rect 20315 15685 20320 15715
rect 20280 15680 20320 15685
rect 20360 15715 20400 15720
rect 20360 15685 20365 15715
rect 20395 15685 20400 15715
rect 20360 15680 20400 15685
rect 20440 15715 20480 15720
rect 20440 15685 20445 15715
rect 20475 15685 20480 15715
rect 20440 15680 20480 15685
rect 20520 15715 20560 15720
rect 20520 15685 20525 15715
rect 20555 15685 20560 15715
rect 20520 15680 20560 15685
rect 20600 15715 20640 15720
rect 20600 15685 20605 15715
rect 20635 15685 20640 15715
rect 20600 15680 20640 15685
rect 20680 15715 20720 15720
rect 20680 15685 20685 15715
rect 20715 15685 20720 15715
rect 20680 15680 20720 15685
rect 20760 15715 20800 15720
rect 20760 15685 20765 15715
rect 20795 15685 20800 15715
rect 20760 15680 20800 15685
rect 20840 15715 20880 15720
rect 20840 15685 20845 15715
rect 20875 15685 20880 15715
rect 20840 15680 20880 15685
rect 20920 15715 20960 15720
rect 20920 15685 20925 15715
rect 20955 15685 20960 15715
rect 20920 15680 20960 15685
rect 0 15555 40 15560
rect 0 15525 5 15555
rect 35 15525 40 15555
rect 0 15520 40 15525
rect 80 15555 120 15560
rect 80 15525 85 15555
rect 115 15525 120 15555
rect 80 15520 120 15525
rect 160 15555 200 15560
rect 160 15525 165 15555
rect 195 15525 200 15555
rect 160 15520 200 15525
rect 240 15555 280 15560
rect 240 15525 245 15555
rect 275 15525 280 15555
rect 240 15520 280 15525
rect 320 15555 360 15560
rect 320 15525 325 15555
rect 355 15525 360 15555
rect 320 15520 360 15525
rect 400 15555 440 15560
rect 400 15525 405 15555
rect 435 15525 440 15555
rect 400 15520 440 15525
rect 480 15555 520 15560
rect 480 15525 485 15555
rect 515 15525 520 15555
rect 480 15520 520 15525
rect 560 15555 600 15560
rect 560 15525 565 15555
rect 595 15525 600 15555
rect 560 15520 600 15525
rect 640 15555 680 15560
rect 640 15525 645 15555
rect 675 15525 680 15555
rect 640 15520 680 15525
rect 720 15555 760 15560
rect 720 15525 725 15555
rect 755 15525 760 15555
rect 720 15520 760 15525
rect 800 15555 840 15560
rect 800 15525 805 15555
rect 835 15525 840 15555
rect 800 15520 840 15525
rect 880 15555 920 15560
rect 880 15525 885 15555
rect 915 15525 920 15555
rect 880 15520 920 15525
rect 960 15555 1000 15560
rect 960 15525 965 15555
rect 995 15525 1000 15555
rect 960 15520 1000 15525
rect 1040 15555 1080 15560
rect 1040 15525 1045 15555
rect 1075 15525 1080 15555
rect 1040 15520 1080 15525
rect 1120 15555 1160 15560
rect 1120 15525 1125 15555
rect 1155 15525 1160 15555
rect 1120 15520 1160 15525
rect 1200 15555 1240 15560
rect 1200 15525 1205 15555
rect 1235 15525 1240 15555
rect 1200 15520 1240 15525
rect 1280 15555 1320 15560
rect 1280 15525 1285 15555
rect 1315 15525 1320 15555
rect 1280 15520 1320 15525
rect 1360 15555 1400 15560
rect 1360 15525 1365 15555
rect 1395 15525 1400 15555
rect 1360 15520 1400 15525
rect 1440 15555 1480 15560
rect 1440 15525 1445 15555
rect 1475 15525 1480 15555
rect 1440 15520 1480 15525
rect 1520 15555 1560 15560
rect 1520 15525 1525 15555
rect 1555 15525 1560 15555
rect 1520 15520 1560 15525
rect 1600 15555 1640 15560
rect 1600 15525 1605 15555
rect 1635 15525 1640 15555
rect 1600 15520 1640 15525
rect 1680 15555 1720 15560
rect 1680 15525 1685 15555
rect 1715 15525 1720 15555
rect 1680 15520 1720 15525
rect 1760 15555 1800 15560
rect 1760 15525 1765 15555
rect 1795 15525 1800 15555
rect 1760 15520 1800 15525
rect 1840 15555 1880 15560
rect 1840 15525 1845 15555
rect 1875 15525 1880 15555
rect 1840 15520 1880 15525
rect 1920 15555 1960 15560
rect 1920 15525 1925 15555
rect 1955 15525 1960 15555
rect 1920 15520 1960 15525
rect 2000 15555 2040 15560
rect 2000 15525 2005 15555
rect 2035 15525 2040 15555
rect 2000 15520 2040 15525
rect 2080 15555 2120 15560
rect 2080 15525 2085 15555
rect 2115 15525 2120 15555
rect 2080 15520 2120 15525
rect 2160 15555 2200 15560
rect 2160 15525 2165 15555
rect 2195 15525 2200 15555
rect 2160 15520 2200 15525
rect 2240 15555 2280 15560
rect 2240 15525 2245 15555
rect 2275 15525 2280 15555
rect 2240 15520 2280 15525
rect 2320 15555 2360 15560
rect 2320 15525 2325 15555
rect 2355 15525 2360 15555
rect 2320 15520 2360 15525
rect 2400 15555 2440 15560
rect 2400 15525 2405 15555
rect 2435 15525 2440 15555
rect 2400 15520 2440 15525
rect 2480 15555 2520 15560
rect 2480 15525 2485 15555
rect 2515 15525 2520 15555
rect 2480 15520 2520 15525
rect 2560 15555 2600 15560
rect 2560 15525 2565 15555
rect 2595 15525 2600 15555
rect 2560 15520 2600 15525
rect 2640 15555 2680 15560
rect 2640 15525 2645 15555
rect 2675 15525 2680 15555
rect 2640 15520 2680 15525
rect 2720 15555 2760 15560
rect 2720 15525 2725 15555
rect 2755 15525 2760 15555
rect 2720 15520 2760 15525
rect 2800 15555 2840 15560
rect 2800 15525 2805 15555
rect 2835 15525 2840 15555
rect 2800 15520 2840 15525
rect 2880 15555 2920 15560
rect 2880 15525 2885 15555
rect 2915 15525 2920 15555
rect 2880 15520 2920 15525
rect 2960 15555 3000 15560
rect 2960 15525 2965 15555
rect 2995 15525 3000 15555
rect 2960 15520 3000 15525
rect 3040 15555 3080 15560
rect 3040 15525 3045 15555
rect 3075 15525 3080 15555
rect 3040 15520 3080 15525
rect 3120 15555 3160 15560
rect 3120 15525 3125 15555
rect 3155 15525 3160 15555
rect 3120 15520 3160 15525
rect 3200 15555 3240 15560
rect 3200 15525 3205 15555
rect 3235 15525 3240 15555
rect 3200 15520 3240 15525
rect 3280 15555 3320 15560
rect 3280 15525 3285 15555
rect 3315 15525 3320 15555
rect 3280 15520 3320 15525
rect 3360 15555 3400 15560
rect 3360 15525 3365 15555
rect 3395 15525 3400 15555
rect 3360 15520 3400 15525
rect 3440 15555 3480 15560
rect 3440 15525 3445 15555
rect 3475 15525 3480 15555
rect 3440 15520 3480 15525
rect 3520 15555 3560 15560
rect 3520 15525 3525 15555
rect 3555 15525 3560 15555
rect 3520 15520 3560 15525
rect 3600 15555 3640 15560
rect 3600 15525 3605 15555
rect 3635 15525 3640 15555
rect 3600 15520 3640 15525
rect 3680 15555 3720 15560
rect 3680 15525 3685 15555
rect 3715 15525 3720 15555
rect 3680 15520 3720 15525
rect 3760 15555 3800 15560
rect 3760 15525 3765 15555
rect 3795 15525 3800 15555
rect 3760 15520 3800 15525
rect 3840 15555 3880 15560
rect 3840 15525 3845 15555
rect 3875 15525 3880 15555
rect 3840 15520 3880 15525
rect 3920 15555 3960 15560
rect 3920 15525 3925 15555
rect 3955 15525 3960 15555
rect 3920 15520 3960 15525
rect 4000 15555 4040 15560
rect 4000 15525 4005 15555
rect 4035 15525 4040 15555
rect 4000 15520 4040 15525
rect 4080 15555 4120 15560
rect 4080 15525 4085 15555
rect 4115 15525 4120 15555
rect 4080 15520 4120 15525
rect 4160 15555 4200 15560
rect 4160 15525 4165 15555
rect 4195 15525 4200 15555
rect 4160 15520 4200 15525
rect 6240 15555 6280 15560
rect 6240 15525 6245 15555
rect 6275 15525 6280 15555
rect 6240 15520 6280 15525
rect 6320 15555 6360 15560
rect 6320 15525 6325 15555
rect 6355 15525 6360 15555
rect 6320 15520 6360 15525
rect 6400 15555 6440 15560
rect 6400 15525 6405 15555
rect 6435 15525 6440 15555
rect 6400 15520 6440 15525
rect 6480 15555 6520 15560
rect 6480 15525 6485 15555
rect 6515 15525 6520 15555
rect 6480 15520 6520 15525
rect 6560 15555 6600 15560
rect 6560 15525 6565 15555
rect 6595 15525 6600 15555
rect 6560 15520 6600 15525
rect 6640 15555 6680 15560
rect 6640 15525 6645 15555
rect 6675 15525 6680 15555
rect 6640 15520 6680 15525
rect 6720 15555 6760 15560
rect 6720 15525 6725 15555
rect 6755 15525 6760 15555
rect 6720 15520 6760 15525
rect 6800 15555 6840 15560
rect 6800 15525 6805 15555
rect 6835 15525 6840 15555
rect 6800 15520 6840 15525
rect 6880 15555 6920 15560
rect 6880 15525 6885 15555
rect 6915 15525 6920 15555
rect 6880 15520 6920 15525
rect 6960 15555 7000 15560
rect 6960 15525 6965 15555
rect 6995 15525 7000 15555
rect 6960 15520 7000 15525
rect 7040 15555 7080 15560
rect 7040 15525 7045 15555
rect 7075 15525 7080 15555
rect 7040 15520 7080 15525
rect 7120 15555 7160 15560
rect 7120 15525 7125 15555
rect 7155 15525 7160 15555
rect 7120 15520 7160 15525
rect 7200 15555 7240 15560
rect 7200 15525 7205 15555
rect 7235 15525 7240 15555
rect 7200 15520 7240 15525
rect 7280 15555 7320 15560
rect 7280 15525 7285 15555
rect 7315 15525 7320 15555
rect 7280 15520 7320 15525
rect 7360 15555 7400 15560
rect 7360 15525 7365 15555
rect 7395 15525 7400 15555
rect 7360 15520 7400 15525
rect 7440 15555 7480 15560
rect 7440 15525 7445 15555
rect 7475 15525 7480 15555
rect 7440 15520 7480 15525
rect 7520 15555 7560 15560
rect 7520 15525 7525 15555
rect 7555 15525 7560 15555
rect 7520 15520 7560 15525
rect 7600 15555 7640 15560
rect 7600 15525 7605 15555
rect 7635 15525 7640 15555
rect 7600 15520 7640 15525
rect 7680 15555 7720 15560
rect 7680 15525 7685 15555
rect 7715 15525 7720 15555
rect 7680 15520 7720 15525
rect 7760 15555 7800 15560
rect 7760 15525 7765 15555
rect 7795 15525 7800 15555
rect 7760 15520 7800 15525
rect 7840 15555 7880 15560
rect 7840 15525 7845 15555
rect 7875 15525 7880 15555
rect 7840 15520 7880 15525
rect 7920 15555 7960 15560
rect 7920 15525 7925 15555
rect 7955 15525 7960 15555
rect 7920 15520 7960 15525
rect 8000 15555 8040 15560
rect 8000 15525 8005 15555
rect 8035 15525 8040 15555
rect 8000 15520 8040 15525
rect 8080 15555 8120 15560
rect 8080 15525 8085 15555
rect 8115 15525 8120 15555
rect 8080 15520 8120 15525
rect 8160 15555 8200 15560
rect 8160 15525 8165 15555
rect 8195 15525 8200 15555
rect 8160 15520 8200 15525
rect 8240 15555 8280 15560
rect 8240 15525 8245 15555
rect 8275 15525 8280 15555
rect 8240 15520 8280 15525
rect 8320 15555 8360 15560
rect 8320 15525 8325 15555
rect 8355 15525 8360 15555
rect 8320 15520 8360 15525
rect 8400 15555 8440 15560
rect 8400 15525 8405 15555
rect 8435 15525 8440 15555
rect 8400 15520 8440 15525
rect 8480 15555 8520 15560
rect 8480 15525 8485 15555
rect 8515 15525 8520 15555
rect 8480 15520 8520 15525
rect 8560 15555 8600 15560
rect 8560 15525 8565 15555
rect 8595 15525 8600 15555
rect 8560 15520 8600 15525
rect 8640 15555 8680 15560
rect 8640 15525 8645 15555
rect 8675 15525 8680 15555
rect 8640 15520 8680 15525
rect 8720 15555 8760 15560
rect 8720 15525 8725 15555
rect 8755 15525 8760 15555
rect 8720 15520 8760 15525
rect 8800 15555 8840 15560
rect 8800 15525 8805 15555
rect 8835 15525 8840 15555
rect 8800 15520 8840 15525
rect 8880 15555 8920 15560
rect 8880 15525 8885 15555
rect 8915 15525 8920 15555
rect 8880 15520 8920 15525
rect 8960 15555 9000 15560
rect 8960 15525 8965 15555
rect 8995 15525 9000 15555
rect 8960 15520 9000 15525
rect 9040 15555 9080 15560
rect 9040 15525 9045 15555
rect 9075 15525 9080 15555
rect 9040 15520 9080 15525
rect 9120 15555 9160 15560
rect 9120 15525 9125 15555
rect 9155 15525 9160 15555
rect 9120 15520 9160 15525
rect 9200 15555 9240 15560
rect 9200 15525 9205 15555
rect 9235 15525 9240 15555
rect 9200 15520 9240 15525
rect 9280 15555 9320 15560
rect 9280 15525 9285 15555
rect 9315 15525 9320 15555
rect 9280 15520 9320 15525
rect 9360 15555 9400 15560
rect 9360 15525 9365 15555
rect 9395 15525 9400 15555
rect 9360 15520 9400 15525
rect 9440 15555 9480 15560
rect 9440 15525 9445 15555
rect 9475 15525 9480 15555
rect 9440 15520 9480 15525
rect 11560 15555 11600 15560
rect 11560 15525 11565 15555
rect 11595 15525 11600 15555
rect 11560 15520 11600 15525
rect 11640 15555 11680 15560
rect 11640 15525 11645 15555
rect 11675 15525 11680 15555
rect 11640 15520 11680 15525
rect 11720 15555 11760 15560
rect 11720 15525 11725 15555
rect 11755 15525 11760 15555
rect 11720 15520 11760 15525
rect 11800 15555 11840 15560
rect 11800 15525 11805 15555
rect 11835 15525 11840 15555
rect 11800 15520 11840 15525
rect 11880 15555 11920 15560
rect 11880 15525 11885 15555
rect 11915 15525 11920 15555
rect 11880 15520 11920 15525
rect 11960 15555 12000 15560
rect 11960 15525 11965 15555
rect 11995 15525 12000 15555
rect 11960 15520 12000 15525
rect 12040 15555 12080 15560
rect 12040 15525 12045 15555
rect 12075 15525 12080 15555
rect 12040 15520 12080 15525
rect 12120 15555 12160 15560
rect 12120 15525 12125 15555
rect 12155 15525 12160 15555
rect 12120 15520 12160 15525
rect 12200 15555 12240 15560
rect 12200 15525 12205 15555
rect 12235 15525 12240 15555
rect 12200 15520 12240 15525
rect 12280 15555 12320 15560
rect 12280 15525 12285 15555
rect 12315 15525 12320 15555
rect 12280 15520 12320 15525
rect 12360 15555 12400 15560
rect 12360 15525 12365 15555
rect 12395 15525 12400 15555
rect 12360 15520 12400 15525
rect 12440 15555 12480 15560
rect 12440 15525 12445 15555
rect 12475 15525 12480 15555
rect 12440 15520 12480 15525
rect 12520 15555 12560 15560
rect 12520 15525 12525 15555
rect 12555 15525 12560 15555
rect 12520 15520 12560 15525
rect 12600 15555 12640 15560
rect 12600 15525 12605 15555
rect 12635 15525 12640 15555
rect 12600 15520 12640 15525
rect 12680 15555 12720 15560
rect 12680 15525 12685 15555
rect 12715 15525 12720 15555
rect 12680 15520 12720 15525
rect 12760 15555 12800 15560
rect 12760 15525 12765 15555
rect 12795 15525 12800 15555
rect 12760 15520 12800 15525
rect 12840 15555 12880 15560
rect 12840 15525 12845 15555
rect 12875 15525 12880 15555
rect 12840 15520 12880 15525
rect 12920 15555 12960 15560
rect 12920 15525 12925 15555
rect 12955 15525 12960 15555
rect 12920 15520 12960 15525
rect 13000 15555 13040 15560
rect 13000 15525 13005 15555
rect 13035 15525 13040 15555
rect 13000 15520 13040 15525
rect 13080 15555 13120 15560
rect 13080 15525 13085 15555
rect 13115 15525 13120 15555
rect 13080 15520 13120 15525
rect 13160 15555 13200 15560
rect 13160 15525 13165 15555
rect 13195 15525 13200 15555
rect 13160 15520 13200 15525
rect 13240 15555 13280 15560
rect 13240 15525 13245 15555
rect 13275 15525 13280 15555
rect 13240 15520 13280 15525
rect 13320 15555 13360 15560
rect 13320 15525 13325 15555
rect 13355 15525 13360 15555
rect 13320 15520 13360 15525
rect 13400 15555 13440 15560
rect 13400 15525 13405 15555
rect 13435 15525 13440 15555
rect 13400 15520 13440 15525
rect 13480 15555 13520 15560
rect 13480 15525 13485 15555
rect 13515 15525 13520 15555
rect 13480 15520 13520 15525
rect 13560 15555 13600 15560
rect 13560 15525 13565 15555
rect 13595 15525 13600 15555
rect 13560 15520 13600 15525
rect 13640 15555 13680 15560
rect 13640 15525 13645 15555
rect 13675 15525 13680 15555
rect 13640 15520 13680 15525
rect 13720 15555 13760 15560
rect 13720 15525 13725 15555
rect 13755 15525 13760 15555
rect 13720 15520 13760 15525
rect 13800 15555 13840 15560
rect 13800 15525 13805 15555
rect 13835 15525 13840 15555
rect 13800 15520 13840 15525
rect 13880 15555 13920 15560
rect 13880 15525 13885 15555
rect 13915 15525 13920 15555
rect 13880 15520 13920 15525
rect 13960 15555 14000 15560
rect 13960 15525 13965 15555
rect 13995 15525 14000 15555
rect 13960 15520 14000 15525
rect 14040 15555 14080 15560
rect 14040 15525 14045 15555
rect 14075 15525 14080 15555
rect 14040 15520 14080 15525
rect 14120 15555 14160 15560
rect 14120 15525 14125 15555
rect 14155 15525 14160 15555
rect 14120 15520 14160 15525
rect 14200 15555 14240 15560
rect 14200 15525 14205 15555
rect 14235 15525 14240 15555
rect 14200 15520 14240 15525
rect 14280 15555 14320 15560
rect 14280 15525 14285 15555
rect 14315 15525 14320 15555
rect 14280 15520 14320 15525
rect 14360 15555 14400 15560
rect 14360 15525 14365 15555
rect 14395 15525 14400 15555
rect 14360 15520 14400 15525
rect 14440 15555 14480 15560
rect 14440 15525 14445 15555
rect 14475 15525 14480 15555
rect 14440 15520 14480 15525
rect 14520 15555 14560 15560
rect 14520 15525 14525 15555
rect 14555 15525 14560 15555
rect 14520 15520 14560 15525
rect 14600 15555 14640 15560
rect 14600 15525 14605 15555
rect 14635 15525 14640 15555
rect 14600 15520 14640 15525
rect 14680 15555 14720 15560
rect 14680 15525 14685 15555
rect 14715 15525 14720 15555
rect 14680 15520 14720 15525
rect 16760 15555 16800 15560
rect 16760 15525 16765 15555
rect 16795 15525 16800 15555
rect 16760 15520 16800 15525
rect 16840 15555 16880 15560
rect 16840 15525 16845 15555
rect 16875 15525 16880 15555
rect 16840 15520 16880 15525
rect 16920 15555 16960 15560
rect 16920 15525 16925 15555
rect 16955 15525 16960 15555
rect 16920 15520 16960 15525
rect 17000 15555 17040 15560
rect 17000 15525 17005 15555
rect 17035 15525 17040 15555
rect 17000 15520 17040 15525
rect 17080 15555 17120 15560
rect 17080 15525 17085 15555
rect 17115 15525 17120 15555
rect 17080 15520 17120 15525
rect 17160 15555 17200 15560
rect 17160 15525 17165 15555
rect 17195 15525 17200 15555
rect 17160 15520 17200 15525
rect 17240 15555 17280 15560
rect 17240 15525 17245 15555
rect 17275 15525 17280 15555
rect 17240 15520 17280 15525
rect 17320 15555 17360 15560
rect 17320 15525 17325 15555
rect 17355 15525 17360 15555
rect 17320 15520 17360 15525
rect 17400 15555 17440 15560
rect 17400 15525 17405 15555
rect 17435 15525 17440 15555
rect 17400 15520 17440 15525
rect 17480 15555 17520 15560
rect 17480 15525 17485 15555
rect 17515 15525 17520 15555
rect 17480 15520 17520 15525
rect 17560 15555 17600 15560
rect 17560 15525 17565 15555
rect 17595 15525 17600 15555
rect 17560 15520 17600 15525
rect 17640 15555 17680 15560
rect 17640 15525 17645 15555
rect 17675 15525 17680 15555
rect 17640 15520 17680 15525
rect 17720 15555 17760 15560
rect 17720 15525 17725 15555
rect 17755 15525 17760 15555
rect 17720 15520 17760 15525
rect 17800 15555 17840 15560
rect 17800 15525 17805 15555
rect 17835 15525 17840 15555
rect 17800 15520 17840 15525
rect 17880 15555 17920 15560
rect 17880 15525 17885 15555
rect 17915 15525 17920 15555
rect 17880 15520 17920 15525
rect 17960 15555 18000 15560
rect 17960 15525 17965 15555
rect 17995 15525 18000 15555
rect 17960 15520 18000 15525
rect 18040 15555 18080 15560
rect 18040 15525 18045 15555
rect 18075 15525 18080 15555
rect 18040 15520 18080 15525
rect 18120 15555 18160 15560
rect 18120 15525 18125 15555
rect 18155 15525 18160 15555
rect 18120 15520 18160 15525
rect 18200 15555 18240 15560
rect 18200 15525 18205 15555
rect 18235 15525 18240 15555
rect 18200 15520 18240 15525
rect 18280 15555 18320 15560
rect 18280 15525 18285 15555
rect 18315 15525 18320 15555
rect 18280 15520 18320 15525
rect 18360 15555 18400 15560
rect 18360 15525 18365 15555
rect 18395 15525 18400 15555
rect 18360 15520 18400 15525
rect 18440 15555 18480 15560
rect 18440 15525 18445 15555
rect 18475 15525 18480 15555
rect 18440 15520 18480 15525
rect 18520 15555 18560 15560
rect 18520 15525 18525 15555
rect 18555 15525 18560 15555
rect 18520 15520 18560 15525
rect 18600 15555 18640 15560
rect 18600 15525 18605 15555
rect 18635 15525 18640 15555
rect 18600 15520 18640 15525
rect 18680 15555 18720 15560
rect 18680 15525 18685 15555
rect 18715 15525 18720 15555
rect 18680 15520 18720 15525
rect 18760 15555 18800 15560
rect 18760 15525 18765 15555
rect 18795 15525 18800 15555
rect 18760 15520 18800 15525
rect 18840 15555 18880 15560
rect 18840 15525 18845 15555
rect 18875 15525 18880 15555
rect 18840 15520 18880 15525
rect 18920 15555 18960 15560
rect 18920 15525 18925 15555
rect 18955 15525 18960 15555
rect 18920 15520 18960 15525
rect 19000 15555 19040 15560
rect 19000 15525 19005 15555
rect 19035 15525 19040 15555
rect 19000 15520 19040 15525
rect 19080 15555 19120 15560
rect 19080 15525 19085 15555
rect 19115 15525 19120 15555
rect 19080 15520 19120 15525
rect 19160 15555 19200 15560
rect 19160 15525 19165 15555
rect 19195 15525 19200 15555
rect 19160 15520 19200 15525
rect 19240 15555 19280 15560
rect 19240 15525 19245 15555
rect 19275 15525 19280 15555
rect 19240 15520 19280 15525
rect 19320 15555 19360 15560
rect 19320 15525 19325 15555
rect 19355 15525 19360 15555
rect 19320 15520 19360 15525
rect 19400 15555 19440 15560
rect 19400 15525 19405 15555
rect 19435 15525 19440 15555
rect 19400 15520 19440 15525
rect 19480 15555 19520 15560
rect 19480 15525 19485 15555
rect 19515 15525 19520 15555
rect 19480 15520 19520 15525
rect 19560 15555 19600 15560
rect 19560 15525 19565 15555
rect 19595 15525 19600 15555
rect 19560 15520 19600 15525
rect 19640 15555 19680 15560
rect 19640 15525 19645 15555
rect 19675 15525 19680 15555
rect 19640 15520 19680 15525
rect 19720 15555 19760 15560
rect 19720 15525 19725 15555
rect 19755 15525 19760 15555
rect 19720 15520 19760 15525
rect 19800 15555 19840 15560
rect 19800 15525 19805 15555
rect 19835 15525 19840 15555
rect 19800 15520 19840 15525
rect 19880 15555 19920 15560
rect 19880 15525 19885 15555
rect 19915 15525 19920 15555
rect 19880 15520 19920 15525
rect 19960 15555 20000 15560
rect 19960 15525 19965 15555
rect 19995 15525 20000 15555
rect 19960 15520 20000 15525
rect 20040 15555 20080 15560
rect 20040 15525 20045 15555
rect 20075 15525 20080 15555
rect 20040 15520 20080 15525
rect 20120 15555 20160 15560
rect 20120 15525 20125 15555
rect 20155 15525 20160 15555
rect 20120 15520 20160 15525
rect 20200 15555 20240 15560
rect 20200 15525 20205 15555
rect 20235 15525 20240 15555
rect 20200 15520 20240 15525
rect 20280 15555 20320 15560
rect 20280 15525 20285 15555
rect 20315 15525 20320 15555
rect 20280 15520 20320 15525
rect 20360 15555 20400 15560
rect 20360 15525 20365 15555
rect 20395 15525 20400 15555
rect 20360 15520 20400 15525
rect 20440 15555 20480 15560
rect 20440 15525 20445 15555
rect 20475 15525 20480 15555
rect 20440 15520 20480 15525
rect 20520 15555 20560 15560
rect 20520 15525 20525 15555
rect 20555 15525 20560 15555
rect 20520 15520 20560 15525
rect 20600 15555 20640 15560
rect 20600 15525 20605 15555
rect 20635 15525 20640 15555
rect 20600 15520 20640 15525
rect 20680 15555 20720 15560
rect 20680 15525 20685 15555
rect 20715 15525 20720 15555
rect 20680 15520 20720 15525
rect 20760 15555 20800 15560
rect 20760 15525 20765 15555
rect 20795 15525 20800 15555
rect 20760 15520 20800 15525
rect 20840 15555 20880 15560
rect 20840 15525 20845 15555
rect 20875 15525 20880 15555
rect 20840 15520 20880 15525
rect 20920 15555 20960 15560
rect 20920 15525 20925 15555
rect 20955 15525 20960 15555
rect 20920 15520 20960 15525
rect 0 15395 40 15400
rect 0 15365 5 15395
rect 35 15365 40 15395
rect 0 15360 40 15365
rect 80 15395 120 15400
rect 80 15365 85 15395
rect 115 15365 120 15395
rect 80 15360 120 15365
rect 160 15395 200 15400
rect 160 15365 165 15395
rect 195 15365 200 15395
rect 160 15360 200 15365
rect 240 15395 280 15400
rect 240 15365 245 15395
rect 275 15365 280 15395
rect 240 15360 280 15365
rect 320 15395 360 15400
rect 320 15365 325 15395
rect 355 15365 360 15395
rect 320 15360 360 15365
rect 400 15395 440 15400
rect 400 15365 405 15395
rect 435 15365 440 15395
rect 400 15360 440 15365
rect 480 15395 520 15400
rect 480 15365 485 15395
rect 515 15365 520 15395
rect 480 15360 520 15365
rect 560 15395 600 15400
rect 560 15365 565 15395
rect 595 15365 600 15395
rect 560 15360 600 15365
rect 640 15395 680 15400
rect 640 15365 645 15395
rect 675 15365 680 15395
rect 640 15360 680 15365
rect 720 15395 760 15400
rect 720 15365 725 15395
rect 755 15365 760 15395
rect 720 15360 760 15365
rect 800 15395 840 15400
rect 800 15365 805 15395
rect 835 15365 840 15395
rect 800 15360 840 15365
rect 880 15395 920 15400
rect 880 15365 885 15395
rect 915 15365 920 15395
rect 880 15360 920 15365
rect 960 15395 1000 15400
rect 960 15365 965 15395
rect 995 15365 1000 15395
rect 960 15360 1000 15365
rect 1040 15395 1080 15400
rect 1040 15365 1045 15395
rect 1075 15365 1080 15395
rect 1040 15360 1080 15365
rect 1120 15395 1160 15400
rect 1120 15365 1125 15395
rect 1155 15365 1160 15395
rect 1120 15360 1160 15365
rect 1200 15395 1240 15400
rect 1200 15365 1205 15395
rect 1235 15365 1240 15395
rect 1200 15360 1240 15365
rect 1280 15395 1320 15400
rect 1280 15365 1285 15395
rect 1315 15365 1320 15395
rect 1280 15360 1320 15365
rect 1360 15395 1400 15400
rect 1360 15365 1365 15395
rect 1395 15365 1400 15395
rect 1360 15360 1400 15365
rect 1440 15395 1480 15400
rect 1440 15365 1445 15395
rect 1475 15365 1480 15395
rect 1440 15360 1480 15365
rect 1520 15395 1560 15400
rect 1520 15365 1525 15395
rect 1555 15365 1560 15395
rect 1520 15360 1560 15365
rect 1600 15395 1640 15400
rect 1600 15365 1605 15395
rect 1635 15365 1640 15395
rect 1600 15360 1640 15365
rect 1680 15395 1720 15400
rect 1680 15365 1685 15395
rect 1715 15365 1720 15395
rect 1680 15360 1720 15365
rect 1760 15395 1800 15400
rect 1760 15365 1765 15395
rect 1795 15365 1800 15395
rect 1760 15360 1800 15365
rect 1840 15395 1880 15400
rect 1840 15365 1845 15395
rect 1875 15365 1880 15395
rect 1840 15360 1880 15365
rect 1920 15395 1960 15400
rect 1920 15365 1925 15395
rect 1955 15365 1960 15395
rect 1920 15360 1960 15365
rect 2000 15395 2040 15400
rect 2000 15365 2005 15395
rect 2035 15365 2040 15395
rect 2000 15360 2040 15365
rect 2080 15395 2120 15400
rect 2080 15365 2085 15395
rect 2115 15365 2120 15395
rect 2080 15360 2120 15365
rect 2160 15395 2200 15400
rect 2160 15365 2165 15395
rect 2195 15365 2200 15395
rect 2160 15360 2200 15365
rect 2240 15395 2280 15400
rect 2240 15365 2245 15395
rect 2275 15365 2280 15395
rect 2240 15360 2280 15365
rect 2320 15395 2360 15400
rect 2320 15365 2325 15395
rect 2355 15365 2360 15395
rect 2320 15360 2360 15365
rect 2400 15395 2440 15400
rect 2400 15365 2405 15395
rect 2435 15365 2440 15395
rect 2400 15360 2440 15365
rect 2480 15395 2520 15400
rect 2480 15365 2485 15395
rect 2515 15365 2520 15395
rect 2480 15360 2520 15365
rect 2560 15395 2600 15400
rect 2560 15365 2565 15395
rect 2595 15365 2600 15395
rect 2560 15360 2600 15365
rect 2640 15395 2680 15400
rect 2640 15365 2645 15395
rect 2675 15365 2680 15395
rect 2640 15360 2680 15365
rect 2720 15395 2760 15400
rect 2720 15365 2725 15395
rect 2755 15365 2760 15395
rect 2720 15360 2760 15365
rect 2800 15395 2840 15400
rect 2800 15365 2805 15395
rect 2835 15365 2840 15395
rect 2800 15360 2840 15365
rect 2880 15395 2920 15400
rect 2880 15365 2885 15395
rect 2915 15365 2920 15395
rect 2880 15360 2920 15365
rect 2960 15395 3000 15400
rect 2960 15365 2965 15395
rect 2995 15365 3000 15395
rect 2960 15360 3000 15365
rect 3040 15395 3080 15400
rect 3040 15365 3045 15395
rect 3075 15365 3080 15395
rect 3040 15360 3080 15365
rect 3120 15395 3160 15400
rect 3120 15365 3125 15395
rect 3155 15365 3160 15395
rect 3120 15360 3160 15365
rect 3200 15395 3240 15400
rect 3200 15365 3205 15395
rect 3235 15365 3240 15395
rect 3200 15360 3240 15365
rect 3280 15395 3320 15400
rect 3280 15365 3285 15395
rect 3315 15365 3320 15395
rect 3280 15360 3320 15365
rect 3360 15395 3400 15400
rect 3360 15365 3365 15395
rect 3395 15365 3400 15395
rect 3360 15360 3400 15365
rect 3440 15395 3480 15400
rect 3440 15365 3445 15395
rect 3475 15365 3480 15395
rect 3440 15360 3480 15365
rect 3520 15395 3560 15400
rect 3520 15365 3525 15395
rect 3555 15365 3560 15395
rect 3520 15360 3560 15365
rect 3600 15395 3640 15400
rect 3600 15365 3605 15395
rect 3635 15365 3640 15395
rect 3600 15360 3640 15365
rect 3680 15395 3720 15400
rect 3680 15365 3685 15395
rect 3715 15365 3720 15395
rect 3680 15360 3720 15365
rect 3760 15395 3800 15400
rect 3760 15365 3765 15395
rect 3795 15365 3800 15395
rect 3760 15360 3800 15365
rect 3840 15395 3880 15400
rect 3840 15365 3845 15395
rect 3875 15365 3880 15395
rect 3840 15360 3880 15365
rect 3920 15395 3960 15400
rect 3920 15365 3925 15395
rect 3955 15365 3960 15395
rect 3920 15360 3960 15365
rect 4000 15395 4040 15400
rect 4000 15365 4005 15395
rect 4035 15365 4040 15395
rect 4000 15360 4040 15365
rect 4080 15395 4120 15400
rect 4080 15365 4085 15395
rect 4115 15365 4120 15395
rect 4080 15360 4120 15365
rect 4160 15395 4200 15400
rect 4160 15365 4165 15395
rect 4195 15365 4200 15395
rect 4160 15360 4200 15365
rect 6240 15395 6280 15400
rect 6240 15365 6245 15395
rect 6275 15365 6280 15395
rect 6240 15360 6280 15365
rect 6320 15395 6360 15400
rect 6320 15365 6325 15395
rect 6355 15365 6360 15395
rect 6320 15360 6360 15365
rect 6400 15395 6440 15400
rect 6400 15365 6405 15395
rect 6435 15365 6440 15395
rect 6400 15360 6440 15365
rect 6480 15395 6520 15400
rect 6480 15365 6485 15395
rect 6515 15365 6520 15395
rect 6480 15360 6520 15365
rect 6560 15395 6600 15400
rect 6560 15365 6565 15395
rect 6595 15365 6600 15395
rect 6560 15360 6600 15365
rect 6640 15395 6680 15400
rect 6640 15365 6645 15395
rect 6675 15365 6680 15395
rect 6640 15360 6680 15365
rect 6720 15395 6760 15400
rect 6720 15365 6725 15395
rect 6755 15365 6760 15395
rect 6720 15360 6760 15365
rect 6800 15395 6840 15400
rect 6800 15365 6805 15395
rect 6835 15365 6840 15395
rect 6800 15360 6840 15365
rect 6880 15395 6920 15400
rect 6880 15365 6885 15395
rect 6915 15365 6920 15395
rect 6880 15360 6920 15365
rect 6960 15395 7000 15400
rect 6960 15365 6965 15395
rect 6995 15365 7000 15395
rect 6960 15360 7000 15365
rect 7040 15395 7080 15400
rect 7040 15365 7045 15395
rect 7075 15365 7080 15395
rect 7040 15360 7080 15365
rect 7120 15395 7160 15400
rect 7120 15365 7125 15395
rect 7155 15365 7160 15395
rect 7120 15360 7160 15365
rect 7200 15395 7240 15400
rect 7200 15365 7205 15395
rect 7235 15365 7240 15395
rect 7200 15360 7240 15365
rect 7280 15395 7320 15400
rect 7280 15365 7285 15395
rect 7315 15365 7320 15395
rect 7280 15360 7320 15365
rect 7360 15395 7400 15400
rect 7360 15365 7365 15395
rect 7395 15365 7400 15395
rect 7360 15360 7400 15365
rect 7440 15395 7480 15400
rect 7440 15365 7445 15395
rect 7475 15365 7480 15395
rect 7440 15360 7480 15365
rect 7520 15395 7560 15400
rect 7520 15365 7525 15395
rect 7555 15365 7560 15395
rect 7520 15360 7560 15365
rect 7600 15395 7640 15400
rect 7600 15365 7605 15395
rect 7635 15365 7640 15395
rect 7600 15360 7640 15365
rect 7680 15395 7720 15400
rect 7680 15365 7685 15395
rect 7715 15365 7720 15395
rect 7680 15360 7720 15365
rect 7760 15395 7800 15400
rect 7760 15365 7765 15395
rect 7795 15365 7800 15395
rect 7760 15360 7800 15365
rect 7840 15395 7880 15400
rect 7840 15365 7845 15395
rect 7875 15365 7880 15395
rect 7840 15360 7880 15365
rect 7920 15395 7960 15400
rect 7920 15365 7925 15395
rect 7955 15365 7960 15395
rect 7920 15360 7960 15365
rect 8000 15395 8040 15400
rect 8000 15365 8005 15395
rect 8035 15365 8040 15395
rect 8000 15360 8040 15365
rect 8080 15395 8120 15400
rect 8080 15365 8085 15395
rect 8115 15365 8120 15395
rect 8080 15360 8120 15365
rect 8160 15395 8200 15400
rect 8160 15365 8165 15395
rect 8195 15365 8200 15395
rect 8160 15360 8200 15365
rect 8240 15395 8280 15400
rect 8240 15365 8245 15395
rect 8275 15365 8280 15395
rect 8240 15360 8280 15365
rect 8320 15395 8360 15400
rect 8320 15365 8325 15395
rect 8355 15365 8360 15395
rect 8320 15360 8360 15365
rect 8400 15395 8440 15400
rect 8400 15365 8405 15395
rect 8435 15365 8440 15395
rect 8400 15360 8440 15365
rect 8480 15395 8520 15400
rect 8480 15365 8485 15395
rect 8515 15365 8520 15395
rect 8480 15360 8520 15365
rect 8560 15395 8600 15400
rect 8560 15365 8565 15395
rect 8595 15365 8600 15395
rect 8560 15360 8600 15365
rect 8640 15395 8680 15400
rect 8640 15365 8645 15395
rect 8675 15365 8680 15395
rect 8640 15360 8680 15365
rect 8720 15395 8760 15400
rect 8720 15365 8725 15395
rect 8755 15365 8760 15395
rect 8720 15360 8760 15365
rect 8800 15395 8840 15400
rect 8800 15365 8805 15395
rect 8835 15365 8840 15395
rect 8800 15360 8840 15365
rect 8880 15395 8920 15400
rect 8880 15365 8885 15395
rect 8915 15365 8920 15395
rect 8880 15360 8920 15365
rect 8960 15395 9000 15400
rect 8960 15365 8965 15395
rect 8995 15365 9000 15395
rect 8960 15360 9000 15365
rect 9040 15395 9080 15400
rect 9040 15365 9045 15395
rect 9075 15365 9080 15395
rect 9040 15360 9080 15365
rect 9120 15395 9160 15400
rect 9120 15365 9125 15395
rect 9155 15365 9160 15395
rect 9120 15360 9160 15365
rect 9200 15395 9240 15400
rect 9200 15365 9205 15395
rect 9235 15365 9240 15395
rect 9200 15360 9240 15365
rect 9280 15395 9320 15400
rect 9280 15365 9285 15395
rect 9315 15365 9320 15395
rect 9280 15360 9320 15365
rect 9360 15395 9400 15400
rect 9360 15365 9365 15395
rect 9395 15365 9400 15395
rect 9360 15360 9400 15365
rect 9440 15395 9480 15400
rect 9440 15365 9445 15395
rect 9475 15365 9480 15395
rect 9440 15360 9480 15365
rect 11560 15395 11600 15400
rect 11560 15365 11565 15395
rect 11595 15365 11600 15395
rect 11560 15360 11600 15365
rect 11640 15395 11680 15400
rect 11640 15365 11645 15395
rect 11675 15365 11680 15395
rect 11640 15360 11680 15365
rect 11720 15395 11760 15400
rect 11720 15365 11725 15395
rect 11755 15365 11760 15395
rect 11720 15360 11760 15365
rect 11800 15395 11840 15400
rect 11800 15365 11805 15395
rect 11835 15365 11840 15395
rect 11800 15360 11840 15365
rect 11880 15395 11920 15400
rect 11880 15365 11885 15395
rect 11915 15365 11920 15395
rect 11880 15360 11920 15365
rect 11960 15395 12000 15400
rect 11960 15365 11965 15395
rect 11995 15365 12000 15395
rect 11960 15360 12000 15365
rect 12040 15395 12080 15400
rect 12040 15365 12045 15395
rect 12075 15365 12080 15395
rect 12040 15360 12080 15365
rect 12120 15395 12160 15400
rect 12120 15365 12125 15395
rect 12155 15365 12160 15395
rect 12120 15360 12160 15365
rect 12200 15395 12240 15400
rect 12200 15365 12205 15395
rect 12235 15365 12240 15395
rect 12200 15360 12240 15365
rect 12280 15395 12320 15400
rect 12280 15365 12285 15395
rect 12315 15365 12320 15395
rect 12280 15360 12320 15365
rect 12360 15395 12400 15400
rect 12360 15365 12365 15395
rect 12395 15365 12400 15395
rect 12360 15360 12400 15365
rect 12440 15395 12480 15400
rect 12440 15365 12445 15395
rect 12475 15365 12480 15395
rect 12440 15360 12480 15365
rect 12520 15395 12560 15400
rect 12520 15365 12525 15395
rect 12555 15365 12560 15395
rect 12520 15360 12560 15365
rect 12600 15395 12640 15400
rect 12600 15365 12605 15395
rect 12635 15365 12640 15395
rect 12600 15360 12640 15365
rect 12680 15395 12720 15400
rect 12680 15365 12685 15395
rect 12715 15365 12720 15395
rect 12680 15360 12720 15365
rect 12760 15395 12800 15400
rect 12760 15365 12765 15395
rect 12795 15365 12800 15395
rect 12760 15360 12800 15365
rect 12840 15395 12880 15400
rect 12840 15365 12845 15395
rect 12875 15365 12880 15395
rect 12840 15360 12880 15365
rect 12920 15395 12960 15400
rect 12920 15365 12925 15395
rect 12955 15365 12960 15395
rect 12920 15360 12960 15365
rect 13000 15395 13040 15400
rect 13000 15365 13005 15395
rect 13035 15365 13040 15395
rect 13000 15360 13040 15365
rect 13080 15395 13120 15400
rect 13080 15365 13085 15395
rect 13115 15365 13120 15395
rect 13080 15360 13120 15365
rect 13160 15395 13200 15400
rect 13160 15365 13165 15395
rect 13195 15365 13200 15395
rect 13160 15360 13200 15365
rect 13240 15395 13280 15400
rect 13240 15365 13245 15395
rect 13275 15365 13280 15395
rect 13240 15360 13280 15365
rect 13320 15395 13360 15400
rect 13320 15365 13325 15395
rect 13355 15365 13360 15395
rect 13320 15360 13360 15365
rect 13400 15395 13440 15400
rect 13400 15365 13405 15395
rect 13435 15365 13440 15395
rect 13400 15360 13440 15365
rect 13480 15395 13520 15400
rect 13480 15365 13485 15395
rect 13515 15365 13520 15395
rect 13480 15360 13520 15365
rect 13560 15395 13600 15400
rect 13560 15365 13565 15395
rect 13595 15365 13600 15395
rect 13560 15360 13600 15365
rect 13640 15395 13680 15400
rect 13640 15365 13645 15395
rect 13675 15365 13680 15395
rect 13640 15360 13680 15365
rect 13720 15395 13760 15400
rect 13720 15365 13725 15395
rect 13755 15365 13760 15395
rect 13720 15360 13760 15365
rect 13800 15395 13840 15400
rect 13800 15365 13805 15395
rect 13835 15365 13840 15395
rect 13800 15360 13840 15365
rect 13880 15395 13920 15400
rect 13880 15365 13885 15395
rect 13915 15365 13920 15395
rect 13880 15360 13920 15365
rect 13960 15395 14000 15400
rect 13960 15365 13965 15395
rect 13995 15365 14000 15395
rect 13960 15360 14000 15365
rect 14040 15395 14080 15400
rect 14040 15365 14045 15395
rect 14075 15365 14080 15395
rect 14040 15360 14080 15365
rect 14120 15395 14160 15400
rect 14120 15365 14125 15395
rect 14155 15365 14160 15395
rect 14120 15360 14160 15365
rect 14200 15395 14240 15400
rect 14200 15365 14205 15395
rect 14235 15365 14240 15395
rect 14200 15360 14240 15365
rect 14280 15395 14320 15400
rect 14280 15365 14285 15395
rect 14315 15365 14320 15395
rect 14280 15360 14320 15365
rect 14360 15395 14400 15400
rect 14360 15365 14365 15395
rect 14395 15365 14400 15395
rect 14360 15360 14400 15365
rect 14440 15395 14480 15400
rect 14440 15365 14445 15395
rect 14475 15365 14480 15395
rect 14440 15360 14480 15365
rect 14520 15395 14560 15400
rect 14520 15365 14525 15395
rect 14555 15365 14560 15395
rect 14520 15360 14560 15365
rect 14600 15395 14640 15400
rect 14600 15365 14605 15395
rect 14635 15365 14640 15395
rect 14600 15360 14640 15365
rect 14680 15395 14720 15400
rect 14680 15365 14685 15395
rect 14715 15365 14720 15395
rect 14680 15360 14720 15365
rect 16760 15395 16800 15400
rect 16760 15365 16765 15395
rect 16795 15365 16800 15395
rect 16760 15360 16800 15365
rect 16840 15395 16880 15400
rect 16840 15365 16845 15395
rect 16875 15365 16880 15395
rect 16840 15360 16880 15365
rect 16920 15395 16960 15400
rect 16920 15365 16925 15395
rect 16955 15365 16960 15395
rect 16920 15360 16960 15365
rect 17000 15395 17040 15400
rect 17000 15365 17005 15395
rect 17035 15365 17040 15395
rect 17000 15360 17040 15365
rect 17080 15395 17120 15400
rect 17080 15365 17085 15395
rect 17115 15365 17120 15395
rect 17080 15360 17120 15365
rect 17160 15395 17200 15400
rect 17160 15365 17165 15395
rect 17195 15365 17200 15395
rect 17160 15360 17200 15365
rect 17240 15395 17280 15400
rect 17240 15365 17245 15395
rect 17275 15365 17280 15395
rect 17240 15360 17280 15365
rect 17320 15395 17360 15400
rect 17320 15365 17325 15395
rect 17355 15365 17360 15395
rect 17320 15360 17360 15365
rect 17400 15395 17440 15400
rect 17400 15365 17405 15395
rect 17435 15365 17440 15395
rect 17400 15360 17440 15365
rect 17480 15395 17520 15400
rect 17480 15365 17485 15395
rect 17515 15365 17520 15395
rect 17480 15360 17520 15365
rect 17560 15395 17600 15400
rect 17560 15365 17565 15395
rect 17595 15365 17600 15395
rect 17560 15360 17600 15365
rect 17640 15395 17680 15400
rect 17640 15365 17645 15395
rect 17675 15365 17680 15395
rect 17640 15360 17680 15365
rect 17720 15395 17760 15400
rect 17720 15365 17725 15395
rect 17755 15365 17760 15395
rect 17720 15360 17760 15365
rect 17800 15395 17840 15400
rect 17800 15365 17805 15395
rect 17835 15365 17840 15395
rect 17800 15360 17840 15365
rect 17880 15395 17920 15400
rect 17880 15365 17885 15395
rect 17915 15365 17920 15395
rect 17880 15360 17920 15365
rect 17960 15395 18000 15400
rect 17960 15365 17965 15395
rect 17995 15365 18000 15395
rect 17960 15360 18000 15365
rect 18040 15395 18080 15400
rect 18040 15365 18045 15395
rect 18075 15365 18080 15395
rect 18040 15360 18080 15365
rect 18120 15395 18160 15400
rect 18120 15365 18125 15395
rect 18155 15365 18160 15395
rect 18120 15360 18160 15365
rect 18200 15395 18240 15400
rect 18200 15365 18205 15395
rect 18235 15365 18240 15395
rect 18200 15360 18240 15365
rect 18280 15395 18320 15400
rect 18280 15365 18285 15395
rect 18315 15365 18320 15395
rect 18280 15360 18320 15365
rect 18360 15395 18400 15400
rect 18360 15365 18365 15395
rect 18395 15365 18400 15395
rect 18360 15360 18400 15365
rect 18440 15395 18480 15400
rect 18440 15365 18445 15395
rect 18475 15365 18480 15395
rect 18440 15360 18480 15365
rect 18520 15395 18560 15400
rect 18520 15365 18525 15395
rect 18555 15365 18560 15395
rect 18520 15360 18560 15365
rect 18600 15395 18640 15400
rect 18600 15365 18605 15395
rect 18635 15365 18640 15395
rect 18600 15360 18640 15365
rect 18680 15395 18720 15400
rect 18680 15365 18685 15395
rect 18715 15365 18720 15395
rect 18680 15360 18720 15365
rect 18760 15395 18800 15400
rect 18760 15365 18765 15395
rect 18795 15365 18800 15395
rect 18760 15360 18800 15365
rect 18840 15395 18880 15400
rect 18840 15365 18845 15395
rect 18875 15365 18880 15395
rect 18840 15360 18880 15365
rect 18920 15395 18960 15400
rect 18920 15365 18925 15395
rect 18955 15365 18960 15395
rect 18920 15360 18960 15365
rect 19000 15395 19040 15400
rect 19000 15365 19005 15395
rect 19035 15365 19040 15395
rect 19000 15360 19040 15365
rect 19080 15395 19120 15400
rect 19080 15365 19085 15395
rect 19115 15365 19120 15395
rect 19080 15360 19120 15365
rect 19160 15395 19200 15400
rect 19160 15365 19165 15395
rect 19195 15365 19200 15395
rect 19160 15360 19200 15365
rect 19240 15395 19280 15400
rect 19240 15365 19245 15395
rect 19275 15365 19280 15395
rect 19240 15360 19280 15365
rect 19320 15395 19360 15400
rect 19320 15365 19325 15395
rect 19355 15365 19360 15395
rect 19320 15360 19360 15365
rect 19400 15395 19440 15400
rect 19400 15365 19405 15395
rect 19435 15365 19440 15395
rect 19400 15360 19440 15365
rect 19480 15395 19520 15400
rect 19480 15365 19485 15395
rect 19515 15365 19520 15395
rect 19480 15360 19520 15365
rect 19560 15395 19600 15400
rect 19560 15365 19565 15395
rect 19595 15365 19600 15395
rect 19560 15360 19600 15365
rect 19640 15395 19680 15400
rect 19640 15365 19645 15395
rect 19675 15365 19680 15395
rect 19640 15360 19680 15365
rect 19720 15395 19760 15400
rect 19720 15365 19725 15395
rect 19755 15365 19760 15395
rect 19720 15360 19760 15365
rect 19800 15395 19840 15400
rect 19800 15365 19805 15395
rect 19835 15365 19840 15395
rect 19800 15360 19840 15365
rect 19880 15395 19920 15400
rect 19880 15365 19885 15395
rect 19915 15365 19920 15395
rect 19880 15360 19920 15365
rect 19960 15395 20000 15400
rect 19960 15365 19965 15395
rect 19995 15365 20000 15395
rect 19960 15360 20000 15365
rect 20040 15395 20080 15400
rect 20040 15365 20045 15395
rect 20075 15365 20080 15395
rect 20040 15360 20080 15365
rect 20120 15395 20160 15400
rect 20120 15365 20125 15395
rect 20155 15365 20160 15395
rect 20120 15360 20160 15365
rect 20200 15395 20240 15400
rect 20200 15365 20205 15395
rect 20235 15365 20240 15395
rect 20200 15360 20240 15365
rect 20280 15395 20320 15400
rect 20280 15365 20285 15395
rect 20315 15365 20320 15395
rect 20280 15360 20320 15365
rect 20360 15395 20400 15400
rect 20360 15365 20365 15395
rect 20395 15365 20400 15395
rect 20360 15360 20400 15365
rect 20440 15395 20480 15400
rect 20440 15365 20445 15395
rect 20475 15365 20480 15395
rect 20440 15360 20480 15365
rect 20520 15395 20560 15400
rect 20520 15365 20525 15395
rect 20555 15365 20560 15395
rect 20520 15360 20560 15365
rect 20600 15395 20640 15400
rect 20600 15365 20605 15395
rect 20635 15365 20640 15395
rect 20600 15360 20640 15365
rect 20680 15395 20720 15400
rect 20680 15365 20685 15395
rect 20715 15365 20720 15395
rect 20680 15360 20720 15365
rect 20760 15395 20800 15400
rect 20760 15365 20765 15395
rect 20795 15365 20800 15395
rect 20760 15360 20800 15365
rect 20840 15395 20880 15400
rect 20840 15365 20845 15395
rect 20875 15365 20880 15395
rect 20840 15360 20880 15365
rect 20920 15395 20960 15400
rect 20920 15365 20925 15395
rect 20955 15365 20960 15395
rect 20920 15360 20960 15365
rect 0 15235 40 15240
rect 0 15205 5 15235
rect 35 15205 40 15235
rect 0 15200 40 15205
rect 80 15235 120 15240
rect 80 15205 85 15235
rect 115 15205 120 15235
rect 80 15200 120 15205
rect 160 15235 200 15240
rect 160 15205 165 15235
rect 195 15205 200 15235
rect 160 15200 200 15205
rect 240 15235 280 15240
rect 240 15205 245 15235
rect 275 15205 280 15235
rect 240 15200 280 15205
rect 320 15235 360 15240
rect 320 15205 325 15235
rect 355 15205 360 15235
rect 320 15200 360 15205
rect 400 15235 440 15240
rect 400 15205 405 15235
rect 435 15205 440 15235
rect 400 15200 440 15205
rect 480 15235 520 15240
rect 480 15205 485 15235
rect 515 15205 520 15235
rect 480 15200 520 15205
rect 560 15235 600 15240
rect 560 15205 565 15235
rect 595 15205 600 15235
rect 560 15200 600 15205
rect 640 15235 680 15240
rect 640 15205 645 15235
rect 675 15205 680 15235
rect 640 15200 680 15205
rect 720 15235 760 15240
rect 720 15205 725 15235
rect 755 15205 760 15235
rect 720 15200 760 15205
rect 800 15235 840 15240
rect 800 15205 805 15235
rect 835 15205 840 15235
rect 800 15200 840 15205
rect 880 15235 920 15240
rect 880 15205 885 15235
rect 915 15205 920 15235
rect 880 15200 920 15205
rect 960 15235 1000 15240
rect 960 15205 965 15235
rect 995 15205 1000 15235
rect 960 15200 1000 15205
rect 1040 15235 1080 15240
rect 1040 15205 1045 15235
rect 1075 15205 1080 15235
rect 1040 15200 1080 15205
rect 1120 15235 1160 15240
rect 1120 15205 1125 15235
rect 1155 15205 1160 15235
rect 1120 15200 1160 15205
rect 1200 15235 1240 15240
rect 1200 15205 1205 15235
rect 1235 15205 1240 15235
rect 1200 15200 1240 15205
rect 1280 15235 1320 15240
rect 1280 15205 1285 15235
rect 1315 15205 1320 15235
rect 1280 15200 1320 15205
rect 1360 15235 1400 15240
rect 1360 15205 1365 15235
rect 1395 15205 1400 15235
rect 1360 15200 1400 15205
rect 1440 15235 1480 15240
rect 1440 15205 1445 15235
rect 1475 15205 1480 15235
rect 1440 15200 1480 15205
rect 1520 15235 1560 15240
rect 1520 15205 1525 15235
rect 1555 15205 1560 15235
rect 1520 15200 1560 15205
rect 1600 15235 1640 15240
rect 1600 15205 1605 15235
rect 1635 15205 1640 15235
rect 1600 15200 1640 15205
rect 1680 15235 1720 15240
rect 1680 15205 1685 15235
rect 1715 15205 1720 15235
rect 1680 15200 1720 15205
rect 1760 15235 1800 15240
rect 1760 15205 1765 15235
rect 1795 15205 1800 15235
rect 1760 15200 1800 15205
rect 1840 15235 1880 15240
rect 1840 15205 1845 15235
rect 1875 15205 1880 15235
rect 1840 15200 1880 15205
rect 1920 15235 1960 15240
rect 1920 15205 1925 15235
rect 1955 15205 1960 15235
rect 1920 15200 1960 15205
rect 2000 15235 2040 15240
rect 2000 15205 2005 15235
rect 2035 15205 2040 15235
rect 2000 15200 2040 15205
rect 2080 15235 2120 15240
rect 2080 15205 2085 15235
rect 2115 15205 2120 15235
rect 2080 15200 2120 15205
rect 2160 15235 2200 15240
rect 2160 15205 2165 15235
rect 2195 15205 2200 15235
rect 2160 15200 2200 15205
rect 2240 15235 2280 15240
rect 2240 15205 2245 15235
rect 2275 15205 2280 15235
rect 2240 15200 2280 15205
rect 2320 15235 2360 15240
rect 2320 15205 2325 15235
rect 2355 15205 2360 15235
rect 2320 15200 2360 15205
rect 2400 15235 2440 15240
rect 2400 15205 2405 15235
rect 2435 15205 2440 15235
rect 2400 15200 2440 15205
rect 2480 15235 2520 15240
rect 2480 15205 2485 15235
rect 2515 15205 2520 15235
rect 2480 15200 2520 15205
rect 2560 15235 2600 15240
rect 2560 15205 2565 15235
rect 2595 15205 2600 15235
rect 2560 15200 2600 15205
rect 2640 15235 2680 15240
rect 2640 15205 2645 15235
rect 2675 15205 2680 15235
rect 2640 15200 2680 15205
rect 2720 15235 2760 15240
rect 2720 15205 2725 15235
rect 2755 15205 2760 15235
rect 2720 15200 2760 15205
rect 2800 15235 2840 15240
rect 2800 15205 2805 15235
rect 2835 15205 2840 15235
rect 2800 15200 2840 15205
rect 2880 15235 2920 15240
rect 2880 15205 2885 15235
rect 2915 15205 2920 15235
rect 2880 15200 2920 15205
rect 2960 15235 3000 15240
rect 2960 15205 2965 15235
rect 2995 15205 3000 15235
rect 2960 15200 3000 15205
rect 3040 15235 3080 15240
rect 3040 15205 3045 15235
rect 3075 15205 3080 15235
rect 3040 15200 3080 15205
rect 3120 15235 3160 15240
rect 3120 15205 3125 15235
rect 3155 15205 3160 15235
rect 3120 15200 3160 15205
rect 3200 15235 3240 15240
rect 3200 15205 3205 15235
rect 3235 15205 3240 15235
rect 3200 15200 3240 15205
rect 3280 15235 3320 15240
rect 3280 15205 3285 15235
rect 3315 15205 3320 15235
rect 3280 15200 3320 15205
rect 3360 15235 3400 15240
rect 3360 15205 3365 15235
rect 3395 15205 3400 15235
rect 3360 15200 3400 15205
rect 3440 15235 3480 15240
rect 3440 15205 3445 15235
rect 3475 15205 3480 15235
rect 3440 15200 3480 15205
rect 3520 15235 3560 15240
rect 3520 15205 3525 15235
rect 3555 15205 3560 15235
rect 3520 15200 3560 15205
rect 3600 15235 3640 15240
rect 3600 15205 3605 15235
rect 3635 15205 3640 15235
rect 3600 15200 3640 15205
rect 3680 15235 3720 15240
rect 3680 15205 3685 15235
rect 3715 15205 3720 15235
rect 3680 15200 3720 15205
rect 3760 15235 3800 15240
rect 3760 15205 3765 15235
rect 3795 15205 3800 15235
rect 3760 15200 3800 15205
rect 3840 15235 3880 15240
rect 3840 15205 3845 15235
rect 3875 15205 3880 15235
rect 3840 15200 3880 15205
rect 3920 15235 3960 15240
rect 3920 15205 3925 15235
rect 3955 15205 3960 15235
rect 3920 15200 3960 15205
rect 4000 15235 4040 15240
rect 4000 15205 4005 15235
rect 4035 15205 4040 15235
rect 4000 15200 4040 15205
rect 4080 15235 4120 15240
rect 4080 15205 4085 15235
rect 4115 15205 4120 15235
rect 4080 15200 4120 15205
rect 4160 15235 4200 15240
rect 4160 15205 4165 15235
rect 4195 15205 4200 15235
rect 4160 15200 4200 15205
rect 6240 15235 6280 15240
rect 6240 15205 6245 15235
rect 6275 15205 6280 15235
rect 6240 15200 6280 15205
rect 6320 15235 6360 15240
rect 6320 15205 6325 15235
rect 6355 15205 6360 15235
rect 6320 15200 6360 15205
rect 6400 15235 6440 15240
rect 6400 15205 6405 15235
rect 6435 15205 6440 15235
rect 6400 15200 6440 15205
rect 6480 15235 6520 15240
rect 6480 15205 6485 15235
rect 6515 15205 6520 15235
rect 6480 15200 6520 15205
rect 6560 15235 6600 15240
rect 6560 15205 6565 15235
rect 6595 15205 6600 15235
rect 6560 15200 6600 15205
rect 6640 15235 6680 15240
rect 6640 15205 6645 15235
rect 6675 15205 6680 15235
rect 6640 15200 6680 15205
rect 6720 15235 6760 15240
rect 6720 15205 6725 15235
rect 6755 15205 6760 15235
rect 6720 15200 6760 15205
rect 6800 15235 6840 15240
rect 6800 15205 6805 15235
rect 6835 15205 6840 15235
rect 6800 15200 6840 15205
rect 6880 15235 6920 15240
rect 6880 15205 6885 15235
rect 6915 15205 6920 15235
rect 6880 15200 6920 15205
rect 6960 15235 7000 15240
rect 6960 15205 6965 15235
rect 6995 15205 7000 15235
rect 6960 15200 7000 15205
rect 7040 15235 7080 15240
rect 7040 15205 7045 15235
rect 7075 15205 7080 15235
rect 7040 15200 7080 15205
rect 7120 15235 7160 15240
rect 7120 15205 7125 15235
rect 7155 15205 7160 15235
rect 7120 15200 7160 15205
rect 7200 15235 7240 15240
rect 7200 15205 7205 15235
rect 7235 15205 7240 15235
rect 7200 15200 7240 15205
rect 7280 15235 7320 15240
rect 7280 15205 7285 15235
rect 7315 15205 7320 15235
rect 7280 15200 7320 15205
rect 7360 15235 7400 15240
rect 7360 15205 7365 15235
rect 7395 15205 7400 15235
rect 7360 15200 7400 15205
rect 7440 15235 7480 15240
rect 7440 15205 7445 15235
rect 7475 15205 7480 15235
rect 7440 15200 7480 15205
rect 7520 15235 7560 15240
rect 7520 15205 7525 15235
rect 7555 15205 7560 15235
rect 7520 15200 7560 15205
rect 7600 15235 7640 15240
rect 7600 15205 7605 15235
rect 7635 15205 7640 15235
rect 7600 15200 7640 15205
rect 7680 15235 7720 15240
rect 7680 15205 7685 15235
rect 7715 15205 7720 15235
rect 7680 15200 7720 15205
rect 7760 15235 7800 15240
rect 7760 15205 7765 15235
rect 7795 15205 7800 15235
rect 7760 15200 7800 15205
rect 7840 15235 7880 15240
rect 7840 15205 7845 15235
rect 7875 15205 7880 15235
rect 7840 15200 7880 15205
rect 7920 15235 7960 15240
rect 7920 15205 7925 15235
rect 7955 15205 7960 15235
rect 7920 15200 7960 15205
rect 8000 15235 8040 15240
rect 8000 15205 8005 15235
rect 8035 15205 8040 15235
rect 8000 15200 8040 15205
rect 8080 15235 8120 15240
rect 8080 15205 8085 15235
rect 8115 15205 8120 15235
rect 8080 15200 8120 15205
rect 8160 15235 8200 15240
rect 8160 15205 8165 15235
rect 8195 15205 8200 15235
rect 8160 15200 8200 15205
rect 8240 15235 8280 15240
rect 8240 15205 8245 15235
rect 8275 15205 8280 15235
rect 8240 15200 8280 15205
rect 8320 15235 8360 15240
rect 8320 15205 8325 15235
rect 8355 15205 8360 15235
rect 8320 15200 8360 15205
rect 8400 15235 8440 15240
rect 8400 15205 8405 15235
rect 8435 15205 8440 15235
rect 8400 15200 8440 15205
rect 8480 15235 8520 15240
rect 8480 15205 8485 15235
rect 8515 15205 8520 15235
rect 8480 15200 8520 15205
rect 8560 15235 8600 15240
rect 8560 15205 8565 15235
rect 8595 15205 8600 15235
rect 8560 15200 8600 15205
rect 8640 15235 8680 15240
rect 8640 15205 8645 15235
rect 8675 15205 8680 15235
rect 8640 15200 8680 15205
rect 8720 15235 8760 15240
rect 8720 15205 8725 15235
rect 8755 15205 8760 15235
rect 8720 15200 8760 15205
rect 8800 15235 8840 15240
rect 8800 15205 8805 15235
rect 8835 15205 8840 15235
rect 8800 15200 8840 15205
rect 8880 15235 8920 15240
rect 8880 15205 8885 15235
rect 8915 15205 8920 15235
rect 8880 15200 8920 15205
rect 8960 15235 9000 15240
rect 8960 15205 8965 15235
rect 8995 15205 9000 15235
rect 8960 15200 9000 15205
rect 9040 15235 9080 15240
rect 9040 15205 9045 15235
rect 9075 15205 9080 15235
rect 9040 15200 9080 15205
rect 9120 15235 9160 15240
rect 9120 15205 9125 15235
rect 9155 15205 9160 15235
rect 9120 15200 9160 15205
rect 9200 15235 9240 15240
rect 9200 15205 9205 15235
rect 9235 15205 9240 15235
rect 9200 15200 9240 15205
rect 9280 15235 9320 15240
rect 9280 15205 9285 15235
rect 9315 15205 9320 15235
rect 9280 15200 9320 15205
rect 9360 15235 9400 15240
rect 9360 15205 9365 15235
rect 9395 15205 9400 15235
rect 9360 15200 9400 15205
rect 9440 15235 9480 15240
rect 9440 15205 9445 15235
rect 9475 15205 9480 15235
rect 9440 15200 9480 15205
rect 11560 15235 11600 15240
rect 11560 15205 11565 15235
rect 11595 15205 11600 15235
rect 11560 15200 11600 15205
rect 11640 15235 11680 15240
rect 11640 15205 11645 15235
rect 11675 15205 11680 15235
rect 11640 15200 11680 15205
rect 11720 15235 11760 15240
rect 11720 15205 11725 15235
rect 11755 15205 11760 15235
rect 11720 15200 11760 15205
rect 11800 15235 11840 15240
rect 11800 15205 11805 15235
rect 11835 15205 11840 15235
rect 11800 15200 11840 15205
rect 11880 15235 11920 15240
rect 11880 15205 11885 15235
rect 11915 15205 11920 15235
rect 11880 15200 11920 15205
rect 11960 15235 12000 15240
rect 11960 15205 11965 15235
rect 11995 15205 12000 15235
rect 11960 15200 12000 15205
rect 12040 15235 12080 15240
rect 12040 15205 12045 15235
rect 12075 15205 12080 15235
rect 12040 15200 12080 15205
rect 12120 15235 12160 15240
rect 12120 15205 12125 15235
rect 12155 15205 12160 15235
rect 12120 15200 12160 15205
rect 12200 15235 12240 15240
rect 12200 15205 12205 15235
rect 12235 15205 12240 15235
rect 12200 15200 12240 15205
rect 12280 15235 12320 15240
rect 12280 15205 12285 15235
rect 12315 15205 12320 15235
rect 12280 15200 12320 15205
rect 12360 15235 12400 15240
rect 12360 15205 12365 15235
rect 12395 15205 12400 15235
rect 12360 15200 12400 15205
rect 12440 15235 12480 15240
rect 12440 15205 12445 15235
rect 12475 15205 12480 15235
rect 12440 15200 12480 15205
rect 12520 15235 12560 15240
rect 12520 15205 12525 15235
rect 12555 15205 12560 15235
rect 12520 15200 12560 15205
rect 12600 15235 12640 15240
rect 12600 15205 12605 15235
rect 12635 15205 12640 15235
rect 12600 15200 12640 15205
rect 12680 15235 12720 15240
rect 12680 15205 12685 15235
rect 12715 15205 12720 15235
rect 12680 15200 12720 15205
rect 12760 15235 12800 15240
rect 12760 15205 12765 15235
rect 12795 15205 12800 15235
rect 12760 15200 12800 15205
rect 12840 15235 12880 15240
rect 12840 15205 12845 15235
rect 12875 15205 12880 15235
rect 12840 15200 12880 15205
rect 12920 15235 12960 15240
rect 12920 15205 12925 15235
rect 12955 15205 12960 15235
rect 12920 15200 12960 15205
rect 13000 15235 13040 15240
rect 13000 15205 13005 15235
rect 13035 15205 13040 15235
rect 13000 15200 13040 15205
rect 13080 15235 13120 15240
rect 13080 15205 13085 15235
rect 13115 15205 13120 15235
rect 13080 15200 13120 15205
rect 13160 15235 13200 15240
rect 13160 15205 13165 15235
rect 13195 15205 13200 15235
rect 13160 15200 13200 15205
rect 13240 15235 13280 15240
rect 13240 15205 13245 15235
rect 13275 15205 13280 15235
rect 13240 15200 13280 15205
rect 13320 15235 13360 15240
rect 13320 15205 13325 15235
rect 13355 15205 13360 15235
rect 13320 15200 13360 15205
rect 13400 15235 13440 15240
rect 13400 15205 13405 15235
rect 13435 15205 13440 15235
rect 13400 15200 13440 15205
rect 13480 15235 13520 15240
rect 13480 15205 13485 15235
rect 13515 15205 13520 15235
rect 13480 15200 13520 15205
rect 13560 15235 13600 15240
rect 13560 15205 13565 15235
rect 13595 15205 13600 15235
rect 13560 15200 13600 15205
rect 13640 15235 13680 15240
rect 13640 15205 13645 15235
rect 13675 15205 13680 15235
rect 13640 15200 13680 15205
rect 13720 15235 13760 15240
rect 13720 15205 13725 15235
rect 13755 15205 13760 15235
rect 13720 15200 13760 15205
rect 13800 15235 13840 15240
rect 13800 15205 13805 15235
rect 13835 15205 13840 15235
rect 13800 15200 13840 15205
rect 13880 15235 13920 15240
rect 13880 15205 13885 15235
rect 13915 15205 13920 15235
rect 13880 15200 13920 15205
rect 13960 15235 14000 15240
rect 13960 15205 13965 15235
rect 13995 15205 14000 15235
rect 13960 15200 14000 15205
rect 14040 15235 14080 15240
rect 14040 15205 14045 15235
rect 14075 15205 14080 15235
rect 14040 15200 14080 15205
rect 14120 15235 14160 15240
rect 14120 15205 14125 15235
rect 14155 15205 14160 15235
rect 14120 15200 14160 15205
rect 14200 15235 14240 15240
rect 14200 15205 14205 15235
rect 14235 15205 14240 15235
rect 14200 15200 14240 15205
rect 14280 15235 14320 15240
rect 14280 15205 14285 15235
rect 14315 15205 14320 15235
rect 14280 15200 14320 15205
rect 14360 15235 14400 15240
rect 14360 15205 14365 15235
rect 14395 15205 14400 15235
rect 14360 15200 14400 15205
rect 14440 15235 14480 15240
rect 14440 15205 14445 15235
rect 14475 15205 14480 15235
rect 14440 15200 14480 15205
rect 14520 15235 14560 15240
rect 14520 15205 14525 15235
rect 14555 15205 14560 15235
rect 14520 15200 14560 15205
rect 14600 15235 14640 15240
rect 14600 15205 14605 15235
rect 14635 15205 14640 15235
rect 14600 15200 14640 15205
rect 14680 15235 14720 15240
rect 14680 15205 14685 15235
rect 14715 15205 14720 15235
rect 14680 15200 14720 15205
rect 16760 15235 16800 15240
rect 16760 15205 16765 15235
rect 16795 15205 16800 15235
rect 16760 15200 16800 15205
rect 16840 15235 16880 15240
rect 16840 15205 16845 15235
rect 16875 15205 16880 15235
rect 16840 15200 16880 15205
rect 16920 15235 16960 15240
rect 16920 15205 16925 15235
rect 16955 15205 16960 15235
rect 16920 15200 16960 15205
rect 17000 15235 17040 15240
rect 17000 15205 17005 15235
rect 17035 15205 17040 15235
rect 17000 15200 17040 15205
rect 17080 15235 17120 15240
rect 17080 15205 17085 15235
rect 17115 15205 17120 15235
rect 17080 15200 17120 15205
rect 17160 15235 17200 15240
rect 17160 15205 17165 15235
rect 17195 15205 17200 15235
rect 17160 15200 17200 15205
rect 17240 15235 17280 15240
rect 17240 15205 17245 15235
rect 17275 15205 17280 15235
rect 17240 15200 17280 15205
rect 17320 15235 17360 15240
rect 17320 15205 17325 15235
rect 17355 15205 17360 15235
rect 17320 15200 17360 15205
rect 17400 15235 17440 15240
rect 17400 15205 17405 15235
rect 17435 15205 17440 15235
rect 17400 15200 17440 15205
rect 17480 15235 17520 15240
rect 17480 15205 17485 15235
rect 17515 15205 17520 15235
rect 17480 15200 17520 15205
rect 17560 15235 17600 15240
rect 17560 15205 17565 15235
rect 17595 15205 17600 15235
rect 17560 15200 17600 15205
rect 17640 15235 17680 15240
rect 17640 15205 17645 15235
rect 17675 15205 17680 15235
rect 17640 15200 17680 15205
rect 17720 15235 17760 15240
rect 17720 15205 17725 15235
rect 17755 15205 17760 15235
rect 17720 15200 17760 15205
rect 17800 15235 17840 15240
rect 17800 15205 17805 15235
rect 17835 15205 17840 15235
rect 17800 15200 17840 15205
rect 17880 15235 17920 15240
rect 17880 15205 17885 15235
rect 17915 15205 17920 15235
rect 17880 15200 17920 15205
rect 17960 15235 18000 15240
rect 17960 15205 17965 15235
rect 17995 15205 18000 15235
rect 17960 15200 18000 15205
rect 18040 15235 18080 15240
rect 18040 15205 18045 15235
rect 18075 15205 18080 15235
rect 18040 15200 18080 15205
rect 18120 15235 18160 15240
rect 18120 15205 18125 15235
rect 18155 15205 18160 15235
rect 18120 15200 18160 15205
rect 18200 15235 18240 15240
rect 18200 15205 18205 15235
rect 18235 15205 18240 15235
rect 18200 15200 18240 15205
rect 18280 15235 18320 15240
rect 18280 15205 18285 15235
rect 18315 15205 18320 15235
rect 18280 15200 18320 15205
rect 18360 15235 18400 15240
rect 18360 15205 18365 15235
rect 18395 15205 18400 15235
rect 18360 15200 18400 15205
rect 18440 15235 18480 15240
rect 18440 15205 18445 15235
rect 18475 15205 18480 15235
rect 18440 15200 18480 15205
rect 18520 15235 18560 15240
rect 18520 15205 18525 15235
rect 18555 15205 18560 15235
rect 18520 15200 18560 15205
rect 18600 15235 18640 15240
rect 18600 15205 18605 15235
rect 18635 15205 18640 15235
rect 18600 15200 18640 15205
rect 18680 15235 18720 15240
rect 18680 15205 18685 15235
rect 18715 15205 18720 15235
rect 18680 15200 18720 15205
rect 18760 15235 18800 15240
rect 18760 15205 18765 15235
rect 18795 15205 18800 15235
rect 18760 15200 18800 15205
rect 18840 15235 18880 15240
rect 18840 15205 18845 15235
rect 18875 15205 18880 15235
rect 18840 15200 18880 15205
rect 18920 15235 18960 15240
rect 18920 15205 18925 15235
rect 18955 15205 18960 15235
rect 18920 15200 18960 15205
rect 19000 15235 19040 15240
rect 19000 15205 19005 15235
rect 19035 15205 19040 15235
rect 19000 15200 19040 15205
rect 19080 15235 19120 15240
rect 19080 15205 19085 15235
rect 19115 15205 19120 15235
rect 19080 15200 19120 15205
rect 19160 15235 19200 15240
rect 19160 15205 19165 15235
rect 19195 15205 19200 15235
rect 19160 15200 19200 15205
rect 19240 15235 19280 15240
rect 19240 15205 19245 15235
rect 19275 15205 19280 15235
rect 19240 15200 19280 15205
rect 19320 15235 19360 15240
rect 19320 15205 19325 15235
rect 19355 15205 19360 15235
rect 19320 15200 19360 15205
rect 19400 15235 19440 15240
rect 19400 15205 19405 15235
rect 19435 15205 19440 15235
rect 19400 15200 19440 15205
rect 19480 15235 19520 15240
rect 19480 15205 19485 15235
rect 19515 15205 19520 15235
rect 19480 15200 19520 15205
rect 19560 15235 19600 15240
rect 19560 15205 19565 15235
rect 19595 15205 19600 15235
rect 19560 15200 19600 15205
rect 19640 15235 19680 15240
rect 19640 15205 19645 15235
rect 19675 15205 19680 15235
rect 19640 15200 19680 15205
rect 19720 15235 19760 15240
rect 19720 15205 19725 15235
rect 19755 15205 19760 15235
rect 19720 15200 19760 15205
rect 19800 15235 19840 15240
rect 19800 15205 19805 15235
rect 19835 15205 19840 15235
rect 19800 15200 19840 15205
rect 19880 15235 19920 15240
rect 19880 15205 19885 15235
rect 19915 15205 19920 15235
rect 19880 15200 19920 15205
rect 19960 15235 20000 15240
rect 19960 15205 19965 15235
rect 19995 15205 20000 15235
rect 19960 15200 20000 15205
rect 20040 15235 20080 15240
rect 20040 15205 20045 15235
rect 20075 15205 20080 15235
rect 20040 15200 20080 15205
rect 20120 15235 20160 15240
rect 20120 15205 20125 15235
rect 20155 15205 20160 15235
rect 20120 15200 20160 15205
rect 20200 15235 20240 15240
rect 20200 15205 20205 15235
rect 20235 15205 20240 15235
rect 20200 15200 20240 15205
rect 20280 15235 20320 15240
rect 20280 15205 20285 15235
rect 20315 15205 20320 15235
rect 20280 15200 20320 15205
rect 20360 15235 20400 15240
rect 20360 15205 20365 15235
rect 20395 15205 20400 15235
rect 20360 15200 20400 15205
rect 20440 15235 20480 15240
rect 20440 15205 20445 15235
rect 20475 15205 20480 15235
rect 20440 15200 20480 15205
rect 20520 15235 20560 15240
rect 20520 15205 20525 15235
rect 20555 15205 20560 15235
rect 20520 15200 20560 15205
rect 20600 15235 20640 15240
rect 20600 15205 20605 15235
rect 20635 15205 20640 15235
rect 20600 15200 20640 15205
rect 20680 15235 20720 15240
rect 20680 15205 20685 15235
rect 20715 15205 20720 15235
rect 20680 15200 20720 15205
rect 20760 15235 20800 15240
rect 20760 15205 20765 15235
rect 20795 15205 20800 15235
rect 20760 15200 20800 15205
rect 20840 15235 20880 15240
rect 20840 15205 20845 15235
rect 20875 15205 20880 15235
rect 20840 15200 20880 15205
rect 20920 15235 20960 15240
rect 20920 15205 20925 15235
rect 20955 15205 20960 15235
rect 20920 15200 20960 15205
rect 0 15155 40 15160
rect 0 15125 5 15155
rect 35 15125 40 15155
rect 0 15120 40 15125
rect 80 15155 120 15160
rect 80 15125 85 15155
rect 115 15125 120 15155
rect 80 15120 120 15125
rect 160 15155 200 15160
rect 160 15125 165 15155
rect 195 15125 200 15155
rect 160 15120 200 15125
rect 240 15155 280 15160
rect 240 15125 245 15155
rect 275 15125 280 15155
rect 240 15120 280 15125
rect 320 15155 360 15160
rect 320 15125 325 15155
rect 355 15125 360 15155
rect 320 15120 360 15125
rect 400 15155 440 15160
rect 400 15125 405 15155
rect 435 15125 440 15155
rect 400 15120 440 15125
rect 480 15155 520 15160
rect 480 15125 485 15155
rect 515 15125 520 15155
rect 480 15120 520 15125
rect 560 15155 600 15160
rect 560 15125 565 15155
rect 595 15125 600 15155
rect 560 15120 600 15125
rect 640 15155 680 15160
rect 640 15125 645 15155
rect 675 15125 680 15155
rect 640 15120 680 15125
rect 720 15155 760 15160
rect 720 15125 725 15155
rect 755 15125 760 15155
rect 720 15120 760 15125
rect 800 15155 840 15160
rect 800 15125 805 15155
rect 835 15125 840 15155
rect 800 15120 840 15125
rect 880 15155 920 15160
rect 880 15125 885 15155
rect 915 15125 920 15155
rect 880 15120 920 15125
rect 960 15155 1000 15160
rect 960 15125 965 15155
rect 995 15125 1000 15155
rect 960 15120 1000 15125
rect 1040 15155 1080 15160
rect 1040 15125 1045 15155
rect 1075 15125 1080 15155
rect 1040 15120 1080 15125
rect 1120 15155 1160 15160
rect 1120 15125 1125 15155
rect 1155 15125 1160 15155
rect 1120 15120 1160 15125
rect 1200 15155 1240 15160
rect 1200 15125 1205 15155
rect 1235 15125 1240 15155
rect 1200 15120 1240 15125
rect 1280 15155 1320 15160
rect 1280 15125 1285 15155
rect 1315 15125 1320 15155
rect 1280 15120 1320 15125
rect 1360 15155 1400 15160
rect 1360 15125 1365 15155
rect 1395 15125 1400 15155
rect 1360 15120 1400 15125
rect 1440 15155 1480 15160
rect 1440 15125 1445 15155
rect 1475 15125 1480 15155
rect 1440 15120 1480 15125
rect 1520 15155 1560 15160
rect 1520 15125 1525 15155
rect 1555 15125 1560 15155
rect 1520 15120 1560 15125
rect 1600 15155 1640 15160
rect 1600 15125 1605 15155
rect 1635 15125 1640 15155
rect 1600 15120 1640 15125
rect 1680 15155 1720 15160
rect 1680 15125 1685 15155
rect 1715 15125 1720 15155
rect 1680 15120 1720 15125
rect 1760 15155 1800 15160
rect 1760 15125 1765 15155
rect 1795 15125 1800 15155
rect 1760 15120 1800 15125
rect 1840 15155 1880 15160
rect 1840 15125 1845 15155
rect 1875 15125 1880 15155
rect 1840 15120 1880 15125
rect 1920 15155 1960 15160
rect 1920 15125 1925 15155
rect 1955 15125 1960 15155
rect 1920 15120 1960 15125
rect 2000 15155 2040 15160
rect 2000 15125 2005 15155
rect 2035 15125 2040 15155
rect 2000 15120 2040 15125
rect 2080 15155 2120 15160
rect 2080 15125 2085 15155
rect 2115 15125 2120 15155
rect 2080 15120 2120 15125
rect 2160 15155 2200 15160
rect 2160 15125 2165 15155
rect 2195 15125 2200 15155
rect 2160 15120 2200 15125
rect 2240 15155 2280 15160
rect 2240 15125 2245 15155
rect 2275 15125 2280 15155
rect 2240 15120 2280 15125
rect 2320 15155 2360 15160
rect 2320 15125 2325 15155
rect 2355 15125 2360 15155
rect 2320 15120 2360 15125
rect 2400 15155 2440 15160
rect 2400 15125 2405 15155
rect 2435 15125 2440 15155
rect 2400 15120 2440 15125
rect 2480 15155 2520 15160
rect 2480 15125 2485 15155
rect 2515 15125 2520 15155
rect 2480 15120 2520 15125
rect 2560 15155 2600 15160
rect 2560 15125 2565 15155
rect 2595 15125 2600 15155
rect 2560 15120 2600 15125
rect 2640 15155 2680 15160
rect 2640 15125 2645 15155
rect 2675 15125 2680 15155
rect 2640 15120 2680 15125
rect 2720 15155 2760 15160
rect 2720 15125 2725 15155
rect 2755 15125 2760 15155
rect 2720 15120 2760 15125
rect 2800 15155 2840 15160
rect 2800 15125 2805 15155
rect 2835 15125 2840 15155
rect 2800 15120 2840 15125
rect 2880 15155 2920 15160
rect 2880 15125 2885 15155
rect 2915 15125 2920 15155
rect 2880 15120 2920 15125
rect 2960 15155 3000 15160
rect 2960 15125 2965 15155
rect 2995 15125 3000 15155
rect 2960 15120 3000 15125
rect 3040 15155 3080 15160
rect 3040 15125 3045 15155
rect 3075 15125 3080 15155
rect 3040 15120 3080 15125
rect 3120 15155 3160 15160
rect 3120 15125 3125 15155
rect 3155 15125 3160 15155
rect 3120 15120 3160 15125
rect 3200 15155 3240 15160
rect 3200 15125 3205 15155
rect 3235 15125 3240 15155
rect 3200 15120 3240 15125
rect 3280 15155 3320 15160
rect 3280 15125 3285 15155
rect 3315 15125 3320 15155
rect 3280 15120 3320 15125
rect 3360 15155 3400 15160
rect 3360 15125 3365 15155
rect 3395 15125 3400 15155
rect 3360 15120 3400 15125
rect 3440 15155 3480 15160
rect 3440 15125 3445 15155
rect 3475 15125 3480 15155
rect 3440 15120 3480 15125
rect 3520 15155 3560 15160
rect 3520 15125 3525 15155
rect 3555 15125 3560 15155
rect 3520 15120 3560 15125
rect 3600 15155 3640 15160
rect 3600 15125 3605 15155
rect 3635 15125 3640 15155
rect 3600 15120 3640 15125
rect 3680 15155 3720 15160
rect 3680 15125 3685 15155
rect 3715 15125 3720 15155
rect 3680 15120 3720 15125
rect 3760 15155 3800 15160
rect 3760 15125 3765 15155
rect 3795 15125 3800 15155
rect 3760 15120 3800 15125
rect 3840 15155 3880 15160
rect 3840 15125 3845 15155
rect 3875 15125 3880 15155
rect 3840 15120 3880 15125
rect 3920 15155 3960 15160
rect 3920 15125 3925 15155
rect 3955 15125 3960 15155
rect 3920 15120 3960 15125
rect 4000 15155 4040 15160
rect 4000 15125 4005 15155
rect 4035 15125 4040 15155
rect 4000 15120 4040 15125
rect 4080 15155 4120 15160
rect 4080 15125 4085 15155
rect 4115 15125 4120 15155
rect 4080 15120 4120 15125
rect 4160 15155 4200 15160
rect 4160 15125 4165 15155
rect 4195 15125 4200 15155
rect 4160 15120 4200 15125
rect 6240 15155 6280 15160
rect 6240 15125 6245 15155
rect 6275 15125 6280 15155
rect 6240 15120 6280 15125
rect 6320 15155 6360 15160
rect 6320 15125 6325 15155
rect 6355 15125 6360 15155
rect 6320 15120 6360 15125
rect 6400 15155 6440 15160
rect 6400 15125 6405 15155
rect 6435 15125 6440 15155
rect 6400 15120 6440 15125
rect 6480 15155 6520 15160
rect 6480 15125 6485 15155
rect 6515 15125 6520 15155
rect 6480 15120 6520 15125
rect 6560 15155 6600 15160
rect 6560 15125 6565 15155
rect 6595 15125 6600 15155
rect 6560 15120 6600 15125
rect 6640 15155 6680 15160
rect 6640 15125 6645 15155
rect 6675 15125 6680 15155
rect 6640 15120 6680 15125
rect 6720 15155 6760 15160
rect 6720 15125 6725 15155
rect 6755 15125 6760 15155
rect 6720 15120 6760 15125
rect 6800 15155 6840 15160
rect 6800 15125 6805 15155
rect 6835 15125 6840 15155
rect 6800 15120 6840 15125
rect 6880 15155 6920 15160
rect 6880 15125 6885 15155
rect 6915 15125 6920 15155
rect 6880 15120 6920 15125
rect 6960 15155 7000 15160
rect 6960 15125 6965 15155
rect 6995 15125 7000 15155
rect 6960 15120 7000 15125
rect 7040 15155 7080 15160
rect 7040 15125 7045 15155
rect 7075 15125 7080 15155
rect 7040 15120 7080 15125
rect 7120 15155 7160 15160
rect 7120 15125 7125 15155
rect 7155 15125 7160 15155
rect 7120 15120 7160 15125
rect 7200 15155 7240 15160
rect 7200 15125 7205 15155
rect 7235 15125 7240 15155
rect 7200 15120 7240 15125
rect 7280 15155 7320 15160
rect 7280 15125 7285 15155
rect 7315 15125 7320 15155
rect 7280 15120 7320 15125
rect 7360 15155 7400 15160
rect 7360 15125 7365 15155
rect 7395 15125 7400 15155
rect 7360 15120 7400 15125
rect 7440 15155 7480 15160
rect 7440 15125 7445 15155
rect 7475 15125 7480 15155
rect 7440 15120 7480 15125
rect 7520 15155 7560 15160
rect 7520 15125 7525 15155
rect 7555 15125 7560 15155
rect 7520 15120 7560 15125
rect 7600 15155 7640 15160
rect 7600 15125 7605 15155
rect 7635 15125 7640 15155
rect 7600 15120 7640 15125
rect 7680 15155 7720 15160
rect 7680 15125 7685 15155
rect 7715 15125 7720 15155
rect 7680 15120 7720 15125
rect 7760 15155 7800 15160
rect 7760 15125 7765 15155
rect 7795 15125 7800 15155
rect 7760 15120 7800 15125
rect 7840 15155 7880 15160
rect 7840 15125 7845 15155
rect 7875 15125 7880 15155
rect 7840 15120 7880 15125
rect 7920 15155 7960 15160
rect 7920 15125 7925 15155
rect 7955 15125 7960 15155
rect 7920 15120 7960 15125
rect 8000 15155 8040 15160
rect 8000 15125 8005 15155
rect 8035 15125 8040 15155
rect 8000 15120 8040 15125
rect 8080 15155 8120 15160
rect 8080 15125 8085 15155
rect 8115 15125 8120 15155
rect 8080 15120 8120 15125
rect 8160 15155 8200 15160
rect 8160 15125 8165 15155
rect 8195 15125 8200 15155
rect 8160 15120 8200 15125
rect 8240 15155 8280 15160
rect 8240 15125 8245 15155
rect 8275 15125 8280 15155
rect 8240 15120 8280 15125
rect 8320 15155 8360 15160
rect 8320 15125 8325 15155
rect 8355 15125 8360 15155
rect 8320 15120 8360 15125
rect 8400 15155 8440 15160
rect 8400 15125 8405 15155
rect 8435 15125 8440 15155
rect 8400 15120 8440 15125
rect 8480 15155 8520 15160
rect 8480 15125 8485 15155
rect 8515 15125 8520 15155
rect 8480 15120 8520 15125
rect 8560 15155 8600 15160
rect 8560 15125 8565 15155
rect 8595 15125 8600 15155
rect 8560 15120 8600 15125
rect 8640 15155 8680 15160
rect 8640 15125 8645 15155
rect 8675 15125 8680 15155
rect 8640 15120 8680 15125
rect 8720 15155 8760 15160
rect 8720 15125 8725 15155
rect 8755 15125 8760 15155
rect 8720 15120 8760 15125
rect 8800 15155 8840 15160
rect 8800 15125 8805 15155
rect 8835 15125 8840 15155
rect 8800 15120 8840 15125
rect 8880 15155 8920 15160
rect 8880 15125 8885 15155
rect 8915 15125 8920 15155
rect 8880 15120 8920 15125
rect 8960 15155 9000 15160
rect 8960 15125 8965 15155
rect 8995 15125 9000 15155
rect 8960 15120 9000 15125
rect 9040 15155 9080 15160
rect 9040 15125 9045 15155
rect 9075 15125 9080 15155
rect 9040 15120 9080 15125
rect 9120 15155 9160 15160
rect 9120 15125 9125 15155
rect 9155 15125 9160 15155
rect 9120 15120 9160 15125
rect 9200 15155 9240 15160
rect 9200 15125 9205 15155
rect 9235 15125 9240 15155
rect 9200 15120 9240 15125
rect 9280 15155 9320 15160
rect 9280 15125 9285 15155
rect 9315 15125 9320 15155
rect 9280 15120 9320 15125
rect 9360 15155 9400 15160
rect 9360 15125 9365 15155
rect 9395 15125 9400 15155
rect 9360 15120 9400 15125
rect 9440 15155 9480 15160
rect 9440 15125 9445 15155
rect 9475 15125 9480 15155
rect 9440 15120 9480 15125
rect 11560 15155 11600 15160
rect 11560 15125 11565 15155
rect 11595 15125 11600 15155
rect 11560 15120 11600 15125
rect 11640 15155 11680 15160
rect 11640 15125 11645 15155
rect 11675 15125 11680 15155
rect 11640 15120 11680 15125
rect 11720 15155 11760 15160
rect 11720 15125 11725 15155
rect 11755 15125 11760 15155
rect 11720 15120 11760 15125
rect 11800 15155 11840 15160
rect 11800 15125 11805 15155
rect 11835 15125 11840 15155
rect 11800 15120 11840 15125
rect 11880 15155 11920 15160
rect 11880 15125 11885 15155
rect 11915 15125 11920 15155
rect 11880 15120 11920 15125
rect 11960 15155 12000 15160
rect 11960 15125 11965 15155
rect 11995 15125 12000 15155
rect 11960 15120 12000 15125
rect 12040 15155 12080 15160
rect 12040 15125 12045 15155
rect 12075 15125 12080 15155
rect 12040 15120 12080 15125
rect 12120 15155 12160 15160
rect 12120 15125 12125 15155
rect 12155 15125 12160 15155
rect 12120 15120 12160 15125
rect 12200 15155 12240 15160
rect 12200 15125 12205 15155
rect 12235 15125 12240 15155
rect 12200 15120 12240 15125
rect 12280 15155 12320 15160
rect 12280 15125 12285 15155
rect 12315 15125 12320 15155
rect 12280 15120 12320 15125
rect 12360 15155 12400 15160
rect 12360 15125 12365 15155
rect 12395 15125 12400 15155
rect 12360 15120 12400 15125
rect 12440 15155 12480 15160
rect 12440 15125 12445 15155
rect 12475 15125 12480 15155
rect 12440 15120 12480 15125
rect 12520 15155 12560 15160
rect 12520 15125 12525 15155
rect 12555 15125 12560 15155
rect 12520 15120 12560 15125
rect 12600 15155 12640 15160
rect 12600 15125 12605 15155
rect 12635 15125 12640 15155
rect 12600 15120 12640 15125
rect 12680 15155 12720 15160
rect 12680 15125 12685 15155
rect 12715 15125 12720 15155
rect 12680 15120 12720 15125
rect 12760 15155 12800 15160
rect 12760 15125 12765 15155
rect 12795 15125 12800 15155
rect 12760 15120 12800 15125
rect 12840 15155 12880 15160
rect 12840 15125 12845 15155
rect 12875 15125 12880 15155
rect 12840 15120 12880 15125
rect 12920 15155 12960 15160
rect 12920 15125 12925 15155
rect 12955 15125 12960 15155
rect 12920 15120 12960 15125
rect 13000 15155 13040 15160
rect 13000 15125 13005 15155
rect 13035 15125 13040 15155
rect 13000 15120 13040 15125
rect 13080 15155 13120 15160
rect 13080 15125 13085 15155
rect 13115 15125 13120 15155
rect 13080 15120 13120 15125
rect 13160 15155 13200 15160
rect 13160 15125 13165 15155
rect 13195 15125 13200 15155
rect 13160 15120 13200 15125
rect 13240 15155 13280 15160
rect 13240 15125 13245 15155
rect 13275 15125 13280 15155
rect 13240 15120 13280 15125
rect 13320 15155 13360 15160
rect 13320 15125 13325 15155
rect 13355 15125 13360 15155
rect 13320 15120 13360 15125
rect 13400 15155 13440 15160
rect 13400 15125 13405 15155
rect 13435 15125 13440 15155
rect 13400 15120 13440 15125
rect 13480 15155 13520 15160
rect 13480 15125 13485 15155
rect 13515 15125 13520 15155
rect 13480 15120 13520 15125
rect 13560 15155 13600 15160
rect 13560 15125 13565 15155
rect 13595 15125 13600 15155
rect 13560 15120 13600 15125
rect 13640 15155 13680 15160
rect 13640 15125 13645 15155
rect 13675 15125 13680 15155
rect 13640 15120 13680 15125
rect 13720 15155 13760 15160
rect 13720 15125 13725 15155
rect 13755 15125 13760 15155
rect 13720 15120 13760 15125
rect 13800 15155 13840 15160
rect 13800 15125 13805 15155
rect 13835 15125 13840 15155
rect 13800 15120 13840 15125
rect 13880 15155 13920 15160
rect 13880 15125 13885 15155
rect 13915 15125 13920 15155
rect 13880 15120 13920 15125
rect 13960 15155 14000 15160
rect 13960 15125 13965 15155
rect 13995 15125 14000 15155
rect 13960 15120 14000 15125
rect 14040 15155 14080 15160
rect 14040 15125 14045 15155
rect 14075 15125 14080 15155
rect 14040 15120 14080 15125
rect 14120 15155 14160 15160
rect 14120 15125 14125 15155
rect 14155 15125 14160 15155
rect 14120 15120 14160 15125
rect 14200 15155 14240 15160
rect 14200 15125 14205 15155
rect 14235 15125 14240 15155
rect 14200 15120 14240 15125
rect 14280 15155 14320 15160
rect 14280 15125 14285 15155
rect 14315 15125 14320 15155
rect 14280 15120 14320 15125
rect 14360 15155 14400 15160
rect 14360 15125 14365 15155
rect 14395 15125 14400 15155
rect 14360 15120 14400 15125
rect 14440 15155 14480 15160
rect 14440 15125 14445 15155
rect 14475 15125 14480 15155
rect 14440 15120 14480 15125
rect 14520 15155 14560 15160
rect 14520 15125 14525 15155
rect 14555 15125 14560 15155
rect 14520 15120 14560 15125
rect 14600 15155 14640 15160
rect 14600 15125 14605 15155
rect 14635 15125 14640 15155
rect 14600 15120 14640 15125
rect 14680 15155 14720 15160
rect 14680 15125 14685 15155
rect 14715 15125 14720 15155
rect 14680 15120 14720 15125
rect 16760 15155 16800 15160
rect 16760 15125 16765 15155
rect 16795 15125 16800 15155
rect 16760 15120 16800 15125
rect 16840 15155 16880 15160
rect 16840 15125 16845 15155
rect 16875 15125 16880 15155
rect 16840 15120 16880 15125
rect 16920 15155 16960 15160
rect 16920 15125 16925 15155
rect 16955 15125 16960 15155
rect 16920 15120 16960 15125
rect 17000 15155 17040 15160
rect 17000 15125 17005 15155
rect 17035 15125 17040 15155
rect 17000 15120 17040 15125
rect 17080 15155 17120 15160
rect 17080 15125 17085 15155
rect 17115 15125 17120 15155
rect 17080 15120 17120 15125
rect 17160 15155 17200 15160
rect 17160 15125 17165 15155
rect 17195 15125 17200 15155
rect 17160 15120 17200 15125
rect 17240 15155 17280 15160
rect 17240 15125 17245 15155
rect 17275 15125 17280 15155
rect 17240 15120 17280 15125
rect 17320 15155 17360 15160
rect 17320 15125 17325 15155
rect 17355 15125 17360 15155
rect 17320 15120 17360 15125
rect 17400 15155 17440 15160
rect 17400 15125 17405 15155
rect 17435 15125 17440 15155
rect 17400 15120 17440 15125
rect 17480 15155 17520 15160
rect 17480 15125 17485 15155
rect 17515 15125 17520 15155
rect 17480 15120 17520 15125
rect 17560 15155 17600 15160
rect 17560 15125 17565 15155
rect 17595 15125 17600 15155
rect 17560 15120 17600 15125
rect 17640 15155 17680 15160
rect 17640 15125 17645 15155
rect 17675 15125 17680 15155
rect 17640 15120 17680 15125
rect 17720 15155 17760 15160
rect 17720 15125 17725 15155
rect 17755 15125 17760 15155
rect 17720 15120 17760 15125
rect 17800 15155 17840 15160
rect 17800 15125 17805 15155
rect 17835 15125 17840 15155
rect 17800 15120 17840 15125
rect 17880 15155 17920 15160
rect 17880 15125 17885 15155
rect 17915 15125 17920 15155
rect 17880 15120 17920 15125
rect 17960 15155 18000 15160
rect 17960 15125 17965 15155
rect 17995 15125 18000 15155
rect 17960 15120 18000 15125
rect 18040 15155 18080 15160
rect 18040 15125 18045 15155
rect 18075 15125 18080 15155
rect 18040 15120 18080 15125
rect 18120 15155 18160 15160
rect 18120 15125 18125 15155
rect 18155 15125 18160 15155
rect 18120 15120 18160 15125
rect 18200 15155 18240 15160
rect 18200 15125 18205 15155
rect 18235 15125 18240 15155
rect 18200 15120 18240 15125
rect 18280 15155 18320 15160
rect 18280 15125 18285 15155
rect 18315 15125 18320 15155
rect 18280 15120 18320 15125
rect 18360 15155 18400 15160
rect 18360 15125 18365 15155
rect 18395 15125 18400 15155
rect 18360 15120 18400 15125
rect 18440 15155 18480 15160
rect 18440 15125 18445 15155
rect 18475 15125 18480 15155
rect 18440 15120 18480 15125
rect 18520 15155 18560 15160
rect 18520 15125 18525 15155
rect 18555 15125 18560 15155
rect 18520 15120 18560 15125
rect 18600 15155 18640 15160
rect 18600 15125 18605 15155
rect 18635 15125 18640 15155
rect 18600 15120 18640 15125
rect 18680 15155 18720 15160
rect 18680 15125 18685 15155
rect 18715 15125 18720 15155
rect 18680 15120 18720 15125
rect 18760 15155 18800 15160
rect 18760 15125 18765 15155
rect 18795 15125 18800 15155
rect 18760 15120 18800 15125
rect 18840 15155 18880 15160
rect 18840 15125 18845 15155
rect 18875 15125 18880 15155
rect 18840 15120 18880 15125
rect 18920 15155 18960 15160
rect 18920 15125 18925 15155
rect 18955 15125 18960 15155
rect 18920 15120 18960 15125
rect 19000 15155 19040 15160
rect 19000 15125 19005 15155
rect 19035 15125 19040 15155
rect 19000 15120 19040 15125
rect 19080 15155 19120 15160
rect 19080 15125 19085 15155
rect 19115 15125 19120 15155
rect 19080 15120 19120 15125
rect 19160 15155 19200 15160
rect 19160 15125 19165 15155
rect 19195 15125 19200 15155
rect 19160 15120 19200 15125
rect 19240 15155 19280 15160
rect 19240 15125 19245 15155
rect 19275 15125 19280 15155
rect 19240 15120 19280 15125
rect 19320 15155 19360 15160
rect 19320 15125 19325 15155
rect 19355 15125 19360 15155
rect 19320 15120 19360 15125
rect 19400 15155 19440 15160
rect 19400 15125 19405 15155
rect 19435 15125 19440 15155
rect 19400 15120 19440 15125
rect 19480 15155 19520 15160
rect 19480 15125 19485 15155
rect 19515 15125 19520 15155
rect 19480 15120 19520 15125
rect 19560 15155 19600 15160
rect 19560 15125 19565 15155
rect 19595 15125 19600 15155
rect 19560 15120 19600 15125
rect 19640 15155 19680 15160
rect 19640 15125 19645 15155
rect 19675 15125 19680 15155
rect 19640 15120 19680 15125
rect 19720 15155 19760 15160
rect 19720 15125 19725 15155
rect 19755 15125 19760 15155
rect 19720 15120 19760 15125
rect 19800 15155 19840 15160
rect 19800 15125 19805 15155
rect 19835 15125 19840 15155
rect 19800 15120 19840 15125
rect 19880 15155 19920 15160
rect 19880 15125 19885 15155
rect 19915 15125 19920 15155
rect 19880 15120 19920 15125
rect 19960 15155 20000 15160
rect 19960 15125 19965 15155
rect 19995 15125 20000 15155
rect 19960 15120 20000 15125
rect 20040 15155 20080 15160
rect 20040 15125 20045 15155
rect 20075 15125 20080 15155
rect 20040 15120 20080 15125
rect 20120 15155 20160 15160
rect 20120 15125 20125 15155
rect 20155 15125 20160 15155
rect 20120 15120 20160 15125
rect 20200 15155 20240 15160
rect 20200 15125 20205 15155
rect 20235 15125 20240 15155
rect 20200 15120 20240 15125
rect 20280 15155 20320 15160
rect 20280 15125 20285 15155
rect 20315 15125 20320 15155
rect 20280 15120 20320 15125
rect 20360 15155 20400 15160
rect 20360 15125 20365 15155
rect 20395 15125 20400 15155
rect 20360 15120 20400 15125
rect 20440 15155 20480 15160
rect 20440 15125 20445 15155
rect 20475 15125 20480 15155
rect 20440 15120 20480 15125
rect 20520 15155 20560 15160
rect 20520 15125 20525 15155
rect 20555 15125 20560 15155
rect 20520 15120 20560 15125
rect 20600 15155 20640 15160
rect 20600 15125 20605 15155
rect 20635 15125 20640 15155
rect 20600 15120 20640 15125
rect 20680 15155 20720 15160
rect 20680 15125 20685 15155
rect 20715 15125 20720 15155
rect 20680 15120 20720 15125
rect 20760 15155 20800 15160
rect 20760 15125 20765 15155
rect 20795 15125 20800 15155
rect 20760 15120 20800 15125
rect 20840 15155 20880 15160
rect 20840 15125 20845 15155
rect 20875 15125 20880 15155
rect 20840 15120 20880 15125
rect 20920 15155 20960 15160
rect 20920 15125 20925 15155
rect 20955 15125 20960 15155
rect 20920 15120 20960 15125
rect 0 14995 40 15000
rect 0 14965 5 14995
rect 35 14965 40 14995
rect 0 14960 40 14965
rect 80 14995 120 15000
rect 80 14965 85 14995
rect 115 14965 120 14995
rect 80 14960 120 14965
rect 160 14995 200 15000
rect 160 14965 165 14995
rect 195 14965 200 14995
rect 160 14960 200 14965
rect 240 14995 280 15000
rect 240 14965 245 14995
rect 275 14965 280 14995
rect 240 14960 280 14965
rect 320 14995 360 15000
rect 320 14965 325 14995
rect 355 14965 360 14995
rect 320 14960 360 14965
rect 400 14995 440 15000
rect 400 14965 405 14995
rect 435 14965 440 14995
rect 400 14960 440 14965
rect 480 14995 520 15000
rect 480 14965 485 14995
rect 515 14965 520 14995
rect 480 14960 520 14965
rect 560 14995 600 15000
rect 560 14965 565 14995
rect 595 14965 600 14995
rect 560 14960 600 14965
rect 640 14995 680 15000
rect 640 14965 645 14995
rect 675 14965 680 14995
rect 640 14960 680 14965
rect 720 14995 760 15000
rect 720 14965 725 14995
rect 755 14965 760 14995
rect 720 14960 760 14965
rect 800 14995 840 15000
rect 800 14965 805 14995
rect 835 14965 840 14995
rect 800 14960 840 14965
rect 880 14995 920 15000
rect 880 14965 885 14995
rect 915 14965 920 14995
rect 880 14960 920 14965
rect 960 14995 1000 15000
rect 960 14965 965 14995
rect 995 14965 1000 14995
rect 960 14960 1000 14965
rect 1040 14995 1080 15000
rect 1040 14965 1045 14995
rect 1075 14965 1080 14995
rect 1040 14960 1080 14965
rect 1120 14995 1160 15000
rect 1120 14965 1125 14995
rect 1155 14965 1160 14995
rect 1120 14960 1160 14965
rect 1200 14995 1240 15000
rect 1200 14965 1205 14995
rect 1235 14965 1240 14995
rect 1200 14960 1240 14965
rect 1280 14995 1320 15000
rect 1280 14965 1285 14995
rect 1315 14965 1320 14995
rect 1280 14960 1320 14965
rect 1360 14995 1400 15000
rect 1360 14965 1365 14995
rect 1395 14965 1400 14995
rect 1360 14960 1400 14965
rect 1440 14995 1480 15000
rect 1440 14965 1445 14995
rect 1475 14965 1480 14995
rect 1440 14960 1480 14965
rect 1520 14995 1560 15000
rect 1520 14965 1525 14995
rect 1555 14965 1560 14995
rect 1520 14960 1560 14965
rect 1600 14995 1640 15000
rect 1600 14965 1605 14995
rect 1635 14965 1640 14995
rect 1600 14960 1640 14965
rect 1680 14995 1720 15000
rect 1680 14965 1685 14995
rect 1715 14965 1720 14995
rect 1680 14960 1720 14965
rect 1760 14995 1800 15000
rect 1760 14965 1765 14995
rect 1795 14965 1800 14995
rect 1760 14960 1800 14965
rect 1840 14995 1880 15000
rect 1840 14965 1845 14995
rect 1875 14965 1880 14995
rect 1840 14960 1880 14965
rect 1920 14995 1960 15000
rect 1920 14965 1925 14995
rect 1955 14965 1960 14995
rect 1920 14960 1960 14965
rect 2000 14995 2040 15000
rect 2000 14965 2005 14995
rect 2035 14965 2040 14995
rect 2000 14960 2040 14965
rect 2080 14995 2120 15000
rect 2080 14965 2085 14995
rect 2115 14965 2120 14995
rect 2080 14960 2120 14965
rect 2160 14995 2200 15000
rect 2160 14965 2165 14995
rect 2195 14965 2200 14995
rect 2160 14960 2200 14965
rect 2240 14995 2280 15000
rect 2240 14965 2245 14995
rect 2275 14965 2280 14995
rect 2240 14960 2280 14965
rect 2320 14995 2360 15000
rect 2320 14965 2325 14995
rect 2355 14965 2360 14995
rect 2320 14960 2360 14965
rect 2400 14995 2440 15000
rect 2400 14965 2405 14995
rect 2435 14965 2440 14995
rect 2400 14960 2440 14965
rect 2480 14995 2520 15000
rect 2480 14965 2485 14995
rect 2515 14965 2520 14995
rect 2480 14960 2520 14965
rect 2560 14995 2600 15000
rect 2560 14965 2565 14995
rect 2595 14965 2600 14995
rect 2560 14960 2600 14965
rect 2640 14995 2680 15000
rect 2640 14965 2645 14995
rect 2675 14965 2680 14995
rect 2640 14960 2680 14965
rect 2720 14995 2760 15000
rect 2720 14965 2725 14995
rect 2755 14965 2760 14995
rect 2720 14960 2760 14965
rect 2800 14995 2840 15000
rect 2800 14965 2805 14995
rect 2835 14965 2840 14995
rect 2800 14960 2840 14965
rect 2880 14995 2920 15000
rect 2880 14965 2885 14995
rect 2915 14965 2920 14995
rect 2880 14960 2920 14965
rect 2960 14995 3000 15000
rect 2960 14965 2965 14995
rect 2995 14965 3000 14995
rect 2960 14960 3000 14965
rect 3040 14995 3080 15000
rect 3040 14965 3045 14995
rect 3075 14965 3080 14995
rect 3040 14960 3080 14965
rect 3120 14995 3160 15000
rect 3120 14965 3125 14995
rect 3155 14965 3160 14995
rect 3120 14960 3160 14965
rect 3200 14995 3240 15000
rect 3200 14965 3205 14995
rect 3235 14965 3240 14995
rect 3200 14960 3240 14965
rect 3280 14995 3320 15000
rect 3280 14965 3285 14995
rect 3315 14965 3320 14995
rect 3280 14960 3320 14965
rect 3360 14995 3400 15000
rect 3360 14965 3365 14995
rect 3395 14965 3400 14995
rect 3360 14960 3400 14965
rect 3440 14995 3480 15000
rect 3440 14965 3445 14995
rect 3475 14965 3480 14995
rect 3440 14960 3480 14965
rect 3520 14995 3560 15000
rect 3520 14965 3525 14995
rect 3555 14965 3560 14995
rect 3520 14960 3560 14965
rect 3600 14995 3640 15000
rect 3600 14965 3605 14995
rect 3635 14965 3640 14995
rect 3600 14960 3640 14965
rect 3680 14995 3720 15000
rect 3680 14965 3685 14995
rect 3715 14965 3720 14995
rect 3680 14960 3720 14965
rect 3760 14995 3800 15000
rect 3760 14965 3765 14995
rect 3795 14965 3800 14995
rect 3760 14960 3800 14965
rect 3840 14995 3880 15000
rect 3840 14965 3845 14995
rect 3875 14965 3880 14995
rect 3840 14960 3880 14965
rect 3920 14995 3960 15000
rect 3920 14965 3925 14995
rect 3955 14965 3960 14995
rect 3920 14960 3960 14965
rect 4000 14995 4040 15000
rect 4000 14965 4005 14995
rect 4035 14965 4040 14995
rect 4000 14960 4040 14965
rect 4080 14995 4120 15000
rect 4080 14965 4085 14995
rect 4115 14965 4120 14995
rect 4080 14960 4120 14965
rect 4160 14995 4200 15000
rect 4160 14965 4165 14995
rect 4195 14965 4200 14995
rect 4160 14960 4200 14965
rect 6240 14995 6280 15000
rect 6240 14965 6245 14995
rect 6275 14965 6280 14995
rect 6240 14960 6280 14965
rect 6320 14995 6360 15000
rect 6320 14965 6325 14995
rect 6355 14965 6360 14995
rect 6320 14960 6360 14965
rect 6400 14995 6440 15000
rect 6400 14965 6405 14995
rect 6435 14965 6440 14995
rect 6400 14960 6440 14965
rect 6480 14995 6520 15000
rect 6480 14965 6485 14995
rect 6515 14965 6520 14995
rect 6480 14960 6520 14965
rect 6560 14995 6600 15000
rect 6560 14965 6565 14995
rect 6595 14965 6600 14995
rect 6560 14960 6600 14965
rect 6640 14995 6680 15000
rect 6640 14965 6645 14995
rect 6675 14965 6680 14995
rect 6640 14960 6680 14965
rect 6720 14995 6760 15000
rect 6720 14965 6725 14995
rect 6755 14965 6760 14995
rect 6720 14960 6760 14965
rect 6800 14995 6840 15000
rect 6800 14965 6805 14995
rect 6835 14965 6840 14995
rect 6800 14960 6840 14965
rect 6880 14995 6920 15000
rect 6880 14965 6885 14995
rect 6915 14965 6920 14995
rect 6880 14960 6920 14965
rect 6960 14995 7000 15000
rect 6960 14965 6965 14995
rect 6995 14965 7000 14995
rect 6960 14960 7000 14965
rect 7040 14995 7080 15000
rect 7040 14965 7045 14995
rect 7075 14965 7080 14995
rect 7040 14960 7080 14965
rect 7120 14995 7160 15000
rect 7120 14965 7125 14995
rect 7155 14965 7160 14995
rect 7120 14960 7160 14965
rect 7200 14995 7240 15000
rect 7200 14965 7205 14995
rect 7235 14965 7240 14995
rect 7200 14960 7240 14965
rect 7280 14995 7320 15000
rect 7280 14965 7285 14995
rect 7315 14965 7320 14995
rect 7280 14960 7320 14965
rect 7360 14995 7400 15000
rect 7360 14965 7365 14995
rect 7395 14965 7400 14995
rect 7360 14960 7400 14965
rect 7440 14995 7480 15000
rect 7440 14965 7445 14995
rect 7475 14965 7480 14995
rect 7440 14960 7480 14965
rect 7520 14995 7560 15000
rect 7520 14965 7525 14995
rect 7555 14965 7560 14995
rect 7520 14960 7560 14965
rect 7600 14995 7640 15000
rect 7600 14965 7605 14995
rect 7635 14965 7640 14995
rect 7600 14960 7640 14965
rect 7680 14995 7720 15000
rect 7680 14965 7685 14995
rect 7715 14965 7720 14995
rect 7680 14960 7720 14965
rect 7760 14995 7800 15000
rect 7760 14965 7765 14995
rect 7795 14965 7800 14995
rect 7760 14960 7800 14965
rect 7840 14995 7880 15000
rect 7840 14965 7845 14995
rect 7875 14965 7880 14995
rect 7840 14960 7880 14965
rect 7920 14995 7960 15000
rect 7920 14965 7925 14995
rect 7955 14965 7960 14995
rect 7920 14960 7960 14965
rect 8000 14995 8040 15000
rect 8000 14965 8005 14995
rect 8035 14965 8040 14995
rect 8000 14960 8040 14965
rect 8080 14995 8120 15000
rect 8080 14965 8085 14995
rect 8115 14965 8120 14995
rect 8080 14960 8120 14965
rect 8160 14995 8200 15000
rect 8160 14965 8165 14995
rect 8195 14965 8200 14995
rect 8160 14960 8200 14965
rect 8240 14995 8280 15000
rect 8240 14965 8245 14995
rect 8275 14965 8280 14995
rect 8240 14960 8280 14965
rect 8320 14995 8360 15000
rect 8320 14965 8325 14995
rect 8355 14965 8360 14995
rect 8320 14960 8360 14965
rect 8400 14995 8440 15000
rect 8400 14965 8405 14995
rect 8435 14965 8440 14995
rect 8400 14960 8440 14965
rect 8480 14995 8520 15000
rect 8480 14965 8485 14995
rect 8515 14965 8520 14995
rect 8480 14960 8520 14965
rect 8560 14995 8600 15000
rect 8560 14965 8565 14995
rect 8595 14965 8600 14995
rect 8560 14960 8600 14965
rect 8640 14995 8680 15000
rect 8640 14965 8645 14995
rect 8675 14965 8680 14995
rect 8640 14960 8680 14965
rect 8720 14995 8760 15000
rect 8720 14965 8725 14995
rect 8755 14965 8760 14995
rect 8720 14960 8760 14965
rect 8800 14995 8840 15000
rect 8800 14965 8805 14995
rect 8835 14965 8840 14995
rect 8800 14960 8840 14965
rect 8880 14995 8920 15000
rect 8880 14965 8885 14995
rect 8915 14965 8920 14995
rect 8880 14960 8920 14965
rect 8960 14995 9000 15000
rect 8960 14965 8965 14995
rect 8995 14965 9000 14995
rect 8960 14960 9000 14965
rect 9040 14995 9080 15000
rect 9040 14965 9045 14995
rect 9075 14965 9080 14995
rect 9040 14960 9080 14965
rect 9120 14995 9160 15000
rect 9120 14965 9125 14995
rect 9155 14965 9160 14995
rect 9120 14960 9160 14965
rect 9200 14995 9240 15000
rect 9200 14965 9205 14995
rect 9235 14965 9240 14995
rect 9200 14960 9240 14965
rect 9280 14995 9320 15000
rect 9280 14965 9285 14995
rect 9315 14965 9320 14995
rect 9280 14960 9320 14965
rect 9360 14995 9400 15000
rect 9360 14965 9365 14995
rect 9395 14965 9400 14995
rect 9360 14960 9400 14965
rect 9440 14995 9480 15000
rect 9440 14965 9445 14995
rect 9475 14965 9480 14995
rect 9440 14960 9480 14965
rect 11560 14995 11600 15000
rect 11560 14965 11565 14995
rect 11595 14965 11600 14995
rect 11560 14960 11600 14965
rect 11640 14995 11680 15000
rect 11640 14965 11645 14995
rect 11675 14965 11680 14995
rect 11640 14960 11680 14965
rect 11720 14995 11760 15000
rect 11720 14965 11725 14995
rect 11755 14965 11760 14995
rect 11720 14960 11760 14965
rect 11800 14995 11840 15000
rect 11800 14965 11805 14995
rect 11835 14965 11840 14995
rect 11800 14960 11840 14965
rect 11880 14995 11920 15000
rect 11880 14965 11885 14995
rect 11915 14965 11920 14995
rect 11880 14960 11920 14965
rect 11960 14995 12000 15000
rect 11960 14965 11965 14995
rect 11995 14965 12000 14995
rect 11960 14960 12000 14965
rect 12040 14995 12080 15000
rect 12040 14965 12045 14995
rect 12075 14965 12080 14995
rect 12040 14960 12080 14965
rect 12120 14995 12160 15000
rect 12120 14965 12125 14995
rect 12155 14965 12160 14995
rect 12120 14960 12160 14965
rect 12200 14995 12240 15000
rect 12200 14965 12205 14995
rect 12235 14965 12240 14995
rect 12200 14960 12240 14965
rect 12280 14995 12320 15000
rect 12280 14965 12285 14995
rect 12315 14965 12320 14995
rect 12280 14960 12320 14965
rect 12360 14995 12400 15000
rect 12360 14965 12365 14995
rect 12395 14965 12400 14995
rect 12360 14960 12400 14965
rect 12440 14995 12480 15000
rect 12440 14965 12445 14995
rect 12475 14965 12480 14995
rect 12440 14960 12480 14965
rect 12520 14995 12560 15000
rect 12520 14965 12525 14995
rect 12555 14965 12560 14995
rect 12520 14960 12560 14965
rect 12600 14995 12640 15000
rect 12600 14965 12605 14995
rect 12635 14965 12640 14995
rect 12600 14960 12640 14965
rect 12680 14995 12720 15000
rect 12680 14965 12685 14995
rect 12715 14965 12720 14995
rect 12680 14960 12720 14965
rect 12760 14995 12800 15000
rect 12760 14965 12765 14995
rect 12795 14965 12800 14995
rect 12760 14960 12800 14965
rect 12840 14995 12880 15000
rect 12840 14965 12845 14995
rect 12875 14965 12880 14995
rect 12840 14960 12880 14965
rect 12920 14995 12960 15000
rect 12920 14965 12925 14995
rect 12955 14965 12960 14995
rect 12920 14960 12960 14965
rect 13000 14995 13040 15000
rect 13000 14965 13005 14995
rect 13035 14965 13040 14995
rect 13000 14960 13040 14965
rect 13080 14995 13120 15000
rect 13080 14965 13085 14995
rect 13115 14965 13120 14995
rect 13080 14960 13120 14965
rect 13160 14995 13200 15000
rect 13160 14965 13165 14995
rect 13195 14965 13200 14995
rect 13160 14960 13200 14965
rect 13240 14995 13280 15000
rect 13240 14965 13245 14995
rect 13275 14965 13280 14995
rect 13240 14960 13280 14965
rect 13320 14995 13360 15000
rect 13320 14965 13325 14995
rect 13355 14965 13360 14995
rect 13320 14960 13360 14965
rect 13400 14995 13440 15000
rect 13400 14965 13405 14995
rect 13435 14965 13440 14995
rect 13400 14960 13440 14965
rect 13480 14995 13520 15000
rect 13480 14965 13485 14995
rect 13515 14965 13520 14995
rect 13480 14960 13520 14965
rect 13560 14995 13600 15000
rect 13560 14965 13565 14995
rect 13595 14965 13600 14995
rect 13560 14960 13600 14965
rect 13640 14995 13680 15000
rect 13640 14965 13645 14995
rect 13675 14965 13680 14995
rect 13640 14960 13680 14965
rect 13720 14995 13760 15000
rect 13720 14965 13725 14995
rect 13755 14965 13760 14995
rect 13720 14960 13760 14965
rect 13800 14995 13840 15000
rect 13800 14965 13805 14995
rect 13835 14965 13840 14995
rect 13800 14960 13840 14965
rect 13880 14995 13920 15000
rect 13880 14965 13885 14995
rect 13915 14965 13920 14995
rect 13880 14960 13920 14965
rect 13960 14995 14000 15000
rect 13960 14965 13965 14995
rect 13995 14965 14000 14995
rect 13960 14960 14000 14965
rect 14040 14995 14080 15000
rect 14040 14965 14045 14995
rect 14075 14965 14080 14995
rect 14040 14960 14080 14965
rect 14120 14995 14160 15000
rect 14120 14965 14125 14995
rect 14155 14965 14160 14995
rect 14120 14960 14160 14965
rect 14200 14995 14240 15000
rect 14200 14965 14205 14995
rect 14235 14965 14240 14995
rect 14200 14960 14240 14965
rect 14280 14995 14320 15000
rect 14280 14965 14285 14995
rect 14315 14965 14320 14995
rect 14280 14960 14320 14965
rect 14360 14995 14400 15000
rect 14360 14965 14365 14995
rect 14395 14965 14400 14995
rect 14360 14960 14400 14965
rect 14440 14995 14480 15000
rect 14440 14965 14445 14995
rect 14475 14965 14480 14995
rect 14440 14960 14480 14965
rect 14520 14995 14560 15000
rect 14520 14965 14525 14995
rect 14555 14965 14560 14995
rect 14520 14960 14560 14965
rect 14600 14995 14640 15000
rect 14600 14965 14605 14995
rect 14635 14965 14640 14995
rect 14600 14960 14640 14965
rect 14680 14995 14720 15000
rect 14680 14965 14685 14995
rect 14715 14965 14720 14995
rect 14680 14960 14720 14965
rect 16760 14995 16800 15000
rect 16760 14965 16765 14995
rect 16795 14965 16800 14995
rect 16760 14960 16800 14965
rect 16840 14995 16880 15000
rect 16840 14965 16845 14995
rect 16875 14965 16880 14995
rect 16840 14960 16880 14965
rect 16920 14995 16960 15000
rect 16920 14965 16925 14995
rect 16955 14965 16960 14995
rect 16920 14960 16960 14965
rect 17000 14995 17040 15000
rect 17000 14965 17005 14995
rect 17035 14965 17040 14995
rect 17000 14960 17040 14965
rect 17080 14995 17120 15000
rect 17080 14965 17085 14995
rect 17115 14965 17120 14995
rect 17080 14960 17120 14965
rect 17160 14995 17200 15000
rect 17160 14965 17165 14995
rect 17195 14965 17200 14995
rect 17160 14960 17200 14965
rect 17240 14995 17280 15000
rect 17240 14965 17245 14995
rect 17275 14965 17280 14995
rect 17240 14960 17280 14965
rect 17320 14995 17360 15000
rect 17320 14965 17325 14995
rect 17355 14965 17360 14995
rect 17320 14960 17360 14965
rect 17400 14995 17440 15000
rect 17400 14965 17405 14995
rect 17435 14965 17440 14995
rect 17400 14960 17440 14965
rect 17480 14995 17520 15000
rect 17480 14965 17485 14995
rect 17515 14965 17520 14995
rect 17480 14960 17520 14965
rect 17560 14995 17600 15000
rect 17560 14965 17565 14995
rect 17595 14965 17600 14995
rect 17560 14960 17600 14965
rect 17640 14995 17680 15000
rect 17640 14965 17645 14995
rect 17675 14965 17680 14995
rect 17640 14960 17680 14965
rect 17720 14995 17760 15000
rect 17720 14965 17725 14995
rect 17755 14965 17760 14995
rect 17720 14960 17760 14965
rect 17800 14995 17840 15000
rect 17800 14965 17805 14995
rect 17835 14965 17840 14995
rect 17800 14960 17840 14965
rect 17880 14995 17920 15000
rect 17880 14965 17885 14995
rect 17915 14965 17920 14995
rect 17880 14960 17920 14965
rect 17960 14995 18000 15000
rect 17960 14965 17965 14995
rect 17995 14965 18000 14995
rect 17960 14960 18000 14965
rect 18040 14995 18080 15000
rect 18040 14965 18045 14995
rect 18075 14965 18080 14995
rect 18040 14960 18080 14965
rect 18120 14995 18160 15000
rect 18120 14965 18125 14995
rect 18155 14965 18160 14995
rect 18120 14960 18160 14965
rect 18200 14995 18240 15000
rect 18200 14965 18205 14995
rect 18235 14965 18240 14995
rect 18200 14960 18240 14965
rect 18280 14995 18320 15000
rect 18280 14965 18285 14995
rect 18315 14965 18320 14995
rect 18280 14960 18320 14965
rect 18360 14995 18400 15000
rect 18360 14965 18365 14995
rect 18395 14965 18400 14995
rect 18360 14960 18400 14965
rect 18440 14995 18480 15000
rect 18440 14965 18445 14995
rect 18475 14965 18480 14995
rect 18440 14960 18480 14965
rect 18520 14995 18560 15000
rect 18520 14965 18525 14995
rect 18555 14965 18560 14995
rect 18520 14960 18560 14965
rect 18600 14995 18640 15000
rect 18600 14965 18605 14995
rect 18635 14965 18640 14995
rect 18600 14960 18640 14965
rect 18680 14995 18720 15000
rect 18680 14965 18685 14995
rect 18715 14965 18720 14995
rect 18680 14960 18720 14965
rect 18760 14995 18800 15000
rect 18760 14965 18765 14995
rect 18795 14965 18800 14995
rect 18760 14960 18800 14965
rect 18840 14995 18880 15000
rect 18840 14965 18845 14995
rect 18875 14965 18880 14995
rect 18840 14960 18880 14965
rect 18920 14995 18960 15000
rect 18920 14965 18925 14995
rect 18955 14965 18960 14995
rect 18920 14960 18960 14965
rect 19000 14995 19040 15000
rect 19000 14965 19005 14995
rect 19035 14965 19040 14995
rect 19000 14960 19040 14965
rect 19080 14995 19120 15000
rect 19080 14965 19085 14995
rect 19115 14965 19120 14995
rect 19080 14960 19120 14965
rect 19160 14995 19200 15000
rect 19160 14965 19165 14995
rect 19195 14965 19200 14995
rect 19160 14960 19200 14965
rect 19240 14995 19280 15000
rect 19240 14965 19245 14995
rect 19275 14965 19280 14995
rect 19240 14960 19280 14965
rect 19320 14995 19360 15000
rect 19320 14965 19325 14995
rect 19355 14965 19360 14995
rect 19320 14960 19360 14965
rect 19400 14995 19440 15000
rect 19400 14965 19405 14995
rect 19435 14965 19440 14995
rect 19400 14960 19440 14965
rect 19480 14995 19520 15000
rect 19480 14965 19485 14995
rect 19515 14965 19520 14995
rect 19480 14960 19520 14965
rect 19560 14995 19600 15000
rect 19560 14965 19565 14995
rect 19595 14965 19600 14995
rect 19560 14960 19600 14965
rect 19640 14995 19680 15000
rect 19640 14965 19645 14995
rect 19675 14965 19680 14995
rect 19640 14960 19680 14965
rect 19720 14995 19760 15000
rect 19720 14965 19725 14995
rect 19755 14965 19760 14995
rect 19720 14960 19760 14965
rect 19800 14995 19840 15000
rect 19800 14965 19805 14995
rect 19835 14965 19840 14995
rect 19800 14960 19840 14965
rect 19880 14995 19920 15000
rect 19880 14965 19885 14995
rect 19915 14965 19920 14995
rect 19880 14960 19920 14965
rect 19960 14995 20000 15000
rect 19960 14965 19965 14995
rect 19995 14965 20000 14995
rect 19960 14960 20000 14965
rect 20040 14995 20080 15000
rect 20040 14965 20045 14995
rect 20075 14965 20080 14995
rect 20040 14960 20080 14965
rect 20120 14995 20160 15000
rect 20120 14965 20125 14995
rect 20155 14965 20160 14995
rect 20120 14960 20160 14965
rect 20200 14995 20240 15000
rect 20200 14965 20205 14995
rect 20235 14965 20240 14995
rect 20200 14960 20240 14965
rect 20280 14995 20320 15000
rect 20280 14965 20285 14995
rect 20315 14965 20320 14995
rect 20280 14960 20320 14965
rect 20360 14995 20400 15000
rect 20360 14965 20365 14995
rect 20395 14965 20400 14995
rect 20360 14960 20400 14965
rect 20440 14995 20480 15000
rect 20440 14965 20445 14995
rect 20475 14965 20480 14995
rect 20440 14960 20480 14965
rect 20520 14995 20560 15000
rect 20520 14965 20525 14995
rect 20555 14965 20560 14995
rect 20520 14960 20560 14965
rect 20600 14995 20640 15000
rect 20600 14965 20605 14995
rect 20635 14965 20640 14995
rect 20600 14960 20640 14965
rect 20680 14995 20720 15000
rect 20680 14965 20685 14995
rect 20715 14965 20720 14995
rect 20680 14960 20720 14965
rect 20760 14995 20800 15000
rect 20760 14965 20765 14995
rect 20795 14965 20800 14995
rect 20760 14960 20800 14965
rect 20840 14995 20880 15000
rect 20840 14965 20845 14995
rect 20875 14965 20880 14995
rect 20840 14960 20880 14965
rect 20920 14995 20960 15000
rect 20920 14965 20925 14995
rect 20955 14965 20960 14995
rect 20920 14960 20960 14965
rect 0 14915 40 14920
rect 0 14885 5 14915
rect 35 14885 40 14915
rect 0 14880 40 14885
rect 80 14915 120 14920
rect 80 14885 85 14915
rect 115 14885 120 14915
rect 80 14880 120 14885
rect 160 14915 200 14920
rect 160 14885 165 14915
rect 195 14885 200 14915
rect 160 14880 200 14885
rect 240 14915 280 14920
rect 240 14885 245 14915
rect 275 14885 280 14915
rect 240 14880 280 14885
rect 320 14915 360 14920
rect 320 14885 325 14915
rect 355 14885 360 14915
rect 320 14880 360 14885
rect 400 14915 440 14920
rect 400 14885 405 14915
rect 435 14885 440 14915
rect 400 14880 440 14885
rect 480 14915 520 14920
rect 480 14885 485 14915
rect 515 14885 520 14915
rect 480 14880 520 14885
rect 560 14915 600 14920
rect 560 14885 565 14915
rect 595 14885 600 14915
rect 560 14880 600 14885
rect 640 14915 680 14920
rect 640 14885 645 14915
rect 675 14885 680 14915
rect 640 14880 680 14885
rect 720 14915 760 14920
rect 720 14885 725 14915
rect 755 14885 760 14915
rect 720 14880 760 14885
rect 800 14915 840 14920
rect 800 14885 805 14915
rect 835 14885 840 14915
rect 800 14880 840 14885
rect 880 14915 920 14920
rect 880 14885 885 14915
rect 915 14885 920 14915
rect 880 14880 920 14885
rect 960 14915 1000 14920
rect 960 14885 965 14915
rect 995 14885 1000 14915
rect 960 14880 1000 14885
rect 1040 14915 1080 14920
rect 1040 14885 1045 14915
rect 1075 14885 1080 14915
rect 1040 14880 1080 14885
rect 1120 14915 1160 14920
rect 1120 14885 1125 14915
rect 1155 14885 1160 14915
rect 1120 14880 1160 14885
rect 1200 14915 1240 14920
rect 1200 14885 1205 14915
rect 1235 14885 1240 14915
rect 1200 14880 1240 14885
rect 1280 14915 1320 14920
rect 1280 14885 1285 14915
rect 1315 14885 1320 14915
rect 1280 14880 1320 14885
rect 1360 14915 1400 14920
rect 1360 14885 1365 14915
rect 1395 14885 1400 14915
rect 1360 14880 1400 14885
rect 1440 14915 1480 14920
rect 1440 14885 1445 14915
rect 1475 14885 1480 14915
rect 1440 14880 1480 14885
rect 1520 14915 1560 14920
rect 1520 14885 1525 14915
rect 1555 14885 1560 14915
rect 1520 14880 1560 14885
rect 1600 14915 1640 14920
rect 1600 14885 1605 14915
rect 1635 14885 1640 14915
rect 1600 14880 1640 14885
rect 1680 14915 1720 14920
rect 1680 14885 1685 14915
rect 1715 14885 1720 14915
rect 1680 14880 1720 14885
rect 1760 14915 1800 14920
rect 1760 14885 1765 14915
rect 1795 14885 1800 14915
rect 1760 14880 1800 14885
rect 1840 14915 1880 14920
rect 1840 14885 1845 14915
rect 1875 14885 1880 14915
rect 1840 14880 1880 14885
rect 1920 14915 1960 14920
rect 1920 14885 1925 14915
rect 1955 14885 1960 14915
rect 1920 14880 1960 14885
rect 2000 14915 2040 14920
rect 2000 14885 2005 14915
rect 2035 14885 2040 14915
rect 2000 14880 2040 14885
rect 2080 14915 2120 14920
rect 2080 14885 2085 14915
rect 2115 14885 2120 14915
rect 2080 14880 2120 14885
rect 2160 14915 2200 14920
rect 2160 14885 2165 14915
rect 2195 14885 2200 14915
rect 2160 14880 2200 14885
rect 2240 14915 2280 14920
rect 2240 14885 2245 14915
rect 2275 14885 2280 14915
rect 2240 14880 2280 14885
rect 2320 14915 2360 14920
rect 2320 14885 2325 14915
rect 2355 14885 2360 14915
rect 2320 14880 2360 14885
rect 2400 14915 2440 14920
rect 2400 14885 2405 14915
rect 2435 14885 2440 14915
rect 2400 14880 2440 14885
rect 2480 14915 2520 14920
rect 2480 14885 2485 14915
rect 2515 14885 2520 14915
rect 2480 14880 2520 14885
rect 2560 14915 2600 14920
rect 2560 14885 2565 14915
rect 2595 14885 2600 14915
rect 2560 14880 2600 14885
rect 2640 14915 2680 14920
rect 2640 14885 2645 14915
rect 2675 14885 2680 14915
rect 2640 14880 2680 14885
rect 2720 14915 2760 14920
rect 2720 14885 2725 14915
rect 2755 14885 2760 14915
rect 2720 14880 2760 14885
rect 2800 14915 2840 14920
rect 2800 14885 2805 14915
rect 2835 14885 2840 14915
rect 2800 14880 2840 14885
rect 2880 14915 2920 14920
rect 2880 14885 2885 14915
rect 2915 14885 2920 14915
rect 2880 14880 2920 14885
rect 2960 14915 3000 14920
rect 2960 14885 2965 14915
rect 2995 14885 3000 14915
rect 2960 14880 3000 14885
rect 3040 14915 3080 14920
rect 3040 14885 3045 14915
rect 3075 14885 3080 14915
rect 3040 14880 3080 14885
rect 3120 14915 3160 14920
rect 3120 14885 3125 14915
rect 3155 14885 3160 14915
rect 3120 14880 3160 14885
rect 3200 14915 3240 14920
rect 3200 14885 3205 14915
rect 3235 14885 3240 14915
rect 3200 14880 3240 14885
rect 3280 14915 3320 14920
rect 3280 14885 3285 14915
rect 3315 14885 3320 14915
rect 3280 14880 3320 14885
rect 3360 14915 3400 14920
rect 3360 14885 3365 14915
rect 3395 14885 3400 14915
rect 3360 14880 3400 14885
rect 3440 14915 3480 14920
rect 3440 14885 3445 14915
rect 3475 14885 3480 14915
rect 3440 14880 3480 14885
rect 3520 14915 3560 14920
rect 3520 14885 3525 14915
rect 3555 14885 3560 14915
rect 3520 14880 3560 14885
rect 3600 14915 3640 14920
rect 3600 14885 3605 14915
rect 3635 14885 3640 14915
rect 3600 14880 3640 14885
rect 3680 14915 3720 14920
rect 3680 14885 3685 14915
rect 3715 14885 3720 14915
rect 3680 14880 3720 14885
rect 3760 14915 3800 14920
rect 3760 14885 3765 14915
rect 3795 14885 3800 14915
rect 3760 14880 3800 14885
rect 3840 14915 3880 14920
rect 3840 14885 3845 14915
rect 3875 14885 3880 14915
rect 3840 14880 3880 14885
rect 3920 14915 3960 14920
rect 3920 14885 3925 14915
rect 3955 14885 3960 14915
rect 3920 14880 3960 14885
rect 4000 14915 4040 14920
rect 4000 14885 4005 14915
rect 4035 14885 4040 14915
rect 4000 14880 4040 14885
rect 4080 14915 4120 14920
rect 4080 14885 4085 14915
rect 4115 14885 4120 14915
rect 4080 14880 4120 14885
rect 4160 14915 4200 14920
rect 4160 14885 4165 14915
rect 4195 14885 4200 14915
rect 4160 14880 4200 14885
rect 6240 14915 6280 14920
rect 6240 14885 6245 14915
rect 6275 14885 6280 14915
rect 6240 14880 6280 14885
rect 6320 14915 6360 14920
rect 6320 14885 6325 14915
rect 6355 14885 6360 14915
rect 6320 14880 6360 14885
rect 6400 14915 6440 14920
rect 6400 14885 6405 14915
rect 6435 14885 6440 14915
rect 6400 14880 6440 14885
rect 6480 14915 6520 14920
rect 6480 14885 6485 14915
rect 6515 14885 6520 14915
rect 6480 14880 6520 14885
rect 6560 14915 6600 14920
rect 6560 14885 6565 14915
rect 6595 14885 6600 14915
rect 6560 14880 6600 14885
rect 6640 14915 6680 14920
rect 6640 14885 6645 14915
rect 6675 14885 6680 14915
rect 6640 14880 6680 14885
rect 6720 14915 6760 14920
rect 6720 14885 6725 14915
rect 6755 14885 6760 14915
rect 6720 14880 6760 14885
rect 6800 14915 6840 14920
rect 6800 14885 6805 14915
rect 6835 14885 6840 14915
rect 6800 14880 6840 14885
rect 6880 14915 6920 14920
rect 6880 14885 6885 14915
rect 6915 14885 6920 14915
rect 6880 14880 6920 14885
rect 6960 14915 7000 14920
rect 6960 14885 6965 14915
rect 6995 14885 7000 14915
rect 6960 14880 7000 14885
rect 7040 14915 7080 14920
rect 7040 14885 7045 14915
rect 7075 14885 7080 14915
rect 7040 14880 7080 14885
rect 7120 14915 7160 14920
rect 7120 14885 7125 14915
rect 7155 14885 7160 14915
rect 7120 14880 7160 14885
rect 7200 14915 7240 14920
rect 7200 14885 7205 14915
rect 7235 14885 7240 14915
rect 7200 14880 7240 14885
rect 7280 14915 7320 14920
rect 7280 14885 7285 14915
rect 7315 14885 7320 14915
rect 7280 14880 7320 14885
rect 7360 14915 7400 14920
rect 7360 14885 7365 14915
rect 7395 14885 7400 14915
rect 7360 14880 7400 14885
rect 7440 14915 7480 14920
rect 7440 14885 7445 14915
rect 7475 14885 7480 14915
rect 7440 14880 7480 14885
rect 7520 14915 7560 14920
rect 7520 14885 7525 14915
rect 7555 14885 7560 14915
rect 7520 14880 7560 14885
rect 7600 14915 7640 14920
rect 7600 14885 7605 14915
rect 7635 14885 7640 14915
rect 7600 14880 7640 14885
rect 7680 14915 7720 14920
rect 7680 14885 7685 14915
rect 7715 14885 7720 14915
rect 7680 14880 7720 14885
rect 7760 14915 7800 14920
rect 7760 14885 7765 14915
rect 7795 14885 7800 14915
rect 7760 14880 7800 14885
rect 7840 14915 7880 14920
rect 7840 14885 7845 14915
rect 7875 14885 7880 14915
rect 7840 14880 7880 14885
rect 7920 14915 7960 14920
rect 7920 14885 7925 14915
rect 7955 14885 7960 14915
rect 7920 14880 7960 14885
rect 8000 14915 8040 14920
rect 8000 14885 8005 14915
rect 8035 14885 8040 14915
rect 8000 14880 8040 14885
rect 8080 14915 8120 14920
rect 8080 14885 8085 14915
rect 8115 14885 8120 14915
rect 8080 14880 8120 14885
rect 8160 14915 8200 14920
rect 8160 14885 8165 14915
rect 8195 14885 8200 14915
rect 8160 14880 8200 14885
rect 8240 14915 8280 14920
rect 8240 14885 8245 14915
rect 8275 14885 8280 14915
rect 8240 14880 8280 14885
rect 8320 14915 8360 14920
rect 8320 14885 8325 14915
rect 8355 14885 8360 14915
rect 8320 14880 8360 14885
rect 8400 14915 8440 14920
rect 8400 14885 8405 14915
rect 8435 14885 8440 14915
rect 8400 14880 8440 14885
rect 8480 14915 8520 14920
rect 8480 14885 8485 14915
rect 8515 14885 8520 14915
rect 8480 14880 8520 14885
rect 8560 14915 8600 14920
rect 8560 14885 8565 14915
rect 8595 14885 8600 14915
rect 8560 14880 8600 14885
rect 8640 14915 8680 14920
rect 8640 14885 8645 14915
rect 8675 14885 8680 14915
rect 8640 14880 8680 14885
rect 8720 14915 8760 14920
rect 8720 14885 8725 14915
rect 8755 14885 8760 14915
rect 8720 14880 8760 14885
rect 8800 14915 8840 14920
rect 8800 14885 8805 14915
rect 8835 14885 8840 14915
rect 8800 14880 8840 14885
rect 8880 14915 8920 14920
rect 8880 14885 8885 14915
rect 8915 14885 8920 14915
rect 8880 14880 8920 14885
rect 8960 14915 9000 14920
rect 8960 14885 8965 14915
rect 8995 14885 9000 14915
rect 8960 14880 9000 14885
rect 9040 14915 9080 14920
rect 9040 14885 9045 14915
rect 9075 14885 9080 14915
rect 9040 14880 9080 14885
rect 9120 14915 9160 14920
rect 9120 14885 9125 14915
rect 9155 14885 9160 14915
rect 9120 14880 9160 14885
rect 9200 14915 9240 14920
rect 9200 14885 9205 14915
rect 9235 14885 9240 14915
rect 9200 14880 9240 14885
rect 9280 14915 9320 14920
rect 9280 14885 9285 14915
rect 9315 14885 9320 14915
rect 9280 14880 9320 14885
rect 9360 14915 9400 14920
rect 9360 14885 9365 14915
rect 9395 14885 9400 14915
rect 9360 14880 9400 14885
rect 9440 14915 9480 14920
rect 9440 14885 9445 14915
rect 9475 14885 9480 14915
rect 9440 14880 9480 14885
rect 11560 14915 11600 14920
rect 11560 14885 11565 14915
rect 11595 14885 11600 14915
rect 11560 14880 11600 14885
rect 11640 14915 11680 14920
rect 11640 14885 11645 14915
rect 11675 14885 11680 14915
rect 11640 14880 11680 14885
rect 11720 14915 11760 14920
rect 11720 14885 11725 14915
rect 11755 14885 11760 14915
rect 11720 14880 11760 14885
rect 11800 14915 11840 14920
rect 11800 14885 11805 14915
rect 11835 14885 11840 14915
rect 11800 14880 11840 14885
rect 11880 14915 11920 14920
rect 11880 14885 11885 14915
rect 11915 14885 11920 14915
rect 11880 14880 11920 14885
rect 11960 14915 12000 14920
rect 11960 14885 11965 14915
rect 11995 14885 12000 14915
rect 11960 14880 12000 14885
rect 12040 14915 12080 14920
rect 12040 14885 12045 14915
rect 12075 14885 12080 14915
rect 12040 14880 12080 14885
rect 12120 14915 12160 14920
rect 12120 14885 12125 14915
rect 12155 14885 12160 14915
rect 12120 14880 12160 14885
rect 12200 14915 12240 14920
rect 12200 14885 12205 14915
rect 12235 14885 12240 14915
rect 12200 14880 12240 14885
rect 12280 14915 12320 14920
rect 12280 14885 12285 14915
rect 12315 14885 12320 14915
rect 12280 14880 12320 14885
rect 12360 14915 12400 14920
rect 12360 14885 12365 14915
rect 12395 14885 12400 14915
rect 12360 14880 12400 14885
rect 12440 14915 12480 14920
rect 12440 14885 12445 14915
rect 12475 14885 12480 14915
rect 12440 14880 12480 14885
rect 12520 14915 12560 14920
rect 12520 14885 12525 14915
rect 12555 14885 12560 14915
rect 12520 14880 12560 14885
rect 12600 14915 12640 14920
rect 12600 14885 12605 14915
rect 12635 14885 12640 14915
rect 12600 14880 12640 14885
rect 12680 14915 12720 14920
rect 12680 14885 12685 14915
rect 12715 14885 12720 14915
rect 12680 14880 12720 14885
rect 12760 14915 12800 14920
rect 12760 14885 12765 14915
rect 12795 14885 12800 14915
rect 12760 14880 12800 14885
rect 12840 14915 12880 14920
rect 12840 14885 12845 14915
rect 12875 14885 12880 14915
rect 12840 14880 12880 14885
rect 12920 14915 12960 14920
rect 12920 14885 12925 14915
rect 12955 14885 12960 14915
rect 12920 14880 12960 14885
rect 13000 14915 13040 14920
rect 13000 14885 13005 14915
rect 13035 14885 13040 14915
rect 13000 14880 13040 14885
rect 13080 14915 13120 14920
rect 13080 14885 13085 14915
rect 13115 14885 13120 14915
rect 13080 14880 13120 14885
rect 13160 14915 13200 14920
rect 13160 14885 13165 14915
rect 13195 14885 13200 14915
rect 13160 14880 13200 14885
rect 13240 14915 13280 14920
rect 13240 14885 13245 14915
rect 13275 14885 13280 14915
rect 13240 14880 13280 14885
rect 13320 14915 13360 14920
rect 13320 14885 13325 14915
rect 13355 14885 13360 14915
rect 13320 14880 13360 14885
rect 13400 14915 13440 14920
rect 13400 14885 13405 14915
rect 13435 14885 13440 14915
rect 13400 14880 13440 14885
rect 13480 14915 13520 14920
rect 13480 14885 13485 14915
rect 13515 14885 13520 14915
rect 13480 14880 13520 14885
rect 13560 14915 13600 14920
rect 13560 14885 13565 14915
rect 13595 14885 13600 14915
rect 13560 14880 13600 14885
rect 13640 14915 13680 14920
rect 13640 14885 13645 14915
rect 13675 14885 13680 14915
rect 13640 14880 13680 14885
rect 13720 14915 13760 14920
rect 13720 14885 13725 14915
rect 13755 14885 13760 14915
rect 13720 14880 13760 14885
rect 13800 14915 13840 14920
rect 13800 14885 13805 14915
rect 13835 14885 13840 14915
rect 13800 14880 13840 14885
rect 13880 14915 13920 14920
rect 13880 14885 13885 14915
rect 13915 14885 13920 14915
rect 13880 14880 13920 14885
rect 13960 14915 14000 14920
rect 13960 14885 13965 14915
rect 13995 14885 14000 14915
rect 13960 14880 14000 14885
rect 14040 14915 14080 14920
rect 14040 14885 14045 14915
rect 14075 14885 14080 14915
rect 14040 14880 14080 14885
rect 14120 14915 14160 14920
rect 14120 14885 14125 14915
rect 14155 14885 14160 14915
rect 14120 14880 14160 14885
rect 14200 14915 14240 14920
rect 14200 14885 14205 14915
rect 14235 14885 14240 14915
rect 14200 14880 14240 14885
rect 14280 14915 14320 14920
rect 14280 14885 14285 14915
rect 14315 14885 14320 14915
rect 14280 14880 14320 14885
rect 14360 14915 14400 14920
rect 14360 14885 14365 14915
rect 14395 14885 14400 14915
rect 14360 14880 14400 14885
rect 14440 14915 14480 14920
rect 14440 14885 14445 14915
rect 14475 14885 14480 14915
rect 14440 14880 14480 14885
rect 14520 14915 14560 14920
rect 14520 14885 14525 14915
rect 14555 14885 14560 14915
rect 14520 14880 14560 14885
rect 14600 14915 14640 14920
rect 14600 14885 14605 14915
rect 14635 14885 14640 14915
rect 14600 14880 14640 14885
rect 14680 14915 14720 14920
rect 14680 14885 14685 14915
rect 14715 14885 14720 14915
rect 14680 14880 14720 14885
rect 16760 14915 16800 14920
rect 16760 14885 16765 14915
rect 16795 14885 16800 14915
rect 16760 14880 16800 14885
rect 16840 14915 16880 14920
rect 16840 14885 16845 14915
rect 16875 14885 16880 14915
rect 16840 14880 16880 14885
rect 16920 14915 16960 14920
rect 16920 14885 16925 14915
rect 16955 14885 16960 14915
rect 16920 14880 16960 14885
rect 17000 14915 17040 14920
rect 17000 14885 17005 14915
rect 17035 14885 17040 14915
rect 17000 14880 17040 14885
rect 17080 14915 17120 14920
rect 17080 14885 17085 14915
rect 17115 14885 17120 14915
rect 17080 14880 17120 14885
rect 17160 14915 17200 14920
rect 17160 14885 17165 14915
rect 17195 14885 17200 14915
rect 17160 14880 17200 14885
rect 17240 14915 17280 14920
rect 17240 14885 17245 14915
rect 17275 14885 17280 14915
rect 17240 14880 17280 14885
rect 17320 14915 17360 14920
rect 17320 14885 17325 14915
rect 17355 14885 17360 14915
rect 17320 14880 17360 14885
rect 17400 14915 17440 14920
rect 17400 14885 17405 14915
rect 17435 14885 17440 14915
rect 17400 14880 17440 14885
rect 17480 14915 17520 14920
rect 17480 14885 17485 14915
rect 17515 14885 17520 14915
rect 17480 14880 17520 14885
rect 17560 14915 17600 14920
rect 17560 14885 17565 14915
rect 17595 14885 17600 14915
rect 17560 14880 17600 14885
rect 17640 14915 17680 14920
rect 17640 14885 17645 14915
rect 17675 14885 17680 14915
rect 17640 14880 17680 14885
rect 17720 14915 17760 14920
rect 17720 14885 17725 14915
rect 17755 14885 17760 14915
rect 17720 14880 17760 14885
rect 17800 14915 17840 14920
rect 17800 14885 17805 14915
rect 17835 14885 17840 14915
rect 17800 14880 17840 14885
rect 17880 14915 17920 14920
rect 17880 14885 17885 14915
rect 17915 14885 17920 14915
rect 17880 14880 17920 14885
rect 17960 14915 18000 14920
rect 17960 14885 17965 14915
rect 17995 14885 18000 14915
rect 17960 14880 18000 14885
rect 18040 14915 18080 14920
rect 18040 14885 18045 14915
rect 18075 14885 18080 14915
rect 18040 14880 18080 14885
rect 18120 14915 18160 14920
rect 18120 14885 18125 14915
rect 18155 14885 18160 14915
rect 18120 14880 18160 14885
rect 18200 14915 18240 14920
rect 18200 14885 18205 14915
rect 18235 14885 18240 14915
rect 18200 14880 18240 14885
rect 18280 14915 18320 14920
rect 18280 14885 18285 14915
rect 18315 14885 18320 14915
rect 18280 14880 18320 14885
rect 18360 14915 18400 14920
rect 18360 14885 18365 14915
rect 18395 14885 18400 14915
rect 18360 14880 18400 14885
rect 18440 14915 18480 14920
rect 18440 14885 18445 14915
rect 18475 14885 18480 14915
rect 18440 14880 18480 14885
rect 18520 14915 18560 14920
rect 18520 14885 18525 14915
rect 18555 14885 18560 14915
rect 18520 14880 18560 14885
rect 18600 14915 18640 14920
rect 18600 14885 18605 14915
rect 18635 14885 18640 14915
rect 18600 14880 18640 14885
rect 18680 14915 18720 14920
rect 18680 14885 18685 14915
rect 18715 14885 18720 14915
rect 18680 14880 18720 14885
rect 18760 14915 18800 14920
rect 18760 14885 18765 14915
rect 18795 14885 18800 14915
rect 18760 14880 18800 14885
rect 18840 14915 18880 14920
rect 18840 14885 18845 14915
rect 18875 14885 18880 14915
rect 18840 14880 18880 14885
rect 18920 14915 18960 14920
rect 18920 14885 18925 14915
rect 18955 14885 18960 14915
rect 18920 14880 18960 14885
rect 19000 14915 19040 14920
rect 19000 14885 19005 14915
rect 19035 14885 19040 14915
rect 19000 14880 19040 14885
rect 19080 14915 19120 14920
rect 19080 14885 19085 14915
rect 19115 14885 19120 14915
rect 19080 14880 19120 14885
rect 19160 14915 19200 14920
rect 19160 14885 19165 14915
rect 19195 14885 19200 14915
rect 19160 14880 19200 14885
rect 19240 14915 19280 14920
rect 19240 14885 19245 14915
rect 19275 14885 19280 14915
rect 19240 14880 19280 14885
rect 19320 14915 19360 14920
rect 19320 14885 19325 14915
rect 19355 14885 19360 14915
rect 19320 14880 19360 14885
rect 19400 14915 19440 14920
rect 19400 14885 19405 14915
rect 19435 14885 19440 14915
rect 19400 14880 19440 14885
rect 19480 14915 19520 14920
rect 19480 14885 19485 14915
rect 19515 14885 19520 14915
rect 19480 14880 19520 14885
rect 19560 14915 19600 14920
rect 19560 14885 19565 14915
rect 19595 14885 19600 14915
rect 19560 14880 19600 14885
rect 19640 14915 19680 14920
rect 19640 14885 19645 14915
rect 19675 14885 19680 14915
rect 19640 14880 19680 14885
rect 19720 14915 19760 14920
rect 19720 14885 19725 14915
rect 19755 14885 19760 14915
rect 19720 14880 19760 14885
rect 19800 14915 19840 14920
rect 19800 14885 19805 14915
rect 19835 14885 19840 14915
rect 19800 14880 19840 14885
rect 19880 14915 19920 14920
rect 19880 14885 19885 14915
rect 19915 14885 19920 14915
rect 19880 14880 19920 14885
rect 19960 14915 20000 14920
rect 19960 14885 19965 14915
rect 19995 14885 20000 14915
rect 19960 14880 20000 14885
rect 20040 14915 20080 14920
rect 20040 14885 20045 14915
rect 20075 14885 20080 14915
rect 20040 14880 20080 14885
rect 20120 14915 20160 14920
rect 20120 14885 20125 14915
rect 20155 14885 20160 14915
rect 20120 14880 20160 14885
rect 20200 14915 20240 14920
rect 20200 14885 20205 14915
rect 20235 14885 20240 14915
rect 20200 14880 20240 14885
rect 20280 14915 20320 14920
rect 20280 14885 20285 14915
rect 20315 14885 20320 14915
rect 20280 14880 20320 14885
rect 20360 14915 20400 14920
rect 20360 14885 20365 14915
rect 20395 14885 20400 14915
rect 20360 14880 20400 14885
rect 20440 14915 20480 14920
rect 20440 14885 20445 14915
rect 20475 14885 20480 14915
rect 20440 14880 20480 14885
rect 20520 14915 20560 14920
rect 20520 14885 20525 14915
rect 20555 14885 20560 14915
rect 20520 14880 20560 14885
rect 20600 14915 20640 14920
rect 20600 14885 20605 14915
rect 20635 14885 20640 14915
rect 20600 14880 20640 14885
rect 20680 14915 20720 14920
rect 20680 14885 20685 14915
rect 20715 14885 20720 14915
rect 20680 14880 20720 14885
rect 20760 14915 20800 14920
rect 20760 14885 20765 14915
rect 20795 14885 20800 14915
rect 20760 14880 20800 14885
rect 20840 14915 20880 14920
rect 20840 14885 20845 14915
rect 20875 14885 20880 14915
rect 20840 14880 20880 14885
rect 20920 14915 20960 14920
rect 20920 14885 20925 14915
rect 20955 14885 20960 14915
rect 20920 14880 20960 14885
rect 0 14755 40 14760
rect 0 14725 5 14755
rect 35 14725 40 14755
rect 0 14720 40 14725
rect 80 14755 120 14760
rect 80 14725 85 14755
rect 115 14725 120 14755
rect 80 14720 120 14725
rect 160 14755 200 14760
rect 160 14725 165 14755
rect 195 14725 200 14755
rect 160 14720 200 14725
rect 240 14755 280 14760
rect 240 14725 245 14755
rect 275 14725 280 14755
rect 240 14720 280 14725
rect 320 14755 360 14760
rect 320 14725 325 14755
rect 355 14725 360 14755
rect 320 14720 360 14725
rect 400 14755 440 14760
rect 400 14725 405 14755
rect 435 14725 440 14755
rect 400 14720 440 14725
rect 480 14755 520 14760
rect 480 14725 485 14755
rect 515 14725 520 14755
rect 480 14720 520 14725
rect 560 14755 600 14760
rect 560 14725 565 14755
rect 595 14725 600 14755
rect 560 14720 600 14725
rect 640 14755 680 14760
rect 640 14725 645 14755
rect 675 14725 680 14755
rect 640 14720 680 14725
rect 720 14755 760 14760
rect 720 14725 725 14755
rect 755 14725 760 14755
rect 720 14720 760 14725
rect 800 14755 840 14760
rect 800 14725 805 14755
rect 835 14725 840 14755
rect 800 14720 840 14725
rect 880 14755 920 14760
rect 880 14725 885 14755
rect 915 14725 920 14755
rect 880 14720 920 14725
rect 960 14755 1000 14760
rect 960 14725 965 14755
rect 995 14725 1000 14755
rect 960 14720 1000 14725
rect 1040 14755 1080 14760
rect 1040 14725 1045 14755
rect 1075 14725 1080 14755
rect 1040 14720 1080 14725
rect 1120 14755 1160 14760
rect 1120 14725 1125 14755
rect 1155 14725 1160 14755
rect 1120 14720 1160 14725
rect 1200 14755 1240 14760
rect 1200 14725 1205 14755
rect 1235 14725 1240 14755
rect 1200 14720 1240 14725
rect 1280 14755 1320 14760
rect 1280 14725 1285 14755
rect 1315 14725 1320 14755
rect 1280 14720 1320 14725
rect 1360 14755 1400 14760
rect 1360 14725 1365 14755
rect 1395 14725 1400 14755
rect 1360 14720 1400 14725
rect 1440 14755 1480 14760
rect 1440 14725 1445 14755
rect 1475 14725 1480 14755
rect 1440 14720 1480 14725
rect 1520 14755 1560 14760
rect 1520 14725 1525 14755
rect 1555 14725 1560 14755
rect 1520 14720 1560 14725
rect 1600 14755 1640 14760
rect 1600 14725 1605 14755
rect 1635 14725 1640 14755
rect 1600 14720 1640 14725
rect 1680 14755 1720 14760
rect 1680 14725 1685 14755
rect 1715 14725 1720 14755
rect 1680 14720 1720 14725
rect 1760 14755 1800 14760
rect 1760 14725 1765 14755
rect 1795 14725 1800 14755
rect 1760 14720 1800 14725
rect 1840 14755 1880 14760
rect 1840 14725 1845 14755
rect 1875 14725 1880 14755
rect 1840 14720 1880 14725
rect 1920 14755 1960 14760
rect 1920 14725 1925 14755
rect 1955 14725 1960 14755
rect 1920 14720 1960 14725
rect 2000 14755 2040 14760
rect 2000 14725 2005 14755
rect 2035 14725 2040 14755
rect 2000 14720 2040 14725
rect 2080 14755 2120 14760
rect 2080 14725 2085 14755
rect 2115 14725 2120 14755
rect 2080 14720 2120 14725
rect 2160 14755 2200 14760
rect 2160 14725 2165 14755
rect 2195 14725 2200 14755
rect 2160 14720 2200 14725
rect 2240 14755 2280 14760
rect 2240 14725 2245 14755
rect 2275 14725 2280 14755
rect 2240 14720 2280 14725
rect 2320 14755 2360 14760
rect 2320 14725 2325 14755
rect 2355 14725 2360 14755
rect 2320 14720 2360 14725
rect 2400 14755 2440 14760
rect 2400 14725 2405 14755
rect 2435 14725 2440 14755
rect 2400 14720 2440 14725
rect 2480 14755 2520 14760
rect 2480 14725 2485 14755
rect 2515 14725 2520 14755
rect 2480 14720 2520 14725
rect 2560 14755 2600 14760
rect 2560 14725 2565 14755
rect 2595 14725 2600 14755
rect 2560 14720 2600 14725
rect 2640 14755 2680 14760
rect 2640 14725 2645 14755
rect 2675 14725 2680 14755
rect 2640 14720 2680 14725
rect 2720 14755 2760 14760
rect 2720 14725 2725 14755
rect 2755 14725 2760 14755
rect 2720 14720 2760 14725
rect 2800 14755 2840 14760
rect 2800 14725 2805 14755
rect 2835 14725 2840 14755
rect 2800 14720 2840 14725
rect 2880 14755 2920 14760
rect 2880 14725 2885 14755
rect 2915 14725 2920 14755
rect 2880 14720 2920 14725
rect 2960 14755 3000 14760
rect 2960 14725 2965 14755
rect 2995 14725 3000 14755
rect 2960 14720 3000 14725
rect 3040 14755 3080 14760
rect 3040 14725 3045 14755
rect 3075 14725 3080 14755
rect 3040 14720 3080 14725
rect 3120 14755 3160 14760
rect 3120 14725 3125 14755
rect 3155 14725 3160 14755
rect 3120 14720 3160 14725
rect 3200 14755 3240 14760
rect 3200 14725 3205 14755
rect 3235 14725 3240 14755
rect 3200 14720 3240 14725
rect 3280 14755 3320 14760
rect 3280 14725 3285 14755
rect 3315 14725 3320 14755
rect 3280 14720 3320 14725
rect 3360 14755 3400 14760
rect 3360 14725 3365 14755
rect 3395 14725 3400 14755
rect 3360 14720 3400 14725
rect 3440 14755 3480 14760
rect 3440 14725 3445 14755
rect 3475 14725 3480 14755
rect 3440 14720 3480 14725
rect 3520 14755 3560 14760
rect 3520 14725 3525 14755
rect 3555 14725 3560 14755
rect 3520 14720 3560 14725
rect 3600 14755 3640 14760
rect 3600 14725 3605 14755
rect 3635 14725 3640 14755
rect 3600 14720 3640 14725
rect 3680 14755 3720 14760
rect 3680 14725 3685 14755
rect 3715 14725 3720 14755
rect 3680 14720 3720 14725
rect 3760 14755 3800 14760
rect 3760 14725 3765 14755
rect 3795 14725 3800 14755
rect 3760 14720 3800 14725
rect 3840 14755 3880 14760
rect 3840 14725 3845 14755
rect 3875 14725 3880 14755
rect 3840 14720 3880 14725
rect 3920 14755 3960 14760
rect 3920 14725 3925 14755
rect 3955 14725 3960 14755
rect 3920 14720 3960 14725
rect 4000 14755 4040 14760
rect 4000 14725 4005 14755
rect 4035 14725 4040 14755
rect 4000 14720 4040 14725
rect 4080 14755 4120 14760
rect 4080 14725 4085 14755
rect 4115 14725 4120 14755
rect 4080 14720 4120 14725
rect 4160 14755 4200 14760
rect 4160 14725 4165 14755
rect 4195 14725 4200 14755
rect 4160 14720 4200 14725
rect 6240 14755 6280 14760
rect 6240 14725 6245 14755
rect 6275 14725 6280 14755
rect 6240 14720 6280 14725
rect 6320 14755 6360 14760
rect 6320 14725 6325 14755
rect 6355 14725 6360 14755
rect 6320 14720 6360 14725
rect 6400 14755 6440 14760
rect 6400 14725 6405 14755
rect 6435 14725 6440 14755
rect 6400 14720 6440 14725
rect 6480 14755 6520 14760
rect 6480 14725 6485 14755
rect 6515 14725 6520 14755
rect 6480 14720 6520 14725
rect 6560 14755 6600 14760
rect 6560 14725 6565 14755
rect 6595 14725 6600 14755
rect 6560 14720 6600 14725
rect 6640 14755 6680 14760
rect 6640 14725 6645 14755
rect 6675 14725 6680 14755
rect 6640 14720 6680 14725
rect 6720 14755 6760 14760
rect 6720 14725 6725 14755
rect 6755 14725 6760 14755
rect 6720 14720 6760 14725
rect 6800 14755 6840 14760
rect 6800 14725 6805 14755
rect 6835 14725 6840 14755
rect 6800 14720 6840 14725
rect 6880 14755 6920 14760
rect 6880 14725 6885 14755
rect 6915 14725 6920 14755
rect 6880 14720 6920 14725
rect 6960 14755 7000 14760
rect 6960 14725 6965 14755
rect 6995 14725 7000 14755
rect 6960 14720 7000 14725
rect 7040 14755 7080 14760
rect 7040 14725 7045 14755
rect 7075 14725 7080 14755
rect 7040 14720 7080 14725
rect 7120 14755 7160 14760
rect 7120 14725 7125 14755
rect 7155 14725 7160 14755
rect 7120 14720 7160 14725
rect 7200 14755 7240 14760
rect 7200 14725 7205 14755
rect 7235 14725 7240 14755
rect 7200 14720 7240 14725
rect 7280 14755 7320 14760
rect 7280 14725 7285 14755
rect 7315 14725 7320 14755
rect 7280 14720 7320 14725
rect 7360 14755 7400 14760
rect 7360 14725 7365 14755
rect 7395 14725 7400 14755
rect 7360 14720 7400 14725
rect 7440 14755 7480 14760
rect 7440 14725 7445 14755
rect 7475 14725 7480 14755
rect 7440 14720 7480 14725
rect 7520 14755 7560 14760
rect 7520 14725 7525 14755
rect 7555 14725 7560 14755
rect 7520 14720 7560 14725
rect 7600 14755 7640 14760
rect 7600 14725 7605 14755
rect 7635 14725 7640 14755
rect 7600 14720 7640 14725
rect 7680 14755 7720 14760
rect 7680 14725 7685 14755
rect 7715 14725 7720 14755
rect 7680 14720 7720 14725
rect 7760 14755 7800 14760
rect 7760 14725 7765 14755
rect 7795 14725 7800 14755
rect 7760 14720 7800 14725
rect 7840 14755 7880 14760
rect 7840 14725 7845 14755
rect 7875 14725 7880 14755
rect 7840 14720 7880 14725
rect 7920 14755 7960 14760
rect 7920 14725 7925 14755
rect 7955 14725 7960 14755
rect 7920 14720 7960 14725
rect 8000 14755 8040 14760
rect 8000 14725 8005 14755
rect 8035 14725 8040 14755
rect 8000 14720 8040 14725
rect 8080 14755 8120 14760
rect 8080 14725 8085 14755
rect 8115 14725 8120 14755
rect 8080 14720 8120 14725
rect 8160 14755 8200 14760
rect 8160 14725 8165 14755
rect 8195 14725 8200 14755
rect 8160 14720 8200 14725
rect 8240 14755 8280 14760
rect 8240 14725 8245 14755
rect 8275 14725 8280 14755
rect 8240 14720 8280 14725
rect 8320 14755 8360 14760
rect 8320 14725 8325 14755
rect 8355 14725 8360 14755
rect 8320 14720 8360 14725
rect 8400 14755 8440 14760
rect 8400 14725 8405 14755
rect 8435 14725 8440 14755
rect 8400 14720 8440 14725
rect 8480 14755 8520 14760
rect 8480 14725 8485 14755
rect 8515 14725 8520 14755
rect 8480 14720 8520 14725
rect 8560 14755 8600 14760
rect 8560 14725 8565 14755
rect 8595 14725 8600 14755
rect 8560 14720 8600 14725
rect 8640 14755 8680 14760
rect 8640 14725 8645 14755
rect 8675 14725 8680 14755
rect 8640 14720 8680 14725
rect 8720 14755 8760 14760
rect 8720 14725 8725 14755
rect 8755 14725 8760 14755
rect 8720 14720 8760 14725
rect 8800 14755 8840 14760
rect 8800 14725 8805 14755
rect 8835 14725 8840 14755
rect 8800 14720 8840 14725
rect 8880 14755 8920 14760
rect 8880 14725 8885 14755
rect 8915 14725 8920 14755
rect 8880 14720 8920 14725
rect 8960 14755 9000 14760
rect 8960 14725 8965 14755
rect 8995 14725 9000 14755
rect 8960 14720 9000 14725
rect 9040 14755 9080 14760
rect 9040 14725 9045 14755
rect 9075 14725 9080 14755
rect 9040 14720 9080 14725
rect 9120 14755 9160 14760
rect 9120 14725 9125 14755
rect 9155 14725 9160 14755
rect 9120 14720 9160 14725
rect 9200 14755 9240 14760
rect 9200 14725 9205 14755
rect 9235 14725 9240 14755
rect 9200 14720 9240 14725
rect 9280 14755 9320 14760
rect 9280 14725 9285 14755
rect 9315 14725 9320 14755
rect 9280 14720 9320 14725
rect 9360 14755 9400 14760
rect 9360 14725 9365 14755
rect 9395 14725 9400 14755
rect 9360 14720 9400 14725
rect 9440 14755 9480 14760
rect 9440 14725 9445 14755
rect 9475 14725 9480 14755
rect 9440 14720 9480 14725
rect 11560 14755 11600 14760
rect 11560 14725 11565 14755
rect 11595 14725 11600 14755
rect 11560 14720 11600 14725
rect 11640 14755 11680 14760
rect 11640 14725 11645 14755
rect 11675 14725 11680 14755
rect 11640 14720 11680 14725
rect 11720 14755 11760 14760
rect 11720 14725 11725 14755
rect 11755 14725 11760 14755
rect 11720 14720 11760 14725
rect 11800 14755 11840 14760
rect 11800 14725 11805 14755
rect 11835 14725 11840 14755
rect 11800 14720 11840 14725
rect 11880 14755 11920 14760
rect 11880 14725 11885 14755
rect 11915 14725 11920 14755
rect 11880 14720 11920 14725
rect 11960 14755 12000 14760
rect 11960 14725 11965 14755
rect 11995 14725 12000 14755
rect 11960 14720 12000 14725
rect 12040 14755 12080 14760
rect 12040 14725 12045 14755
rect 12075 14725 12080 14755
rect 12040 14720 12080 14725
rect 12120 14755 12160 14760
rect 12120 14725 12125 14755
rect 12155 14725 12160 14755
rect 12120 14720 12160 14725
rect 12200 14755 12240 14760
rect 12200 14725 12205 14755
rect 12235 14725 12240 14755
rect 12200 14720 12240 14725
rect 12280 14755 12320 14760
rect 12280 14725 12285 14755
rect 12315 14725 12320 14755
rect 12280 14720 12320 14725
rect 12360 14755 12400 14760
rect 12360 14725 12365 14755
rect 12395 14725 12400 14755
rect 12360 14720 12400 14725
rect 12440 14755 12480 14760
rect 12440 14725 12445 14755
rect 12475 14725 12480 14755
rect 12440 14720 12480 14725
rect 12520 14755 12560 14760
rect 12520 14725 12525 14755
rect 12555 14725 12560 14755
rect 12520 14720 12560 14725
rect 12600 14755 12640 14760
rect 12600 14725 12605 14755
rect 12635 14725 12640 14755
rect 12600 14720 12640 14725
rect 12680 14755 12720 14760
rect 12680 14725 12685 14755
rect 12715 14725 12720 14755
rect 12680 14720 12720 14725
rect 12760 14755 12800 14760
rect 12760 14725 12765 14755
rect 12795 14725 12800 14755
rect 12760 14720 12800 14725
rect 12840 14755 12880 14760
rect 12840 14725 12845 14755
rect 12875 14725 12880 14755
rect 12840 14720 12880 14725
rect 12920 14755 12960 14760
rect 12920 14725 12925 14755
rect 12955 14725 12960 14755
rect 12920 14720 12960 14725
rect 13000 14755 13040 14760
rect 13000 14725 13005 14755
rect 13035 14725 13040 14755
rect 13000 14720 13040 14725
rect 13080 14755 13120 14760
rect 13080 14725 13085 14755
rect 13115 14725 13120 14755
rect 13080 14720 13120 14725
rect 13160 14755 13200 14760
rect 13160 14725 13165 14755
rect 13195 14725 13200 14755
rect 13160 14720 13200 14725
rect 13240 14755 13280 14760
rect 13240 14725 13245 14755
rect 13275 14725 13280 14755
rect 13240 14720 13280 14725
rect 13320 14755 13360 14760
rect 13320 14725 13325 14755
rect 13355 14725 13360 14755
rect 13320 14720 13360 14725
rect 13400 14755 13440 14760
rect 13400 14725 13405 14755
rect 13435 14725 13440 14755
rect 13400 14720 13440 14725
rect 13480 14755 13520 14760
rect 13480 14725 13485 14755
rect 13515 14725 13520 14755
rect 13480 14720 13520 14725
rect 13560 14755 13600 14760
rect 13560 14725 13565 14755
rect 13595 14725 13600 14755
rect 13560 14720 13600 14725
rect 13640 14755 13680 14760
rect 13640 14725 13645 14755
rect 13675 14725 13680 14755
rect 13640 14720 13680 14725
rect 13720 14755 13760 14760
rect 13720 14725 13725 14755
rect 13755 14725 13760 14755
rect 13720 14720 13760 14725
rect 13800 14755 13840 14760
rect 13800 14725 13805 14755
rect 13835 14725 13840 14755
rect 13800 14720 13840 14725
rect 13880 14755 13920 14760
rect 13880 14725 13885 14755
rect 13915 14725 13920 14755
rect 13880 14720 13920 14725
rect 13960 14755 14000 14760
rect 13960 14725 13965 14755
rect 13995 14725 14000 14755
rect 13960 14720 14000 14725
rect 14040 14755 14080 14760
rect 14040 14725 14045 14755
rect 14075 14725 14080 14755
rect 14040 14720 14080 14725
rect 14120 14755 14160 14760
rect 14120 14725 14125 14755
rect 14155 14725 14160 14755
rect 14120 14720 14160 14725
rect 14200 14755 14240 14760
rect 14200 14725 14205 14755
rect 14235 14725 14240 14755
rect 14200 14720 14240 14725
rect 14280 14755 14320 14760
rect 14280 14725 14285 14755
rect 14315 14725 14320 14755
rect 14280 14720 14320 14725
rect 14360 14755 14400 14760
rect 14360 14725 14365 14755
rect 14395 14725 14400 14755
rect 14360 14720 14400 14725
rect 14440 14755 14480 14760
rect 14440 14725 14445 14755
rect 14475 14725 14480 14755
rect 14440 14720 14480 14725
rect 14520 14755 14560 14760
rect 14520 14725 14525 14755
rect 14555 14725 14560 14755
rect 14520 14720 14560 14725
rect 14600 14755 14640 14760
rect 14600 14725 14605 14755
rect 14635 14725 14640 14755
rect 14600 14720 14640 14725
rect 14680 14755 14720 14760
rect 14680 14725 14685 14755
rect 14715 14725 14720 14755
rect 14680 14720 14720 14725
rect 16760 14755 16800 14760
rect 16760 14725 16765 14755
rect 16795 14725 16800 14755
rect 16760 14720 16800 14725
rect 16840 14755 16880 14760
rect 16840 14725 16845 14755
rect 16875 14725 16880 14755
rect 16840 14720 16880 14725
rect 16920 14755 16960 14760
rect 16920 14725 16925 14755
rect 16955 14725 16960 14755
rect 16920 14720 16960 14725
rect 17000 14755 17040 14760
rect 17000 14725 17005 14755
rect 17035 14725 17040 14755
rect 17000 14720 17040 14725
rect 17080 14755 17120 14760
rect 17080 14725 17085 14755
rect 17115 14725 17120 14755
rect 17080 14720 17120 14725
rect 17160 14755 17200 14760
rect 17160 14725 17165 14755
rect 17195 14725 17200 14755
rect 17160 14720 17200 14725
rect 17240 14755 17280 14760
rect 17240 14725 17245 14755
rect 17275 14725 17280 14755
rect 17240 14720 17280 14725
rect 17320 14755 17360 14760
rect 17320 14725 17325 14755
rect 17355 14725 17360 14755
rect 17320 14720 17360 14725
rect 17400 14755 17440 14760
rect 17400 14725 17405 14755
rect 17435 14725 17440 14755
rect 17400 14720 17440 14725
rect 17480 14755 17520 14760
rect 17480 14725 17485 14755
rect 17515 14725 17520 14755
rect 17480 14720 17520 14725
rect 17560 14755 17600 14760
rect 17560 14725 17565 14755
rect 17595 14725 17600 14755
rect 17560 14720 17600 14725
rect 17640 14755 17680 14760
rect 17640 14725 17645 14755
rect 17675 14725 17680 14755
rect 17640 14720 17680 14725
rect 17720 14755 17760 14760
rect 17720 14725 17725 14755
rect 17755 14725 17760 14755
rect 17720 14720 17760 14725
rect 17800 14755 17840 14760
rect 17800 14725 17805 14755
rect 17835 14725 17840 14755
rect 17800 14720 17840 14725
rect 17880 14755 17920 14760
rect 17880 14725 17885 14755
rect 17915 14725 17920 14755
rect 17880 14720 17920 14725
rect 17960 14755 18000 14760
rect 17960 14725 17965 14755
rect 17995 14725 18000 14755
rect 17960 14720 18000 14725
rect 18040 14755 18080 14760
rect 18040 14725 18045 14755
rect 18075 14725 18080 14755
rect 18040 14720 18080 14725
rect 18120 14755 18160 14760
rect 18120 14725 18125 14755
rect 18155 14725 18160 14755
rect 18120 14720 18160 14725
rect 18200 14755 18240 14760
rect 18200 14725 18205 14755
rect 18235 14725 18240 14755
rect 18200 14720 18240 14725
rect 18280 14755 18320 14760
rect 18280 14725 18285 14755
rect 18315 14725 18320 14755
rect 18280 14720 18320 14725
rect 18360 14755 18400 14760
rect 18360 14725 18365 14755
rect 18395 14725 18400 14755
rect 18360 14720 18400 14725
rect 18440 14755 18480 14760
rect 18440 14725 18445 14755
rect 18475 14725 18480 14755
rect 18440 14720 18480 14725
rect 18520 14755 18560 14760
rect 18520 14725 18525 14755
rect 18555 14725 18560 14755
rect 18520 14720 18560 14725
rect 18600 14755 18640 14760
rect 18600 14725 18605 14755
rect 18635 14725 18640 14755
rect 18600 14720 18640 14725
rect 18680 14755 18720 14760
rect 18680 14725 18685 14755
rect 18715 14725 18720 14755
rect 18680 14720 18720 14725
rect 18760 14755 18800 14760
rect 18760 14725 18765 14755
rect 18795 14725 18800 14755
rect 18760 14720 18800 14725
rect 18840 14755 18880 14760
rect 18840 14725 18845 14755
rect 18875 14725 18880 14755
rect 18840 14720 18880 14725
rect 18920 14755 18960 14760
rect 18920 14725 18925 14755
rect 18955 14725 18960 14755
rect 18920 14720 18960 14725
rect 19000 14755 19040 14760
rect 19000 14725 19005 14755
rect 19035 14725 19040 14755
rect 19000 14720 19040 14725
rect 19080 14755 19120 14760
rect 19080 14725 19085 14755
rect 19115 14725 19120 14755
rect 19080 14720 19120 14725
rect 19160 14755 19200 14760
rect 19160 14725 19165 14755
rect 19195 14725 19200 14755
rect 19160 14720 19200 14725
rect 19240 14755 19280 14760
rect 19240 14725 19245 14755
rect 19275 14725 19280 14755
rect 19240 14720 19280 14725
rect 19320 14755 19360 14760
rect 19320 14725 19325 14755
rect 19355 14725 19360 14755
rect 19320 14720 19360 14725
rect 19400 14755 19440 14760
rect 19400 14725 19405 14755
rect 19435 14725 19440 14755
rect 19400 14720 19440 14725
rect 19480 14755 19520 14760
rect 19480 14725 19485 14755
rect 19515 14725 19520 14755
rect 19480 14720 19520 14725
rect 19560 14755 19600 14760
rect 19560 14725 19565 14755
rect 19595 14725 19600 14755
rect 19560 14720 19600 14725
rect 19640 14755 19680 14760
rect 19640 14725 19645 14755
rect 19675 14725 19680 14755
rect 19640 14720 19680 14725
rect 19720 14755 19760 14760
rect 19720 14725 19725 14755
rect 19755 14725 19760 14755
rect 19720 14720 19760 14725
rect 19800 14755 19840 14760
rect 19800 14725 19805 14755
rect 19835 14725 19840 14755
rect 19800 14720 19840 14725
rect 19880 14755 19920 14760
rect 19880 14725 19885 14755
rect 19915 14725 19920 14755
rect 19880 14720 19920 14725
rect 19960 14755 20000 14760
rect 19960 14725 19965 14755
rect 19995 14725 20000 14755
rect 19960 14720 20000 14725
rect 20040 14755 20080 14760
rect 20040 14725 20045 14755
rect 20075 14725 20080 14755
rect 20040 14720 20080 14725
rect 20120 14755 20160 14760
rect 20120 14725 20125 14755
rect 20155 14725 20160 14755
rect 20120 14720 20160 14725
rect 20200 14755 20240 14760
rect 20200 14725 20205 14755
rect 20235 14725 20240 14755
rect 20200 14720 20240 14725
rect 20280 14755 20320 14760
rect 20280 14725 20285 14755
rect 20315 14725 20320 14755
rect 20280 14720 20320 14725
rect 20360 14755 20400 14760
rect 20360 14725 20365 14755
rect 20395 14725 20400 14755
rect 20360 14720 20400 14725
rect 20440 14755 20480 14760
rect 20440 14725 20445 14755
rect 20475 14725 20480 14755
rect 20440 14720 20480 14725
rect 20520 14755 20560 14760
rect 20520 14725 20525 14755
rect 20555 14725 20560 14755
rect 20520 14720 20560 14725
rect 20600 14755 20640 14760
rect 20600 14725 20605 14755
rect 20635 14725 20640 14755
rect 20600 14720 20640 14725
rect 20680 14755 20720 14760
rect 20680 14725 20685 14755
rect 20715 14725 20720 14755
rect 20680 14720 20720 14725
rect 20760 14755 20800 14760
rect 20760 14725 20765 14755
rect 20795 14725 20800 14755
rect 20760 14720 20800 14725
rect 20840 14755 20880 14760
rect 20840 14725 20845 14755
rect 20875 14725 20880 14755
rect 20840 14720 20880 14725
rect 20920 14755 20960 14760
rect 20920 14725 20925 14755
rect 20955 14725 20960 14755
rect 20920 14720 20960 14725
<< via1 >>
rect 5 18670 35 18675
rect 5 18650 10 18670
rect 10 18650 30 18670
rect 30 18650 35 18670
rect 5 18645 35 18650
rect 85 18670 115 18675
rect 85 18650 90 18670
rect 90 18650 110 18670
rect 110 18650 115 18670
rect 85 18645 115 18650
rect 165 18670 195 18675
rect 165 18650 170 18670
rect 170 18650 190 18670
rect 190 18650 195 18670
rect 165 18645 195 18650
rect 245 18670 275 18675
rect 245 18650 250 18670
rect 250 18650 270 18670
rect 270 18650 275 18670
rect 245 18645 275 18650
rect 325 18670 355 18675
rect 325 18650 330 18670
rect 330 18650 350 18670
rect 350 18650 355 18670
rect 325 18645 355 18650
rect 405 18670 435 18675
rect 405 18650 410 18670
rect 410 18650 430 18670
rect 430 18650 435 18670
rect 405 18645 435 18650
rect 485 18670 515 18675
rect 485 18650 490 18670
rect 490 18650 510 18670
rect 510 18650 515 18670
rect 485 18645 515 18650
rect 565 18670 595 18675
rect 565 18650 570 18670
rect 570 18650 590 18670
rect 590 18650 595 18670
rect 565 18645 595 18650
rect 645 18670 675 18675
rect 645 18650 650 18670
rect 650 18650 670 18670
rect 670 18650 675 18670
rect 645 18645 675 18650
rect 725 18670 755 18675
rect 725 18650 730 18670
rect 730 18650 750 18670
rect 750 18650 755 18670
rect 725 18645 755 18650
rect 805 18670 835 18675
rect 805 18650 810 18670
rect 810 18650 830 18670
rect 830 18650 835 18670
rect 805 18645 835 18650
rect 885 18670 915 18675
rect 885 18650 890 18670
rect 890 18650 910 18670
rect 910 18650 915 18670
rect 885 18645 915 18650
rect 965 18670 995 18675
rect 965 18650 970 18670
rect 970 18650 990 18670
rect 990 18650 995 18670
rect 965 18645 995 18650
rect 1045 18670 1075 18675
rect 1045 18650 1050 18670
rect 1050 18650 1070 18670
rect 1070 18650 1075 18670
rect 1045 18645 1075 18650
rect 1125 18670 1155 18675
rect 1125 18650 1130 18670
rect 1130 18650 1150 18670
rect 1150 18650 1155 18670
rect 1125 18645 1155 18650
rect 1205 18670 1235 18675
rect 1205 18650 1210 18670
rect 1210 18650 1230 18670
rect 1230 18650 1235 18670
rect 1205 18645 1235 18650
rect 1285 18670 1315 18675
rect 1285 18650 1290 18670
rect 1290 18650 1310 18670
rect 1310 18650 1315 18670
rect 1285 18645 1315 18650
rect 1365 18670 1395 18675
rect 1365 18650 1370 18670
rect 1370 18650 1390 18670
rect 1390 18650 1395 18670
rect 1365 18645 1395 18650
rect 1445 18670 1475 18675
rect 1445 18650 1450 18670
rect 1450 18650 1470 18670
rect 1470 18650 1475 18670
rect 1445 18645 1475 18650
rect 1525 18670 1555 18675
rect 1525 18650 1530 18670
rect 1530 18650 1550 18670
rect 1550 18650 1555 18670
rect 1525 18645 1555 18650
rect 1605 18670 1635 18675
rect 1605 18650 1610 18670
rect 1610 18650 1630 18670
rect 1630 18650 1635 18670
rect 1605 18645 1635 18650
rect 1685 18670 1715 18675
rect 1685 18650 1690 18670
rect 1690 18650 1710 18670
rect 1710 18650 1715 18670
rect 1685 18645 1715 18650
rect 1765 18670 1795 18675
rect 1765 18650 1770 18670
rect 1770 18650 1790 18670
rect 1790 18650 1795 18670
rect 1765 18645 1795 18650
rect 1845 18670 1875 18675
rect 1845 18650 1850 18670
rect 1850 18650 1870 18670
rect 1870 18650 1875 18670
rect 1845 18645 1875 18650
rect 1925 18670 1955 18675
rect 1925 18650 1930 18670
rect 1930 18650 1950 18670
rect 1950 18650 1955 18670
rect 1925 18645 1955 18650
rect 2005 18670 2035 18675
rect 2005 18650 2010 18670
rect 2010 18650 2030 18670
rect 2030 18650 2035 18670
rect 2005 18645 2035 18650
rect 2085 18670 2115 18675
rect 2085 18650 2090 18670
rect 2090 18650 2110 18670
rect 2110 18650 2115 18670
rect 2085 18645 2115 18650
rect 2165 18670 2195 18675
rect 2165 18650 2170 18670
rect 2170 18650 2190 18670
rect 2190 18650 2195 18670
rect 2165 18645 2195 18650
rect 2245 18670 2275 18675
rect 2245 18650 2250 18670
rect 2250 18650 2270 18670
rect 2270 18650 2275 18670
rect 2245 18645 2275 18650
rect 2325 18670 2355 18675
rect 2325 18650 2330 18670
rect 2330 18650 2350 18670
rect 2350 18650 2355 18670
rect 2325 18645 2355 18650
rect 2405 18670 2435 18675
rect 2405 18650 2410 18670
rect 2410 18650 2430 18670
rect 2430 18650 2435 18670
rect 2405 18645 2435 18650
rect 2485 18670 2515 18675
rect 2485 18650 2490 18670
rect 2490 18650 2510 18670
rect 2510 18650 2515 18670
rect 2485 18645 2515 18650
rect 2565 18670 2595 18675
rect 2565 18650 2570 18670
rect 2570 18650 2590 18670
rect 2590 18650 2595 18670
rect 2565 18645 2595 18650
rect 2645 18670 2675 18675
rect 2645 18650 2650 18670
rect 2650 18650 2670 18670
rect 2670 18650 2675 18670
rect 2645 18645 2675 18650
rect 2725 18670 2755 18675
rect 2725 18650 2730 18670
rect 2730 18650 2750 18670
rect 2750 18650 2755 18670
rect 2725 18645 2755 18650
rect 2805 18670 2835 18675
rect 2805 18650 2810 18670
rect 2810 18650 2830 18670
rect 2830 18650 2835 18670
rect 2805 18645 2835 18650
rect 2885 18670 2915 18675
rect 2885 18650 2890 18670
rect 2890 18650 2910 18670
rect 2910 18650 2915 18670
rect 2885 18645 2915 18650
rect 2965 18670 2995 18675
rect 2965 18650 2970 18670
rect 2970 18650 2990 18670
rect 2990 18650 2995 18670
rect 2965 18645 2995 18650
rect 3045 18670 3075 18675
rect 3045 18650 3050 18670
rect 3050 18650 3070 18670
rect 3070 18650 3075 18670
rect 3045 18645 3075 18650
rect 3125 18670 3155 18675
rect 3125 18650 3130 18670
rect 3130 18650 3150 18670
rect 3150 18650 3155 18670
rect 3125 18645 3155 18650
rect 3205 18670 3235 18675
rect 3205 18650 3210 18670
rect 3210 18650 3230 18670
rect 3230 18650 3235 18670
rect 3205 18645 3235 18650
rect 3285 18670 3315 18675
rect 3285 18650 3290 18670
rect 3290 18650 3310 18670
rect 3310 18650 3315 18670
rect 3285 18645 3315 18650
rect 3365 18670 3395 18675
rect 3365 18650 3370 18670
rect 3370 18650 3390 18670
rect 3390 18650 3395 18670
rect 3365 18645 3395 18650
rect 3445 18670 3475 18675
rect 3445 18650 3450 18670
rect 3450 18650 3470 18670
rect 3470 18650 3475 18670
rect 3445 18645 3475 18650
rect 3525 18670 3555 18675
rect 3525 18650 3530 18670
rect 3530 18650 3550 18670
rect 3550 18650 3555 18670
rect 3525 18645 3555 18650
rect 3605 18670 3635 18675
rect 3605 18650 3610 18670
rect 3610 18650 3630 18670
rect 3630 18650 3635 18670
rect 3605 18645 3635 18650
rect 3685 18670 3715 18675
rect 3685 18650 3690 18670
rect 3690 18650 3710 18670
rect 3710 18650 3715 18670
rect 3685 18645 3715 18650
rect 3765 18670 3795 18675
rect 3765 18650 3770 18670
rect 3770 18650 3790 18670
rect 3790 18650 3795 18670
rect 3765 18645 3795 18650
rect 3845 18670 3875 18675
rect 3845 18650 3850 18670
rect 3850 18650 3870 18670
rect 3870 18650 3875 18670
rect 3845 18645 3875 18650
rect 3925 18670 3955 18675
rect 3925 18650 3930 18670
rect 3930 18650 3950 18670
rect 3950 18650 3955 18670
rect 3925 18645 3955 18650
rect 4005 18670 4035 18675
rect 4005 18650 4010 18670
rect 4010 18650 4030 18670
rect 4030 18650 4035 18670
rect 4005 18645 4035 18650
rect 4085 18670 4115 18675
rect 4085 18650 4090 18670
rect 4090 18650 4110 18670
rect 4110 18650 4115 18670
rect 4085 18645 4115 18650
rect 4165 18670 4195 18675
rect 4165 18650 4170 18670
rect 4170 18650 4190 18670
rect 4190 18650 4195 18670
rect 4165 18645 4195 18650
rect 6245 18670 6275 18675
rect 6245 18650 6250 18670
rect 6250 18650 6270 18670
rect 6270 18650 6275 18670
rect 6245 18645 6275 18650
rect 6325 18670 6355 18675
rect 6325 18650 6330 18670
rect 6330 18650 6350 18670
rect 6350 18650 6355 18670
rect 6325 18645 6355 18650
rect 6405 18670 6435 18675
rect 6405 18650 6410 18670
rect 6410 18650 6430 18670
rect 6430 18650 6435 18670
rect 6405 18645 6435 18650
rect 6485 18670 6515 18675
rect 6485 18650 6490 18670
rect 6490 18650 6510 18670
rect 6510 18650 6515 18670
rect 6485 18645 6515 18650
rect 6565 18670 6595 18675
rect 6565 18650 6570 18670
rect 6570 18650 6590 18670
rect 6590 18650 6595 18670
rect 6565 18645 6595 18650
rect 6645 18670 6675 18675
rect 6645 18650 6650 18670
rect 6650 18650 6670 18670
rect 6670 18650 6675 18670
rect 6645 18645 6675 18650
rect 6725 18670 6755 18675
rect 6725 18650 6730 18670
rect 6730 18650 6750 18670
rect 6750 18650 6755 18670
rect 6725 18645 6755 18650
rect 6805 18670 6835 18675
rect 6805 18650 6810 18670
rect 6810 18650 6830 18670
rect 6830 18650 6835 18670
rect 6805 18645 6835 18650
rect 6885 18670 6915 18675
rect 6885 18650 6890 18670
rect 6890 18650 6910 18670
rect 6910 18650 6915 18670
rect 6885 18645 6915 18650
rect 6965 18670 6995 18675
rect 6965 18650 6970 18670
rect 6970 18650 6990 18670
rect 6990 18650 6995 18670
rect 6965 18645 6995 18650
rect 7045 18670 7075 18675
rect 7045 18650 7050 18670
rect 7050 18650 7070 18670
rect 7070 18650 7075 18670
rect 7045 18645 7075 18650
rect 7125 18670 7155 18675
rect 7125 18650 7130 18670
rect 7130 18650 7150 18670
rect 7150 18650 7155 18670
rect 7125 18645 7155 18650
rect 7205 18670 7235 18675
rect 7205 18650 7210 18670
rect 7210 18650 7230 18670
rect 7230 18650 7235 18670
rect 7205 18645 7235 18650
rect 7285 18670 7315 18675
rect 7285 18650 7290 18670
rect 7290 18650 7310 18670
rect 7310 18650 7315 18670
rect 7285 18645 7315 18650
rect 7365 18670 7395 18675
rect 7365 18650 7370 18670
rect 7370 18650 7390 18670
rect 7390 18650 7395 18670
rect 7365 18645 7395 18650
rect 7445 18670 7475 18675
rect 7445 18650 7450 18670
rect 7450 18650 7470 18670
rect 7470 18650 7475 18670
rect 7445 18645 7475 18650
rect 7525 18670 7555 18675
rect 7525 18650 7530 18670
rect 7530 18650 7550 18670
rect 7550 18650 7555 18670
rect 7525 18645 7555 18650
rect 7605 18670 7635 18675
rect 7605 18650 7610 18670
rect 7610 18650 7630 18670
rect 7630 18650 7635 18670
rect 7605 18645 7635 18650
rect 7685 18670 7715 18675
rect 7685 18650 7690 18670
rect 7690 18650 7710 18670
rect 7710 18650 7715 18670
rect 7685 18645 7715 18650
rect 7765 18670 7795 18675
rect 7765 18650 7770 18670
rect 7770 18650 7790 18670
rect 7790 18650 7795 18670
rect 7765 18645 7795 18650
rect 7845 18670 7875 18675
rect 7845 18650 7850 18670
rect 7850 18650 7870 18670
rect 7870 18650 7875 18670
rect 7845 18645 7875 18650
rect 7925 18670 7955 18675
rect 7925 18650 7930 18670
rect 7930 18650 7950 18670
rect 7950 18650 7955 18670
rect 7925 18645 7955 18650
rect 8005 18670 8035 18675
rect 8005 18650 8010 18670
rect 8010 18650 8030 18670
rect 8030 18650 8035 18670
rect 8005 18645 8035 18650
rect 8085 18670 8115 18675
rect 8085 18650 8090 18670
rect 8090 18650 8110 18670
rect 8110 18650 8115 18670
rect 8085 18645 8115 18650
rect 8165 18670 8195 18675
rect 8165 18650 8170 18670
rect 8170 18650 8190 18670
rect 8190 18650 8195 18670
rect 8165 18645 8195 18650
rect 8245 18670 8275 18675
rect 8245 18650 8250 18670
rect 8250 18650 8270 18670
rect 8270 18650 8275 18670
rect 8245 18645 8275 18650
rect 8325 18670 8355 18675
rect 8325 18650 8330 18670
rect 8330 18650 8350 18670
rect 8350 18650 8355 18670
rect 8325 18645 8355 18650
rect 8405 18670 8435 18675
rect 8405 18650 8410 18670
rect 8410 18650 8430 18670
rect 8430 18650 8435 18670
rect 8405 18645 8435 18650
rect 8485 18670 8515 18675
rect 8485 18650 8490 18670
rect 8490 18650 8510 18670
rect 8510 18650 8515 18670
rect 8485 18645 8515 18650
rect 8565 18670 8595 18675
rect 8565 18650 8570 18670
rect 8570 18650 8590 18670
rect 8590 18650 8595 18670
rect 8565 18645 8595 18650
rect 8645 18670 8675 18675
rect 8645 18650 8650 18670
rect 8650 18650 8670 18670
rect 8670 18650 8675 18670
rect 8645 18645 8675 18650
rect 8725 18670 8755 18675
rect 8725 18650 8730 18670
rect 8730 18650 8750 18670
rect 8750 18650 8755 18670
rect 8725 18645 8755 18650
rect 8805 18670 8835 18675
rect 8805 18650 8810 18670
rect 8810 18650 8830 18670
rect 8830 18650 8835 18670
rect 8805 18645 8835 18650
rect 8885 18670 8915 18675
rect 8885 18650 8890 18670
rect 8890 18650 8910 18670
rect 8910 18650 8915 18670
rect 8885 18645 8915 18650
rect 8965 18670 8995 18675
rect 8965 18650 8970 18670
rect 8970 18650 8990 18670
rect 8990 18650 8995 18670
rect 8965 18645 8995 18650
rect 9045 18670 9075 18675
rect 9045 18650 9050 18670
rect 9050 18650 9070 18670
rect 9070 18650 9075 18670
rect 9045 18645 9075 18650
rect 9125 18670 9155 18675
rect 9125 18650 9130 18670
rect 9130 18650 9150 18670
rect 9150 18650 9155 18670
rect 9125 18645 9155 18650
rect 9205 18670 9235 18675
rect 9205 18650 9210 18670
rect 9210 18650 9230 18670
rect 9230 18650 9235 18670
rect 9205 18645 9235 18650
rect 9285 18670 9315 18675
rect 9285 18650 9290 18670
rect 9290 18650 9310 18670
rect 9310 18650 9315 18670
rect 9285 18645 9315 18650
rect 9365 18670 9395 18675
rect 9365 18650 9370 18670
rect 9370 18650 9390 18670
rect 9390 18650 9395 18670
rect 9365 18645 9395 18650
rect 9445 18670 9475 18675
rect 9445 18650 9450 18670
rect 9450 18650 9470 18670
rect 9470 18650 9475 18670
rect 9445 18645 9475 18650
rect 11565 18670 11595 18675
rect 11565 18650 11570 18670
rect 11570 18650 11590 18670
rect 11590 18650 11595 18670
rect 11565 18645 11595 18650
rect 11645 18670 11675 18675
rect 11645 18650 11650 18670
rect 11650 18650 11670 18670
rect 11670 18650 11675 18670
rect 11645 18645 11675 18650
rect 11725 18670 11755 18675
rect 11725 18650 11730 18670
rect 11730 18650 11750 18670
rect 11750 18650 11755 18670
rect 11725 18645 11755 18650
rect 11805 18670 11835 18675
rect 11805 18650 11810 18670
rect 11810 18650 11830 18670
rect 11830 18650 11835 18670
rect 11805 18645 11835 18650
rect 11885 18670 11915 18675
rect 11885 18650 11890 18670
rect 11890 18650 11910 18670
rect 11910 18650 11915 18670
rect 11885 18645 11915 18650
rect 11965 18670 11995 18675
rect 11965 18650 11970 18670
rect 11970 18650 11990 18670
rect 11990 18650 11995 18670
rect 11965 18645 11995 18650
rect 12045 18670 12075 18675
rect 12045 18650 12050 18670
rect 12050 18650 12070 18670
rect 12070 18650 12075 18670
rect 12045 18645 12075 18650
rect 12125 18670 12155 18675
rect 12125 18650 12130 18670
rect 12130 18650 12150 18670
rect 12150 18650 12155 18670
rect 12125 18645 12155 18650
rect 12205 18670 12235 18675
rect 12205 18650 12210 18670
rect 12210 18650 12230 18670
rect 12230 18650 12235 18670
rect 12205 18645 12235 18650
rect 12285 18670 12315 18675
rect 12285 18650 12290 18670
rect 12290 18650 12310 18670
rect 12310 18650 12315 18670
rect 12285 18645 12315 18650
rect 12365 18670 12395 18675
rect 12365 18650 12370 18670
rect 12370 18650 12390 18670
rect 12390 18650 12395 18670
rect 12365 18645 12395 18650
rect 12445 18670 12475 18675
rect 12445 18650 12450 18670
rect 12450 18650 12470 18670
rect 12470 18650 12475 18670
rect 12445 18645 12475 18650
rect 12525 18670 12555 18675
rect 12525 18650 12530 18670
rect 12530 18650 12550 18670
rect 12550 18650 12555 18670
rect 12525 18645 12555 18650
rect 12605 18670 12635 18675
rect 12605 18650 12610 18670
rect 12610 18650 12630 18670
rect 12630 18650 12635 18670
rect 12605 18645 12635 18650
rect 12685 18670 12715 18675
rect 12685 18650 12690 18670
rect 12690 18650 12710 18670
rect 12710 18650 12715 18670
rect 12685 18645 12715 18650
rect 12765 18670 12795 18675
rect 12765 18650 12770 18670
rect 12770 18650 12790 18670
rect 12790 18650 12795 18670
rect 12765 18645 12795 18650
rect 12845 18670 12875 18675
rect 12845 18650 12850 18670
rect 12850 18650 12870 18670
rect 12870 18650 12875 18670
rect 12845 18645 12875 18650
rect 12925 18670 12955 18675
rect 12925 18650 12930 18670
rect 12930 18650 12950 18670
rect 12950 18650 12955 18670
rect 12925 18645 12955 18650
rect 13005 18670 13035 18675
rect 13005 18650 13010 18670
rect 13010 18650 13030 18670
rect 13030 18650 13035 18670
rect 13005 18645 13035 18650
rect 13085 18670 13115 18675
rect 13085 18650 13090 18670
rect 13090 18650 13110 18670
rect 13110 18650 13115 18670
rect 13085 18645 13115 18650
rect 13165 18670 13195 18675
rect 13165 18650 13170 18670
rect 13170 18650 13190 18670
rect 13190 18650 13195 18670
rect 13165 18645 13195 18650
rect 13245 18670 13275 18675
rect 13245 18650 13250 18670
rect 13250 18650 13270 18670
rect 13270 18650 13275 18670
rect 13245 18645 13275 18650
rect 13325 18670 13355 18675
rect 13325 18650 13330 18670
rect 13330 18650 13350 18670
rect 13350 18650 13355 18670
rect 13325 18645 13355 18650
rect 13405 18670 13435 18675
rect 13405 18650 13410 18670
rect 13410 18650 13430 18670
rect 13430 18650 13435 18670
rect 13405 18645 13435 18650
rect 13485 18670 13515 18675
rect 13485 18650 13490 18670
rect 13490 18650 13510 18670
rect 13510 18650 13515 18670
rect 13485 18645 13515 18650
rect 13565 18670 13595 18675
rect 13565 18650 13570 18670
rect 13570 18650 13590 18670
rect 13590 18650 13595 18670
rect 13565 18645 13595 18650
rect 13645 18670 13675 18675
rect 13645 18650 13650 18670
rect 13650 18650 13670 18670
rect 13670 18650 13675 18670
rect 13645 18645 13675 18650
rect 13725 18670 13755 18675
rect 13725 18650 13730 18670
rect 13730 18650 13750 18670
rect 13750 18650 13755 18670
rect 13725 18645 13755 18650
rect 13805 18670 13835 18675
rect 13805 18650 13810 18670
rect 13810 18650 13830 18670
rect 13830 18650 13835 18670
rect 13805 18645 13835 18650
rect 13885 18670 13915 18675
rect 13885 18650 13890 18670
rect 13890 18650 13910 18670
rect 13910 18650 13915 18670
rect 13885 18645 13915 18650
rect 13965 18670 13995 18675
rect 13965 18650 13970 18670
rect 13970 18650 13990 18670
rect 13990 18650 13995 18670
rect 13965 18645 13995 18650
rect 14045 18670 14075 18675
rect 14045 18650 14050 18670
rect 14050 18650 14070 18670
rect 14070 18650 14075 18670
rect 14045 18645 14075 18650
rect 14125 18670 14155 18675
rect 14125 18650 14130 18670
rect 14130 18650 14150 18670
rect 14150 18650 14155 18670
rect 14125 18645 14155 18650
rect 14205 18670 14235 18675
rect 14205 18650 14210 18670
rect 14210 18650 14230 18670
rect 14230 18650 14235 18670
rect 14205 18645 14235 18650
rect 14285 18670 14315 18675
rect 14285 18650 14290 18670
rect 14290 18650 14310 18670
rect 14310 18650 14315 18670
rect 14285 18645 14315 18650
rect 14365 18670 14395 18675
rect 14365 18650 14370 18670
rect 14370 18650 14390 18670
rect 14390 18650 14395 18670
rect 14365 18645 14395 18650
rect 14445 18670 14475 18675
rect 14445 18650 14450 18670
rect 14450 18650 14470 18670
rect 14470 18650 14475 18670
rect 14445 18645 14475 18650
rect 14525 18670 14555 18675
rect 14525 18650 14530 18670
rect 14530 18650 14550 18670
rect 14550 18650 14555 18670
rect 14525 18645 14555 18650
rect 14605 18670 14635 18675
rect 14605 18650 14610 18670
rect 14610 18650 14630 18670
rect 14630 18650 14635 18670
rect 14605 18645 14635 18650
rect 14685 18670 14715 18675
rect 14685 18650 14690 18670
rect 14690 18650 14710 18670
rect 14710 18650 14715 18670
rect 14685 18645 14715 18650
rect 16765 18670 16795 18675
rect 16765 18650 16770 18670
rect 16770 18650 16790 18670
rect 16790 18650 16795 18670
rect 16765 18645 16795 18650
rect 16845 18670 16875 18675
rect 16845 18650 16850 18670
rect 16850 18650 16870 18670
rect 16870 18650 16875 18670
rect 16845 18645 16875 18650
rect 16925 18670 16955 18675
rect 16925 18650 16930 18670
rect 16930 18650 16950 18670
rect 16950 18650 16955 18670
rect 16925 18645 16955 18650
rect 17005 18670 17035 18675
rect 17005 18650 17010 18670
rect 17010 18650 17030 18670
rect 17030 18650 17035 18670
rect 17005 18645 17035 18650
rect 17085 18670 17115 18675
rect 17085 18650 17090 18670
rect 17090 18650 17110 18670
rect 17110 18650 17115 18670
rect 17085 18645 17115 18650
rect 17165 18670 17195 18675
rect 17165 18650 17170 18670
rect 17170 18650 17190 18670
rect 17190 18650 17195 18670
rect 17165 18645 17195 18650
rect 17245 18670 17275 18675
rect 17245 18650 17250 18670
rect 17250 18650 17270 18670
rect 17270 18650 17275 18670
rect 17245 18645 17275 18650
rect 17325 18670 17355 18675
rect 17325 18650 17330 18670
rect 17330 18650 17350 18670
rect 17350 18650 17355 18670
rect 17325 18645 17355 18650
rect 17405 18670 17435 18675
rect 17405 18650 17410 18670
rect 17410 18650 17430 18670
rect 17430 18650 17435 18670
rect 17405 18645 17435 18650
rect 17485 18670 17515 18675
rect 17485 18650 17490 18670
rect 17490 18650 17510 18670
rect 17510 18650 17515 18670
rect 17485 18645 17515 18650
rect 17565 18670 17595 18675
rect 17565 18650 17570 18670
rect 17570 18650 17590 18670
rect 17590 18650 17595 18670
rect 17565 18645 17595 18650
rect 17645 18670 17675 18675
rect 17645 18650 17650 18670
rect 17650 18650 17670 18670
rect 17670 18650 17675 18670
rect 17645 18645 17675 18650
rect 17725 18670 17755 18675
rect 17725 18650 17730 18670
rect 17730 18650 17750 18670
rect 17750 18650 17755 18670
rect 17725 18645 17755 18650
rect 17805 18670 17835 18675
rect 17805 18650 17810 18670
rect 17810 18650 17830 18670
rect 17830 18650 17835 18670
rect 17805 18645 17835 18650
rect 17885 18670 17915 18675
rect 17885 18650 17890 18670
rect 17890 18650 17910 18670
rect 17910 18650 17915 18670
rect 17885 18645 17915 18650
rect 17965 18670 17995 18675
rect 17965 18650 17970 18670
rect 17970 18650 17990 18670
rect 17990 18650 17995 18670
rect 17965 18645 17995 18650
rect 18045 18670 18075 18675
rect 18045 18650 18050 18670
rect 18050 18650 18070 18670
rect 18070 18650 18075 18670
rect 18045 18645 18075 18650
rect 18125 18670 18155 18675
rect 18125 18650 18130 18670
rect 18130 18650 18150 18670
rect 18150 18650 18155 18670
rect 18125 18645 18155 18650
rect 18205 18670 18235 18675
rect 18205 18650 18210 18670
rect 18210 18650 18230 18670
rect 18230 18650 18235 18670
rect 18205 18645 18235 18650
rect 18285 18670 18315 18675
rect 18285 18650 18290 18670
rect 18290 18650 18310 18670
rect 18310 18650 18315 18670
rect 18285 18645 18315 18650
rect 18365 18670 18395 18675
rect 18365 18650 18370 18670
rect 18370 18650 18390 18670
rect 18390 18650 18395 18670
rect 18365 18645 18395 18650
rect 18445 18670 18475 18675
rect 18445 18650 18450 18670
rect 18450 18650 18470 18670
rect 18470 18650 18475 18670
rect 18445 18645 18475 18650
rect 18525 18670 18555 18675
rect 18525 18650 18530 18670
rect 18530 18650 18550 18670
rect 18550 18650 18555 18670
rect 18525 18645 18555 18650
rect 18605 18670 18635 18675
rect 18605 18650 18610 18670
rect 18610 18650 18630 18670
rect 18630 18650 18635 18670
rect 18605 18645 18635 18650
rect 18685 18670 18715 18675
rect 18685 18650 18690 18670
rect 18690 18650 18710 18670
rect 18710 18650 18715 18670
rect 18685 18645 18715 18650
rect 18765 18670 18795 18675
rect 18765 18650 18770 18670
rect 18770 18650 18790 18670
rect 18790 18650 18795 18670
rect 18765 18645 18795 18650
rect 18845 18670 18875 18675
rect 18845 18650 18850 18670
rect 18850 18650 18870 18670
rect 18870 18650 18875 18670
rect 18845 18645 18875 18650
rect 18925 18670 18955 18675
rect 18925 18650 18930 18670
rect 18930 18650 18950 18670
rect 18950 18650 18955 18670
rect 18925 18645 18955 18650
rect 19005 18670 19035 18675
rect 19005 18650 19010 18670
rect 19010 18650 19030 18670
rect 19030 18650 19035 18670
rect 19005 18645 19035 18650
rect 19085 18670 19115 18675
rect 19085 18650 19090 18670
rect 19090 18650 19110 18670
rect 19110 18650 19115 18670
rect 19085 18645 19115 18650
rect 19165 18670 19195 18675
rect 19165 18650 19170 18670
rect 19170 18650 19190 18670
rect 19190 18650 19195 18670
rect 19165 18645 19195 18650
rect 19245 18670 19275 18675
rect 19245 18650 19250 18670
rect 19250 18650 19270 18670
rect 19270 18650 19275 18670
rect 19245 18645 19275 18650
rect 19325 18670 19355 18675
rect 19325 18650 19330 18670
rect 19330 18650 19350 18670
rect 19350 18650 19355 18670
rect 19325 18645 19355 18650
rect 19405 18670 19435 18675
rect 19405 18650 19410 18670
rect 19410 18650 19430 18670
rect 19430 18650 19435 18670
rect 19405 18645 19435 18650
rect 19485 18670 19515 18675
rect 19485 18650 19490 18670
rect 19490 18650 19510 18670
rect 19510 18650 19515 18670
rect 19485 18645 19515 18650
rect 19565 18670 19595 18675
rect 19565 18650 19570 18670
rect 19570 18650 19590 18670
rect 19590 18650 19595 18670
rect 19565 18645 19595 18650
rect 19645 18670 19675 18675
rect 19645 18650 19650 18670
rect 19650 18650 19670 18670
rect 19670 18650 19675 18670
rect 19645 18645 19675 18650
rect 19725 18670 19755 18675
rect 19725 18650 19730 18670
rect 19730 18650 19750 18670
rect 19750 18650 19755 18670
rect 19725 18645 19755 18650
rect 19805 18670 19835 18675
rect 19805 18650 19810 18670
rect 19810 18650 19830 18670
rect 19830 18650 19835 18670
rect 19805 18645 19835 18650
rect 19885 18670 19915 18675
rect 19885 18650 19890 18670
rect 19890 18650 19910 18670
rect 19910 18650 19915 18670
rect 19885 18645 19915 18650
rect 19965 18670 19995 18675
rect 19965 18650 19970 18670
rect 19970 18650 19990 18670
rect 19990 18650 19995 18670
rect 19965 18645 19995 18650
rect 20045 18670 20075 18675
rect 20045 18650 20050 18670
rect 20050 18650 20070 18670
rect 20070 18650 20075 18670
rect 20045 18645 20075 18650
rect 20125 18670 20155 18675
rect 20125 18650 20130 18670
rect 20130 18650 20150 18670
rect 20150 18650 20155 18670
rect 20125 18645 20155 18650
rect 20205 18670 20235 18675
rect 20205 18650 20210 18670
rect 20210 18650 20230 18670
rect 20230 18650 20235 18670
rect 20205 18645 20235 18650
rect 20285 18670 20315 18675
rect 20285 18650 20290 18670
rect 20290 18650 20310 18670
rect 20310 18650 20315 18670
rect 20285 18645 20315 18650
rect 20365 18670 20395 18675
rect 20365 18650 20370 18670
rect 20370 18650 20390 18670
rect 20390 18650 20395 18670
rect 20365 18645 20395 18650
rect 20445 18670 20475 18675
rect 20445 18650 20450 18670
rect 20450 18650 20470 18670
rect 20470 18650 20475 18670
rect 20445 18645 20475 18650
rect 20525 18670 20555 18675
rect 20525 18650 20530 18670
rect 20530 18650 20550 18670
rect 20550 18650 20555 18670
rect 20525 18645 20555 18650
rect 20605 18670 20635 18675
rect 20605 18650 20610 18670
rect 20610 18650 20630 18670
rect 20630 18650 20635 18670
rect 20605 18645 20635 18650
rect 20685 18670 20715 18675
rect 20685 18650 20690 18670
rect 20690 18650 20710 18670
rect 20710 18650 20715 18670
rect 20685 18645 20715 18650
rect 20765 18670 20795 18675
rect 20765 18650 20770 18670
rect 20770 18650 20790 18670
rect 20790 18650 20795 18670
rect 20765 18645 20795 18650
rect 20845 18670 20875 18675
rect 20845 18650 20850 18670
rect 20850 18650 20870 18670
rect 20870 18650 20875 18670
rect 20845 18645 20875 18650
rect 20925 18670 20955 18675
rect 20925 18650 20930 18670
rect 20930 18650 20950 18670
rect 20950 18650 20955 18670
rect 20925 18645 20955 18650
rect 5 18510 35 18515
rect 5 18490 10 18510
rect 10 18490 30 18510
rect 30 18490 35 18510
rect 5 18485 35 18490
rect 85 18510 115 18515
rect 85 18490 90 18510
rect 90 18490 110 18510
rect 110 18490 115 18510
rect 85 18485 115 18490
rect 165 18510 195 18515
rect 165 18490 170 18510
rect 170 18490 190 18510
rect 190 18490 195 18510
rect 165 18485 195 18490
rect 245 18510 275 18515
rect 245 18490 250 18510
rect 250 18490 270 18510
rect 270 18490 275 18510
rect 245 18485 275 18490
rect 325 18510 355 18515
rect 325 18490 330 18510
rect 330 18490 350 18510
rect 350 18490 355 18510
rect 325 18485 355 18490
rect 405 18510 435 18515
rect 405 18490 410 18510
rect 410 18490 430 18510
rect 430 18490 435 18510
rect 405 18485 435 18490
rect 485 18510 515 18515
rect 485 18490 490 18510
rect 490 18490 510 18510
rect 510 18490 515 18510
rect 485 18485 515 18490
rect 565 18510 595 18515
rect 565 18490 570 18510
rect 570 18490 590 18510
rect 590 18490 595 18510
rect 565 18485 595 18490
rect 645 18510 675 18515
rect 645 18490 650 18510
rect 650 18490 670 18510
rect 670 18490 675 18510
rect 645 18485 675 18490
rect 725 18510 755 18515
rect 725 18490 730 18510
rect 730 18490 750 18510
rect 750 18490 755 18510
rect 725 18485 755 18490
rect 805 18510 835 18515
rect 805 18490 810 18510
rect 810 18490 830 18510
rect 830 18490 835 18510
rect 805 18485 835 18490
rect 885 18510 915 18515
rect 885 18490 890 18510
rect 890 18490 910 18510
rect 910 18490 915 18510
rect 885 18485 915 18490
rect 965 18510 995 18515
rect 965 18490 970 18510
rect 970 18490 990 18510
rect 990 18490 995 18510
rect 965 18485 995 18490
rect 1045 18510 1075 18515
rect 1045 18490 1050 18510
rect 1050 18490 1070 18510
rect 1070 18490 1075 18510
rect 1045 18485 1075 18490
rect 1125 18510 1155 18515
rect 1125 18490 1130 18510
rect 1130 18490 1150 18510
rect 1150 18490 1155 18510
rect 1125 18485 1155 18490
rect 1205 18510 1235 18515
rect 1205 18490 1210 18510
rect 1210 18490 1230 18510
rect 1230 18490 1235 18510
rect 1205 18485 1235 18490
rect 1285 18510 1315 18515
rect 1285 18490 1290 18510
rect 1290 18490 1310 18510
rect 1310 18490 1315 18510
rect 1285 18485 1315 18490
rect 1365 18510 1395 18515
rect 1365 18490 1370 18510
rect 1370 18490 1390 18510
rect 1390 18490 1395 18510
rect 1365 18485 1395 18490
rect 1445 18510 1475 18515
rect 1445 18490 1450 18510
rect 1450 18490 1470 18510
rect 1470 18490 1475 18510
rect 1445 18485 1475 18490
rect 1525 18510 1555 18515
rect 1525 18490 1530 18510
rect 1530 18490 1550 18510
rect 1550 18490 1555 18510
rect 1525 18485 1555 18490
rect 1605 18510 1635 18515
rect 1605 18490 1610 18510
rect 1610 18490 1630 18510
rect 1630 18490 1635 18510
rect 1605 18485 1635 18490
rect 1685 18510 1715 18515
rect 1685 18490 1690 18510
rect 1690 18490 1710 18510
rect 1710 18490 1715 18510
rect 1685 18485 1715 18490
rect 1765 18510 1795 18515
rect 1765 18490 1770 18510
rect 1770 18490 1790 18510
rect 1790 18490 1795 18510
rect 1765 18485 1795 18490
rect 1845 18510 1875 18515
rect 1845 18490 1850 18510
rect 1850 18490 1870 18510
rect 1870 18490 1875 18510
rect 1845 18485 1875 18490
rect 1925 18510 1955 18515
rect 1925 18490 1930 18510
rect 1930 18490 1950 18510
rect 1950 18490 1955 18510
rect 1925 18485 1955 18490
rect 2005 18510 2035 18515
rect 2005 18490 2010 18510
rect 2010 18490 2030 18510
rect 2030 18490 2035 18510
rect 2005 18485 2035 18490
rect 2085 18510 2115 18515
rect 2085 18490 2090 18510
rect 2090 18490 2110 18510
rect 2110 18490 2115 18510
rect 2085 18485 2115 18490
rect 2165 18510 2195 18515
rect 2165 18490 2170 18510
rect 2170 18490 2190 18510
rect 2190 18490 2195 18510
rect 2165 18485 2195 18490
rect 2245 18510 2275 18515
rect 2245 18490 2250 18510
rect 2250 18490 2270 18510
rect 2270 18490 2275 18510
rect 2245 18485 2275 18490
rect 2325 18510 2355 18515
rect 2325 18490 2330 18510
rect 2330 18490 2350 18510
rect 2350 18490 2355 18510
rect 2325 18485 2355 18490
rect 2405 18510 2435 18515
rect 2405 18490 2410 18510
rect 2410 18490 2430 18510
rect 2430 18490 2435 18510
rect 2405 18485 2435 18490
rect 2485 18510 2515 18515
rect 2485 18490 2490 18510
rect 2490 18490 2510 18510
rect 2510 18490 2515 18510
rect 2485 18485 2515 18490
rect 2565 18510 2595 18515
rect 2565 18490 2570 18510
rect 2570 18490 2590 18510
rect 2590 18490 2595 18510
rect 2565 18485 2595 18490
rect 2645 18510 2675 18515
rect 2645 18490 2650 18510
rect 2650 18490 2670 18510
rect 2670 18490 2675 18510
rect 2645 18485 2675 18490
rect 2725 18510 2755 18515
rect 2725 18490 2730 18510
rect 2730 18490 2750 18510
rect 2750 18490 2755 18510
rect 2725 18485 2755 18490
rect 2805 18510 2835 18515
rect 2805 18490 2810 18510
rect 2810 18490 2830 18510
rect 2830 18490 2835 18510
rect 2805 18485 2835 18490
rect 2885 18510 2915 18515
rect 2885 18490 2890 18510
rect 2890 18490 2910 18510
rect 2910 18490 2915 18510
rect 2885 18485 2915 18490
rect 2965 18510 2995 18515
rect 2965 18490 2970 18510
rect 2970 18490 2990 18510
rect 2990 18490 2995 18510
rect 2965 18485 2995 18490
rect 3045 18510 3075 18515
rect 3045 18490 3050 18510
rect 3050 18490 3070 18510
rect 3070 18490 3075 18510
rect 3045 18485 3075 18490
rect 3125 18510 3155 18515
rect 3125 18490 3130 18510
rect 3130 18490 3150 18510
rect 3150 18490 3155 18510
rect 3125 18485 3155 18490
rect 3205 18510 3235 18515
rect 3205 18490 3210 18510
rect 3210 18490 3230 18510
rect 3230 18490 3235 18510
rect 3205 18485 3235 18490
rect 3285 18510 3315 18515
rect 3285 18490 3290 18510
rect 3290 18490 3310 18510
rect 3310 18490 3315 18510
rect 3285 18485 3315 18490
rect 3365 18510 3395 18515
rect 3365 18490 3370 18510
rect 3370 18490 3390 18510
rect 3390 18490 3395 18510
rect 3365 18485 3395 18490
rect 3445 18510 3475 18515
rect 3445 18490 3450 18510
rect 3450 18490 3470 18510
rect 3470 18490 3475 18510
rect 3445 18485 3475 18490
rect 3525 18510 3555 18515
rect 3525 18490 3530 18510
rect 3530 18490 3550 18510
rect 3550 18490 3555 18510
rect 3525 18485 3555 18490
rect 3605 18510 3635 18515
rect 3605 18490 3610 18510
rect 3610 18490 3630 18510
rect 3630 18490 3635 18510
rect 3605 18485 3635 18490
rect 3685 18510 3715 18515
rect 3685 18490 3690 18510
rect 3690 18490 3710 18510
rect 3710 18490 3715 18510
rect 3685 18485 3715 18490
rect 3765 18510 3795 18515
rect 3765 18490 3770 18510
rect 3770 18490 3790 18510
rect 3790 18490 3795 18510
rect 3765 18485 3795 18490
rect 3845 18510 3875 18515
rect 3845 18490 3850 18510
rect 3850 18490 3870 18510
rect 3870 18490 3875 18510
rect 3845 18485 3875 18490
rect 3925 18510 3955 18515
rect 3925 18490 3930 18510
rect 3930 18490 3950 18510
rect 3950 18490 3955 18510
rect 3925 18485 3955 18490
rect 4005 18510 4035 18515
rect 4005 18490 4010 18510
rect 4010 18490 4030 18510
rect 4030 18490 4035 18510
rect 4005 18485 4035 18490
rect 4085 18510 4115 18515
rect 4085 18490 4090 18510
rect 4090 18490 4110 18510
rect 4110 18490 4115 18510
rect 4085 18485 4115 18490
rect 4165 18510 4195 18515
rect 4165 18490 4170 18510
rect 4170 18490 4190 18510
rect 4190 18490 4195 18510
rect 4165 18485 4195 18490
rect 6245 18510 6275 18515
rect 6245 18490 6250 18510
rect 6250 18490 6270 18510
rect 6270 18490 6275 18510
rect 6245 18485 6275 18490
rect 6325 18510 6355 18515
rect 6325 18490 6330 18510
rect 6330 18490 6350 18510
rect 6350 18490 6355 18510
rect 6325 18485 6355 18490
rect 6405 18510 6435 18515
rect 6405 18490 6410 18510
rect 6410 18490 6430 18510
rect 6430 18490 6435 18510
rect 6405 18485 6435 18490
rect 6485 18510 6515 18515
rect 6485 18490 6490 18510
rect 6490 18490 6510 18510
rect 6510 18490 6515 18510
rect 6485 18485 6515 18490
rect 6565 18510 6595 18515
rect 6565 18490 6570 18510
rect 6570 18490 6590 18510
rect 6590 18490 6595 18510
rect 6565 18485 6595 18490
rect 6645 18510 6675 18515
rect 6645 18490 6650 18510
rect 6650 18490 6670 18510
rect 6670 18490 6675 18510
rect 6645 18485 6675 18490
rect 6725 18510 6755 18515
rect 6725 18490 6730 18510
rect 6730 18490 6750 18510
rect 6750 18490 6755 18510
rect 6725 18485 6755 18490
rect 6805 18510 6835 18515
rect 6805 18490 6810 18510
rect 6810 18490 6830 18510
rect 6830 18490 6835 18510
rect 6805 18485 6835 18490
rect 6885 18510 6915 18515
rect 6885 18490 6890 18510
rect 6890 18490 6910 18510
rect 6910 18490 6915 18510
rect 6885 18485 6915 18490
rect 6965 18510 6995 18515
rect 6965 18490 6970 18510
rect 6970 18490 6990 18510
rect 6990 18490 6995 18510
rect 6965 18485 6995 18490
rect 7045 18510 7075 18515
rect 7045 18490 7050 18510
rect 7050 18490 7070 18510
rect 7070 18490 7075 18510
rect 7045 18485 7075 18490
rect 7125 18510 7155 18515
rect 7125 18490 7130 18510
rect 7130 18490 7150 18510
rect 7150 18490 7155 18510
rect 7125 18485 7155 18490
rect 7205 18510 7235 18515
rect 7205 18490 7210 18510
rect 7210 18490 7230 18510
rect 7230 18490 7235 18510
rect 7205 18485 7235 18490
rect 7285 18510 7315 18515
rect 7285 18490 7290 18510
rect 7290 18490 7310 18510
rect 7310 18490 7315 18510
rect 7285 18485 7315 18490
rect 7365 18510 7395 18515
rect 7365 18490 7370 18510
rect 7370 18490 7390 18510
rect 7390 18490 7395 18510
rect 7365 18485 7395 18490
rect 7445 18510 7475 18515
rect 7445 18490 7450 18510
rect 7450 18490 7470 18510
rect 7470 18490 7475 18510
rect 7445 18485 7475 18490
rect 7525 18510 7555 18515
rect 7525 18490 7530 18510
rect 7530 18490 7550 18510
rect 7550 18490 7555 18510
rect 7525 18485 7555 18490
rect 7605 18510 7635 18515
rect 7605 18490 7610 18510
rect 7610 18490 7630 18510
rect 7630 18490 7635 18510
rect 7605 18485 7635 18490
rect 7685 18510 7715 18515
rect 7685 18490 7690 18510
rect 7690 18490 7710 18510
rect 7710 18490 7715 18510
rect 7685 18485 7715 18490
rect 7765 18510 7795 18515
rect 7765 18490 7770 18510
rect 7770 18490 7790 18510
rect 7790 18490 7795 18510
rect 7765 18485 7795 18490
rect 7845 18510 7875 18515
rect 7845 18490 7850 18510
rect 7850 18490 7870 18510
rect 7870 18490 7875 18510
rect 7845 18485 7875 18490
rect 7925 18510 7955 18515
rect 7925 18490 7930 18510
rect 7930 18490 7950 18510
rect 7950 18490 7955 18510
rect 7925 18485 7955 18490
rect 8005 18510 8035 18515
rect 8005 18490 8010 18510
rect 8010 18490 8030 18510
rect 8030 18490 8035 18510
rect 8005 18485 8035 18490
rect 8085 18510 8115 18515
rect 8085 18490 8090 18510
rect 8090 18490 8110 18510
rect 8110 18490 8115 18510
rect 8085 18485 8115 18490
rect 8165 18510 8195 18515
rect 8165 18490 8170 18510
rect 8170 18490 8190 18510
rect 8190 18490 8195 18510
rect 8165 18485 8195 18490
rect 8245 18510 8275 18515
rect 8245 18490 8250 18510
rect 8250 18490 8270 18510
rect 8270 18490 8275 18510
rect 8245 18485 8275 18490
rect 8325 18510 8355 18515
rect 8325 18490 8330 18510
rect 8330 18490 8350 18510
rect 8350 18490 8355 18510
rect 8325 18485 8355 18490
rect 8405 18510 8435 18515
rect 8405 18490 8410 18510
rect 8410 18490 8430 18510
rect 8430 18490 8435 18510
rect 8405 18485 8435 18490
rect 8485 18510 8515 18515
rect 8485 18490 8490 18510
rect 8490 18490 8510 18510
rect 8510 18490 8515 18510
rect 8485 18485 8515 18490
rect 8565 18510 8595 18515
rect 8565 18490 8570 18510
rect 8570 18490 8590 18510
rect 8590 18490 8595 18510
rect 8565 18485 8595 18490
rect 8645 18510 8675 18515
rect 8645 18490 8650 18510
rect 8650 18490 8670 18510
rect 8670 18490 8675 18510
rect 8645 18485 8675 18490
rect 8725 18510 8755 18515
rect 8725 18490 8730 18510
rect 8730 18490 8750 18510
rect 8750 18490 8755 18510
rect 8725 18485 8755 18490
rect 8805 18510 8835 18515
rect 8805 18490 8810 18510
rect 8810 18490 8830 18510
rect 8830 18490 8835 18510
rect 8805 18485 8835 18490
rect 8885 18510 8915 18515
rect 8885 18490 8890 18510
rect 8890 18490 8910 18510
rect 8910 18490 8915 18510
rect 8885 18485 8915 18490
rect 8965 18510 8995 18515
rect 8965 18490 8970 18510
rect 8970 18490 8990 18510
rect 8990 18490 8995 18510
rect 8965 18485 8995 18490
rect 9045 18510 9075 18515
rect 9045 18490 9050 18510
rect 9050 18490 9070 18510
rect 9070 18490 9075 18510
rect 9045 18485 9075 18490
rect 9125 18510 9155 18515
rect 9125 18490 9130 18510
rect 9130 18490 9150 18510
rect 9150 18490 9155 18510
rect 9125 18485 9155 18490
rect 9205 18510 9235 18515
rect 9205 18490 9210 18510
rect 9210 18490 9230 18510
rect 9230 18490 9235 18510
rect 9205 18485 9235 18490
rect 9285 18510 9315 18515
rect 9285 18490 9290 18510
rect 9290 18490 9310 18510
rect 9310 18490 9315 18510
rect 9285 18485 9315 18490
rect 9365 18510 9395 18515
rect 9365 18490 9370 18510
rect 9370 18490 9390 18510
rect 9390 18490 9395 18510
rect 9365 18485 9395 18490
rect 9445 18510 9475 18515
rect 9445 18490 9450 18510
rect 9450 18490 9470 18510
rect 9470 18490 9475 18510
rect 9445 18485 9475 18490
rect 11565 18510 11595 18515
rect 11565 18490 11570 18510
rect 11570 18490 11590 18510
rect 11590 18490 11595 18510
rect 11565 18485 11595 18490
rect 11645 18510 11675 18515
rect 11645 18490 11650 18510
rect 11650 18490 11670 18510
rect 11670 18490 11675 18510
rect 11645 18485 11675 18490
rect 11725 18510 11755 18515
rect 11725 18490 11730 18510
rect 11730 18490 11750 18510
rect 11750 18490 11755 18510
rect 11725 18485 11755 18490
rect 11805 18510 11835 18515
rect 11805 18490 11810 18510
rect 11810 18490 11830 18510
rect 11830 18490 11835 18510
rect 11805 18485 11835 18490
rect 11885 18510 11915 18515
rect 11885 18490 11890 18510
rect 11890 18490 11910 18510
rect 11910 18490 11915 18510
rect 11885 18485 11915 18490
rect 11965 18510 11995 18515
rect 11965 18490 11970 18510
rect 11970 18490 11990 18510
rect 11990 18490 11995 18510
rect 11965 18485 11995 18490
rect 12045 18510 12075 18515
rect 12045 18490 12050 18510
rect 12050 18490 12070 18510
rect 12070 18490 12075 18510
rect 12045 18485 12075 18490
rect 12125 18510 12155 18515
rect 12125 18490 12130 18510
rect 12130 18490 12150 18510
rect 12150 18490 12155 18510
rect 12125 18485 12155 18490
rect 12205 18510 12235 18515
rect 12205 18490 12210 18510
rect 12210 18490 12230 18510
rect 12230 18490 12235 18510
rect 12205 18485 12235 18490
rect 12285 18510 12315 18515
rect 12285 18490 12290 18510
rect 12290 18490 12310 18510
rect 12310 18490 12315 18510
rect 12285 18485 12315 18490
rect 12365 18510 12395 18515
rect 12365 18490 12370 18510
rect 12370 18490 12390 18510
rect 12390 18490 12395 18510
rect 12365 18485 12395 18490
rect 12445 18510 12475 18515
rect 12445 18490 12450 18510
rect 12450 18490 12470 18510
rect 12470 18490 12475 18510
rect 12445 18485 12475 18490
rect 12525 18510 12555 18515
rect 12525 18490 12530 18510
rect 12530 18490 12550 18510
rect 12550 18490 12555 18510
rect 12525 18485 12555 18490
rect 12605 18510 12635 18515
rect 12605 18490 12610 18510
rect 12610 18490 12630 18510
rect 12630 18490 12635 18510
rect 12605 18485 12635 18490
rect 12685 18510 12715 18515
rect 12685 18490 12690 18510
rect 12690 18490 12710 18510
rect 12710 18490 12715 18510
rect 12685 18485 12715 18490
rect 12765 18510 12795 18515
rect 12765 18490 12770 18510
rect 12770 18490 12790 18510
rect 12790 18490 12795 18510
rect 12765 18485 12795 18490
rect 12845 18510 12875 18515
rect 12845 18490 12850 18510
rect 12850 18490 12870 18510
rect 12870 18490 12875 18510
rect 12845 18485 12875 18490
rect 12925 18510 12955 18515
rect 12925 18490 12930 18510
rect 12930 18490 12950 18510
rect 12950 18490 12955 18510
rect 12925 18485 12955 18490
rect 13005 18510 13035 18515
rect 13005 18490 13010 18510
rect 13010 18490 13030 18510
rect 13030 18490 13035 18510
rect 13005 18485 13035 18490
rect 13085 18510 13115 18515
rect 13085 18490 13090 18510
rect 13090 18490 13110 18510
rect 13110 18490 13115 18510
rect 13085 18485 13115 18490
rect 13165 18510 13195 18515
rect 13165 18490 13170 18510
rect 13170 18490 13190 18510
rect 13190 18490 13195 18510
rect 13165 18485 13195 18490
rect 13245 18510 13275 18515
rect 13245 18490 13250 18510
rect 13250 18490 13270 18510
rect 13270 18490 13275 18510
rect 13245 18485 13275 18490
rect 13325 18510 13355 18515
rect 13325 18490 13330 18510
rect 13330 18490 13350 18510
rect 13350 18490 13355 18510
rect 13325 18485 13355 18490
rect 13405 18510 13435 18515
rect 13405 18490 13410 18510
rect 13410 18490 13430 18510
rect 13430 18490 13435 18510
rect 13405 18485 13435 18490
rect 13485 18510 13515 18515
rect 13485 18490 13490 18510
rect 13490 18490 13510 18510
rect 13510 18490 13515 18510
rect 13485 18485 13515 18490
rect 13565 18510 13595 18515
rect 13565 18490 13570 18510
rect 13570 18490 13590 18510
rect 13590 18490 13595 18510
rect 13565 18485 13595 18490
rect 13645 18510 13675 18515
rect 13645 18490 13650 18510
rect 13650 18490 13670 18510
rect 13670 18490 13675 18510
rect 13645 18485 13675 18490
rect 13725 18510 13755 18515
rect 13725 18490 13730 18510
rect 13730 18490 13750 18510
rect 13750 18490 13755 18510
rect 13725 18485 13755 18490
rect 13805 18510 13835 18515
rect 13805 18490 13810 18510
rect 13810 18490 13830 18510
rect 13830 18490 13835 18510
rect 13805 18485 13835 18490
rect 13885 18510 13915 18515
rect 13885 18490 13890 18510
rect 13890 18490 13910 18510
rect 13910 18490 13915 18510
rect 13885 18485 13915 18490
rect 13965 18510 13995 18515
rect 13965 18490 13970 18510
rect 13970 18490 13990 18510
rect 13990 18490 13995 18510
rect 13965 18485 13995 18490
rect 14045 18510 14075 18515
rect 14045 18490 14050 18510
rect 14050 18490 14070 18510
rect 14070 18490 14075 18510
rect 14045 18485 14075 18490
rect 14125 18510 14155 18515
rect 14125 18490 14130 18510
rect 14130 18490 14150 18510
rect 14150 18490 14155 18510
rect 14125 18485 14155 18490
rect 14205 18510 14235 18515
rect 14205 18490 14210 18510
rect 14210 18490 14230 18510
rect 14230 18490 14235 18510
rect 14205 18485 14235 18490
rect 14285 18510 14315 18515
rect 14285 18490 14290 18510
rect 14290 18490 14310 18510
rect 14310 18490 14315 18510
rect 14285 18485 14315 18490
rect 14365 18510 14395 18515
rect 14365 18490 14370 18510
rect 14370 18490 14390 18510
rect 14390 18490 14395 18510
rect 14365 18485 14395 18490
rect 14445 18510 14475 18515
rect 14445 18490 14450 18510
rect 14450 18490 14470 18510
rect 14470 18490 14475 18510
rect 14445 18485 14475 18490
rect 14525 18510 14555 18515
rect 14525 18490 14530 18510
rect 14530 18490 14550 18510
rect 14550 18490 14555 18510
rect 14525 18485 14555 18490
rect 14605 18510 14635 18515
rect 14605 18490 14610 18510
rect 14610 18490 14630 18510
rect 14630 18490 14635 18510
rect 14605 18485 14635 18490
rect 14685 18510 14715 18515
rect 14685 18490 14690 18510
rect 14690 18490 14710 18510
rect 14710 18490 14715 18510
rect 14685 18485 14715 18490
rect 16765 18510 16795 18515
rect 16765 18490 16770 18510
rect 16770 18490 16790 18510
rect 16790 18490 16795 18510
rect 16765 18485 16795 18490
rect 16845 18510 16875 18515
rect 16845 18490 16850 18510
rect 16850 18490 16870 18510
rect 16870 18490 16875 18510
rect 16845 18485 16875 18490
rect 16925 18510 16955 18515
rect 16925 18490 16930 18510
rect 16930 18490 16950 18510
rect 16950 18490 16955 18510
rect 16925 18485 16955 18490
rect 17005 18510 17035 18515
rect 17005 18490 17010 18510
rect 17010 18490 17030 18510
rect 17030 18490 17035 18510
rect 17005 18485 17035 18490
rect 17085 18510 17115 18515
rect 17085 18490 17090 18510
rect 17090 18490 17110 18510
rect 17110 18490 17115 18510
rect 17085 18485 17115 18490
rect 17165 18510 17195 18515
rect 17165 18490 17170 18510
rect 17170 18490 17190 18510
rect 17190 18490 17195 18510
rect 17165 18485 17195 18490
rect 17245 18510 17275 18515
rect 17245 18490 17250 18510
rect 17250 18490 17270 18510
rect 17270 18490 17275 18510
rect 17245 18485 17275 18490
rect 17325 18510 17355 18515
rect 17325 18490 17330 18510
rect 17330 18490 17350 18510
rect 17350 18490 17355 18510
rect 17325 18485 17355 18490
rect 17405 18510 17435 18515
rect 17405 18490 17410 18510
rect 17410 18490 17430 18510
rect 17430 18490 17435 18510
rect 17405 18485 17435 18490
rect 17485 18510 17515 18515
rect 17485 18490 17490 18510
rect 17490 18490 17510 18510
rect 17510 18490 17515 18510
rect 17485 18485 17515 18490
rect 17565 18510 17595 18515
rect 17565 18490 17570 18510
rect 17570 18490 17590 18510
rect 17590 18490 17595 18510
rect 17565 18485 17595 18490
rect 17645 18510 17675 18515
rect 17645 18490 17650 18510
rect 17650 18490 17670 18510
rect 17670 18490 17675 18510
rect 17645 18485 17675 18490
rect 17725 18510 17755 18515
rect 17725 18490 17730 18510
rect 17730 18490 17750 18510
rect 17750 18490 17755 18510
rect 17725 18485 17755 18490
rect 17805 18510 17835 18515
rect 17805 18490 17810 18510
rect 17810 18490 17830 18510
rect 17830 18490 17835 18510
rect 17805 18485 17835 18490
rect 17885 18510 17915 18515
rect 17885 18490 17890 18510
rect 17890 18490 17910 18510
rect 17910 18490 17915 18510
rect 17885 18485 17915 18490
rect 17965 18510 17995 18515
rect 17965 18490 17970 18510
rect 17970 18490 17990 18510
rect 17990 18490 17995 18510
rect 17965 18485 17995 18490
rect 18045 18510 18075 18515
rect 18045 18490 18050 18510
rect 18050 18490 18070 18510
rect 18070 18490 18075 18510
rect 18045 18485 18075 18490
rect 18125 18510 18155 18515
rect 18125 18490 18130 18510
rect 18130 18490 18150 18510
rect 18150 18490 18155 18510
rect 18125 18485 18155 18490
rect 18205 18510 18235 18515
rect 18205 18490 18210 18510
rect 18210 18490 18230 18510
rect 18230 18490 18235 18510
rect 18205 18485 18235 18490
rect 18285 18510 18315 18515
rect 18285 18490 18290 18510
rect 18290 18490 18310 18510
rect 18310 18490 18315 18510
rect 18285 18485 18315 18490
rect 18365 18510 18395 18515
rect 18365 18490 18370 18510
rect 18370 18490 18390 18510
rect 18390 18490 18395 18510
rect 18365 18485 18395 18490
rect 18445 18510 18475 18515
rect 18445 18490 18450 18510
rect 18450 18490 18470 18510
rect 18470 18490 18475 18510
rect 18445 18485 18475 18490
rect 18525 18510 18555 18515
rect 18525 18490 18530 18510
rect 18530 18490 18550 18510
rect 18550 18490 18555 18510
rect 18525 18485 18555 18490
rect 18605 18510 18635 18515
rect 18605 18490 18610 18510
rect 18610 18490 18630 18510
rect 18630 18490 18635 18510
rect 18605 18485 18635 18490
rect 18685 18510 18715 18515
rect 18685 18490 18690 18510
rect 18690 18490 18710 18510
rect 18710 18490 18715 18510
rect 18685 18485 18715 18490
rect 18765 18510 18795 18515
rect 18765 18490 18770 18510
rect 18770 18490 18790 18510
rect 18790 18490 18795 18510
rect 18765 18485 18795 18490
rect 18845 18510 18875 18515
rect 18845 18490 18850 18510
rect 18850 18490 18870 18510
rect 18870 18490 18875 18510
rect 18845 18485 18875 18490
rect 18925 18510 18955 18515
rect 18925 18490 18930 18510
rect 18930 18490 18950 18510
rect 18950 18490 18955 18510
rect 18925 18485 18955 18490
rect 19005 18510 19035 18515
rect 19005 18490 19010 18510
rect 19010 18490 19030 18510
rect 19030 18490 19035 18510
rect 19005 18485 19035 18490
rect 19085 18510 19115 18515
rect 19085 18490 19090 18510
rect 19090 18490 19110 18510
rect 19110 18490 19115 18510
rect 19085 18485 19115 18490
rect 19165 18510 19195 18515
rect 19165 18490 19170 18510
rect 19170 18490 19190 18510
rect 19190 18490 19195 18510
rect 19165 18485 19195 18490
rect 19245 18510 19275 18515
rect 19245 18490 19250 18510
rect 19250 18490 19270 18510
rect 19270 18490 19275 18510
rect 19245 18485 19275 18490
rect 19325 18510 19355 18515
rect 19325 18490 19330 18510
rect 19330 18490 19350 18510
rect 19350 18490 19355 18510
rect 19325 18485 19355 18490
rect 19405 18510 19435 18515
rect 19405 18490 19410 18510
rect 19410 18490 19430 18510
rect 19430 18490 19435 18510
rect 19405 18485 19435 18490
rect 19485 18510 19515 18515
rect 19485 18490 19490 18510
rect 19490 18490 19510 18510
rect 19510 18490 19515 18510
rect 19485 18485 19515 18490
rect 19565 18510 19595 18515
rect 19565 18490 19570 18510
rect 19570 18490 19590 18510
rect 19590 18490 19595 18510
rect 19565 18485 19595 18490
rect 19645 18510 19675 18515
rect 19645 18490 19650 18510
rect 19650 18490 19670 18510
rect 19670 18490 19675 18510
rect 19645 18485 19675 18490
rect 19725 18510 19755 18515
rect 19725 18490 19730 18510
rect 19730 18490 19750 18510
rect 19750 18490 19755 18510
rect 19725 18485 19755 18490
rect 19805 18510 19835 18515
rect 19805 18490 19810 18510
rect 19810 18490 19830 18510
rect 19830 18490 19835 18510
rect 19805 18485 19835 18490
rect 19885 18510 19915 18515
rect 19885 18490 19890 18510
rect 19890 18490 19910 18510
rect 19910 18490 19915 18510
rect 19885 18485 19915 18490
rect 19965 18510 19995 18515
rect 19965 18490 19970 18510
rect 19970 18490 19990 18510
rect 19990 18490 19995 18510
rect 19965 18485 19995 18490
rect 20045 18510 20075 18515
rect 20045 18490 20050 18510
rect 20050 18490 20070 18510
rect 20070 18490 20075 18510
rect 20045 18485 20075 18490
rect 20125 18510 20155 18515
rect 20125 18490 20130 18510
rect 20130 18490 20150 18510
rect 20150 18490 20155 18510
rect 20125 18485 20155 18490
rect 20205 18510 20235 18515
rect 20205 18490 20210 18510
rect 20210 18490 20230 18510
rect 20230 18490 20235 18510
rect 20205 18485 20235 18490
rect 20285 18510 20315 18515
rect 20285 18490 20290 18510
rect 20290 18490 20310 18510
rect 20310 18490 20315 18510
rect 20285 18485 20315 18490
rect 20365 18510 20395 18515
rect 20365 18490 20370 18510
rect 20370 18490 20390 18510
rect 20390 18490 20395 18510
rect 20365 18485 20395 18490
rect 20445 18510 20475 18515
rect 20445 18490 20450 18510
rect 20450 18490 20470 18510
rect 20470 18490 20475 18510
rect 20445 18485 20475 18490
rect 20525 18510 20555 18515
rect 20525 18490 20530 18510
rect 20530 18490 20550 18510
rect 20550 18490 20555 18510
rect 20525 18485 20555 18490
rect 20605 18510 20635 18515
rect 20605 18490 20610 18510
rect 20610 18490 20630 18510
rect 20630 18490 20635 18510
rect 20605 18485 20635 18490
rect 20685 18510 20715 18515
rect 20685 18490 20690 18510
rect 20690 18490 20710 18510
rect 20710 18490 20715 18510
rect 20685 18485 20715 18490
rect 20765 18510 20795 18515
rect 20765 18490 20770 18510
rect 20770 18490 20790 18510
rect 20790 18490 20795 18510
rect 20765 18485 20795 18490
rect 20845 18510 20875 18515
rect 20845 18490 20850 18510
rect 20850 18490 20870 18510
rect 20870 18490 20875 18510
rect 20845 18485 20875 18490
rect 20925 18510 20955 18515
rect 20925 18490 20930 18510
rect 20930 18490 20950 18510
rect 20950 18490 20955 18510
rect 20925 18485 20955 18490
rect 5 18430 35 18435
rect 5 18410 10 18430
rect 10 18410 30 18430
rect 30 18410 35 18430
rect 5 18405 35 18410
rect 85 18430 115 18435
rect 85 18410 90 18430
rect 90 18410 110 18430
rect 110 18410 115 18430
rect 85 18405 115 18410
rect 165 18430 195 18435
rect 165 18410 170 18430
rect 170 18410 190 18430
rect 190 18410 195 18430
rect 165 18405 195 18410
rect 245 18430 275 18435
rect 245 18410 250 18430
rect 250 18410 270 18430
rect 270 18410 275 18430
rect 245 18405 275 18410
rect 325 18430 355 18435
rect 325 18410 330 18430
rect 330 18410 350 18430
rect 350 18410 355 18430
rect 325 18405 355 18410
rect 405 18430 435 18435
rect 405 18410 410 18430
rect 410 18410 430 18430
rect 430 18410 435 18430
rect 405 18405 435 18410
rect 485 18430 515 18435
rect 485 18410 490 18430
rect 490 18410 510 18430
rect 510 18410 515 18430
rect 485 18405 515 18410
rect 565 18430 595 18435
rect 565 18410 570 18430
rect 570 18410 590 18430
rect 590 18410 595 18430
rect 565 18405 595 18410
rect 645 18430 675 18435
rect 645 18410 650 18430
rect 650 18410 670 18430
rect 670 18410 675 18430
rect 645 18405 675 18410
rect 725 18430 755 18435
rect 725 18410 730 18430
rect 730 18410 750 18430
rect 750 18410 755 18430
rect 725 18405 755 18410
rect 805 18430 835 18435
rect 805 18410 810 18430
rect 810 18410 830 18430
rect 830 18410 835 18430
rect 805 18405 835 18410
rect 885 18430 915 18435
rect 885 18410 890 18430
rect 890 18410 910 18430
rect 910 18410 915 18430
rect 885 18405 915 18410
rect 965 18430 995 18435
rect 965 18410 970 18430
rect 970 18410 990 18430
rect 990 18410 995 18430
rect 965 18405 995 18410
rect 1045 18430 1075 18435
rect 1045 18410 1050 18430
rect 1050 18410 1070 18430
rect 1070 18410 1075 18430
rect 1045 18405 1075 18410
rect 1125 18430 1155 18435
rect 1125 18410 1130 18430
rect 1130 18410 1150 18430
rect 1150 18410 1155 18430
rect 1125 18405 1155 18410
rect 1205 18430 1235 18435
rect 1205 18410 1210 18430
rect 1210 18410 1230 18430
rect 1230 18410 1235 18430
rect 1205 18405 1235 18410
rect 1285 18430 1315 18435
rect 1285 18410 1290 18430
rect 1290 18410 1310 18430
rect 1310 18410 1315 18430
rect 1285 18405 1315 18410
rect 1365 18430 1395 18435
rect 1365 18410 1370 18430
rect 1370 18410 1390 18430
rect 1390 18410 1395 18430
rect 1365 18405 1395 18410
rect 1445 18430 1475 18435
rect 1445 18410 1450 18430
rect 1450 18410 1470 18430
rect 1470 18410 1475 18430
rect 1445 18405 1475 18410
rect 1525 18430 1555 18435
rect 1525 18410 1530 18430
rect 1530 18410 1550 18430
rect 1550 18410 1555 18430
rect 1525 18405 1555 18410
rect 1605 18430 1635 18435
rect 1605 18410 1610 18430
rect 1610 18410 1630 18430
rect 1630 18410 1635 18430
rect 1605 18405 1635 18410
rect 1685 18430 1715 18435
rect 1685 18410 1690 18430
rect 1690 18410 1710 18430
rect 1710 18410 1715 18430
rect 1685 18405 1715 18410
rect 1765 18430 1795 18435
rect 1765 18410 1770 18430
rect 1770 18410 1790 18430
rect 1790 18410 1795 18430
rect 1765 18405 1795 18410
rect 1845 18430 1875 18435
rect 1845 18410 1850 18430
rect 1850 18410 1870 18430
rect 1870 18410 1875 18430
rect 1845 18405 1875 18410
rect 1925 18430 1955 18435
rect 1925 18410 1930 18430
rect 1930 18410 1950 18430
rect 1950 18410 1955 18430
rect 1925 18405 1955 18410
rect 2005 18430 2035 18435
rect 2005 18410 2010 18430
rect 2010 18410 2030 18430
rect 2030 18410 2035 18430
rect 2005 18405 2035 18410
rect 2085 18430 2115 18435
rect 2085 18410 2090 18430
rect 2090 18410 2110 18430
rect 2110 18410 2115 18430
rect 2085 18405 2115 18410
rect 2165 18430 2195 18435
rect 2165 18410 2170 18430
rect 2170 18410 2190 18430
rect 2190 18410 2195 18430
rect 2165 18405 2195 18410
rect 2245 18430 2275 18435
rect 2245 18410 2250 18430
rect 2250 18410 2270 18430
rect 2270 18410 2275 18430
rect 2245 18405 2275 18410
rect 2325 18430 2355 18435
rect 2325 18410 2330 18430
rect 2330 18410 2350 18430
rect 2350 18410 2355 18430
rect 2325 18405 2355 18410
rect 2405 18430 2435 18435
rect 2405 18410 2410 18430
rect 2410 18410 2430 18430
rect 2430 18410 2435 18430
rect 2405 18405 2435 18410
rect 2485 18430 2515 18435
rect 2485 18410 2490 18430
rect 2490 18410 2510 18430
rect 2510 18410 2515 18430
rect 2485 18405 2515 18410
rect 2565 18430 2595 18435
rect 2565 18410 2570 18430
rect 2570 18410 2590 18430
rect 2590 18410 2595 18430
rect 2565 18405 2595 18410
rect 2645 18430 2675 18435
rect 2645 18410 2650 18430
rect 2650 18410 2670 18430
rect 2670 18410 2675 18430
rect 2645 18405 2675 18410
rect 2725 18430 2755 18435
rect 2725 18410 2730 18430
rect 2730 18410 2750 18430
rect 2750 18410 2755 18430
rect 2725 18405 2755 18410
rect 2805 18430 2835 18435
rect 2805 18410 2810 18430
rect 2810 18410 2830 18430
rect 2830 18410 2835 18430
rect 2805 18405 2835 18410
rect 2885 18430 2915 18435
rect 2885 18410 2890 18430
rect 2890 18410 2910 18430
rect 2910 18410 2915 18430
rect 2885 18405 2915 18410
rect 2965 18430 2995 18435
rect 2965 18410 2970 18430
rect 2970 18410 2990 18430
rect 2990 18410 2995 18430
rect 2965 18405 2995 18410
rect 3045 18430 3075 18435
rect 3045 18410 3050 18430
rect 3050 18410 3070 18430
rect 3070 18410 3075 18430
rect 3045 18405 3075 18410
rect 3125 18430 3155 18435
rect 3125 18410 3130 18430
rect 3130 18410 3150 18430
rect 3150 18410 3155 18430
rect 3125 18405 3155 18410
rect 3205 18430 3235 18435
rect 3205 18410 3210 18430
rect 3210 18410 3230 18430
rect 3230 18410 3235 18430
rect 3205 18405 3235 18410
rect 3285 18430 3315 18435
rect 3285 18410 3290 18430
rect 3290 18410 3310 18430
rect 3310 18410 3315 18430
rect 3285 18405 3315 18410
rect 3365 18430 3395 18435
rect 3365 18410 3370 18430
rect 3370 18410 3390 18430
rect 3390 18410 3395 18430
rect 3365 18405 3395 18410
rect 3445 18430 3475 18435
rect 3445 18410 3450 18430
rect 3450 18410 3470 18430
rect 3470 18410 3475 18430
rect 3445 18405 3475 18410
rect 3525 18430 3555 18435
rect 3525 18410 3530 18430
rect 3530 18410 3550 18430
rect 3550 18410 3555 18430
rect 3525 18405 3555 18410
rect 3605 18430 3635 18435
rect 3605 18410 3610 18430
rect 3610 18410 3630 18430
rect 3630 18410 3635 18430
rect 3605 18405 3635 18410
rect 3685 18430 3715 18435
rect 3685 18410 3690 18430
rect 3690 18410 3710 18430
rect 3710 18410 3715 18430
rect 3685 18405 3715 18410
rect 3765 18430 3795 18435
rect 3765 18410 3770 18430
rect 3770 18410 3790 18430
rect 3790 18410 3795 18430
rect 3765 18405 3795 18410
rect 3845 18430 3875 18435
rect 3845 18410 3850 18430
rect 3850 18410 3870 18430
rect 3870 18410 3875 18430
rect 3845 18405 3875 18410
rect 3925 18430 3955 18435
rect 3925 18410 3930 18430
rect 3930 18410 3950 18430
rect 3950 18410 3955 18430
rect 3925 18405 3955 18410
rect 4005 18430 4035 18435
rect 4005 18410 4010 18430
rect 4010 18410 4030 18430
rect 4030 18410 4035 18430
rect 4005 18405 4035 18410
rect 4085 18430 4115 18435
rect 4085 18410 4090 18430
rect 4090 18410 4110 18430
rect 4110 18410 4115 18430
rect 4085 18405 4115 18410
rect 4165 18430 4195 18435
rect 4165 18410 4170 18430
rect 4170 18410 4190 18430
rect 4190 18410 4195 18430
rect 4165 18405 4195 18410
rect 6245 18430 6275 18435
rect 6245 18410 6250 18430
rect 6250 18410 6270 18430
rect 6270 18410 6275 18430
rect 6245 18405 6275 18410
rect 6325 18430 6355 18435
rect 6325 18410 6330 18430
rect 6330 18410 6350 18430
rect 6350 18410 6355 18430
rect 6325 18405 6355 18410
rect 6405 18430 6435 18435
rect 6405 18410 6410 18430
rect 6410 18410 6430 18430
rect 6430 18410 6435 18430
rect 6405 18405 6435 18410
rect 6485 18430 6515 18435
rect 6485 18410 6490 18430
rect 6490 18410 6510 18430
rect 6510 18410 6515 18430
rect 6485 18405 6515 18410
rect 6565 18430 6595 18435
rect 6565 18410 6570 18430
rect 6570 18410 6590 18430
rect 6590 18410 6595 18430
rect 6565 18405 6595 18410
rect 6645 18430 6675 18435
rect 6645 18410 6650 18430
rect 6650 18410 6670 18430
rect 6670 18410 6675 18430
rect 6645 18405 6675 18410
rect 6725 18430 6755 18435
rect 6725 18410 6730 18430
rect 6730 18410 6750 18430
rect 6750 18410 6755 18430
rect 6725 18405 6755 18410
rect 6805 18430 6835 18435
rect 6805 18410 6810 18430
rect 6810 18410 6830 18430
rect 6830 18410 6835 18430
rect 6805 18405 6835 18410
rect 6885 18430 6915 18435
rect 6885 18410 6890 18430
rect 6890 18410 6910 18430
rect 6910 18410 6915 18430
rect 6885 18405 6915 18410
rect 6965 18430 6995 18435
rect 6965 18410 6970 18430
rect 6970 18410 6990 18430
rect 6990 18410 6995 18430
rect 6965 18405 6995 18410
rect 7045 18430 7075 18435
rect 7045 18410 7050 18430
rect 7050 18410 7070 18430
rect 7070 18410 7075 18430
rect 7045 18405 7075 18410
rect 7125 18430 7155 18435
rect 7125 18410 7130 18430
rect 7130 18410 7150 18430
rect 7150 18410 7155 18430
rect 7125 18405 7155 18410
rect 7205 18430 7235 18435
rect 7205 18410 7210 18430
rect 7210 18410 7230 18430
rect 7230 18410 7235 18430
rect 7205 18405 7235 18410
rect 7285 18430 7315 18435
rect 7285 18410 7290 18430
rect 7290 18410 7310 18430
rect 7310 18410 7315 18430
rect 7285 18405 7315 18410
rect 7365 18430 7395 18435
rect 7365 18410 7370 18430
rect 7370 18410 7390 18430
rect 7390 18410 7395 18430
rect 7365 18405 7395 18410
rect 7445 18430 7475 18435
rect 7445 18410 7450 18430
rect 7450 18410 7470 18430
rect 7470 18410 7475 18430
rect 7445 18405 7475 18410
rect 7525 18430 7555 18435
rect 7525 18410 7530 18430
rect 7530 18410 7550 18430
rect 7550 18410 7555 18430
rect 7525 18405 7555 18410
rect 7605 18430 7635 18435
rect 7605 18410 7610 18430
rect 7610 18410 7630 18430
rect 7630 18410 7635 18430
rect 7605 18405 7635 18410
rect 7685 18430 7715 18435
rect 7685 18410 7690 18430
rect 7690 18410 7710 18430
rect 7710 18410 7715 18430
rect 7685 18405 7715 18410
rect 7765 18430 7795 18435
rect 7765 18410 7770 18430
rect 7770 18410 7790 18430
rect 7790 18410 7795 18430
rect 7765 18405 7795 18410
rect 7845 18430 7875 18435
rect 7845 18410 7850 18430
rect 7850 18410 7870 18430
rect 7870 18410 7875 18430
rect 7845 18405 7875 18410
rect 7925 18430 7955 18435
rect 7925 18410 7930 18430
rect 7930 18410 7950 18430
rect 7950 18410 7955 18430
rect 7925 18405 7955 18410
rect 8005 18430 8035 18435
rect 8005 18410 8010 18430
rect 8010 18410 8030 18430
rect 8030 18410 8035 18430
rect 8005 18405 8035 18410
rect 8085 18430 8115 18435
rect 8085 18410 8090 18430
rect 8090 18410 8110 18430
rect 8110 18410 8115 18430
rect 8085 18405 8115 18410
rect 8165 18430 8195 18435
rect 8165 18410 8170 18430
rect 8170 18410 8190 18430
rect 8190 18410 8195 18430
rect 8165 18405 8195 18410
rect 8245 18430 8275 18435
rect 8245 18410 8250 18430
rect 8250 18410 8270 18430
rect 8270 18410 8275 18430
rect 8245 18405 8275 18410
rect 8325 18430 8355 18435
rect 8325 18410 8330 18430
rect 8330 18410 8350 18430
rect 8350 18410 8355 18430
rect 8325 18405 8355 18410
rect 8405 18430 8435 18435
rect 8405 18410 8410 18430
rect 8410 18410 8430 18430
rect 8430 18410 8435 18430
rect 8405 18405 8435 18410
rect 8485 18430 8515 18435
rect 8485 18410 8490 18430
rect 8490 18410 8510 18430
rect 8510 18410 8515 18430
rect 8485 18405 8515 18410
rect 8565 18430 8595 18435
rect 8565 18410 8570 18430
rect 8570 18410 8590 18430
rect 8590 18410 8595 18430
rect 8565 18405 8595 18410
rect 8645 18430 8675 18435
rect 8645 18410 8650 18430
rect 8650 18410 8670 18430
rect 8670 18410 8675 18430
rect 8645 18405 8675 18410
rect 8725 18430 8755 18435
rect 8725 18410 8730 18430
rect 8730 18410 8750 18430
rect 8750 18410 8755 18430
rect 8725 18405 8755 18410
rect 8805 18430 8835 18435
rect 8805 18410 8810 18430
rect 8810 18410 8830 18430
rect 8830 18410 8835 18430
rect 8805 18405 8835 18410
rect 8885 18430 8915 18435
rect 8885 18410 8890 18430
rect 8890 18410 8910 18430
rect 8910 18410 8915 18430
rect 8885 18405 8915 18410
rect 8965 18430 8995 18435
rect 8965 18410 8970 18430
rect 8970 18410 8990 18430
rect 8990 18410 8995 18430
rect 8965 18405 8995 18410
rect 9045 18430 9075 18435
rect 9045 18410 9050 18430
rect 9050 18410 9070 18430
rect 9070 18410 9075 18430
rect 9045 18405 9075 18410
rect 9125 18430 9155 18435
rect 9125 18410 9130 18430
rect 9130 18410 9150 18430
rect 9150 18410 9155 18430
rect 9125 18405 9155 18410
rect 9205 18430 9235 18435
rect 9205 18410 9210 18430
rect 9210 18410 9230 18430
rect 9230 18410 9235 18430
rect 9205 18405 9235 18410
rect 9285 18430 9315 18435
rect 9285 18410 9290 18430
rect 9290 18410 9310 18430
rect 9310 18410 9315 18430
rect 9285 18405 9315 18410
rect 9365 18430 9395 18435
rect 9365 18410 9370 18430
rect 9370 18410 9390 18430
rect 9390 18410 9395 18430
rect 9365 18405 9395 18410
rect 9445 18430 9475 18435
rect 9445 18410 9450 18430
rect 9450 18410 9470 18430
rect 9470 18410 9475 18430
rect 9445 18405 9475 18410
rect 11565 18430 11595 18435
rect 11565 18410 11570 18430
rect 11570 18410 11590 18430
rect 11590 18410 11595 18430
rect 11565 18405 11595 18410
rect 11645 18430 11675 18435
rect 11645 18410 11650 18430
rect 11650 18410 11670 18430
rect 11670 18410 11675 18430
rect 11645 18405 11675 18410
rect 11725 18430 11755 18435
rect 11725 18410 11730 18430
rect 11730 18410 11750 18430
rect 11750 18410 11755 18430
rect 11725 18405 11755 18410
rect 11805 18430 11835 18435
rect 11805 18410 11810 18430
rect 11810 18410 11830 18430
rect 11830 18410 11835 18430
rect 11805 18405 11835 18410
rect 11885 18430 11915 18435
rect 11885 18410 11890 18430
rect 11890 18410 11910 18430
rect 11910 18410 11915 18430
rect 11885 18405 11915 18410
rect 11965 18430 11995 18435
rect 11965 18410 11970 18430
rect 11970 18410 11990 18430
rect 11990 18410 11995 18430
rect 11965 18405 11995 18410
rect 12045 18430 12075 18435
rect 12045 18410 12050 18430
rect 12050 18410 12070 18430
rect 12070 18410 12075 18430
rect 12045 18405 12075 18410
rect 12125 18430 12155 18435
rect 12125 18410 12130 18430
rect 12130 18410 12150 18430
rect 12150 18410 12155 18430
rect 12125 18405 12155 18410
rect 12205 18430 12235 18435
rect 12205 18410 12210 18430
rect 12210 18410 12230 18430
rect 12230 18410 12235 18430
rect 12205 18405 12235 18410
rect 12285 18430 12315 18435
rect 12285 18410 12290 18430
rect 12290 18410 12310 18430
rect 12310 18410 12315 18430
rect 12285 18405 12315 18410
rect 12365 18430 12395 18435
rect 12365 18410 12370 18430
rect 12370 18410 12390 18430
rect 12390 18410 12395 18430
rect 12365 18405 12395 18410
rect 12445 18430 12475 18435
rect 12445 18410 12450 18430
rect 12450 18410 12470 18430
rect 12470 18410 12475 18430
rect 12445 18405 12475 18410
rect 12525 18430 12555 18435
rect 12525 18410 12530 18430
rect 12530 18410 12550 18430
rect 12550 18410 12555 18430
rect 12525 18405 12555 18410
rect 12605 18430 12635 18435
rect 12605 18410 12610 18430
rect 12610 18410 12630 18430
rect 12630 18410 12635 18430
rect 12605 18405 12635 18410
rect 12685 18430 12715 18435
rect 12685 18410 12690 18430
rect 12690 18410 12710 18430
rect 12710 18410 12715 18430
rect 12685 18405 12715 18410
rect 12765 18430 12795 18435
rect 12765 18410 12770 18430
rect 12770 18410 12790 18430
rect 12790 18410 12795 18430
rect 12765 18405 12795 18410
rect 12845 18430 12875 18435
rect 12845 18410 12850 18430
rect 12850 18410 12870 18430
rect 12870 18410 12875 18430
rect 12845 18405 12875 18410
rect 12925 18430 12955 18435
rect 12925 18410 12930 18430
rect 12930 18410 12950 18430
rect 12950 18410 12955 18430
rect 12925 18405 12955 18410
rect 13005 18430 13035 18435
rect 13005 18410 13010 18430
rect 13010 18410 13030 18430
rect 13030 18410 13035 18430
rect 13005 18405 13035 18410
rect 13085 18430 13115 18435
rect 13085 18410 13090 18430
rect 13090 18410 13110 18430
rect 13110 18410 13115 18430
rect 13085 18405 13115 18410
rect 13165 18430 13195 18435
rect 13165 18410 13170 18430
rect 13170 18410 13190 18430
rect 13190 18410 13195 18430
rect 13165 18405 13195 18410
rect 13245 18430 13275 18435
rect 13245 18410 13250 18430
rect 13250 18410 13270 18430
rect 13270 18410 13275 18430
rect 13245 18405 13275 18410
rect 13325 18430 13355 18435
rect 13325 18410 13330 18430
rect 13330 18410 13350 18430
rect 13350 18410 13355 18430
rect 13325 18405 13355 18410
rect 13405 18430 13435 18435
rect 13405 18410 13410 18430
rect 13410 18410 13430 18430
rect 13430 18410 13435 18430
rect 13405 18405 13435 18410
rect 13485 18430 13515 18435
rect 13485 18410 13490 18430
rect 13490 18410 13510 18430
rect 13510 18410 13515 18430
rect 13485 18405 13515 18410
rect 13565 18430 13595 18435
rect 13565 18410 13570 18430
rect 13570 18410 13590 18430
rect 13590 18410 13595 18430
rect 13565 18405 13595 18410
rect 13645 18430 13675 18435
rect 13645 18410 13650 18430
rect 13650 18410 13670 18430
rect 13670 18410 13675 18430
rect 13645 18405 13675 18410
rect 13725 18430 13755 18435
rect 13725 18410 13730 18430
rect 13730 18410 13750 18430
rect 13750 18410 13755 18430
rect 13725 18405 13755 18410
rect 13805 18430 13835 18435
rect 13805 18410 13810 18430
rect 13810 18410 13830 18430
rect 13830 18410 13835 18430
rect 13805 18405 13835 18410
rect 13885 18430 13915 18435
rect 13885 18410 13890 18430
rect 13890 18410 13910 18430
rect 13910 18410 13915 18430
rect 13885 18405 13915 18410
rect 13965 18430 13995 18435
rect 13965 18410 13970 18430
rect 13970 18410 13990 18430
rect 13990 18410 13995 18430
rect 13965 18405 13995 18410
rect 14045 18430 14075 18435
rect 14045 18410 14050 18430
rect 14050 18410 14070 18430
rect 14070 18410 14075 18430
rect 14045 18405 14075 18410
rect 14125 18430 14155 18435
rect 14125 18410 14130 18430
rect 14130 18410 14150 18430
rect 14150 18410 14155 18430
rect 14125 18405 14155 18410
rect 14205 18430 14235 18435
rect 14205 18410 14210 18430
rect 14210 18410 14230 18430
rect 14230 18410 14235 18430
rect 14205 18405 14235 18410
rect 14285 18430 14315 18435
rect 14285 18410 14290 18430
rect 14290 18410 14310 18430
rect 14310 18410 14315 18430
rect 14285 18405 14315 18410
rect 14365 18430 14395 18435
rect 14365 18410 14370 18430
rect 14370 18410 14390 18430
rect 14390 18410 14395 18430
rect 14365 18405 14395 18410
rect 14445 18430 14475 18435
rect 14445 18410 14450 18430
rect 14450 18410 14470 18430
rect 14470 18410 14475 18430
rect 14445 18405 14475 18410
rect 14525 18430 14555 18435
rect 14525 18410 14530 18430
rect 14530 18410 14550 18430
rect 14550 18410 14555 18430
rect 14525 18405 14555 18410
rect 14605 18430 14635 18435
rect 14605 18410 14610 18430
rect 14610 18410 14630 18430
rect 14630 18410 14635 18430
rect 14605 18405 14635 18410
rect 14685 18430 14715 18435
rect 14685 18410 14690 18430
rect 14690 18410 14710 18430
rect 14710 18410 14715 18430
rect 14685 18405 14715 18410
rect 16765 18430 16795 18435
rect 16765 18410 16770 18430
rect 16770 18410 16790 18430
rect 16790 18410 16795 18430
rect 16765 18405 16795 18410
rect 16845 18430 16875 18435
rect 16845 18410 16850 18430
rect 16850 18410 16870 18430
rect 16870 18410 16875 18430
rect 16845 18405 16875 18410
rect 16925 18430 16955 18435
rect 16925 18410 16930 18430
rect 16930 18410 16950 18430
rect 16950 18410 16955 18430
rect 16925 18405 16955 18410
rect 17005 18430 17035 18435
rect 17005 18410 17010 18430
rect 17010 18410 17030 18430
rect 17030 18410 17035 18430
rect 17005 18405 17035 18410
rect 17085 18430 17115 18435
rect 17085 18410 17090 18430
rect 17090 18410 17110 18430
rect 17110 18410 17115 18430
rect 17085 18405 17115 18410
rect 17165 18430 17195 18435
rect 17165 18410 17170 18430
rect 17170 18410 17190 18430
rect 17190 18410 17195 18430
rect 17165 18405 17195 18410
rect 17245 18430 17275 18435
rect 17245 18410 17250 18430
rect 17250 18410 17270 18430
rect 17270 18410 17275 18430
rect 17245 18405 17275 18410
rect 17325 18430 17355 18435
rect 17325 18410 17330 18430
rect 17330 18410 17350 18430
rect 17350 18410 17355 18430
rect 17325 18405 17355 18410
rect 17405 18430 17435 18435
rect 17405 18410 17410 18430
rect 17410 18410 17430 18430
rect 17430 18410 17435 18430
rect 17405 18405 17435 18410
rect 17485 18430 17515 18435
rect 17485 18410 17490 18430
rect 17490 18410 17510 18430
rect 17510 18410 17515 18430
rect 17485 18405 17515 18410
rect 17565 18430 17595 18435
rect 17565 18410 17570 18430
rect 17570 18410 17590 18430
rect 17590 18410 17595 18430
rect 17565 18405 17595 18410
rect 17645 18430 17675 18435
rect 17645 18410 17650 18430
rect 17650 18410 17670 18430
rect 17670 18410 17675 18430
rect 17645 18405 17675 18410
rect 17725 18430 17755 18435
rect 17725 18410 17730 18430
rect 17730 18410 17750 18430
rect 17750 18410 17755 18430
rect 17725 18405 17755 18410
rect 17805 18430 17835 18435
rect 17805 18410 17810 18430
rect 17810 18410 17830 18430
rect 17830 18410 17835 18430
rect 17805 18405 17835 18410
rect 17885 18430 17915 18435
rect 17885 18410 17890 18430
rect 17890 18410 17910 18430
rect 17910 18410 17915 18430
rect 17885 18405 17915 18410
rect 17965 18430 17995 18435
rect 17965 18410 17970 18430
rect 17970 18410 17990 18430
rect 17990 18410 17995 18430
rect 17965 18405 17995 18410
rect 18045 18430 18075 18435
rect 18045 18410 18050 18430
rect 18050 18410 18070 18430
rect 18070 18410 18075 18430
rect 18045 18405 18075 18410
rect 18125 18430 18155 18435
rect 18125 18410 18130 18430
rect 18130 18410 18150 18430
rect 18150 18410 18155 18430
rect 18125 18405 18155 18410
rect 18205 18430 18235 18435
rect 18205 18410 18210 18430
rect 18210 18410 18230 18430
rect 18230 18410 18235 18430
rect 18205 18405 18235 18410
rect 18285 18430 18315 18435
rect 18285 18410 18290 18430
rect 18290 18410 18310 18430
rect 18310 18410 18315 18430
rect 18285 18405 18315 18410
rect 18365 18430 18395 18435
rect 18365 18410 18370 18430
rect 18370 18410 18390 18430
rect 18390 18410 18395 18430
rect 18365 18405 18395 18410
rect 18445 18430 18475 18435
rect 18445 18410 18450 18430
rect 18450 18410 18470 18430
rect 18470 18410 18475 18430
rect 18445 18405 18475 18410
rect 18525 18430 18555 18435
rect 18525 18410 18530 18430
rect 18530 18410 18550 18430
rect 18550 18410 18555 18430
rect 18525 18405 18555 18410
rect 18605 18430 18635 18435
rect 18605 18410 18610 18430
rect 18610 18410 18630 18430
rect 18630 18410 18635 18430
rect 18605 18405 18635 18410
rect 18685 18430 18715 18435
rect 18685 18410 18690 18430
rect 18690 18410 18710 18430
rect 18710 18410 18715 18430
rect 18685 18405 18715 18410
rect 18765 18430 18795 18435
rect 18765 18410 18770 18430
rect 18770 18410 18790 18430
rect 18790 18410 18795 18430
rect 18765 18405 18795 18410
rect 18845 18430 18875 18435
rect 18845 18410 18850 18430
rect 18850 18410 18870 18430
rect 18870 18410 18875 18430
rect 18845 18405 18875 18410
rect 18925 18430 18955 18435
rect 18925 18410 18930 18430
rect 18930 18410 18950 18430
rect 18950 18410 18955 18430
rect 18925 18405 18955 18410
rect 19005 18430 19035 18435
rect 19005 18410 19010 18430
rect 19010 18410 19030 18430
rect 19030 18410 19035 18430
rect 19005 18405 19035 18410
rect 19085 18430 19115 18435
rect 19085 18410 19090 18430
rect 19090 18410 19110 18430
rect 19110 18410 19115 18430
rect 19085 18405 19115 18410
rect 19165 18430 19195 18435
rect 19165 18410 19170 18430
rect 19170 18410 19190 18430
rect 19190 18410 19195 18430
rect 19165 18405 19195 18410
rect 19245 18430 19275 18435
rect 19245 18410 19250 18430
rect 19250 18410 19270 18430
rect 19270 18410 19275 18430
rect 19245 18405 19275 18410
rect 19325 18430 19355 18435
rect 19325 18410 19330 18430
rect 19330 18410 19350 18430
rect 19350 18410 19355 18430
rect 19325 18405 19355 18410
rect 19405 18430 19435 18435
rect 19405 18410 19410 18430
rect 19410 18410 19430 18430
rect 19430 18410 19435 18430
rect 19405 18405 19435 18410
rect 19485 18430 19515 18435
rect 19485 18410 19490 18430
rect 19490 18410 19510 18430
rect 19510 18410 19515 18430
rect 19485 18405 19515 18410
rect 19565 18430 19595 18435
rect 19565 18410 19570 18430
rect 19570 18410 19590 18430
rect 19590 18410 19595 18430
rect 19565 18405 19595 18410
rect 19645 18430 19675 18435
rect 19645 18410 19650 18430
rect 19650 18410 19670 18430
rect 19670 18410 19675 18430
rect 19645 18405 19675 18410
rect 19725 18430 19755 18435
rect 19725 18410 19730 18430
rect 19730 18410 19750 18430
rect 19750 18410 19755 18430
rect 19725 18405 19755 18410
rect 19805 18430 19835 18435
rect 19805 18410 19810 18430
rect 19810 18410 19830 18430
rect 19830 18410 19835 18430
rect 19805 18405 19835 18410
rect 19885 18430 19915 18435
rect 19885 18410 19890 18430
rect 19890 18410 19910 18430
rect 19910 18410 19915 18430
rect 19885 18405 19915 18410
rect 19965 18430 19995 18435
rect 19965 18410 19970 18430
rect 19970 18410 19990 18430
rect 19990 18410 19995 18430
rect 19965 18405 19995 18410
rect 20045 18430 20075 18435
rect 20045 18410 20050 18430
rect 20050 18410 20070 18430
rect 20070 18410 20075 18430
rect 20045 18405 20075 18410
rect 20125 18430 20155 18435
rect 20125 18410 20130 18430
rect 20130 18410 20150 18430
rect 20150 18410 20155 18430
rect 20125 18405 20155 18410
rect 20205 18430 20235 18435
rect 20205 18410 20210 18430
rect 20210 18410 20230 18430
rect 20230 18410 20235 18430
rect 20205 18405 20235 18410
rect 20285 18430 20315 18435
rect 20285 18410 20290 18430
rect 20290 18410 20310 18430
rect 20310 18410 20315 18430
rect 20285 18405 20315 18410
rect 20365 18430 20395 18435
rect 20365 18410 20370 18430
rect 20370 18410 20390 18430
rect 20390 18410 20395 18430
rect 20365 18405 20395 18410
rect 20445 18430 20475 18435
rect 20445 18410 20450 18430
rect 20450 18410 20470 18430
rect 20470 18410 20475 18430
rect 20445 18405 20475 18410
rect 20525 18430 20555 18435
rect 20525 18410 20530 18430
rect 20530 18410 20550 18430
rect 20550 18410 20555 18430
rect 20525 18405 20555 18410
rect 20605 18430 20635 18435
rect 20605 18410 20610 18430
rect 20610 18410 20630 18430
rect 20630 18410 20635 18430
rect 20605 18405 20635 18410
rect 20685 18430 20715 18435
rect 20685 18410 20690 18430
rect 20690 18410 20710 18430
rect 20710 18410 20715 18430
rect 20685 18405 20715 18410
rect 20765 18430 20795 18435
rect 20765 18410 20770 18430
rect 20770 18410 20790 18430
rect 20790 18410 20795 18430
rect 20765 18405 20795 18410
rect 20845 18430 20875 18435
rect 20845 18410 20850 18430
rect 20850 18410 20870 18430
rect 20870 18410 20875 18430
rect 20845 18405 20875 18410
rect 20925 18430 20955 18435
rect 20925 18410 20930 18430
rect 20930 18410 20950 18430
rect 20950 18410 20955 18430
rect 20925 18405 20955 18410
rect 5 18270 35 18275
rect 5 18250 10 18270
rect 10 18250 30 18270
rect 30 18250 35 18270
rect 5 18245 35 18250
rect 85 18270 115 18275
rect 85 18250 90 18270
rect 90 18250 110 18270
rect 110 18250 115 18270
rect 85 18245 115 18250
rect 165 18270 195 18275
rect 165 18250 170 18270
rect 170 18250 190 18270
rect 190 18250 195 18270
rect 165 18245 195 18250
rect 245 18270 275 18275
rect 245 18250 250 18270
rect 250 18250 270 18270
rect 270 18250 275 18270
rect 245 18245 275 18250
rect 325 18270 355 18275
rect 325 18250 330 18270
rect 330 18250 350 18270
rect 350 18250 355 18270
rect 325 18245 355 18250
rect 405 18270 435 18275
rect 405 18250 410 18270
rect 410 18250 430 18270
rect 430 18250 435 18270
rect 405 18245 435 18250
rect 485 18270 515 18275
rect 485 18250 490 18270
rect 490 18250 510 18270
rect 510 18250 515 18270
rect 485 18245 515 18250
rect 565 18270 595 18275
rect 565 18250 570 18270
rect 570 18250 590 18270
rect 590 18250 595 18270
rect 565 18245 595 18250
rect 645 18270 675 18275
rect 645 18250 650 18270
rect 650 18250 670 18270
rect 670 18250 675 18270
rect 645 18245 675 18250
rect 725 18270 755 18275
rect 725 18250 730 18270
rect 730 18250 750 18270
rect 750 18250 755 18270
rect 725 18245 755 18250
rect 805 18270 835 18275
rect 805 18250 810 18270
rect 810 18250 830 18270
rect 830 18250 835 18270
rect 805 18245 835 18250
rect 885 18270 915 18275
rect 885 18250 890 18270
rect 890 18250 910 18270
rect 910 18250 915 18270
rect 885 18245 915 18250
rect 965 18270 995 18275
rect 965 18250 970 18270
rect 970 18250 990 18270
rect 990 18250 995 18270
rect 965 18245 995 18250
rect 1045 18270 1075 18275
rect 1045 18250 1050 18270
rect 1050 18250 1070 18270
rect 1070 18250 1075 18270
rect 1045 18245 1075 18250
rect 1125 18270 1155 18275
rect 1125 18250 1130 18270
rect 1130 18250 1150 18270
rect 1150 18250 1155 18270
rect 1125 18245 1155 18250
rect 1205 18270 1235 18275
rect 1205 18250 1210 18270
rect 1210 18250 1230 18270
rect 1230 18250 1235 18270
rect 1205 18245 1235 18250
rect 1285 18270 1315 18275
rect 1285 18250 1290 18270
rect 1290 18250 1310 18270
rect 1310 18250 1315 18270
rect 1285 18245 1315 18250
rect 1365 18270 1395 18275
rect 1365 18250 1370 18270
rect 1370 18250 1390 18270
rect 1390 18250 1395 18270
rect 1365 18245 1395 18250
rect 1445 18270 1475 18275
rect 1445 18250 1450 18270
rect 1450 18250 1470 18270
rect 1470 18250 1475 18270
rect 1445 18245 1475 18250
rect 1525 18270 1555 18275
rect 1525 18250 1530 18270
rect 1530 18250 1550 18270
rect 1550 18250 1555 18270
rect 1525 18245 1555 18250
rect 1605 18270 1635 18275
rect 1605 18250 1610 18270
rect 1610 18250 1630 18270
rect 1630 18250 1635 18270
rect 1605 18245 1635 18250
rect 1685 18270 1715 18275
rect 1685 18250 1690 18270
rect 1690 18250 1710 18270
rect 1710 18250 1715 18270
rect 1685 18245 1715 18250
rect 1765 18270 1795 18275
rect 1765 18250 1770 18270
rect 1770 18250 1790 18270
rect 1790 18250 1795 18270
rect 1765 18245 1795 18250
rect 1845 18270 1875 18275
rect 1845 18250 1850 18270
rect 1850 18250 1870 18270
rect 1870 18250 1875 18270
rect 1845 18245 1875 18250
rect 1925 18270 1955 18275
rect 1925 18250 1930 18270
rect 1930 18250 1950 18270
rect 1950 18250 1955 18270
rect 1925 18245 1955 18250
rect 2005 18270 2035 18275
rect 2005 18250 2010 18270
rect 2010 18250 2030 18270
rect 2030 18250 2035 18270
rect 2005 18245 2035 18250
rect 2085 18270 2115 18275
rect 2085 18250 2090 18270
rect 2090 18250 2110 18270
rect 2110 18250 2115 18270
rect 2085 18245 2115 18250
rect 2165 18270 2195 18275
rect 2165 18250 2170 18270
rect 2170 18250 2190 18270
rect 2190 18250 2195 18270
rect 2165 18245 2195 18250
rect 2245 18270 2275 18275
rect 2245 18250 2250 18270
rect 2250 18250 2270 18270
rect 2270 18250 2275 18270
rect 2245 18245 2275 18250
rect 2325 18270 2355 18275
rect 2325 18250 2330 18270
rect 2330 18250 2350 18270
rect 2350 18250 2355 18270
rect 2325 18245 2355 18250
rect 2405 18270 2435 18275
rect 2405 18250 2410 18270
rect 2410 18250 2430 18270
rect 2430 18250 2435 18270
rect 2405 18245 2435 18250
rect 2485 18270 2515 18275
rect 2485 18250 2490 18270
rect 2490 18250 2510 18270
rect 2510 18250 2515 18270
rect 2485 18245 2515 18250
rect 2565 18270 2595 18275
rect 2565 18250 2570 18270
rect 2570 18250 2590 18270
rect 2590 18250 2595 18270
rect 2565 18245 2595 18250
rect 2645 18270 2675 18275
rect 2645 18250 2650 18270
rect 2650 18250 2670 18270
rect 2670 18250 2675 18270
rect 2645 18245 2675 18250
rect 2725 18270 2755 18275
rect 2725 18250 2730 18270
rect 2730 18250 2750 18270
rect 2750 18250 2755 18270
rect 2725 18245 2755 18250
rect 2805 18270 2835 18275
rect 2805 18250 2810 18270
rect 2810 18250 2830 18270
rect 2830 18250 2835 18270
rect 2805 18245 2835 18250
rect 2885 18270 2915 18275
rect 2885 18250 2890 18270
rect 2890 18250 2910 18270
rect 2910 18250 2915 18270
rect 2885 18245 2915 18250
rect 2965 18270 2995 18275
rect 2965 18250 2970 18270
rect 2970 18250 2990 18270
rect 2990 18250 2995 18270
rect 2965 18245 2995 18250
rect 3045 18270 3075 18275
rect 3045 18250 3050 18270
rect 3050 18250 3070 18270
rect 3070 18250 3075 18270
rect 3045 18245 3075 18250
rect 3125 18270 3155 18275
rect 3125 18250 3130 18270
rect 3130 18250 3150 18270
rect 3150 18250 3155 18270
rect 3125 18245 3155 18250
rect 3205 18270 3235 18275
rect 3205 18250 3210 18270
rect 3210 18250 3230 18270
rect 3230 18250 3235 18270
rect 3205 18245 3235 18250
rect 3285 18270 3315 18275
rect 3285 18250 3290 18270
rect 3290 18250 3310 18270
rect 3310 18250 3315 18270
rect 3285 18245 3315 18250
rect 3365 18270 3395 18275
rect 3365 18250 3370 18270
rect 3370 18250 3390 18270
rect 3390 18250 3395 18270
rect 3365 18245 3395 18250
rect 3445 18270 3475 18275
rect 3445 18250 3450 18270
rect 3450 18250 3470 18270
rect 3470 18250 3475 18270
rect 3445 18245 3475 18250
rect 3525 18270 3555 18275
rect 3525 18250 3530 18270
rect 3530 18250 3550 18270
rect 3550 18250 3555 18270
rect 3525 18245 3555 18250
rect 3605 18270 3635 18275
rect 3605 18250 3610 18270
rect 3610 18250 3630 18270
rect 3630 18250 3635 18270
rect 3605 18245 3635 18250
rect 3685 18270 3715 18275
rect 3685 18250 3690 18270
rect 3690 18250 3710 18270
rect 3710 18250 3715 18270
rect 3685 18245 3715 18250
rect 3765 18270 3795 18275
rect 3765 18250 3770 18270
rect 3770 18250 3790 18270
rect 3790 18250 3795 18270
rect 3765 18245 3795 18250
rect 3845 18270 3875 18275
rect 3845 18250 3850 18270
rect 3850 18250 3870 18270
rect 3870 18250 3875 18270
rect 3845 18245 3875 18250
rect 3925 18270 3955 18275
rect 3925 18250 3930 18270
rect 3930 18250 3950 18270
rect 3950 18250 3955 18270
rect 3925 18245 3955 18250
rect 4005 18270 4035 18275
rect 4005 18250 4010 18270
rect 4010 18250 4030 18270
rect 4030 18250 4035 18270
rect 4005 18245 4035 18250
rect 4085 18270 4115 18275
rect 4085 18250 4090 18270
rect 4090 18250 4110 18270
rect 4110 18250 4115 18270
rect 4085 18245 4115 18250
rect 4165 18270 4195 18275
rect 4165 18250 4170 18270
rect 4170 18250 4190 18270
rect 4190 18250 4195 18270
rect 4165 18245 4195 18250
rect 6245 18270 6275 18275
rect 6245 18250 6250 18270
rect 6250 18250 6270 18270
rect 6270 18250 6275 18270
rect 6245 18245 6275 18250
rect 6325 18270 6355 18275
rect 6325 18250 6330 18270
rect 6330 18250 6350 18270
rect 6350 18250 6355 18270
rect 6325 18245 6355 18250
rect 6405 18270 6435 18275
rect 6405 18250 6410 18270
rect 6410 18250 6430 18270
rect 6430 18250 6435 18270
rect 6405 18245 6435 18250
rect 6485 18270 6515 18275
rect 6485 18250 6490 18270
rect 6490 18250 6510 18270
rect 6510 18250 6515 18270
rect 6485 18245 6515 18250
rect 6565 18270 6595 18275
rect 6565 18250 6570 18270
rect 6570 18250 6590 18270
rect 6590 18250 6595 18270
rect 6565 18245 6595 18250
rect 6645 18270 6675 18275
rect 6645 18250 6650 18270
rect 6650 18250 6670 18270
rect 6670 18250 6675 18270
rect 6645 18245 6675 18250
rect 6725 18270 6755 18275
rect 6725 18250 6730 18270
rect 6730 18250 6750 18270
rect 6750 18250 6755 18270
rect 6725 18245 6755 18250
rect 6805 18270 6835 18275
rect 6805 18250 6810 18270
rect 6810 18250 6830 18270
rect 6830 18250 6835 18270
rect 6805 18245 6835 18250
rect 6885 18270 6915 18275
rect 6885 18250 6890 18270
rect 6890 18250 6910 18270
rect 6910 18250 6915 18270
rect 6885 18245 6915 18250
rect 6965 18270 6995 18275
rect 6965 18250 6970 18270
rect 6970 18250 6990 18270
rect 6990 18250 6995 18270
rect 6965 18245 6995 18250
rect 7045 18270 7075 18275
rect 7045 18250 7050 18270
rect 7050 18250 7070 18270
rect 7070 18250 7075 18270
rect 7045 18245 7075 18250
rect 7125 18270 7155 18275
rect 7125 18250 7130 18270
rect 7130 18250 7150 18270
rect 7150 18250 7155 18270
rect 7125 18245 7155 18250
rect 7205 18270 7235 18275
rect 7205 18250 7210 18270
rect 7210 18250 7230 18270
rect 7230 18250 7235 18270
rect 7205 18245 7235 18250
rect 7285 18270 7315 18275
rect 7285 18250 7290 18270
rect 7290 18250 7310 18270
rect 7310 18250 7315 18270
rect 7285 18245 7315 18250
rect 7365 18270 7395 18275
rect 7365 18250 7370 18270
rect 7370 18250 7390 18270
rect 7390 18250 7395 18270
rect 7365 18245 7395 18250
rect 7445 18270 7475 18275
rect 7445 18250 7450 18270
rect 7450 18250 7470 18270
rect 7470 18250 7475 18270
rect 7445 18245 7475 18250
rect 7525 18270 7555 18275
rect 7525 18250 7530 18270
rect 7530 18250 7550 18270
rect 7550 18250 7555 18270
rect 7525 18245 7555 18250
rect 7605 18270 7635 18275
rect 7605 18250 7610 18270
rect 7610 18250 7630 18270
rect 7630 18250 7635 18270
rect 7605 18245 7635 18250
rect 7685 18270 7715 18275
rect 7685 18250 7690 18270
rect 7690 18250 7710 18270
rect 7710 18250 7715 18270
rect 7685 18245 7715 18250
rect 7765 18270 7795 18275
rect 7765 18250 7770 18270
rect 7770 18250 7790 18270
rect 7790 18250 7795 18270
rect 7765 18245 7795 18250
rect 7845 18270 7875 18275
rect 7845 18250 7850 18270
rect 7850 18250 7870 18270
rect 7870 18250 7875 18270
rect 7845 18245 7875 18250
rect 7925 18270 7955 18275
rect 7925 18250 7930 18270
rect 7930 18250 7950 18270
rect 7950 18250 7955 18270
rect 7925 18245 7955 18250
rect 8005 18270 8035 18275
rect 8005 18250 8010 18270
rect 8010 18250 8030 18270
rect 8030 18250 8035 18270
rect 8005 18245 8035 18250
rect 8085 18270 8115 18275
rect 8085 18250 8090 18270
rect 8090 18250 8110 18270
rect 8110 18250 8115 18270
rect 8085 18245 8115 18250
rect 8165 18270 8195 18275
rect 8165 18250 8170 18270
rect 8170 18250 8190 18270
rect 8190 18250 8195 18270
rect 8165 18245 8195 18250
rect 8245 18270 8275 18275
rect 8245 18250 8250 18270
rect 8250 18250 8270 18270
rect 8270 18250 8275 18270
rect 8245 18245 8275 18250
rect 8325 18270 8355 18275
rect 8325 18250 8330 18270
rect 8330 18250 8350 18270
rect 8350 18250 8355 18270
rect 8325 18245 8355 18250
rect 8405 18270 8435 18275
rect 8405 18250 8410 18270
rect 8410 18250 8430 18270
rect 8430 18250 8435 18270
rect 8405 18245 8435 18250
rect 8485 18270 8515 18275
rect 8485 18250 8490 18270
rect 8490 18250 8510 18270
rect 8510 18250 8515 18270
rect 8485 18245 8515 18250
rect 8565 18270 8595 18275
rect 8565 18250 8570 18270
rect 8570 18250 8590 18270
rect 8590 18250 8595 18270
rect 8565 18245 8595 18250
rect 8645 18270 8675 18275
rect 8645 18250 8650 18270
rect 8650 18250 8670 18270
rect 8670 18250 8675 18270
rect 8645 18245 8675 18250
rect 8725 18270 8755 18275
rect 8725 18250 8730 18270
rect 8730 18250 8750 18270
rect 8750 18250 8755 18270
rect 8725 18245 8755 18250
rect 8805 18270 8835 18275
rect 8805 18250 8810 18270
rect 8810 18250 8830 18270
rect 8830 18250 8835 18270
rect 8805 18245 8835 18250
rect 8885 18270 8915 18275
rect 8885 18250 8890 18270
rect 8890 18250 8910 18270
rect 8910 18250 8915 18270
rect 8885 18245 8915 18250
rect 8965 18270 8995 18275
rect 8965 18250 8970 18270
rect 8970 18250 8990 18270
rect 8990 18250 8995 18270
rect 8965 18245 8995 18250
rect 9045 18270 9075 18275
rect 9045 18250 9050 18270
rect 9050 18250 9070 18270
rect 9070 18250 9075 18270
rect 9045 18245 9075 18250
rect 9125 18270 9155 18275
rect 9125 18250 9130 18270
rect 9130 18250 9150 18270
rect 9150 18250 9155 18270
rect 9125 18245 9155 18250
rect 9205 18270 9235 18275
rect 9205 18250 9210 18270
rect 9210 18250 9230 18270
rect 9230 18250 9235 18270
rect 9205 18245 9235 18250
rect 9285 18270 9315 18275
rect 9285 18250 9290 18270
rect 9290 18250 9310 18270
rect 9310 18250 9315 18270
rect 9285 18245 9315 18250
rect 9365 18270 9395 18275
rect 9365 18250 9370 18270
rect 9370 18250 9390 18270
rect 9390 18250 9395 18270
rect 9365 18245 9395 18250
rect 9445 18270 9475 18275
rect 9445 18250 9450 18270
rect 9450 18250 9470 18270
rect 9470 18250 9475 18270
rect 9445 18245 9475 18250
rect 11565 18270 11595 18275
rect 11565 18250 11570 18270
rect 11570 18250 11590 18270
rect 11590 18250 11595 18270
rect 11565 18245 11595 18250
rect 11645 18270 11675 18275
rect 11645 18250 11650 18270
rect 11650 18250 11670 18270
rect 11670 18250 11675 18270
rect 11645 18245 11675 18250
rect 11725 18270 11755 18275
rect 11725 18250 11730 18270
rect 11730 18250 11750 18270
rect 11750 18250 11755 18270
rect 11725 18245 11755 18250
rect 11805 18270 11835 18275
rect 11805 18250 11810 18270
rect 11810 18250 11830 18270
rect 11830 18250 11835 18270
rect 11805 18245 11835 18250
rect 11885 18270 11915 18275
rect 11885 18250 11890 18270
rect 11890 18250 11910 18270
rect 11910 18250 11915 18270
rect 11885 18245 11915 18250
rect 11965 18270 11995 18275
rect 11965 18250 11970 18270
rect 11970 18250 11990 18270
rect 11990 18250 11995 18270
rect 11965 18245 11995 18250
rect 12045 18270 12075 18275
rect 12045 18250 12050 18270
rect 12050 18250 12070 18270
rect 12070 18250 12075 18270
rect 12045 18245 12075 18250
rect 12125 18270 12155 18275
rect 12125 18250 12130 18270
rect 12130 18250 12150 18270
rect 12150 18250 12155 18270
rect 12125 18245 12155 18250
rect 12205 18270 12235 18275
rect 12205 18250 12210 18270
rect 12210 18250 12230 18270
rect 12230 18250 12235 18270
rect 12205 18245 12235 18250
rect 12285 18270 12315 18275
rect 12285 18250 12290 18270
rect 12290 18250 12310 18270
rect 12310 18250 12315 18270
rect 12285 18245 12315 18250
rect 12365 18270 12395 18275
rect 12365 18250 12370 18270
rect 12370 18250 12390 18270
rect 12390 18250 12395 18270
rect 12365 18245 12395 18250
rect 12445 18270 12475 18275
rect 12445 18250 12450 18270
rect 12450 18250 12470 18270
rect 12470 18250 12475 18270
rect 12445 18245 12475 18250
rect 12525 18270 12555 18275
rect 12525 18250 12530 18270
rect 12530 18250 12550 18270
rect 12550 18250 12555 18270
rect 12525 18245 12555 18250
rect 12605 18270 12635 18275
rect 12605 18250 12610 18270
rect 12610 18250 12630 18270
rect 12630 18250 12635 18270
rect 12605 18245 12635 18250
rect 12685 18270 12715 18275
rect 12685 18250 12690 18270
rect 12690 18250 12710 18270
rect 12710 18250 12715 18270
rect 12685 18245 12715 18250
rect 12765 18270 12795 18275
rect 12765 18250 12770 18270
rect 12770 18250 12790 18270
rect 12790 18250 12795 18270
rect 12765 18245 12795 18250
rect 12845 18270 12875 18275
rect 12845 18250 12850 18270
rect 12850 18250 12870 18270
rect 12870 18250 12875 18270
rect 12845 18245 12875 18250
rect 12925 18270 12955 18275
rect 12925 18250 12930 18270
rect 12930 18250 12950 18270
rect 12950 18250 12955 18270
rect 12925 18245 12955 18250
rect 13005 18270 13035 18275
rect 13005 18250 13010 18270
rect 13010 18250 13030 18270
rect 13030 18250 13035 18270
rect 13005 18245 13035 18250
rect 13085 18270 13115 18275
rect 13085 18250 13090 18270
rect 13090 18250 13110 18270
rect 13110 18250 13115 18270
rect 13085 18245 13115 18250
rect 13165 18270 13195 18275
rect 13165 18250 13170 18270
rect 13170 18250 13190 18270
rect 13190 18250 13195 18270
rect 13165 18245 13195 18250
rect 13245 18270 13275 18275
rect 13245 18250 13250 18270
rect 13250 18250 13270 18270
rect 13270 18250 13275 18270
rect 13245 18245 13275 18250
rect 13325 18270 13355 18275
rect 13325 18250 13330 18270
rect 13330 18250 13350 18270
rect 13350 18250 13355 18270
rect 13325 18245 13355 18250
rect 13405 18270 13435 18275
rect 13405 18250 13410 18270
rect 13410 18250 13430 18270
rect 13430 18250 13435 18270
rect 13405 18245 13435 18250
rect 13485 18270 13515 18275
rect 13485 18250 13490 18270
rect 13490 18250 13510 18270
rect 13510 18250 13515 18270
rect 13485 18245 13515 18250
rect 13565 18270 13595 18275
rect 13565 18250 13570 18270
rect 13570 18250 13590 18270
rect 13590 18250 13595 18270
rect 13565 18245 13595 18250
rect 13645 18270 13675 18275
rect 13645 18250 13650 18270
rect 13650 18250 13670 18270
rect 13670 18250 13675 18270
rect 13645 18245 13675 18250
rect 13725 18270 13755 18275
rect 13725 18250 13730 18270
rect 13730 18250 13750 18270
rect 13750 18250 13755 18270
rect 13725 18245 13755 18250
rect 13805 18270 13835 18275
rect 13805 18250 13810 18270
rect 13810 18250 13830 18270
rect 13830 18250 13835 18270
rect 13805 18245 13835 18250
rect 13885 18270 13915 18275
rect 13885 18250 13890 18270
rect 13890 18250 13910 18270
rect 13910 18250 13915 18270
rect 13885 18245 13915 18250
rect 13965 18270 13995 18275
rect 13965 18250 13970 18270
rect 13970 18250 13990 18270
rect 13990 18250 13995 18270
rect 13965 18245 13995 18250
rect 14045 18270 14075 18275
rect 14045 18250 14050 18270
rect 14050 18250 14070 18270
rect 14070 18250 14075 18270
rect 14045 18245 14075 18250
rect 14125 18270 14155 18275
rect 14125 18250 14130 18270
rect 14130 18250 14150 18270
rect 14150 18250 14155 18270
rect 14125 18245 14155 18250
rect 14205 18270 14235 18275
rect 14205 18250 14210 18270
rect 14210 18250 14230 18270
rect 14230 18250 14235 18270
rect 14205 18245 14235 18250
rect 14285 18270 14315 18275
rect 14285 18250 14290 18270
rect 14290 18250 14310 18270
rect 14310 18250 14315 18270
rect 14285 18245 14315 18250
rect 14365 18270 14395 18275
rect 14365 18250 14370 18270
rect 14370 18250 14390 18270
rect 14390 18250 14395 18270
rect 14365 18245 14395 18250
rect 14445 18270 14475 18275
rect 14445 18250 14450 18270
rect 14450 18250 14470 18270
rect 14470 18250 14475 18270
rect 14445 18245 14475 18250
rect 14525 18270 14555 18275
rect 14525 18250 14530 18270
rect 14530 18250 14550 18270
rect 14550 18250 14555 18270
rect 14525 18245 14555 18250
rect 14605 18270 14635 18275
rect 14605 18250 14610 18270
rect 14610 18250 14630 18270
rect 14630 18250 14635 18270
rect 14605 18245 14635 18250
rect 14685 18270 14715 18275
rect 14685 18250 14690 18270
rect 14690 18250 14710 18270
rect 14710 18250 14715 18270
rect 14685 18245 14715 18250
rect 16765 18270 16795 18275
rect 16765 18250 16770 18270
rect 16770 18250 16790 18270
rect 16790 18250 16795 18270
rect 16765 18245 16795 18250
rect 16845 18270 16875 18275
rect 16845 18250 16850 18270
rect 16850 18250 16870 18270
rect 16870 18250 16875 18270
rect 16845 18245 16875 18250
rect 16925 18270 16955 18275
rect 16925 18250 16930 18270
rect 16930 18250 16950 18270
rect 16950 18250 16955 18270
rect 16925 18245 16955 18250
rect 17005 18270 17035 18275
rect 17005 18250 17010 18270
rect 17010 18250 17030 18270
rect 17030 18250 17035 18270
rect 17005 18245 17035 18250
rect 17085 18270 17115 18275
rect 17085 18250 17090 18270
rect 17090 18250 17110 18270
rect 17110 18250 17115 18270
rect 17085 18245 17115 18250
rect 17165 18270 17195 18275
rect 17165 18250 17170 18270
rect 17170 18250 17190 18270
rect 17190 18250 17195 18270
rect 17165 18245 17195 18250
rect 17245 18270 17275 18275
rect 17245 18250 17250 18270
rect 17250 18250 17270 18270
rect 17270 18250 17275 18270
rect 17245 18245 17275 18250
rect 17325 18270 17355 18275
rect 17325 18250 17330 18270
rect 17330 18250 17350 18270
rect 17350 18250 17355 18270
rect 17325 18245 17355 18250
rect 17405 18270 17435 18275
rect 17405 18250 17410 18270
rect 17410 18250 17430 18270
rect 17430 18250 17435 18270
rect 17405 18245 17435 18250
rect 17485 18270 17515 18275
rect 17485 18250 17490 18270
rect 17490 18250 17510 18270
rect 17510 18250 17515 18270
rect 17485 18245 17515 18250
rect 17565 18270 17595 18275
rect 17565 18250 17570 18270
rect 17570 18250 17590 18270
rect 17590 18250 17595 18270
rect 17565 18245 17595 18250
rect 17645 18270 17675 18275
rect 17645 18250 17650 18270
rect 17650 18250 17670 18270
rect 17670 18250 17675 18270
rect 17645 18245 17675 18250
rect 17725 18270 17755 18275
rect 17725 18250 17730 18270
rect 17730 18250 17750 18270
rect 17750 18250 17755 18270
rect 17725 18245 17755 18250
rect 17805 18270 17835 18275
rect 17805 18250 17810 18270
rect 17810 18250 17830 18270
rect 17830 18250 17835 18270
rect 17805 18245 17835 18250
rect 17885 18270 17915 18275
rect 17885 18250 17890 18270
rect 17890 18250 17910 18270
rect 17910 18250 17915 18270
rect 17885 18245 17915 18250
rect 17965 18270 17995 18275
rect 17965 18250 17970 18270
rect 17970 18250 17990 18270
rect 17990 18250 17995 18270
rect 17965 18245 17995 18250
rect 18045 18270 18075 18275
rect 18045 18250 18050 18270
rect 18050 18250 18070 18270
rect 18070 18250 18075 18270
rect 18045 18245 18075 18250
rect 18125 18270 18155 18275
rect 18125 18250 18130 18270
rect 18130 18250 18150 18270
rect 18150 18250 18155 18270
rect 18125 18245 18155 18250
rect 18205 18270 18235 18275
rect 18205 18250 18210 18270
rect 18210 18250 18230 18270
rect 18230 18250 18235 18270
rect 18205 18245 18235 18250
rect 18285 18270 18315 18275
rect 18285 18250 18290 18270
rect 18290 18250 18310 18270
rect 18310 18250 18315 18270
rect 18285 18245 18315 18250
rect 18365 18270 18395 18275
rect 18365 18250 18370 18270
rect 18370 18250 18390 18270
rect 18390 18250 18395 18270
rect 18365 18245 18395 18250
rect 18445 18270 18475 18275
rect 18445 18250 18450 18270
rect 18450 18250 18470 18270
rect 18470 18250 18475 18270
rect 18445 18245 18475 18250
rect 18525 18270 18555 18275
rect 18525 18250 18530 18270
rect 18530 18250 18550 18270
rect 18550 18250 18555 18270
rect 18525 18245 18555 18250
rect 18605 18270 18635 18275
rect 18605 18250 18610 18270
rect 18610 18250 18630 18270
rect 18630 18250 18635 18270
rect 18605 18245 18635 18250
rect 18685 18270 18715 18275
rect 18685 18250 18690 18270
rect 18690 18250 18710 18270
rect 18710 18250 18715 18270
rect 18685 18245 18715 18250
rect 18765 18270 18795 18275
rect 18765 18250 18770 18270
rect 18770 18250 18790 18270
rect 18790 18250 18795 18270
rect 18765 18245 18795 18250
rect 18845 18270 18875 18275
rect 18845 18250 18850 18270
rect 18850 18250 18870 18270
rect 18870 18250 18875 18270
rect 18845 18245 18875 18250
rect 18925 18270 18955 18275
rect 18925 18250 18930 18270
rect 18930 18250 18950 18270
rect 18950 18250 18955 18270
rect 18925 18245 18955 18250
rect 19005 18270 19035 18275
rect 19005 18250 19010 18270
rect 19010 18250 19030 18270
rect 19030 18250 19035 18270
rect 19005 18245 19035 18250
rect 19085 18270 19115 18275
rect 19085 18250 19090 18270
rect 19090 18250 19110 18270
rect 19110 18250 19115 18270
rect 19085 18245 19115 18250
rect 19165 18270 19195 18275
rect 19165 18250 19170 18270
rect 19170 18250 19190 18270
rect 19190 18250 19195 18270
rect 19165 18245 19195 18250
rect 19245 18270 19275 18275
rect 19245 18250 19250 18270
rect 19250 18250 19270 18270
rect 19270 18250 19275 18270
rect 19245 18245 19275 18250
rect 19325 18270 19355 18275
rect 19325 18250 19330 18270
rect 19330 18250 19350 18270
rect 19350 18250 19355 18270
rect 19325 18245 19355 18250
rect 19405 18270 19435 18275
rect 19405 18250 19410 18270
rect 19410 18250 19430 18270
rect 19430 18250 19435 18270
rect 19405 18245 19435 18250
rect 19485 18270 19515 18275
rect 19485 18250 19490 18270
rect 19490 18250 19510 18270
rect 19510 18250 19515 18270
rect 19485 18245 19515 18250
rect 19565 18270 19595 18275
rect 19565 18250 19570 18270
rect 19570 18250 19590 18270
rect 19590 18250 19595 18270
rect 19565 18245 19595 18250
rect 19645 18270 19675 18275
rect 19645 18250 19650 18270
rect 19650 18250 19670 18270
rect 19670 18250 19675 18270
rect 19645 18245 19675 18250
rect 19725 18270 19755 18275
rect 19725 18250 19730 18270
rect 19730 18250 19750 18270
rect 19750 18250 19755 18270
rect 19725 18245 19755 18250
rect 19805 18270 19835 18275
rect 19805 18250 19810 18270
rect 19810 18250 19830 18270
rect 19830 18250 19835 18270
rect 19805 18245 19835 18250
rect 19885 18270 19915 18275
rect 19885 18250 19890 18270
rect 19890 18250 19910 18270
rect 19910 18250 19915 18270
rect 19885 18245 19915 18250
rect 19965 18270 19995 18275
rect 19965 18250 19970 18270
rect 19970 18250 19990 18270
rect 19990 18250 19995 18270
rect 19965 18245 19995 18250
rect 20045 18270 20075 18275
rect 20045 18250 20050 18270
rect 20050 18250 20070 18270
rect 20070 18250 20075 18270
rect 20045 18245 20075 18250
rect 20125 18270 20155 18275
rect 20125 18250 20130 18270
rect 20130 18250 20150 18270
rect 20150 18250 20155 18270
rect 20125 18245 20155 18250
rect 20205 18270 20235 18275
rect 20205 18250 20210 18270
rect 20210 18250 20230 18270
rect 20230 18250 20235 18270
rect 20205 18245 20235 18250
rect 20285 18270 20315 18275
rect 20285 18250 20290 18270
rect 20290 18250 20310 18270
rect 20310 18250 20315 18270
rect 20285 18245 20315 18250
rect 20365 18270 20395 18275
rect 20365 18250 20370 18270
rect 20370 18250 20390 18270
rect 20390 18250 20395 18270
rect 20365 18245 20395 18250
rect 20445 18270 20475 18275
rect 20445 18250 20450 18270
rect 20450 18250 20470 18270
rect 20470 18250 20475 18270
rect 20445 18245 20475 18250
rect 20525 18270 20555 18275
rect 20525 18250 20530 18270
rect 20530 18250 20550 18270
rect 20550 18250 20555 18270
rect 20525 18245 20555 18250
rect 20605 18270 20635 18275
rect 20605 18250 20610 18270
rect 20610 18250 20630 18270
rect 20630 18250 20635 18270
rect 20605 18245 20635 18250
rect 20685 18270 20715 18275
rect 20685 18250 20690 18270
rect 20690 18250 20710 18270
rect 20710 18250 20715 18270
rect 20685 18245 20715 18250
rect 20765 18270 20795 18275
rect 20765 18250 20770 18270
rect 20770 18250 20790 18270
rect 20790 18250 20795 18270
rect 20765 18245 20795 18250
rect 20845 18270 20875 18275
rect 20845 18250 20850 18270
rect 20850 18250 20870 18270
rect 20870 18250 20875 18270
rect 20845 18245 20875 18250
rect 20925 18270 20955 18275
rect 20925 18250 20930 18270
rect 20930 18250 20950 18270
rect 20950 18250 20955 18270
rect 20925 18245 20955 18250
rect 5 18190 35 18195
rect 5 18170 10 18190
rect 10 18170 30 18190
rect 30 18170 35 18190
rect 5 18165 35 18170
rect 85 18190 115 18195
rect 85 18170 90 18190
rect 90 18170 110 18190
rect 110 18170 115 18190
rect 85 18165 115 18170
rect 165 18190 195 18195
rect 165 18170 170 18190
rect 170 18170 190 18190
rect 190 18170 195 18190
rect 165 18165 195 18170
rect 245 18190 275 18195
rect 245 18170 250 18190
rect 250 18170 270 18190
rect 270 18170 275 18190
rect 245 18165 275 18170
rect 325 18190 355 18195
rect 325 18170 330 18190
rect 330 18170 350 18190
rect 350 18170 355 18190
rect 325 18165 355 18170
rect 405 18190 435 18195
rect 405 18170 410 18190
rect 410 18170 430 18190
rect 430 18170 435 18190
rect 405 18165 435 18170
rect 485 18190 515 18195
rect 485 18170 490 18190
rect 490 18170 510 18190
rect 510 18170 515 18190
rect 485 18165 515 18170
rect 565 18190 595 18195
rect 565 18170 570 18190
rect 570 18170 590 18190
rect 590 18170 595 18190
rect 565 18165 595 18170
rect 645 18190 675 18195
rect 645 18170 650 18190
rect 650 18170 670 18190
rect 670 18170 675 18190
rect 645 18165 675 18170
rect 725 18190 755 18195
rect 725 18170 730 18190
rect 730 18170 750 18190
rect 750 18170 755 18190
rect 725 18165 755 18170
rect 805 18190 835 18195
rect 805 18170 810 18190
rect 810 18170 830 18190
rect 830 18170 835 18190
rect 805 18165 835 18170
rect 885 18190 915 18195
rect 885 18170 890 18190
rect 890 18170 910 18190
rect 910 18170 915 18190
rect 885 18165 915 18170
rect 965 18190 995 18195
rect 965 18170 970 18190
rect 970 18170 990 18190
rect 990 18170 995 18190
rect 965 18165 995 18170
rect 1045 18190 1075 18195
rect 1045 18170 1050 18190
rect 1050 18170 1070 18190
rect 1070 18170 1075 18190
rect 1045 18165 1075 18170
rect 1125 18190 1155 18195
rect 1125 18170 1130 18190
rect 1130 18170 1150 18190
rect 1150 18170 1155 18190
rect 1125 18165 1155 18170
rect 1205 18190 1235 18195
rect 1205 18170 1210 18190
rect 1210 18170 1230 18190
rect 1230 18170 1235 18190
rect 1205 18165 1235 18170
rect 1285 18190 1315 18195
rect 1285 18170 1290 18190
rect 1290 18170 1310 18190
rect 1310 18170 1315 18190
rect 1285 18165 1315 18170
rect 1365 18190 1395 18195
rect 1365 18170 1370 18190
rect 1370 18170 1390 18190
rect 1390 18170 1395 18190
rect 1365 18165 1395 18170
rect 1445 18190 1475 18195
rect 1445 18170 1450 18190
rect 1450 18170 1470 18190
rect 1470 18170 1475 18190
rect 1445 18165 1475 18170
rect 1525 18190 1555 18195
rect 1525 18170 1530 18190
rect 1530 18170 1550 18190
rect 1550 18170 1555 18190
rect 1525 18165 1555 18170
rect 1605 18190 1635 18195
rect 1605 18170 1610 18190
rect 1610 18170 1630 18190
rect 1630 18170 1635 18190
rect 1605 18165 1635 18170
rect 1685 18190 1715 18195
rect 1685 18170 1690 18190
rect 1690 18170 1710 18190
rect 1710 18170 1715 18190
rect 1685 18165 1715 18170
rect 1765 18190 1795 18195
rect 1765 18170 1770 18190
rect 1770 18170 1790 18190
rect 1790 18170 1795 18190
rect 1765 18165 1795 18170
rect 1845 18190 1875 18195
rect 1845 18170 1850 18190
rect 1850 18170 1870 18190
rect 1870 18170 1875 18190
rect 1845 18165 1875 18170
rect 1925 18190 1955 18195
rect 1925 18170 1930 18190
rect 1930 18170 1950 18190
rect 1950 18170 1955 18190
rect 1925 18165 1955 18170
rect 2005 18190 2035 18195
rect 2005 18170 2010 18190
rect 2010 18170 2030 18190
rect 2030 18170 2035 18190
rect 2005 18165 2035 18170
rect 2085 18190 2115 18195
rect 2085 18170 2090 18190
rect 2090 18170 2110 18190
rect 2110 18170 2115 18190
rect 2085 18165 2115 18170
rect 2165 18190 2195 18195
rect 2165 18170 2170 18190
rect 2170 18170 2190 18190
rect 2190 18170 2195 18190
rect 2165 18165 2195 18170
rect 2245 18190 2275 18195
rect 2245 18170 2250 18190
rect 2250 18170 2270 18190
rect 2270 18170 2275 18190
rect 2245 18165 2275 18170
rect 2325 18190 2355 18195
rect 2325 18170 2330 18190
rect 2330 18170 2350 18190
rect 2350 18170 2355 18190
rect 2325 18165 2355 18170
rect 2405 18190 2435 18195
rect 2405 18170 2410 18190
rect 2410 18170 2430 18190
rect 2430 18170 2435 18190
rect 2405 18165 2435 18170
rect 2485 18190 2515 18195
rect 2485 18170 2490 18190
rect 2490 18170 2510 18190
rect 2510 18170 2515 18190
rect 2485 18165 2515 18170
rect 2565 18190 2595 18195
rect 2565 18170 2570 18190
rect 2570 18170 2590 18190
rect 2590 18170 2595 18190
rect 2565 18165 2595 18170
rect 2645 18190 2675 18195
rect 2645 18170 2650 18190
rect 2650 18170 2670 18190
rect 2670 18170 2675 18190
rect 2645 18165 2675 18170
rect 2725 18190 2755 18195
rect 2725 18170 2730 18190
rect 2730 18170 2750 18190
rect 2750 18170 2755 18190
rect 2725 18165 2755 18170
rect 2805 18190 2835 18195
rect 2805 18170 2810 18190
rect 2810 18170 2830 18190
rect 2830 18170 2835 18190
rect 2805 18165 2835 18170
rect 2885 18190 2915 18195
rect 2885 18170 2890 18190
rect 2890 18170 2910 18190
rect 2910 18170 2915 18190
rect 2885 18165 2915 18170
rect 2965 18190 2995 18195
rect 2965 18170 2970 18190
rect 2970 18170 2990 18190
rect 2990 18170 2995 18190
rect 2965 18165 2995 18170
rect 3045 18190 3075 18195
rect 3045 18170 3050 18190
rect 3050 18170 3070 18190
rect 3070 18170 3075 18190
rect 3045 18165 3075 18170
rect 3125 18190 3155 18195
rect 3125 18170 3130 18190
rect 3130 18170 3150 18190
rect 3150 18170 3155 18190
rect 3125 18165 3155 18170
rect 3205 18190 3235 18195
rect 3205 18170 3210 18190
rect 3210 18170 3230 18190
rect 3230 18170 3235 18190
rect 3205 18165 3235 18170
rect 3285 18190 3315 18195
rect 3285 18170 3290 18190
rect 3290 18170 3310 18190
rect 3310 18170 3315 18190
rect 3285 18165 3315 18170
rect 3365 18190 3395 18195
rect 3365 18170 3370 18190
rect 3370 18170 3390 18190
rect 3390 18170 3395 18190
rect 3365 18165 3395 18170
rect 3445 18190 3475 18195
rect 3445 18170 3450 18190
rect 3450 18170 3470 18190
rect 3470 18170 3475 18190
rect 3445 18165 3475 18170
rect 3525 18190 3555 18195
rect 3525 18170 3530 18190
rect 3530 18170 3550 18190
rect 3550 18170 3555 18190
rect 3525 18165 3555 18170
rect 3605 18190 3635 18195
rect 3605 18170 3610 18190
rect 3610 18170 3630 18190
rect 3630 18170 3635 18190
rect 3605 18165 3635 18170
rect 3685 18190 3715 18195
rect 3685 18170 3690 18190
rect 3690 18170 3710 18190
rect 3710 18170 3715 18190
rect 3685 18165 3715 18170
rect 3765 18190 3795 18195
rect 3765 18170 3770 18190
rect 3770 18170 3790 18190
rect 3790 18170 3795 18190
rect 3765 18165 3795 18170
rect 3845 18190 3875 18195
rect 3845 18170 3850 18190
rect 3850 18170 3870 18190
rect 3870 18170 3875 18190
rect 3845 18165 3875 18170
rect 3925 18190 3955 18195
rect 3925 18170 3930 18190
rect 3930 18170 3950 18190
rect 3950 18170 3955 18190
rect 3925 18165 3955 18170
rect 4005 18190 4035 18195
rect 4005 18170 4010 18190
rect 4010 18170 4030 18190
rect 4030 18170 4035 18190
rect 4005 18165 4035 18170
rect 4085 18190 4115 18195
rect 4085 18170 4090 18190
rect 4090 18170 4110 18190
rect 4110 18170 4115 18190
rect 4085 18165 4115 18170
rect 4165 18190 4195 18195
rect 4165 18170 4170 18190
rect 4170 18170 4190 18190
rect 4190 18170 4195 18190
rect 4165 18165 4195 18170
rect 6245 18190 6275 18195
rect 6245 18170 6250 18190
rect 6250 18170 6270 18190
rect 6270 18170 6275 18190
rect 6245 18165 6275 18170
rect 6325 18190 6355 18195
rect 6325 18170 6330 18190
rect 6330 18170 6350 18190
rect 6350 18170 6355 18190
rect 6325 18165 6355 18170
rect 6405 18190 6435 18195
rect 6405 18170 6410 18190
rect 6410 18170 6430 18190
rect 6430 18170 6435 18190
rect 6405 18165 6435 18170
rect 6485 18190 6515 18195
rect 6485 18170 6490 18190
rect 6490 18170 6510 18190
rect 6510 18170 6515 18190
rect 6485 18165 6515 18170
rect 6565 18190 6595 18195
rect 6565 18170 6570 18190
rect 6570 18170 6590 18190
rect 6590 18170 6595 18190
rect 6565 18165 6595 18170
rect 6645 18190 6675 18195
rect 6645 18170 6650 18190
rect 6650 18170 6670 18190
rect 6670 18170 6675 18190
rect 6645 18165 6675 18170
rect 6725 18190 6755 18195
rect 6725 18170 6730 18190
rect 6730 18170 6750 18190
rect 6750 18170 6755 18190
rect 6725 18165 6755 18170
rect 6805 18190 6835 18195
rect 6805 18170 6810 18190
rect 6810 18170 6830 18190
rect 6830 18170 6835 18190
rect 6805 18165 6835 18170
rect 6885 18190 6915 18195
rect 6885 18170 6890 18190
rect 6890 18170 6910 18190
rect 6910 18170 6915 18190
rect 6885 18165 6915 18170
rect 6965 18190 6995 18195
rect 6965 18170 6970 18190
rect 6970 18170 6990 18190
rect 6990 18170 6995 18190
rect 6965 18165 6995 18170
rect 7045 18190 7075 18195
rect 7045 18170 7050 18190
rect 7050 18170 7070 18190
rect 7070 18170 7075 18190
rect 7045 18165 7075 18170
rect 7125 18190 7155 18195
rect 7125 18170 7130 18190
rect 7130 18170 7150 18190
rect 7150 18170 7155 18190
rect 7125 18165 7155 18170
rect 7205 18190 7235 18195
rect 7205 18170 7210 18190
rect 7210 18170 7230 18190
rect 7230 18170 7235 18190
rect 7205 18165 7235 18170
rect 7285 18190 7315 18195
rect 7285 18170 7290 18190
rect 7290 18170 7310 18190
rect 7310 18170 7315 18190
rect 7285 18165 7315 18170
rect 7365 18190 7395 18195
rect 7365 18170 7370 18190
rect 7370 18170 7390 18190
rect 7390 18170 7395 18190
rect 7365 18165 7395 18170
rect 7445 18190 7475 18195
rect 7445 18170 7450 18190
rect 7450 18170 7470 18190
rect 7470 18170 7475 18190
rect 7445 18165 7475 18170
rect 7525 18190 7555 18195
rect 7525 18170 7530 18190
rect 7530 18170 7550 18190
rect 7550 18170 7555 18190
rect 7525 18165 7555 18170
rect 7605 18190 7635 18195
rect 7605 18170 7610 18190
rect 7610 18170 7630 18190
rect 7630 18170 7635 18190
rect 7605 18165 7635 18170
rect 7685 18190 7715 18195
rect 7685 18170 7690 18190
rect 7690 18170 7710 18190
rect 7710 18170 7715 18190
rect 7685 18165 7715 18170
rect 7765 18190 7795 18195
rect 7765 18170 7770 18190
rect 7770 18170 7790 18190
rect 7790 18170 7795 18190
rect 7765 18165 7795 18170
rect 7845 18190 7875 18195
rect 7845 18170 7850 18190
rect 7850 18170 7870 18190
rect 7870 18170 7875 18190
rect 7845 18165 7875 18170
rect 7925 18190 7955 18195
rect 7925 18170 7930 18190
rect 7930 18170 7950 18190
rect 7950 18170 7955 18190
rect 7925 18165 7955 18170
rect 8005 18190 8035 18195
rect 8005 18170 8010 18190
rect 8010 18170 8030 18190
rect 8030 18170 8035 18190
rect 8005 18165 8035 18170
rect 8085 18190 8115 18195
rect 8085 18170 8090 18190
rect 8090 18170 8110 18190
rect 8110 18170 8115 18190
rect 8085 18165 8115 18170
rect 8165 18190 8195 18195
rect 8165 18170 8170 18190
rect 8170 18170 8190 18190
rect 8190 18170 8195 18190
rect 8165 18165 8195 18170
rect 8245 18190 8275 18195
rect 8245 18170 8250 18190
rect 8250 18170 8270 18190
rect 8270 18170 8275 18190
rect 8245 18165 8275 18170
rect 8325 18190 8355 18195
rect 8325 18170 8330 18190
rect 8330 18170 8350 18190
rect 8350 18170 8355 18190
rect 8325 18165 8355 18170
rect 8405 18190 8435 18195
rect 8405 18170 8410 18190
rect 8410 18170 8430 18190
rect 8430 18170 8435 18190
rect 8405 18165 8435 18170
rect 8485 18190 8515 18195
rect 8485 18170 8490 18190
rect 8490 18170 8510 18190
rect 8510 18170 8515 18190
rect 8485 18165 8515 18170
rect 8565 18190 8595 18195
rect 8565 18170 8570 18190
rect 8570 18170 8590 18190
rect 8590 18170 8595 18190
rect 8565 18165 8595 18170
rect 8645 18190 8675 18195
rect 8645 18170 8650 18190
rect 8650 18170 8670 18190
rect 8670 18170 8675 18190
rect 8645 18165 8675 18170
rect 8725 18190 8755 18195
rect 8725 18170 8730 18190
rect 8730 18170 8750 18190
rect 8750 18170 8755 18190
rect 8725 18165 8755 18170
rect 8805 18190 8835 18195
rect 8805 18170 8810 18190
rect 8810 18170 8830 18190
rect 8830 18170 8835 18190
rect 8805 18165 8835 18170
rect 8885 18190 8915 18195
rect 8885 18170 8890 18190
rect 8890 18170 8910 18190
rect 8910 18170 8915 18190
rect 8885 18165 8915 18170
rect 8965 18190 8995 18195
rect 8965 18170 8970 18190
rect 8970 18170 8990 18190
rect 8990 18170 8995 18190
rect 8965 18165 8995 18170
rect 9045 18190 9075 18195
rect 9045 18170 9050 18190
rect 9050 18170 9070 18190
rect 9070 18170 9075 18190
rect 9045 18165 9075 18170
rect 9125 18190 9155 18195
rect 9125 18170 9130 18190
rect 9130 18170 9150 18190
rect 9150 18170 9155 18190
rect 9125 18165 9155 18170
rect 9205 18190 9235 18195
rect 9205 18170 9210 18190
rect 9210 18170 9230 18190
rect 9230 18170 9235 18190
rect 9205 18165 9235 18170
rect 9285 18190 9315 18195
rect 9285 18170 9290 18190
rect 9290 18170 9310 18190
rect 9310 18170 9315 18190
rect 9285 18165 9315 18170
rect 9365 18190 9395 18195
rect 9365 18170 9370 18190
rect 9370 18170 9390 18190
rect 9390 18170 9395 18190
rect 9365 18165 9395 18170
rect 9445 18190 9475 18195
rect 9445 18170 9450 18190
rect 9450 18170 9470 18190
rect 9470 18170 9475 18190
rect 9445 18165 9475 18170
rect 11565 18190 11595 18195
rect 11565 18170 11570 18190
rect 11570 18170 11590 18190
rect 11590 18170 11595 18190
rect 11565 18165 11595 18170
rect 11645 18190 11675 18195
rect 11645 18170 11650 18190
rect 11650 18170 11670 18190
rect 11670 18170 11675 18190
rect 11645 18165 11675 18170
rect 11725 18190 11755 18195
rect 11725 18170 11730 18190
rect 11730 18170 11750 18190
rect 11750 18170 11755 18190
rect 11725 18165 11755 18170
rect 11805 18190 11835 18195
rect 11805 18170 11810 18190
rect 11810 18170 11830 18190
rect 11830 18170 11835 18190
rect 11805 18165 11835 18170
rect 11885 18190 11915 18195
rect 11885 18170 11890 18190
rect 11890 18170 11910 18190
rect 11910 18170 11915 18190
rect 11885 18165 11915 18170
rect 11965 18190 11995 18195
rect 11965 18170 11970 18190
rect 11970 18170 11990 18190
rect 11990 18170 11995 18190
rect 11965 18165 11995 18170
rect 12045 18190 12075 18195
rect 12045 18170 12050 18190
rect 12050 18170 12070 18190
rect 12070 18170 12075 18190
rect 12045 18165 12075 18170
rect 12125 18190 12155 18195
rect 12125 18170 12130 18190
rect 12130 18170 12150 18190
rect 12150 18170 12155 18190
rect 12125 18165 12155 18170
rect 12205 18190 12235 18195
rect 12205 18170 12210 18190
rect 12210 18170 12230 18190
rect 12230 18170 12235 18190
rect 12205 18165 12235 18170
rect 12285 18190 12315 18195
rect 12285 18170 12290 18190
rect 12290 18170 12310 18190
rect 12310 18170 12315 18190
rect 12285 18165 12315 18170
rect 12365 18190 12395 18195
rect 12365 18170 12370 18190
rect 12370 18170 12390 18190
rect 12390 18170 12395 18190
rect 12365 18165 12395 18170
rect 12445 18190 12475 18195
rect 12445 18170 12450 18190
rect 12450 18170 12470 18190
rect 12470 18170 12475 18190
rect 12445 18165 12475 18170
rect 12525 18190 12555 18195
rect 12525 18170 12530 18190
rect 12530 18170 12550 18190
rect 12550 18170 12555 18190
rect 12525 18165 12555 18170
rect 12605 18190 12635 18195
rect 12605 18170 12610 18190
rect 12610 18170 12630 18190
rect 12630 18170 12635 18190
rect 12605 18165 12635 18170
rect 12685 18190 12715 18195
rect 12685 18170 12690 18190
rect 12690 18170 12710 18190
rect 12710 18170 12715 18190
rect 12685 18165 12715 18170
rect 12765 18190 12795 18195
rect 12765 18170 12770 18190
rect 12770 18170 12790 18190
rect 12790 18170 12795 18190
rect 12765 18165 12795 18170
rect 12845 18190 12875 18195
rect 12845 18170 12850 18190
rect 12850 18170 12870 18190
rect 12870 18170 12875 18190
rect 12845 18165 12875 18170
rect 12925 18190 12955 18195
rect 12925 18170 12930 18190
rect 12930 18170 12950 18190
rect 12950 18170 12955 18190
rect 12925 18165 12955 18170
rect 13005 18190 13035 18195
rect 13005 18170 13010 18190
rect 13010 18170 13030 18190
rect 13030 18170 13035 18190
rect 13005 18165 13035 18170
rect 13085 18190 13115 18195
rect 13085 18170 13090 18190
rect 13090 18170 13110 18190
rect 13110 18170 13115 18190
rect 13085 18165 13115 18170
rect 13165 18190 13195 18195
rect 13165 18170 13170 18190
rect 13170 18170 13190 18190
rect 13190 18170 13195 18190
rect 13165 18165 13195 18170
rect 13245 18190 13275 18195
rect 13245 18170 13250 18190
rect 13250 18170 13270 18190
rect 13270 18170 13275 18190
rect 13245 18165 13275 18170
rect 13325 18190 13355 18195
rect 13325 18170 13330 18190
rect 13330 18170 13350 18190
rect 13350 18170 13355 18190
rect 13325 18165 13355 18170
rect 13405 18190 13435 18195
rect 13405 18170 13410 18190
rect 13410 18170 13430 18190
rect 13430 18170 13435 18190
rect 13405 18165 13435 18170
rect 13485 18190 13515 18195
rect 13485 18170 13490 18190
rect 13490 18170 13510 18190
rect 13510 18170 13515 18190
rect 13485 18165 13515 18170
rect 13565 18190 13595 18195
rect 13565 18170 13570 18190
rect 13570 18170 13590 18190
rect 13590 18170 13595 18190
rect 13565 18165 13595 18170
rect 13645 18190 13675 18195
rect 13645 18170 13650 18190
rect 13650 18170 13670 18190
rect 13670 18170 13675 18190
rect 13645 18165 13675 18170
rect 13725 18190 13755 18195
rect 13725 18170 13730 18190
rect 13730 18170 13750 18190
rect 13750 18170 13755 18190
rect 13725 18165 13755 18170
rect 13805 18190 13835 18195
rect 13805 18170 13810 18190
rect 13810 18170 13830 18190
rect 13830 18170 13835 18190
rect 13805 18165 13835 18170
rect 13885 18190 13915 18195
rect 13885 18170 13890 18190
rect 13890 18170 13910 18190
rect 13910 18170 13915 18190
rect 13885 18165 13915 18170
rect 13965 18190 13995 18195
rect 13965 18170 13970 18190
rect 13970 18170 13990 18190
rect 13990 18170 13995 18190
rect 13965 18165 13995 18170
rect 14045 18190 14075 18195
rect 14045 18170 14050 18190
rect 14050 18170 14070 18190
rect 14070 18170 14075 18190
rect 14045 18165 14075 18170
rect 14125 18190 14155 18195
rect 14125 18170 14130 18190
rect 14130 18170 14150 18190
rect 14150 18170 14155 18190
rect 14125 18165 14155 18170
rect 14205 18190 14235 18195
rect 14205 18170 14210 18190
rect 14210 18170 14230 18190
rect 14230 18170 14235 18190
rect 14205 18165 14235 18170
rect 14285 18190 14315 18195
rect 14285 18170 14290 18190
rect 14290 18170 14310 18190
rect 14310 18170 14315 18190
rect 14285 18165 14315 18170
rect 14365 18190 14395 18195
rect 14365 18170 14370 18190
rect 14370 18170 14390 18190
rect 14390 18170 14395 18190
rect 14365 18165 14395 18170
rect 14445 18190 14475 18195
rect 14445 18170 14450 18190
rect 14450 18170 14470 18190
rect 14470 18170 14475 18190
rect 14445 18165 14475 18170
rect 14525 18190 14555 18195
rect 14525 18170 14530 18190
rect 14530 18170 14550 18190
rect 14550 18170 14555 18190
rect 14525 18165 14555 18170
rect 14605 18190 14635 18195
rect 14605 18170 14610 18190
rect 14610 18170 14630 18190
rect 14630 18170 14635 18190
rect 14605 18165 14635 18170
rect 14685 18190 14715 18195
rect 14685 18170 14690 18190
rect 14690 18170 14710 18190
rect 14710 18170 14715 18190
rect 14685 18165 14715 18170
rect 16765 18190 16795 18195
rect 16765 18170 16770 18190
rect 16770 18170 16790 18190
rect 16790 18170 16795 18190
rect 16765 18165 16795 18170
rect 16845 18190 16875 18195
rect 16845 18170 16850 18190
rect 16850 18170 16870 18190
rect 16870 18170 16875 18190
rect 16845 18165 16875 18170
rect 16925 18190 16955 18195
rect 16925 18170 16930 18190
rect 16930 18170 16950 18190
rect 16950 18170 16955 18190
rect 16925 18165 16955 18170
rect 17005 18190 17035 18195
rect 17005 18170 17010 18190
rect 17010 18170 17030 18190
rect 17030 18170 17035 18190
rect 17005 18165 17035 18170
rect 17085 18190 17115 18195
rect 17085 18170 17090 18190
rect 17090 18170 17110 18190
rect 17110 18170 17115 18190
rect 17085 18165 17115 18170
rect 17165 18190 17195 18195
rect 17165 18170 17170 18190
rect 17170 18170 17190 18190
rect 17190 18170 17195 18190
rect 17165 18165 17195 18170
rect 17245 18190 17275 18195
rect 17245 18170 17250 18190
rect 17250 18170 17270 18190
rect 17270 18170 17275 18190
rect 17245 18165 17275 18170
rect 17325 18190 17355 18195
rect 17325 18170 17330 18190
rect 17330 18170 17350 18190
rect 17350 18170 17355 18190
rect 17325 18165 17355 18170
rect 17405 18190 17435 18195
rect 17405 18170 17410 18190
rect 17410 18170 17430 18190
rect 17430 18170 17435 18190
rect 17405 18165 17435 18170
rect 17485 18190 17515 18195
rect 17485 18170 17490 18190
rect 17490 18170 17510 18190
rect 17510 18170 17515 18190
rect 17485 18165 17515 18170
rect 17565 18190 17595 18195
rect 17565 18170 17570 18190
rect 17570 18170 17590 18190
rect 17590 18170 17595 18190
rect 17565 18165 17595 18170
rect 17645 18190 17675 18195
rect 17645 18170 17650 18190
rect 17650 18170 17670 18190
rect 17670 18170 17675 18190
rect 17645 18165 17675 18170
rect 17725 18190 17755 18195
rect 17725 18170 17730 18190
rect 17730 18170 17750 18190
rect 17750 18170 17755 18190
rect 17725 18165 17755 18170
rect 17805 18190 17835 18195
rect 17805 18170 17810 18190
rect 17810 18170 17830 18190
rect 17830 18170 17835 18190
rect 17805 18165 17835 18170
rect 17885 18190 17915 18195
rect 17885 18170 17890 18190
rect 17890 18170 17910 18190
rect 17910 18170 17915 18190
rect 17885 18165 17915 18170
rect 17965 18190 17995 18195
rect 17965 18170 17970 18190
rect 17970 18170 17990 18190
rect 17990 18170 17995 18190
rect 17965 18165 17995 18170
rect 18045 18190 18075 18195
rect 18045 18170 18050 18190
rect 18050 18170 18070 18190
rect 18070 18170 18075 18190
rect 18045 18165 18075 18170
rect 18125 18190 18155 18195
rect 18125 18170 18130 18190
rect 18130 18170 18150 18190
rect 18150 18170 18155 18190
rect 18125 18165 18155 18170
rect 18205 18190 18235 18195
rect 18205 18170 18210 18190
rect 18210 18170 18230 18190
rect 18230 18170 18235 18190
rect 18205 18165 18235 18170
rect 18285 18190 18315 18195
rect 18285 18170 18290 18190
rect 18290 18170 18310 18190
rect 18310 18170 18315 18190
rect 18285 18165 18315 18170
rect 18365 18190 18395 18195
rect 18365 18170 18370 18190
rect 18370 18170 18390 18190
rect 18390 18170 18395 18190
rect 18365 18165 18395 18170
rect 18445 18190 18475 18195
rect 18445 18170 18450 18190
rect 18450 18170 18470 18190
rect 18470 18170 18475 18190
rect 18445 18165 18475 18170
rect 18525 18190 18555 18195
rect 18525 18170 18530 18190
rect 18530 18170 18550 18190
rect 18550 18170 18555 18190
rect 18525 18165 18555 18170
rect 18605 18190 18635 18195
rect 18605 18170 18610 18190
rect 18610 18170 18630 18190
rect 18630 18170 18635 18190
rect 18605 18165 18635 18170
rect 18685 18190 18715 18195
rect 18685 18170 18690 18190
rect 18690 18170 18710 18190
rect 18710 18170 18715 18190
rect 18685 18165 18715 18170
rect 18765 18190 18795 18195
rect 18765 18170 18770 18190
rect 18770 18170 18790 18190
rect 18790 18170 18795 18190
rect 18765 18165 18795 18170
rect 18845 18190 18875 18195
rect 18845 18170 18850 18190
rect 18850 18170 18870 18190
rect 18870 18170 18875 18190
rect 18845 18165 18875 18170
rect 18925 18190 18955 18195
rect 18925 18170 18930 18190
rect 18930 18170 18950 18190
rect 18950 18170 18955 18190
rect 18925 18165 18955 18170
rect 19005 18190 19035 18195
rect 19005 18170 19010 18190
rect 19010 18170 19030 18190
rect 19030 18170 19035 18190
rect 19005 18165 19035 18170
rect 19085 18190 19115 18195
rect 19085 18170 19090 18190
rect 19090 18170 19110 18190
rect 19110 18170 19115 18190
rect 19085 18165 19115 18170
rect 19165 18190 19195 18195
rect 19165 18170 19170 18190
rect 19170 18170 19190 18190
rect 19190 18170 19195 18190
rect 19165 18165 19195 18170
rect 19245 18190 19275 18195
rect 19245 18170 19250 18190
rect 19250 18170 19270 18190
rect 19270 18170 19275 18190
rect 19245 18165 19275 18170
rect 19325 18190 19355 18195
rect 19325 18170 19330 18190
rect 19330 18170 19350 18190
rect 19350 18170 19355 18190
rect 19325 18165 19355 18170
rect 19405 18190 19435 18195
rect 19405 18170 19410 18190
rect 19410 18170 19430 18190
rect 19430 18170 19435 18190
rect 19405 18165 19435 18170
rect 19485 18190 19515 18195
rect 19485 18170 19490 18190
rect 19490 18170 19510 18190
rect 19510 18170 19515 18190
rect 19485 18165 19515 18170
rect 19565 18190 19595 18195
rect 19565 18170 19570 18190
rect 19570 18170 19590 18190
rect 19590 18170 19595 18190
rect 19565 18165 19595 18170
rect 19645 18190 19675 18195
rect 19645 18170 19650 18190
rect 19650 18170 19670 18190
rect 19670 18170 19675 18190
rect 19645 18165 19675 18170
rect 19725 18190 19755 18195
rect 19725 18170 19730 18190
rect 19730 18170 19750 18190
rect 19750 18170 19755 18190
rect 19725 18165 19755 18170
rect 19805 18190 19835 18195
rect 19805 18170 19810 18190
rect 19810 18170 19830 18190
rect 19830 18170 19835 18190
rect 19805 18165 19835 18170
rect 19885 18190 19915 18195
rect 19885 18170 19890 18190
rect 19890 18170 19910 18190
rect 19910 18170 19915 18190
rect 19885 18165 19915 18170
rect 19965 18190 19995 18195
rect 19965 18170 19970 18190
rect 19970 18170 19990 18190
rect 19990 18170 19995 18190
rect 19965 18165 19995 18170
rect 20045 18190 20075 18195
rect 20045 18170 20050 18190
rect 20050 18170 20070 18190
rect 20070 18170 20075 18190
rect 20045 18165 20075 18170
rect 20125 18190 20155 18195
rect 20125 18170 20130 18190
rect 20130 18170 20150 18190
rect 20150 18170 20155 18190
rect 20125 18165 20155 18170
rect 20205 18190 20235 18195
rect 20205 18170 20210 18190
rect 20210 18170 20230 18190
rect 20230 18170 20235 18190
rect 20205 18165 20235 18170
rect 20285 18190 20315 18195
rect 20285 18170 20290 18190
rect 20290 18170 20310 18190
rect 20310 18170 20315 18190
rect 20285 18165 20315 18170
rect 20365 18190 20395 18195
rect 20365 18170 20370 18190
rect 20370 18170 20390 18190
rect 20390 18170 20395 18190
rect 20365 18165 20395 18170
rect 20445 18190 20475 18195
rect 20445 18170 20450 18190
rect 20450 18170 20470 18190
rect 20470 18170 20475 18190
rect 20445 18165 20475 18170
rect 20525 18190 20555 18195
rect 20525 18170 20530 18190
rect 20530 18170 20550 18190
rect 20550 18170 20555 18190
rect 20525 18165 20555 18170
rect 20605 18190 20635 18195
rect 20605 18170 20610 18190
rect 20610 18170 20630 18190
rect 20630 18170 20635 18190
rect 20605 18165 20635 18170
rect 20685 18190 20715 18195
rect 20685 18170 20690 18190
rect 20690 18170 20710 18190
rect 20710 18170 20715 18190
rect 20685 18165 20715 18170
rect 20765 18190 20795 18195
rect 20765 18170 20770 18190
rect 20770 18170 20790 18190
rect 20790 18170 20795 18190
rect 20765 18165 20795 18170
rect 20845 18190 20875 18195
rect 20845 18170 20850 18190
rect 20850 18170 20870 18190
rect 20870 18170 20875 18190
rect 20845 18165 20875 18170
rect 20925 18190 20955 18195
rect 20925 18170 20930 18190
rect 20930 18170 20950 18190
rect 20950 18170 20955 18190
rect 20925 18165 20955 18170
rect 5 18030 35 18035
rect 5 18010 10 18030
rect 10 18010 30 18030
rect 30 18010 35 18030
rect 5 18005 35 18010
rect 85 18030 115 18035
rect 85 18010 90 18030
rect 90 18010 110 18030
rect 110 18010 115 18030
rect 85 18005 115 18010
rect 165 18030 195 18035
rect 165 18010 170 18030
rect 170 18010 190 18030
rect 190 18010 195 18030
rect 165 18005 195 18010
rect 245 18030 275 18035
rect 245 18010 250 18030
rect 250 18010 270 18030
rect 270 18010 275 18030
rect 245 18005 275 18010
rect 325 18030 355 18035
rect 325 18010 330 18030
rect 330 18010 350 18030
rect 350 18010 355 18030
rect 325 18005 355 18010
rect 405 18030 435 18035
rect 405 18010 410 18030
rect 410 18010 430 18030
rect 430 18010 435 18030
rect 405 18005 435 18010
rect 485 18030 515 18035
rect 485 18010 490 18030
rect 490 18010 510 18030
rect 510 18010 515 18030
rect 485 18005 515 18010
rect 565 18030 595 18035
rect 565 18010 570 18030
rect 570 18010 590 18030
rect 590 18010 595 18030
rect 565 18005 595 18010
rect 645 18030 675 18035
rect 645 18010 650 18030
rect 650 18010 670 18030
rect 670 18010 675 18030
rect 645 18005 675 18010
rect 725 18030 755 18035
rect 725 18010 730 18030
rect 730 18010 750 18030
rect 750 18010 755 18030
rect 725 18005 755 18010
rect 805 18030 835 18035
rect 805 18010 810 18030
rect 810 18010 830 18030
rect 830 18010 835 18030
rect 805 18005 835 18010
rect 885 18030 915 18035
rect 885 18010 890 18030
rect 890 18010 910 18030
rect 910 18010 915 18030
rect 885 18005 915 18010
rect 965 18030 995 18035
rect 965 18010 970 18030
rect 970 18010 990 18030
rect 990 18010 995 18030
rect 965 18005 995 18010
rect 1045 18030 1075 18035
rect 1045 18010 1050 18030
rect 1050 18010 1070 18030
rect 1070 18010 1075 18030
rect 1045 18005 1075 18010
rect 1125 18030 1155 18035
rect 1125 18010 1130 18030
rect 1130 18010 1150 18030
rect 1150 18010 1155 18030
rect 1125 18005 1155 18010
rect 1205 18030 1235 18035
rect 1205 18010 1210 18030
rect 1210 18010 1230 18030
rect 1230 18010 1235 18030
rect 1205 18005 1235 18010
rect 1285 18030 1315 18035
rect 1285 18010 1290 18030
rect 1290 18010 1310 18030
rect 1310 18010 1315 18030
rect 1285 18005 1315 18010
rect 1365 18030 1395 18035
rect 1365 18010 1370 18030
rect 1370 18010 1390 18030
rect 1390 18010 1395 18030
rect 1365 18005 1395 18010
rect 1445 18030 1475 18035
rect 1445 18010 1450 18030
rect 1450 18010 1470 18030
rect 1470 18010 1475 18030
rect 1445 18005 1475 18010
rect 1525 18030 1555 18035
rect 1525 18010 1530 18030
rect 1530 18010 1550 18030
rect 1550 18010 1555 18030
rect 1525 18005 1555 18010
rect 1605 18030 1635 18035
rect 1605 18010 1610 18030
rect 1610 18010 1630 18030
rect 1630 18010 1635 18030
rect 1605 18005 1635 18010
rect 1685 18030 1715 18035
rect 1685 18010 1690 18030
rect 1690 18010 1710 18030
rect 1710 18010 1715 18030
rect 1685 18005 1715 18010
rect 1765 18030 1795 18035
rect 1765 18010 1770 18030
rect 1770 18010 1790 18030
rect 1790 18010 1795 18030
rect 1765 18005 1795 18010
rect 1845 18030 1875 18035
rect 1845 18010 1850 18030
rect 1850 18010 1870 18030
rect 1870 18010 1875 18030
rect 1845 18005 1875 18010
rect 1925 18030 1955 18035
rect 1925 18010 1930 18030
rect 1930 18010 1950 18030
rect 1950 18010 1955 18030
rect 1925 18005 1955 18010
rect 2005 18030 2035 18035
rect 2005 18010 2010 18030
rect 2010 18010 2030 18030
rect 2030 18010 2035 18030
rect 2005 18005 2035 18010
rect 2085 18030 2115 18035
rect 2085 18010 2090 18030
rect 2090 18010 2110 18030
rect 2110 18010 2115 18030
rect 2085 18005 2115 18010
rect 2165 18030 2195 18035
rect 2165 18010 2170 18030
rect 2170 18010 2190 18030
rect 2190 18010 2195 18030
rect 2165 18005 2195 18010
rect 2245 18030 2275 18035
rect 2245 18010 2250 18030
rect 2250 18010 2270 18030
rect 2270 18010 2275 18030
rect 2245 18005 2275 18010
rect 2325 18030 2355 18035
rect 2325 18010 2330 18030
rect 2330 18010 2350 18030
rect 2350 18010 2355 18030
rect 2325 18005 2355 18010
rect 2405 18030 2435 18035
rect 2405 18010 2410 18030
rect 2410 18010 2430 18030
rect 2430 18010 2435 18030
rect 2405 18005 2435 18010
rect 2485 18030 2515 18035
rect 2485 18010 2490 18030
rect 2490 18010 2510 18030
rect 2510 18010 2515 18030
rect 2485 18005 2515 18010
rect 2565 18030 2595 18035
rect 2565 18010 2570 18030
rect 2570 18010 2590 18030
rect 2590 18010 2595 18030
rect 2565 18005 2595 18010
rect 2645 18030 2675 18035
rect 2645 18010 2650 18030
rect 2650 18010 2670 18030
rect 2670 18010 2675 18030
rect 2645 18005 2675 18010
rect 2725 18030 2755 18035
rect 2725 18010 2730 18030
rect 2730 18010 2750 18030
rect 2750 18010 2755 18030
rect 2725 18005 2755 18010
rect 2805 18030 2835 18035
rect 2805 18010 2810 18030
rect 2810 18010 2830 18030
rect 2830 18010 2835 18030
rect 2805 18005 2835 18010
rect 2885 18030 2915 18035
rect 2885 18010 2890 18030
rect 2890 18010 2910 18030
rect 2910 18010 2915 18030
rect 2885 18005 2915 18010
rect 2965 18030 2995 18035
rect 2965 18010 2970 18030
rect 2970 18010 2990 18030
rect 2990 18010 2995 18030
rect 2965 18005 2995 18010
rect 3045 18030 3075 18035
rect 3045 18010 3050 18030
rect 3050 18010 3070 18030
rect 3070 18010 3075 18030
rect 3045 18005 3075 18010
rect 3125 18030 3155 18035
rect 3125 18010 3130 18030
rect 3130 18010 3150 18030
rect 3150 18010 3155 18030
rect 3125 18005 3155 18010
rect 3205 18030 3235 18035
rect 3205 18010 3210 18030
rect 3210 18010 3230 18030
rect 3230 18010 3235 18030
rect 3205 18005 3235 18010
rect 3285 18030 3315 18035
rect 3285 18010 3290 18030
rect 3290 18010 3310 18030
rect 3310 18010 3315 18030
rect 3285 18005 3315 18010
rect 3365 18030 3395 18035
rect 3365 18010 3370 18030
rect 3370 18010 3390 18030
rect 3390 18010 3395 18030
rect 3365 18005 3395 18010
rect 3445 18030 3475 18035
rect 3445 18010 3450 18030
rect 3450 18010 3470 18030
rect 3470 18010 3475 18030
rect 3445 18005 3475 18010
rect 3525 18030 3555 18035
rect 3525 18010 3530 18030
rect 3530 18010 3550 18030
rect 3550 18010 3555 18030
rect 3525 18005 3555 18010
rect 3605 18030 3635 18035
rect 3605 18010 3610 18030
rect 3610 18010 3630 18030
rect 3630 18010 3635 18030
rect 3605 18005 3635 18010
rect 3685 18030 3715 18035
rect 3685 18010 3690 18030
rect 3690 18010 3710 18030
rect 3710 18010 3715 18030
rect 3685 18005 3715 18010
rect 3765 18030 3795 18035
rect 3765 18010 3770 18030
rect 3770 18010 3790 18030
rect 3790 18010 3795 18030
rect 3765 18005 3795 18010
rect 3845 18030 3875 18035
rect 3845 18010 3850 18030
rect 3850 18010 3870 18030
rect 3870 18010 3875 18030
rect 3845 18005 3875 18010
rect 3925 18030 3955 18035
rect 3925 18010 3930 18030
rect 3930 18010 3950 18030
rect 3950 18010 3955 18030
rect 3925 18005 3955 18010
rect 4005 18030 4035 18035
rect 4005 18010 4010 18030
rect 4010 18010 4030 18030
rect 4030 18010 4035 18030
rect 4005 18005 4035 18010
rect 4085 18030 4115 18035
rect 4085 18010 4090 18030
rect 4090 18010 4110 18030
rect 4110 18010 4115 18030
rect 4085 18005 4115 18010
rect 4165 18030 4195 18035
rect 4165 18010 4170 18030
rect 4170 18010 4190 18030
rect 4190 18010 4195 18030
rect 4165 18005 4195 18010
rect 6245 18030 6275 18035
rect 6245 18010 6250 18030
rect 6250 18010 6270 18030
rect 6270 18010 6275 18030
rect 6245 18005 6275 18010
rect 6325 18030 6355 18035
rect 6325 18010 6330 18030
rect 6330 18010 6350 18030
rect 6350 18010 6355 18030
rect 6325 18005 6355 18010
rect 6405 18030 6435 18035
rect 6405 18010 6410 18030
rect 6410 18010 6430 18030
rect 6430 18010 6435 18030
rect 6405 18005 6435 18010
rect 6485 18030 6515 18035
rect 6485 18010 6490 18030
rect 6490 18010 6510 18030
rect 6510 18010 6515 18030
rect 6485 18005 6515 18010
rect 6565 18030 6595 18035
rect 6565 18010 6570 18030
rect 6570 18010 6590 18030
rect 6590 18010 6595 18030
rect 6565 18005 6595 18010
rect 6645 18030 6675 18035
rect 6645 18010 6650 18030
rect 6650 18010 6670 18030
rect 6670 18010 6675 18030
rect 6645 18005 6675 18010
rect 6725 18030 6755 18035
rect 6725 18010 6730 18030
rect 6730 18010 6750 18030
rect 6750 18010 6755 18030
rect 6725 18005 6755 18010
rect 6805 18030 6835 18035
rect 6805 18010 6810 18030
rect 6810 18010 6830 18030
rect 6830 18010 6835 18030
rect 6805 18005 6835 18010
rect 6885 18030 6915 18035
rect 6885 18010 6890 18030
rect 6890 18010 6910 18030
rect 6910 18010 6915 18030
rect 6885 18005 6915 18010
rect 6965 18030 6995 18035
rect 6965 18010 6970 18030
rect 6970 18010 6990 18030
rect 6990 18010 6995 18030
rect 6965 18005 6995 18010
rect 7045 18030 7075 18035
rect 7045 18010 7050 18030
rect 7050 18010 7070 18030
rect 7070 18010 7075 18030
rect 7045 18005 7075 18010
rect 7125 18030 7155 18035
rect 7125 18010 7130 18030
rect 7130 18010 7150 18030
rect 7150 18010 7155 18030
rect 7125 18005 7155 18010
rect 7205 18030 7235 18035
rect 7205 18010 7210 18030
rect 7210 18010 7230 18030
rect 7230 18010 7235 18030
rect 7205 18005 7235 18010
rect 7285 18030 7315 18035
rect 7285 18010 7290 18030
rect 7290 18010 7310 18030
rect 7310 18010 7315 18030
rect 7285 18005 7315 18010
rect 7365 18030 7395 18035
rect 7365 18010 7370 18030
rect 7370 18010 7390 18030
rect 7390 18010 7395 18030
rect 7365 18005 7395 18010
rect 7445 18030 7475 18035
rect 7445 18010 7450 18030
rect 7450 18010 7470 18030
rect 7470 18010 7475 18030
rect 7445 18005 7475 18010
rect 7525 18030 7555 18035
rect 7525 18010 7530 18030
rect 7530 18010 7550 18030
rect 7550 18010 7555 18030
rect 7525 18005 7555 18010
rect 7605 18030 7635 18035
rect 7605 18010 7610 18030
rect 7610 18010 7630 18030
rect 7630 18010 7635 18030
rect 7605 18005 7635 18010
rect 7685 18030 7715 18035
rect 7685 18010 7690 18030
rect 7690 18010 7710 18030
rect 7710 18010 7715 18030
rect 7685 18005 7715 18010
rect 7765 18030 7795 18035
rect 7765 18010 7770 18030
rect 7770 18010 7790 18030
rect 7790 18010 7795 18030
rect 7765 18005 7795 18010
rect 7845 18030 7875 18035
rect 7845 18010 7850 18030
rect 7850 18010 7870 18030
rect 7870 18010 7875 18030
rect 7845 18005 7875 18010
rect 7925 18030 7955 18035
rect 7925 18010 7930 18030
rect 7930 18010 7950 18030
rect 7950 18010 7955 18030
rect 7925 18005 7955 18010
rect 8005 18030 8035 18035
rect 8005 18010 8010 18030
rect 8010 18010 8030 18030
rect 8030 18010 8035 18030
rect 8005 18005 8035 18010
rect 8085 18030 8115 18035
rect 8085 18010 8090 18030
rect 8090 18010 8110 18030
rect 8110 18010 8115 18030
rect 8085 18005 8115 18010
rect 8165 18030 8195 18035
rect 8165 18010 8170 18030
rect 8170 18010 8190 18030
rect 8190 18010 8195 18030
rect 8165 18005 8195 18010
rect 8245 18030 8275 18035
rect 8245 18010 8250 18030
rect 8250 18010 8270 18030
rect 8270 18010 8275 18030
rect 8245 18005 8275 18010
rect 8325 18030 8355 18035
rect 8325 18010 8330 18030
rect 8330 18010 8350 18030
rect 8350 18010 8355 18030
rect 8325 18005 8355 18010
rect 8405 18030 8435 18035
rect 8405 18010 8410 18030
rect 8410 18010 8430 18030
rect 8430 18010 8435 18030
rect 8405 18005 8435 18010
rect 8485 18030 8515 18035
rect 8485 18010 8490 18030
rect 8490 18010 8510 18030
rect 8510 18010 8515 18030
rect 8485 18005 8515 18010
rect 8565 18030 8595 18035
rect 8565 18010 8570 18030
rect 8570 18010 8590 18030
rect 8590 18010 8595 18030
rect 8565 18005 8595 18010
rect 8645 18030 8675 18035
rect 8645 18010 8650 18030
rect 8650 18010 8670 18030
rect 8670 18010 8675 18030
rect 8645 18005 8675 18010
rect 8725 18030 8755 18035
rect 8725 18010 8730 18030
rect 8730 18010 8750 18030
rect 8750 18010 8755 18030
rect 8725 18005 8755 18010
rect 8805 18030 8835 18035
rect 8805 18010 8810 18030
rect 8810 18010 8830 18030
rect 8830 18010 8835 18030
rect 8805 18005 8835 18010
rect 8885 18030 8915 18035
rect 8885 18010 8890 18030
rect 8890 18010 8910 18030
rect 8910 18010 8915 18030
rect 8885 18005 8915 18010
rect 8965 18030 8995 18035
rect 8965 18010 8970 18030
rect 8970 18010 8990 18030
rect 8990 18010 8995 18030
rect 8965 18005 8995 18010
rect 9045 18030 9075 18035
rect 9045 18010 9050 18030
rect 9050 18010 9070 18030
rect 9070 18010 9075 18030
rect 9045 18005 9075 18010
rect 9125 18030 9155 18035
rect 9125 18010 9130 18030
rect 9130 18010 9150 18030
rect 9150 18010 9155 18030
rect 9125 18005 9155 18010
rect 9205 18030 9235 18035
rect 9205 18010 9210 18030
rect 9210 18010 9230 18030
rect 9230 18010 9235 18030
rect 9205 18005 9235 18010
rect 9285 18030 9315 18035
rect 9285 18010 9290 18030
rect 9290 18010 9310 18030
rect 9310 18010 9315 18030
rect 9285 18005 9315 18010
rect 9365 18030 9395 18035
rect 9365 18010 9370 18030
rect 9370 18010 9390 18030
rect 9390 18010 9395 18030
rect 9365 18005 9395 18010
rect 9445 18030 9475 18035
rect 9445 18010 9450 18030
rect 9450 18010 9470 18030
rect 9470 18010 9475 18030
rect 9445 18005 9475 18010
rect 11565 18030 11595 18035
rect 11565 18010 11570 18030
rect 11570 18010 11590 18030
rect 11590 18010 11595 18030
rect 11565 18005 11595 18010
rect 11645 18030 11675 18035
rect 11645 18010 11650 18030
rect 11650 18010 11670 18030
rect 11670 18010 11675 18030
rect 11645 18005 11675 18010
rect 11725 18030 11755 18035
rect 11725 18010 11730 18030
rect 11730 18010 11750 18030
rect 11750 18010 11755 18030
rect 11725 18005 11755 18010
rect 11805 18030 11835 18035
rect 11805 18010 11810 18030
rect 11810 18010 11830 18030
rect 11830 18010 11835 18030
rect 11805 18005 11835 18010
rect 11885 18030 11915 18035
rect 11885 18010 11890 18030
rect 11890 18010 11910 18030
rect 11910 18010 11915 18030
rect 11885 18005 11915 18010
rect 11965 18030 11995 18035
rect 11965 18010 11970 18030
rect 11970 18010 11990 18030
rect 11990 18010 11995 18030
rect 11965 18005 11995 18010
rect 12045 18030 12075 18035
rect 12045 18010 12050 18030
rect 12050 18010 12070 18030
rect 12070 18010 12075 18030
rect 12045 18005 12075 18010
rect 12125 18030 12155 18035
rect 12125 18010 12130 18030
rect 12130 18010 12150 18030
rect 12150 18010 12155 18030
rect 12125 18005 12155 18010
rect 12205 18030 12235 18035
rect 12205 18010 12210 18030
rect 12210 18010 12230 18030
rect 12230 18010 12235 18030
rect 12205 18005 12235 18010
rect 12285 18030 12315 18035
rect 12285 18010 12290 18030
rect 12290 18010 12310 18030
rect 12310 18010 12315 18030
rect 12285 18005 12315 18010
rect 12365 18030 12395 18035
rect 12365 18010 12370 18030
rect 12370 18010 12390 18030
rect 12390 18010 12395 18030
rect 12365 18005 12395 18010
rect 12445 18030 12475 18035
rect 12445 18010 12450 18030
rect 12450 18010 12470 18030
rect 12470 18010 12475 18030
rect 12445 18005 12475 18010
rect 12525 18030 12555 18035
rect 12525 18010 12530 18030
rect 12530 18010 12550 18030
rect 12550 18010 12555 18030
rect 12525 18005 12555 18010
rect 12605 18030 12635 18035
rect 12605 18010 12610 18030
rect 12610 18010 12630 18030
rect 12630 18010 12635 18030
rect 12605 18005 12635 18010
rect 12685 18030 12715 18035
rect 12685 18010 12690 18030
rect 12690 18010 12710 18030
rect 12710 18010 12715 18030
rect 12685 18005 12715 18010
rect 12765 18030 12795 18035
rect 12765 18010 12770 18030
rect 12770 18010 12790 18030
rect 12790 18010 12795 18030
rect 12765 18005 12795 18010
rect 12845 18030 12875 18035
rect 12845 18010 12850 18030
rect 12850 18010 12870 18030
rect 12870 18010 12875 18030
rect 12845 18005 12875 18010
rect 12925 18030 12955 18035
rect 12925 18010 12930 18030
rect 12930 18010 12950 18030
rect 12950 18010 12955 18030
rect 12925 18005 12955 18010
rect 13005 18030 13035 18035
rect 13005 18010 13010 18030
rect 13010 18010 13030 18030
rect 13030 18010 13035 18030
rect 13005 18005 13035 18010
rect 13085 18030 13115 18035
rect 13085 18010 13090 18030
rect 13090 18010 13110 18030
rect 13110 18010 13115 18030
rect 13085 18005 13115 18010
rect 13165 18030 13195 18035
rect 13165 18010 13170 18030
rect 13170 18010 13190 18030
rect 13190 18010 13195 18030
rect 13165 18005 13195 18010
rect 13245 18030 13275 18035
rect 13245 18010 13250 18030
rect 13250 18010 13270 18030
rect 13270 18010 13275 18030
rect 13245 18005 13275 18010
rect 13325 18030 13355 18035
rect 13325 18010 13330 18030
rect 13330 18010 13350 18030
rect 13350 18010 13355 18030
rect 13325 18005 13355 18010
rect 13405 18030 13435 18035
rect 13405 18010 13410 18030
rect 13410 18010 13430 18030
rect 13430 18010 13435 18030
rect 13405 18005 13435 18010
rect 13485 18030 13515 18035
rect 13485 18010 13490 18030
rect 13490 18010 13510 18030
rect 13510 18010 13515 18030
rect 13485 18005 13515 18010
rect 13565 18030 13595 18035
rect 13565 18010 13570 18030
rect 13570 18010 13590 18030
rect 13590 18010 13595 18030
rect 13565 18005 13595 18010
rect 13645 18030 13675 18035
rect 13645 18010 13650 18030
rect 13650 18010 13670 18030
rect 13670 18010 13675 18030
rect 13645 18005 13675 18010
rect 13725 18030 13755 18035
rect 13725 18010 13730 18030
rect 13730 18010 13750 18030
rect 13750 18010 13755 18030
rect 13725 18005 13755 18010
rect 13805 18030 13835 18035
rect 13805 18010 13810 18030
rect 13810 18010 13830 18030
rect 13830 18010 13835 18030
rect 13805 18005 13835 18010
rect 13885 18030 13915 18035
rect 13885 18010 13890 18030
rect 13890 18010 13910 18030
rect 13910 18010 13915 18030
rect 13885 18005 13915 18010
rect 13965 18030 13995 18035
rect 13965 18010 13970 18030
rect 13970 18010 13990 18030
rect 13990 18010 13995 18030
rect 13965 18005 13995 18010
rect 14045 18030 14075 18035
rect 14045 18010 14050 18030
rect 14050 18010 14070 18030
rect 14070 18010 14075 18030
rect 14045 18005 14075 18010
rect 14125 18030 14155 18035
rect 14125 18010 14130 18030
rect 14130 18010 14150 18030
rect 14150 18010 14155 18030
rect 14125 18005 14155 18010
rect 14205 18030 14235 18035
rect 14205 18010 14210 18030
rect 14210 18010 14230 18030
rect 14230 18010 14235 18030
rect 14205 18005 14235 18010
rect 14285 18030 14315 18035
rect 14285 18010 14290 18030
rect 14290 18010 14310 18030
rect 14310 18010 14315 18030
rect 14285 18005 14315 18010
rect 14365 18030 14395 18035
rect 14365 18010 14370 18030
rect 14370 18010 14390 18030
rect 14390 18010 14395 18030
rect 14365 18005 14395 18010
rect 14445 18030 14475 18035
rect 14445 18010 14450 18030
rect 14450 18010 14470 18030
rect 14470 18010 14475 18030
rect 14445 18005 14475 18010
rect 14525 18030 14555 18035
rect 14525 18010 14530 18030
rect 14530 18010 14550 18030
rect 14550 18010 14555 18030
rect 14525 18005 14555 18010
rect 14605 18030 14635 18035
rect 14605 18010 14610 18030
rect 14610 18010 14630 18030
rect 14630 18010 14635 18030
rect 14605 18005 14635 18010
rect 14685 18030 14715 18035
rect 14685 18010 14690 18030
rect 14690 18010 14710 18030
rect 14710 18010 14715 18030
rect 14685 18005 14715 18010
rect 16765 18030 16795 18035
rect 16765 18010 16770 18030
rect 16770 18010 16790 18030
rect 16790 18010 16795 18030
rect 16765 18005 16795 18010
rect 16845 18030 16875 18035
rect 16845 18010 16850 18030
rect 16850 18010 16870 18030
rect 16870 18010 16875 18030
rect 16845 18005 16875 18010
rect 16925 18030 16955 18035
rect 16925 18010 16930 18030
rect 16930 18010 16950 18030
rect 16950 18010 16955 18030
rect 16925 18005 16955 18010
rect 17005 18030 17035 18035
rect 17005 18010 17010 18030
rect 17010 18010 17030 18030
rect 17030 18010 17035 18030
rect 17005 18005 17035 18010
rect 17085 18030 17115 18035
rect 17085 18010 17090 18030
rect 17090 18010 17110 18030
rect 17110 18010 17115 18030
rect 17085 18005 17115 18010
rect 17165 18030 17195 18035
rect 17165 18010 17170 18030
rect 17170 18010 17190 18030
rect 17190 18010 17195 18030
rect 17165 18005 17195 18010
rect 17245 18030 17275 18035
rect 17245 18010 17250 18030
rect 17250 18010 17270 18030
rect 17270 18010 17275 18030
rect 17245 18005 17275 18010
rect 17325 18030 17355 18035
rect 17325 18010 17330 18030
rect 17330 18010 17350 18030
rect 17350 18010 17355 18030
rect 17325 18005 17355 18010
rect 17405 18030 17435 18035
rect 17405 18010 17410 18030
rect 17410 18010 17430 18030
rect 17430 18010 17435 18030
rect 17405 18005 17435 18010
rect 17485 18030 17515 18035
rect 17485 18010 17490 18030
rect 17490 18010 17510 18030
rect 17510 18010 17515 18030
rect 17485 18005 17515 18010
rect 17565 18030 17595 18035
rect 17565 18010 17570 18030
rect 17570 18010 17590 18030
rect 17590 18010 17595 18030
rect 17565 18005 17595 18010
rect 17645 18030 17675 18035
rect 17645 18010 17650 18030
rect 17650 18010 17670 18030
rect 17670 18010 17675 18030
rect 17645 18005 17675 18010
rect 17725 18030 17755 18035
rect 17725 18010 17730 18030
rect 17730 18010 17750 18030
rect 17750 18010 17755 18030
rect 17725 18005 17755 18010
rect 17805 18030 17835 18035
rect 17805 18010 17810 18030
rect 17810 18010 17830 18030
rect 17830 18010 17835 18030
rect 17805 18005 17835 18010
rect 17885 18030 17915 18035
rect 17885 18010 17890 18030
rect 17890 18010 17910 18030
rect 17910 18010 17915 18030
rect 17885 18005 17915 18010
rect 17965 18030 17995 18035
rect 17965 18010 17970 18030
rect 17970 18010 17990 18030
rect 17990 18010 17995 18030
rect 17965 18005 17995 18010
rect 18045 18030 18075 18035
rect 18045 18010 18050 18030
rect 18050 18010 18070 18030
rect 18070 18010 18075 18030
rect 18045 18005 18075 18010
rect 18125 18030 18155 18035
rect 18125 18010 18130 18030
rect 18130 18010 18150 18030
rect 18150 18010 18155 18030
rect 18125 18005 18155 18010
rect 18205 18030 18235 18035
rect 18205 18010 18210 18030
rect 18210 18010 18230 18030
rect 18230 18010 18235 18030
rect 18205 18005 18235 18010
rect 18285 18030 18315 18035
rect 18285 18010 18290 18030
rect 18290 18010 18310 18030
rect 18310 18010 18315 18030
rect 18285 18005 18315 18010
rect 18365 18030 18395 18035
rect 18365 18010 18370 18030
rect 18370 18010 18390 18030
rect 18390 18010 18395 18030
rect 18365 18005 18395 18010
rect 18445 18030 18475 18035
rect 18445 18010 18450 18030
rect 18450 18010 18470 18030
rect 18470 18010 18475 18030
rect 18445 18005 18475 18010
rect 18525 18030 18555 18035
rect 18525 18010 18530 18030
rect 18530 18010 18550 18030
rect 18550 18010 18555 18030
rect 18525 18005 18555 18010
rect 18605 18030 18635 18035
rect 18605 18010 18610 18030
rect 18610 18010 18630 18030
rect 18630 18010 18635 18030
rect 18605 18005 18635 18010
rect 18685 18030 18715 18035
rect 18685 18010 18690 18030
rect 18690 18010 18710 18030
rect 18710 18010 18715 18030
rect 18685 18005 18715 18010
rect 18765 18030 18795 18035
rect 18765 18010 18770 18030
rect 18770 18010 18790 18030
rect 18790 18010 18795 18030
rect 18765 18005 18795 18010
rect 18845 18030 18875 18035
rect 18845 18010 18850 18030
rect 18850 18010 18870 18030
rect 18870 18010 18875 18030
rect 18845 18005 18875 18010
rect 18925 18030 18955 18035
rect 18925 18010 18930 18030
rect 18930 18010 18950 18030
rect 18950 18010 18955 18030
rect 18925 18005 18955 18010
rect 19005 18030 19035 18035
rect 19005 18010 19010 18030
rect 19010 18010 19030 18030
rect 19030 18010 19035 18030
rect 19005 18005 19035 18010
rect 19085 18030 19115 18035
rect 19085 18010 19090 18030
rect 19090 18010 19110 18030
rect 19110 18010 19115 18030
rect 19085 18005 19115 18010
rect 19165 18030 19195 18035
rect 19165 18010 19170 18030
rect 19170 18010 19190 18030
rect 19190 18010 19195 18030
rect 19165 18005 19195 18010
rect 19245 18030 19275 18035
rect 19245 18010 19250 18030
rect 19250 18010 19270 18030
rect 19270 18010 19275 18030
rect 19245 18005 19275 18010
rect 19325 18030 19355 18035
rect 19325 18010 19330 18030
rect 19330 18010 19350 18030
rect 19350 18010 19355 18030
rect 19325 18005 19355 18010
rect 19405 18030 19435 18035
rect 19405 18010 19410 18030
rect 19410 18010 19430 18030
rect 19430 18010 19435 18030
rect 19405 18005 19435 18010
rect 19485 18030 19515 18035
rect 19485 18010 19490 18030
rect 19490 18010 19510 18030
rect 19510 18010 19515 18030
rect 19485 18005 19515 18010
rect 19565 18030 19595 18035
rect 19565 18010 19570 18030
rect 19570 18010 19590 18030
rect 19590 18010 19595 18030
rect 19565 18005 19595 18010
rect 19645 18030 19675 18035
rect 19645 18010 19650 18030
rect 19650 18010 19670 18030
rect 19670 18010 19675 18030
rect 19645 18005 19675 18010
rect 19725 18030 19755 18035
rect 19725 18010 19730 18030
rect 19730 18010 19750 18030
rect 19750 18010 19755 18030
rect 19725 18005 19755 18010
rect 19805 18030 19835 18035
rect 19805 18010 19810 18030
rect 19810 18010 19830 18030
rect 19830 18010 19835 18030
rect 19805 18005 19835 18010
rect 19885 18030 19915 18035
rect 19885 18010 19890 18030
rect 19890 18010 19910 18030
rect 19910 18010 19915 18030
rect 19885 18005 19915 18010
rect 19965 18030 19995 18035
rect 19965 18010 19970 18030
rect 19970 18010 19990 18030
rect 19990 18010 19995 18030
rect 19965 18005 19995 18010
rect 20045 18030 20075 18035
rect 20045 18010 20050 18030
rect 20050 18010 20070 18030
rect 20070 18010 20075 18030
rect 20045 18005 20075 18010
rect 20125 18030 20155 18035
rect 20125 18010 20130 18030
rect 20130 18010 20150 18030
rect 20150 18010 20155 18030
rect 20125 18005 20155 18010
rect 20205 18030 20235 18035
rect 20205 18010 20210 18030
rect 20210 18010 20230 18030
rect 20230 18010 20235 18030
rect 20205 18005 20235 18010
rect 20285 18030 20315 18035
rect 20285 18010 20290 18030
rect 20290 18010 20310 18030
rect 20310 18010 20315 18030
rect 20285 18005 20315 18010
rect 20365 18030 20395 18035
rect 20365 18010 20370 18030
rect 20370 18010 20390 18030
rect 20390 18010 20395 18030
rect 20365 18005 20395 18010
rect 20445 18030 20475 18035
rect 20445 18010 20450 18030
rect 20450 18010 20470 18030
rect 20470 18010 20475 18030
rect 20445 18005 20475 18010
rect 20525 18030 20555 18035
rect 20525 18010 20530 18030
rect 20530 18010 20550 18030
rect 20550 18010 20555 18030
rect 20525 18005 20555 18010
rect 20605 18030 20635 18035
rect 20605 18010 20610 18030
rect 20610 18010 20630 18030
rect 20630 18010 20635 18030
rect 20605 18005 20635 18010
rect 20685 18030 20715 18035
rect 20685 18010 20690 18030
rect 20690 18010 20710 18030
rect 20710 18010 20715 18030
rect 20685 18005 20715 18010
rect 20765 18030 20795 18035
rect 20765 18010 20770 18030
rect 20770 18010 20790 18030
rect 20790 18010 20795 18030
rect 20765 18005 20795 18010
rect 20845 18030 20875 18035
rect 20845 18010 20850 18030
rect 20850 18010 20870 18030
rect 20870 18010 20875 18030
rect 20845 18005 20875 18010
rect 20925 18030 20955 18035
rect 20925 18010 20930 18030
rect 20930 18010 20950 18030
rect 20950 18010 20955 18030
rect 20925 18005 20955 18010
rect 5 17870 35 17875
rect 5 17850 10 17870
rect 10 17850 30 17870
rect 30 17850 35 17870
rect 5 17845 35 17850
rect 85 17870 115 17875
rect 85 17850 90 17870
rect 90 17850 110 17870
rect 110 17850 115 17870
rect 85 17845 115 17850
rect 165 17870 195 17875
rect 165 17850 170 17870
rect 170 17850 190 17870
rect 190 17850 195 17870
rect 165 17845 195 17850
rect 245 17870 275 17875
rect 245 17850 250 17870
rect 250 17850 270 17870
rect 270 17850 275 17870
rect 245 17845 275 17850
rect 325 17870 355 17875
rect 325 17850 330 17870
rect 330 17850 350 17870
rect 350 17850 355 17870
rect 325 17845 355 17850
rect 405 17870 435 17875
rect 405 17850 410 17870
rect 410 17850 430 17870
rect 430 17850 435 17870
rect 405 17845 435 17850
rect 485 17870 515 17875
rect 485 17850 490 17870
rect 490 17850 510 17870
rect 510 17850 515 17870
rect 485 17845 515 17850
rect 565 17870 595 17875
rect 565 17850 570 17870
rect 570 17850 590 17870
rect 590 17850 595 17870
rect 565 17845 595 17850
rect 645 17870 675 17875
rect 645 17850 650 17870
rect 650 17850 670 17870
rect 670 17850 675 17870
rect 645 17845 675 17850
rect 725 17870 755 17875
rect 725 17850 730 17870
rect 730 17850 750 17870
rect 750 17850 755 17870
rect 725 17845 755 17850
rect 805 17870 835 17875
rect 805 17850 810 17870
rect 810 17850 830 17870
rect 830 17850 835 17870
rect 805 17845 835 17850
rect 885 17870 915 17875
rect 885 17850 890 17870
rect 890 17850 910 17870
rect 910 17850 915 17870
rect 885 17845 915 17850
rect 965 17870 995 17875
rect 965 17850 970 17870
rect 970 17850 990 17870
rect 990 17850 995 17870
rect 965 17845 995 17850
rect 1045 17870 1075 17875
rect 1045 17850 1050 17870
rect 1050 17850 1070 17870
rect 1070 17850 1075 17870
rect 1045 17845 1075 17850
rect 1125 17870 1155 17875
rect 1125 17850 1130 17870
rect 1130 17850 1150 17870
rect 1150 17850 1155 17870
rect 1125 17845 1155 17850
rect 1205 17870 1235 17875
rect 1205 17850 1210 17870
rect 1210 17850 1230 17870
rect 1230 17850 1235 17870
rect 1205 17845 1235 17850
rect 1285 17870 1315 17875
rect 1285 17850 1290 17870
rect 1290 17850 1310 17870
rect 1310 17850 1315 17870
rect 1285 17845 1315 17850
rect 1365 17870 1395 17875
rect 1365 17850 1370 17870
rect 1370 17850 1390 17870
rect 1390 17850 1395 17870
rect 1365 17845 1395 17850
rect 1445 17870 1475 17875
rect 1445 17850 1450 17870
rect 1450 17850 1470 17870
rect 1470 17850 1475 17870
rect 1445 17845 1475 17850
rect 1525 17870 1555 17875
rect 1525 17850 1530 17870
rect 1530 17850 1550 17870
rect 1550 17850 1555 17870
rect 1525 17845 1555 17850
rect 1605 17870 1635 17875
rect 1605 17850 1610 17870
rect 1610 17850 1630 17870
rect 1630 17850 1635 17870
rect 1605 17845 1635 17850
rect 1685 17870 1715 17875
rect 1685 17850 1690 17870
rect 1690 17850 1710 17870
rect 1710 17850 1715 17870
rect 1685 17845 1715 17850
rect 1765 17870 1795 17875
rect 1765 17850 1770 17870
rect 1770 17850 1790 17870
rect 1790 17850 1795 17870
rect 1765 17845 1795 17850
rect 1845 17870 1875 17875
rect 1845 17850 1850 17870
rect 1850 17850 1870 17870
rect 1870 17850 1875 17870
rect 1845 17845 1875 17850
rect 1925 17870 1955 17875
rect 1925 17850 1930 17870
rect 1930 17850 1950 17870
rect 1950 17850 1955 17870
rect 1925 17845 1955 17850
rect 2005 17870 2035 17875
rect 2005 17850 2010 17870
rect 2010 17850 2030 17870
rect 2030 17850 2035 17870
rect 2005 17845 2035 17850
rect 2085 17870 2115 17875
rect 2085 17850 2090 17870
rect 2090 17850 2110 17870
rect 2110 17850 2115 17870
rect 2085 17845 2115 17850
rect 2165 17870 2195 17875
rect 2165 17850 2170 17870
rect 2170 17850 2190 17870
rect 2190 17850 2195 17870
rect 2165 17845 2195 17850
rect 2245 17870 2275 17875
rect 2245 17850 2250 17870
rect 2250 17850 2270 17870
rect 2270 17850 2275 17870
rect 2245 17845 2275 17850
rect 2325 17870 2355 17875
rect 2325 17850 2330 17870
rect 2330 17850 2350 17870
rect 2350 17850 2355 17870
rect 2325 17845 2355 17850
rect 2405 17870 2435 17875
rect 2405 17850 2410 17870
rect 2410 17850 2430 17870
rect 2430 17850 2435 17870
rect 2405 17845 2435 17850
rect 2485 17870 2515 17875
rect 2485 17850 2490 17870
rect 2490 17850 2510 17870
rect 2510 17850 2515 17870
rect 2485 17845 2515 17850
rect 2565 17870 2595 17875
rect 2565 17850 2570 17870
rect 2570 17850 2590 17870
rect 2590 17850 2595 17870
rect 2565 17845 2595 17850
rect 2645 17870 2675 17875
rect 2645 17850 2650 17870
rect 2650 17850 2670 17870
rect 2670 17850 2675 17870
rect 2645 17845 2675 17850
rect 2725 17870 2755 17875
rect 2725 17850 2730 17870
rect 2730 17850 2750 17870
rect 2750 17850 2755 17870
rect 2725 17845 2755 17850
rect 2805 17870 2835 17875
rect 2805 17850 2810 17870
rect 2810 17850 2830 17870
rect 2830 17850 2835 17870
rect 2805 17845 2835 17850
rect 2885 17870 2915 17875
rect 2885 17850 2890 17870
rect 2890 17850 2910 17870
rect 2910 17850 2915 17870
rect 2885 17845 2915 17850
rect 2965 17870 2995 17875
rect 2965 17850 2970 17870
rect 2970 17850 2990 17870
rect 2990 17850 2995 17870
rect 2965 17845 2995 17850
rect 3045 17870 3075 17875
rect 3045 17850 3050 17870
rect 3050 17850 3070 17870
rect 3070 17850 3075 17870
rect 3045 17845 3075 17850
rect 3125 17870 3155 17875
rect 3125 17850 3130 17870
rect 3130 17850 3150 17870
rect 3150 17850 3155 17870
rect 3125 17845 3155 17850
rect 3205 17870 3235 17875
rect 3205 17850 3210 17870
rect 3210 17850 3230 17870
rect 3230 17850 3235 17870
rect 3205 17845 3235 17850
rect 3285 17870 3315 17875
rect 3285 17850 3290 17870
rect 3290 17850 3310 17870
rect 3310 17850 3315 17870
rect 3285 17845 3315 17850
rect 3365 17870 3395 17875
rect 3365 17850 3370 17870
rect 3370 17850 3390 17870
rect 3390 17850 3395 17870
rect 3365 17845 3395 17850
rect 3445 17870 3475 17875
rect 3445 17850 3450 17870
rect 3450 17850 3470 17870
rect 3470 17850 3475 17870
rect 3445 17845 3475 17850
rect 3525 17870 3555 17875
rect 3525 17850 3530 17870
rect 3530 17850 3550 17870
rect 3550 17850 3555 17870
rect 3525 17845 3555 17850
rect 3605 17870 3635 17875
rect 3605 17850 3610 17870
rect 3610 17850 3630 17870
rect 3630 17850 3635 17870
rect 3605 17845 3635 17850
rect 3685 17870 3715 17875
rect 3685 17850 3690 17870
rect 3690 17850 3710 17870
rect 3710 17850 3715 17870
rect 3685 17845 3715 17850
rect 3765 17870 3795 17875
rect 3765 17850 3770 17870
rect 3770 17850 3790 17870
rect 3790 17850 3795 17870
rect 3765 17845 3795 17850
rect 3845 17870 3875 17875
rect 3845 17850 3850 17870
rect 3850 17850 3870 17870
rect 3870 17850 3875 17870
rect 3845 17845 3875 17850
rect 3925 17870 3955 17875
rect 3925 17850 3930 17870
rect 3930 17850 3950 17870
rect 3950 17850 3955 17870
rect 3925 17845 3955 17850
rect 4005 17870 4035 17875
rect 4005 17850 4010 17870
rect 4010 17850 4030 17870
rect 4030 17850 4035 17870
rect 4005 17845 4035 17850
rect 4085 17870 4115 17875
rect 4085 17850 4090 17870
rect 4090 17850 4110 17870
rect 4110 17850 4115 17870
rect 4085 17845 4115 17850
rect 4165 17870 4195 17875
rect 4165 17850 4170 17870
rect 4170 17850 4190 17870
rect 4190 17850 4195 17870
rect 4165 17845 4195 17850
rect 6245 17870 6275 17875
rect 6245 17850 6250 17870
rect 6250 17850 6270 17870
rect 6270 17850 6275 17870
rect 6245 17845 6275 17850
rect 6325 17870 6355 17875
rect 6325 17850 6330 17870
rect 6330 17850 6350 17870
rect 6350 17850 6355 17870
rect 6325 17845 6355 17850
rect 6405 17870 6435 17875
rect 6405 17850 6410 17870
rect 6410 17850 6430 17870
rect 6430 17850 6435 17870
rect 6405 17845 6435 17850
rect 6485 17870 6515 17875
rect 6485 17850 6490 17870
rect 6490 17850 6510 17870
rect 6510 17850 6515 17870
rect 6485 17845 6515 17850
rect 6565 17870 6595 17875
rect 6565 17850 6570 17870
rect 6570 17850 6590 17870
rect 6590 17850 6595 17870
rect 6565 17845 6595 17850
rect 6645 17870 6675 17875
rect 6645 17850 6650 17870
rect 6650 17850 6670 17870
rect 6670 17850 6675 17870
rect 6645 17845 6675 17850
rect 6725 17870 6755 17875
rect 6725 17850 6730 17870
rect 6730 17850 6750 17870
rect 6750 17850 6755 17870
rect 6725 17845 6755 17850
rect 6805 17870 6835 17875
rect 6805 17850 6810 17870
rect 6810 17850 6830 17870
rect 6830 17850 6835 17870
rect 6805 17845 6835 17850
rect 6885 17870 6915 17875
rect 6885 17850 6890 17870
rect 6890 17850 6910 17870
rect 6910 17850 6915 17870
rect 6885 17845 6915 17850
rect 6965 17870 6995 17875
rect 6965 17850 6970 17870
rect 6970 17850 6990 17870
rect 6990 17850 6995 17870
rect 6965 17845 6995 17850
rect 7045 17870 7075 17875
rect 7045 17850 7050 17870
rect 7050 17850 7070 17870
rect 7070 17850 7075 17870
rect 7045 17845 7075 17850
rect 7125 17870 7155 17875
rect 7125 17850 7130 17870
rect 7130 17850 7150 17870
rect 7150 17850 7155 17870
rect 7125 17845 7155 17850
rect 7205 17870 7235 17875
rect 7205 17850 7210 17870
rect 7210 17850 7230 17870
rect 7230 17850 7235 17870
rect 7205 17845 7235 17850
rect 7285 17870 7315 17875
rect 7285 17850 7290 17870
rect 7290 17850 7310 17870
rect 7310 17850 7315 17870
rect 7285 17845 7315 17850
rect 7365 17870 7395 17875
rect 7365 17850 7370 17870
rect 7370 17850 7390 17870
rect 7390 17850 7395 17870
rect 7365 17845 7395 17850
rect 7445 17870 7475 17875
rect 7445 17850 7450 17870
rect 7450 17850 7470 17870
rect 7470 17850 7475 17870
rect 7445 17845 7475 17850
rect 7525 17870 7555 17875
rect 7525 17850 7530 17870
rect 7530 17850 7550 17870
rect 7550 17850 7555 17870
rect 7525 17845 7555 17850
rect 7605 17870 7635 17875
rect 7605 17850 7610 17870
rect 7610 17850 7630 17870
rect 7630 17850 7635 17870
rect 7605 17845 7635 17850
rect 7685 17870 7715 17875
rect 7685 17850 7690 17870
rect 7690 17850 7710 17870
rect 7710 17850 7715 17870
rect 7685 17845 7715 17850
rect 7765 17870 7795 17875
rect 7765 17850 7770 17870
rect 7770 17850 7790 17870
rect 7790 17850 7795 17870
rect 7765 17845 7795 17850
rect 7845 17870 7875 17875
rect 7845 17850 7850 17870
rect 7850 17850 7870 17870
rect 7870 17850 7875 17870
rect 7845 17845 7875 17850
rect 7925 17870 7955 17875
rect 7925 17850 7930 17870
rect 7930 17850 7950 17870
rect 7950 17850 7955 17870
rect 7925 17845 7955 17850
rect 8005 17870 8035 17875
rect 8005 17850 8010 17870
rect 8010 17850 8030 17870
rect 8030 17850 8035 17870
rect 8005 17845 8035 17850
rect 8085 17870 8115 17875
rect 8085 17850 8090 17870
rect 8090 17850 8110 17870
rect 8110 17850 8115 17870
rect 8085 17845 8115 17850
rect 8165 17870 8195 17875
rect 8165 17850 8170 17870
rect 8170 17850 8190 17870
rect 8190 17850 8195 17870
rect 8165 17845 8195 17850
rect 8245 17870 8275 17875
rect 8245 17850 8250 17870
rect 8250 17850 8270 17870
rect 8270 17850 8275 17870
rect 8245 17845 8275 17850
rect 8325 17870 8355 17875
rect 8325 17850 8330 17870
rect 8330 17850 8350 17870
rect 8350 17850 8355 17870
rect 8325 17845 8355 17850
rect 8405 17870 8435 17875
rect 8405 17850 8410 17870
rect 8410 17850 8430 17870
rect 8430 17850 8435 17870
rect 8405 17845 8435 17850
rect 8485 17870 8515 17875
rect 8485 17850 8490 17870
rect 8490 17850 8510 17870
rect 8510 17850 8515 17870
rect 8485 17845 8515 17850
rect 8565 17870 8595 17875
rect 8565 17850 8570 17870
rect 8570 17850 8590 17870
rect 8590 17850 8595 17870
rect 8565 17845 8595 17850
rect 8645 17870 8675 17875
rect 8645 17850 8650 17870
rect 8650 17850 8670 17870
rect 8670 17850 8675 17870
rect 8645 17845 8675 17850
rect 8725 17870 8755 17875
rect 8725 17850 8730 17870
rect 8730 17850 8750 17870
rect 8750 17850 8755 17870
rect 8725 17845 8755 17850
rect 8805 17870 8835 17875
rect 8805 17850 8810 17870
rect 8810 17850 8830 17870
rect 8830 17850 8835 17870
rect 8805 17845 8835 17850
rect 8885 17870 8915 17875
rect 8885 17850 8890 17870
rect 8890 17850 8910 17870
rect 8910 17850 8915 17870
rect 8885 17845 8915 17850
rect 8965 17870 8995 17875
rect 8965 17850 8970 17870
rect 8970 17850 8990 17870
rect 8990 17850 8995 17870
rect 8965 17845 8995 17850
rect 9045 17870 9075 17875
rect 9045 17850 9050 17870
rect 9050 17850 9070 17870
rect 9070 17850 9075 17870
rect 9045 17845 9075 17850
rect 9125 17870 9155 17875
rect 9125 17850 9130 17870
rect 9130 17850 9150 17870
rect 9150 17850 9155 17870
rect 9125 17845 9155 17850
rect 9205 17870 9235 17875
rect 9205 17850 9210 17870
rect 9210 17850 9230 17870
rect 9230 17850 9235 17870
rect 9205 17845 9235 17850
rect 9285 17870 9315 17875
rect 9285 17850 9290 17870
rect 9290 17850 9310 17870
rect 9310 17850 9315 17870
rect 9285 17845 9315 17850
rect 9365 17870 9395 17875
rect 9365 17850 9370 17870
rect 9370 17850 9390 17870
rect 9390 17850 9395 17870
rect 9365 17845 9395 17850
rect 9445 17870 9475 17875
rect 9445 17850 9450 17870
rect 9450 17850 9470 17870
rect 9470 17850 9475 17870
rect 9445 17845 9475 17850
rect 11565 17870 11595 17875
rect 11565 17850 11570 17870
rect 11570 17850 11590 17870
rect 11590 17850 11595 17870
rect 11565 17845 11595 17850
rect 11645 17870 11675 17875
rect 11645 17850 11650 17870
rect 11650 17850 11670 17870
rect 11670 17850 11675 17870
rect 11645 17845 11675 17850
rect 11725 17870 11755 17875
rect 11725 17850 11730 17870
rect 11730 17850 11750 17870
rect 11750 17850 11755 17870
rect 11725 17845 11755 17850
rect 11805 17870 11835 17875
rect 11805 17850 11810 17870
rect 11810 17850 11830 17870
rect 11830 17850 11835 17870
rect 11805 17845 11835 17850
rect 11885 17870 11915 17875
rect 11885 17850 11890 17870
rect 11890 17850 11910 17870
rect 11910 17850 11915 17870
rect 11885 17845 11915 17850
rect 11965 17870 11995 17875
rect 11965 17850 11970 17870
rect 11970 17850 11990 17870
rect 11990 17850 11995 17870
rect 11965 17845 11995 17850
rect 12045 17870 12075 17875
rect 12045 17850 12050 17870
rect 12050 17850 12070 17870
rect 12070 17850 12075 17870
rect 12045 17845 12075 17850
rect 12125 17870 12155 17875
rect 12125 17850 12130 17870
rect 12130 17850 12150 17870
rect 12150 17850 12155 17870
rect 12125 17845 12155 17850
rect 12205 17870 12235 17875
rect 12205 17850 12210 17870
rect 12210 17850 12230 17870
rect 12230 17850 12235 17870
rect 12205 17845 12235 17850
rect 12285 17870 12315 17875
rect 12285 17850 12290 17870
rect 12290 17850 12310 17870
rect 12310 17850 12315 17870
rect 12285 17845 12315 17850
rect 12365 17870 12395 17875
rect 12365 17850 12370 17870
rect 12370 17850 12390 17870
rect 12390 17850 12395 17870
rect 12365 17845 12395 17850
rect 12445 17870 12475 17875
rect 12445 17850 12450 17870
rect 12450 17850 12470 17870
rect 12470 17850 12475 17870
rect 12445 17845 12475 17850
rect 12525 17870 12555 17875
rect 12525 17850 12530 17870
rect 12530 17850 12550 17870
rect 12550 17850 12555 17870
rect 12525 17845 12555 17850
rect 12605 17870 12635 17875
rect 12605 17850 12610 17870
rect 12610 17850 12630 17870
rect 12630 17850 12635 17870
rect 12605 17845 12635 17850
rect 12685 17870 12715 17875
rect 12685 17850 12690 17870
rect 12690 17850 12710 17870
rect 12710 17850 12715 17870
rect 12685 17845 12715 17850
rect 12765 17870 12795 17875
rect 12765 17850 12770 17870
rect 12770 17850 12790 17870
rect 12790 17850 12795 17870
rect 12765 17845 12795 17850
rect 12845 17870 12875 17875
rect 12845 17850 12850 17870
rect 12850 17850 12870 17870
rect 12870 17850 12875 17870
rect 12845 17845 12875 17850
rect 12925 17870 12955 17875
rect 12925 17850 12930 17870
rect 12930 17850 12950 17870
rect 12950 17850 12955 17870
rect 12925 17845 12955 17850
rect 13005 17870 13035 17875
rect 13005 17850 13010 17870
rect 13010 17850 13030 17870
rect 13030 17850 13035 17870
rect 13005 17845 13035 17850
rect 13085 17870 13115 17875
rect 13085 17850 13090 17870
rect 13090 17850 13110 17870
rect 13110 17850 13115 17870
rect 13085 17845 13115 17850
rect 13165 17870 13195 17875
rect 13165 17850 13170 17870
rect 13170 17850 13190 17870
rect 13190 17850 13195 17870
rect 13165 17845 13195 17850
rect 13245 17870 13275 17875
rect 13245 17850 13250 17870
rect 13250 17850 13270 17870
rect 13270 17850 13275 17870
rect 13245 17845 13275 17850
rect 13325 17870 13355 17875
rect 13325 17850 13330 17870
rect 13330 17850 13350 17870
rect 13350 17850 13355 17870
rect 13325 17845 13355 17850
rect 13405 17870 13435 17875
rect 13405 17850 13410 17870
rect 13410 17850 13430 17870
rect 13430 17850 13435 17870
rect 13405 17845 13435 17850
rect 13485 17870 13515 17875
rect 13485 17850 13490 17870
rect 13490 17850 13510 17870
rect 13510 17850 13515 17870
rect 13485 17845 13515 17850
rect 13565 17870 13595 17875
rect 13565 17850 13570 17870
rect 13570 17850 13590 17870
rect 13590 17850 13595 17870
rect 13565 17845 13595 17850
rect 13645 17870 13675 17875
rect 13645 17850 13650 17870
rect 13650 17850 13670 17870
rect 13670 17850 13675 17870
rect 13645 17845 13675 17850
rect 13725 17870 13755 17875
rect 13725 17850 13730 17870
rect 13730 17850 13750 17870
rect 13750 17850 13755 17870
rect 13725 17845 13755 17850
rect 13805 17870 13835 17875
rect 13805 17850 13810 17870
rect 13810 17850 13830 17870
rect 13830 17850 13835 17870
rect 13805 17845 13835 17850
rect 13885 17870 13915 17875
rect 13885 17850 13890 17870
rect 13890 17850 13910 17870
rect 13910 17850 13915 17870
rect 13885 17845 13915 17850
rect 13965 17870 13995 17875
rect 13965 17850 13970 17870
rect 13970 17850 13990 17870
rect 13990 17850 13995 17870
rect 13965 17845 13995 17850
rect 14045 17870 14075 17875
rect 14045 17850 14050 17870
rect 14050 17850 14070 17870
rect 14070 17850 14075 17870
rect 14045 17845 14075 17850
rect 14125 17870 14155 17875
rect 14125 17850 14130 17870
rect 14130 17850 14150 17870
rect 14150 17850 14155 17870
rect 14125 17845 14155 17850
rect 14205 17870 14235 17875
rect 14205 17850 14210 17870
rect 14210 17850 14230 17870
rect 14230 17850 14235 17870
rect 14205 17845 14235 17850
rect 14285 17870 14315 17875
rect 14285 17850 14290 17870
rect 14290 17850 14310 17870
rect 14310 17850 14315 17870
rect 14285 17845 14315 17850
rect 14365 17870 14395 17875
rect 14365 17850 14370 17870
rect 14370 17850 14390 17870
rect 14390 17850 14395 17870
rect 14365 17845 14395 17850
rect 14445 17870 14475 17875
rect 14445 17850 14450 17870
rect 14450 17850 14470 17870
rect 14470 17850 14475 17870
rect 14445 17845 14475 17850
rect 14525 17870 14555 17875
rect 14525 17850 14530 17870
rect 14530 17850 14550 17870
rect 14550 17850 14555 17870
rect 14525 17845 14555 17850
rect 14605 17870 14635 17875
rect 14605 17850 14610 17870
rect 14610 17850 14630 17870
rect 14630 17850 14635 17870
rect 14605 17845 14635 17850
rect 14685 17870 14715 17875
rect 14685 17850 14690 17870
rect 14690 17850 14710 17870
rect 14710 17850 14715 17870
rect 14685 17845 14715 17850
rect 16765 17870 16795 17875
rect 16765 17850 16770 17870
rect 16770 17850 16790 17870
rect 16790 17850 16795 17870
rect 16765 17845 16795 17850
rect 16845 17870 16875 17875
rect 16845 17850 16850 17870
rect 16850 17850 16870 17870
rect 16870 17850 16875 17870
rect 16845 17845 16875 17850
rect 16925 17870 16955 17875
rect 16925 17850 16930 17870
rect 16930 17850 16950 17870
rect 16950 17850 16955 17870
rect 16925 17845 16955 17850
rect 17005 17870 17035 17875
rect 17005 17850 17010 17870
rect 17010 17850 17030 17870
rect 17030 17850 17035 17870
rect 17005 17845 17035 17850
rect 17085 17870 17115 17875
rect 17085 17850 17090 17870
rect 17090 17850 17110 17870
rect 17110 17850 17115 17870
rect 17085 17845 17115 17850
rect 17165 17870 17195 17875
rect 17165 17850 17170 17870
rect 17170 17850 17190 17870
rect 17190 17850 17195 17870
rect 17165 17845 17195 17850
rect 17245 17870 17275 17875
rect 17245 17850 17250 17870
rect 17250 17850 17270 17870
rect 17270 17850 17275 17870
rect 17245 17845 17275 17850
rect 17325 17870 17355 17875
rect 17325 17850 17330 17870
rect 17330 17850 17350 17870
rect 17350 17850 17355 17870
rect 17325 17845 17355 17850
rect 17405 17870 17435 17875
rect 17405 17850 17410 17870
rect 17410 17850 17430 17870
rect 17430 17850 17435 17870
rect 17405 17845 17435 17850
rect 17485 17870 17515 17875
rect 17485 17850 17490 17870
rect 17490 17850 17510 17870
rect 17510 17850 17515 17870
rect 17485 17845 17515 17850
rect 17565 17870 17595 17875
rect 17565 17850 17570 17870
rect 17570 17850 17590 17870
rect 17590 17850 17595 17870
rect 17565 17845 17595 17850
rect 17645 17870 17675 17875
rect 17645 17850 17650 17870
rect 17650 17850 17670 17870
rect 17670 17850 17675 17870
rect 17645 17845 17675 17850
rect 17725 17870 17755 17875
rect 17725 17850 17730 17870
rect 17730 17850 17750 17870
rect 17750 17850 17755 17870
rect 17725 17845 17755 17850
rect 17805 17870 17835 17875
rect 17805 17850 17810 17870
rect 17810 17850 17830 17870
rect 17830 17850 17835 17870
rect 17805 17845 17835 17850
rect 17885 17870 17915 17875
rect 17885 17850 17890 17870
rect 17890 17850 17910 17870
rect 17910 17850 17915 17870
rect 17885 17845 17915 17850
rect 17965 17870 17995 17875
rect 17965 17850 17970 17870
rect 17970 17850 17990 17870
rect 17990 17850 17995 17870
rect 17965 17845 17995 17850
rect 18045 17870 18075 17875
rect 18045 17850 18050 17870
rect 18050 17850 18070 17870
rect 18070 17850 18075 17870
rect 18045 17845 18075 17850
rect 18125 17870 18155 17875
rect 18125 17850 18130 17870
rect 18130 17850 18150 17870
rect 18150 17850 18155 17870
rect 18125 17845 18155 17850
rect 18205 17870 18235 17875
rect 18205 17850 18210 17870
rect 18210 17850 18230 17870
rect 18230 17850 18235 17870
rect 18205 17845 18235 17850
rect 18285 17870 18315 17875
rect 18285 17850 18290 17870
rect 18290 17850 18310 17870
rect 18310 17850 18315 17870
rect 18285 17845 18315 17850
rect 18365 17870 18395 17875
rect 18365 17850 18370 17870
rect 18370 17850 18390 17870
rect 18390 17850 18395 17870
rect 18365 17845 18395 17850
rect 18445 17870 18475 17875
rect 18445 17850 18450 17870
rect 18450 17850 18470 17870
rect 18470 17850 18475 17870
rect 18445 17845 18475 17850
rect 18525 17870 18555 17875
rect 18525 17850 18530 17870
rect 18530 17850 18550 17870
rect 18550 17850 18555 17870
rect 18525 17845 18555 17850
rect 18605 17870 18635 17875
rect 18605 17850 18610 17870
rect 18610 17850 18630 17870
rect 18630 17850 18635 17870
rect 18605 17845 18635 17850
rect 18685 17870 18715 17875
rect 18685 17850 18690 17870
rect 18690 17850 18710 17870
rect 18710 17850 18715 17870
rect 18685 17845 18715 17850
rect 18765 17870 18795 17875
rect 18765 17850 18770 17870
rect 18770 17850 18790 17870
rect 18790 17850 18795 17870
rect 18765 17845 18795 17850
rect 18845 17870 18875 17875
rect 18845 17850 18850 17870
rect 18850 17850 18870 17870
rect 18870 17850 18875 17870
rect 18845 17845 18875 17850
rect 18925 17870 18955 17875
rect 18925 17850 18930 17870
rect 18930 17850 18950 17870
rect 18950 17850 18955 17870
rect 18925 17845 18955 17850
rect 19005 17870 19035 17875
rect 19005 17850 19010 17870
rect 19010 17850 19030 17870
rect 19030 17850 19035 17870
rect 19005 17845 19035 17850
rect 19085 17870 19115 17875
rect 19085 17850 19090 17870
rect 19090 17850 19110 17870
rect 19110 17850 19115 17870
rect 19085 17845 19115 17850
rect 19165 17870 19195 17875
rect 19165 17850 19170 17870
rect 19170 17850 19190 17870
rect 19190 17850 19195 17870
rect 19165 17845 19195 17850
rect 19245 17870 19275 17875
rect 19245 17850 19250 17870
rect 19250 17850 19270 17870
rect 19270 17850 19275 17870
rect 19245 17845 19275 17850
rect 19325 17870 19355 17875
rect 19325 17850 19330 17870
rect 19330 17850 19350 17870
rect 19350 17850 19355 17870
rect 19325 17845 19355 17850
rect 19405 17870 19435 17875
rect 19405 17850 19410 17870
rect 19410 17850 19430 17870
rect 19430 17850 19435 17870
rect 19405 17845 19435 17850
rect 19485 17870 19515 17875
rect 19485 17850 19490 17870
rect 19490 17850 19510 17870
rect 19510 17850 19515 17870
rect 19485 17845 19515 17850
rect 19565 17870 19595 17875
rect 19565 17850 19570 17870
rect 19570 17850 19590 17870
rect 19590 17850 19595 17870
rect 19565 17845 19595 17850
rect 19645 17870 19675 17875
rect 19645 17850 19650 17870
rect 19650 17850 19670 17870
rect 19670 17850 19675 17870
rect 19645 17845 19675 17850
rect 19725 17870 19755 17875
rect 19725 17850 19730 17870
rect 19730 17850 19750 17870
rect 19750 17850 19755 17870
rect 19725 17845 19755 17850
rect 19805 17870 19835 17875
rect 19805 17850 19810 17870
rect 19810 17850 19830 17870
rect 19830 17850 19835 17870
rect 19805 17845 19835 17850
rect 19885 17870 19915 17875
rect 19885 17850 19890 17870
rect 19890 17850 19910 17870
rect 19910 17850 19915 17870
rect 19885 17845 19915 17850
rect 19965 17870 19995 17875
rect 19965 17850 19970 17870
rect 19970 17850 19990 17870
rect 19990 17850 19995 17870
rect 19965 17845 19995 17850
rect 20045 17870 20075 17875
rect 20045 17850 20050 17870
rect 20050 17850 20070 17870
rect 20070 17850 20075 17870
rect 20045 17845 20075 17850
rect 20125 17870 20155 17875
rect 20125 17850 20130 17870
rect 20130 17850 20150 17870
rect 20150 17850 20155 17870
rect 20125 17845 20155 17850
rect 20205 17870 20235 17875
rect 20205 17850 20210 17870
rect 20210 17850 20230 17870
rect 20230 17850 20235 17870
rect 20205 17845 20235 17850
rect 20285 17870 20315 17875
rect 20285 17850 20290 17870
rect 20290 17850 20310 17870
rect 20310 17850 20315 17870
rect 20285 17845 20315 17850
rect 20365 17870 20395 17875
rect 20365 17850 20370 17870
rect 20370 17850 20390 17870
rect 20390 17850 20395 17870
rect 20365 17845 20395 17850
rect 20445 17870 20475 17875
rect 20445 17850 20450 17870
rect 20450 17850 20470 17870
rect 20470 17850 20475 17870
rect 20445 17845 20475 17850
rect 20525 17870 20555 17875
rect 20525 17850 20530 17870
rect 20530 17850 20550 17870
rect 20550 17850 20555 17870
rect 20525 17845 20555 17850
rect 20605 17870 20635 17875
rect 20605 17850 20610 17870
rect 20610 17850 20630 17870
rect 20630 17850 20635 17870
rect 20605 17845 20635 17850
rect 20685 17870 20715 17875
rect 20685 17850 20690 17870
rect 20690 17850 20710 17870
rect 20710 17850 20715 17870
rect 20685 17845 20715 17850
rect 20765 17870 20795 17875
rect 20765 17850 20770 17870
rect 20770 17850 20790 17870
rect 20790 17850 20795 17870
rect 20765 17845 20795 17850
rect 20845 17870 20875 17875
rect 20845 17850 20850 17870
rect 20850 17850 20870 17870
rect 20870 17850 20875 17870
rect 20845 17845 20875 17850
rect 20925 17870 20955 17875
rect 20925 17850 20930 17870
rect 20930 17850 20950 17870
rect 20950 17850 20955 17870
rect 20925 17845 20955 17850
rect 5 17710 35 17715
rect 5 17690 10 17710
rect 10 17690 30 17710
rect 30 17690 35 17710
rect 5 17685 35 17690
rect 85 17710 115 17715
rect 85 17690 90 17710
rect 90 17690 110 17710
rect 110 17690 115 17710
rect 85 17685 115 17690
rect 165 17710 195 17715
rect 165 17690 170 17710
rect 170 17690 190 17710
rect 190 17690 195 17710
rect 165 17685 195 17690
rect 245 17710 275 17715
rect 245 17690 250 17710
rect 250 17690 270 17710
rect 270 17690 275 17710
rect 245 17685 275 17690
rect 325 17710 355 17715
rect 325 17690 330 17710
rect 330 17690 350 17710
rect 350 17690 355 17710
rect 325 17685 355 17690
rect 405 17710 435 17715
rect 405 17690 410 17710
rect 410 17690 430 17710
rect 430 17690 435 17710
rect 405 17685 435 17690
rect 485 17710 515 17715
rect 485 17690 490 17710
rect 490 17690 510 17710
rect 510 17690 515 17710
rect 485 17685 515 17690
rect 565 17710 595 17715
rect 565 17690 570 17710
rect 570 17690 590 17710
rect 590 17690 595 17710
rect 565 17685 595 17690
rect 645 17710 675 17715
rect 645 17690 650 17710
rect 650 17690 670 17710
rect 670 17690 675 17710
rect 645 17685 675 17690
rect 725 17710 755 17715
rect 725 17690 730 17710
rect 730 17690 750 17710
rect 750 17690 755 17710
rect 725 17685 755 17690
rect 805 17710 835 17715
rect 805 17690 810 17710
rect 810 17690 830 17710
rect 830 17690 835 17710
rect 805 17685 835 17690
rect 885 17710 915 17715
rect 885 17690 890 17710
rect 890 17690 910 17710
rect 910 17690 915 17710
rect 885 17685 915 17690
rect 965 17710 995 17715
rect 965 17690 970 17710
rect 970 17690 990 17710
rect 990 17690 995 17710
rect 965 17685 995 17690
rect 1045 17710 1075 17715
rect 1045 17690 1050 17710
rect 1050 17690 1070 17710
rect 1070 17690 1075 17710
rect 1045 17685 1075 17690
rect 1125 17710 1155 17715
rect 1125 17690 1130 17710
rect 1130 17690 1150 17710
rect 1150 17690 1155 17710
rect 1125 17685 1155 17690
rect 1205 17710 1235 17715
rect 1205 17690 1210 17710
rect 1210 17690 1230 17710
rect 1230 17690 1235 17710
rect 1205 17685 1235 17690
rect 1285 17710 1315 17715
rect 1285 17690 1290 17710
rect 1290 17690 1310 17710
rect 1310 17690 1315 17710
rect 1285 17685 1315 17690
rect 1365 17710 1395 17715
rect 1365 17690 1370 17710
rect 1370 17690 1390 17710
rect 1390 17690 1395 17710
rect 1365 17685 1395 17690
rect 1445 17710 1475 17715
rect 1445 17690 1450 17710
rect 1450 17690 1470 17710
rect 1470 17690 1475 17710
rect 1445 17685 1475 17690
rect 1525 17710 1555 17715
rect 1525 17690 1530 17710
rect 1530 17690 1550 17710
rect 1550 17690 1555 17710
rect 1525 17685 1555 17690
rect 1605 17710 1635 17715
rect 1605 17690 1610 17710
rect 1610 17690 1630 17710
rect 1630 17690 1635 17710
rect 1605 17685 1635 17690
rect 1685 17710 1715 17715
rect 1685 17690 1690 17710
rect 1690 17690 1710 17710
rect 1710 17690 1715 17710
rect 1685 17685 1715 17690
rect 1765 17710 1795 17715
rect 1765 17690 1770 17710
rect 1770 17690 1790 17710
rect 1790 17690 1795 17710
rect 1765 17685 1795 17690
rect 1845 17710 1875 17715
rect 1845 17690 1850 17710
rect 1850 17690 1870 17710
rect 1870 17690 1875 17710
rect 1845 17685 1875 17690
rect 1925 17710 1955 17715
rect 1925 17690 1930 17710
rect 1930 17690 1950 17710
rect 1950 17690 1955 17710
rect 1925 17685 1955 17690
rect 2005 17710 2035 17715
rect 2005 17690 2010 17710
rect 2010 17690 2030 17710
rect 2030 17690 2035 17710
rect 2005 17685 2035 17690
rect 2085 17710 2115 17715
rect 2085 17690 2090 17710
rect 2090 17690 2110 17710
rect 2110 17690 2115 17710
rect 2085 17685 2115 17690
rect 2165 17710 2195 17715
rect 2165 17690 2170 17710
rect 2170 17690 2190 17710
rect 2190 17690 2195 17710
rect 2165 17685 2195 17690
rect 2245 17710 2275 17715
rect 2245 17690 2250 17710
rect 2250 17690 2270 17710
rect 2270 17690 2275 17710
rect 2245 17685 2275 17690
rect 2325 17710 2355 17715
rect 2325 17690 2330 17710
rect 2330 17690 2350 17710
rect 2350 17690 2355 17710
rect 2325 17685 2355 17690
rect 2405 17710 2435 17715
rect 2405 17690 2410 17710
rect 2410 17690 2430 17710
rect 2430 17690 2435 17710
rect 2405 17685 2435 17690
rect 2485 17710 2515 17715
rect 2485 17690 2490 17710
rect 2490 17690 2510 17710
rect 2510 17690 2515 17710
rect 2485 17685 2515 17690
rect 2565 17710 2595 17715
rect 2565 17690 2570 17710
rect 2570 17690 2590 17710
rect 2590 17690 2595 17710
rect 2565 17685 2595 17690
rect 2645 17710 2675 17715
rect 2645 17690 2650 17710
rect 2650 17690 2670 17710
rect 2670 17690 2675 17710
rect 2645 17685 2675 17690
rect 2725 17710 2755 17715
rect 2725 17690 2730 17710
rect 2730 17690 2750 17710
rect 2750 17690 2755 17710
rect 2725 17685 2755 17690
rect 2805 17710 2835 17715
rect 2805 17690 2810 17710
rect 2810 17690 2830 17710
rect 2830 17690 2835 17710
rect 2805 17685 2835 17690
rect 2885 17710 2915 17715
rect 2885 17690 2890 17710
rect 2890 17690 2910 17710
rect 2910 17690 2915 17710
rect 2885 17685 2915 17690
rect 2965 17710 2995 17715
rect 2965 17690 2970 17710
rect 2970 17690 2990 17710
rect 2990 17690 2995 17710
rect 2965 17685 2995 17690
rect 3045 17710 3075 17715
rect 3045 17690 3050 17710
rect 3050 17690 3070 17710
rect 3070 17690 3075 17710
rect 3045 17685 3075 17690
rect 3125 17710 3155 17715
rect 3125 17690 3130 17710
rect 3130 17690 3150 17710
rect 3150 17690 3155 17710
rect 3125 17685 3155 17690
rect 3205 17710 3235 17715
rect 3205 17690 3210 17710
rect 3210 17690 3230 17710
rect 3230 17690 3235 17710
rect 3205 17685 3235 17690
rect 3285 17710 3315 17715
rect 3285 17690 3290 17710
rect 3290 17690 3310 17710
rect 3310 17690 3315 17710
rect 3285 17685 3315 17690
rect 3365 17710 3395 17715
rect 3365 17690 3370 17710
rect 3370 17690 3390 17710
rect 3390 17690 3395 17710
rect 3365 17685 3395 17690
rect 3445 17710 3475 17715
rect 3445 17690 3450 17710
rect 3450 17690 3470 17710
rect 3470 17690 3475 17710
rect 3445 17685 3475 17690
rect 3525 17710 3555 17715
rect 3525 17690 3530 17710
rect 3530 17690 3550 17710
rect 3550 17690 3555 17710
rect 3525 17685 3555 17690
rect 3605 17710 3635 17715
rect 3605 17690 3610 17710
rect 3610 17690 3630 17710
rect 3630 17690 3635 17710
rect 3605 17685 3635 17690
rect 3685 17710 3715 17715
rect 3685 17690 3690 17710
rect 3690 17690 3710 17710
rect 3710 17690 3715 17710
rect 3685 17685 3715 17690
rect 3765 17710 3795 17715
rect 3765 17690 3770 17710
rect 3770 17690 3790 17710
rect 3790 17690 3795 17710
rect 3765 17685 3795 17690
rect 3845 17710 3875 17715
rect 3845 17690 3850 17710
rect 3850 17690 3870 17710
rect 3870 17690 3875 17710
rect 3845 17685 3875 17690
rect 3925 17710 3955 17715
rect 3925 17690 3930 17710
rect 3930 17690 3950 17710
rect 3950 17690 3955 17710
rect 3925 17685 3955 17690
rect 4005 17710 4035 17715
rect 4005 17690 4010 17710
rect 4010 17690 4030 17710
rect 4030 17690 4035 17710
rect 4005 17685 4035 17690
rect 4085 17710 4115 17715
rect 4085 17690 4090 17710
rect 4090 17690 4110 17710
rect 4110 17690 4115 17710
rect 4085 17685 4115 17690
rect 4165 17710 4195 17715
rect 4165 17690 4170 17710
rect 4170 17690 4190 17710
rect 4190 17690 4195 17710
rect 4165 17685 4195 17690
rect 6245 17710 6275 17715
rect 6245 17690 6250 17710
rect 6250 17690 6270 17710
rect 6270 17690 6275 17710
rect 6245 17685 6275 17690
rect 6325 17710 6355 17715
rect 6325 17690 6330 17710
rect 6330 17690 6350 17710
rect 6350 17690 6355 17710
rect 6325 17685 6355 17690
rect 6405 17710 6435 17715
rect 6405 17690 6410 17710
rect 6410 17690 6430 17710
rect 6430 17690 6435 17710
rect 6405 17685 6435 17690
rect 6485 17710 6515 17715
rect 6485 17690 6490 17710
rect 6490 17690 6510 17710
rect 6510 17690 6515 17710
rect 6485 17685 6515 17690
rect 6565 17710 6595 17715
rect 6565 17690 6570 17710
rect 6570 17690 6590 17710
rect 6590 17690 6595 17710
rect 6565 17685 6595 17690
rect 6645 17710 6675 17715
rect 6645 17690 6650 17710
rect 6650 17690 6670 17710
rect 6670 17690 6675 17710
rect 6645 17685 6675 17690
rect 6725 17710 6755 17715
rect 6725 17690 6730 17710
rect 6730 17690 6750 17710
rect 6750 17690 6755 17710
rect 6725 17685 6755 17690
rect 6805 17710 6835 17715
rect 6805 17690 6810 17710
rect 6810 17690 6830 17710
rect 6830 17690 6835 17710
rect 6805 17685 6835 17690
rect 6885 17710 6915 17715
rect 6885 17690 6890 17710
rect 6890 17690 6910 17710
rect 6910 17690 6915 17710
rect 6885 17685 6915 17690
rect 6965 17710 6995 17715
rect 6965 17690 6970 17710
rect 6970 17690 6990 17710
rect 6990 17690 6995 17710
rect 6965 17685 6995 17690
rect 7045 17710 7075 17715
rect 7045 17690 7050 17710
rect 7050 17690 7070 17710
rect 7070 17690 7075 17710
rect 7045 17685 7075 17690
rect 7125 17710 7155 17715
rect 7125 17690 7130 17710
rect 7130 17690 7150 17710
rect 7150 17690 7155 17710
rect 7125 17685 7155 17690
rect 7205 17710 7235 17715
rect 7205 17690 7210 17710
rect 7210 17690 7230 17710
rect 7230 17690 7235 17710
rect 7205 17685 7235 17690
rect 7285 17710 7315 17715
rect 7285 17690 7290 17710
rect 7290 17690 7310 17710
rect 7310 17690 7315 17710
rect 7285 17685 7315 17690
rect 7365 17710 7395 17715
rect 7365 17690 7370 17710
rect 7370 17690 7390 17710
rect 7390 17690 7395 17710
rect 7365 17685 7395 17690
rect 7445 17710 7475 17715
rect 7445 17690 7450 17710
rect 7450 17690 7470 17710
rect 7470 17690 7475 17710
rect 7445 17685 7475 17690
rect 7525 17710 7555 17715
rect 7525 17690 7530 17710
rect 7530 17690 7550 17710
rect 7550 17690 7555 17710
rect 7525 17685 7555 17690
rect 7605 17710 7635 17715
rect 7605 17690 7610 17710
rect 7610 17690 7630 17710
rect 7630 17690 7635 17710
rect 7605 17685 7635 17690
rect 7685 17710 7715 17715
rect 7685 17690 7690 17710
rect 7690 17690 7710 17710
rect 7710 17690 7715 17710
rect 7685 17685 7715 17690
rect 7765 17710 7795 17715
rect 7765 17690 7770 17710
rect 7770 17690 7790 17710
rect 7790 17690 7795 17710
rect 7765 17685 7795 17690
rect 7845 17710 7875 17715
rect 7845 17690 7850 17710
rect 7850 17690 7870 17710
rect 7870 17690 7875 17710
rect 7845 17685 7875 17690
rect 7925 17710 7955 17715
rect 7925 17690 7930 17710
rect 7930 17690 7950 17710
rect 7950 17690 7955 17710
rect 7925 17685 7955 17690
rect 8005 17710 8035 17715
rect 8005 17690 8010 17710
rect 8010 17690 8030 17710
rect 8030 17690 8035 17710
rect 8005 17685 8035 17690
rect 8085 17710 8115 17715
rect 8085 17690 8090 17710
rect 8090 17690 8110 17710
rect 8110 17690 8115 17710
rect 8085 17685 8115 17690
rect 8165 17710 8195 17715
rect 8165 17690 8170 17710
rect 8170 17690 8190 17710
rect 8190 17690 8195 17710
rect 8165 17685 8195 17690
rect 8245 17710 8275 17715
rect 8245 17690 8250 17710
rect 8250 17690 8270 17710
rect 8270 17690 8275 17710
rect 8245 17685 8275 17690
rect 8325 17710 8355 17715
rect 8325 17690 8330 17710
rect 8330 17690 8350 17710
rect 8350 17690 8355 17710
rect 8325 17685 8355 17690
rect 8405 17710 8435 17715
rect 8405 17690 8410 17710
rect 8410 17690 8430 17710
rect 8430 17690 8435 17710
rect 8405 17685 8435 17690
rect 8485 17710 8515 17715
rect 8485 17690 8490 17710
rect 8490 17690 8510 17710
rect 8510 17690 8515 17710
rect 8485 17685 8515 17690
rect 8565 17710 8595 17715
rect 8565 17690 8570 17710
rect 8570 17690 8590 17710
rect 8590 17690 8595 17710
rect 8565 17685 8595 17690
rect 8645 17710 8675 17715
rect 8645 17690 8650 17710
rect 8650 17690 8670 17710
rect 8670 17690 8675 17710
rect 8645 17685 8675 17690
rect 8725 17710 8755 17715
rect 8725 17690 8730 17710
rect 8730 17690 8750 17710
rect 8750 17690 8755 17710
rect 8725 17685 8755 17690
rect 8805 17710 8835 17715
rect 8805 17690 8810 17710
rect 8810 17690 8830 17710
rect 8830 17690 8835 17710
rect 8805 17685 8835 17690
rect 8885 17710 8915 17715
rect 8885 17690 8890 17710
rect 8890 17690 8910 17710
rect 8910 17690 8915 17710
rect 8885 17685 8915 17690
rect 8965 17710 8995 17715
rect 8965 17690 8970 17710
rect 8970 17690 8990 17710
rect 8990 17690 8995 17710
rect 8965 17685 8995 17690
rect 9045 17710 9075 17715
rect 9045 17690 9050 17710
rect 9050 17690 9070 17710
rect 9070 17690 9075 17710
rect 9045 17685 9075 17690
rect 9125 17710 9155 17715
rect 9125 17690 9130 17710
rect 9130 17690 9150 17710
rect 9150 17690 9155 17710
rect 9125 17685 9155 17690
rect 9205 17710 9235 17715
rect 9205 17690 9210 17710
rect 9210 17690 9230 17710
rect 9230 17690 9235 17710
rect 9205 17685 9235 17690
rect 9285 17710 9315 17715
rect 9285 17690 9290 17710
rect 9290 17690 9310 17710
rect 9310 17690 9315 17710
rect 9285 17685 9315 17690
rect 9365 17710 9395 17715
rect 9365 17690 9370 17710
rect 9370 17690 9390 17710
rect 9390 17690 9395 17710
rect 9365 17685 9395 17690
rect 9445 17710 9475 17715
rect 9445 17690 9450 17710
rect 9450 17690 9470 17710
rect 9470 17690 9475 17710
rect 9445 17685 9475 17690
rect 11565 17710 11595 17715
rect 11565 17690 11570 17710
rect 11570 17690 11590 17710
rect 11590 17690 11595 17710
rect 11565 17685 11595 17690
rect 11645 17710 11675 17715
rect 11645 17690 11650 17710
rect 11650 17690 11670 17710
rect 11670 17690 11675 17710
rect 11645 17685 11675 17690
rect 11725 17710 11755 17715
rect 11725 17690 11730 17710
rect 11730 17690 11750 17710
rect 11750 17690 11755 17710
rect 11725 17685 11755 17690
rect 11805 17710 11835 17715
rect 11805 17690 11810 17710
rect 11810 17690 11830 17710
rect 11830 17690 11835 17710
rect 11805 17685 11835 17690
rect 11885 17710 11915 17715
rect 11885 17690 11890 17710
rect 11890 17690 11910 17710
rect 11910 17690 11915 17710
rect 11885 17685 11915 17690
rect 11965 17710 11995 17715
rect 11965 17690 11970 17710
rect 11970 17690 11990 17710
rect 11990 17690 11995 17710
rect 11965 17685 11995 17690
rect 12045 17710 12075 17715
rect 12045 17690 12050 17710
rect 12050 17690 12070 17710
rect 12070 17690 12075 17710
rect 12045 17685 12075 17690
rect 12125 17710 12155 17715
rect 12125 17690 12130 17710
rect 12130 17690 12150 17710
rect 12150 17690 12155 17710
rect 12125 17685 12155 17690
rect 12205 17710 12235 17715
rect 12205 17690 12210 17710
rect 12210 17690 12230 17710
rect 12230 17690 12235 17710
rect 12205 17685 12235 17690
rect 12285 17710 12315 17715
rect 12285 17690 12290 17710
rect 12290 17690 12310 17710
rect 12310 17690 12315 17710
rect 12285 17685 12315 17690
rect 12365 17710 12395 17715
rect 12365 17690 12370 17710
rect 12370 17690 12390 17710
rect 12390 17690 12395 17710
rect 12365 17685 12395 17690
rect 12445 17710 12475 17715
rect 12445 17690 12450 17710
rect 12450 17690 12470 17710
rect 12470 17690 12475 17710
rect 12445 17685 12475 17690
rect 12525 17710 12555 17715
rect 12525 17690 12530 17710
rect 12530 17690 12550 17710
rect 12550 17690 12555 17710
rect 12525 17685 12555 17690
rect 12605 17710 12635 17715
rect 12605 17690 12610 17710
rect 12610 17690 12630 17710
rect 12630 17690 12635 17710
rect 12605 17685 12635 17690
rect 12685 17710 12715 17715
rect 12685 17690 12690 17710
rect 12690 17690 12710 17710
rect 12710 17690 12715 17710
rect 12685 17685 12715 17690
rect 12765 17710 12795 17715
rect 12765 17690 12770 17710
rect 12770 17690 12790 17710
rect 12790 17690 12795 17710
rect 12765 17685 12795 17690
rect 12845 17710 12875 17715
rect 12845 17690 12850 17710
rect 12850 17690 12870 17710
rect 12870 17690 12875 17710
rect 12845 17685 12875 17690
rect 12925 17710 12955 17715
rect 12925 17690 12930 17710
rect 12930 17690 12950 17710
rect 12950 17690 12955 17710
rect 12925 17685 12955 17690
rect 13005 17710 13035 17715
rect 13005 17690 13010 17710
rect 13010 17690 13030 17710
rect 13030 17690 13035 17710
rect 13005 17685 13035 17690
rect 13085 17710 13115 17715
rect 13085 17690 13090 17710
rect 13090 17690 13110 17710
rect 13110 17690 13115 17710
rect 13085 17685 13115 17690
rect 13165 17710 13195 17715
rect 13165 17690 13170 17710
rect 13170 17690 13190 17710
rect 13190 17690 13195 17710
rect 13165 17685 13195 17690
rect 13245 17710 13275 17715
rect 13245 17690 13250 17710
rect 13250 17690 13270 17710
rect 13270 17690 13275 17710
rect 13245 17685 13275 17690
rect 13325 17710 13355 17715
rect 13325 17690 13330 17710
rect 13330 17690 13350 17710
rect 13350 17690 13355 17710
rect 13325 17685 13355 17690
rect 13405 17710 13435 17715
rect 13405 17690 13410 17710
rect 13410 17690 13430 17710
rect 13430 17690 13435 17710
rect 13405 17685 13435 17690
rect 13485 17710 13515 17715
rect 13485 17690 13490 17710
rect 13490 17690 13510 17710
rect 13510 17690 13515 17710
rect 13485 17685 13515 17690
rect 13565 17710 13595 17715
rect 13565 17690 13570 17710
rect 13570 17690 13590 17710
rect 13590 17690 13595 17710
rect 13565 17685 13595 17690
rect 13645 17710 13675 17715
rect 13645 17690 13650 17710
rect 13650 17690 13670 17710
rect 13670 17690 13675 17710
rect 13645 17685 13675 17690
rect 13725 17710 13755 17715
rect 13725 17690 13730 17710
rect 13730 17690 13750 17710
rect 13750 17690 13755 17710
rect 13725 17685 13755 17690
rect 13805 17710 13835 17715
rect 13805 17690 13810 17710
rect 13810 17690 13830 17710
rect 13830 17690 13835 17710
rect 13805 17685 13835 17690
rect 13885 17710 13915 17715
rect 13885 17690 13890 17710
rect 13890 17690 13910 17710
rect 13910 17690 13915 17710
rect 13885 17685 13915 17690
rect 13965 17710 13995 17715
rect 13965 17690 13970 17710
rect 13970 17690 13990 17710
rect 13990 17690 13995 17710
rect 13965 17685 13995 17690
rect 14045 17710 14075 17715
rect 14045 17690 14050 17710
rect 14050 17690 14070 17710
rect 14070 17690 14075 17710
rect 14045 17685 14075 17690
rect 14125 17710 14155 17715
rect 14125 17690 14130 17710
rect 14130 17690 14150 17710
rect 14150 17690 14155 17710
rect 14125 17685 14155 17690
rect 14205 17710 14235 17715
rect 14205 17690 14210 17710
rect 14210 17690 14230 17710
rect 14230 17690 14235 17710
rect 14205 17685 14235 17690
rect 14285 17710 14315 17715
rect 14285 17690 14290 17710
rect 14290 17690 14310 17710
rect 14310 17690 14315 17710
rect 14285 17685 14315 17690
rect 14365 17710 14395 17715
rect 14365 17690 14370 17710
rect 14370 17690 14390 17710
rect 14390 17690 14395 17710
rect 14365 17685 14395 17690
rect 14445 17710 14475 17715
rect 14445 17690 14450 17710
rect 14450 17690 14470 17710
rect 14470 17690 14475 17710
rect 14445 17685 14475 17690
rect 14525 17710 14555 17715
rect 14525 17690 14530 17710
rect 14530 17690 14550 17710
rect 14550 17690 14555 17710
rect 14525 17685 14555 17690
rect 14605 17710 14635 17715
rect 14605 17690 14610 17710
rect 14610 17690 14630 17710
rect 14630 17690 14635 17710
rect 14605 17685 14635 17690
rect 14685 17710 14715 17715
rect 14685 17690 14690 17710
rect 14690 17690 14710 17710
rect 14710 17690 14715 17710
rect 14685 17685 14715 17690
rect 16765 17710 16795 17715
rect 16765 17690 16770 17710
rect 16770 17690 16790 17710
rect 16790 17690 16795 17710
rect 16765 17685 16795 17690
rect 16845 17710 16875 17715
rect 16845 17690 16850 17710
rect 16850 17690 16870 17710
rect 16870 17690 16875 17710
rect 16845 17685 16875 17690
rect 16925 17710 16955 17715
rect 16925 17690 16930 17710
rect 16930 17690 16950 17710
rect 16950 17690 16955 17710
rect 16925 17685 16955 17690
rect 17005 17710 17035 17715
rect 17005 17690 17010 17710
rect 17010 17690 17030 17710
rect 17030 17690 17035 17710
rect 17005 17685 17035 17690
rect 17085 17710 17115 17715
rect 17085 17690 17090 17710
rect 17090 17690 17110 17710
rect 17110 17690 17115 17710
rect 17085 17685 17115 17690
rect 17165 17710 17195 17715
rect 17165 17690 17170 17710
rect 17170 17690 17190 17710
rect 17190 17690 17195 17710
rect 17165 17685 17195 17690
rect 17245 17710 17275 17715
rect 17245 17690 17250 17710
rect 17250 17690 17270 17710
rect 17270 17690 17275 17710
rect 17245 17685 17275 17690
rect 17325 17710 17355 17715
rect 17325 17690 17330 17710
rect 17330 17690 17350 17710
rect 17350 17690 17355 17710
rect 17325 17685 17355 17690
rect 17405 17710 17435 17715
rect 17405 17690 17410 17710
rect 17410 17690 17430 17710
rect 17430 17690 17435 17710
rect 17405 17685 17435 17690
rect 17485 17710 17515 17715
rect 17485 17690 17490 17710
rect 17490 17690 17510 17710
rect 17510 17690 17515 17710
rect 17485 17685 17515 17690
rect 17565 17710 17595 17715
rect 17565 17690 17570 17710
rect 17570 17690 17590 17710
rect 17590 17690 17595 17710
rect 17565 17685 17595 17690
rect 17645 17710 17675 17715
rect 17645 17690 17650 17710
rect 17650 17690 17670 17710
rect 17670 17690 17675 17710
rect 17645 17685 17675 17690
rect 17725 17710 17755 17715
rect 17725 17690 17730 17710
rect 17730 17690 17750 17710
rect 17750 17690 17755 17710
rect 17725 17685 17755 17690
rect 17805 17710 17835 17715
rect 17805 17690 17810 17710
rect 17810 17690 17830 17710
rect 17830 17690 17835 17710
rect 17805 17685 17835 17690
rect 17885 17710 17915 17715
rect 17885 17690 17890 17710
rect 17890 17690 17910 17710
rect 17910 17690 17915 17710
rect 17885 17685 17915 17690
rect 17965 17710 17995 17715
rect 17965 17690 17970 17710
rect 17970 17690 17990 17710
rect 17990 17690 17995 17710
rect 17965 17685 17995 17690
rect 18045 17710 18075 17715
rect 18045 17690 18050 17710
rect 18050 17690 18070 17710
rect 18070 17690 18075 17710
rect 18045 17685 18075 17690
rect 18125 17710 18155 17715
rect 18125 17690 18130 17710
rect 18130 17690 18150 17710
rect 18150 17690 18155 17710
rect 18125 17685 18155 17690
rect 18205 17710 18235 17715
rect 18205 17690 18210 17710
rect 18210 17690 18230 17710
rect 18230 17690 18235 17710
rect 18205 17685 18235 17690
rect 18285 17710 18315 17715
rect 18285 17690 18290 17710
rect 18290 17690 18310 17710
rect 18310 17690 18315 17710
rect 18285 17685 18315 17690
rect 18365 17710 18395 17715
rect 18365 17690 18370 17710
rect 18370 17690 18390 17710
rect 18390 17690 18395 17710
rect 18365 17685 18395 17690
rect 18445 17710 18475 17715
rect 18445 17690 18450 17710
rect 18450 17690 18470 17710
rect 18470 17690 18475 17710
rect 18445 17685 18475 17690
rect 18525 17710 18555 17715
rect 18525 17690 18530 17710
rect 18530 17690 18550 17710
rect 18550 17690 18555 17710
rect 18525 17685 18555 17690
rect 18605 17710 18635 17715
rect 18605 17690 18610 17710
rect 18610 17690 18630 17710
rect 18630 17690 18635 17710
rect 18605 17685 18635 17690
rect 18685 17710 18715 17715
rect 18685 17690 18690 17710
rect 18690 17690 18710 17710
rect 18710 17690 18715 17710
rect 18685 17685 18715 17690
rect 18765 17710 18795 17715
rect 18765 17690 18770 17710
rect 18770 17690 18790 17710
rect 18790 17690 18795 17710
rect 18765 17685 18795 17690
rect 18845 17710 18875 17715
rect 18845 17690 18850 17710
rect 18850 17690 18870 17710
rect 18870 17690 18875 17710
rect 18845 17685 18875 17690
rect 18925 17710 18955 17715
rect 18925 17690 18930 17710
rect 18930 17690 18950 17710
rect 18950 17690 18955 17710
rect 18925 17685 18955 17690
rect 19005 17710 19035 17715
rect 19005 17690 19010 17710
rect 19010 17690 19030 17710
rect 19030 17690 19035 17710
rect 19005 17685 19035 17690
rect 19085 17710 19115 17715
rect 19085 17690 19090 17710
rect 19090 17690 19110 17710
rect 19110 17690 19115 17710
rect 19085 17685 19115 17690
rect 19165 17710 19195 17715
rect 19165 17690 19170 17710
rect 19170 17690 19190 17710
rect 19190 17690 19195 17710
rect 19165 17685 19195 17690
rect 19245 17710 19275 17715
rect 19245 17690 19250 17710
rect 19250 17690 19270 17710
rect 19270 17690 19275 17710
rect 19245 17685 19275 17690
rect 19325 17710 19355 17715
rect 19325 17690 19330 17710
rect 19330 17690 19350 17710
rect 19350 17690 19355 17710
rect 19325 17685 19355 17690
rect 19405 17710 19435 17715
rect 19405 17690 19410 17710
rect 19410 17690 19430 17710
rect 19430 17690 19435 17710
rect 19405 17685 19435 17690
rect 19485 17710 19515 17715
rect 19485 17690 19490 17710
rect 19490 17690 19510 17710
rect 19510 17690 19515 17710
rect 19485 17685 19515 17690
rect 19565 17710 19595 17715
rect 19565 17690 19570 17710
rect 19570 17690 19590 17710
rect 19590 17690 19595 17710
rect 19565 17685 19595 17690
rect 19645 17710 19675 17715
rect 19645 17690 19650 17710
rect 19650 17690 19670 17710
rect 19670 17690 19675 17710
rect 19645 17685 19675 17690
rect 19725 17710 19755 17715
rect 19725 17690 19730 17710
rect 19730 17690 19750 17710
rect 19750 17690 19755 17710
rect 19725 17685 19755 17690
rect 19805 17710 19835 17715
rect 19805 17690 19810 17710
rect 19810 17690 19830 17710
rect 19830 17690 19835 17710
rect 19805 17685 19835 17690
rect 19885 17710 19915 17715
rect 19885 17690 19890 17710
rect 19890 17690 19910 17710
rect 19910 17690 19915 17710
rect 19885 17685 19915 17690
rect 19965 17710 19995 17715
rect 19965 17690 19970 17710
rect 19970 17690 19990 17710
rect 19990 17690 19995 17710
rect 19965 17685 19995 17690
rect 20045 17710 20075 17715
rect 20045 17690 20050 17710
rect 20050 17690 20070 17710
rect 20070 17690 20075 17710
rect 20045 17685 20075 17690
rect 20125 17710 20155 17715
rect 20125 17690 20130 17710
rect 20130 17690 20150 17710
rect 20150 17690 20155 17710
rect 20125 17685 20155 17690
rect 20205 17710 20235 17715
rect 20205 17690 20210 17710
rect 20210 17690 20230 17710
rect 20230 17690 20235 17710
rect 20205 17685 20235 17690
rect 20285 17710 20315 17715
rect 20285 17690 20290 17710
rect 20290 17690 20310 17710
rect 20310 17690 20315 17710
rect 20285 17685 20315 17690
rect 20365 17710 20395 17715
rect 20365 17690 20370 17710
rect 20370 17690 20390 17710
rect 20390 17690 20395 17710
rect 20365 17685 20395 17690
rect 20445 17710 20475 17715
rect 20445 17690 20450 17710
rect 20450 17690 20470 17710
rect 20470 17690 20475 17710
rect 20445 17685 20475 17690
rect 20525 17710 20555 17715
rect 20525 17690 20530 17710
rect 20530 17690 20550 17710
rect 20550 17690 20555 17710
rect 20525 17685 20555 17690
rect 20605 17710 20635 17715
rect 20605 17690 20610 17710
rect 20610 17690 20630 17710
rect 20630 17690 20635 17710
rect 20605 17685 20635 17690
rect 20685 17710 20715 17715
rect 20685 17690 20690 17710
rect 20690 17690 20710 17710
rect 20710 17690 20715 17710
rect 20685 17685 20715 17690
rect 20765 17710 20795 17715
rect 20765 17690 20770 17710
rect 20770 17690 20790 17710
rect 20790 17690 20795 17710
rect 20765 17685 20795 17690
rect 20845 17710 20875 17715
rect 20845 17690 20850 17710
rect 20850 17690 20870 17710
rect 20870 17690 20875 17710
rect 20845 17685 20875 17690
rect 20925 17710 20955 17715
rect 20925 17690 20930 17710
rect 20930 17690 20950 17710
rect 20950 17690 20955 17710
rect 20925 17685 20955 17690
rect 5 17550 35 17555
rect 5 17530 10 17550
rect 10 17530 30 17550
rect 30 17530 35 17550
rect 5 17525 35 17530
rect 85 17550 115 17555
rect 85 17530 90 17550
rect 90 17530 110 17550
rect 110 17530 115 17550
rect 85 17525 115 17530
rect 165 17550 195 17555
rect 165 17530 170 17550
rect 170 17530 190 17550
rect 190 17530 195 17550
rect 165 17525 195 17530
rect 245 17550 275 17555
rect 245 17530 250 17550
rect 250 17530 270 17550
rect 270 17530 275 17550
rect 245 17525 275 17530
rect 325 17550 355 17555
rect 325 17530 330 17550
rect 330 17530 350 17550
rect 350 17530 355 17550
rect 325 17525 355 17530
rect 405 17550 435 17555
rect 405 17530 410 17550
rect 410 17530 430 17550
rect 430 17530 435 17550
rect 405 17525 435 17530
rect 485 17550 515 17555
rect 485 17530 490 17550
rect 490 17530 510 17550
rect 510 17530 515 17550
rect 485 17525 515 17530
rect 565 17550 595 17555
rect 565 17530 570 17550
rect 570 17530 590 17550
rect 590 17530 595 17550
rect 565 17525 595 17530
rect 645 17550 675 17555
rect 645 17530 650 17550
rect 650 17530 670 17550
rect 670 17530 675 17550
rect 645 17525 675 17530
rect 725 17550 755 17555
rect 725 17530 730 17550
rect 730 17530 750 17550
rect 750 17530 755 17550
rect 725 17525 755 17530
rect 805 17550 835 17555
rect 805 17530 810 17550
rect 810 17530 830 17550
rect 830 17530 835 17550
rect 805 17525 835 17530
rect 885 17550 915 17555
rect 885 17530 890 17550
rect 890 17530 910 17550
rect 910 17530 915 17550
rect 885 17525 915 17530
rect 965 17550 995 17555
rect 965 17530 970 17550
rect 970 17530 990 17550
rect 990 17530 995 17550
rect 965 17525 995 17530
rect 1045 17550 1075 17555
rect 1045 17530 1050 17550
rect 1050 17530 1070 17550
rect 1070 17530 1075 17550
rect 1045 17525 1075 17530
rect 1125 17550 1155 17555
rect 1125 17530 1130 17550
rect 1130 17530 1150 17550
rect 1150 17530 1155 17550
rect 1125 17525 1155 17530
rect 1205 17550 1235 17555
rect 1205 17530 1210 17550
rect 1210 17530 1230 17550
rect 1230 17530 1235 17550
rect 1205 17525 1235 17530
rect 1285 17550 1315 17555
rect 1285 17530 1290 17550
rect 1290 17530 1310 17550
rect 1310 17530 1315 17550
rect 1285 17525 1315 17530
rect 1365 17550 1395 17555
rect 1365 17530 1370 17550
rect 1370 17530 1390 17550
rect 1390 17530 1395 17550
rect 1365 17525 1395 17530
rect 1445 17550 1475 17555
rect 1445 17530 1450 17550
rect 1450 17530 1470 17550
rect 1470 17530 1475 17550
rect 1445 17525 1475 17530
rect 1525 17550 1555 17555
rect 1525 17530 1530 17550
rect 1530 17530 1550 17550
rect 1550 17530 1555 17550
rect 1525 17525 1555 17530
rect 1605 17550 1635 17555
rect 1605 17530 1610 17550
rect 1610 17530 1630 17550
rect 1630 17530 1635 17550
rect 1605 17525 1635 17530
rect 1685 17550 1715 17555
rect 1685 17530 1690 17550
rect 1690 17530 1710 17550
rect 1710 17530 1715 17550
rect 1685 17525 1715 17530
rect 1765 17550 1795 17555
rect 1765 17530 1770 17550
rect 1770 17530 1790 17550
rect 1790 17530 1795 17550
rect 1765 17525 1795 17530
rect 1845 17550 1875 17555
rect 1845 17530 1850 17550
rect 1850 17530 1870 17550
rect 1870 17530 1875 17550
rect 1845 17525 1875 17530
rect 1925 17550 1955 17555
rect 1925 17530 1930 17550
rect 1930 17530 1950 17550
rect 1950 17530 1955 17550
rect 1925 17525 1955 17530
rect 2005 17550 2035 17555
rect 2005 17530 2010 17550
rect 2010 17530 2030 17550
rect 2030 17530 2035 17550
rect 2005 17525 2035 17530
rect 2085 17550 2115 17555
rect 2085 17530 2090 17550
rect 2090 17530 2110 17550
rect 2110 17530 2115 17550
rect 2085 17525 2115 17530
rect 2165 17550 2195 17555
rect 2165 17530 2170 17550
rect 2170 17530 2190 17550
rect 2190 17530 2195 17550
rect 2165 17525 2195 17530
rect 2245 17550 2275 17555
rect 2245 17530 2250 17550
rect 2250 17530 2270 17550
rect 2270 17530 2275 17550
rect 2245 17525 2275 17530
rect 2325 17550 2355 17555
rect 2325 17530 2330 17550
rect 2330 17530 2350 17550
rect 2350 17530 2355 17550
rect 2325 17525 2355 17530
rect 2405 17550 2435 17555
rect 2405 17530 2410 17550
rect 2410 17530 2430 17550
rect 2430 17530 2435 17550
rect 2405 17525 2435 17530
rect 2485 17550 2515 17555
rect 2485 17530 2490 17550
rect 2490 17530 2510 17550
rect 2510 17530 2515 17550
rect 2485 17525 2515 17530
rect 2565 17550 2595 17555
rect 2565 17530 2570 17550
rect 2570 17530 2590 17550
rect 2590 17530 2595 17550
rect 2565 17525 2595 17530
rect 2645 17550 2675 17555
rect 2645 17530 2650 17550
rect 2650 17530 2670 17550
rect 2670 17530 2675 17550
rect 2645 17525 2675 17530
rect 2725 17550 2755 17555
rect 2725 17530 2730 17550
rect 2730 17530 2750 17550
rect 2750 17530 2755 17550
rect 2725 17525 2755 17530
rect 2805 17550 2835 17555
rect 2805 17530 2810 17550
rect 2810 17530 2830 17550
rect 2830 17530 2835 17550
rect 2805 17525 2835 17530
rect 2885 17550 2915 17555
rect 2885 17530 2890 17550
rect 2890 17530 2910 17550
rect 2910 17530 2915 17550
rect 2885 17525 2915 17530
rect 2965 17550 2995 17555
rect 2965 17530 2970 17550
rect 2970 17530 2990 17550
rect 2990 17530 2995 17550
rect 2965 17525 2995 17530
rect 3045 17550 3075 17555
rect 3045 17530 3050 17550
rect 3050 17530 3070 17550
rect 3070 17530 3075 17550
rect 3045 17525 3075 17530
rect 3125 17550 3155 17555
rect 3125 17530 3130 17550
rect 3130 17530 3150 17550
rect 3150 17530 3155 17550
rect 3125 17525 3155 17530
rect 3205 17550 3235 17555
rect 3205 17530 3210 17550
rect 3210 17530 3230 17550
rect 3230 17530 3235 17550
rect 3205 17525 3235 17530
rect 3285 17550 3315 17555
rect 3285 17530 3290 17550
rect 3290 17530 3310 17550
rect 3310 17530 3315 17550
rect 3285 17525 3315 17530
rect 3365 17550 3395 17555
rect 3365 17530 3370 17550
rect 3370 17530 3390 17550
rect 3390 17530 3395 17550
rect 3365 17525 3395 17530
rect 3445 17550 3475 17555
rect 3445 17530 3450 17550
rect 3450 17530 3470 17550
rect 3470 17530 3475 17550
rect 3445 17525 3475 17530
rect 3525 17550 3555 17555
rect 3525 17530 3530 17550
rect 3530 17530 3550 17550
rect 3550 17530 3555 17550
rect 3525 17525 3555 17530
rect 3605 17550 3635 17555
rect 3605 17530 3610 17550
rect 3610 17530 3630 17550
rect 3630 17530 3635 17550
rect 3605 17525 3635 17530
rect 3685 17550 3715 17555
rect 3685 17530 3690 17550
rect 3690 17530 3710 17550
rect 3710 17530 3715 17550
rect 3685 17525 3715 17530
rect 3765 17550 3795 17555
rect 3765 17530 3770 17550
rect 3770 17530 3790 17550
rect 3790 17530 3795 17550
rect 3765 17525 3795 17530
rect 3845 17550 3875 17555
rect 3845 17530 3850 17550
rect 3850 17530 3870 17550
rect 3870 17530 3875 17550
rect 3845 17525 3875 17530
rect 3925 17550 3955 17555
rect 3925 17530 3930 17550
rect 3930 17530 3950 17550
rect 3950 17530 3955 17550
rect 3925 17525 3955 17530
rect 4005 17550 4035 17555
rect 4005 17530 4010 17550
rect 4010 17530 4030 17550
rect 4030 17530 4035 17550
rect 4005 17525 4035 17530
rect 4085 17550 4115 17555
rect 4085 17530 4090 17550
rect 4090 17530 4110 17550
rect 4110 17530 4115 17550
rect 4085 17525 4115 17530
rect 4165 17550 4195 17555
rect 4165 17530 4170 17550
rect 4170 17530 4190 17550
rect 4190 17530 4195 17550
rect 4165 17525 4195 17530
rect 6245 17550 6275 17555
rect 6245 17530 6250 17550
rect 6250 17530 6270 17550
rect 6270 17530 6275 17550
rect 6245 17525 6275 17530
rect 6325 17550 6355 17555
rect 6325 17530 6330 17550
rect 6330 17530 6350 17550
rect 6350 17530 6355 17550
rect 6325 17525 6355 17530
rect 6405 17550 6435 17555
rect 6405 17530 6410 17550
rect 6410 17530 6430 17550
rect 6430 17530 6435 17550
rect 6405 17525 6435 17530
rect 6485 17550 6515 17555
rect 6485 17530 6490 17550
rect 6490 17530 6510 17550
rect 6510 17530 6515 17550
rect 6485 17525 6515 17530
rect 6565 17550 6595 17555
rect 6565 17530 6570 17550
rect 6570 17530 6590 17550
rect 6590 17530 6595 17550
rect 6565 17525 6595 17530
rect 6645 17550 6675 17555
rect 6645 17530 6650 17550
rect 6650 17530 6670 17550
rect 6670 17530 6675 17550
rect 6645 17525 6675 17530
rect 6725 17550 6755 17555
rect 6725 17530 6730 17550
rect 6730 17530 6750 17550
rect 6750 17530 6755 17550
rect 6725 17525 6755 17530
rect 6805 17550 6835 17555
rect 6805 17530 6810 17550
rect 6810 17530 6830 17550
rect 6830 17530 6835 17550
rect 6805 17525 6835 17530
rect 6885 17550 6915 17555
rect 6885 17530 6890 17550
rect 6890 17530 6910 17550
rect 6910 17530 6915 17550
rect 6885 17525 6915 17530
rect 6965 17550 6995 17555
rect 6965 17530 6970 17550
rect 6970 17530 6990 17550
rect 6990 17530 6995 17550
rect 6965 17525 6995 17530
rect 7045 17550 7075 17555
rect 7045 17530 7050 17550
rect 7050 17530 7070 17550
rect 7070 17530 7075 17550
rect 7045 17525 7075 17530
rect 7125 17550 7155 17555
rect 7125 17530 7130 17550
rect 7130 17530 7150 17550
rect 7150 17530 7155 17550
rect 7125 17525 7155 17530
rect 7205 17550 7235 17555
rect 7205 17530 7210 17550
rect 7210 17530 7230 17550
rect 7230 17530 7235 17550
rect 7205 17525 7235 17530
rect 7285 17550 7315 17555
rect 7285 17530 7290 17550
rect 7290 17530 7310 17550
rect 7310 17530 7315 17550
rect 7285 17525 7315 17530
rect 7365 17550 7395 17555
rect 7365 17530 7370 17550
rect 7370 17530 7390 17550
rect 7390 17530 7395 17550
rect 7365 17525 7395 17530
rect 7445 17550 7475 17555
rect 7445 17530 7450 17550
rect 7450 17530 7470 17550
rect 7470 17530 7475 17550
rect 7445 17525 7475 17530
rect 7525 17550 7555 17555
rect 7525 17530 7530 17550
rect 7530 17530 7550 17550
rect 7550 17530 7555 17550
rect 7525 17525 7555 17530
rect 7605 17550 7635 17555
rect 7605 17530 7610 17550
rect 7610 17530 7630 17550
rect 7630 17530 7635 17550
rect 7605 17525 7635 17530
rect 7685 17550 7715 17555
rect 7685 17530 7690 17550
rect 7690 17530 7710 17550
rect 7710 17530 7715 17550
rect 7685 17525 7715 17530
rect 7765 17550 7795 17555
rect 7765 17530 7770 17550
rect 7770 17530 7790 17550
rect 7790 17530 7795 17550
rect 7765 17525 7795 17530
rect 7845 17550 7875 17555
rect 7845 17530 7850 17550
rect 7850 17530 7870 17550
rect 7870 17530 7875 17550
rect 7845 17525 7875 17530
rect 7925 17550 7955 17555
rect 7925 17530 7930 17550
rect 7930 17530 7950 17550
rect 7950 17530 7955 17550
rect 7925 17525 7955 17530
rect 8005 17550 8035 17555
rect 8005 17530 8010 17550
rect 8010 17530 8030 17550
rect 8030 17530 8035 17550
rect 8005 17525 8035 17530
rect 8085 17550 8115 17555
rect 8085 17530 8090 17550
rect 8090 17530 8110 17550
rect 8110 17530 8115 17550
rect 8085 17525 8115 17530
rect 8165 17550 8195 17555
rect 8165 17530 8170 17550
rect 8170 17530 8190 17550
rect 8190 17530 8195 17550
rect 8165 17525 8195 17530
rect 8245 17550 8275 17555
rect 8245 17530 8250 17550
rect 8250 17530 8270 17550
rect 8270 17530 8275 17550
rect 8245 17525 8275 17530
rect 8325 17550 8355 17555
rect 8325 17530 8330 17550
rect 8330 17530 8350 17550
rect 8350 17530 8355 17550
rect 8325 17525 8355 17530
rect 8405 17550 8435 17555
rect 8405 17530 8410 17550
rect 8410 17530 8430 17550
rect 8430 17530 8435 17550
rect 8405 17525 8435 17530
rect 8485 17550 8515 17555
rect 8485 17530 8490 17550
rect 8490 17530 8510 17550
rect 8510 17530 8515 17550
rect 8485 17525 8515 17530
rect 8565 17550 8595 17555
rect 8565 17530 8570 17550
rect 8570 17530 8590 17550
rect 8590 17530 8595 17550
rect 8565 17525 8595 17530
rect 8645 17550 8675 17555
rect 8645 17530 8650 17550
rect 8650 17530 8670 17550
rect 8670 17530 8675 17550
rect 8645 17525 8675 17530
rect 8725 17550 8755 17555
rect 8725 17530 8730 17550
rect 8730 17530 8750 17550
rect 8750 17530 8755 17550
rect 8725 17525 8755 17530
rect 8805 17550 8835 17555
rect 8805 17530 8810 17550
rect 8810 17530 8830 17550
rect 8830 17530 8835 17550
rect 8805 17525 8835 17530
rect 8885 17550 8915 17555
rect 8885 17530 8890 17550
rect 8890 17530 8910 17550
rect 8910 17530 8915 17550
rect 8885 17525 8915 17530
rect 8965 17550 8995 17555
rect 8965 17530 8970 17550
rect 8970 17530 8990 17550
rect 8990 17530 8995 17550
rect 8965 17525 8995 17530
rect 9045 17550 9075 17555
rect 9045 17530 9050 17550
rect 9050 17530 9070 17550
rect 9070 17530 9075 17550
rect 9045 17525 9075 17530
rect 9125 17550 9155 17555
rect 9125 17530 9130 17550
rect 9130 17530 9150 17550
rect 9150 17530 9155 17550
rect 9125 17525 9155 17530
rect 9205 17550 9235 17555
rect 9205 17530 9210 17550
rect 9210 17530 9230 17550
rect 9230 17530 9235 17550
rect 9205 17525 9235 17530
rect 9285 17550 9315 17555
rect 9285 17530 9290 17550
rect 9290 17530 9310 17550
rect 9310 17530 9315 17550
rect 9285 17525 9315 17530
rect 9365 17550 9395 17555
rect 9365 17530 9370 17550
rect 9370 17530 9390 17550
rect 9390 17530 9395 17550
rect 9365 17525 9395 17530
rect 9445 17550 9475 17555
rect 9445 17530 9450 17550
rect 9450 17530 9470 17550
rect 9470 17530 9475 17550
rect 9445 17525 9475 17530
rect 11565 17550 11595 17555
rect 11565 17530 11570 17550
rect 11570 17530 11590 17550
rect 11590 17530 11595 17550
rect 11565 17525 11595 17530
rect 11645 17550 11675 17555
rect 11645 17530 11650 17550
rect 11650 17530 11670 17550
rect 11670 17530 11675 17550
rect 11645 17525 11675 17530
rect 11725 17550 11755 17555
rect 11725 17530 11730 17550
rect 11730 17530 11750 17550
rect 11750 17530 11755 17550
rect 11725 17525 11755 17530
rect 11805 17550 11835 17555
rect 11805 17530 11810 17550
rect 11810 17530 11830 17550
rect 11830 17530 11835 17550
rect 11805 17525 11835 17530
rect 11885 17550 11915 17555
rect 11885 17530 11890 17550
rect 11890 17530 11910 17550
rect 11910 17530 11915 17550
rect 11885 17525 11915 17530
rect 11965 17550 11995 17555
rect 11965 17530 11970 17550
rect 11970 17530 11990 17550
rect 11990 17530 11995 17550
rect 11965 17525 11995 17530
rect 12045 17550 12075 17555
rect 12045 17530 12050 17550
rect 12050 17530 12070 17550
rect 12070 17530 12075 17550
rect 12045 17525 12075 17530
rect 12125 17550 12155 17555
rect 12125 17530 12130 17550
rect 12130 17530 12150 17550
rect 12150 17530 12155 17550
rect 12125 17525 12155 17530
rect 12205 17550 12235 17555
rect 12205 17530 12210 17550
rect 12210 17530 12230 17550
rect 12230 17530 12235 17550
rect 12205 17525 12235 17530
rect 12285 17550 12315 17555
rect 12285 17530 12290 17550
rect 12290 17530 12310 17550
rect 12310 17530 12315 17550
rect 12285 17525 12315 17530
rect 12365 17550 12395 17555
rect 12365 17530 12370 17550
rect 12370 17530 12390 17550
rect 12390 17530 12395 17550
rect 12365 17525 12395 17530
rect 12445 17550 12475 17555
rect 12445 17530 12450 17550
rect 12450 17530 12470 17550
rect 12470 17530 12475 17550
rect 12445 17525 12475 17530
rect 12525 17550 12555 17555
rect 12525 17530 12530 17550
rect 12530 17530 12550 17550
rect 12550 17530 12555 17550
rect 12525 17525 12555 17530
rect 12605 17550 12635 17555
rect 12605 17530 12610 17550
rect 12610 17530 12630 17550
rect 12630 17530 12635 17550
rect 12605 17525 12635 17530
rect 12685 17550 12715 17555
rect 12685 17530 12690 17550
rect 12690 17530 12710 17550
rect 12710 17530 12715 17550
rect 12685 17525 12715 17530
rect 12765 17550 12795 17555
rect 12765 17530 12770 17550
rect 12770 17530 12790 17550
rect 12790 17530 12795 17550
rect 12765 17525 12795 17530
rect 12845 17550 12875 17555
rect 12845 17530 12850 17550
rect 12850 17530 12870 17550
rect 12870 17530 12875 17550
rect 12845 17525 12875 17530
rect 12925 17550 12955 17555
rect 12925 17530 12930 17550
rect 12930 17530 12950 17550
rect 12950 17530 12955 17550
rect 12925 17525 12955 17530
rect 13005 17550 13035 17555
rect 13005 17530 13010 17550
rect 13010 17530 13030 17550
rect 13030 17530 13035 17550
rect 13005 17525 13035 17530
rect 13085 17550 13115 17555
rect 13085 17530 13090 17550
rect 13090 17530 13110 17550
rect 13110 17530 13115 17550
rect 13085 17525 13115 17530
rect 13165 17550 13195 17555
rect 13165 17530 13170 17550
rect 13170 17530 13190 17550
rect 13190 17530 13195 17550
rect 13165 17525 13195 17530
rect 13245 17550 13275 17555
rect 13245 17530 13250 17550
rect 13250 17530 13270 17550
rect 13270 17530 13275 17550
rect 13245 17525 13275 17530
rect 13325 17550 13355 17555
rect 13325 17530 13330 17550
rect 13330 17530 13350 17550
rect 13350 17530 13355 17550
rect 13325 17525 13355 17530
rect 13405 17550 13435 17555
rect 13405 17530 13410 17550
rect 13410 17530 13430 17550
rect 13430 17530 13435 17550
rect 13405 17525 13435 17530
rect 13485 17550 13515 17555
rect 13485 17530 13490 17550
rect 13490 17530 13510 17550
rect 13510 17530 13515 17550
rect 13485 17525 13515 17530
rect 13565 17550 13595 17555
rect 13565 17530 13570 17550
rect 13570 17530 13590 17550
rect 13590 17530 13595 17550
rect 13565 17525 13595 17530
rect 13645 17550 13675 17555
rect 13645 17530 13650 17550
rect 13650 17530 13670 17550
rect 13670 17530 13675 17550
rect 13645 17525 13675 17530
rect 13725 17550 13755 17555
rect 13725 17530 13730 17550
rect 13730 17530 13750 17550
rect 13750 17530 13755 17550
rect 13725 17525 13755 17530
rect 13805 17550 13835 17555
rect 13805 17530 13810 17550
rect 13810 17530 13830 17550
rect 13830 17530 13835 17550
rect 13805 17525 13835 17530
rect 13885 17550 13915 17555
rect 13885 17530 13890 17550
rect 13890 17530 13910 17550
rect 13910 17530 13915 17550
rect 13885 17525 13915 17530
rect 13965 17550 13995 17555
rect 13965 17530 13970 17550
rect 13970 17530 13990 17550
rect 13990 17530 13995 17550
rect 13965 17525 13995 17530
rect 14045 17550 14075 17555
rect 14045 17530 14050 17550
rect 14050 17530 14070 17550
rect 14070 17530 14075 17550
rect 14045 17525 14075 17530
rect 14125 17550 14155 17555
rect 14125 17530 14130 17550
rect 14130 17530 14150 17550
rect 14150 17530 14155 17550
rect 14125 17525 14155 17530
rect 14205 17550 14235 17555
rect 14205 17530 14210 17550
rect 14210 17530 14230 17550
rect 14230 17530 14235 17550
rect 14205 17525 14235 17530
rect 14285 17550 14315 17555
rect 14285 17530 14290 17550
rect 14290 17530 14310 17550
rect 14310 17530 14315 17550
rect 14285 17525 14315 17530
rect 14365 17550 14395 17555
rect 14365 17530 14370 17550
rect 14370 17530 14390 17550
rect 14390 17530 14395 17550
rect 14365 17525 14395 17530
rect 14445 17550 14475 17555
rect 14445 17530 14450 17550
rect 14450 17530 14470 17550
rect 14470 17530 14475 17550
rect 14445 17525 14475 17530
rect 14525 17550 14555 17555
rect 14525 17530 14530 17550
rect 14530 17530 14550 17550
rect 14550 17530 14555 17550
rect 14525 17525 14555 17530
rect 14605 17550 14635 17555
rect 14605 17530 14610 17550
rect 14610 17530 14630 17550
rect 14630 17530 14635 17550
rect 14605 17525 14635 17530
rect 14685 17550 14715 17555
rect 14685 17530 14690 17550
rect 14690 17530 14710 17550
rect 14710 17530 14715 17550
rect 14685 17525 14715 17530
rect 16765 17550 16795 17555
rect 16765 17530 16770 17550
rect 16770 17530 16790 17550
rect 16790 17530 16795 17550
rect 16765 17525 16795 17530
rect 16845 17550 16875 17555
rect 16845 17530 16850 17550
rect 16850 17530 16870 17550
rect 16870 17530 16875 17550
rect 16845 17525 16875 17530
rect 16925 17550 16955 17555
rect 16925 17530 16930 17550
rect 16930 17530 16950 17550
rect 16950 17530 16955 17550
rect 16925 17525 16955 17530
rect 17005 17550 17035 17555
rect 17005 17530 17010 17550
rect 17010 17530 17030 17550
rect 17030 17530 17035 17550
rect 17005 17525 17035 17530
rect 17085 17550 17115 17555
rect 17085 17530 17090 17550
rect 17090 17530 17110 17550
rect 17110 17530 17115 17550
rect 17085 17525 17115 17530
rect 17165 17550 17195 17555
rect 17165 17530 17170 17550
rect 17170 17530 17190 17550
rect 17190 17530 17195 17550
rect 17165 17525 17195 17530
rect 17245 17550 17275 17555
rect 17245 17530 17250 17550
rect 17250 17530 17270 17550
rect 17270 17530 17275 17550
rect 17245 17525 17275 17530
rect 17325 17550 17355 17555
rect 17325 17530 17330 17550
rect 17330 17530 17350 17550
rect 17350 17530 17355 17550
rect 17325 17525 17355 17530
rect 17405 17550 17435 17555
rect 17405 17530 17410 17550
rect 17410 17530 17430 17550
rect 17430 17530 17435 17550
rect 17405 17525 17435 17530
rect 17485 17550 17515 17555
rect 17485 17530 17490 17550
rect 17490 17530 17510 17550
rect 17510 17530 17515 17550
rect 17485 17525 17515 17530
rect 17565 17550 17595 17555
rect 17565 17530 17570 17550
rect 17570 17530 17590 17550
rect 17590 17530 17595 17550
rect 17565 17525 17595 17530
rect 17645 17550 17675 17555
rect 17645 17530 17650 17550
rect 17650 17530 17670 17550
rect 17670 17530 17675 17550
rect 17645 17525 17675 17530
rect 17725 17550 17755 17555
rect 17725 17530 17730 17550
rect 17730 17530 17750 17550
rect 17750 17530 17755 17550
rect 17725 17525 17755 17530
rect 17805 17550 17835 17555
rect 17805 17530 17810 17550
rect 17810 17530 17830 17550
rect 17830 17530 17835 17550
rect 17805 17525 17835 17530
rect 17885 17550 17915 17555
rect 17885 17530 17890 17550
rect 17890 17530 17910 17550
rect 17910 17530 17915 17550
rect 17885 17525 17915 17530
rect 17965 17550 17995 17555
rect 17965 17530 17970 17550
rect 17970 17530 17990 17550
rect 17990 17530 17995 17550
rect 17965 17525 17995 17530
rect 18045 17550 18075 17555
rect 18045 17530 18050 17550
rect 18050 17530 18070 17550
rect 18070 17530 18075 17550
rect 18045 17525 18075 17530
rect 18125 17550 18155 17555
rect 18125 17530 18130 17550
rect 18130 17530 18150 17550
rect 18150 17530 18155 17550
rect 18125 17525 18155 17530
rect 18205 17550 18235 17555
rect 18205 17530 18210 17550
rect 18210 17530 18230 17550
rect 18230 17530 18235 17550
rect 18205 17525 18235 17530
rect 18285 17550 18315 17555
rect 18285 17530 18290 17550
rect 18290 17530 18310 17550
rect 18310 17530 18315 17550
rect 18285 17525 18315 17530
rect 18365 17550 18395 17555
rect 18365 17530 18370 17550
rect 18370 17530 18390 17550
rect 18390 17530 18395 17550
rect 18365 17525 18395 17530
rect 18445 17550 18475 17555
rect 18445 17530 18450 17550
rect 18450 17530 18470 17550
rect 18470 17530 18475 17550
rect 18445 17525 18475 17530
rect 18525 17550 18555 17555
rect 18525 17530 18530 17550
rect 18530 17530 18550 17550
rect 18550 17530 18555 17550
rect 18525 17525 18555 17530
rect 18605 17550 18635 17555
rect 18605 17530 18610 17550
rect 18610 17530 18630 17550
rect 18630 17530 18635 17550
rect 18605 17525 18635 17530
rect 18685 17550 18715 17555
rect 18685 17530 18690 17550
rect 18690 17530 18710 17550
rect 18710 17530 18715 17550
rect 18685 17525 18715 17530
rect 18765 17550 18795 17555
rect 18765 17530 18770 17550
rect 18770 17530 18790 17550
rect 18790 17530 18795 17550
rect 18765 17525 18795 17530
rect 18845 17550 18875 17555
rect 18845 17530 18850 17550
rect 18850 17530 18870 17550
rect 18870 17530 18875 17550
rect 18845 17525 18875 17530
rect 18925 17550 18955 17555
rect 18925 17530 18930 17550
rect 18930 17530 18950 17550
rect 18950 17530 18955 17550
rect 18925 17525 18955 17530
rect 19005 17550 19035 17555
rect 19005 17530 19010 17550
rect 19010 17530 19030 17550
rect 19030 17530 19035 17550
rect 19005 17525 19035 17530
rect 19085 17550 19115 17555
rect 19085 17530 19090 17550
rect 19090 17530 19110 17550
rect 19110 17530 19115 17550
rect 19085 17525 19115 17530
rect 19165 17550 19195 17555
rect 19165 17530 19170 17550
rect 19170 17530 19190 17550
rect 19190 17530 19195 17550
rect 19165 17525 19195 17530
rect 19245 17550 19275 17555
rect 19245 17530 19250 17550
rect 19250 17530 19270 17550
rect 19270 17530 19275 17550
rect 19245 17525 19275 17530
rect 19325 17550 19355 17555
rect 19325 17530 19330 17550
rect 19330 17530 19350 17550
rect 19350 17530 19355 17550
rect 19325 17525 19355 17530
rect 19405 17550 19435 17555
rect 19405 17530 19410 17550
rect 19410 17530 19430 17550
rect 19430 17530 19435 17550
rect 19405 17525 19435 17530
rect 19485 17550 19515 17555
rect 19485 17530 19490 17550
rect 19490 17530 19510 17550
rect 19510 17530 19515 17550
rect 19485 17525 19515 17530
rect 19565 17550 19595 17555
rect 19565 17530 19570 17550
rect 19570 17530 19590 17550
rect 19590 17530 19595 17550
rect 19565 17525 19595 17530
rect 19645 17550 19675 17555
rect 19645 17530 19650 17550
rect 19650 17530 19670 17550
rect 19670 17530 19675 17550
rect 19645 17525 19675 17530
rect 19725 17550 19755 17555
rect 19725 17530 19730 17550
rect 19730 17530 19750 17550
rect 19750 17530 19755 17550
rect 19725 17525 19755 17530
rect 19805 17550 19835 17555
rect 19805 17530 19810 17550
rect 19810 17530 19830 17550
rect 19830 17530 19835 17550
rect 19805 17525 19835 17530
rect 19885 17550 19915 17555
rect 19885 17530 19890 17550
rect 19890 17530 19910 17550
rect 19910 17530 19915 17550
rect 19885 17525 19915 17530
rect 19965 17550 19995 17555
rect 19965 17530 19970 17550
rect 19970 17530 19990 17550
rect 19990 17530 19995 17550
rect 19965 17525 19995 17530
rect 20045 17550 20075 17555
rect 20045 17530 20050 17550
rect 20050 17530 20070 17550
rect 20070 17530 20075 17550
rect 20045 17525 20075 17530
rect 20125 17550 20155 17555
rect 20125 17530 20130 17550
rect 20130 17530 20150 17550
rect 20150 17530 20155 17550
rect 20125 17525 20155 17530
rect 20205 17550 20235 17555
rect 20205 17530 20210 17550
rect 20210 17530 20230 17550
rect 20230 17530 20235 17550
rect 20205 17525 20235 17530
rect 20285 17550 20315 17555
rect 20285 17530 20290 17550
rect 20290 17530 20310 17550
rect 20310 17530 20315 17550
rect 20285 17525 20315 17530
rect 20365 17550 20395 17555
rect 20365 17530 20370 17550
rect 20370 17530 20390 17550
rect 20390 17530 20395 17550
rect 20365 17525 20395 17530
rect 20445 17550 20475 17555
rect 20445 17530 20450 17550
rect 20450 17530 20470 17550
rect 20470 17530 20475 17550
rect 20445 17525 20475 17530
rect 20525 17550 20555 17555
rect 20525 17530 20530 17550
rect 20530 17530 20550 17550
rect 20550 17530 20555 17550
rect 20525 17525 20555 17530
rect 20605 17550 20635 17555
rect 20605 17530 20610 17550
rect 20610 17530 20630 17550
rect 20630 17530 20635 17550
rect 20605 17525 20635 17530
rect 20685 17550 20715 17555
rect 20685 17530 20690 17550
rect 20690 17530 20710 17550
rect 20710 17530 20715 17550
rect 20685 17525 20715 17530
rect 20765 17550 20795 17555
rect 20765 17530 20770 17550
rect 20770 17530 20790 17550
rect 20790 17530 20795 17550
rect 20765 17525 20795 17530
rect 20845 17550 20875 17555
rect 20845 17530 20850 17550
rect 20850 17530 20870 17550
rect 20870 17530 20875 17550
rect 20845 17525 20875 17530
rect 20925 17550 20955 17555
rect 20925 17530 20930 17550
rect 20930 17530 20950 17550
rect 20950 17530 20955 17550
rect 20925 17525 20955 17530
rect 5 17390 35 17395
rect 5 17370 10 17390
rect 10 17370 30 17390
rect 30 17370 35 17390
rect 5 17365 35 17370
rect 85 17390 115 17395
rect 85 17370 90 17390
rect 90 17370 110 17390
rect 110 17370 115 17390
rect 85 17365 115 17370
rect 165 17390 195 17395
rect 165 17370 170 17390
rect 170 17370 190 17390
rect 190 17370 195 17390
rect 165 17365 195 17370
rect 245 17390 275 17395
rect 245 17370 250 17390
rect 250 17370 270 17390
rect 270 17370 275 17390
rect 245 17365 275 17370
rect 325 17390 355 17395
rect 325 17370 330 17390
rect 330 17370 350 17390
rect 350 17370 355 17390
rect 325 17365 355 17370
rect 405 17390 435 17395
rect 405 17370 410 17390
rect 410 17370 430 17390
rect 430 17370 435 17390
rect 405 17365 435 17370
rect 485 17390 515 17395
rect 485 17370 490 17390
rect 490 17370 510 17390
rect 510 17370 515 17390
rect 485 17365 515 17370
rect 565 17390 595 17395
rect 565 17370 570 17390
rect 570 17370 590 17390
rect 590 17370 595 17390
rect 565 17365 595 17370
rect 645 17390 675 17395
rect 645 17370 650 17390
rect 650 17370 670 17390
rect 670 17370 675 17390
rect 645 17365 675 17370
rect 725 17390 755 17395
rect 725 17370 730 17390
rect 730 17370 750 17390
rect 750 17370 755 17390
rect 725 17365 755 17370
rect 805 17390 835 17395
rect 805 17370 810 17390
rect 810 17370 830 17390
rect 830 17370 835 17390
rect 805 17365 835 17370
rect 885 17390 915 17395
rect 885 17370 890 17390
rect 890 17370 910 17390
rect 910 17370 915 17390
rect 885 17365 915 17370
rect 965 17390 995 17395
rect 965 17370 970 17390
rect 970 17370 990 17390
rect 990 17370 995 17390
rect 965 17365 995 17370
rect 1045 17390 1075 17395
rect 1045 17370 1050 17390
rect 1050 17370 1070 17390
rect 1070 17370 1075 17390
rect 1045 17365 1075 17370
rect 1125 17390 1155 17395
rect 1125 17370 1130 17390
rect 1130 17370 1150 17390
rect 1150 17370 1155 17390
rect 1125 17365 1155 17370
rect 1205 17390 1235 17395
rect 1205 17370 1210 17390
rect 1210 17370 1230 17390
rect 1230 17370 1235 17390
rect 1205 17365 1235 17370
rect 1285 17390 1315 17395
rect 1285 17370 1290 17390
rect 1290 17370 1310 17390
rect 1310 17370 1315 17390
rect 1285 17365 1315 17370
rect 1365 17390 1395 17395
rect 1365 17370 1370 17390
rect 1370 17370 1390 17390
rect 1390 17370 1395 17390
rect 1365 17365 1395 17370
rect 1445 17390 1475 17395
rect 1445 17370 1450 17390
rect 1450 17370 1470 17390
rect 1470 17370 1475 17390
rect 1445 17365 1475 17370
rect 1525 17390 1555 17395
rect 1525 17370 1530 17390
rect 1530 17370 1550 17390
rect 1550 17370 1555 17390
rect 1525 17365 1555 17370
rect 1605 17390 1635 17395
rect 1605 17370 1610 17390
rect 1610 17370 1630 17390
rect 1630 17370 1635 17390
rect 1605 17365 1635 17370
rect 1685 17390 1715 17395
rect 1685 17370 1690 17390
rect 1690 17370 1710 17390
rect 1710 17370 1715 17390
rect 1685 17365 1715 17370
rect 1765 17390 1795 17395
rect 1765 17370 1770 17390
rect 1770 17370 1790 17390
rect 1790 17370 1795 17390
rect 1765 17365 1795 17370
rect 1845 17390 1875 17395
rect 1845 17370 1850 17390
rect 1850 17370 1870 17390
rect 1870 17370 1875 17390
rect 1845 17365 1875 17370
rect 1925 17390 1955 17395
rect 1925 17370 1930 17390
rect 1930 17370 1950 17390
rect 1950 17370 1955 17390
rect 1925 17365 1955 17370
rect 2005 17390 2035 17395
rect 2005 17370 2010 17390
rect 2010 17370 2030 17390
rect 2030 17370 2035 17390
rect 2005 17365 2035 17370
rect 2085 17390 2115 17395
rect 2085 17370 2090 17390
rect 2090 17370 2110 17390
rect 2110 17370 2115 17390
rect 2085 17365 2115 17370
rect 2165 17390 2195 17395
rect 2165 17370 2170 17390
rect 2170 17370 2190 17390
rect 2190 17370 2195 17390
rect 2165 17365 2195 17370
rect 2245 17390 2275 17395
rect 2245 17370 2250 17390
rect 2250 17370 2270 17390
rect 2270 17370 2275 17390
rect 2245 17365 2275 17370
rect 2325 17390 2355 17395
rect 2325 17370 2330 17390
rect 2330 17370 2350 17390
rect 2350 17370 2355 17390
rect 2325 17365 2355 17370
rect 2405 17390 2435 17395
rect 2405 17370 2410 17390
rect 2410 17370 2430 17390
rect 2430 17370 2435 17390
rect 2405 17365 2435 17370
rect 2485 17390 2515 17395
rect 2485 17370 2490 17390
rect 2490 17370 2510 17390
rect 2510 17370 2515 17390
rect 2485 17365 2515 17370
rect 2565 17390 2595 17395
rect 2565 17370 2570 17390
rect 2570 17370 2590 17390
rect 2590 17370 2595 17390
rect 2565 17365 2595 17370
rect 2645 17390 2675 17395
rect 2645 17370 2650 17390
rect 2650 17370 2670 17390
rect 2670 17370 2675 17390
rect 2645 17365 2675 17370
rect 2725 17390 2755 17395
rect 2725 17370 2730 17390
rect 2730 17370 2750 17390
rect 2750 17370 2755 17390
rect 2725 17365 2755 17370
rect 2805 17390 2835 17395
rect 2805 17370 2810 17390
rect 2810 17370 2830 17390
rect 2830 17370 2835 17390
rect 2805 17365 2835 17370
rect 2885 17390 2915 17395
rect 2885 17370 2890 17390
rect 2890 17370 2910 17390
rect 2910 17370 2915 17390
rect 2885 17365 2915 17370
rect 2965 17390 2995 17395
rect 2965 17370 2970 17390
rect 2970 17370 2990 17390
rect 2990 17370 2995 17390
rect 2965 17365 2995 17370
rect 3045 17390 3075 17395
rect 3045 17370 3050 17390
rect 3050 17370 3070 17390
rect 3070 17370 3075 17390
rect 3045 17365 3075 17370
rect 3125 17390 3155 17395
rect 3125 17370 3130 17390
rect 3130 17370 3150 17390
rect 3150 17370 3155 17390
rect 3125 17365 3155 17370
rect 3205 17390 3235 17395
rect 3205 17370 3210 17390
rect 3210 17370 3230 17390
rect 3230 17370 3235 17390
rect 3205 17365 3235 17370
rect 3285 17390 3315 17395
rect 3285 17370 3290 17390
rect 3290 17370 3310 17390
rect 3310 17370 3315 17390
rect 3285 17365 3315 17370
rect 3365 17390 3395 17395
rect 3365 17370 3370 17390
rect 3370 17370 3390 17390
rect 3390 17370 3395 17390
rect 3365 17365 3395 17370
rect 3445 17390 3475 17395
rect 3445 17370 3450 17390
rect 3450 17370 3470 17390
rect 3470 17370 3475 17390
rect 3445 17365 3475 17370
rect 3525 17390 3555 17395
rect 3525 17370 3530 17390
rect 3530 17370 3550 17390
rect 3550 17370 3555 17390
rect 3525 17365 3555 17370
rect 3605 17390 3635 17395
rect 3605 17370 3610 17390
rect 3610 17370 3630 17390
rect 3630 17370 3635 17390
rect 3605 17365 3635 17370
rect 3685 17390 3715 17395
rect 3685 17370 3690 17390
rect 3690 17370 3710 17390
rect 3710 17370 3715 17390
rect 3685 17365 3715 17370
rect 3765 17390 3795 17395
rect 3765 17370 3770 17390
rect 3770 17370 3790 17390
rect 3790 17370 3795 17390
rect 3765 17365 3795 17370
rect 3845 17390 3875 17395
rect 3845 17370 3850 17390
rect 3850 17370 3870 17390
rect 3870 17370 3875 17390
rect 3845 17365 3875 17370
rect 3925 17390 3955 17395
rect 3925 17370 3930 17390
rect 3930 17370 3950 17390
rect 3950 17370 3955 17390
rect 3925 17365 3955 17370
rect 4005 17390 4035 17395
rect 4005 17370 4010 17390
rect 4010 17370 4030 17390
rect 4030 17370 4035 17390
rect 4005 17365 4035 17370
rect 4085 17390 4115 17395
rect 4085 17370 4090 17390
rect 4090 17370 4110 17390
rect 4110 17370 4115 17390
rect 4085 17365 4115 17370
rect 4165 17390 4195 17395
rect 4165 17370 4170 17390
rect 4170 17370 4190 17390
rect 4190 17370 4195 17390
rect 4165 17365 4195 17370
rect 6245 17390 6275 17395
rect 6245 17370 6250 17390
rect 6250 17370 6270 17390
rect 6270 17370 6275 17390
rect 6245 17365 6275 17370
rect 6325 17390 6355 17395
rect 6325 17370 6330 17390
rect 6330 17370 6350 17390
rect 6350 17370 6355 17390
rect 6325 17365 6355 17370
rect 6405 17390 6435 17395
rect 6405 17370 6410 17390
rect 6410 17370 6430 17390
rect 6430 17370 6435 17390
rect 6405 17365 6435 17370
rect 6485 17390 6515 17395
rect 6485 17370 6490 17390
rect 6490 17370 6510 17390
rect 6510 17370 6515 17390
rect 6485 17365 6515 17370
rect 6565 17390 6595 17395
rect 6565 17370 6570 17390
rect 6570 17370 6590 17390
rect 6590 17370 6595 17390
rect 6565 17365 6595 17370
rect 6645 17390 6675 17395
rect 6645 17370 6650 17390
rect 6650 17370 6670 17390
rect 6670 17370 6675 17390
rect 6645 17365 6675 17370
rect 6725 17390 6755 17395
rect 6725 17370 6730 17390
rect 6730 17370 6750 17390
rect 6750 17370 6755 17390
rect 6725 17365 6755 17370
rect 6805 17390 6835 17395
rect 6805 17370 6810 17390
rect 6810 17370 6830 17390
rect 6830 17370 6835 17390
rect 6805 17365 6835 17370
rect 6885 17390 6915 17395
rect 6885 17370 6890 17390
rect 6890 17370 6910 17390
rect 6910 17370 6915 17390
rect 6885 17365 6915 17370
rect 6965 17390 6995 17395
rect 6965 17370 6970 17390
rect 6970 17370 6990 17390
rect 6990 17370 6995 17390
rect 6965 17365 6995 17370
rect 7045 17390 7075 17395
rect 7045 17370 7050 17390
rect 7050 17370 7070 17390
rect 7070 17370 7075 17390
rect 7045 17365 7075 17370
rect 7125 17390 7155 17395
rect 7125 17370 7130 17390
rect 7130 17370 7150 17390
rect 7150 17370 7155 17390
rect 7125 17365 7155 17370
rect 7205 17390 7235 17395
rect 7205 17370 7210 17390
rect 7210 17370 7230 17390
rect 7230 17370 7235 17390
rect 7205 17365 7235 17370
rect 7285 17390 7315 17395
rect 7285 17370 7290 17390
rect 7290 17370 7310 17390
rect 7310 17370 7315 17390
rect 7285 17365 7315 17370
rect 7365 17390 7395 17395
rect 7365 17370 7370 17390
rect 7370 17370 7390 17390
rect 7390 17370 7395 17390
rect 7365 17365 7395 17370
rect 7445 17390 7475 17395
rect 7445 17370 7450 17390
rect 7450 17370 7470 17390
rect 7470 17370 7475 17390
rect 7445 17365 7475 17370
rect 7525 17390 7555 17395
rect 7525 17370 7530 17390
rect 7530 17370 7550 17390
rect 7550 17370 7555 17390
rect 7525 17365 7555 17370
rect 7605 17390 7635 17395
rect 7605 17370 7610 17390
rect 7610 17370 7630 17390
rect 7630 17370 7635 17390
rect 7605 17365 7635 17370
rect 7685 17390 7715 17395
rect 7685 17370 7690 17390
rect 7690 17370 7710 17390
rect 7710 17370 7715 17390
rect 7685 17365 7715 17370
rect 7765 17390 7795 17395
rect 7765 17370 7770 17390
rect 7770 17370 7790 17390
rect 7790 17370 7795 17390
rect 7765 17365 7795 17370
rect 7845 17390 7875 17395
rect 7845 17370 7850 17390
rect 7850 17370 7870 17390
rect 7870 17370 7875 17390
rect 7845 17365 7875 17370
rect 7925 17390 7955 17395
rect 7925 17370 7930 17390
rect 7930 17370 7950 17390
rect 7950 17370 7955 17390
rect 7925 17365 7955 17370
rect 8005 17390 8035 17395
rect 8005 17370 8010 17390
rect 8010 17370 8030 17390
rect 8030 17370 8035 17390
rect 8005 17365 8035 17370
rect 8085 17390 8115 17395
rect 8085 17370 8090 17390
rect 8090 17370 8110 17390
rect 8110 17370 8115 17390
rect 8085 17365 8115 17370
rect 8165 17390 8195 17395
rect 8165 17370 8170 17390
rect 8170 17370 8190 17390
rect 8190 17370 8195 17390
rect 8165 17365 8195 17370
rect 8245 17390 8275 17395
rect 8245 17370 8250 17390
rect 8250 17370 8270 17390
rect 8270 17370 8275 17390
rect 8245 17365 8275 17370
rect 8325 17390 8355 17395
rect 8325 17370 8330 17390
rect 8330 17370 8350 17390
rect 8350 17370 8355 17390
rect 8325 17365 8355 17370
rect 8405 17390 8435 17395
rect 8405 17370 8410 17390
rect 8410 17370 8430 17390
rect 8430 17370 8435 17390
rect 8405 17365 8435 17370
rect 8485 17390 8515 17395
rect 8485 17370 8490 17390
rect 8490 17370 8510 17390
rect 8510 17370 8515 17390
rect 8485 17365 8515 17370
rect 8565 17390 8595 17395
rect 8565 17370 8570 17390
rect 8570 17370 8590 17390
rect 8590 17370 8595 17390
rect 8565 17365 8595 17370
rect 8645 17390 8675 17395
rect 8645 17370 8650 17390
rect 8650 17370 8670 17390
rect 8670 17370 8675 17390
rect 8645 17365 8675 17370
rect 8725 17390 8755 17395
rect 8725 17370 8730 17390
rect 8730 17370 8750 17390
rect 8750 17370 8755 17390
rect 8725 17365 8755 17370
rect 8805 17390 8835 17395
rect 8805 17370 8810 17390
rect 8810 17370 8830 17390
rect 8830 17370 8835 17390
rect 8805 17365 8835 17370
rect 8885 17390 8915 17395
rect 8885 17370 8890 17390
rect 8890 17370 8910 17390
rect 8910 17370 8915 17390
rect 8885 17365 8915 17370
rect 8965 17390 8995 17395
rect 8965 17370 8970 17390
rect 8970 17370 8990 17390
rect 8990 17370 8995 17390
rect 8965 17365 8995 17370
rect 9045 17390 9075 17395
rect 9045 17370 9050 17390
rect 9050 17370 9070 17390
rect 9070 17370 9075 17390
rect 9045 17365 9075 17370
rect 9125 17390 9155 17395
rect 9125 17370 9130 17390
rect 9130 17370 9150 17390
rect 9150 17370 9155 17390
rect 9125 17365 9155 17370
rect 9205 17390 9235 17395
rect 9205 17370 9210 17390
rect 9210 17370 9230 17390
rect 9230 17370 9235 17390
rect 9205 17365 9235 17370
rect 9285 17390 9315 17395
rect 9285 17370 9290 17390
rect 9290 17370 9310 17390
rect 9310 17370 9315 17390
rect 9285 17365 9315 17370
rect 9365 17390 9395 17395
rect 9365 17370 9370 17390
rect 9370 17370 9390 17390
rect 9390 17370 9395 17390
rect 9365 17365 9395 17370
rect 9445 17390 9475 17395
rect 9445 17370 9450 17390
rect 9450 17370 9470 17390
rect 9470 17370 9475 17390
rect 9445 17365 9475 17370
rect 11565 17390 11595 17395
rect 11565 17370 11570 17390
rect 11570 17370 11590 17390
rect 11590 17370 11595 17390
rect 11565 17365 11595 17370
rect 11645 17390 11675 17395
rect 11645 17370 11650 17390
rect 11650 17370 11670 17390
rect 11670 17370 11675 17390
rect 11645 17365 11675 17370
rect 11725 17390 11755 17395
rect 11725 17370 11730 17390
rect 11730 17370 11750 17390
rect 11750 17370 11755 17390
rect 11725 17365 11755 17370
rect 11805 17390 11835 17395
rect 11805 17370 11810 17390
rect 11810 17370 11830 17390
rect 11830 17370 11835 17390
rect 11805 17365 11835 17370
rect 11885 17390 11915 17395
rect 11885 17370 11890 17390
rect 11890 17370 11910 17390
rect 11910 17370 11915 17390
rect 11885 17365 11915 17370
rect 11965 17390 11995 17395
rect 11965 17370 11970 17390
rect 11970 17370 11990 17390
rect 11990 17370 11995 17390
rect 11965 17365 11995 17370
rect 12045 17390 12075 17395
rect 12045 17370 12050 17390
rect 12050 17370 12070 17390
rect 12070 17370 12075 17390
rect 12045 17365 12075 17370
rect 12125 17390 12155 17395
rect 12125 17370 12130 17390
rect 12130 17370 12150 17390
rect 12150 17370 12155 17390
rect 12125 17365 12155 17370
rect 12205 17390 12235 17395
rect 12205 17370 12210 17390
rect 12210 17370 12230 17390
rect 12230 17370 12235 17390
rect 12205 17365 12235 17370
rect 12285 17390 12315 17395
rect 12285 17370 12290 17390
rect 12290 17370 12310 17390
rect 12310 17370 12315 17390
rect 12285 17365 12315 17370
rect 12365 17390 12395 17395
rect 12365 17370 12370 17390
rect 12370 17370 12390 17390
rect 12390 17370 12395 17390
rect 12365 17365 12395 17370
rect 12445 17390 12475 17395
rect 12445 17370 12450 17390
rect 12450 17370 12470 17390
rect 12470 17370 12475 17390
rect 12445 17365 12475 17370
rect 12525 17390 12555 17395
rect 12525 17370 12530 17390
rect 12530 17370 12550 17390
rect 12550 17370 12555 17390
rect 12525 17365 12555 17370
rect 12605 17390 12635 17395
rect 12605 17370 12610 17390
rect 12610 17370 12630 17390
rect 12630 17370 12635 17390
rect 12605 17365 12635 17370
rect 12685 17390 12715 17395
rect 12685 17370 12690 17390
rect 12690 17370 12710 17390
rect 12710 17370 12715 17390
rect 12685 17365 12715 17370
rect 12765 17390 12795 17395
rect 12765 17370 12770 17390
rect 12770 17370 12790 17390
rect 12790 17370 12795 17390
rect 12765 17365 12795 17370
rect 12845 17390 12875 17395
rect 12845 17370 12850 17390
rect 12850 17370 12870 17390
rect 12870 17370 12875 17390
rect 12845 17365 12875 17370
rect 12925 17390 12955 17395
rect 12925 17370 12930 17390
rect 12930 17370 12950 17390
rect 12950 17370 12955 17390
rect 12925 17365 12955 17370
rect 13005 17390 13035 17395
rect 13005 17370 13010 17390
rect 13010 17370 13030 17390
rect 13030 17370 13035 17390
rect 13005 17365 13035 17370
rect 13085 17390 13115 17395
rect 13085 17370 13090 17390
rect 13090 17370 13110 17390
rect 13110 17370 13115 17390
rect 13085 17365 13115 17370
rect 13165 17390 13195 17395
rect 13165 17370 13170 17390
rect 13170 17370 13190 17390
rect 13190 17370 13195 17390
rect 13165 17365 13195 17370
rect 13245 17390 13275 17395
rect 13245 17370 13250 17390
rect 13250 17370 13270 17390
rect 13270 17370 13275 17390
rect 13245 17365 13275 17370
rect 13325 17390 13355 17395
rect 13325 17370 13330 17390
rect 13330 17370 13350 17390
rect 13350 17370 13355 17390
rect 13325 17365 13355 17370
rect 13405 17390 13435 17395
rect 13405 17370 13410 17390
rect 13410 17370 13430 17390
rect 13430 17370 13435 17390
rect 13405 17365 13435 17370
rect 13485 17390 13515 17395
rect 13485 17370 13490 17390
rect 13490 17370 13510 17390
rect 13510 17370 13515 17390
rect 13485 17365 13515 17370
rect 13565 17390 13595 17395
rect 13565 17370 13570 17390
rect 13570 17370 13590 17390
rect 13590 17370 13595 17390
rect 13565 17365 13595 17370
rect 13645 17390 13675 17395
rect 13645 17370 13650 17390
rect 13650 17370 13670 17390
rect 13670 17370 13675 17390
rect 13645 17365 13675 17370
rect 13725 17390 13755 17395
rect 13725 17370 13730 17390
rect 13730 17370 13750 17390
rect 13750 17370 13755 17390
rect 13725 17365 13755 17370
rect 13805 17390 13835 17395
rect 13805 17370 13810 17390
rect 13810 17370 13830 17390
rect 13830 17370 13835 17390
rect 13805 17365 13835 17370
rect 13885 17390 13915 17395
rect 13885 17370 13890 17390
rect 13890 17370 13910 17390
rect 13910 17370 13915 17390
rect 13885 17365 13915 17370
rect 13965 17390 13995 17395
rect 13965 17370 13970 17390
rect 13970 17370 13990 17390
rect 13990 17370 13995 17390
rect 13965 17365 13995 17370
rect 14045 17390 14075 17395
rect 14045 17370 14050 17390
rect 14050 17370 14070 17390
rect 14070 17370 14075 17390
rect 14045 17365 14075 17370
rect 14125 17390 14155 17395
rect 14125 17370 14130 17390
rect 14130 17370 14150 17390
rect 14150 17370 14155 17390
rect 14125 17365 14155 17370
rect 14205 17390 14235 17395
rect 14205 17370 14210 17390
rect 14210 17370 14230 17390
rect 14230 17370 14235 17390
rect 14205 17365 14235 17370
rect 14285 17390 14315 17395
rect 14285 17370 14290 17390
rect 14290 17370 14310 17390
rect 14310 17370 14315 17390
rect 14285 17365 14315 17370
rect 14365 17390 14395 17395
rect 14365 17370 14370 17390
rect 14370 17370 14390 17390
rect 14390 17370 14395 17390
rect 14365 17365 14395 17370
rect 14445 17390 14475 17395
rect 14445 17370 14450 17390
rect 14450 17370 14470 17390
rect 14470 17370 14475 17390
rect 14445 17365 14475 17370
rect 14525 17390 14555 17395
rect 14525 17370 14530 17390
rect 14530 17370 14550 17390
rect 14550 17370 14555 17390
rect 14525 17365 14555 17370
rect 14605 17390 14635 17395
rect 14605 17370 14610 17390
rect 14610 17370 14630 17390
rect 14630 17370 14635 17390
rect 14605 17365 14635 17370
rect 14685 17390 14715 17395
rect 14685 17370 14690 17390
rect 14690 17370 14710 17390
rect 14710 17370 14715 17390
rect 14685 17365 14715 17370
rect 16765 17390 16795 17395
rect 16765 17370 16770 17390
rect 16770 17370 16790 17390
rect 16790 17370 16795 17390
rect 16765 17365 16795 17370
rect 16845 17390 16875 17395
rect 16845 17370 16850 17390
rect 16850 17370 16870 17390
rect 16870 17370 16875 17390
rect 16845 17365 16875 17370
rect 16925 17390 16955 17395
rect 16925 17370 16930 17390
rect 16930 17370 16950 17390
rect 16950 17370 16955 17390
rect 16925 17365 16955 17370
rect 17005 17390 17035 17395
rect 17005 17370 17010 17390
rect 17010 17370 17030 17390
rect 17030 17370 17035 17390
rect 17005 17365 17035 17370
rect 17085 17390 17115 17395
rect 17085 17370 17090 17390
rect 17090 17370 17110 17390
rect 17110 17370 17115 17390
rect 17085 17365 17115 17370
rect 17165 17390 17195 17395
rect 17165 17370 17170 17390
rect 17170 17370 17190 17390
rect 17190 17370 17195 17390
rect 17165 17365 17195 17370
rect 17245 17390 17275 17395
rect 17245 17370 17250 17390
rect 17250 17370 17270 17390
rect 17270 17370 17275 17390
rect 17245 17365 17275 17370
rect 17325 17390 17355 17395
rect 17325 17370 17330 17390
rect 17330 17370 17350 17390
rect 17350 17370 17355 17390
rect 17325 17365 17355 17370
rect 17405 17390 17435 17395
rect 17405 17370 17410 17390
rect 17410 17370 17430 17390
rect 17430 17370 17435 17390
rect 17405 17365 17435 17370
rect 17485 17390 17515 17395
rect 17485 17370 17490 17390
rect 17490 17370 17510 17390
rect 17510 17370 17515 17390
rect 17485 17365 17515 17370
rect 17565 17390 17595 17395
rect 17565 17370 17570 17390
rect 17570 17370 17590 17390
rect 17590 17370 17595 17390
rect 17565 17365 17595 17370
rect 17645 17390 17675 17395
rect 17645 17370 17650 17390
rect 17650 17370 17670 17390
rect 17670 17370 17675 17390
rect 17645 17365 17675 17370
rect 17725 17390 17755 17395
rect 17725 17370 17730 17390
rect 17730 17370 17750 17390
rect 17750 17370 17755 17390
rect 17725 17365 17755 17370
rect 17805 17390 17835 17395
rect 17805 17370 17810 17390
rect 17810 17370 17830 17390
rect 17830 17370 17835 17390
rect 17805 17365 17835 17370
rect 17885 17390 17915 17395
rect 17885 17370 17890 17390
rect 17890 17370 17910 17390
rect 17910 17370 17915 17390
rect 17885 17365 17915 17370
rect 17965 17390 17995 17395
rect 17965 17370 17970 17390
rect 17970 17370 17990 17390
rect 17990 17370 17995 17390
rect 17965 17365 17995 17370
rect 18045 17390 18075 17395
rect 18045 17370 18050 17390
rect 18050 17370 18070 17390
rect 18070 17370 18075 17390
rect 18045 17365 18075 17370
rect 18125 17390 18155 17395
rect 18125 17370 18130 17390
rect 18130 17370 18150 17390
rect 18150 17370 18155 17390
rect 18125 17365 18155 17370
rect 18205 17390 18235 17395
rect 18205 17370 18210 17390
rect 18210 17370 18230 17390
rect 18230 17370 18235 17390
rect 18205 17365 18235 17370
rect 18285 17390 18315 17395
rect 18285 17370 18290 17390
rect 18290 17370 18310 17390
rect 18310 17370 18315 17390
rect 18285 17365 18315 17370
rect 18365 17390 18395 17395
rect 18365 17370 18370 17390
rect 18370 17370 18390 17390
rect 18390 17370 18395 17390
rect 18365 17365 18395 17370
rect 18445 17390 18475 17395
rect 18445 17370 18450 17390
rect 18450 17370 18470 17390
rect 18470 17370 18475 17390
rect 18445 17365 18475 17370
rect 18525 17390 18555 17395
rect 18525 17370 18530 17390
rect 18530 17370 18550 17390
rect 18550 17370 18555 17390
rect 18525 17365 18555 17370
rect 18605 17390 18635 17395
rect 18605 17370 18610 17390
rect 18610 17370 18630 17390
rect 18630 17370 18635 17390
rect 18605 17365 18635 17370
rect 18685 17390 18715 17395
rect 18685 17370 18690 17390
rect 18690 17370 18710 17390
rect 18710 17370 18715 17390
rect 18685 17365 18715 17370
rect 18765 17390 18795 17395
rect 18765 17370 18770 17390
rect 18770 17370 18790 17390
rect 18790 17370 18795 17390
rect 18765 17365 18795 17370
rect 18845 17390 18875 17395
rect 18845 17370 18850 17390
rect 18850 17370 18870 17390
rect 18870 17370 18875 17390
rect 18845 17365 18875 17370
rect 18925 17390 18955 17395
rect 18925 17370 18930 17390
rect 18930 17370 18950 17390
rect 18950 17370 18955 17390
rect 18925 17365 18955 17370
rect 19005 17390 19035 17395
rect 19005 17370 19010 17390
rect 19010 17370 19030 17390
rect 19030 17370 19035 17390
rect 19005 17365 19035 17370
rect 19085 17390 19115 17395
rect 19085 17370 19090 17390
rect 19090 17370 19110 17390
rect 19110 17370 19115 17390
rect 19085 17365 19115 17370
rect 19165 17390 19195 17395
rect 19165 17370 19170 17390
rect 19170 17370 19190 17390
rect 19190 17370 19195 17390
rect 19165 17365 19195 17370
rect 19245 17390 19275 17395
rect 19245 17370 19250 17390
rect 19250 17370 19270 17390
rect 19270 17370 19275 17390
rect 19245 17365 19275 17370
rect 19325 17390 19355 17395
rect 19325 17370 19330 17390
rect 19330 17370 19350 17390
rect 19350 17370 19355 17390
rect 19325 17365 19355 17370
rect 19405 17390 19435 17395
rect 19405 17370 19410 17390
rect 19410 17370 19430 17390
rect 19430 17370 19435 17390
rect 19405 17365 19435 17370
rect 19485 17390 19515 17395
rect 19485 17370 19490 17390
rect 19490 17370 19510 17390
rect 19510 17370 19515 17390
rect 19485 17365 19515 17370
rect 19565 17390 19595 17395
rect 19565 17370 19570 17390
rect 19570 17370 19590 17390
rect 19590 17370 19595 17390
rect 19565 17365 19595 17370
rect 19645 17390 19675 17395
rect 19645 17370 19650 17390
rect 19650 17370 19670 17390
rect 19670 17370 19675 17390
rect 19645 17365 19675 17370
rect 19725 17390 19755 17395
rect 19725 17370 19730 17390
rect 19730 17370 19750 17390
rect 19750 17370 19755 17390
rect 19725 17365 19755 17370
rect 19805 17390 19835 17395
rect 19805 17370 19810 17390
rect 19810 17370 19830 17390
rect 19830 17370 19835 17390
rect 19805 17365 19835 17370
rect 19885 17390 19915 17395
rect 19885 17370 19890 17390
rect 19890 17370 19910 17390
rect 19910 17370 19915 17390
rect 19885 17365 19915 17370
rect 19965 17390 19995 17395
rect 19965 17370 19970 17390
rect 19970 17370 19990 17390
rect 19990 17370 19995 17390
rect 19965 17365 19995 17370
rect 20045 17390 20075 17395
rect 20045 17370 20050 17390
rect 20050 17370 20070 17390
rect 20070 17370 20075 17390
rect 20045 17365 20075 17370
rect 20125 17390 20155 17395
rect 20125 17370 20130 17390
rect 20130 17370 20150 17390
rect 20150 17370 20155 17390
rect 20125 17365 20155 17370
rect 20205 17390 20235 17395
rect 20205 17370 20210 17390
rect 20210 17370 20230 17390
rect 20230 17370 20235 17390
rect 20205 17365 20235 17370
rect 20285 17390 20315 17395
rect 20285 17370 20290 17390
rect 20290 17370 20310 17390
rect 20310 17370 20315 17390
rect 20285 17365 20315 17370
rect 20365 17390 20395 17395
rect 20365 17370 20370 17390
rect 20370 17370 20390 17390
rect 20390 17370 20395 17390
rect 20365 17365 20395 17370
rect 20445 17390 20475 17395
rect 20445 17370 20450 17390
rect 20450 17370 20470 17390
rect 20470 17370 20475 17390
rect 20445 17365 20475 17370
rect 20525 17390 20555 17395
rect 20525 17370 20530 17390
rect 20530 17370 20550 17390
rect 20550 17370 20555 17390
rect 20525 17365 20555 17370
rect 20605 17390 20635 17395
rect 20605 17370 20610 17390
rect 20610 17370 20630 17390
rect 20630 17370 20635 17390
rect 20605 17365 20635 17370
rect 20685 17390 20715 17395
rect 20685 17370 20690 17390
rect 20690 17370 20710 17390
rect 20710 17370 20715 17390
rect 20685 17365 20715 17370
rect 20765 17390 20795 17395
rect 20765 17370 20770 17390
rect 20770 17370 20790 17390
rect 20790 17370 20795 17390
rect 20765 17365 20795 17370
rect 20845 17390 20875 17395
rect 20845 17370 20850 17390
rect 20850 17370 20870 17390
rect 20870 17370 20875 17390
rect 20845 17365 20875 17370
rect 20925 17390 20955 17395
rect 20925 17370 20930 17390
rect 20930 17370 20950 17390
rect 20950 17370 20955 17390
rect 20925 17365 20955 17370
rect 5 17230 35 17235
rect 5 17210 10 17230
rect 10 17210 30 17230
rect 30 17210 35 17230
rect 5 17205 35 17210
rect 85 17230 115 17235
rect 85 17210 90 17230
rect 90 17210 110 17230
rect 110 17210 115 17230
rect 85 17205 115 17210
rect 165 17230 195 17235
rect 165 17210 170 17230
rect 170 17210 190 17230
rect 190 17210 195 17230
rect 165 17205 195 17210
rect 245 17230 275 17235
rect 245 17210 250 17230
rect 250 17210 270 17230
rect 270 17210 275 17230
rect 245 17205 275 17210
rect 325 17230 355 17235
rect 325 17210 330 17230
rect 330 17210 350 17230
rect 350 17210 355 17230
rect 325 17205 355 17210
rect 405 17230 435 17235
rect 405 17210 410 17230
rect 410 17210 430 17230
rect 430 17210 435 17230
rect 405 17205 435 17210
rect 485 17230 515 17235
rect 485 17210 490 17230
rect 490 17210 510 17230
rect 510 17210 515 17230
rect 485 17205 515 17210
rect 565 17230 595 17235
rect 565 17210 570 17230
rect 570 17210 590 17230
rect 590 17210 595 17230
rect 565 17205 595 17210
rect 645 17230 675 17235
rect 645 17210 650 17230
rect 650 17210 670 17230
rect 670 17210 675 17230
rect 645 17205 675 17210
rect 725 17230 755 17235
rect 725 17210 730 17230
rect 730 17210 750 17230
rect 750 17210 755 17230
rect 725 17205 755 17210
rect 805 17230 835 17235
rect 805 17210 810 17230
rect 810 17210 830 17230
rect 830 17210 835 17230
rect 805 17205 835 17210
rect 885 17230 915 17235
rect 885 17210 890 17230
rect 890 17210 910 17230
rect 910 17210 915 17230
rect 885 17205 915 17210
rect 965 17230 995 17235
rect 965 17210 970 17230
rect 970 17210 990 17230
rect 990 17210 995 17230
rect 965 17205 995 17210
rect 1045 17230 1075 17235
rect 1045 17210 1050 17230
rect 1050 17210 1070 17230
rect 1070 17210 1075 17230
rect 1045 17205 1075 17210
rect 1125 17230 1155 17235
rect 1125 17210 1130 17230
rect 1130 17210 1150 17230
rect 1150 17210 1155 17230
rect 1125 17205 1155 17210
rect 1205 17230 1235 17235
rect 1205 17210 1210 17230
rect 1210 17210 1230 17230
rect 1230 17210 1235 17230
rect 1205 17205 1235 17210
rect 1285 17230 1315 17235
rect 1285 17210 1290 17230
rect 1290 17210 1310 17230
rect 1310 17210 1315 17230
rect 1285 17205 1315 17210
rect 1365 17230 1395 17235
rect 1365 17210 1370 17230
rect 1370 17210 1390 17230
rect 1390 17210 1395 17230
rect 1365 17205 1395 17210
rect 1445 17230 1475 17235
rect 1445 17210 1450 17230
rect 1450 17210 1470 17230
rect 1470 17210 1475 17230
rect 1445 17205 1475 17210
rect 1525 17230 1555 17235
rect 1525 17210 1530 17230
rect 1530 17210 1550 17230
rect 1550 17210 1555 17230
rect 1525 17205 1555 17210
rect 1605 17230 1635 17235
rect 1605 17210 1610 17230
rect 1610 17210 1630 17230
rect 1630 17210 1635 17230
rect 1605 17205 1635 17210
rect 1685 17230 1715 17235
rect 1685 17210 1690 17230
rect 1690 17210 1710 17230
rect 1710 17210 1715 17230
rect 1685 17205 1715 17210
rect 1765 17230 1795 17235
rect 1765 17210 1770 17230
rect 1770 17210 1790 17230
rect 1790 17210 1795 17230
rect 1765 17205 1795 17210
rect 1845 17230 1875 17235
rect 1845 17210 1850 17230
rect 1850 17210 1870 17230
rect 1870 17210 1875 17230
rect 1845 17205 1875 17210
rect 1925 17230 1955 17235
rect 1925 17210 1930 17230
rect 1930 17210 1950 17230
rect 1950 17210 1955 17230
rect 1925 17205 1955 17210
rect 2005 17230 2035 17235
rect 2005 17210 2010 17230
rect 2010 17210 2030 17230
rect 2030 17210 2035 17230
rect 2005 17205 2035 17210
rect 2085 17230 2115 17235
rect 2085 17210 2090 17230
rect 2090 17210 2110 17230
rect 2110 17210 2115 17230
rect 2085 17205 2115 17210
rect 2165 17230 2195 17235
rect 2165 17210 2170 17230
rect 2170 17210 2190 17230
rect 2190 17210 2195 17230
rect 2165 17205 2195 17210
rect 2245 17230 2275 17235
rect 2245 17210 2250 17230
rect 2250 17210 2270 17230
rect 2270 17210 2275 17230
rect 2245 17205 2275 17210
rect 2325 17230 2355 17235
rect 2325 17210 2330 17230
rect 2330 17210 2350 17230
rect 2350 17210 2355 17230
rect 2325 17205 2355 17210
rect 2405 17230 2435 17235
rect 2405 17210 2410 17230
rect 2410 17210 2430 17230
rect 2430 17210 2435 17230
rect 2405 17205 2435 17210
rect 2485 17230 2515 17235
rect 2485 17210 2490 17230
rect 2490 17210 2510 17230
rect 2510 17210 2515 17230
rect 2485 17205 2515 17210
rect 2565 17230 2595 17235
rect 2565 17210 2570 17230
rect 2570 17210 2590 17230
rect 2590 17210 2595 17230
rect 2565 17205 2595 17210
rect 2645 17230 2675 17235
rect 2645 17210 2650 17230
rect 2650 17210 2670 17230
rect 2670 17210 2675 17230
rect 2645 17205 2675 17210
rect 2725 17230 2755 17235
rect 2725 17210 2730 17230
rect 2730 17210 2750 17230
rect 2750 17210 2755 17230
rect 2725 17205 2755 17210
rect 2805 17230 2835 17235
rect 2805 17210 2810 17230
rect 2810 17210 2830 17230
rect 2830 17210 2835 17230
rect 2805 17205 2835 17210
rect 2885 17230 2915 17235
rect 2885 17210 2890 17230
rect 2890 17210 2910 17230
rect 2910 17210 2915 17230
rect 2885 17205 2915 17210
rect 2965 17230 2995 17235
rect 2965 17210 2970 17230
rect 2970 17210 2990 17230
rect 2990 17210 2995 17230
rect 2965 17205 2995 17210
rect 3045 17230 3075 17235
rect 3045 17210 3050 17230
rect 3050 17210 3070 17230
rect 3070 17210 3075 17230
rect 3045 17205 3075 17210
rect 3125 17230 3155 17235
rect 3125 17210 3130 17230
rect 3130 17210 3150 17230
rect 3150 17210 3155 17230
rect 3125 17205 3155 17210
rect 3205 17230 3235 17235
rect 3205 17210 3210 17230
rect 3210 17210 3230 17230
rect 3230 17210 3235 17230
rect 3205 17205 3235 17210
rect 3285 17230 3315 17235
rect 3285 17210 3290 17230
rect 3290 17210 3310 17230
rect 3310 17210 3315 17230
rect 3285 17205 3315 17210
rect 3365 17230 3395 17235
rect 3365 17210 3370 17230
rect 3370 17210 3390 17230
rect 3390 17210 3395 17230
rect 3365 17205 3395 17210
rect 3445 17230 3475 17235
rect 3445 17210 3450 17230
rect 3450 17210 3470 17230
rect 3470 17210 3475 17230
rect 3445 17205 3475 17210
rect 3525 17230 3555 17235
rect 3525 17210 3530 17230
rect 3530 17210 3550 17230
rect 3550 17210 3555 17230
rect 3525 17205 3555 17210
rect 3605 17230 3635 17235
rect 3605 17210 3610 17230
rect 3610 17210 3630 17230
rect 3630 17210 3635 17230
rect 3605 17205 3635 17210
rect 3685 17230 3715 17235
rect 3685 17210 3690 17230
rect 3690 17210 3710 17230
rect 3710 17210 3715 17230
rect 3685 17205 3715 17210
rect 3765 17230 3795 17235
rect 3765 17210 3770 17230
rect 3770 17210 3790 17230
rect 3790 17210 3795 17230
rect 3765 17205 3795 17210
rect 3845 17230 3875 17235
rect 3845 17210 3850 17230
rect 3850 17210 3870 17230
rect 3870 17210 3875 17230
rect 3845 17205 3875 17210
rect 3925 17230 3955 17235
rect 3925 17210 3930 17230
rect 3930 17210 3950 17230
rect 3950 17210 3955 17230
rect 3925 17205 3955 17210
rect 4005 17230 4035 17235
rect 4005 17210 4010 17230
rect 4010 17210 4030 17230
rect 4030 17210 4035 17230
rect 4005 17205 4035 17210
rect 4085 17230 4115 17235
rect 4085 17210 4090 17230
rect 4090 17210 4110 17230
rect 4110 17210 4115 17230
rect 4085 17205 4115 17210
rect 4165 17230 4195 17235
rect 4165 17210 4170 17230
rect 4170 17210 4190 17230
rect 4190 17210 4195 17230
rect 4165 17205 4195 17210
rect 6245 17230 6275 17235
rect 6245 17210 6250 17230
rect 6250 17210 6270 17230
rect 6270 17210 6275 17230
rect 6245 17205 6275 17210
rect 6325 17230 6355 17235
rect 6325 17210 6330 17230
rect 6330 17210 6350 17230
rect 6350 17210 6355 17230
rect 6325 17205 6355 17210
rect 6405 17230 6435 17235
rect 6405 17210 6410 17230
rect 6410 17210 6430 17230
rect 6430 17210 6435 17230
rect 6405 17205 6435 17210
rect 6485 17230 6515 17235
rect 6485 17210 6490 17230
rect 6490 17210 6510 17230
rect 6510 17210 6515 17230
rect 6485 17205 6515 17210
rect 6565 17230 6595 17235
rect 6565 17210 6570 17230
rect 6570 17210 6590 17230
rect 6590 17210 6595 17230
rect 6565 17205 6595 17210
rect 6645 17230 6675 17235
rect 6645 17210 6650 17230
rect 6650 17210 6670 17230
rect 6670 17210 6675 17230
rect 6645 17205 6675 17210
rect 6725 17230 6755 17235
rect 6725 17210 6730 17230
rect 6730 17210 6750 17230
rect 6750 17210 6755 17230
rect 6725 17205 6755 17210
rect 6805 17230 6835 17235
rect 6805 17210 6810 17230
rect 6810 17210 6830 17230
rect 6830 17210 6835 17230
rect 6805 17205 6835 17210
rect 6885 17230 6915 17235
rect 6885 17210 6890 17230
rect 6890 17210 6910 17230
rect 6910 17210 6915 17230
rect 6885 17205 6915 17210
rect 6965 17230 6995 17235
rect 6965 17210 6970 17230
rect 6970 17210 6990 17230
rect 6990 17210 6995 17230
rect 6965 17205 6995 17210
rect 7045 17230 7075 17235
rect 7045 17210 7050 17230
rect 7050 17210 7070 17230
rect 7070 17210 7075 17230
rect 7045 17205 7075 17210
rect 7125 17230 7155 17235
rect 7125 17210 7130 17230
rect 7130 17210 7150 17230
rect 7150 17210 7155 17230
rect 7125 17205 7155 17210
rect 7205 17230 7235 17235
rect 7205 17210 7210 17230
rect 7210 17210 7230 17230
rect 7230 17210 7235 17230
rect 7205 17205 7235 17210
rect 7285 17230 7315 17235
rect 7285 17210 7290 17230
rect 7290 17210 7310 17230
rect 7310 17210 7315 17230
rect 7285 17205 7315 17210
rect 7365 17230 7395 17235
rect 7365 17210 7370 17230
rect 7370 17210 7390 17230
rect 7390 17210 7395 17230
rect 7365 17205 7395 17210
rect 7445 17230 7475 17235
rect 7445 17210 7450 17230
rect 7450 17210 7470 17230
rect 7470 17210 7475 17230
rect 7445 17205 7475 17210
rect 7525 17230 7555 17235
rect 7525 17210 7530 17230
rect 7530 17210 7550 17230
rect 7550 17210 7555 17230
rect 7525 17205 7555 17210
rect 7605 17230 7635 17235
rect 7605 17210 7610 17230
rect 7610 17210 7630 17230
rect 7630 17210 7635 17230
rect 7605 17205 7635 17210
rect 7685 17230 7715 17235
rect 7685 17210 7690 17230
rect 7690 17210 7710 17230
rect 7710 17210 7715 17230
rect 7685 17205 7715 17210
rect 7765 17230 7795 17235
rect 7765 17210 7770 17230
rect 7770 17210 7790 17230
rect 7790 17210 7795 17230
rect 7765 17205 7795 17210
rect 7845 17230 7875 17235
rect 7845 17210 7850 17230
rect 7850 17210 7870 17230
rect 7870 17210 7875 17230
rect 7845 17205 7875 17210
rect 7925 17230 7955 17235
rect 7925 17210 7930 17230
rect 7930 17210 7950 17230
rect 7950 17210 7955 17230
rect 7925 17205 7955 17210
rect 8005 17230 8035 17235
rect 8005 17210 8010 17230
rect 8010 17210 8030 17230
rect 8030 17210 8035 17230
rect 8005 17205 8035 17210
rect 8085 17230 8115 17235
rect 8085 17210 8090 17230
rect 8090 17210 8110 17230
rect 8110 17210 8115 17230
rect 8085 17205 8115 17210
rect 8165 17230 8195 17235
rect 8165 17210 8170 17230
rect 8170 17210 8190 17230
rect 8190 17210 8195 17230
rect 8165 17205 8195 17210
rect 8245 17230 8275 17235
rect 8245 17210 8250 17230
rect 8250 17210 8270 17230
rect 8270 17210 8275 17230
rect 8245 17205 8275 17210
rect 8325 17230 8355 17235
rect 8325 17210 8330 17230
rect 8330 17210 8350 17230
rect 8350 17210 8355 17230
rect 8325 17205 8355 17210
rect 8405 17230 8435 17235
rect 8405 17210 8410 17230
rect 8410 17210 8430 17230
rect 8430 17210 8435 17230
rect 8405 17205 8435 17210
rect 8485 17230 8515 17235
rect 8485 17210 8490 17230
rect 8490 17210 8510 17230
rect 8510 17210 8515 17230
rect 8485 17205 8515 17210
rect 8565 17230 8595 17235
rect 8565 17210 8570 17230
rect 8570 17210 8590 17230
rect 8590 17210 8595 17230
rect 8565 17205 8595 17210
rect 8645 17230 8675 17235
rect 8645 17210 8650 17230
rect 8650 17210 8670 17230
rect 8670 17210 8675 17230
rect 8645 17205 8675 17210
rect 8725 17230 8755 17235
rect 8725 17210 8730 17230
rect 8730 17210 8750 17230
rect 8750 17210 8755 17230
rect 8725 17205 8755 17210
rect 8805 17230 8835 17235
rect 8805 17210 8810 17230
rect 8810 17210 8830 17230
rect 8830 17210 8835 17230
rect 8805 17205 8835 17210
rect 8885 17230 8915 17235
rect 8885 17210 8890 17230
rect 8890 17210 8910 17230
rect 8910 17210 8915 17230
rect 8885 17205 8915 17210
rect 8965 17230 8995 17235
rect 8965 17210 8970 17230
rect 8970 17210 8990 17230
rect 8990 17210 8995 17230
rect 8965 17205 8995 17210
rect 9045 17230 9075 17235
rect 9045 17210 9050 17230
rect 9050 17210 9070 17230
rect 9070 17210 9075 17230
rect 9045 17205 9075 17210
rect 9125 17230 9155 17235
rect 9125 17210 9130 17230
rect 9130 17210 9150 17230
rect 9150 17210 9155 17230
rect 9125 17205 9155 17210
rect 9205 17230 9235 17235
rect 9205 17210 9210 17230
rect 9210 17210 9230 17230
rect 9230 17210 9235 17230
rect 9205 17205 9235 17210
rect 9285 17230 9315 17235
rect 9285 17210 9290 17230
rect 9290 17210 9310 17230
rect 9310 17210 9315 17230
rect 9285 17205 9315 17210
rect 9365 17230 9395 17235
rect 9365 17210 9370 17230
rect 9370 17210 9390 17230
rect 9390 17210 9395 17230
rect 9365 17205 9395 17210
rect 9445 17230 9475 17235
rect 9445 17210 9450 17230
rect 9450 17210 9470 17230
rect 9470 17210 9475 17230
rect 9445 17205 9475 17210
rect 11565 17230 11595 17235
rect 11565 17210 11570 17230
rect 11570 17210 11590 17230
rect 11590 17210 11595 17230
rect 11565 17205 11595 17210
rect 11645 17230 11675 17235
rect 11645 17210 11650 17230
rect 11650 17210 11670 17230
rect 11670 17210 11675 17230
rect 11645 17205 11675 17210
rect 11725 17230 11755 17235
rect 11725 17210 11730 17230
rect 11730 17210 11750 17230
rect 11750 17210 11755 17230
rect 11725 17205 11755 17210
rect 11805 17230 11835 17235
rect 11805 17210 11810 17230
rect 11810 17210 11830 17230
rect 11830 17210 11835 17230
rect 11805 17205 11835 17210
rect 11885 17230 11915 17235
rect 11885 17210 11890 17230
rect 11890 17210 11910 17230
rect 11910 17210 11915 17230
rect 11885 17205 11915 17210
rect 11965 17230 11995 17235
rect 11965 17210 11970 17230
rect 11970 17210 11990 17230
rect 11990 17210 11995 17230
rect 11965 17205 11995 17210
rect 12045 17230 12075 17235
rect 12045 17210 12050 17230
rect 12050 17210 12070 17230
rect 12070 17210 12075 17230
rect 12045 17205 12075 17210
rect 12125 17230 12155 17235
rect 12125 17210 12130 17230
rect 12130 17210 12150 17230
rect 12150 17210 12155 17230
rect 12125 17205 12155 17210
rect 12205 17230 12235 17235
rect 12205 17210 12210 17230
rect 12210 17210 12230 17230
rect 12230 17210 12235 17230
rect 12205 17205 12235 17210
rect 12285 17230 12315 17235
rect 12285 17210 12290 17230
rect 12290 17210 12310 17230
rect 12310 17210 12315 17230
rect 12285 17205 12315 17210
rect 12365 17230 12395 17235
rect 12365 17210 12370 17230
rect 12370 17210 12390 17230
rect 12390 17210 12395 17230
rect 12365 17205 12395 17210
rect 12445 17230 12475 17235
rect 12445 17210 12450 17230
rect 12450 17210 12470 17230
rect 12470 17210 12475 17230
rect 12445 17205 12475 17210
rect 12525 17230 12555 17235
rect 12525 17210 12530 17230
rect 12530 17210 12550 17230
rect 12550 17210 12555 17230
rect 12525 17205 12555 17210
rect 12605 17230 12635 17235
rect 12605 17210 12610 17230
rect 12610 17210 12630 17230
rect 12630 17210 12635 17230
rect 12605 17205 12635 17210
rect 12685 17230 12715 17235
rect 12685 17210 12690 17230
rect 12690 17210 12710 17230
rect 12710 17210 12715 17230
rect 12685 17205 12715 17210
rect 12765 17230 12795 17235
rect 12765 17210 12770 17230
rect 12770 17210 12790 17230
rect 12790 17210 12795 17230
rect 12765 17205 12795 17210
rect 12845 17230 12875 17235
rect 12845 17210 12850 17230
rect 12850 17210 12870 17230
rect 12870 17210 12875 17230
rect 12845 17205 12875 17210
rect 12925 17230 12955 17235
rect 12925 17210 12930 17230
rect 12930 17210 12950 17230
rect 12950 17210 12955 17230
rect 12925 17205 12955 17210
rect 13005 17230 13035 17235
rect 13005 17210 13010 17230
rect 13010 17210 13030 17230
rect 13030 17210 13035 17230
rect 13005 17205 13035 17210
rect 13085 17230 13115 17235
rect 13085 17210 13090 17230
rect 13090 17210 13110 17230
rect 13110 17210 13115 17230
rect 13085 17205 13115 17210
rect 13165 17230 13195 17235
rect 13165 17210 13170 17230
rect 13170 17210 13190 17230
rect 13190 17210 13195 17230
rect 13165 17205 13195 17210
rect 13245 17230 13275 17235
rect 13245 17210 13250 17230
rect 13250 17210 13270 17230
rect 13270 17210 13275 17230
rect 13245 17205 13275 17210
rect 13325 17230 13355 17235
rect 13325 17210 13330 17230
rect 13330 17210 13350 17230
rect 13350 17210 13355 17230
rect 13325 17205 13355 17210
rect 13405 17230 13435 17235
rect 13405 17210 13410 17230
rect 13410 17210 13430 17230
rect 13430 17210 13435 17230
rect 13405 17205 13435 17210
rect 13485 17230 13515 17235
rect 13485 17210 13490 17230
rect 13490 17210 13510 17230
rect 13510 17210 13515 17230
rect 13485 17205 13515 17210
rect 13565 17230 13595 17235
rect 13565 17210 13570 17230
rect 13570 17210 13590 17230
rect 13590 17210 13595 17230
rect 13565 17205 13595 17210
rect 13645 17230 13675 17235
rect 13645 17210 13650 17230
rect 13650 17210 13670 17230
rect 13670 17210 13675 17230
rect 13645 17205 13675 17210
rect 13725 17230 13755 17235
rect 13725 17210 13730 17230
rect 13730 17210 13750 17230
rect 13750 17210 13755 17230
rect 13725 17205 13755 17210
rect 13805 17230 13835 17235
rect 13805 17210 13810 17230
rect 13810 17210 13830 17230
rect 13830 17210 13835 17230
rect 13805 17205 13835 17210
rect 13885 17230 13915 17235
rect 13885 17210 13890 17230
rect 13890 17210 13910 17230
rect 13910 17210 13915 17230
rect 13885 17205 13915 17210
rect 13965 17230 13995 17235
rect 13965 17210 13970 17230
rect 13970 17210 13990 17230
rect 13990 17210 13995 17230
rect 13965 17205 13995 17210
rect 14045 17230 14075 17235
rect 14045 17210 14050 17230
rect 14050 17210 14070 17230
rect 14070 17210 14075 17230
rect 14045 17205 14075 17210
rect 14125 17230 14155 17235
rect 14125 17210 14130 17230
rect 14130 17210 14150 17230
rect 14150 17210 14155 17230
rect 14125 17205 14155 17210
rect 14205 17230 14235 17235
rect 14205 17210 14210 17230
rect 14210 17210 14230 17230
rect 14230 17210 14235 17230
rect 14205 17205 14235 17210
rect 14285 17230 14315 17235
rect 14285 17210 14290 17230
rect 14290 17210 14310 17230
rect 14310 17210 14315 17230
rect 14285 17205 14315 17210
rect 14365 17230 14395 17235
rect 14365 17210 14370 17230
rect 14370 17210 14390 17230
rect 14390 17210 14395 17230
rect 14365 17205 14395 17210
rect 14445 17230 14475 17235
rect 14445 17210 14450 17230
rect 14450 17210 14470 17230
rect 14470 17210 14475 17230
rect 14445 17205 14475 17210
rect 14525 17230 14555 17235
rect 14525 17210 14530 17230
rect 14530 17210 14550 17230
rect 14550 17210 14555 17230
rect 14525 17205 14555 17210
rect 14605 17230 14635 17235
rect 14605 17210 14610 17230
rect 14610 17210 14630 17230
rect 14630 17210 14635 17230
rect 14605 17205 14635 17210
rect 14685 17230 14715 17235
rect 14685 17210 14690 17230
rect 14690 17210 14710 17230
rect 14710 17210 14715 17230
rect 14685 17205 14715 17210
rect 16765 17230 16795 17235
rect 16765 17210 16770 17230
rect 16770 17210 16790 17230
rect 16790 17210 16795 17230
rect 16765 17205 16795 17210
rect 16845 17230 16875 17235
rect 16845 17210 16850 17230
rect 16850 17210 16870 17230
rect 16870 17210 16875 17230
rect 16845 17205 16875 17210
rect 16925 17230 16955 17235
rect 16925 17210 16930 17230
rect 16930 17210 16950 17230
rect 16950 17210 16955 17230
rect 16925 17205 16955 17210
rect 17005 17230 17035 17235
rect 17005 17210 17010 17230
rect 17010 17210 17030 17230
rect 17030 17210 17035 17230
rect 17005 17205 17035 17210
rect 17085 17230 17115 17235
rect 17085 17210 17090 17230
rect 17090 17210 17110 17230
rect 17110 17210 17115 17230
rect 17085 17205 17115 17210
rect 17165 17230 17195 17235
rect 17165 17210 17170 17230
rect 17170 17210 17190 17230
rect 17190 17210 17195 17230
rect 17165 17205 17195 17210
rect 17245 17230 17275 17235
rect 17245 17210 17250 17230
rect 17250 17210 17270 17230
rect 17270 17210 17275 17230
rect 17245 17205 17275 17210
rect 17325 17230 17355 17235
rect 17325 17210 17330 17230
rect 17330 17210 17350 17230
rect 17350 17210 17355 17230
rect 17325 17205 17355 17210
rect 17405 17230 17435 17235
rect 17405 17210 17410 17230
rect 17410 17210 17430 17230
rect 17430 17210 17435 17230
rect 17405 17205 17435 17210
rect 17485 17230 17515 17235
rect 17485 17210 17490 17230
rect 17490 17210 17510 17230
rect 17510 17210 17515 17230
rect 17485 17205 17515 17210
rect 17565 17230 17595 17235
rect 17565 17210 17570 17230
rect 17570 17210 17590 17230
rect 17590 17210 17595 17230
rect 17565 17205 17595 17210
rect 17645 17230 17675 17235
rect 17645 17210 17650 17230
rect 17650 17210 17670 17230
rect 17670 17210 17675 17230
rect 17645 17205 17675 17210
rect 17725 17230 17755 17235
rect 17725 17210 17730 17230
rect 17730 17210 17750 17230
rect 17750 17210 17755 17230
rect 17725 17205 17755 17210
rect 17805 17230 17835 17235
rect 17805 17210 17810 17230
rect 17810 17210 17830 17230
rect 17830 17210 17835 17230
rect 17805 17205 17835 17210
rect 17885 17230 17915 17235
rect 17885 17210 17890 17230
rect 17890 17210 17910 17230
rect 17910 17210 17915 17230
rect 17885 17205 17915 17210
rect 17965 17230 17995 17235
rect 17965 17210 17970 17230
rect 17970 17210 17990 17230
rect 17990 17210 17995 17230
rect 17965 17205 17995 17210
rect 18045 17230 18075 17235
rect 18045 17210 18050 17230
rect 18050 17210 18070 17230
rect 18070 17210 18075 17230
rect 18045 17205 18075 17210
rect 18125 17230 18155 17235
rect 18125 17210 18130 17230
rect 18130 17210 18150 17230
rect 18150 17210 18155 17230
rect 18125 17205 18155 17210
rect 18205 17230 18235 17235
rect 18205 17210 18210 17230
rect 18210 17210 18230 17230
rect 18230 17210 18235 17230
rect 18205 17205 18235 17210
rect 18285 17230 18315 17235
rect 18285 17210 18290 17230
rect 18290 17210 18310 17230
rect 18310 17210 18315 17230
rect 18285 17205 18315 17210
rect 18365 17230 18395 17235
rect 18365 17210 18370 17230
rect 18370 17210 18390 17230
rect 18390 17210 18395 17230
rect 18365 17205 18395 17210
rect 18445 17230 18475 17235
rect 18445 17210 18450 17230
rect 18450 17210 18470 17230
rect 18470 17210 18475 17230
rect 18445 17205 18475 17210
rect 18525 17230 18555 17235
rect 18525 17210 18530 17230
rect 18530 17210 18550 17230
rect 18550 17210 18555 17230
rect 18525 17205 18555 17210
rect 18605 17230 18635 17235
rect 18605 17210 18610 17230
rect 18610 17210 18630 17230
rect 18630 17210 18635 17230
rect 18605 17205 18635 17210
rect 18685 17230 18715 17235
rect 18685 17210 18690 17230
rect 18690 17210 18710 17230
rect 18710 17210 18715 17230
rect 18685 17205 18715 17210
rect 18765 17230 18795 17235
rect 18765 17210 18770 17230
rect 18770 17210 18790 17230
rect 18790 17210 18795 17230
rect 18765 17205 18795 17210
rect 18845 17230 18875 17235
rect 18845 17210 18850 17230
rect 18850 17210 18870 17230
rect 18870 17210 18875 17230
rect 18845 17205 18875 17210
rect 18925 17230 18955 17235
rect 18925 17210 18930 17230
rect 18930 17210 18950 17230
rect 18950 17210 18955 17230
rect 18925 17205 18955 17210
rect 19005 17230 19035 17235
rect 19005 17210 19010 17230
rect 19010 17210 19030 17230
rect 19030 17210 19035 17230
rect 19005 17205 19035 17210
rect 19085 17230 19115 17235
rect 19085 17210 19090 17230
rect 19090 17210 19110 17230
rect 19110 17210 19115 17230
rect 19085 17205 19115 17210
rect 19165 17230 19195 17235
rect 19165 17210 19170 17230
rect 19170 17210 19190 17230
rect 19190 17210 19195 17230
rect 19165 17205 19195 17210
rect 19245 17230 19275 17235
rect 19245 17210 19250 17230
rect 19250 17210 19270 17230
rect 19270 17210 19275 17230
rect 19245 17205 19275 17210
rect 19325 17230 19355 17235
rect 19325 17210 19330 17230
rect 19330 17210 19350 17230
rect 19350 17210 19355 17230
rect 19325 17205 19355 17210
rect 19405 17230 19435 17235
rect 19405 17210 19410 17230
rect 19410 17210 19430 17230
rect 19430 17210 19435 17230
rect 19405 17205 19435 17210
rect 19485 17230 19515 17235
rect 19485 17210 19490 17230
rect 19490 17210 19510 17230
rect 19510 17210 19515 17230
rect 19485 17205 19515 17210
rect 19565 17230 19595 17235
rect 19565 17210 19570 17230
rect 19570 17210 19590 17230
rect 19590 17210 19595 17230
rect 19565 17205 19595 17210
rect 19645 17230 19675 17235
rect 19645 17210 19650 17230
rect 19650 17210 19670 17230
rect 19670 17210 19675 17230
rect 19645 17205 19675 17210
rect 19725 17230 19755 17235
rect 19725 17210 19730 17230
rect 19730 17210 19750 17230
rect 19750 17210 19755 17230
rect 19725 17205 19755 17210
rect 19805 17230 19835 17235
rect 19805 17210 19810 17230
rect 19810 17210 19830 17230
rect 19830 17210 19835 17230
rect 19805 17205 19835 17210
rect 19885 17230 19915 17235
rect 19885 17210 19890 17230
rect 19890 17210 19910 17230
rect 19910 17210 19915 17230
rect 19885 17205 19915 17210
rect 19965 17230 19995 17235
rect 19965 17210 19970 17230
rect 19970 17210 19990 17230
rect 19990 17210 19995 17230
rect 19965 17205 19995 17210
rect 20045 17230 20075 17235
rect 20045 17210 20050 17230
rect 20050 17210 20070 17230
rect 20070 17210 20075 17230
rect 20045 17205 20075 17210
rect 20125 17230 20155 17235
rect 20125 17210 20130 17230
rect 20130 17210 20150 17230
rect 20150 17210 20155 17230
rect 20125 17205 20155 17210
rect 20205 17230 20235 17235
rect 20205 17210 20210 17230
rect 20210 17210 20230 17230
rect 20230 17210 20235 17230
rect 20205 17205 20235 17210
rect 20285 17230 20315 17235
rect 20285 17210 20290 17230
rect 20290 17210 20310 17230
rect 20310 17210 20315 17230
rect 20285 17205 20315 17210
rect 20365 17230 20395 17235
rect 20365 17210 20370 17230
rect 20370 17210 20390 17230
rect 20390 17210 20395 17230
rect 20365 17205 20395 17210
rect 20445 17230 20475 17235
rect 20445 17210 20450 17230
rect 20450 17210 20470 17230
rect 20470 17210 20475 17230
rect 20445 17205 20475 17210
rect 20525 17230 20555 17235
rect 20525 17210 20530 17230
rect 20530 17210 20550 17230
rect 20550 17210 20555 17230
rect 20525 17205 20555 17210
rect 20605 17230 20635 17235
rect 20605 17210 20610 17230
rect 20610 17210 20630 17230
rect 20630 17210 20635 17230
rect 20605 17205 20635 17210
rect 20685 17230 20715 17235
rect 20685 17210 20690 17230
rect 20690 17210 20710 17230
rect 20710 17210 20715 17230
rect 20685 17205 20715 17210
rect 20765 17230 20795 17235
rect 20765 17210 20770 17230
rect 20770 17210 20790 17230
rect 20790 17210 20795 17230
rect 20765 17205 20795 17210
rect 20845 17230 20875 17235
rect 20845 17210 20850 17230
rect 20850 17210 20870 17230
rect 20870 17210 20875 17230
rect 20845 17205 20875 17210
rect 20925 17230 20955 17235
rect 20925 17210 20930 17230
rect 20930 17210 20950 17230
rect 20950 17210 20955 17230
rect 20925 17205 20955 17210
rect 5 17150 35 17155
rect 5 17130 10 17150
rect 10 17130 30 17150
rect 30 17130 35 17150
rect 5 17125 35 17130
rect 85 17150 115 17155
rect 85 17130 90 17150
rect 90 17130 110 17150
rect 110 17130 115 17150
rect 85 17125 115 17130
rect 165 17150 195 17155
rect 165 17130 170 17150
rect 170 17130 190 17150
rect 190 17130 195 17150
rect 165 17125 195 17130
rect 245 17150 275 17155
rect 245 17130 250 17150
rect 250 17130 270 17150
rect 270 17130 275 17150
rect 245 17125 275 17130
rect 325 17150 355 17155
rect 325 17130 330 17150
rect 330 17130 350 17150
rect 350 17130 355 17150
rect 325 17125 355 17130
rect 405 17150 435 17155
rect 405 17130 410 17150
rect 410 17130 430 17150
rect 430 17130 435 17150
rect 405 17125 435 17130
rect 485 17150 515 17155
rect 485 17130 490 17150
rect 490 17130 510 17150
rect 510 17130 515 17150
rect 485 17125 515 17130
rect 565 17150 595 17155
rect 565 17130 570 17150
rect 570 17130 590 17150
rect 590 17130 595 17150
rect 565 17125 595 17130
rect 645 17150 675 17155
rect 645 17130 650 17150
rect 650 17130 670 17150
rect 670 17130 675 17150
rect 645 17125 675 17130
rect 725 17150 755 17155
rect 725 17130 730 17150
rect 730 17130 750 17150
rect 750 17130 755 17150
rect 725 17125 755 17130
rect 805 17150 835 17155
rect 805 17130 810 17150
rect 810 17130 830 17150
rect 830 17130 835 17150
rect 805 17125 835 17130
rect 885 17150 915 17155
rect 885 17130 890 17150
rect 890 17130 910 17150
rect 910 17130 915 17150
rect 885 17125 915 17130
rect 965 17150 995 17155
rect 965 17130 970 17150
rect 970 17130 990 17150
rect 990 17130 995 17150
rect 965 17125 995 17130
rect 1045 17150 1075 17155
rect 1045 17130 1050 17150
rect 1050 17130 1070 17150
rect 1070 17130 1075 17150
rect 1045 17125 1075 17130
rect 1125 17150 1155 17155
rect 1125 17130 1130 17150
rect 1130 17130 1150 17150
rect 1150 17130 1155 17150
rect 1125 17125 1155 17130
rect 1205 17150 1235 17155
rect 1205 17130 1210 17150
rect 1210 17130 1230 17150
rect 1230 17130 1235 17150
rect 1205 17125 1235 17130
rect 1285 17150 1315 17155
rect 1285 17130 1290 17150
rect 1290 17130 1310 17150
rect 1310 17130 1315 17150
rect 1285 17125 1315 17130
rect 1365 17150 1395 17155
rect 1365 17130 1370 17150
rect 1370 17130 1390 17150
rect 1390 17130 1395 17150
rect 1365 17125 1395 17130
rect 1445 17150 1475 17155
rect 1445 17130 1450 17150
rect 1450 17130 1470 17150
rect 1470 17130 1475 17150
rect 1445 17125 1475 17130
rect 1525 17150 1555 17155
rect 1525 17130 1530 17150
rect 1530 17130 1550 17150
rect 1550 17130 1555 17150
rect 1525 17125 1555 17130
rect 1605 17150 1635 17155
rect 1605 17130 1610 17150
rect 1610 17130 1630 17150
rect 1630 17130 1635 17150
rect 1605 17125 1635 17130
rect 1685 17150 1715 17155
rect 1685 17130 1690 17150
rect 1690 17130 1710 17150
rect 1710 17130 1715 17150
rect 1685 17125 1715 17130
rect 1765 17150 1795 17155
rect 1765 17130 1770 17150
rect 1770 17130 1790 17150
rect 1790 17130 1795 17150
rect 1765 17125 1795 17130
rect 1845 17150 1875 17155
rect 1845 17130 1850 17150
rect 1850 17130 1870 17150
rect 1870 17130 1875 17150
rect 1845 17125 1875 17130
rect 1925 17150 1955 17155
rect 1925 17130 1930 17150
rect 1930 17130 1950 17150
rect 1950 17130 1955 17150
rect 1925 17125 1955 17130
rect 2005 17150 2035 17155
rect 2005 17130 2010 17150
rect 2010 17130 2030 17150
rect 2030 17130 2035 17150
rect 2005 17125 2035 17130
rect 2085 17150 2115 17155
rect 2085 17130 2090 17150
rect 2090 17130 2110 17150
rect 2110 17130 2115 17150
rect 2085 17125 2115 17130
rect 2165 17150 2195 17155
rect 2165 17130 2170 17150
rect 2170 17130 2190 17150
rect 2190 17130 2195 17150
rect 2165 17125 2195 17130
rect 2245 17150 2275 17155
rect 2245 17130 2250 17150
rect 2250 17130 2270 17150
rect 2270 17130 2275 17150
rect 2245 17125 2275 17130
rect 2325 17150 2355 17155
rect 2325 17130 2330 17150
rect 2330 17130 2350 17150
rect 2350 17130 2355 17150
rect 2325 17125 2355 17130
rect 2405 17150 2435 17155
rect 2405 17130 2410 17150
rect 2410 17130 2430 17150
rect 2430 17130 2435 17150
rect 2405 17125 2435 17130
rect 2485 17150 2515 17155
rect 2485 17130 2490 17150
rect 2490 17130 2510 17150
rect 2510 17130 2515 17150
rect 2485 17125 2515 17130
rect 2565 17150 2595 17155
rect 2565 17130 2570 17150
rect 2570 17130 2590 17150
rect 2590 17130 2595 17150
rect 2565 17125 2595 17130
rect 2645 17150 2675 17155
rect 2645 17130 2650 17150
rect 2650 17130 2670 17150
rect 2670 17130 2675 17150
rect 2645 17125 2675 17130
rect 2725 17150 2755 17155
rect 2725 17130 2730 17150
rect 2730 17130 2750 17150
rect 2750 17130 2755 17150
rect 2725 17125 2755 17130
rect 2805 17150 2835 17155
rect 2805 17130 2810 17150
rect 2810 17130 2830 17150
rect 2830 17130 2835 17150
rect 2805 17125 2835 17130
rect 2885 17150 2915 17155
rect 2885 17130 2890 17150
rect 2890 17130 2910 17150
rect 2910 17130 2915 17150
rect 2885 17125 2915 17130
rect 2965 17150 2995 17155
rect 2965 17130 2970 17150
rect 2970 17130 2990 17150
rect 2990 17130 2995 17150
rect 2965 17125 2995 17130
rect 3045 17150 3075 17155
rect 3045 17130 3050 17150
rect 3050 17130 3070 17150
rect 3070 17130 3075 17150
rect 3045 17125 3075 17130
rect 3125 17150 3155 17155
rect 3125 17130 3130 17150
rect 3130 17130 3150 17150
rect 3150 17130 3155 17150
rect 3125 17125 3155 17130
rect 3205 17150 3235 17155
rect 3205 17130 3210 17150
rect 3210 17130 3230 17150
rect 3230 17130 3235 17150
rect 3205 17125 3235 17130
rect 3285 17150 3315 17155
rect 3285 17130 3290 17150
rect 3290 17130 3310 17150
rect 3310 17130 3315 17150
rect 3285 17125 3315 17130
rect 3365 17150 3395 17155
rect 3365 17130 3370 17150
rect 3370 17130 3390 17150
rect 3390 17130 3395 17150
rect 3365 17125 3395 17130
rect 3445 17150 3475 17155
rect 3445 17130 3450 17150
rect 3450 17130 3470 17150
rect 3470 17130 3475 17150
rect 3445 17125 3475 17130
rect 3525 17150 3555 17155
rect 3525 17130 3530 17150
rect 3530 17130 3550 17150
rect 3550 17130 3555 17150
rect 3525 17125 3555 17130
rect 3605 17150 3635 17155
rect 3605 17130 3610 17150
rect 3610 17130 3630 17150
rect 3630 17130 3635 17150
rect 3605 17125 3635 17130
rect 3685 17150 3715 17155
rect 3685 17130 3690 17150
rect 3690 17130 3710 17150
rect 3710 17130 3715 17150
rect 3685 17125 3715 17130
rect 3765 17150 3795 17155
rect 3765 17130 3770 17150
rect 3770 17130 3790 17150
rect 3790 17130 3795 17150
rect 3765 17125 3795 17130
rect 3845 17150 3875 17155
rect 3845 17130 3850 17150
rect 3850 17130 3870 17150
rect 3870 17130 3875 17150
rect 3845 17125 3875 17130
rect 3925 17150 3955 17155
rect 3925 17130 3930 17150
rect 3930 17130 3950 17150
rect 3950 17130 3955 17150
rect 3925 17125 3955 17130
rect 4005 17150 4035 17155
rect 4005 17130 4010 17150
rect 4010 17130 4030 17150
rect 4030 17130 4035 17150
rect 4005 17125 4035 17130
rect 4085 17150 4115 17155
rect 4085 17130 4090 17150
rect 4090 17130 4110 17150
rect 4110 17130 4115 17150
rect 4085 17125 4115 17130
rect 4165 17150 4195 17155
rect 4165 17130 4170 17150
rect 4170 17130 4190 17150
rect 4190 17130 4195 17150
rect 4165 17125 4195 17130
rect 6245 17150 6275 17155
rect 6245 17130 6250 17150
rect 6250 17130 6270 17150
rect 6270 17130 6275 17150
rect 6245 17125 6275 17130
rect 6325 17150 6355 17155
rect 6325 17130 6330 17150
rect 6330 17130 6350 17150
rect 6350 17130 6355 17150
rect 6325 17125 6355 17130
rect 6405 17150 6435 17155
rect 6405 17130 6410 17150
rect 6410 17130 6430 17150
rect 6430 17130 6435 17150
rect 6405 17125 6435 17130
rect 6485 17150 6515 17155
rect 6485 17130 6490 17150
rect 6490 17130 6510 17150
rect 6510 17130 6515 17150
rect 6485 17125 6515 17130
rect 6565 17150 6595 17155
rect 6565 17130 6570 17150
rect 6570 17130 6590 17150
rect 6590 17130 6595 17150
rect 6565 17125 6595 17130
rect 6645 17150 6675 17155
rect 6645 17130 6650 17150
rect 6650 17130 6670 17150
rect 6670 17130 6675 17150
rect 6645 17125 6675 17130
rect 6725 17150 6755 17155
rect 6725 17130 6730 17150
rect 6730 17130 6750 17150
rect 6750 17130 6755 17150
rect 6725 17125 6755 17130
rect 6805 17150 6835 17155
rect 6805 17130 6810 17150
rect 6810 17130 6830 17150
rect 6830 17130 6835 17150
rect 6805 17125 6835 17130
rect 6885 17150 6915 17155
rect 6885 17130 6890 17150
rect 6890 17130 6910 17150
rect 6910 17130 6915 17150
rect 6885 17125 6915 17130
rect 6965 17150 6995 17155
rect 6965 17130 6970 17150
rect 6970 17130 6990 17150
rect 6990 17130 6995 17150
rect 6965 17125 6995 17130
rect 7045 17150 7075 17155
rect 7045 17130 7050 17150
rect 7050 17130 7070 17150
rect 7070 17130 7075 17150
rect 7045 17125 7075 17130
rect 7125 17150 7155 17155
rect 7125 17130 7130 17150
rect 7130 17130 7150 17150
rect 7150 17130 7155 17150
rect 7125 17125 7155 17130
rect 7205 17150 7235 17155
rect 7205 17130 7210 17150
rect 7210 17130 7230 17150
rect 7230 17130 7235 17150
rect 7205 17125 7235 17130
rect 7285 17150 7315 17155
rect 7285 17130 7290 17150
rect 7290 17130 7310 17150
rect 7310 17130 7315 17150
rect 7285 17125 7315 17130
rect 7365 17150 7395 17155
rect 7365 17130 7370 17150
rect 7370 17130 7390 17150
rect 7390 17130 7395 17150
rect 7365 17125 7395 17130
rect 7445 17150 7475 17155
rect 7445 17130 7450 17150
rect 7450 17130 7470 17150
rect 7470 17130 7475 17150
rect 7445 17125 7475 17130
rect 7525 17150 7555 17155
rect 7525 17130 7530 17150
rect 7530 17130 7550 17150
rect 7550 17130 7555 17150
rect 7525 17125 7555 17130
rect 7605 17150 7635 17155
rect 7605 17130 7610 17150
rect 7610 17130 7630 17150
rect 7630 17130 7635 17150
rect 7605 17125 7635 17130
rect 7685 17150 7715 17155
rect 7685 17130 7690 17150
rect 7690 17130 7710 17150
rect 7710 17130 7715 17150
rect 7685 17125 7715 17130
rect 7765 17150 7795 17155
rect 7765 17130 7770 17150
rect 7770 17130 7790 17150
rect 7790 17130 7795 17150
rect 7765 17125 7795 17130
rect 7845 17150 7875 17155
rect 7845 17130 7850 17150
rect 7850 17130 7870 17150
rect 7870 17130 7875 17150
rect 7845 17125 7875 17130
rect 7925 17150 7955 17155
rect 7925 17130 7930 17150
rect 7930 17130 7950 17150
rect 7950 17130 7955 17150
rect 7925 17125 7955 17130
rect 8005 17150 8035 17155
rect 8005 17130 8010 17150
rect 8010 17130 8030 17150
rect 8030 17130 8035 17150
rect 8005 17125 8035 17130
rect 8085 17150 8115 17155
rect 8085 17130 8090 17150
rect 8090 17130 8110 17150
rect 8110 17130 8115 17150
rect 8085 17125 8115 17130
rect 8165 17150 8195 17155
rect 8165 17130 8170 17150
rect 8170 17130 8190 17150
rect 8190 17130 8195 17150
rect 8165 17125 8195 17130
rect 8245 17150 8275 17155
rect 8245 17130 8250 17150
rect 8250 17130 8270 17150
rect 8270 17130 8275 17150
rect 8245 17125 8275 17130
rect 8325 17150 8355 17155
rect 8325 17130 8330 17150
rect 8330 17130 8350 17150
rect 8350 17130 8355 17150
rect 8325 17125 8355 17130
rect 8405 17150 8435 17155
rect 8405 17130 8410 17150
rect 8410 17130 8430 17150
rect 8430 17130 8435 17150
rect 8405 17125 8435 17130
rect 8485 17150 8515 17155
rect 8485 17130 8490 17150
rect 8490 17130 8510 17150
rect 8510 17130 8515 17150
rect 8485 17125 8515 17130
rect 8565 17150 8595 17155
rect 8565 17130 8570 17150
rect 8570 17130 8590 17150
rect 8590 17130 8595 17150
rect 8565 17125 8595 17130
rect 8645 17150 8675 17155
rect 8645 17130 8650 17150
rect 8650 17130 8670 17150
rect 8670 17130 8675 17150
rect 8645 17125 8675 17130
rect 8725 17150 8755 17155
rect 8725 17130 8730 17150
rect 8730 17130 8750 17150
rect 8750 17130 8755 17150
rect 8725 17125 8755 17130
rect 8805 17150 8835 17155
rect 8805 17130 8810 17150
rect 8810 17130 8830 17150
rect 8830 17130 8835 17150
rect 8805 17125 8835 17130
rect 8885 17150 8915 17155
rect 8885 17130 8890 17150
rect 8890 17130 8910 17150
rect 8910 17130 8915 17150
rect 8885 17125 8915 17130
rect 8965 17150 8995 17155
rect 8965 17130 8970 17150
rect 8970 17130 8990 17150
rect 8990 17130 8995 17150
rect 8965 17125 8995 17130
rect 9045 17150 9075 17155
rect 9045 17130 9050 17150
rect 9050 17130 9070 17150
rect 9070 17130 9075 17150
rect 9045 17125 9075 17130
rect 9125 17150 9155 17155
rect 9125 17130 9130 17150
rect 9130 17130 9150 17150
rect 9150 17130 9155 17150
rect 9125 17125 9155 17130
rect 9205 17150 9235 17155
rect 9205 17130 9210 17150
rect 9210 17130 9230 17150
rect 9230 17130 9235 17150
rect 9205 17125 9235 17130
rect 9285 17150 9315 17155
rect 9285 17130 9290 17150
rect 9290 17130 9310 17150
rect 9310 17130 9315 17150
rect 9285 17125 9315 17130
rect 9365 17150 9395 17155
rect 9365 17130 9370 17150
rect 9370 17130 9390 17150
rect 9390 17130 9395 17150
rect 9365 17125 9395 17130
rect 9445 17150 9475 17155
rect 9445 17130 9450 17150
rect 9450 17130 9470 17150
rect 9470 17130 9475 17150
rect 9445 17125 9475 17130
rect 11565 17150 11595 17155
rect 11565 17130 11570 17150
rect 11570 17130 11590 17150
rect 11590 17130 11595 17150
rect 11565 17125 11595 17130
rect 11645 17150 11675 17155
rect 11645 17130 11650 17150
rect 11650 17130 11670 17150
rect 11670 17130 11675 17150
rect 11645 17125 11675 17130
rect 11725 17150 11755 17155
rect 11725 17130 11730 17150
rect 11730 17130 11750 17150
rect 11750 17130 11755 17150
rect 11725 17125 11755 17130
rect 11805 17150 11835 17155
rect 11805 17130 11810 17150
rect 11810 17130 11830 17150
rect 11830 17130 11835 17150
rect 11805 17125 11835 17130
rect 11885 17150 11915 17155
rect 11885 17130 11890 17150
rect 11890 17130 11910 17150
rect 11910 17130 11915 17150
rect 11885 17125 11915 17130
rect 11965 17150 11995 17155
rect 11965 17130 11970 17150
rect 11970 17130 11990 17150
rect 11990 17130 11995 17150
rect 11965 17125 11995 17130
rect 12045 17150 12075 17155
rect 12045 17130 12050 17150
rect 12050 17130 12070 17150
rect 12070 17130 12075 17150
rect 12045 17125 12075 17130
rect 12125 17150 12155 17155
rect 12125 17130 12130 17150
rect 12130 17130 12150 17150
rect 12150 17130 12155 17150
rect 12125 17125 12155 17130
rect 12205 17150 12235 17155
rect 12205 17130 12210 17150
rect 12210 17130 12230 17150
rect 12230 17130 12235 17150
rect 12205 17125 12235 17130
rect 12285 17150 12315 17155
rect 12285 17130 12290 17150
rect 12290 17130 12310 17150
rect 12310 17130 12315 17150
rect 12285 17125 12315 17130
rect 12365 17150 12395 17155
rect 12365 17130 12370 17150
rect 12370 17130 12390 17150
rect 12390 17130 12395 17150
rect 12365 17125 12395 17130
rect 12445 17150 12475 17155
rect 12445 17130 12450 17150
rect 12450 17130 12470 17150
rect 12470 17130 12475 17150
rect 12445 17125 12475 17130
rect 12525 17150 12555 17155
rect 12525 17130 12530 17150
rect 12530 17130 12550 17150
rect 12550 17130 12555 17150
rect 12525 17125 12555 17130
rect 12605 17150 12635 17155
rect 12605 17130 12610 17150
rect 12610 17130 12630 17150
rect 12630 17130 12635 17150
rect 12605 17125 12635 17130
rect 12685 17150 12715 17155
rect 12685 17130 12690 17150
rect 12690 17130 12710 17150
rect 12710 17130 12715 17150
rect 12685 17125 12715 17130
rect 12765 17150 12795 17155
rect 12765 17130 12770 17150
rect 12770 17130 12790 17150
rect 12790 17130 12795 17150
rect 12765 17125 12795 17130
rect 12845 17150 12875 17155
rect 12845 17130 12850 17150
rect 12850 17130 12870 17150
rect 12870 17130 12875 17150
rect 12845 17125 12875 17130
rect 12925 17150 12955 17155
rect 12925 17130 12930 17150
rect 12930 17130 12950 17150
rect 12950 17130 12955 17150
rect 12925 17125 12955 17130
rect 13005 17150 13035 17155
rect 13005 17130 13010 17150
rect 13010 17130 13030 17150
rect 13030 17130 13035 17150
rect 13005 17125 13035 17130
rect 13085 17150 13115 17155
rect 13085 17130 13090 17150
rect 13090 17130 13110 17150
rect 13110 17130 13115 17150
rect 13085 17125 13115 17130
rect 13165 17150 13195 17155
rect 13165 17130 13170 17150
rect 13170 17130 13190 17150
rect 13190 17130 13195 17150
rect 13165 17125 13195 17130
rect 13245 17150 13275 17155
rect 13245 17130 13250 17150
rect 13250 17130 13270 17150
rect 13270 17130 13275 17150
rect 13245 17125 13275 17130
rect 13325 17150 13355 17155
rect 13325 17130 13330 17150
rect 13330 17130 13350 17150
rect 13350 17130 13355 17150
rect 13325 17125 13355 17130
rect 13405 17150 13435 17155
rect 13405 17130 13410 17150
rect 13410 17130 13430 17150
rect 13430 17130 13435 17150
rect 13405 17125 13435 17130
rect 13485 17150 13515 17155
rect 13485 17130 13490 17150
rect 13490 17130 13510 17150
rect 13510 17130 13515 17150
rect 13485 17125 13515 17130
rect 13565 17150 13595 17155
rect 13565 17130 13570 17150
rect 13570 17130 13590 17150
rect 13590 17130 13595 17150
rect 13565 17125 13595 17130
rect 13645 17150 13675 17155
rect 13645 17130 13650 17150
rect 13650 17130 13670 17150
rect 13670 17130 13675 17150
rect 13645 17125 13675 17130
rect 13725 17150 13755 17155
rect 13725 17130 13730 17150
rect 13730 17130 13750 17150
rect 13750 17130 13755 17150
rect 13725 17125 13755 17130
rect 13805 17150 13835 17155
rect 13805 17130 13810 17150
rect 13810 17130 13830 17150
rect 13830 17130 13835 17150
rect 13805 17125 13835 17130
rect 13885 17150 13915 17155
rect 13885 17130 13890 17150
rect 13890 17130 13910 17150
rect 13910 17130 13915 17150
rect 13885 17125 13915 17130
rect 13965 17150 13995 17155
rect 13965 17130 13970 17150
rect 13970 17130 13990 17150
rect 13990 17130 13995 17150
rect 13965 17125 13995 17130
rect 14045 17150 14075 17155
rect 14045 17130 14050 17150
rect 14050 17130 14070 17150
rect 14070 17130 14075 17150
rect 14045 17125 14075 17130
rect 14125 17150 14155 17155
rect 14125 17130 14130 17150
rect 14130 17130 14150 17150
rect 14150 17130 14155 17150
rect 14125 17125 14155 17130
rect 14205 17150 14235 17155
rect 14205 17130 14210 17150
rect 14210 17130 14230 17150
rect 14230 17130 14235 17150
rect 14205 17125 14235 17130
rect 14285 17150 14315 17155
rect 14285 17130 14290 17150
rect 14290 17130 14310 17150
rect 14310 17130 14315 17150
rect 14285 17125 14315 17130
rect 14365 17150 14395 17155
rect 14365 17130 14370 17150
rect 14370 17130 14390 17150
rect 14390 17130 14395 17150
rect 14365 17125 14395 17130
rect 14445 17150 14475 17155
rect 14445 17130 14450 17150
rect 14450 17130 14470 17150
rect 14470 17130 14475 17150
rect 14445 17125 14475 17130
rect 14525 17150 14555 17155
rect 14525 17130 14530 17150
rect 14530 17130 14550 17150
rect 14550 17130 14555 17150
rect 14525 17125 14555 17130
rect 14605 17150 14635 17155
rect 14605 17130 14610 17150
rect 14610 17130 14630 17150
rect 14630 17130 14635 17150
rect 14605 17125 14635 17130
rect 14685 17150 14715 17155
rect 14685 17130 14690 17150
rect 14690 17130 14710 17150
rect 14710 17130 14715 17150
rect 14685 17125 14715 17130
rect 16765 17150 16795 17155
rect 16765 17130 16770 17150
rect 16770 17130 16790 17150
rect 16790 17130 16795 17150
rect 16765 17125 16795 17130
rect 16845 17150 16875 17155
rect 16845 17130 16850 17150
rect 16850 17130 16870 17150
rect 16870 17130 16875 17150
rect 16845 17125 16875 17130
rect 16925 17150 16955 17155
rect 16925 17130 16930 17150
rect 16930 17130 16950 17150
rect 16950 17130 16955 17150
rect 16925 17125 16955 17130
rect 17005 17150 17035 17155
rect 17005 17130 17010 17150
rect 17010 17130 17030 17150
rect 17030 17130 17035 17150
rect 17005 17125 17035 17130
rect 17085 17150 17115 17155
rect 17085 17130 17090 17150
rect 17090 17130 17110 17150
rect 17110 17130 17115 17150
rect 17085 17125 17115 17130
rect 17165 17150 17195 17155
rect 17165 17130 17170 17150
rect 17170 17130 17190 17150
rect 17190 17130 17195 17150
rect 17165 17125 17195 17130
rect 17245 17150 17275 17155
rect 17245 17130 17250 17150
rect 17250 17130 17270 17150
rect 17270 17130 17275 17150
rect 17245 17125 17275 17130
rect 17325 17150 17355 17155
rect 17325 17130 17330 17150
rect 17330 17130 17350 17150
rect 17350 17130 17355 17150
rect 17325 17125 17355 17130
rect 17405 17150 17435 17155
rect 17405 17130 17410 17150
rect 17410 17130 17430 17150
rect 17430 17130 17435 17150
rect 17405 17125 17435 17130
rect 17485 17150 17515 17155
rect 17485 17130 17490 17150
rect 17490 17130 17510 17150
rect 17510 17130 17515 17150
rect 17485 17125 17515 17130
rect 17565 17150 17595 17155
rect 17565 17130 17570 17150
rect 17570 17130 17590 17150
rect 17590 17130 17595 17150
rect 17565 17125 17595 17130
rect 17645 17150 17675 17155
rect 17645 17130 17650 17150
rect 17650 17130 17670 17150
rect 17670 17130 17675 17150
rect 17645 17125 17675 17130
rect 17725 17150 17755 17155
rect 17725 17130 17730 17150
rect 17730 17130 17750 17150
rect 17750 17130 17755 17150
rect 17725 17125 17755 17130
rect 17805 17150 17835 17155
rect 17805 17130 17810 17150
rect 17810 17130 17830 17150
rect 17830 17130 17835 17150
rect 17805 17125 17835 17130
rect 17885 17150 17915 17155
rect 17885 17130 17890 17150
rect 17890 17130 17910 17150
rect 17910 17130 17915 17150
rect 17885 17125 17915 17130
rect 17965 17150 17995 17155
rect 17965 17130 17970 17150
rect 17970 17130 17990 17150
rect 17990 17130 17995 17150
rect 17965 17125 17995 17130
rect 18045 17150 18075 17155
rect 18045 17130 18050 17150
rect 18050 17130 18070 17150
rect 18070 17130 18075 17150
rect 18045 17125 18075 17130
rect 18125 17150 18155 17155
rect 18125 17130 18130 17150
rect 18130 17130 18150 17150
rect 18150 17130 18155 17150
rect 18125 17125 18155 17130
rect 18205 17150 18235 17155
rect 18205 17130 18210 17150
rect 18210 17130 18230 17150
rect 18230 17130 18235 17150
rect 18205 17125 18235 17130
rect 18285 17150 18315 17155
rect 18285 17130 18290 17150
rect 18290 17130 18310 17150
rect 18310 17130 18315 17150
rect 18285 17125 18315 17130
rect 18365 17150 18395 17155
rect 18365 17130 18370 17150
rect 18370 17130 18390 17150
rect 18390 17130 18395 17150
rect 18365 17125 18395 17130
rect 18445 17150 18475 17155
rect 18445 17130 18450 17150
rect 18450 17130 18470 17150
rect 18470 17130 18475 17150
rect 18445 17125 18475 17130
rect 18525 17150 18555 17155
rect 18525 17130 18530 17150
rect 18530 17130 18550 17150
rect 18550 17130 18555 17150
rect 18525 17125 18555 17130
rect 18605 17150 18635 17155
rect 18605 17130 18610 17150
rect 18610 17130 18630 17150
rect 18630 17130 18635 17150
rect 18605 17125 18635 17130
rect 18685 17150 18715 17155
rect 18685 17130 18690 17150
rect 18690 17130 18710 17150
rect 18710 17130 18715 17150
rect 18685 17125 18715 17130
rect 18765 17150 18795 17155
rect 18765 17130 18770 17150
rect 18770 17130 18790 17150
rect 18790 17130 18795 17150
rect 18765 17125 18795 17130
rect 18845 17150 18875 17155
rect 18845 17130 18850 17150
rect 18850 17130 18870 17150
rect 18870 17130 18875 17150
rect 18845 17125 18875 17130
rect 18925 17150 18955 17155
rect 18925 17130 18930 17150
rect 18930 17130 18950 17150
rect 18950 17130 18955 17150
rect 18925 17125 18955 17130
rect 19005 17150 19035 17155
rect 19005 17130 19010 17150
rect 19010 17130 19030 17150
rect 19030 17130 19035 17150
rect 19005 17125 19035 17130
rect 19085 17150 19115 17155
rect 19085 17130 19090 17150
rect 19090 17130 19110 17150
rect 19110 17130 19115 17150
rect 19085 17125 19115 17130
rect 19165 17150 19195 17155
rect 19165 17130 19170 17150
rect 19170 17130 19190 17150
rect 19190 17130 19195 17150
rect 19165 17125 19195 17130
rect 19245 17150 19275 17155
rect 19245 17130 19250 17150
rect 19250 17130 19270 17150
rect 19270 17130 19275 17150
rect 19245 17125 19275 17130
rect 19325 17150 19355 17155
rect 19325 17130 19330 17150
rect 19330 17130 19350 17150
rect 19350 17130 19355 17150
rect 19325 17125 19355 17130
rect 19405 17150 19435 17155
rect 19405 17130 19410 17150
rect 19410 17130 19430 17150
rect 19430 17130 19435 17150
rect 19405 17125 19435 17130
rect 19485 17150 19515 17155
rect 19485 17130 19490 17150
rect 19490 17130 19510 17150
rect 19510 17130 19515 17150
rect 19485 17125 19515 17130
rect 19565 17150 19595 17155
rect 19565 17130 19570 17150
rect 19570 17130 19590 17150
rect 19590 17130 19595 17150
rect 19565 17125 19595 17130
rect 19645 17150 19675 17155
rect 19645 17130 19650 17150
rect 19650 17130 19670 17150
rect 19670 17130 19675 17150
rect 19645 17125 19675 17130
rect 19725 17150 19755 17155
rect 19725 17130 19730 17150
rect 19730 17130 19750 17150
rect 19750 17130 19755 17150
rect 19725 17125 19755 17130
rect 19805 17150 19835 17155
rect 19805 17130 19810 17150
rect 19810 17130 19830 17150
rect 19830 17130 19835 17150
rect 19805 17125 19835 17130
rect 19885 17150 19915 17155
rect 19885 17130 19890 17150
rect 19890 17130 19910 17150
rect 19910 17130 19915 17150
rect 19885 17125 19915 17130
rect 19965 17150 19995 17155
rect 19965 17130 19970 17150
rect 19970 17130 19990 17150
rect 19990 17130 19995 17150
rect 19965 17125 19995 17130
rect 20045 17150 20075 17155
rect 20045 17130 20050 17150
rect 20050 17130 20070 17150
rect 20070 17130 20075 17150
rect 20045 17125 20075 17130
rect 20125 17150 20155 17155
rect 20125 17130 20130 17150
rect 20130 17130 20150 17150
rect 20150 17130 20155 17150
rect 20125 17125 20155 17130
rect 20205 17150 20235 17155
rect 20205 17130 20210 17150
rect 20210 17130 20230 17150
rect 20230 17130 20235 17150
rect 20205 17125 20235 17130
rect 20285 17150 20315 17155
rect 20285 17130 20290 17150
rect 20290 17130 20310 17150
rect 20310 17130 20315 17150
rect 20285 17125 20315 17130
rect 20365 17150 20395 17155
rect 20365 17130 20370 17150
rect 20370 17130 20390 17150
rect 20390 17130 20395 17150
rect 20365 17125 20395 17130
rect 20445 17150 20475 17155
rect 20445 17130 20450 17150
rect 20450 17130 20470 17150
rect 20470 17130 20475 17150
rect 20445 17125 20475 17130
rect 20525 17150 20555 17155
rect 20525 17130 20530 17150
rect 20530 17130 20550 17150
rect 20550 17130 20555 17150
rect 20525 17125 20555 17130
rect 20605 17150 20635 17155
rect 20605 17130 20610 17150
rect 20610 17130 20630 17150
rect 20630 17130 20635 17150
rect 20605 17125 20635 17130
rect 20685 17150 20715 17155
rect 20685 17130 20690 17150
rect 20690 17130 20710 17150
rect 20710 17130 20715 17150
rect 20685 17125 20715 17130
rect 20765 17150 20795 17155
rect 20765 17130 20770 17150
rect 20770 17130 20790 17150
rect 20790 17130 20795 17150
rect 20765 17125 20795 17130
rect 20845 17150 20875 17155
rect 20845 17130 20850 17150
rect 20850 17130 20870 17150
rect 20870 17130 20875 17150
rect 20845 17125 20875 17130
rect 20925 17150 20955 17155
rect 20925 17130 20930 17150
rect 20930 17130 20950 17150
rect 20950 17130 20955 17150
rect 20925 17125 20955 17130
rect 5 16990 35 16995
rect 5 16970 10 16990
rect 10 16970 30 16990
rect 30 16970 35 16990
rect 5 16965 35 16970
rect 85 16990 115 16995
rect 85 16970 90 16990
rect 90 16970 110 16990
rect 110 16970 115 16990
rect 85 16965 115 16970
rect 165 16990 195 16995
rect 165 16970 170 16990
rect 170 16970 190 16990
rect 190 16970 195 16990
rect 165 16965 195 16970
rect 245 16990 275 16995
rect 245 16970 250 16990
rect 250 16970 270 16990
rect 270 16970 275 16990
rect 245 16965 275 16970
rect 325 16990 355 16995
rect 325 16970 330 16990
rect 330 16970 350 16990
rect 350 16970 355 16990
rect 325 16965 355 16970
rect 405 16990 435 16995
rect 405 16970 410 16990
rect 410 16970 430 16990
rect 430 16970 435 16990
rect 405 16965 435 16970
rect 485 16990 515 16995
rect 485 16970 490 16990
rect 490 16970 510 16990
rect 510 16970 515 16990
rect 485 16965 515 16970
rect 565 16990 595 16995
rect 565 16970 570 16990
rect 570 16970 590 16990
rect 590 16970 595 16990
rect 565 16965 595 16970
rect 645 16990 675 16995
rect 645 16970 650 16990
rect 650 16970 670 16990
rect 670 16970 675 16990
rect 645 16965 675 16970
rect 725 16990 755 16995
rect 725 16970 730 16990
rect 730 16970 750 16990
rect 750 16970 755 16990
rect 725 16965 755 16970
rect 805 16990 835 16995
rect 805 16970 810 16990
rect 810 16970 830 16990
rect 830 16970 835 16990
rect 805 16965 835 16970
rect 885 16990 915 16995
rect 885 16970 890 16990
rect 890 16970 910 16990
rect 910 16970 915 16990
rect 885 16965 915 16970
rect 965 16990 995 16995
rect 965 16970 970 16990
rect 970 16970 990 16990
rect 990 16970 995 16990
rect 965 16965 995 16970
rect 1045 16990 1075 16995
rect 1045 16970 1050 16990
rect 1050 16970 1070 16990
rect 1070 16970 1075 16990
rect 1045 16965 1075 16970
rect 1125 16990 1155 16995
rect 1125 16970 1130 16990
rect 1130 16970 1150 16990
rect 1150 16970 1155 16990
rect 1125 16965 1155 16970
rect 1205 16990 1235 16995
rect 1205 16970 1210 16990
rect 1210 16970 1230 16990
rect 1230 16970 1235 16990
rect 1205 16965 1235 16970
rect 1285 16990 1315 16995
rect 1285 16970 1290 16990
rect 1290 16970 1310 16990
rect 1310 16970 1315 16990
rect 1285 16965 1315 16970
rect 1365 16990 1395 16995
rect 1365 16970 1370 16990
rect 1370 16970 1390 16990
rect 1390 16970 1395 16990
rect 1365 16965 1395 16970
rect 1445 16990 1475 16995
rect 1445 16970 1450 16990
rect 1450 16970 1470 16990
rect 1470 16970 1475 16990
rect 1445 16965 1475 16970
rect 1525 16990 1555 16995
rect 1525 16970 1530 16990
rect 1530 16970 1550 16990
rect 1550 16970 1555 16990
rect 1525 16965 1555 16970
rect 1605 16990 1635 16995
rect 1605 16970 1610 16990
rect 1610 16970 1630 16990
rect 1630 16970 1635 16990
rect 1605 16965 1635 16970
rect 1685 16990 1715 16995
rect 1685 16970 1690 16990
rect 1690 16970 1710 16990
rect 1710 16970 1715 16990
rect 1685 16965 1715 16970
rect 1765 16990 1795 16995
rect 1765 16970 1770 16990
rect 1770 16970 1790 16990
rect 1790 16970 1795 16990
rect 1765 16965 1795 16970
rect 1845 16990 1875 16995
rect 1845 16970 1850 16990
rect 1850 16970 1870 16990
rect 1870 16970 1875 16990
rect 1845 16965 1875 16970
rect 1925 16990 1955 16995
rect 1925 16970 1930 16990
rect 1930 16970 1950 16990
rect 1950 16970 1955 16990
rect 1925 16965 1955 16970
rect 2005 16990 2035 16995
rect 2005 16970 2010 16990
rect 2010 16970 2030 16990
rect 2030 16970 2035 16990
rect 2005 16965 2035 16970
rect 2085 16990 2115 16995
rect 2085 16970 2090 16990
rect 2090 16970 2110 16990
rect 2110 16970 2115 16990
rect 2085 16965 2115 16970
rect 2165 16990 2195 16995
rect 2165 16970 2170 16990
rect 2170 16970 2190 16990
rect 2190 16970 2195 16990
rect 2165 16965 2195 16970
rect 2245 16990 2275 16995
rect 2245 16970 2250 16990
rect 2250 16970 2270 16990
rect 2270 16970 2275 16990
rect 2245 16965 2275 16970
rect 2325 16990 2355 16995
rect 2325 16970 2330 16990
rect 2330 16970 2350 16990
rect 2350 16970 2355 16990
rect 2325 16965 2355 16970
rect 2405 16990 2435 16995
rect 2405 16970 2410 16990
rect 2410 16970 2430 16990
rect 2430 16970 2435 16990
rect 2405 16965 2435 16970
rect 2485 16990 2515 16995
rect 2485 16970 2490 16990
rect 2490 16970 2510 16990
rect 2510 16970 2515 16990
rect 2485 16965 2515 16970
rect 2565 16990 2595 16995
rect 2565 16970 2570 16990
rect 2570 16970 2590 16990
rect 2590 16970 2595 16990
rect 2565 16965 2595 16970
rect 2645 16990 2675 16995
rect 2645 16970 2650 16990
rect 2650 16970 2670 16990
rect 2670 16970 2675 16990
rect 2645 16965 2675 16970
rect 2725 16990 2755 16995
rect 2725 16970 2730 16990
rect 2730 16970 2750 16990
rect 2750 16970 2755 16990
rect 2725 16965 2755 16970
rect 2805 16990 2835 16995
rect 2805 16970 2810 16990
rect 2810 16970 2830 16990
rect 2830 16970 2835 16990
rect 2805 16965 2835 16970
rect 2885 16990 2915 16995
rect 2885 16970 2890 16990
rect 2890 16970 2910 16990
rect 2910 16970 2915 16990
rect 2885 16965 2915 16970
rect 2965 16990 2995 16995
rect 2965 16970 2970 16990
rect 2970 16970 2990 16990
rect 2990 16970 2995 16990
rect 2965 16965 2995 16970
rect 3045 16990 3075 16995
rect 3045 16970 3050 16990
rect 3050 16970 3070 16990
rect 3070 16970 3075 16990
rect 3045 16965 3075 16970
rect 3125 16990 3155 16995
rect 3125 16970 3130 16990
rect 3130 16970 3150 16990
rect 3150 16970 3155 16990
rect 3125 16965 3155 16970
rect 3205 16990 3235 16995
rect 3205 16970 3210 16990
rect 3210 16970 3230 16990
rect 3230 16970 3235 16990
rect 3205 16965 3235 16970
rect 3285 16990 3315 16995
rect 3285 16970 3290 16990
rect 3290 16970 3310 16990
rect 3310 16970 3315 16990
rect 3285 16965 3315 16970
rect 3365 16990 3395 16995
rect 3365 16970 3370 16990
rect 3370 16970 3390 16990
rect 3390 16970 3395 16990
rect 3365 16965 3395 16970
rect 3445 16990 3475 16995
rect 3445 16970 3450 16990
rect 3450 16970 3470 16990
rect 3470 16970 3475 16990
rect 3445 16965 3475 16970
rect 3525 16990 3555 16995
rect 3525 16970 3530 16990
rect 3530 16970 3550 16990
rect 3550 16970 3555 16990
rect 3525 16965 3555 16970
rect 3605 16990 3635 16995
rect 3605 16970 3610 16990
rect 3610 16970 3630 16990
rect 3630 16970 3635 16990
rect 3605 16965 3635 16970
rect 3685 16990 3715 16995
rect 3685 16970 3690 16990
rect 3690 16970 3710 16990
rect 3710 16970 3715 16990
rect 3685 16965 3715 16970
rect 3765 16990 3795 16995
rect 3765 16970 3770 16990
rect 3770 16970 3790 16990
rect 3790 16970 3795 16990
rect 3765 16965 3795 16970
rect 3845 16990 3875 16995
rect 3845 16970 3850 16990
rect 3850 16970 3870 16990
rect 3870 16970 3875 16990
rect 3845 16965 3875 16970
rect 3925 16990 3955 16995
rect 3925 16970 3930 16990
rect 3930 16970 3950 16990
rect 3950 16970 3955 16990
rect 3925 16965 3955 16970
rect 4005 16990 4035 16995
rect 4005 16970 4010 16990
rect 4010 16970 4030 16990
rect 4030 16970 4035 16990
rect 4005 16965 4035 16970
rect 4085 16990 4115 16995
rect 4085 16970 4090 16990
rect 4090 16970 4110 16990
rect 4110 16970 4115 16990
rect 4085 16965 4115 16970
rect 4165 16990 4195 16995
rect 4165 16970 4170 16990
rect 4170 16970 4190 16990
rect 4190 16970 4195 16990
rect 4165 16965 4195 16970
rect 6245 16990 6275 16995
rect 6245 16970 6250 16990
rect 6250 16970 6270 16990
rect 6270 16970 6275 16990
rect 6245 16965 6275 16970
rect 6325 16990 6355 16995
rect 6325 16970 6330 16990
rect 6330 16970 6350 16990
rect 6350 16970 6355 16990
rect 6325 16965 6355 16970
rect 6405 16990 6435 16995
rect 6405 16970 6410 16990
rect 6410 16970 6430 16990
rect 6430 16970 6435 16990
rect 6405 16965 6435 16970
rect 6485 16990 6515 16995
rect 6485 16970 6490 16990
rect 6490 16970 6510 16990
rect 6510 16970 6515 16990
rect 6485 16965 6515 16970
rect 6565 16990 6595 16995
rect 6565 16970 6570 16990
rect 6570 16970 6590 16990
rect 6590 16970 6595 16990
rect 6565 16965 6595 16970
rect 6645 16990 6675 16995
rect 6645 16970 6650 16990
rect 6650 16970 6670 16990
rect 6670 16970 6675 16990
rect 6645 16965 6675 16970
rect 6725 16990 6755 16995
rect 6725 16970 6730 16990
rect 6730 16970 6750 16990
rect 6750 16970 6755 16990
rect 6725 16965 6755 16970
rect 6805 16990 6835 16995
rect 6805 16970 6810 16990
rect 6810 16970 6830 16990
rect 6830 16970 6835 16990
rect 6805 16965 6835 16970
rect 6885 16990 6915 16995
rect 6885 16970 6890 16990
rect 6890 16970 6910 16990
rect 6910 16970 6915 16990
rect 6885 16965 6915 16970
rect 6965 16990 6995 16995
rect 6965 16970 6970 16990
rect 6970 16970 6990 16990
rect 6990 16970 6995 16990
rect 6965 16965 6995 16970
rect 7045 16990 7075 16995
rect 7045 16970 7050 16990
rect 7050 16970 7070 16990
rect 7070 16970 7075 16990
rect 7045 16965 7075 16970
rect 7125 16990 7155 16995
rect 7125 16970 7130 16990
rect 7130 16970 7150 16990
rect 7150 16970 7155 16990
rect 7125 16965 7155 16970
rect 7205 16990 7235 16995
rect 7205 16970 7210 16990
rect 7210 16970 7230 16990
rect 7230 16970 7235 16990
rect 7205 16965 7235 16970
rect 7285 16990 7315 16995
rect 7285 16970 7290 16990
rect 7290 16970 7310 16990
rect 7310 16970 7315 16990
rect 7285 16965 7315 16970
rect 7365 16990 7395 16995
rect 7365 16970 7370 16990
rect 7370 16970 7390 16990
rect 7390 16970 7395 16990
rect 7365 16965 7395 16970
rect 7445 16990 7475 16995
rect 7445 16970 7450 16990
rect 7450 16970 7470 16990
rect 7470 16970 7475 16990
rect 7445 16965 7475 16970
rect 7525 16990 7555 16995
rect 7525 16970 7530 16990
rect 7530 16970 7550 16990
rect 7550 16970 7555 16990
rect 7525 16965 7555 16970
rect 7605 16990 7635 16995
rect 7605 16970 7610 16990
rect 7610 16970 7630 16990
rect 7630 16970 7635 16990
rect 7605 16965 7635 16970
rect 7685 16990 7715 16995
rect 7685 16970 7690 16990
rect 7690 16970 7710 16990
rect 7710 16970 7715 16990
rect 7685 16965 7715 16970
rect 7765 16990 7795 16995
rect 7765 16970 7770 16990
rect 7770 16970 7790 16990
rect 7790 16970 7795 16990
rect 7765 16965 7795 16970
rect 7845 16990 7875 16995
rect 7845 16970 7850 16990
rect 7850 16970 7870 16990
rect 7870 16970 7875 16990
rect 7845 16965 7875 16970
rect 7925 16990 7955 16995
rect 7925 16970 7930 16990
rect 7930 16970 7950 16990
rect 7950 16970 7955 16990
rect 7925 16965 7955 16970
rect 8005 16990 8035 16995
rect 8005 16970 8010 16990
rect 8010 16970 8030 16990
rect 8030 16970 8035 16990
rect 8005 16965 8035 16970
rect 8085 16990 8115 16995
rect 8085 16970 8090 16990
rect 8090 16970 8110 16990
rect 8110 16970 8115 16990
rect 8085 16965 8115 16970
rect 8165 16990 8195 16995
rect 8165 16970 8170 16990
rect 8170 16970 8190 16990
rect 8190 16970 8195 16990
rect 8165 16965 8195 16970
rect 8245 16990 8275 16995
rect 8245 16970 8250 16990
rect 8250 16970 8270 16990
rect 8270 16970 8275 16990
rect 8245 16965 8275 16970
rect 8325 16990 8355 16995
rect 8325 16970 8330 16990
rect 8330 16970 8350 16990
rect 8350 16970 8355 16990
rect 8325 16965 8355 16970
rect 8405 16990 8435 16995
rect 8405 16970 8410 16990
rect 8410 16970 8430 16990
rect 8430 16970 8435 16990
rect 8405 16965 8435 16970
rect 8485 16990 8515 16995
rect 8485 16970 8490 16990
rect 8490 16970 8510 16990
rect 8510 16970 8515 16990
rect 8485 16965 8515 16970
rect 8565 16990 8595 16995
rect 8565 16970 8570 16990
rect 8570 16970 8590 16990
rect 8590 16970 8595 16990
rect 8565 16965 8595 16970
rect 8645 16990 8675 16995
rect 8645 16970 8650 16990
rect 8650 16970 8670 16990
rect 8670 16970 8675 16990
rect 8645 16965 8675 16970
rect 8725 16990 8755 16995
rect 8725 16970 8730 16990
rect 8730 16970 8750 16990
rect 8750 16970 8755 16990
rect 8725 16965 8755 16970
rect 8805 16990 8835 16995
rect 8805 16970 8810 16990
rect 8810 16970 8830 16990
rect 8830 16970 8835 16990
rect 8805 16965 8835 16970
rect 8885 16990 8915 16995
rect 8885 16970 8890 16990
rect 8890 16970 8910 16990
rect 8910 16970 8915 16990
rect 8885 16965 8915 16970
rect 8965 16990 8995 16995
rect 8965 16970 8970 16990
rect 8970 16970 8990 16990
rect 8990 16970 8995 16990
rect 8965 16965 8995 16970
rect 9045 16990 9075 16995
rect 9045 16970 9050 16990
rect 9050 16970 9070 16990
rect 9070 16970 9075 16990
rect 9045 16965 9075 16970
rect 9125 16990 9155 16995
rect 9125 16970 9130 16990
rect 9130 16970 9150 16990
rect 9150 16970 9155 16990
rect 9125 16965 9155 16970
rect 9205 16990 9235 16995
rect 9205 16970 9210 16990
rect 9210 16970 9230 16990
rect 9230 16970 9235 16990
rect 9205 16965 9235 16970
rect 9285 16990 9315 16995
rect 9285 16970 9290 16990
rect 9290 16970 9310 16990
rect 9310 16970 9315 16990
rect 9285 16965 9315 16970
rect 9365 16990 9395 16995
rect 9365 16970 9370 16990
rect 9370 16970 9390 16990
rect 9390 16970 9395 16990
rect 9365 16965 9395 16970
rect 9445 16990 9475 16995
rect 9445 16970 9450 16990
rect 9450 16970 9470 16990
rect 9470 16970 9475 16990
rect 9445 16965 9475 16970
rect 11565 16990 11595 16995
rect 11565 16970 11570 16990
rect 11570 16970 11590 16990
rect 11590 16970 11595 16990
rect 11565 16965 11595 16970
rect 11645 16990 11675 16995
rect 11645 16970 11650 16990
rect 11650 16970 11670 16990
rect 11670 16970 11675 16990
rect 11645 16965 11675 16970
rect 11725 16990 11755 16995
rect 11725 16970 11730 16990
rect 11730 16970 11750 16990
rect 11750 16970 11755 16990
rect 11725 16965 11755 16970
rect 11805 16990 11835 16995
rect 11805 16970 11810 16990
rect 11810 16970 11830 16990
rect 11830 16970 11835 16990
rect 11805 16965 11835 16970
rect 11885 16990 11915 16995
rect 11885 16970 11890 16990
rect 11890 16970 11910 16990
rect 11910 16970 11915 16990
rect 11885 16965 11915 16970
rect 11965 16990 11995 16995
rect 11965 16970 11970 16990
rect 11970 16970 11990 16990
rect 11990 16970 11995 16990
rect 11965 16965 11995 16970
rect 12045 16990 12075 16995
rect 12045 16970 12050 16990
rect 12050 16970 12070 16990
rect 12070 16970 12075 16990
rect 12045 16965 12075 16970
rect 12125 16990 12155 16995
rect 12125 16970 12130 16990
rect 12130 16970 12150 16990
rect 12150 16970 12155 16990
rect 12125 16965 12155 16970
rect 12205 16990 12235 16995
rect 12205 16970 12210 16990
rect 12210 16970 12230 16990
rect 12230 16970 12235 16990
rect 12205 16965 12235 16970
rect 12285 16990 12315 16995
rect 12285 16970 12290 16990
rect 12290 16970 12310 16990
rect 12310 16970 12315 16990
rect 12285 16965 12315 16970
rect 12365 16990 12395 16995
rect 12365 16970 12370 16990
rect 12370 16970 12390 16990
rect 12390 16970 12395 16990
rect 12365 16965 12395 16970
rect 12445 16990 12475 16995
rect 12445 16970 12450 16990
rect 12450 16970 12470 16990
rect 12470 16970 12475 16990
rect 12445 16965 12475 16970
rect 12525 16990 12555 16995
rect 12525 16970 12530 16990
rect 12530 16970 12550 16990
rect 12550 16970 12555 16990
rect 12525 16965 12555 16970
rect 12605 16990 12635 16995
rect 12605 16970 12610 16990
rect 12610 16970 12630 16990
rect 12630 16970 12635 16990
rect 12605 16965 12635 16970
rect 12685 16990 12715 16995
rect 12685 16970 12690 16990
rect 12690 16970 12710 16990
rect 12710 16970 12715 16990
rect 12685 16965 12715 16970
rect 12765 16990 12795 16995
rect 12765 16970 12770 16990
rect 12770 16970 12790 16990
rect 12790 16970 12795 16990
rect 12765 16965 12795 16970
rect 12845 16990 12875 16995
rect 12845 16970 12850 16990
rect 12850 16970 12870 16990
rect 12870 16970 12875 16990
rect 12845 16965 12875 16970
rect 12925 16990 12955 16995
rect 12925 16970 12930 16990
rect 12930 16970 12950 16990
rect 12950 16970 12955 16990
rect 12925 16965 12955 16970
rect 13005 16990 13035 16995
rect 13005 16970 13010 16990
rect 13010 16970 13030 16990
rect 13030 16970 13035 16990
rect 13005 16965 13035 16970
rect 13085 16990 13115 16995
rect 13085 16970 13090 16990
rect 13090 16970 13110 16990
rect 13110 16970 13115 16990
rect 13085 16965 13115 16970
rect 13165 16990 13195 16995
rect 13165 16970 13170 16990
rect 13170 16970 13190 16990
rect 13190 16970 13195 16990
rect 13165 16965 13195 16970
rect 13245 16990 13275 16995
rect 13245 16970 13250 16990
rect 13250 16970 13270 16990
rect 13270 16970 13275 16990
rect 13245 16965 13275 16970
rect 13325 16990 13355 16995
rect 13325 16970 13330 16990
rect 13330 16970 13350 16990
rect 13350 16970 13355 16990
rect 13325 16965 13355 16970
rect 13405 16990 13435 16995
rect 13405 16970 13410 16990
rect 13410 16970 13430 16990
rect 13430 16970 13435 16990
rect 13405 16965 13435 16970
rect 13485 16990 13515 16995
rect 13485 16970 13490 16990
rect 13490 16970 13510 16990
rect 13510 16970 13515 16990
rect 13485 16965 13515 16970
rect 13565 16990 13595 16995
rect 13565 16970 13570 16990
rect 13570 16970 13590 16990
rect 13590 16970 13595 16990
rect 13565 16965 13595 16970
rect 13645 16990 13675 16995
rect 13645 16970 13650 16990
rect 13650 16970 13670 16990
rect 13670 16970 13675 16990
rect 13645 16965 13675 16970
rect 13725 16990 13755 16995
rect 13725 16970 13730 16990
rect 13730 16970 13750 16990
rect 13750 16970 13755 16990
rect 13725 16965 13755 16970
rect 13805 16990 13835 16995
rect 13805 16970 13810 16990
rect 13810 16970 13830 16990
rect 13830 16970 13835 16990
rect 13805 16965 13835 16970
rect 13885 16990 13915 16995
rect 13885 16970 13890 16990
rect 13890 16970 13910 16990
rect 13910 16970 13915 16990
rect 13885 16965 13915 16970
rect 13965 16990 13995 16995
rect 13965 16970 13970 16990
rect 13970 16970 13990 16990
rect 13990 16970 13995 16990
rect 13965 16965 13995 16970
rect 14045 16990 14075 16995
rect 14045 16970 14050 16990
rect 14050 16970 14070 16990
rect 14070 16970 14075 16990
rect 14045 16965 14075 16970
rect 14125 16990 14155 16995
rect 14125 16970 14130 16990
rect 14130 16970 14150 16990
rect 14150 16970 14155 16990
rect 14125 16965 14155 16970
rect 14205 16990 14235 16995
rect 14205 16970 14210 16990
rect 14210 16970 14230 16990
rect 14230 16970 14235 16990
rect 14205 16965 14235 16970
rect 14285 16990 14315 16995
rect 14285 16970 14290 16990
rect 14290 16970 14310 16990
rect 14310 16970 14315 16990
rect 14285 16965 14315 16970
rect 14365 16990 14395 16995
rect 14365 16970 14370 16990
rect 14370 16970 14390 16990
rect 14390 16970 14395 16990
rect 14365 16965 14395 16970
rect 14445 16990 14475 16995
rect 14445 16970 14450 16990
rect 14450 16970 14470 16990
rect 14470 16970 14475 16990
rect 14445 16965 14475 16970
rect 14525 16990 14555 16995
rect 14525 16970 14530 16990
rect 14530 16970 14550 16990
rect 14550 16970 14555 16990
rect 14525 16965 14555 16970
rect 14605 16990 14635 16995
rect 14605 16970 14610 16990
rect 14610 16970 14630 16990
rect 14630 16970 14635 16990
rect 14605 16965 14635 16970
rect 14685 16990 14715 16995
rect 14685 16970 14690 16990
rect 14690 16970 14710 16990
rect 14710 16970 14715 16990
rect 14685 16965 14715 16970
rect 16765 16990 16795 16995
rect 16765 16970 16770 16990
rect 16770 16970 16790 16990
rect 16790 16970 16795 16990
rect 16765 16965 16795 16970
rect 16845 16990 16875 16995
rect 16845 16970 16850 16990
rect 16850 16970 16870 16990
rect 16870 16970 16875 16990
rect 16845 16965 16875 16970
rect 16925 16990 16955 16995
rect 16925 16970 16930 16990
rect 16930 16970 16950 16990
rect 16950 16970 16955 16990
rect 16925 16965 16955 16970
rect 17005 16990 17035 16995
rect 17005 16970 17010 16990
rect 17010 16970 17030 16990
rect 17030 16970 17035 16990
rect 17005 16965 17035 16970
rect 17085 16990 17115 16995
rect 17085 16970 17090 16990
rect 17090 16970 17110 16990
rect 17110 16970 17115 16990
rect 17085 16965 17115 16970
rect 17165 16990 17195 16995
rect 17165 16970 17170 16990
rect 17170 16970 17190 16990
rect 17190 16970 17195 16990
rect 17165 16965 17195 16970
rect 17245 16990 17275 16995
rect 17245 16970 17250 16990
rect 17250 16970 17270 16990
rect 17270 16970 17275 16990
rect 17245 16965 17275 16970
rect 17325 16990 17355 16995
rect 17325 16970 17330 16990
rect 17330 16970 17350 16990
rect 17350 16970 17355 16990
rect 17325 16965 17355 16970
rect 17405 16990 17435 16995
rect 17405 16970 17410 16990
rect 17410 16970 17430 16990
rect 17430 16970 17435 16990
rect 17405 16965 17435 16970
rect 17485 16990 17515 16995
rect 17485 16970 17490 16990
rect 17490 16970 17510 16990
rect 17510 16970 17515 16990
rect 17485 16965 17515 16970
rect 17565 16990 17595 16995
rect 17565 16970 17570 16990
rect 17570 16970 17590 16990
rect 17590 16970 17595 16990
rect 17565 16965 17595 16970
rect 17645 16990 17675 16995
rect 17645 16970 17650 16990
rect 17650 16970 17670 16990
rect 17670 16970 17675 16990
rect 17645 16965 17675 16970
rect 17725 16990 17755 16995
rect 17725 16970 17730 16990
rect 17730 16970 17750 16990
rect 17750 16970 17755 16990
rect 17725 16965 17755 16970
rect 17805 16990 17835 16995
rect 17805 16970 17810 16990
rect 17810 16970 17830 16990
rect 17830 16970 17835 16990
rect 17805 16965 17835 16970
rect 17885 16990 17915 16995
rect 17885 16970 17890 16990
rect 17890 16970 17910 16990
rect 17910 16970 17915 16990
rect 17885 16965 17915 16970
rect 17965 16990 17995 16995
rect 17965 16970 17970 16990
rect 17970 16970 17990 16990
rect 17990 16970 17995 16990
rect 17965 16965 17995 16970
rect 18045 16990 18075 16995
rect 18045 16970 18050 16990
rect 18050 16970 18070 16990
rect 18070 16970 18075 16990
rect 18045 16965 18075 16970
rect 18125 16990 18155 16995
rect 18125 16970 18130 16990
rect 18130 16970 18150 16990
rect 18150 16970 18155 16990
rect 18125 16965 18155 16970
rect 18205 16990 18235 16995
rect 18205 16970 18210 16990
rect 18210 16970 18230 16990
rect 18230 16970 18235 16990
rect 18205 16965 18235 16970
rect 18285 16990 18315 16995
rect 18285 16970 18290 16990
rect 18290 16970 18310 16990
rect 18310 16970 18315 16990
rect 18285 16965 18315 16970
rect 18365 16990 18395 16995
rect 18365 16970 18370 16990
rect 18370 16970 18390 16990
rect 18390 16970 18395 16990
rect 18365 16965 18395 16970
rect 18445 16990 18475 16995
rect 18445 16970 18450 16990
rect 18450 16970 18470 16990
rect 18470 16970 18475 16990
rect 18445 16965 18475 16970
rect 18525 16990 18555 16995
rect 18525 16970 18530 16990
rect 18530 16970 18550 16990
rect 18550 16970 18555 16990
rect 18525 16965 18555 16970
rect 18605 16990 18635 16995
rect 18605 16970 18610 16990
rect 18610 16970 18630 16990
rect 18630 16970 18635 16990
rect 18605 16965 18635 16970
rect 18685 16990 18715 16995
rect 18685 16970 18690 16990
rect 18690 16970 18710 16990
rect 18710 16970 18715 16990
rect 18685 16965 18715 16970
rect 18765 16990 18795 16995
rect 18765 16970 18770 16990
rect 18770 16970 18790 16990
rect 18790 16970 18795 16990
rect 18765 16965 18795 16970
rect 18845 16990 18875 16995
rect 18845 16970 18850 16990
rect 18850 16970 18870 16990
rect 18870 16970 18875 16990
rect 18845 16965 18875 16970
rect 18925 16990 18955 16995
rect 18925 16970 18930 16990
rect 18930 16970 18950 16990
rect 18950 16970 18955 16990
rect 18925 16965 18955 16970
rect 19005 16990 19035 16995
rect 19005 16970 19010 16990
rect 19010 16970 19030 16990
rect 19030 16970 19035 16990
rect 19005 16965 19035 16970
rect 19085 16990 19115 16995
rect 19085 16970 19090 16990
rect 19090 16970 19110 16990
rect 19110 16970 19115 16990
rect 19085 16965 19115 16970
rect 19165 16990 19195 16995
rect 19165 16970 19170 16990
rect 19170 16970 19190 16990
rect 19190 16970 19195 16990
rect 19165 16965 19195 16970
rect 19245 16990 19275 16995
rect 19245 16970 19250 16990
rect 19250 16970 19270 16990
rect 19270 16970 19275 16990
rect 19245 16965 19275 16970
rect 19325 16990 19355 16995
rect 19325 16970 19330 16990
rect 19330 16970 19350 16990
rect 19350 16970 19355 16990
rect 19325 16965 19355 16970
rect 19405 16990 19435 16995
rect 19405 16970 19410 16990
rect 19410 16970 19430 16990
rect 19430 16970 19435 16990
rect 19405 16965 19435 16970
rect 19485 16990 19515 16995
rect 19485 16970 19490 16990
rect 19490 16970 19510 16990
rect 19510 16970 19515 16990
rect 19485 16965 19515 16970
rect 19565 16990 19595 16995
rect 19565 16970 19570 16990
rect 19570 16970 19590 16990
rect 19590 16970 19595 16990
rect 19565 16965 19595 16970
rect 19645 16990 19675 16995
rect 19645 16970 19650 16990
rect 19650 16970 19670 16990
rect 19670 16970 19675 16990
rect 19645 16965 19675 16970
rect 19725 16990 19755 16995
rect 19725 16970 19730 16990
rect 19730 16970 19750 16990
rect 19750 16970 19755 16990
rect 19725 16965 19755 16970
rect 19805 16990 19835 16995
rect 19805 16970 19810 16990
rect 19810 16970 19830 16990
rect 19830 16970 19835 16990
rect 19805 16965 19835 16970
rect 19885 16990 19915 16995
rect 19885 16970 19890 16990
rect 19890 16970 19910 16990
rect 19910 16970 19915 16990
rect 19885 16965 19915 16970
rect 19965 16990 19995 16995
rect 19965 16970 19970 16990
rect 19970 16970 19990 16990
rect 19990 16970 19995 16990
rect 19965 16965 19995 16970
rect 20045 16990 20075 16995
rect 20045 16970 20050 16990
rect 20050 16970 20070 16990
rect 20070 16970 20075 16990
rect 20045 16965 20075 16970
rect 20125 16990 20155 16995
rect 20125 16970 20130 16990
rect 20130 16970 20150 16990
rect 20150 16970 20155 16990
rect 20125 16965 20155 16970
rect 20205 16990 20235 16995
rect 20205 16970 20210 16990
rect 20210 16970 20230 16990
rect 20230 16970 20235 16990
rect 20205 16965 20235 16970
rect 20285 16990 20315 16995
rect 20285 16970 20290 16990
rect 20290 16970 20310 16990
rect 20310 16970 20315 16990
rect 20285 16965 20315 16970
rect 20365 16990 20395 16995
rect 20365 16970 20370 16990
rect 20370 16970 20390 16990
rect 20390 16970 20395 16990
rect 20365 16965 20395 16970
rect 20445 16990 20475 16995
rect 20445 16970 20450 16990
rect 20450 16970 20470 16990
rect 20470 16970 20475 16990
rect 20445 16965 20475 16970
rect 20525 16990 20555 16995
rect 20525 16970 20530 16990
rect 20530 16970 20550 16990
rect 20550 16970 20555 16990
rect 20525 16965 20555 16970
rect 20605 16990 20635 16995
rect 20605 16970 20610 16990
rect 20610 16970 20630 16990
rect 20630 16970 20635 16990
rect 20605 16965 20635 16970
rect 20685 16990 20715 16995
rect 20685 16970 20690 16990
rect 20690 16970 20710 16990
rect 20710 16970 20715 16990
rect 20685 16965 20715 16970
rect 20765 16990 20795 16995
rect 20765 16970 20770 16990
rect 20770 16970 20790 16990
rect 20790 16970 20795 16990
rect 20765 16965 20795 16970
rect 20845 16990 20875 16995
rect 20845 16970 20850 16990
rect 20850 16970 20870 16990
rect 20870 16970 20875 16990
rect 20845 16965 20875 16970
rect 20925 16990 20955 16995
rect 20925 16970 20930 16990
rect 20930 16970 20950 16990
rect 20950 16970 20955 16990
rect 20925 16965 20955 16970
rect 5 16910 35 16915
rect 5 16890 10 16910
rect 10 16890 30 16910
rect 30 16890 35 16910
rect 5 16885 35 16890
rect 85 16910 115 16915
rect 85 16890 90 16910
rect 90 16890 110 16910
rect 110 16890 115 16910
rect 85 16885 115 16890
rect 165 16910 195 16915
rect 165 16890 170 16910
rect 170 16890 190 16910
rect 190 16890 195 16910
rect 165 16885 195 16890
rect 245 16910 275 16915
rect 245 16890 250 16910
rect 250 16890 270 16910
rect 270 16890 275 16910
rect 245 16885 275 16890
rect 325 16910 355 16915
rect 325 16890 330 16910
rect 330 16890 350 16910
rect 350 16890 355 16910
rect 325 16885 355 16890
rect 405 16910 435 16915
rect 405 16890 410 16910
rect 410 16890 430 16910
rect 430 16890 435 16910
rect 405 16885 435 16890
rect 485 16910 515 16915
rect 485 16890 490 16910
rect 490 16890 510 16910
rect 510 16890 515 16910
rect 485 16885 515 16890
rect 565 16910 595 16915
rect 565 16890 570 16910
rect 570 16890 590 16910
rect 590 16890 595 16910
rect 565 16885 595 16890
rect 645 16910 675 16915
rect 645 16890 650 16910
rect 650 16890 670 16910
rect 670 16890 675 16910
rect 645 16885 675 16890
rect 725 16910 755 16915
rect 725 16890 730 16910
rect 730 16890 750 16910
rect 750 16890 755 16910
rect 725 16885 755 16890
rect 805 16910 835 16915
rect 805 16890 810 16910
rect 810 16890 830 16910
rect 830 16890 835 16910
rect 805 16885 835 16890
rect 885 16910 915 16915
rect 885 16890 890 16910
rect 890 16890 910 16910
rect 910 16890 915 16910
rect 885 16885 915 16890
rect 965 16910 995 16915
rect 965 16890 970 16910
rect 970 16890 990 16910
rect 990 16890 995 16910
rect 965 16885 995 16890
rect 1045 16910 1075 16915
rect 1045 16890 1050 16910
rect 1050 16890 1070 16910
rect 1070 16890 1075 16910
rect 1045 16885 1075 16890
rect 1125 16910 1155 16915
rect 1125 16890 1130 16910
rect 1130 16890 1150 16910
rect 1150 16890 1155 16910
rect 1125 16885 1155 16890
rect 1205 16910 1235 16915
rect 1205 16890 1210 16910
rect 1210 16890 1230 16910
rect 1230 16890 1235 16910
rect 1205 16885 1235 16890
rect 1285 16910 1315 16915
rect 1285 16890 1290 16910
rect 1290 16890 1310 16910
rect 1310 16890 1315 16910
rect 1285 16885 1315 16890
rect 1365 16910 1395 16915
rect 1365 16890 1370 16910
rect 1370 16890 1390 16910
rect 1390 16890 1395 16910
rect 1365 16885 1395 16890
rect 1445 16910 1475 16915
rect 1445 16890 1450 16910
rect 1450 16890 1470 16910
rect 1470 16890 1475 16910
rect 1445 16885 1475 16890
rect 1525 16910 1555 16915
rect 1525 16890 1530 16910
rect 1530 16890 1550 16910
rect 1550 16890 1555 16910
rect 1525 16885 1555 16890
rect 1605 16910 1635 16915
rect 1605 16890 1610 16910
rect 1610 16890 1630 16910
rect 1630 16890 1635 16910
rect 1605 16885 1635 16890
rect 1685 16910 1715 16915
rect 1685 16890 1690 16910
rect 1690 16890 1710 16910
rect 1710 16890 1715 16910
rect 1685 16885 1715 16890
rect 1765 16910 1795 16915
rect 1765 16890 1770 16910
rect 1770 16890 1790 16910
rect 1790 16890 1795 16910
rect 1765 16885 1795 16890
rect 1845 16910 1875 16915
rect 1845 16890 1850 16910
rect 1850 16890 1870 16910
rect 1870 16890 1875 16910
rect 1845 16885 1875 16890
rect 1925 16910 1955 16915
rect 1925 16890 1930 16910
rect 1930 16890 1950 16910
rect 1950 16890 1955 16910
rect 1925 16885 1955 16890
rect 2005 16910 2035 16915
rect 2005 16890 2010 16910
rect 2010 16890 2030 16910
rect 2030 16890 2035 16910
rect 2005 16885 2035 16890
rect 2085 16910 2115 16915
rect 2085 16890 2090 16910
rect 2090 16890 2110 16910
rect 2110 16890 2115 16910
rect 2085 16885 2115 16890
rect 2165 16910 2195 16915
rect 2165 16890 2170 16910
rect 2170 16890 2190 16910
rect 2190 16890 2195 16910
rect 2165 16885 2195 16890
rect 2245 16910 2275 16915
rect 2245 16890 2250 16910
rect 2250 16890 2270 16910
rect 2270 16890 2275 16910
rect 2245 16885 2275 16890
rect 2325 16910 2355 16915
rect 2325 16890 2330 16910
rect 2330 16890 2350 16910
rect 2350 16890 2355 16910
rect 2325 16885 2355 16890
rect 2405 16910 2435 16915
rect 2405 16890 2410 16910
rect 2410 16890 2430 16910
rect 2430 16890 2435 16910
rect 2405 16885 2435 16890
rect 2485 16910 2515 16915
rect 2485 16890 2490 16910
rect 2490 16890 2510 16910
rect 2510 16890 2515 16910
rect 2485 16885 2515 16890
rect 2565 16910 2595 16915
rect 2565 16890 2570 16910
rect 2570 16890 2590 16910
rect 2590 16890 2595 16910
rect 2565 16885 2595 16890
rect 2645 16910 2675 16915
rect 2645 16890 2650 16910
rect 2650 16890 2670 16910
rect 2670 16890 2675 16910
rect 2645 16885 2675 16890
rect 2725 16910 2755 16915
rect 2725 16890 2730 16910
rect 2730 16890 2750 16910
rect 2750 16890 2755 16910
rect 2725 16885 2755 16890
rect 2805 16910 2835 16915
rect 2805 16890 2810 16910
rect 2810 16890 2830 16910
rect 2830 16890 2835 16910
rect 2805 16885 2835 16890
rect 2885 16910 2915 16915
rect 2885 16890 2890 16910
rect 2890 16890 2910 16910
rect 2910 16890 2915 16910
rect 2885 16885 2915 16890
rect 2965 16910 2995 16915
rect 2965 16890 2970 16910
rect 2970 16890 2990 16910
rect 2990 16890 2995 16910
rect 2965 16885 2995 16890
rect 3045 16910 3075 16915
rect 3045 16890 3050 16910
rect 3050 16890 3070 16910
rect 3070 16890 3075 16910
rect 3045 16885 3075 16890
rect 3125 16910 3155 16915
rect 3125 16890 3130 16910
rect 3130 16890 3150 16910
rect 3150 16890 3155 16910
rect 3125 16885 3155 16890
rect 3205 16910 3235 16915
rect 3205 16890 3210 16910
rect 3210 16890 3230 16910
rect 3230 16890 3235 16910
rect 3205 16885 3235 16890
rect 3285 16910 3315 16915
rect 3285 16890 3290 16910
rect 3290 16890 3310 16910
rect 3310 16890 3315 16910
rect 3285 16885 3315 16890
rect 3365 16910 3395 16915
rect 3365 16890 3370 16910
rect 3370 16890 3390 16910
rect 3390 16890 3395 16910
rect 3365 16885 3395 16890
rect 3445 16910 3475 16915
rect 3445 16890 3450 16910
rect 3450 16890 3470 16910
rect 3470 16890 3475 16910
rect 3445 16885 3475 16890
rect 3525 16910 3555 16915
rect 3525 16890 3530 16910
rect 3530 16890 3550 16910
rect 3550 16890 3555 16910
rect 3525 16885 3555 16890
rect 3605 16910 3635 16915
rect 3605 16890 3610 16910
rect 3610 16890 3630 16910
rect 3630 16890 3635 16910
rect 3605 16885 3635 16890
rect 3685 16910 3715 16915
rect 3685 16890 3690 16910
rect 3690 16890 3710 16910
rect 3710 16890 3715 16910
rect 3685 16885 3715 16890
rect 3765 16910 3795 16915
rect 3765 16890 3770 16910
rect 3770 16890 3790 16910
rect 3790 16890 3795 16910
rect 3765 16885 3795 16890
rect 3845 16910 3875 16915
rect 3845 16890 3850 16910
rect 3850 16890 3870 16910
rect 3870 16890 3875 16910
rect 3845 16885 3875 16890
rect 3925 16910 3955 16915
rect 3925 16890 3930 16910
rect 3930 16890 3950 16910
rect 3950 16890 3955 16910
rect 3925 16885 3955 16890
rect 4005 16910 4035 16915
rect 4005 16890 4010 16910
rect 4010 16890 4030 16910
rect 4030 16890 4035 16910
rect 4005 16885 4035 16890
rect 4085 16910 4115 16915
rect 4085 16890 4090 16910
rect 4090 16890 4110 16910
rect 4110 16890 4115 16910
rect 4085 16885 4115 16890
rect 4165 16910 4195 16915
rect 4165 16890 4170 16910
rect 4170 16890 4190 16910
rect 4190 16890 4195 16910
rect 4165 16885 4195 16890
rect 6245 16910 6275 16915
rect 6245 16890 6250 16910
rect 6250 16890 6270 16910
rect 6270 16890 6275 16910
rect 6245 16885 6275 16890
rect 6325 16910 6355 16915
rect 6325 16890 6330 16910
rect 6330 16890 6350 16910
rect 6350 16890 6355 16910
rect 6325 16885 6355 16890
rect 6405 16910 6435 16915
rect 6405 16890 6410 16910
rect 6410 16890 6430 16910
rect 6430 16890 6435 16910
rect 6405 16885 6435 16890
rect 6485 16910 6515 16915
rect 6485 16890 6490 16910
rect 6490 16890 6510 16910
rect 6510 16890 6515 16910
rect 6485 16885 6515 16890
rect 6565 16910 6595 16915
rect 6565 16890 6570 16910
rect 6570 16890 6590 16910
rect 6590 16890 6595 16910
rect 6565 16885 6595 16890
rect 6645 16910 6675 16915
rect 6645 16890 6650 16910
rect 6650 16890 6670 16910
rect 6670 16890 6675 16910
rect 6645 16885 6675 16890
rect 6725 16910 6755 16915
rect 6725 16890 6730 16910
rect 6730 16890 6750 16910
rect 6750 16890 6755 16910
rect 6725 16885 6755 16890
rect 6805 16910 6835 16915
rect 6805 16890 6810 16910
rect 6810 16890 6830 16910
rect 6830 16890 6835 16910
rect 6805 16885 6835 16890
rect 6885 16910 6915 16915
rect 6885 16890 6890 16910
rect 6890 16890 6910 16910
rect 6910 16890 6915 16910
rect 6885 16885 6915 16890
rect 6965 16910 6995 16915
rect 6965 16890 6970 16910
rect 6970 16890 6990 16910
rect 6990 16890 6995 16910
rect 6965 16885 6995 16890
rect 7045 16910 7075 16915
rect 7045 16890 7050 16910
rect 7050 16890 7070 16910
rect 7070 16890 7075 16910
rect 7045 16885 7075 16890
rect 7125 16910 7155 16915
rect 7125 16890 7130 16910
rect 7130 16890 7150 16910
rect 7150 16890 7155 16910
rect 7125 16885 7155 16890
rect 7205 16910 7235 16915
rect 7205 16890 7210 16910
rect 7210 16890 7230 16910
rect 7230 16890 7235 16910
rect 7205 16885 7235 16890
rect 7285 16910 7315 16915
rect 7285 16890 7290 16910
rect 7290 16890 7310 16910
rect 7310 16890 7315 16910
rect 7285 16885 7315 16890
rect 7365 16910 7395 16915
rect 7365 16890 7370 16910
rect 7370 16890 7390 16910
rect 7390 16890 7395 16910
rect 7365 16885 7395 16890
rect 7445 16910 7475 16915
rect 7445 16890 7450 16910
rect 7450 16890 7470 16910
rect 7470 16890 7475 16910
rect 7445 16885 7475 16890
rect 7525 16910 7555 16915
rect 7525 16890 7530 16910
rect 7530 16890 7550 16910
rect 7550 16890 7555 16910
rect 7525 16885 7555 16890
rect 7605 16910 7635 16915
rect 7605 16890 7610 16910
rect 7610 16890 7630 16910
rect 7630 16890 7635 16910
rect 7605 16885 7635 16890
rect 7685 16910 7715 16915
rect 7685 16890 7690 16910
rect 7690 16890 7710 16910
rect 7710 16890 7715 16910
rect 7685 16885 7715 16890
rect 7765 16910 7795 16915
rect 7765 16890 7770 16910
rect 7770 16890 7790 16910
rect 7790 16890 7795 16910
rect 7765 16885 7795 16890
rect 7845 16910 7875 16915
rect 7845 16890 7850 16910
rect 7850 16890 7870 16910
rect 7870 16890 7875 16910
rect 7845 16885 7875 16890
rect 7925 16910 7955 16915
rect 7925 16890 7930 16910
rect 7930 16890 7950 16910
rect 7950 16890 7955 16910
rect 7925 16885 7955 16890
rect 8005 16910 8035 16915
rect 8005 16890 8010 16910
rect 8010 16890 8030 16910
rect 8030 16890 8035 16910
rect 8005 16885 8035 16890
rect 8085 16910 8115 16915
rect 8085 16890 8090 16910
rect 8090 16890 8110 16910
rect 8110 16890 8115 16910
rect 8085 16885 8115 16890
rect 8165 16910 8195 16915
rect 8165 16890 8170 16910
rect 8170 16890 8190 16910
rect 8190 16890 8195 16910
rect 8165 16885 8195 16890
rect 8245 16910 8275 16915
rect 8245 16890 8250 16910
rect 8250 16890 8270 16910
rect 8270 16890 8275 16910
rect 8245 16885 8275 16890
rect 8325 16910 8355 16915
rect 8325 16890 8330 16910
rect 8330 16890 8350 16910
rect 8350 16890 8355 16910
rect 8325 16885 8355 16890
rect 8405 16910 8435 16915
rect 8405 16890 8410 16910
rect 8410 16890 8430 16910
rect 8430 16890 8435 16910
rect 8405 16885 8435 16890
rect 8485 16910 8515 16915
rect 8485 16890 8490 16910
rect 8490 16890 8510 16910
rect 8510 16890 8515 16910
rect 8485 16885 8515 16890
rect 8565 16910 8595 16915
rect 8565 16890 8570 16910
rect 8570 16890 8590 16910
rect 8590 16890 8595 16910
rect 8565 16885 8595 16890
rect 8645 16910 8675 16915
rect 8645 16890 8650 16910
rect 8650 16890 8670 16910
rect 8670 16890 8675 16910
rect 8645 16885 8675 16890
rect 8725 16910 8755 16915
rect 8725 16890 8730 16910
rect 8730 16890 8750 16910
rect 8750 16890 8755 16910
rect 8725 16885 8755 16890
rect 8805 16910 8835 16915
rect 8805 16890 8810 16910
rect 8810 16890 8830 16910
rect 8830 16890 8835 16910
rect 8805 16885 8835 16890
rect 8885 16910 8915 16915
rect 8885 16890 8890 16910
rect 8890 16890 8910 16910
rect 8910 16890 8915 16910
rect 8885 16885 8915 16890
rect 8965 16910 8995 16915
rect 8965 16890 8970 16910
rect 8970 16890 8990 16910
rect 8990 16890 8995 16910
rect 8965 16885 8995 16890
rect 9045 16910 9075 16915
rect 9045 16890 9050 16910
rect 9050 16890 9070 16910
rect 9070 16890 9075 16910
rect 9045 16885 9075 16890
rect 9125 16910 9155 16915
rect 9125 16890 9130 16910
rect 9130 16890 9150 16910
rect 9150 16890 9155 16910
rect 9125 16885 9155 16890
rect 9205 16910 9235 16915
rect 9205 16890 9210 16910
rect 9210 16890 9230 16910
rect 9230 16890 9235 16910
rect 9205 16885 9235 16890
rect 9285 16910 9315 16915
rect 9285 16890 9290 16910
rect 9290 16890 9310 16910
rect 9310 16890 9315 16910
rect 9285 16885 9315 16890
rect 9365 16910 9395 16915
rect 9365 16890 9370 16910
rect 9370 16890 9390 16910
rect 9390 16890 9395 16910
rect 9365 16885 9395 16890
rect 9445 16910 9475 16915
rect 9445 16890 9450 16910
rect 9450 16890 9470 16910
rect 9470 16890 9475 16910
rect 9445 16885 9475 16890
rect 11565 16910 11595 16915
rect 11565 16890 11570 16910
rect 11570 16890 11590 16910
rect 11590 16890 11595 16910
rect 11565 16885 11595 16890
rect 11645 16910 11675 16915
rect 11645 16890 11650 16910
rect 11650 16890 11670 16910
rect 11670 16890 11675 16910
rect 11645 16885 11675 16890
rect 11725 16910 11755 16915
rect 11725 16890 11730 16910
rect 11730 16890 11750 16910
rect 11750 16890 11755 16910
rect 11725 16885 11755 16890
rect 11805 16910 11835 16915
rect 11805 16890 11810 16910
rect 11810 16890 11830 16910
rect 11830 16890 11835 16910
rect 11805 16885 11835 16890
rect 11885 16910 11915 16915
rect 11885 16890 11890 16910
rect 11890 16890 11910 16910
rect 11910 16890 11915 16910
rect 11885 16885 11915 16890
rect 11965 16910 11995 16915
rect 11965 16890 11970 16910
rect 11970 16890 11990 16910
rect 11990 16890 11995 16910
rect 11965 16885 11995 16890
rect 12045 16910 12075 16915
rect 12045 16890 12050 16910
rect 12050 16890 12070 16910
rect 12070 16890 12075 16910
rect 12045 16885 12075 16890
rect 12125 16910 12155 16915
rect 12125 16890 12130 16910
rect 12130 16890 12150 16910
rect 12150 16890 12155 16910
rect 12125 16885 12155 16890
rect 12205 16910 12235 16915
rect 12205 16890 12210 16910
rect 12210 16890 12230 16910
rect 12230 16890 12235 16910
rect 12205 16885 12235 16890
rect 12285 16910 12315 16915
rect 12285 16890 12290 16910
rect 12290 16890 12310 16910
rect 12310 16890 12315 16910
rect 12285 16885 12315 16890
rect 12365 16910 12395 16915
rect 12365 16890 12370 16910
rect 12370 16890 12390 16910
rect 12390 16890 12395 16910
rect 12365 16885 12395 16890
rect 12445 16910 12475 16915
rect 12445 16890 12450 16910
rect 12450 16890 12470 16910
rect 12470 16890 12475 16910
rect 12445 16885 12475 16890
rect 12525 16910 12555 16915
rect 12525 16890 12530 16910
rect 12530 16890 12550 16910
rect 12550 16890 12555 16910
rect 12525 16885 12555 16890
rect 12605 16910 12635 16915
rect 12605 16890 12610 16910
rect 12610 16890 12630 16910
rect 12630 16890 12635 16910
rect 12605 16885 12635 16890
rect 12685 16910 12715 16915
rect 12685 16890 12690 16910
rect 12690 16890 12710 16910
rect 12710 16890 12715 16910
rect 12685 16885 12715 16890
rect 12765 16910 12795 16915
rect 12765 16890 12770 16910
rect 12770 16890 12790 16910
rect 12790 16890 12795 16910
rect 12765 16885 12795 16890
rect 12845 16910 12875 16915
rect 12845 16890 12850 16910
rect 12850 16890 12870 16910
rect 12870 16890 12875 16910
rect 12845 16885 12875 16890
rect 12925 16910 12955 16915
rect 12925 16890 12930 16910
rect 12930 16890 12950 16910
rect 12950 16890 12955 16910
rect 12925 16885 12955 16890
rect 13005 16910 13035 16915
rect 13005 16890 13010 16910
rect 13010 16890 13030 16910
rect 13030 16890 13035 16910
rect 13005 16885 13035 16890
rect 13085 16910 13115 16915
rect 13085 16890 13090 16910
rect 13090 16890 13110 16910
rect 13110 16890 13115 16910
rect 13085 16885 13115 16890
rect 13165 16910 13195 16915
rect 13165 16890 13170 16910
rect 13170 16890 13190 16910
rect 13190 16890 13195 16910
rect 13165 16885 13195 16890
rect 13245 16910 13275 16915
rect 13245 16890 13250 16910
rect 13250 16890 13270 16910
rect 13270 16890 13275 16910
rect 13245 16885 13275 16890
rect 13325 16910 13355 16915
rect 13325 16890 13330 16910
rect 13330 16890 13350 16910
rect 13350 16890 13355 16910
rect 13325 16885 13355 16890
rect 13405 16910 13435 16915
rect 13405 16890 13410 16910
rect 13410 16890 13430 16910
rect 13430 16890 13435 16910
rect 13405 16885 13435 16890
rect 13485 16910 13515 16915
rect 13485 16890 13490 16910
rect 13490 16890 13510 16910
rect 13510 16890 13515 16910
rect 13485 16885 13515 16890
rect 13565 16910 13595 16915
rect 13565 16890 13570 16910
rect 13570 16890 13590 16910
rect 13590 16890 13595 16910
rect 13565 16885 13595 16890
rect 13645 16910 13675 16915
rect 13645 16890 13650 16910
rect 13650 16890 13670 16910
rect 13670 16890 13675 16910
rect 13645 16885 13675 16890
rect 13725 16910 13755 16915
rect 13725 16890 13730 16910
rect 13730 16890 13750 16910
rect 13750 16890 13755 16910
rect 13725 16885 13755 16890
rect 13805 16910 13835 16915
rect 13805 16890 13810 16910
rect 13810 16890 13830 16910
rect 13830 16890 13835 16910
rect 13805 16885 13835 16890
rect 13885 16910 13915 16915
rect 13885 16890 13890 16910
rect 13890 16890 13910 16910
rect 13910 16890 13915 16910
rect 13885 16885 13915 16890
rect 13965 16910 13995 16915
rect 13965 16890 13970 16910
rect 13970 16890 13990 16910
rect 13990 16890 13995 16910
rect 13965 16885 13995 16890
rect 14045 16910 14075 16915
rect 14045 16890 14050 16910
rect 14050 16890 14070 16910
rect 14070 16890 14075 16910
rect 14045 16885 14075 16890
rect 14125 16910 14155 16915
rect 14125 16890 14130 16910
rect 14130 16890 14150 16910
rect 14150 16890 14155 16910
rect 14125 16885 14155 16890
rect 14205 16910 14235 16915
rect 14205 16890 14210 16910
rect 14210 16890 14230 16910
rect 14230 16890 14235 16910
rect 14205 16885 14235 16890
rect 14285 16910 14315 16915
rect 14285 16890 14290 16910
rect 14290 16890 14310 16910
rect 14310 16890 14315 16910
rect 14285 16885 14315 16890
rect 14365 16910 14395 16915
rect 14365 16890 14370 16910
rect 14370 16890 14390 16910
rect 14390 16890 14395 16910
rect 14365 16885 14395 16890
rect 14445 16910 14475 16915
rect 14445 16890 14450 16910
rect 14450 16890 14470 16910
rect 14470 16890 14475 16910
rect 14445 16885 14475 16890
rect 14525 16910 14555 16915
rect 14525 16890 14530 16910
rect 14530 16890 14550 16910
rect 14550 16890 14555 16910
rect 14525 16885 14555 16890
rect 14605 16910 14635 16915
rect 14605 16890 14610 16910
rect 14610 16890 14630 16910
rect 14630 16890 14635 16910
rect 14605 16885 14635 16890
rect 14685 16910 14715 16915
rect 14685 16890 14690 16910
rect 14690 16890 14710 16910
rect 14710 16890 14715 16910
rect 14685 16885 14715 16890
rect 16765 16910 16795 16915
rect 16765 16890 16770 16910
rect 16770 16890 16790 16910
rect 16790 16890 16795 16910
rect 16765 16885 16795 16890
rect 16845 16910 16875 16915
rect 16845 16890 16850 16910
rect 16850 16890 16870 16910
rect 16870 16890 16875 16910
rect 16845 16885 16875 16890
rect 16925 16910 16955 16915
rect 16925 16890 16930 16910
rect 16930 16890 16950 16910
rect 16950 16890 16955 16910
rect 16925 16885 16955 16890
rect 17005 16910 17035 16915
rect 17005 16890 17010 16910
rect 17010 16890 17030 16910
rect 17030 16890 17035 16910
rect 17005 16885 17035 16890
rect 17085 16910 17115 16915
rect 17085 16890 17090 16910
rect 17090 16890 17110 16910
rect 17110 16890 17115 16910
rect 17085 16885 17115 16890
rect 17165 16910 17195 16915
rect 17165 16890 17170 16910
rect 17170 16890 17190 16910
rect 17190 16890 17195 16910
rect 17165 16885 17195 16890
rect 17245 16910 17275 16915
rect 17245 16890 17250 16910
rect 17250 16890 17270 16910
rect 17270 16890 17275 16910
rect 17245 16885 17275 16890
rect 17325 16910 17355 16915
rect 17325 16890 17330 16910
rect 17330 16890 17350 16910
rect 17350 16890 17355 16910
rect 17325 16885 17355 16890
rect 17405 16910 17435 16915
rect 17405 16890 17410 16910
rect 17410 16890 17430 16910
rect 17430 16890 17435 16910
rect 17405 16885 17435 16890
rect 17485 16910 17515 16915
rect 17485 16890 17490 16910
rect 17490 16890 17510 16910
rect 17510 16890 17515 16910
rect 17485 16885 17515 16890
rect 17565 16910 17595 16915
rect 17565 16890 17570 16910
rect 17570 16890 17590 16910
rect 17590 16890 17595 16910
rect 17565 16885 17595 16890
rect 17645 16910 17675 16915
rect 17645 16890 17650 16910
rect 17650 16890 17670 16910
rect 17670 16890 17675 16910
rect 17645 16885 17675 16890
rect 17725 16910 17755 16915
rect 17725 16890 17730 16910
rect 17730 16890 17750 16910
rect 17750 16890 17755 16910
rect 17725 16885 17755 16890
rect 17805 16910 17835 16915
rect 17805 16890 17810 16910
rect 17810 16890 17830 16910
rect 17830 16890 17835 16910
rect 17805 16885 17835 16890
rect 17885 16910 17915 16915
rect 17885 16890 17890 16910
rect 17890 16890 17910 16910
rect 17910 16890 17915 16910
rect 17885 16885 17915 16890
rect 17965 16910 17995 16915
rect 17965 16890 17970 16910
rect 17970 16890 17990 16910
rect 17990 16890 17995 16910
rect 17965 16885 17995 16890
rect 18045 16910 18075 16915
rect 18045 16890 18050 16910
rect 18050 16890 18070 16910
rect 18070 16890 18075 16910
rect 18045 16885 18075 16890
rect 18125 16910 18155 16915
rect 18125 16890 18130 16910
rect 18130 16890 18150 16910
rect 18150 16890 18155 16910
rect 18125 16885 18155 16890
rect 18205 16910 18235 16915
rect 18205 16890 18210 16910
rect 18210 16890 18230 16910
rect 18230 16890 18235 16910
rect 18205 16885 18235 16890
rect 18285 16910 18315 16915
rect 18285 16890 18290 16910
rect 18290 16890 18310 16910
rect 18310 16890 18315 16910
rect 18285 16885 18315 16890
rect 18365 16910 18395 16915
rect 18365 16890 18370 16910
rect 18370 16890 18390 16910
rect 18390 16890 18395 16910
rect 18365 16885 18395 16890
rect 18445 16910 18475 16915
rect 18445 16890 18450 16910
rect 18450 16890 18470 16910
rect 18470 16890 18475 16910
rect 18445 16885 18475 16890
rect 18525 16910 18555 16915
rect 18525 16890 18530 16910
rect 18530 16890 18550 16910
rect 18550 16890 18555 16910
rect 18525 16885 18555 16890
rect 18605 16910 18635 16915
rect 18605 16890 18610 16910
rect 18610 16890 18630 16910
rect 18630 16890 18635 16910
rect 18605 16885 18635 16890
rect 18685 16910 18715 16915
rect 18685 16890 18690 16910
rect 18690 16890 18710 16910
rect 18710 16890 18715 16910
rect 18685 16885 18715 16890
rect 18765 16910 18795 16915
rect 18765 16890 18770 16910
rect 18770 16890 18790 16910
rect 18790 16890 18795 16910
rect 18765 16885 18795 16890
rect 18845 16910 18875 16915
rect 18845 16890 18850 16910
rect 18850 16890 18870 16910
rect 18870 16890 18875 16910
rect 18845 16885 18875 16890
rect 18925 16910 18955 16915
rect 18925 16890 18930 16910
rect 18930 16890 18950 16910
rect 18950 16890 18955 16910
rect 18925 16885 18955 16890
rect 19005 16910 19035 16915
rect 19005 16890 19010 16910
rect 19010 16890 19030 16910
rect 19030 16890 19035 16910
rect 19005 16885 19035 16890
rect 19085 16910 19115 16915
rect 19085 16890 19090 16910
rect 19090 16890 19110 16910
rect 19110 16890 19115 16910
rect 19085 16885 19115 16890
rect 19165 16910 19195 16915
rect 19165 16890 19170 16910
rect 19170 16890 19190 16910
rect 19190 16890 19195 16910
rect 19165 16885 19195 16890
rect 19245 16910 19275 16915
rect 19245 16890 19250 16910
rect 19250 16890 19270 16910
rect 19270 16890 19275 16910
rect 19245 16885 19275 16890
rect 19325 16910 19355 16915
rect 19325 16890 19330 16910
rect 19330 16890 19350 16910
rect 19350 16890 19355 16910
rect 19325 16885 19355 16890
rect 19405 16910 19435 16915
rect 19405 16890 19410 16910
rect 19410 16890 19430 16910
rect 19430 16890 19435 16910
rect 19405 16885 19435 16890
rect 19485 16910 19515 16915
rect 19485 16890 19490 16910
rect 19490 16890 19510 16910
rect 19510 16890 19515 16910
rect 19485 16885 19515 16890
rect 19565 16910 19595 16915
rect 19565 16890 19570 16910
rect 19570 16890 19590 16910
rect 19590 16890 19595 16910
rect 19565 16885 19595 16890
rect 19645 16910 19675 16915
rect 19645 16890 19650 16910
rect 19650 16890 19670 16910
rect 19670 16890 19675 16910
rect 19645 16885 19675 16890
rect 19725 16910 19755 16915
rect 19725 16890 19730 16910
rect 19730 16890 19750 16910
rect 19750 16890 19755 16910
rect 19725 16885 19755 16890
rect 19805 16910 19835 16915
rect 19805 16890 19810 16910
rect 19810 16890 19830 16910
rect 19830 16890 19835 16910
rect 19805 16885 19835 16890
rect 19885 16910 19915 16915
rect 19885 16890 19890 16910
rect 19890 16890 19910 16910
rect 19910 16890 19915 16910
rect 19885 16885 19915 16890
rect 19965 16910 19995 16915
rect 19965 16890 19970 16910
rect 19970 16890 19990 16910
rect 19990 16890 19995 16910
rect 19965 16885 19995 16890
rect 20045 16910 20075 16915
rect 20045 16890 20050 16910
rect 20050 16890 20070 16910
rect 20070 16890 20075 16910
rect 20045 16885 20075 16890
rect 20125 16910 20155 16915
rect 20125 16890 20130 16910
rect 20130 16890 20150 16910
rect 20150 16890 20155 16910
rect 20125 16885 20155 16890
rect 20205 16910 20235 16915
rect 20205 16890 20210 16910
rect 20210 16890 20230 16910
rect 20230 16890 20235 16910
rect 20205 16885 20235 16890
rect 20285 16910 20315 16915
rect 20285 16890 20290 16910
rect 20290 16890 20310 16910
rect 20310 16890 20315 16910
rect 20285 16885 20315 16890
rect 20365 16910 20395 16915
rect 20365 16890 20370 16910
rect 20370 16890 20390 16910
rect 20390 16890 20395 16910
rect 20365 16885 20395 16890
rect 20445 16910 20475 16915
rect 20445 16890 20450 16910
rect 20450 16890 20470 16910
rect 20470 16890 20475 16910
rect 20445 16885 20475 16890
rect 20525 16910 20555 16915
rect 20525 16890 20530 16910
rect 20530 16890 20550 16910
rect 20550 16890 20555 16910
rect 20525 16885 20555 16890
rect 20605 16910 20635 16915
rect 20605 16890 20610 16910
rect 20610 16890 20630 16910
rect 20630 16890 20635 16910
rect 20605 16885 20635 16890
rect 20685 16910 20715 16915
rect 20685 16890 20690 16910
rect 20690 16890 20710 16910
rect 20710 16890 20715 16910
rect 20685 16885 20715 16890
rect 20765 16910 20795 16915
rect 20765 16890 20770 16910
rect 20770 16890 20790 16910
rect 20790 16890 20795 16910
rect 20765 16885 20795 16890
rect 20845 16910 20875 16915
rect 20845 16890 20850 16910
rect 20850 16890 20870 16910
rect 20870 16890 20875 16910
rect 20845 16885 20875 16890
rect 20925 16910 20955 16915
rect 20925 16890 20930 16910
rect 20930 16890 20950 16910
rect 20950 16890 20955 16910
rect 20925 16885 20955 16890
rect 5 16750 35 16755
rect 5 16730 10 16750
rect 10 16730 30 16750
rect 30 16730 35 16750
rect 5 16725 35 16730
rect 85 16750 115 16755
rect 85 16730 90 16750
rect 90 16730 110 16750
rect 110 16730 115 16750
rect 85 16725 115 16730
rect 165 16750 195 16755
rect 165 16730 170 16750
rect 170 16730 190 16750
rect 190 16730 195 16750
rect 165 16725 195 16730
rect 245 16750 275 16755
rect 245 16730 250 16750
rect 250 16730 270 16750
rect 270 16730 275 16750
rect 245 16725 275 16730
rect 325 16750 355 16755
rect 325 16730 330 16750
rect 330 16730 350 16750
rect 350 16730 355 16750
rect 325 16725 355 16730
rect 405 16750 435 16755
rect 405 16730 410 16750
rect 410 16730 430 16750
rect 430 16730 435 16750
rect 405 16725 435 16730
rect 485 16750 515 16755
rect 485 16730 490 16750
rect 490 16730 510 16750
rect 510 16730 515 16750
rect 485 16725 515 16730
rect 565 16750 595 16755
rect 565 16730 570 16750
rect 570 16730 590 16750
rect 590 16730 595 16750
rect 565 16725 595 16730
rect 645 16750 675 16755
rect 645 16730 650 16750
rect 650 16730 670 16750
rect 670 16730 675 16750
rect 645 16725 675 16730
rect 725 16750 755 16755
rect 725 16730 730 16750
rect 730 16730 750 16750
rect 750 16730 755 16750
rect 725 16725 755 16730
rect 805 16750 835 16755
rect 805 16730 810 16750
rect 810 16730 830 16750
rect 830 16730 835 16750
rect 805 16725 835 16730
rect 885 16750 915 16755
rect 885 16730 890 16750
rect 890 16730 910 16750
rect 910 16730 915 16750
rect 885 16725 915 16730
rect 965 16750 995 16755
rect 965 16730 970 16750
rect 970 16730 990 16750
rect 990 16730 995 16750
rect 965 16725 995 16730
rect 1045 16750 1075 16755
rect 1045 16730 1050 16750
rect 1050 16730 1070 16750
rect 1070 16730 1075 16750
rect 1045 16725 1075 16730
rect 1125 16750 1155 16755
rect 1125 16730 1130 16750
rect 1130 16730 1150 16750
rect 1150 16730 1155 16750
rect 1125 16725 1155 16730
rect 1205 16750 1235 16755
rect 1205 16730 1210 16750
rect 1210 16730 1230 16750
rect 1230 16730 1235 16750
rect 1205 16725 1235 16730
rect 1285 16750 1315 16755
rect 1285 16730 1290 16750
rect 1290 16730 1310 16750
rect 1310 16730 1315 16750
rect 1285 16725 1315 16730
rect 1365 16750 1395 16755
rect 1365 16730 1370 16750
rect 1370 16730 1390 16750
rect 1390 16730 1395 16750
rect 1365 16725 1395 16730
rect 1445 16750 1475 16755
rect 1445 16730 1450 16750
rect 1450 16730 1470 16750
rect 1470 16730 1475 16750
rect 1445 16725 1475 16730
rect 1525 16750 1555 16755
rect 1525 16730 1530 16750
rect 1530 16730 1550 16750
rect 1550 16730 1555 16750
rect 1525 16725 1555 16730
rect 1605 16750 1635 16755
rect 1605 16730 1610 16750
rect 1610 16730 1630 16750
rect 1630 16730 1635 16750
rect 1605 16725 1635 16730
rect 1685 16750 1715 16755
rect 1685 16730 1690 16750
rect 1690 16730 1710 16750
rect 1710 16730 1715 16750
rect 1685 16725 1715 16730
rect 1765 16750 1795 16755
rect 1765 16730 1770 16750
rect 1770 16730 1790 16750
rect 1790 16730 1795 16750
rect 1765 16725 1795 16730
rect 1845 16750 1875 16755
rect 1845 16730 1850 16750
rect 1850 16730 1870 16750
rect 1870 16730 1875 16750
rect 1845 16725 1875 16730
rect 1925 16750 1955 16755
rect 1925 16730 1930 16750
rect 1930 16730 1950 16750
rect 1950 16730 1955 16750
rect 1925 16725 1955 16730
rect 2005 16750 2035 16755
rect 2005 16730 2010 16750
rect 2010 16730 2030 16750
rect 2030 16730 2035 16750
rect 2005 16725 2035 16730
rect 2085 16750 2115 16755
rect 2085 16730 2090 16750
rect 2090 16730 2110 16750
rect 2110 16730 2115 16750
rect 2085 16725 2115 16730
rect 2165 16750 2195 16755
rect 2165 16730 2170 16750
rect 2170 16730 2190 16750
rect 2190 16730 2195 16750
rect 2165 16725 2195 16730
rect 2245 16750 2275 16755
rect 2245 16730 2250 16750
rect 2250 16730 2270 16750
rect 2270 16730 2275 16750
rect 2245 16725 2275 16730
rect 2325 16750 2355 16755
rect 2325 16730 2330 16750
rect 2330 16730 2350 16750
rect 2350 16730 2355 16750
rect 2325 16725 2355 16730
rect 2405 16750 2435 16755
rect 2405 16730 2410 16750
rect 2410 16730 2430 16750
rect 2430 16730 2435 16750
rect 2405 16725 2435 16730
rect 2485 16750 2515 16755
rect 2485 16730 2490 16750
rect 2490 16730 2510 16750
rect 2510 16730 2515 16750
rect 2485 16725 2515 16730
rect 2565 16750 2595 16755
rect 2565 16730 2570 16750
rect 2570 16730 2590 16750
rect 2590 16730 2595 16750
rect 2565 16725 2595 16730
rect 2645 16750 2675 16755
rect 2645 16730 2650 16750
rect 2650 16730 2670 16750
rect 2670 16730 2675 16750
rect 2645 16725 2675 16730
rect 2725 16750 2755 16755
rect 2725 16730 2730 16750
rect 2730 16730 2750 16750
rect 2750 16730 2755 16750
rect 2725 16725 2755 16730
rect 2805 16750 2835 16755
rect 2805 16730 2810 16750
rect 2810 16730 2830 16750
rect 2830 16730 2835 16750
rect 2805 16725 2835 16730
rect 2885 16750 2915 16755
rect 2885 16730 2890 16750
rect 2890 16730 2910 16750
rect 2910 16730 2915 16750
rect 2885 16725 2915 16730
rect 2965 16750 2995 16755
rect 2965 16730 2970 16750
rect 2970 16730 2990 16750
rect 2990 16730 2995 16750
rect 2965 16725 2995 16730
rect 3045 16750 3075 16755
rect 3045 16730 3050 16750
rect 3050 16730 3070 16750
rect 3070 16730 3075 16750
rect 3045 16725 3075 16730
rect 3125 16750 3155 16755
rect 3125 16730 3130 16750
rect 3130 16730 3150 16750
rect 3150 16730 3155 16750
rect 3125 16725 3155 16730
rect 3205 16750 3235 16755
rect 3205 16730 3210 16750
rect 3210 16730 3230 16750
rect 3230 16730 3235 16750
rect 3205 16725 3235 16730
rect 3285 16750 3315 16755
rect 3285 16730 3290 16750
rect 3290 16730 3310 16750
rect 3310 16730 3315 16750
rect 3285 16725 3315 16730
rect 3365 16750 3395 16755
rect 3365 16730 3370 16750
rect 3370 16730 3390 16750
rect 3390 16730 3395 16750
rect 3365 16725 3395 16730
rect 3445 16750 3475 16755
rect 3445 16730 3450 16750
rect 3450 16730 3470 16750
rect 3470 16730 3475 16750
rect 3445 16725 3475 16730
rect 3525 16750 3555 16755
rect 3525 16730 3530 16750
rect 3530 16730 3550 16750
rect 3550 16730 3555 16750
rect 3525 16725 3555 16730
rect 3605 16750 3635 16755
rect 3605 16730 3610 16750
rect 3610 16730 3630 16750
rect 3630 16730 3635 16750
rect 3605 16725 3635 16730
rect 3685 16750 3715 16755
rect 3685 16730 3690 16750
rect 3690 16730 3710 16750
rect 3710 16730 3715 16750
rect 3685 16725 3715 16730
rect 3765 16750 3795 16755
rect 3765 16730 3770 16750
rect 3770 16730 3790 16750
rect 3790 16730 3795 16750
rect 3765 16725 3795 16730
rect 3845 16750 3875 16755
rect 3845 16730 3850 16750
rect 3850 16730 3870 16750
rect 3870 16730 3875 16750
rect 3845 16725 3875 16730
rect 3925 16750 3955 16755
rect 3925 16730 3930 16750
rect 3930 16730 3950 16750
rect 3950 16730 3955 16750
rect 3925 16725 3955 16730
rect 4005 16750 4035 16755
rect 4005 16730 4010 16750
rect 4010 16730 4030 16750
rect 4030 16730 4035 16750
rect 4005 16725 4035 16730
rect 4085 16750 4115 16755
rect 4085 16730 4090 16750
rect 4090 16730 4110 16750
rect 4110 16730 4115 16750
rect 4085 16725 4115 16730
rect 4165 16750 4195 16755
rect 4165 16730 4170 16750
rect 4170 16730 4190 16750
rect 4190 16730 4195 16750
rect 4165 16725 4195 16730
rect 6245 16750 6275 16755
rect 6245 16730 6250 16750
rect 6250 16730 6270 16750
rect 6270 16730 6275 16750
rect 6245 16725 6275 16730
rect 6325 16750 6355 16755
rect 6325 16730 6330 16750
rect 6330 16730 6350 16750
rect 6350 16730 6355 16750
rect 6325 16725 6355 16730
rect 6405 16750 6435 16755
rect 6405 16730 6410 16750
rect 6410 16730 6430 16750
rect 6430 16730 6435 16750
rect 6405 16725 6435 16730
rect 6485 16750 6515 16755
rect 6485 16730 6490 16750
rect 6490 16730 6510 16750
rect 6510 16730 6515 16750
rect 6485 16725 6515 16730
rect 6565 16750 6595 16755
rect 6565 16730 6570 16750
rect 6570 16730 6590 16750
rect 6590 16730 6595 16750
rect 6565 16725 6595 16730
rect 6645 16750 6675 16755
rect 6645 16730 6650 16750
rect 6650 16730 6670 16750
rect 6670 16730 6675 16750
rect 6645 16725 6675 16730
rect 6725 16750 6755 16755
rect 6725 16730 6730 16750
rect 6730 16730 6750 16750
rect 6750 16730 6755 16750
rect 6725 16725 6755 16730
rect 6805 16750 6835 16755
rect 6805 16730 6810 16750
rect 6810 16730 6830 16750
rect 6830 16730 6835 16750
rect 6805 16725 6835 16730
rect 6885 16750 6915 16755
rect 6885 16730 6890 16750
rect 6890 16730 6910 16750
rect 6910 16730 6915 16750
rect 6885 16725 6915 16730
rect 6965 16750 6995 16755
rect 6965 16730 6970 16750
rect 6970 16730 6990 16750
rect 6990 16730 6995 16750
rect 6965 16725 6995 16730
rect 7045 16750 7075 16755
rect 7045 16730 7050 16750
rect 7050 16730 7070 16750
rect 7070 16730 7075 16750
rect 7045 16725 7075 16730
rect 7125 16750 7155 16755
rect 7125 16730 7130 16750
rect 7130 16730 7150 16750
rect 7150 16730 7155 16750
rect 7125 16725 7155 16730
rect 7205 16750 7235 16755
rect 7205 16730 7210 16750
rect 7210 16730 7230 16750
rect 7230 16730 7235 16750
rect 7205 16725 7235 16730
rect 7285 16750 7315 16755
rect 7285 16730 7290 16750
rect 7290 16730 7310 16750
rect 7310 16730 7315 16750
rect 7285 16725 7315 16730
rect 7365 16750 7395 16755
rect 7365 16730 7370 16750
rect 7370 16730 7390 16750
rect 7390 16730 7395 16750
rect 7365 16725 7395 16730
rect 7445 16750 7475 16755
rect 7445 16730 7450 16750
rect 7450 16730 7470 16750
rect 7470 16730 7475 16750
rect 7445 16725 7475 16730
rect 7525 16750 7555 16755
rect 7525 16730 7530 16750
rect 7530 16730 7550 16750
rect 7550 16730 7555 16750
rect 7525 16725 7555 16730
rect 7605 16750 7635 16755
rect 7605 16730 7610 16750
rect 7610 16730 7630 16750
rect 7630 16730 7635 16750
rect 7605 16725 7635 16730
rect 7685 16750 7715 16755
rect 7685 16730 7690 16750
rect 7690 16730 7710 16750
rect 7710 16730 7715 16750
rect 7685 16725 7715 16730
rect 7765 16750 7795 16755
rect 7765 16730 7770 16750
rect 7770 16730 7790 16750
rect 7790 16730 7795 16750
rect 7765 16725 7795 16730
rect 7845 16750 7875 16755
rect 7845 16730 7850 16750
rect 7850 16730 7870 16750
rect 7870 16730 7875 16750
rect 7845 16725 7875 16730
rect 7925 16750 7955 16755
rect 7925 16730 7930 16750
rect 7930 16730 7950 16750
rect 7950 16730 7955 16750
rect 7925 16725 7955 16730
rect 8005 16750 8035 16755
rect 8005 16730 8010 16750
rect 8010 16730 8030 16750
rect 8030 16730 8035 16750
rect 8005 16725 8035 16730
rect 8085 16750 8115 16755
rect 8085 16730 8090 16750
rect 8090 16730 8110 16750
rect 8110 16730 8115 16750
rect 8085 16725 8115 16730
rect 8165 16750 8195 16755
rect 8165 16730 8170 16750
rect 8170 16730 8190 16750
rect 8190 16730 8195 16750
rect 8165 16725 8195 16730
rect 8245 16750 8275 16755
rect 8245 16730 8250 16750
rect 8250 16730 8270 16750
rect 8270 16730 8275 16750
rect 8245 16725 8275 16730
rect 8325 16750 8355 16755
rect 8325 16730 8330 16750
rect 8330 16730 8350 16750
rect 8350 16730 8355 16750
rect 8325 16725 8355 16730
rect 8405 16750 8435 16755
rect 8405 16730 8410 16750
rect 8410 16730 8430 16750
rect 8430 16730 8435 16750
rect 8405 16725 8435 16730
rect 8485 16750 8515 16755
rect 8485 16730 8490 16750
rect 8490 16730 8510 16750
rect 8510 16730 8515 16750
rect 8485 16725 8515 16730
rect 8565 16750 8595 16755
rect 8565 16730 8570 16750
rect 8570 16730 8590 16750
rect 8590 16730 8595 16750
rect 8565 16725 8595 16730
rect 8645 16750 8675 16755
rect 8645 16730 8650 16750
rect 8650 16730 8670 16750
rect 8670 16730 8675 16750
rect 8645 16725 8675 16730
rect 8725 16750 8755 16755
rect 8725 16730 8730 16750
rect 8730 16730 8750 16750
rect 8750 16730 8755 16750
rect 8725 16725 8755 16730
rect 8805 16750 8835 16755
rect 8805 16730 8810 16750
rect 8810 16730 8830 16750
rect 8830 16730 8835 16750
rect 8805 16725 8835 16730
rect 8885 16750 8915 16755
rect 8885 16730 8890 16750
rect 8890 16730 8910 16750
rect 8910 16730 8915 16750
rect 8885 16725 8915 16730
rect 8965 16750 8995 16755
rect 8965 16730 8970 16750
rect 8970 16730 8990 16750
rect 8990 16730 8995 16750
rect 8965 16725 8995 16730
rect 9045 16750 9075 16755
rect 9045 16730 9050 16750
rect 9050 16730 9070 16750
rect 9070 16730 9075 16750
rect 9045 16725 9075 16730
rect 9125 16750 9155 16755
rect 9125 16730 9130 16750
rect 9130 16730 9150 16750
rect 9150 16730 9155 16750
rect 9125 16725 9155 16730
rect 9205 16750 9235 16755
rect 9205 16730 9210 16750
rect 9210 16730 9230 16750
rect 9230 16730 9235 16750
rect 9205 16725 9235 16730
rect 9285 16750 9315 16755
rect 9285 16730 9290 16750
rect 9290 16730 9310 16750
rect 9310 16730 9315 16750
rect 9285 16725 9315 16730
rect 9365 16750 9395 16755
rect 9365 16730 9370 16750
rect 9370 16730 9390 16750
rect 9390 16730 9395 16750
rect 9365 16725 9395 16730
rect 9445 16750 9475 16755
rect 9445 16730 9450 16750
rect 9450 16730 9470 16750
rect 9470 16730 9475 16750
rect 9445 16725 9475 16730
rect 11565 16750 11595 16755
rect 11565 16730 11570 16750
rect 11570 16730 11590 16750
rect 11590 16730 11595 16750
rect 11565 16725 11595 16730
rect 11645 16750 11675 16755
rect 11645 16730 11650 16750
rect 11650 16730 11670 16750
rect 11670 16730 11675 16750
rect 11645 16725 11675 16730
rect 11725 16750 11755 16755
rect 11725 16730 11730 16750
rect 11730 16730 11750 16750
rect 11750 16730 11755 16750
rect 11725 16725 11755 16730
rect 11805 16750 11835 16755
rect 11805 16730 11810 16750
rect 11810 16730 11830 16750
rect 11830 16730 11835 16750
rect 11805 16725 11835 16730
rect 11885 16750 11915 16755
rect 11885 16730 11890 16750
rect 11890 16730 11910 16750
rect 11910 16730 11915 16750
rect 11885 16725 11915 16730
rect 11965 16750 11995 16755
rect 11965 16730 11970 16750
rect 11970 16730 11990 16750
rect 11990 16730 11995 16750
rect 11965 16725 11995 16730
rect 12045 16750 12075 16755
rect 12045 16730 12050 16750
rect 12050 16730 12070 16750
rect 12070 16730 12075 16750
rect 12045 16725 12075 16730
rect 12125 16750 12155 16755
rect 12125 16730 12130 16750
rect 12130 16730 12150 16750
rect 12150 16730 12155 16750
rect 12125 16725 12155 16730
rect 12205 16750 12235 16755
rect 12205 16730 12210 16750
rect 12210 16730 12230 16750
rect 12230 16730 12235 16750
rect 12205 16725 12235 16730
rect 12285 16750 12315 16755
rect 12285 16730 12290 16750
rect 12290 16730 12310 16750
rect 12310 16730 12315 16750
rect 12285 16725 12315 16730
rect 12365 16750 12395 16755
rect 12365 16730 12370 16750
rect 12370 16730 12390 16750
rect 12390 16730 12395 16750
rect 12365 16725 12395 16730
rect 12445 16750 12475 16755
rect 12445 16730 12450 16750
rect 12450 16730 12470 16750
rect 12470 16730 12475 16750
rect 12445 16725 12475 16730
rect 12525 16750 12555 16755
rect 12525 16730 12530 16750
rect 12530 16730 12550 16750
rect 12550 16730 12555 16750
rect 12525 16725 12555 16730
rect 12605 16750 12635 16755
rect 12605 16730 12610 16750
rect 12610 16730 12630 16750
rect 12630 16730 12635 16750
rect 12605 16725 12635 16730
rect 12685 16750 12715 16755
rect 12685 16730 12690 16750
rect 12690 16730 12710 16750
rect 12710 16730 12715 16750
rect 12685 16725 12715 16730
rect 12765 16750 12795 16755
rect 12765 16730 12770 16750
rect 12770 16730 12790 16750
rect 12790 16730 12795 16750
rect 12765 16725 12795 16730
rect 12845 16750 12875 16755
rect 12845 16730 12850 16750
rect 12850 16730 12870 16750
rect 12870 16730 12875 16750
rect 12845 16725 12875 16730
rect 12925 16750 12955 16755
rect 12925 16730 12930 16750
rect 12930 16730 12950 16750
rect 12950 16730 12955 16750
rect 12925 16725 12955 16730
rect 13005 16750 13035 16755
rect 13005 16730 13010 16750
rect 13010 16730 13030 16750
rect 13030 16730 13035 16750
rect 13005 16725 13035 16730
rect 13085 16750 13115 16755
rect 13085 16730 13090 16750
rect 13090 16730 13110 16750
rect 13110 16730 13115 16750
rect 13085 16725 13115 16730
rect 13165 16750 13195 16755
rect 13165 16730 13170 16750
rect 13170 16730 13190 16750
rect 13190 16730 13195 16750
rect 13165 16725 13195 16730
rect 13245 16750 13275 16755
rect 13245 16730 13250 16750
rect 13250 16730 13270 16750
rect 13270 16730 13275 16750
rect 13245 16725 13275 16730
rect 13325 16750 13355 16755
rect 13325 16730 13330 16750
rect 13330 16730 13350 16750
rect 13350 16730 13355 16750
rect 13325 16725 13355 16730
rect 13405 16750 13435 16755
rect 13405 16730 13410 16750
rect 13410 16730 13430 16750
rect 13430 16730 13435 16750
rect 13405 16725 13435 16730
rect 13485 16750 13515 16755
rect 13485 16730 13490 16750
rect 13490 16730 13510 16750
rect 13510 16730 13515 16750
rect 13485 16725 13515 16730
rect 13565 16750 13595 16755
rect 13565 16730 13570 16750
rect 13570 16730 13590 16750
rect 13590 16730 13595 16750
rect 13565 16725 13595 16730
rect 13645 16750 13675 16755
rect 13645 16730 13650 16750
rect 13650 16730 13670 16750
rect 13670 16730 13675 16750
rect 13645 16725 13675 16730
rect 13725 16750 13755 16755
rect 13725 16730 13730 16750
rect 13730 16730 13750 16750
rect 13750 16730 13755 16750
rect 13725 16725 13755 16730
rect 13805 16750 13835 16755
rect 13805 16730 13810 16750
rect 13810 16730 13830 16750
rect 13830 16730 13835 16750
rect 13805 16725 13835 16730
rect 13885 16750 13915 16755
rect 13885 16730 13890 16750
rect 13890 16730 13910 16750
rect 13910 16730 13915 16750
rect 13885 16725 13915 16730
rect 13965 16750 13995 16755
rect 13965 16730 13970 16750
rect 13970 16730 13990 16750
rect 13990 16730 13995 16750
rect 13965 16725 13995 16730
rect 14045 16750 14075 16755
rect 14045 16730 14050 16750
rect 14050 16730 14070 16750
rect 14070 16730 14075 16750
rect 14045 16725 14075 16730
rect 14125 16750 14155 16755
rect 14125 16730 14130 16750
rect 14130 16730 14150 16750
rect 14150 16730 14155 16750
rect 14125 16725 14155 16730
rect 14205 16750 14235 16755
rect 14205 16730 14210 16750
rect 14210 16730 14230 16750
rect 14230 16730 14235 16750
rect 14205 16725 14235 16730
rect 14285 16750 14315 16755
rect 14285 16730 14290 16750
rect 14290 16730 14310 16750
rect 14310 16730 14315 16750
rect 14285 16725 14315 16730
rect 14365 16750 14395 16755
rect 14365 16730 14370 16750
rect 14370 16730 14390 16750
rect 14390 16730 14395 16750
rect 14365 16725 14395 16730
rect 14445 16750 14475 16755
rect 14445 16730 14450 16750
rect 14450 16730 14470 16750
rect 14470 16730 14475 16750
rect 14445 16725 14475 16730
rect 14525 16750 14555 16755
rect 14525 16730 14530 16750
rect 14530 16730 14550 16750
rect 14550 16730 14555 16750
rect 14525 16725 14555 16730
rect 14605 16750 14635 16755
rect 14605 16730 14610 16750
rect 14610 16730 14630 16750
rect 14630 16730 14635 16750
rect 14605 16725 14635 16730
rect 14685 16750 14715 16755
rect 14685 16730 14690 16750
rect 14690 16730 14710 16750
rect 14710 16730 14715 16750
rect 14685 16725 14715 16730
rect 16765 16750 16795 16755
rect 16765 16730 16770 16750
rect 16770 16730 16790 16750
rect 16790 16730 16795 16750
rect 16765 16725 16795 16730
rect 16845 16750 16875 16755
rect 16845 16730 16850 16750
rect 16850 16730 16870 16750
rect 16870 16730 16875 16750
rect 16845 16725 16875 16730
rect 16925 16750 16955 16755
rect 16925 16730 16930 16750
rect 16930 16730 16950 16750
rect 16950 16730 16955 16750
rect 16925 16725 16955 16730
rect 17005 16750 17035 16755
rect 17005 16730 17010 16750
rect 17010 16730 17030 16750
rect 17030 16730 17035 16750
rect 17005 16725 17035 16730
rect 17085 16750 17115 16755
rect 17085 16730 17090 16750
rect 17090 16730 17110 16750
rect 17110 16730 17115 16750
rect 17085 16725 17115 16730
rect 17165 16750 17195 16755
rect 17165 16730 17170 16750
rect 17170 16730 17190 16750
rect 17190 16730 17195 16750
rect 17165 16725 17195 16730
rect 17245 16750 17275 16755
rect 17245 16730 17250 16750
rect 17250 16730 17270 16750
rect 17270 16730 17275 16750
rect 17245 16725 17275 16730
rect 17325 16750 17355 16755
rect 17325 16730 17330 16750
rect 17330 16730 17350 16750
rect 17350 16730 17355 16750
rect 17325 16725 17355 16730
rect 17405 16750 17435 16755
rect 17405 16730 17410 16750
rect 17410 16730 17430 16750
rect 17430 16730 17435 16750
rect 17405 16725 17435 16730
rect 17485 16750 17515 16755
rect 17485 16730 17490 16750
rect 17490 16730 17510 16750
rect 17510 16730 17515 16750
rect 17485 16725 17515 16730
rect 17565 16750 17595 16755
rect 17565 16730 17570 16750
rect 17570 16730 17590 16750
rect 17590 16730 17595 16750
rect 17565 16725 17595 16730
rect 17645 16750 17675 16755
rect 17645 16730 17650 16750
rect 17650 16730 17670 16750
rect 17670 16730 17675 16750
rect 17645 16725 17675 16730
rect 17725 16750 17755 16755
rect 17725 16730 17730 16750
rect 17730 16730 17750 16750
rect 17750 16730 17755 16750
rect 17725 16725 17755 16730
rect 17805 16750 17835 16755
rect 17805 16730 17810 16750
rect 17810 16730 17830 16750
rect 17830 16730 17835 16750
rect 17805 16725 17835 16730
rect 17885 16750 17915 16755
rect 17885 16730 17890 16750
rect 17890 16730 17910 16750
rect 17910 16730 17915 16750
rect 17885 16725 17915 16730
rect 17965 16750 17995 16755
rect 17965 16730 17970 16750
rect 17970 16730 17990 16750
rect 17990 16730 17995 16750
rect 17965 16725 17995 16730
rect 18045 16750 18075 16755
rect 18045 16730 18050 16750
rect 18050 16730 18070 16750
rect 18070 16730 18075 16750
rect 18045 16725 18075 16730
rect 18125 16750 18155 16755
rect 18125 16730 18130 16750
rect 18130 16730 18150 16750
rect 18150 16730 18155 16750
rect 18125 16725 18155 16730
rect 18205 16750 18235 16755
rect 18205 16730 18210 16750
rect 18210 16730 18230 16750
rect 18230 16730 18235 16750
rect 18205 16725 18235 16730
rect 18285 16750 18315 16755
rect 18285 16730 18290 16750
rect 18290 16730 18310 16750
rect 18310 16730 18315 16750
rect 18285 16725 18315 16730
rect 18365 16750 18395 16755
rect 18365 16730 18370 16750
rect 18370 16730 18390 16750
rect 18390 16730 18395 16750
rect 18365 16725 18395 16730
rect 18445 16750 18475 16755
rect 18445 16730 18450 16750
rect 18450 16730 18470 16750
rect 18470 16730 18475 16750
rect 18445 16725 18475 16730
rect 18525 16750 18555 16755
rect 18525 16730 18530 16750
rect 18530 16730 18550 16750
rect 18550 16730 18555 16750
rect 18525 16725 18555 16730
rect 18605 16750 18635 16755
rect 18605 16730 18610 16750
rect 18610 16730 18630 16750
rect 18630 16730 18635 16750
rect 18605 16725 18635 16730
rect 18685 16750 18715 16755
rect 18685 16730 18690 16750
rect 18690 16730 18710 16750
rect 18710 16730 18715 16750
rect 18685 16725 18715 16730
rect 18765 16750 18795 16755
rect 18765 16730 18770 16750
rect 18770 16730 18790 16750
rect 18790 16730 18795 16750
rect 18765 16725 18795 16730
rect 18845 16750 18875 16755
rect 18845 16730 18850 16750
rect 18850 16730 18870 16750
rect 18870 16730 18875 16750
rect 18845 16725 18875 16730
rect 18925 16750 18955 16755
rect 18925 16730 18930 16750
rect 18930 16730 18950 16750
rect 18950 16730 18955 16750
rect 18925 16725 18955 16730
rect 19005 16750 19035 16755
rect 19005 16730 19010 16750
rect 19010 16730 19030 16750
rect 19030 16730 19035 16750
rect 19005 16725 19035 16730
rect 19085 16750 19115 16755
rect 19085 16730 19090 16750
rect 19090 16730 19110 16750
rect 19110 16730 19115 16750
rect 19085 16725 19115 16730
rect 19165 16750 19195 16755
rect 19165 16730 19170 16750
rect 19170 16730 19190 16750
rect 19190 16730 19195 16750
rect 19165 16725 19195 16730
rect 19245 16750 19275 16755
rect 19245 16730 19250 16750
rect 19250 16730 19270 16750
rect 19270 16730 19275 16750
rect 19245 16725 19275 16730
rect 19325 16750 19355 16755
rect 19325 16730 19330 16750
rect 19330 16730 19350 16750
rect 19350 16730 19355 16750
rect 19325 16725 19355 16730
rect 19405 16750 19435 16755
rect 19405 16730 19410 16750
rect 19410 16730 19430 16750
rect 19430 16730 19435 16750
rect 19405 16725 19435 16730
rect 19485 16750 19515 16755
rect 19485 16730 19490 16750
rect 19490 16730 19510 16750
rect 19510 16730 19515 16750
rect 19485 16725 19515 16730
rect 19565 16750 19595 16755
rect 19565 16730 19570 16750
rect 19570 16730 19590 16750
rect 19590 16730 19595 16750
rect 19565 16725 19595 16730
rect 19645 16750 19675 16755
rect 19645 16730 19650 16750
rect 19650 16730 19670 16750
rect 19670 16730 19675 16750
rect 19645 16725 19675 16730
rect 19725 16750 19755 16755
rect 19725 16730 19730 16750
rect 19730 16730 19750 16750
rect 19750 16730 19755 16750
rect 19725 16725 19755 16730
rect 19805 16750 19835 16755
rect 19805 16730 19810 16750
rect 19810 16730 19830 16750
rect 19830 16730 19835 16750
rect 19805 16725 19835 16730
rect 19885 16750 19915 16755
rect 19885 16730 19890 16750
rect 19890 16730 19910 16750
rect 19910 16730 19915 16750
rect 19885 16725 19915 16730
rect 19965 16750 19995 16755
rect 19965 16730 19970 16750
rect 19970 16730 19990 16750
rect 19990 16730 19995 16750
rect 19965 16725 19995 16730
rect 20045 16750 20075 16755
rect 20045 16730 20050 16750
rect 20050 16730 20070 16750
rect 20070 16730 20075 16750
rect 20045 16725 20075 16730
rect 20125 16750 20155 16755
rect 20125 16730 20130 16750
rect 20130 16730 20150 16750
rect 20150 16730 20155 16750
rect 20125 16725 20155 16730
rect 20205 16750 20235 16755
rect 20205 16730 20210 16750
rect 20210 16730 20230 16750
rect 20230 16730 20235 16750
rect 20205 16725 20235 16730
rect 20285 16750 20315 16755
rect 20285 16730 20290 16750
rect 20290 16730 20310 16750
rect 20310 16730 20315 16750
rect 20285 16725 20315 16730
rect 20365 16750 20395 16755
rect 20365 16730 20370 16750
rect 20370 16730 20390 16750
rect 20390 16730 20395 16750
rect 20365 16725 20395 16730
rect 20445 16750 20475 16755
rect 20445 16730 20450 16750
rect 20450 16730 20470 16750
rect 20470 16730 20475 16750
rect 20445 16725 20475 16730
rect 20525 16750 20555 16755
rect 20525 16730 20530 16750
rect 20530 16730 20550 16750
rect 20550 16730 20555 16750
rect 20525 16725 20555 16730
rect 20605 16750 20635 16755
rect 20605 16730 20610 16750
rect 20610 16730 20630 16750
rect 20630 16730 20635 16750
rect 20605 16725 20635 16730
rect 20685 16750 20715 16755
rect 20685 16730 20690 16750
rect 20690 16730 20710 16750
rect 20710 16730 20715 16750
rect 20685 16725 20715 16730
rect 20765 16750 20795 16755
rect 20765 16730 20770 16750
rect 20770 16730 20790 16750
rect 20790 16730 20795 16750
rect 20765 16725 20795 16730
rect 20845 16750 20875 16755
rect 20845 16730 20850 16750
rect 20850 16730 20870 16750
rect 20870 16730 20875 16750
rect 20845 16725 20875 16730
rect 20925 16750 20955 16755
rect 20925 16730 20930 16750
rect 20930 16730 20950 16750
rect 20950 16730 20955 16750
rect 20925 16725 20955 16730
rect 5 16670 35 16675
rect 5 16650 10 16670
rect 10 16650 30 16670
rect 30 16650 35 16670
rect 5 16645 35 16650
rect 85 16670 115 16675
rect 85 16650 90 16670
rect 90 16650 110 16670
rect 110 16650 115 16670
rect 85 16645 115 16650
rect 165 16670 195 16675
rect 165 16650 170 16670
rect 170 16650 190 16670
rect 190 16650 195 16670
rect 165 16645 195 16650
rect 245 16670 275 16675
rect 245 16650 250 16670
rect 250 16650 270 16670
rect 270 16650 275 16670
rect 245 16645 275 16650
rect 325 16670 355 16675
rect 325 16650 330 16670
rect 330 16650 350 16670
rect 350 16650 355 16670
rect 325 16645 355 16650
rect 405 16670 435 16675
rect 405 16650 410 16670
rect 410 16650 430 16670
rect 430 16650 435 16670
rect 405 16645 435 16650
rect 485 16670 515 16675
rect 485 16650 490 16670
rect 490 16650 510 16670
rect 510 16650 515 16670
rect 485 16645 515 16650
rect 565 16670 595 16675
rect 565 16650 570 16670
rect 570 16650 590 16670
rect 590 16650 595 16670
rect 565 16645 595 16650
rect 645 16670 675 16675
rect 645 16650 650 16670
rect 650 16650 670 16670
rect 670 16650 675 16670
rect 645 16645 675 16650
rect 725 16670 755 16675
rect 725 16650 730 16670
rect 730 16650 750 16670
rect 750 16650 755 16670
rect 725 16645 755 16650
rect 805 16670 835 16675
rect 805 16650 810 16670
rect 810 16650 830 16670
rect 830 16650 835 16670
rect 805 16645 835 16650
rect 885 16670 915 16675
rect 885 16650 890 16670
rect 890 16650 910 16670
rect 910 16650 915 16670
rect 885 16645 915 16650
rect 965 16670 995 16675
rect 965 16650 970 16670
rect 970 16650 990 16670
rect 990 16650 995 16670
rect 965 16645 995 16650
rect 1045 16670 1075 16675
rect 1045 16650 1050 16670
rect 1050 16650 1070 16670
rect 1070 16650 1075 16670
rect 1045 16645 1075 16650
rect 1125 16670 1155 16675
rect 1125 16650 1130 16670
rect 1130 16650 1150 16670
rect 1150 16650 1155 16670
rect 1125 16645 1155 16650
rect 1205 16670 1235 16675
rect 1205 16650 1210 16670
rect 1210 16650 1230 16670
rect 1230 16650 1235 16670
rect 1205 16645 1235 16650
rect 1285 16670 1315 16675
rect 1285 16650 1290 16670
rect 1290 16650 1310 16670
rect 1310 16650 1315 16670
rect 1285 16645 1315 16650
rect 1365 16670 1395 16675
rect 1365 16650 1370 16670
rect 1370 16650 1390 16670
rect 1390 16650 1395 16670
rect 1365 16645 1395 16650
rect 1445 16670 1475 16675
rect 1445 16650 1450 16670
rect 1450 16650 1470 16670
rect 1470 16650 1475 16670
rect 1445 16645 1475 16650
rect 1525 16670 1555 16675
rect 1525 16650 1530 16670
rect 1530 16650 1550 16670
rect 1550 16650 1555 16670
rect 1525 16645 1555 16650
rect 1605 16670 1635 16675
rect 1605 16650 1610 16670
rect 1610 16650 1630 16670
rect 1630 16650 1635 16670
rect 1605 16645 1635 16650
rect 1685 16670 1715 16675
rect 1685 16650 1690 16670
rect 1690 16650 1710 16670
rect 1710 16650 1715 16670
rect 1685 16645 1715 16650
rect 1765 16670 1795 16675
rect 1765 16650 1770 16670
rect 1770 16650 1790 16670
rect 1790 16650 1795 16670
rect 1765 16645 1795 16650
rect 1845 16670 1875 16675
rect 1845 16650 1850 16670
rect 1850 16650 1870 16670
rect 1870 16650 1875 16670
rect 1845 16645 1875 16650
rect 1925 16670 1955 16675
rect 1925 16650 1930 16670
rect 1930 16650 1950 16670
rect 1950 16650 1955 16670
rect 1925 16645 1955 16650
rect 2005 16670 2035 16675
rect 2005 16650 2010 16670
rect 2010 16650 2030 16670
rect 2030 16650 2035 16670
rect 2005 16645 2035 16650
rect 2085 16670 2115 16675
rect 2085 16650 2090 16670
rect 2090 16650 2110 16670
rect 2110 16650 2115 16670
rect 2085 16645 2115 16650
rect 2165 16670 2195 16675
rect 2165 16650 2170 16670
rect 2170 16650 2190 16670
rect 2190 16650 2195 16670
rect 2165 16645 2195 16650
rect 2245 16670 2275 16675
rect 2245 16650 2250 16670
rect 2250 16650 2270 16670
rect 2270 16650 2275 16670
rect 2245 16645 2275 16650
rect 2325 16670 2355 16675
rect 2325 16650 2330 16670
rect 2330 16650 2350 16670
rect 2350 16650 2355 16670
rect 2325 16645 2355 16650
rect 2405 16670 2435 16675
rect 2405 16650 2410 16670
rect 2410 16650 2430 16670
rect 2430 16650 2435 16670
rect 2405 16645 2435 16650
rect 2485 16670 2515 16675
rect 2485 16650 2490 16670
rect 2490 16650 2510 16670
rect 2510 16650 2515 16670
rect 2485 16645 2515 16650
rect 2565 16670 2595 16675
rect 2565 16650 2570 16670
rect 2570 16650 2590 16670
rect 2590 16650 2595 16670
rect 2565 16645 2595 16650
rect 2645 16670 2675 16675
rect 2645 16650 2650 16670
rect 2650 16650 2670 16670
rect 2670 16650 2675 16670
rect 2645 16645 2675 16650
rect 2725 16670 2755 16675
rect 2725 16650 2730 16670
rect 2730 16650 2750 16670
rect 2750 16650 2755 16670
rect 2725 16645 2755 16650
rect 2805 16670 2835 16675
rect 2805 16650 2810 16670
rect 2810 16650 2830 16670
rect 2830 16650 2835 16670
rect 2805 16645 2835 16650
rect 2885 16670 2915 16675
rect 2885 16650 2890 16670
rect 2890 16650 2910 16670
rect 2910 16650 2915 16670
rect 2885 16645 2915 16650
rect 2965 16670 2995 16675
rect 2965 16650 2970 16670
rect 2970 16650 2990 16670
rect 2990 16650 2995 16670
rect 2965 16645 2995 16650
rect 3045 16670 3075 16675
rect 3045 16650 3050 16670
rect 3050 16650 3070 16670
rect 3070 16650 3075 16670
rect 3045 16645 3075 16650
rect 3125 16670 3155 16675
rect 3125 16650 3130 16670
rect 3130 16650 3150 16670
rect 3150 16650 3155 16670
rect 3125 16645 3155 16650
rect 3205 16670 3235 16675
rect 3205 16650 3210 16670
rect 3210 16650 3230 16670
rect 3230 16650 3235 16670
rect 3205 16645 3235 16650
rect 3285 16670 3315 16675
rect 3285 16650 3290 16670
rect 3290 16650 3310 16670
rect 3310 16650 3315 16670
rect 3285 16645 3315 16650
rect 3365 16670 3395 16675
rect 3365 16650 3370 16670
rect 3370 16650 3390 16670
rect 3390 16650 3395 16670
rect 3365 16645 3395 16650
rect 3445 16670 3475 16675
rect 3445 16650 3450 16670
rect 3450 16650 3470 16670
rect 3470 16650 3475 16670
rect 3445 16645 3475 16650
rect 3525 16670 3555 16675
rect 3525 16650 3530 16670
rect 3530 16650 3550 16670
rect 3550 16650 3555 16670
rect 3525 16645 3555 16650
rect 3605 16670 3635 16675
rect 3605 16650 3610 16670
rect 3610 16650 3630 16670
rect 3630 16650 3635 16670
rect 3605 16645 3635 16650
rect 3685 16670 3715 16675
rect 3685 16650 3690 16670
rect 3690 16650 3710 16670
rect 3710 16650 3715 16670
rect 3685 16645 3715 16650
rect 3765 16670 3795 16675
rect 3765 16650 3770 16670
rect 3770 16650 3790 16670
rect 3790 16650 3795 16670
rect 3765 16645 3795 16650
rect 3845 16670 3875 16675
rect 3845 16650 3850 16670
rect 3850 16650 3870 16670
rect 3870 16650 3875 16670
rect 3845 16645 3875 16650
rect 3925 16670 3955 16675
rect 3925 16650 3930 16670
rect 3930 16650 3950 16670
rect 3950 16650 3955 16670
rect 3925 16645 3955 16650
rect 4005 16670 4035 16675
rect 4005 16650 4010 16670
rect 4010 16650 4030 16670
rect 4030 16650 4035 16670
rect 4005 16645 4035 16650
rect 4085 16670 4115 16675
rect 4085 16650 4090 16670
rect 4090 16650 4110 16670
rect 4110 16650 4115 16670
rect 4085 16645 4115 16650
rect 4165 16670 4195 16675
rect 4165 16650 4170 16670
rect 4170 16650 4190 16670
rect 4190 16650 4195 16670
rect 4165 16645 4195 16650
rect 6245 16670 6275 16675
rect 6245 16650 6250 16670
rect 6250 16650 6270 16670
rect 6270 16650 6275 16670
rect 6245 16645 6275 16650
rect 6325 16670 6355 16675
rect 6325 16650 6330 16670
rect 6330 16650 6350 16670
rect 6350 16650 6355 16670
rect 6325 16645 6355 16650
rect 6405 16670 6435 16675
rect 6405 16650 6410 16670
rect 6410 16650 6430 16670
rect 6430 16650 6435 16670
rect 6405 16645 6435 16650
rect 6485 16670 6515 16675
rect 6485 16650 6490 16670
rect 6490 16650 6510 16670
rect 6510 16650 6515 16670
rect 6485 16645 6515 16650
rect 6565 16670 6595 16675
rect 6565 16650 6570 16670
rect 6570 16650 6590 16670
rect 6590 16650 6595 16670
rect 6565 16645 6595 16650
rect 6645 16670 6675 16675
rect 6645 16650 6650 16670
rect 6650 16650 6670 16670
rect 6670 16650 6675 16670
rect 6645 16645 6675 16650
rect 6725 16670 6755 16675
rect 6725 16650 6730 16670
rect 6730 16650 6750 16670
rect 6750 16650 6755 16670
rect 6725 16645 6755 16650
rect 6805 16670 6835 16675
rect 6805 16650 6810 16670
rect 6810 16650 6830 16670
rect 6830 16650 6835 16670
rect 6805 16645 6835 16650
rect 6885 16670 6915 16675
rect 6885 16650 6890 16670
rect 6890 16650 6910 16670
rect 6910 16650 6915 16670
rect 6885 16645 6915 16650
rect 6965 16670 6995 16675
rect 6965 16650 6970 16670
rect 6970 16650 6990 16670
rect 6990 16650 6995 16670
rect 6965 16645 6995 16650
rect 7045 16670 7075 16675
rect 7045 16650 7050 16670
rect 7050 16650 7070 16670
rect 7070 16650 7075 16670
rect 7045 16645 7075 16650
rect 7125 16670 7155 16675
rect 7125 16650 7130 16670
rect 7130 16650 7150 16670
rect 7150 16650 7155 16670
rect 7125 16645 7155 16650
rect 7205 16670 7235 16675
rect 7205 16650 7210 16670
rect 7210 16650 7230 16670
rect 7230 16650 7235 16670
rect 7205 16645 7235 16650
rect 7285 16670 7315 16675
rect 7285 16650 7290 16670
rect 7290 16650 7310 16670
rect 7310 16650 7315 16670
rect 7285 16645 7315 16650
rect 7365 16670 7395 16675
rect 7365 16650 7370 16670
rect 7370 16650 7390 16670
rect 7390 16650 7395 16670
rect 7365 16645 7395 16650
rect 7445 16670 7475 16675
rect 7445 16650 7450 16670
rect 7450 16650 7470 16670
rect 7470 16650 7475 16670
rect 7445 16645 7475 16650
rect 7525 16670 7555 16675
rect 7525 16650 7530 16670
rect 7530 16650 7550 16670
rect 7550 16650 7555 16670
rect 7525 16645 7555 16650
rect 7605 16670 7635 16675
rect 7605 16650 7610 16670
rect 7610 16650 7630 16670
rect 7630 16650 7635 16670
rect 7605 16645 7635 16650
rect 7685 16670 7715 16675
rect 7685 16650 7690 16670
rect 7690 16650 7710 16670
rect 7710 16650 7715 16670
rect 7685 16645 7715 16650
rect 7765 16670 7795 16675
rect 7765 16650 7770 16670
rect 7770 16650 7790 16670
rect 7790 16650 7795 16670
rect 7765 16645 7795 16650
rect 7845 16670 7875 16675
rect 7845 16650 7850 16670
rect 7850 16650 7870 16670
rect 7870 16650 7875 16670
rect 7845 16645 7875 16650
rect 7925 16670 7955 16675
rect 7925 16650 7930 16670
rect 7930 16650 7950 16670
rect 7950 16650 7955 16670
rect 7925 16645 7955 16650
rect 8005 16670 8035 16675
rect 8005 16650 8010 16670
rect 8010 16650 8030 16670
rect 8030 16650 8035 16670
rect 8005 16645 8035 16650
rect 8085 16670 8115 16675
rect 8085 16650 8090 16670
rect 8090 16650 8110 16670
rect 8110 16650 8115 16670
rect 8085 16645 8115 16650
rect 8165 16670 8195 16675
rect 8165 16650 8170 16670
rect 8170 16650 8190 16670
rect 8190 16650 8195 16670
rect 8165 16645 8195 16650
rect 8245 16670 8275 16675
rect 8245 16650 8250 16670
rect 8250 16650 8270 16670
rect 8270 16650 8275 16670
rect 8245 16645 8275 16650
rect 8325 16670 8355 16675
rect 8325 16650 8330 16670
rect 8330 16650 8350 16670
rect 8350 16650 8355 16670
rect 8325 16645 8355 16650
rect 8405 16670 8435 16675
rect 8405 16650 8410 16670
rect 8410 16650 8430 16670
rect 8430 16650 8435 16670
rect 8405 16645 8435 16650
rect 8485 16670 8515 16675
rect 8485 16650 8490 16670
rect 8490 16650 8510 16670
rect 8510 16650 8515 16670
rect 8485 16645 8515 16650
rect 8565 16670 8595 16675
rect 8565 16650 8570 16670
rect 8570 16650 8590 16670
rect 8590 16650 8595 16670
rect 8565 16645 8595 16650
rect 8645 16670 8675 16675
rect 8645 16650 8650 16670
rect 8650 16650 8670 16670
rect 8670 16650 8675 16670
rect 8645 16645 8675 16650
rect 8725 16670 8755 16675
rect 8725 16650 8730 16670
rect 8730 16650 8750 16670
rect 8750 16650 8755 16670
rect 8725 16645 8755 16650
rect 8805 16670 8835 16675
rect 8805 16650 8810 16670
rect 8810 16650 8830 16670
rect 8830 16650 8835 16670
rect 8805 16645 8835 16650
rect 8885 16670 8915 16675
rect 8885 16650 8890 16670
rect 8890 16650 8910 16670
rect 8910 16650 8915 16670
rect 8885 16645 8915 16650
rect 8965 16670 8995 16675
rect 8965 16650 8970 16670
rect 8970 16650 8990 16670
rect 8990 16650 8995 16670
rect 8965 16645 8995 16650
rect 9045 16670 9075 16675
rect 9045 16650 9050 16670
rect 9050 16650 9070 16670
rect 9070 16650 9075 16670
rect 9045 16645 9075 16650
rect 9125 16670 9155 16675
rect 9125 16650 9130 16670
rect 9130 16650 9150 16670
rect 9150 16650 9155 16670
rect 9125 16645 9155 16650
rect 9205 16670 9235 16675
rect 9205 16650 9210 16670
rect 9210 16650 9230 16670
rect 9230 16650 9235 16670
rect 9205 16645 9235 16650
rect 9285 16670 9315 16675
rect 9285 16650 9290 16670
rect 9290 16650 9310 16670
rect 9310 16650 9315 16670
rect 9285 16645 9315 16650
rect 9365 16670 9395 16675
rect 9365 16650 9370 16670
rect 9370 16650 9390 16670
rect 9390 16650 9395 16670
rect 9365 16645 9395 16650
rect 9445 16670 9475 16675
rect 9445 16650 9450 16670
rect 9450 16650 9470 16670
rect 9470 16650 9475 16670
rect 9445 16645 9475 16650
rect 11565 16670 11595 16675
rect 11565 16650 11570 16670
rect 11570 16650 11590 16670
rect 11590 16650 11595 16670
rect 11565 16645 11595 16650
rect 11645 16670 11675 16675
rect 11645 16650 11650 16670
rect 11650 16650 11670 16670
rect 11670 16650 11675 16670
rect 11645 16645 11675 16650
rect 11725 16670 11755 16675
rect 11725 16650 11730 16670
rect 11730 16650 11750 16670
rect 11750 16650 11755 16670
rect 11725 16645 11755 16650
rect 11805 16670 11835 16675
rect 11805 16650 11810 16670
rect 11810 16650 11830 16670
rect 11830 16650 11835 16670
rect 11805 16645 11835 16650
rect 11885 16670 11915 16675
rect 11885 16650 11890 16670
rect 11890 16650 11910 16670
rect 11910 16650 11915 16670
rect 11885 16645 11915 16650
rect 11965 16670 11995 16675
rect 11965 16650 11970 16670
rect 11970 16650 11990 16670
rect 11990 16650 11995 16670
rect 11965 16645 11995 16650
rect 12045 16670 12075 16675
rect 12045 16650 12050 16670
rect 12050 16650 12070 16670
rect 12070 16650 12075 16670
rect 12045 16645 12075 16650
rect 12125 16670 12155 16675
rect 12125 16650 12130 16670
rect 12130 16650 12150 16670
rect 12150 16650 12155 16670
rect 12125 16645 12155 16650
rect 12205 16670 12235 16675
rect 12205 16650 12210 16670
rect 12210 16650 12230 16670
rect 12230 16650 12235 16670
rect 12205 16645 12235 16650
rect 12285 16670 12315 16675
rect 12285 16650 12290 16670
rect 12290 16650 12310 16670
rect 12310 16650 12315 16670
rect 12285 16645 12315 16650
rect 12365 16670 12395 16675
rect 12365 16650 12370 16670
rect 12370 16650 12390 16670
rect 12390 16650 12395 16670
rect 12365 16645 12395 16650
rect 12445 16670 12475 16675
rect 12445 16650 12450 16670
rect 12450 16650 12470 16670
rect 12470 16650 12475 16670
rect 12445 16645 12475 16650
rect 12525 16670 12555 16675
rect 12525 16650 12530 16670
rect 12530 16650 12550 16670
rect 12550 16650 12555 16670
rect 12525 16645 12555 16650
rect 12605 16670 12635 16675
rect 12605 16650 12610 16670
rect 12610 16650 12630 16670
rect 12630 16650 12635 16670
rect 12605 16645 12635 16650
rect 12685 16670 12715 16675
rect 12685 16650 12690 16670
rect 12690 16650 12710 16670
rect 12710 16650 12715 16670
rect 12685 16645 12715 16650
rect 12765 16670 12795 16675
rect 12765 16650 12770 16670
rect 12770 16650 12790 16670
rect 12790 16650 12795 16670
rect 12765 16645 12795 16650
rect 12845 16670 12875 16675
rect 12845 16650 12850 16670
rect 12850 16650 12870 16670
rect 12870 16650 12875 16670
rect 12845 16645 12875 16650
rect 12925 16670 12955 16675
rect 12925 16650 12930 16670
rect 12930 16650 12950 16670
rect 12950 16650 12955 16670
rect 12925 16645 12955 16650
rect 13005 16670 13035 16675
rect 13005 16650 13010 16670
rect 13010 16650 13030 16670
rect 13030 16650 13035 16670
rect 13005 16645 13035 16650
rect 13085 16670 13115 16675
rect 13085 16650 13090 16670
rect 13090 16650 13110 16670
rect 13110 16650 13115 16670
rect 13085 16645 13115 16650
rect 13165 16670 13195 16675
rect 13165 16650 13170 16670
rect 13170 16650 13190 16670
rect 13190 16650 13195 16670
rect 13165 16645 13195 16650
rect 13245 16670 13275 16675
rect 13245 16650 13250 16670
rect 13250 16650 13270 16670
rect 13270 16650 13275 16670
rect 13245 16645 13275 16650
rect 13325 16670 13355 16675
rect 13325 16650 13330 16670
rect 13330 16650 13350 16670
rect 13350 16650 13355 16670
rect 13325 16645 13355 16650
rect 13405 16670 13435 16675
rect 13405 16650 13410 16670
rect 13410 16650 13430 16670
rect 13430 16650 13435 16670
rect 13405 16645 13435 16650
rect 13485 16670 13515 16675
rect 13485 16650 13490 16670
rect 13490 16650 13510 16670
rect 13510 16650 13515 16670
rect 13485 16645 13515 16650
rect 13565 16670 13595 16675
rect 13565 16650 13570 16670
rect 13570 16650 13590 16670
rect 13590 16650 13595 16670
rect 13565 16645 13595 16650
rect 13645 16670 13675 16675
rect 13645 16650 13650 16670
rect 13650 16650 13670 16670
rect 13670 16650 13675 16670
rect 13645 16645 13675 16650
rect 13725 16670 13755 16675
rect 13725 16650 13730 16670
rect 13730 16650 13750 16670
rect 13750 16650 13755 16670
rect 13725 16645 13755 16650
rect 13805 16670 13835 16675
rect 13805 16650 13810 16670
rect 13810 16650 13830 16670
rect 13830 16650 13835 16670
rect 13805 16645 13835 16650
rect 13885 16670 13915 16675
rect 13885 16650 13890 16670
rect 13890 16650 13910 16670
rect 13910 16650 13915 16670
rect 13885 16645 13915 16650
rect 13965 16670 13995 16675
rect 13965 16650 13970 16670
rect 13970 16650 13990 16670
rect 13990 16650 13995 16670
rect 13965 16645 13995 16650
rect 14045 16670 14075 16675
rect 14045 16650 14050 16670
rect 14050 16650 14070 16670
rect 14070 16650 14075 16670
rect 14045 16645 14075 16650
rect 14125 16670 14155 16675
rect 14125 16650 14130 16670
rect 14130 16650 14150 16670
rect 14150 16650 14155 16670
rect 14125 16645 14155 16650
rect 14205 16670 14235 16675
rect 14205 16650 14210 16670
rect 14210 16650 14230 16670
rect 14230 16650 14235 16670
rect 14205 16645 14235 16650
rect 14285 16670 14315 16675
rect 14285 16650 14290 16670
rect 14290 16650 14310 16670
rect 14310 16650 14315 16670
rect 14285 16645 14315 16650
rect 14365 16670 14395 16675
rect 14365 16650 14370 16670
rect 14370 16650 14390 16670
rect 14390 16650 14395 16670
rect 14365 16645 14395 16650
rect 14445 16670 14475 16675
rect 14445 16650 14450 16670
rect 14450 16650 14470 16670
rect 14470 16650 14475 16670
rect 14445 16645 14475 16650
rect 14525 16670 14555 16675
rect 14525 16650 14530 16670
rect 14530 16650 14550 16670
rect 14550 16650 14555 16670
rect 14525 16645 14555 16650
rect 14605 16670 14635 16675
rect 14605 16650 14610 16670
rect 14610 16650 14630 16670
rect 14630 16650 14635 16670
rect 14605 16645 14635 16650
rect 14685 16670 14715 16675
rect 14685 16650 14690 16670
rect 14690 16650 14710 16670
rect 14710 16650 14715 16670
rect 14685 16645 14715 16650
rect 16765 16670 16795 16675
rect 16765 16650 16770 16670
rect 16770 16650 16790 16670
rect 16790 16650 16795 16670
rect 16765 16645 16795 16650
rect 16845 16670 16875 16675
rect 16845 16650 16850 16670
rect 16850 16650 16870 16670
rect 16870 16650 16875 16670
rect 16845 16645 16875 16650
rect 16925 16670 16955 16675
rect 16925 16650 16930 16670
rect 16930 16650 16950 16670
rect 16950 16650 16955 16670
rect 16925 16645 16955 16650
rect 17005 16670 17035 16675
rect 17005 16650 17010 16670
rect 17010 16650 17030 16670
rect 17030 16650 17035 16670
rect 17005 16645 17035 16650
rect 17085 16670 17115 16675
rect 17085 16650 17090 16670
rect 17090 16650 17110 16670
rect 17110 16650 17115 16670
rect 17085 16645 17115 16650
rect 17165 16670 17195 16675
rect 17165 16650 17170 16670
rect 17170 16650 17190 16670
rect 17190 16650 17195 16670
rect 17165 16645 17195 16650
rect 17245 16670 17275 16675
rect 17245 16650 17250 16670
rect 17250 16650 17270 16670
rect 17270 16650 17275 16670
rect 17245 16645 17275 16650
rect 17325 16670 17355 16675
rect 17325 16650 17330 16670
rect 17330 16650 17350 16670
rect 17350 16650 17355 16670
rect 17325 16645 17355 16650
rect 17405 16670 17435 16675
rect 17405 16650 17410 16670
rect 17410 16650 17430 16670
rect 17430 16650 17435 16670
rect 17405 16645 17435 16650
rect 17485 16670 17515 16675
rect 17485 16650 17490 16670
rect 17490 16650 17510 16670
rect 17510 16650 17515 16670
rect 17485 16645 17515 16650
rect 17565 16670 17595 16675
rect 17565 16650 17570 16670
rect 17570 16650 17590 16670
rect 17590 16650 17595 16670
rect 17565 16645 17595 16650
rect 17645 16670 17675 16675
rect 17645 16650 17650 16670
rect 17650 16650 17670 16670
rect 17670 16650 17675 16670
rect 17645 16645 17675 16650
rect 17725 16670 17755 16675
rect 17725 16650 17730 16670
rect 17730 16650 17750 16670
rect 17750 16650 17755 16670
rect 17725 16645 17755 16650
rect 17805 16670 17835 16675
rect 17805 16650 17810 16670
rect 17810 16650 17830 16670
rect 17830 16650 17835 16670
rect 17805 16645 17835 16650
rect 17885 16670 17915 16675
rect 17885 16650 17890 16670
rect 17890 16650 17910 16670
rect 17910 16650 17915 16670
rect 17885 16645 17915 16650
rect 17965 16670 17995 16675
rect 17965 16650 17970 16670
rect 17970 16650 17990 16670
rect 17990 16650 17995 16670
rect 17965 16645 17995 16650
rect 18045 16670 18075 16675
rect 18045 16650 18050 16670
rect 18050 16650 18070 16670
rect 18070 16650 18075 16670
rect 18045 16645 18075 16650
rect 18125 16670 18155 16675
rect 18125 16650 18130 16670
rect 18130 16650 18150 16670
rect 18150 16650 18155 16670
rect 18125 16645 18155 16650
rect 18205 16670 18235 16675
rect 18205 16650 18210 16670
rect 18210 16650 18230 16670
rect 18230 16650 18235 16670
rect 18205 16645 18235 16650
rect 18285 16670 18315 16675
rect 18285 16650 18290 16670
rect 18290 16650 18310 16670
rect 18310 16650 18315 16670
rect 18285 16645 18315 16650
rect 18365 16670 18395 16675
rect 18365 16650 18370 16670
rect 18370 16650 18390 16670
rect 18390 16650 18395 16670
rect 18365 16645 18395 16650
rect 18445 16670 18475 16675
rect 18445 16650 18450 16670
rect 18450 16650 18470 16670
rect 18470 16650 18475 16670
rect 18445 16645 18475 16650
rect 18525 16670 18555 16675
rect 18525 16650 18530 16670
rect 18530 16650 18550 16670
rect 18550 16650 18555 16670
rect 18525 16645 18555 16650
rect 18605 16670 18635 16675
rect 18605 16650 18610 16670
rect 18610 16650 18630 16670
rect 18630 16650 18635 16670
rect 18605 16645 18635 16650
rect 18685 16670 18715 16675
rect 18685 16650 18690 16670
rect 18690 16650 18710 16670
rect 18710 16650 18715 16670
rect 18685 16645 18715 16650
rect 18765 16670 18795 16675
rect 18765 16650 18770 16670
rect 18770 16650 18790 16670
rect 18790 16650 18795 16670
rect 18765 16645 18795 16650
rect 18845 16670 18875 16675
rect 18845 16650 18850 16670
rect 18850 16650 18870 16670
rect 18870 16650 18875 16670
rect 18845 16645 18875 16650
rect 18925 16670 18955 16675
rect 18925 16650 18930 16670
rect 18930 16650 18950 16670
rect 18950 16650 18955 16670
rect 18925 16645 18955 16650
rect 19005 16670 19035 16675
rect 19005 16650 19010 16670
rect 19010 16650 19030 16670
rect 19030 16650 19035 16670
rect 19005 16645 19035 16650
rect 19085 16670 19115 16675
rect 19085 16650 19090 16670
rect 19090 16650 19110 16670
rect 19110 16650 19115 16670
rect 19085 16645 19115 16650
rect 19165 16670 19195 16675
rect 19165 16650 19170 16670
rect 19170 16650 19190 16670
rect 19190 16650 19195 16670
rect 19165 16645 19195 16650
rect 19245 16670 19275 16675
rect 19245 16650 19250 16670
rect 19250 16650 19270 16670
rect 19270 16650 19275 16670
rect 19245 16645 19275 16650
rect 19325 16670 19355 16675
rect 19325 16650 19330 16670
rect 19330 16650 19350 16670
rect 19350 16650 19355 16670
rect 19325 16645 19355 16650
rect 19405 16670 19435 16675
rect 19405 16650 19410 16670
rect 19410 16650 19430 16670
rect 19430 16650 19435 16670
rect 19405 16645 19435 16650
rect 19485 16670 19515 16675
rect 19485 16650 19490 16670
rect 19490 16650 19510 16670
rect 19510 16650 19515 16670
rect 19485 16645 19515 16650
rect 19565 16670 19595 16675
rect 19565 16650 19570 16670
rect 19570 16650 19590 16670
rect 19590 16650 19595 16670
rect 19565 16645 19595 16650
rect 19645 16670 19675 16675
rect 19645 16650 19650 16670
rect 19650 16650 19670 16670
rect 19670 16650 19675 16670
rect 19645 16645 19675 16650
rect 19725 16670 19755 16675
rect 19725 16650 19730 16670
rect 19730 16650 19750 16670
rect 19750 16650 19755 16670
rect 19725 16645 19755 16650
rect 19805 16670 19835 16675
rect 19805 16650 19810 16670
rect 19810 16650 19830 16670
rect 19830 16650 19835 16670
rect 19805 16645 19835 16650
rect 19885 16670 19915 16675
rect 19885 16650 19890 16670
rect 19890 16650 19910 16670
rect 19910 16650 19915 16670
rect 19885 16645 19915 16650
rect 19965 16670 19995 16675
rect 19965 16650 19970 16670
rect 19970 16650 19990 16670
rect 19990 16650 19995 16670
rect 19965 16645 19995 16650
rect 20045 16670 20075 16675
rect 20045 16650 20050 16670
rect 20050 16650 20070 16670
rect 20070 16650 20075 16670
rect 20045 16645 20075 16650
rect 20125 16670 20155 16675
rect 20125 16650 20130 16670
rect 20130 16650 20150 16670
rect 20150 16650 20155 16670
rect 20125 16645 20155 16650
rect 20205 16670 20235 16675
rect 20205 16650 20210 16670
rect 20210 16650 20230 16670
rect 20230 16650 20235 16670
rect 20205 16645 20235 16650
rect 20285 16670 20315 16675
rect 20285 16650 20290 16670
rect 20290 16650 20310 16670
rect 20310 16650 20315 16670
rect 20285 16645 20315 16650
rect 20365 16670 20395 16675
rect 20365 16650 20370 16670
rect 20370 16650 20390 16670
rect 20390 16650 20395 16670
rect 20365 16645 20395 16650
rect 20445 16670 20475 16675
rect 20445 16650 20450 16670
rect 20450 16650 20470 16670
rect 20470 16650 20475 16670
rect 20445 16645 20475 16650
rect 20525 16670 20555 16675
rect 20525 16650 20530 16670
rect 20530 16650 20550 16670
rect 20550 16650 20555 16670
rect 20525 16645 20555 16650
rect 20605 16670 20635 16675
rect 20605 16650 20610 16670
rect 20610 16650 20630 16670
rect 20630 16650 20635 16670
rect 20605 16645 20635 16650
rect 20685 16670 20715 16675
rect 20685 16650 20690 16670
rect 20690 16650 20710 16670
rect 20710 16650 20715 16670
rect 20685 16645 20715 16650
rect 20765 16670 20795 16675
rect 20765 16650 20770 16670
rect 20770 16650 20790 16670
rect 20790 16650 20795 16670
rect 20765 16645 20795 16650
rect 20845 16670 20875 16675
rect 20845 16650 20850 16670
rect 20850 16650 20870 16670
rect 20870 16650 20875 16670
rect 20845 16645 20875 16650
rect 20925 16670 20955 16675
rect 20925 16650 20930 16670
rect 20930 16650 20950 16670
rect 20950 16650 20955 16670
rect 20925 16645 20955 16650
rect 5 16510 35 16515
rect 5 16490 10 16510
rect 10 16490 30 16510
rect 30 16490 35 16510
rect 5 16485 35 16490
rect 85 16510 115 16515
rect 85 16490 90 16510
rect 90 16490 110 16510
rect 110 16490 115 16510
rect 85 16485 115 16490
rect 165 16510 195 16515
rect 165 16490 170 16510
rect 170 16490 190 16510
rect 190 16490 195 16510
rect 165 16485 195 16490
rect 245 16510 275 16515
rect 245 16490 250 16510
rect 250 16490 270 16510
rect 270 16490 275 16510
rect 245 16485 275 16490
rect 325 16510 355 16515
rect 325 16490 330 16510
rect 330 16490 350 16510
rect 350 16490 355 16510
rect 325 16485 355 16490
rect 405 16510 435 16515
rect 405 16490 410 16510
rect 410 16490 430 16510
rect 430 16490 435 16510
rect 405 16485 435 16490
rect 485 16510 515 16515
rect 485 16490 490 16510
rect 490 16490 510 16510
rect 510 16490 515 16510
rect 485 16485 515 16490
rect 565 16510 595 16515
rect 565 16490 570 16510
rect 570 16490 590 16510
rect 590 16490 595 16510
rect 565 16485 595 16490
rect 645 16510 675 16515
rect 645 16490 650 16510
rect 650 16490 670 16510
rect 670 16490 675 16510
rect 645 16485 675 16490
rect 725 16510 755 16515
rect 725 16490 730 16510
rect 730 16490 750 16510
rect 750 16490 755 16510
rect 725 16485 755 16490
rect 805 16510 835 16515
rect 805 16490 810 16510
rect 810 16490 830 16510
rect 830 16490 835 16510
rect 805 16485 835 16490
rect 885 16510 915 16515
rect 885 16490 890 16510
rect 890 16490 910 16510
rect 910 16490 915 16510
rect 885 16485 915 16490
rect 965 16510 995 16515
rect 965 16490 970 16510
rect 970 16490 990 16510
rect 990 16490 995 16510
rect 965 16485 995 16490
rect 1045 16510 1075 16515
rect 1045 16490 1050 16510
rect 1050 16490 1070 16510
rect 1070 16490 1075 16510
rect 1045 16485 1075 16490
rect 1125 16510 1155 16515
rect 1125 16490 1130 16510
rect 1130 16490 1150 16510
rect 1150 16490 1155 16510
rect 1125 16485 1155 16490
rect 1205 16510 1235 16515
rect 1205 16490 1210 16510
rect 1210 16490 1230 16510
rect 1230 16490 1235 16510
rect 1205 16485 1235 16490
rect 1285 16510 1315 16515
rect 1285 16490 1290 16510
rect 1290 16490 1310 16510
rect 1310 16490 1315 16510
rect 1285 16485 1315 16490
rect 1365 16510 1395 16515
rect 1365 16490 1370 16510
rect 1370 16490 1390 16510
rect 1390 16490 1395 16510
rect 1365 16485 1395 16490
rect 1445 16510 1475 16515
rect 1445 16490 1450 16510
rect 1450 16490 1470 16510
rect 1470 16490 1475 16510
rect 1445 16485 1475 16490
rect 1525 16510 1555 16515
rect 1525 16490 1530 16510
rect 1530 16490 1550 16510
rect 1550 16490 1555 16510
rect 1525 16485 1555 16490
rect 1605 16510 1635 16515
rect 1605 16490 1610 16510
rect 1610 16490 1630 16510
rect 1630 16490 1635 16510
rect 1605 16485 1635 16490
rect 1685 16510 1715 16515
rect 1685 16490 1690 16510
rect 1690 16490 1710 16510
rect 1710 16490 1715 16510
rect 1685 16485 1715 16490
rect 1765 16510 1795 16515
rect 1765 16490 1770 16510
rect 1770 16490 1790 16510
rect 1790 16490 1795 16510
rect 1765 16485 1795 16490
rect 1845 16510 1875 16515
rect 1845 16490 1850 16510
rect 1850 16490 1870 16510
rect 1870 16490 1875 16510
rect 1845 16485 1875 16490
rect 1925 16510 1955 16515
rect 1925 16490 1930 16510
rect 1930 16490 1950 16510
rect 1950 16490 1955 16510
rect 1925 16485 1955 16490
rect 2005 16510 2035 16515
rect 2005 16490 2010 16510
rect 2010 16490 2030 16510
rect 2030 16490 2035 16510
rect 2005 16485 2035 16490
rect 2085 16510 2115 16515
rect 2085 16490 2090 16510
rect 2090 16490 2110 16510
rect 2110 16490 2115 16510
rect 2085 16485 2115 16490
rect 2165 16510 2195 16515
rect 2165 16490 2170 16510
rect 2170 16490 2190 16510
rect 2190 16490 2195 16510
rect 2165 16485 2195 16490
rect 2245 16510 2275 16515
rect 2245 16490 2250 16510
rect 2250 16490 2270 16510
rect 2270 16490 2275 16510
rect 2245 16485 2275 16490
rect 2325 16510 2355 16515
rect 2325 16490 2330 16510
rect 2330 16490 2350 16510
rect 2350 16490 2355 16510
rect 2325 16485 2355 16490
rect 2405 16510 2435 16515
rect 2405 16490 2410 16510
rect 2410 16490 2430 16510
rect 2430 16490 2435 16510
rect 2405 16485 2435 16490
rect 2485 16510 2515 16515
rect 2485 16490 2490 16510
rect 2490 16490 2510 16510
rect 2510 16490 2515 16510
rect 2485 16485 2515 16490
rect 2565 16510 2595 16515
rect 2565 16490 2570 16510
rect 2570 16490 2590 16510
rect 2590 16490 2595 16510
rect 2565 16485 2595 16490
rect 2645 16510 2675 16515
rect 2645 16490 2650 16510
rect 2650 16490 2670 16510
rect 2670 16490 2675 16510
rect 2645 16485 2675 16490
rect 2725 16510 2755 16515
rect 2725 16490 2730 16510
rect 2730 16490 2750 16510
rect 2750 16490 2755 16510
rect 2725 16485 2755 16490
rect 2805 16510 2835 16515
rect 2805 16490 2810 16510
rect 2810 16490 2830 16510
rect 2830 16490 2835 16510
rect 2805 16485 2835 16490
rect 2885 16510 2915 16515
rect 2885 16490 2890 16510
rect 2890 16490 2910 16510
rect 2910 16490 2915 16510
rect 2885 16485 2915 16490
rect 2965 16510 2995 16515
rect 2965 16490 2970 16510
rect 2970 16490 2990 16510
rect 2990 16490 2995 16510
rect 2965 16485 2995 16490
rect 3045 16510 3075 16515
rect 3045 16490 3050 16510
rect 3050 16490 3070 16510
rect 3070 16490 3075 16510
rect 3045 16485 3075 16490
rect 3125 16510 3155 16515
rect 3125 16490 3130 16510
rect 3130 16490 3150 16510
rect 3150 16490 3155 16510
rect 3125 16485 3155 16490
rect 3205 16510 3235 16515
rect 3205 16490 3210 16510
rect 3210 16490 3230 16510
rect 3230 16490 3235 16510
rect 3205 16485 3235 16490
rect 3285 16510 3315 16515
rect 3285 16490 3290 16510
rect 3290 16490 3310 16510
rect 3310 16490 3315 16510
rect 3285 16485 3315 16490
rect 3365 16510 3395 16515
rect 3365 16490 3370 16510
rect 3370 16490 3390 16510
rect 3390 16490 3395 16510
rect 3365 16485 3395 16490
rect 3445 16510 3475 16515
rect 3445 16490 3450 16510
rect 3450 16490 3470 16510
rect 3470 16490 3475 16510
rect 3445 16485 3475 16490
rect 3525 16510 3555 16515
rect 3525 16490 3530 16510
rect 3530 16490 3550 16510
rect 3550 16490 3555 16510
rect 3525 16485 3555 16490
rect 3605 16510 3635 16515
rect 3605 16490 3610 16510
rect 3610 16490 3630 16510
rect 3630 16490 3635 16510
rect 3605 16485 3635 16490
rect 3685 16510 3715 16515
rect 3685 16490 3690 16510
rect 3690 16490 3710 16510
rect 3710 16490 3715 16510
rect 3685 16485 3715 16490
rect 3765 16510 3795 16515
rect 3765 16490 3770 16510
rect 3770 16490 3790 16510
rect 3790 16490 3795 16510
rect 3765 16485 3795 16490
rect 3845 16510 3875 16515
rect 3845 16490 3850 16510
rect 3850 16490 3870 16510
rect 3870 16490 3875 16510
rect 3845 16485 3875 16490
rect 3925 16510 3955 16515
rect 3925 16490 3930 16510
rect 3930 16490 3950 16510
rect 3950 16490 3955 16510
rect 3925 16485 3955 16490
rect 4005 16510 4035 16515
rect 4005 16490 4010 16510
rect 4010 16490 4030 16510
rect 4030 16490 4035 16510
rect 4005 16485 4035 16490
rect 4085 16510 4115 16515
rect 4085 16490 4090 16510
rect 4090 16490 4110 16510
rect 4110 16490 4115 16510
rect 4085 16485 4115 16490
rect 4165 16510 4195 16515
rect 4165 16490 4170 16510
rect 4170 16490 4190 16510
rect 4190 16490 4195 16510
rect 4165 16485 4195 16490
rect 6245 16510 6275 16515
rect 6245 16490 6250 16510
rect 6250 16490 6270 16510
rect 6270 16490 6275 16510
rect 6245 16485 6275 16490
rect 6325 16510 6355 16515
rect 6325 16490 6330 16510
rect 6330 16490 6350 16510
rect 6350 16490 6355 16510
rect 6325 16485 6355 16490
rect 6405 16510 6435 16515
rect 6405 16490 6410 16510
rect 6410 16490 6430 16510
rect 6430 16490 6435 16510
rect 6405 16485 6435 16490
rect 6485 16510 6515 16515
rect 6485 16490 6490 16510
rect 6490 16490 6510 16510
rect 6510 16490 6515 16510
rect 6485 16485 6515 16490
rect 6565 16510 6595 16515
rect 6565 16490 6570 16510
rect 6570 16490 6590 16510
rect 6590 16490 6595 16510
rect 6565 16485 6595 16490
rect 6645 16510 6675 16515
rect 6645 16490 6650 16510
rect 6650 16490 6670 16510
rect 6670 16490 6675 16510
rect 6645 16485 6675 16490
rect 6725 16510 6755 16515
rect 6725 16490 6730 16510
rect 6730 16490 6750 16510
rect 6750 16490 6755 16510
rect 6725 16485 6755 16490
rect 6805 16510 6835 16515
rect 6805 16490 6810 16510
rect 6810 16490 6830 16510
rect 6830 16490 6835 16510
rect 6805 16485 6835 16490
rect 6885 16510 6915 16515
rect 6885 16490 6890 16510
rect 6890 16490 6910 16510
rect 6910 16490 6915 16510
rect 6885 16485 6915 16490
rect 6965 16510 6995 16515
rect 6965 16490 6970 16510
rect 6970 16490 6990 16510
rect 6990 16490 6995 16510
rect 6965 16485 6995 16490
rect 7045 16510 7075 16515
rect 7045 16490 7050 16510
rect 7050 16490 7070 16510
rect 7070 16490 7075 16510
rect 7045 16485 7075 16490
rect 7125 16510 7155 16515
rect 7125 16490 7130 16510
rect 7130 16490 7150 16510
rect 7150 16490 7155 16510
rect 7125 16485 7155 16490
rect 7205 16510 7235 16515
rect 7205 16490 7210 16510
rect 7210 16490 7230 16510
rect 7230 16490 7235 16510
rect 7205 16485 7235 16490
rect 7285 16510 7315 16515
rect 7285 16490 7290 16510
rect 7290 16490 7310 16510
rect 7310 16490 7315 16510
rect 7285 16485 7315 16490
rect 7365 16510 7395 16515
rect 7365 16490 7370 16510
rect 7370 16490 7390 16510
rect 7390 16490 7395 16510
rect 7365 16485 7395 16490
rect 7445 16510 7475 16515
rect 7445 16490 7450 16510
rect 7450 16490 7470 16510
rect 7470 16490 7475 16510
rect 7445 16485 7475 16490
rect 7525 16510 7555 16515
rect 7525 16490 7530 16510
rect 7530 16490 7550 16510
rect 7550 16490 7555 16510
rect 7525 16485 7555 16490
rect 7605 16510 7635 16515
rect 7605 16490 7610 16510
rect 7610 16490 7630 16510
rect 7630 16490 7635 16510
rect 7605 16485 7635 16490
rect 7685 16510 7715 16515
rect 7685 16490 7690 16510
rect 7690 16490 7710 16510
rect 7710 16490 7715 16510
rect 7685 16485 7715 16490
rect 7765 16510 7795 16515
rect 7765 16490 7770 16510
rect 7770 16490 7790 16510
rect 7790 16490 7795 16510
rect 7765 16485 7795 16490
rect 7845 16510 7875 16515
rect 7845 16490 7850 16510
rect 7850 16490 7870 16510
rect 7870 16490 7875 16510
rect 7845 16485 7875 16490
rect 7925 16510 7955 16515
rect 7925 16490 7930 16510
rect 7930 16490 7950 16510
rect 7950 16490 7955 16510
rect 7925 16485 7955 16490
rect 8005 16510 8035 16515
rect 8005 16490 8010 16510
rect 8010 16490 8030 16510
rect 8030 16490 8035 16510
rect 8005 16485 8035 16490
rect 8085 16510 8115 16515
rect 8085 16490 8090 16510
rect 8090 16490 8110 16510
rect 8110 16490 8115 16510
rect 8085 16485 8115 16490
rect 8165 16510 8195 16515
rect 8165 16490 8170 16510
rect 8170 16490 8190 16510
rect 8190 16490 8195 16510
rect 8165 16485 8195 16490
rect 8245 16510 8275 16515
rect 8245 16490 8250 16510
rect 8250 16490 8270 16510
rect 8270 16490 8275 16510
rect 8245 16485 8275 16490
rect 8325 16510 8355 16515
rect 8325 16490 8330 16510
rect 8330 16490 8350 16510
rect 8350 16490 8355 16510
rect 8325 16485 8355 16490
rect 8405 16510 8435 16515
rect 8405 16490 8410 16510
rect 8410 16490 8430 16510
rect 8430 16490 8435 16510
rect 8405 16485 8435 16490
rect 8485 16510 8515 16515
rect 8485 16490 8490 16510
rect 8490 16490 8510 16510
rect 8510 16490 8515 16510
rect 8485 16485 8515 16490
rect 8565 16510 8595 16515
rect 8565 16490 8570 16510
rect 8570 16490 8590 16510
rect 8590 16490 8595 16510
rect 8565 16485 8595 16490
rect 8645 16510 8675 16515
rect 8645 16490 8650 16510
rect 8650 16490 8670 16510
rect 8670 16490 8675 16510
rect 8645 16485 8675 16490
rect 8725 16510 8755 16515
rect 8725 16490 8730 16510
rect 8730 16490 8750 16510
rect 8750 16490 8755 16510
rect 8725 16485 8755 16490
rect 8805 16510 8835 16515
rect 8805 16490 8810 16510
rect 8810 16490 8830 16510
rect 8830 16490 8835 16510
rect 8805 16485 8835 16490
rect 8885 16510 8915 16515
rect 8885 16490 8890 16510
rect 8890 16490 8910 16510
rect 8910 16490 8915 16510
rect 8885 16485 8915 16490
rect 8965 16510 8995 16515
rect 8965 16490 8970 16510
rect 8970 16490 8990 16510
rect 8990 16490 8995 16510
rect 8965 16485 8995 16490
rect 9045 16510 9075 16515
rect 9045 16490 9050 16510
rect 9050 16490 9070 16510
rect 9070 16490 9075 16510
rect 9045 16485 9075 16490
rect 9125 16510 9155 16515
rect 9125 16490 9130 16510
rect 9130 16490 9150 16510
rect 9150 16490 9155 16510
rect 9125 16485 9155 16490
rect 9205 16510 9235 16515
rect 9205 16490 9210 16510
rect 9210 16490 9230 16510
rect 9230 16490 9235 16510
rect 9205 16485 9235 16490
rect 9285 16510 9315 16515
rect 9285 16490 9290 16510
rect 9290 16490 9310 16510
rect 9310 16490 9315 16510
rect 9285 16485 9315 16490
rect 9365 16510 9395 16515
rect 9365 16490 9370 16510
rect 9370 16490 9390 16510
rect 9390 16490 9395 16510
rect 9365 16485 9395 16490
rect 9445 16510 9475 16515
rect 9445 16490 9450 16510
rect 9450 16490 9470 16510
rect 9470 16490 9475 16510
rect 9445 16485 9475 16490
rect 11565 16510 11595 16515
rect 11565 16490 11570 16510
rect 11570 16490 11590 16510
rect 11590 16490 11595 16510
rect 11565 16485 11595 16490
rect 11645 16510 11675 16515
rect 11645 16490 11650 16510
rect 11650 16490 11670 16510
rect 11670 16490 11675 16510
rect 11645 16485 11675 16490
rect 11725 16510 11755 16515
rect 11725 16490 11730 16510
rect 11730 16490 11750 16510
rect 11750 16490 11755 16510
rect 11725 16485 11755 16490
rect 11805 16510 11835 16515
rect 11805 16490 11810 16510
rect 11810 16490 11830 16510
rect 11830 16490 11835 16510
rect 11805 16485 11835 16490
rect 11885 16510 11915 16515
rect 11885 16490 11890 16510
rect 11890 16490 11910 16510
rect 11910 16490 11915 16510
rect 11885 16485 11915 16490
rect 11965 16510 11995 16515
rect 11965 16490 11970 16510
rect 11970 16490 11990 16510
rect 11990 16490 11995 16510
rect 11965 16485 11995 16490
rect 12045 16510 12075 16515
rect 12045 16490 12050 16510
rect 12050 16490 12070 16510
rect 12070 16490 12075 16510
rect 12045 16485 12075 16490
rect 12125 16510 12155 16515
rect 12125 16490 12130 16510
rect 12130 16490 12150 16510
rect 12150 16490 12155 16510
rect 12125 16485 12155 16490
rect 12205 16510 12235 16515
rect 12205 16490 12210 16510
rect 12210 16490 12230 16510
rect 12230 16490 12235 16510
rect 12205 16485 12235 16490
rect 12285 16510 12315 16515
rect 12285 16490 12290 16510
rect 12290 16490 12310 16510
rect 12310 16490 12315 16510
rect 12285 16485 12315 16490
rect 12365 16510 12395 16515
rect 12365 16490 12370 16510
rect 12370 16490 12390 16510
rect 12390 16490 12395 16510
rect 12365 16485 12395 16490
rect 12445 16510 12475 16515
rect 12445 16490 12450 16510
rect 12450 16490 12470 16510
rect 12470 16490 12475 16510
rect 12445 16485 12475 16490
rect 12525 16510 12555 16515
rect 12525 16490 12530 16510
rect 12530 16490 12550 16510
rect 12550 16490 12555 16510
rect 12525 16485 12555 16490
rect 12605 16510 12635 16515
rect 12605 16490 12610 16510
rect 12610 16490 12630 16510
rect 12630 16490 12635 16510
rect 12605 16485 12635 16490
rect 12685 16510 12715 16515
rect 12685 16490 12690 16510
rect 12690 16490 12710 16510
rect 12710 16490 12715 16510
rect 12685 16485 12715 16490
rect 12765 16510 12795 16515
rect 12765 16490 12770 16510
rect 12770 16490 12790 16510
rect 12790 16490 12795 16510
rect 12765 16485 12795 16490
rect 12845 16510 12875 16515
rect 12845 16490 12850 16510
rect 12850 16490 12870 16510
rect 12870 16490 12875 16510
rect 12845 16485 12875 16490
rect 12925 16510 12955 16515
rect 12925 16490 12930 16510
rect 12930 16490 12950 16510
rect 12950 16490 12955 16510
rect 12925 16485 12955 16490
rect 13005 16510 13035 16515
rect 13005 16490 13010 16510
rect 13010 16490 13030 16510
rect 13030 16490 13035 16510
rect 13005 16485 13035 16490
rect 13085 16510 13115 16515
rect 13085 16490 13090 16510
rect 13090 16490 13110 16510
rect 13110 16490 13115 16510
rect 13085 16485 13115 16490
rect 13165 16510 13195 16515
rect 13165 16490 13170 16510
rect 13170 16490 13190 16510
rect 13190 16490 13195 16510
rect 13165 16485 13195 16490
rect 13245 16510 13275 16515
rect 13245 16490 13250 16510
rect 13250 16490 13270 16510
rect 13270 16490 13275 16510
rect 13245 16485 13275 16490
rect 13325 16510 13355 16515
rect 13325 16490 13330 16510
rect 13330 16490 13350 16510
rect 13350 16490 13355 16510
rect 13325 16485 13355 16490
rect 13405 16510 13435 16515
rect 13405 16490 13410 16510
rect 13410 16490 13430 16510
rect 13430 16490 13435 16510
rect 13405 16485 13435 16490
rect 13485 16510 13515 16515
rect 13485 16490 13490 16510
rect 13490 16490 13510 16510
rect 13510 16490 13515 16510
rect 13485 16485 13515 16490
rect 13565 16510 13595 16515
rect 13565 16490 13570 16510
rect 13570 16490 13590 16510
rect 13590 16490 13595 16510
rect 13565 16485 13595 16490
rect 13645 16510 13675 16515
rect 13645 16490 13650 16510
rect 13650 16490 13670 16510
rect 13670 16490 13675 16510
rect 13645 16485 13675 16490
rect 13725 16510 13755 16515
rect 13725 16490 13730 16510
rect 13730 16490 13750 16510
rect 13750 16490 13755 16510
rect 13725 16485 13755 16490
rect 13805 16510 13835 16515
rect 13805 16490 13810 16510
rect 13810 16490 13830 16510
rect 13830 16490 13835 16510
rect 13805 16485 13835 16490
rect 13885 16510 13915 16515
rect 13885 16490 13890 16510
rect 13890 16490 13910 16510
rect 13910 16490 13915 16510
rect 13885 16485 13915 16490
rect 13965 16510 13995 16515
rect 13965 16490 13970 16510
rect 13970 16490 13990 16510
rect 13990 16490 13995 16510
rect 13965 16485 13995 16490
rect 14045 16510 14075 16515
rect 14045 16490 14050 16510
rect 14050 16490 14070 16510
rect 14070 16490 14075 16510
rect 14045 16485 14075 16490
rect 14125 16510 14155 16515
rect 14125 16490 14130 16510
rect 14130 16490 14150 16510
rect 14150 16490 14155 16510
rect 14125 16485 14155 16490
rect 14205 16510 14235 16515
rect 14205 16490 14210 16510
rect 14210 16490 14230 16510
rect 14230 16490 14235 16510
rect 14205 16485 14235 16490
rect 14285 16510 14315 16515
rect 14285 16490 14290 16510
rect 14290 16490 14310 16510
rect 14310 16490 14315 16510
rect 14285 16485 14315 16490
rect 14365 16510 14395 16515
rect 14365 16490 14370 16510
rect 14370 16490 14390 16510
rect 14390 16490 14395 16510
rect 14365 16485 14395 16490
rect 14445 16510 14475 16515
rect 14445 16490 14450 16510
rect 14450 16490 14470 16510
rect 14470 16490 14475 16510
rect 14445 16485 14475 16490
rect 14525 16510 14555 16515
rect 14525 16490 14530 16510
rect 14530 16490 14550 16510
rect 14550 16490 14555 16510
rect 14525 16485 14555 16490
rect 14605 16510 14635 16515
rect 14605 16490 14610 16510
rect 14610 16490 14630 16510
rect 14630 16490 14635 16510
rect 14605 16485 14635 16490
rect 14685 16510 14715 16515
rect 14685 16490 14690 16510
rect 14690 16490 14710 16510
rect 14710 16490 14715 16510
rect 14685 16485 14715 16490
rect 16765 16510 16795 16515
rect 16765 16490 16770 16510
rect 16770 16490 16790 16510
rect 16790 16490 16795 16510
rect 16765 16485 16795 16490
rect 16845 16510 16875 16515
rect 16845 16490 16850 16510
rect 16850 16490 16870 16510
rect 16870 16490 16875 16510
rect 16845 16485 16875 16490
rect 16925 16510 16955 16515
rect 16925 16490 16930 16510
rect 16930 16490 16950 16510
rect 16950 16490 16955 16510
rect 16925 16485 16955 16490
rect 17005 16510 17035 16515
rect 17005 16490 17010 16510
rect 17010 16490 17030 16510
rect 17030 16490 17035 16510
rect 17005 16485 17035 16490
rect 17085 16510 17115 16515
rect 17085 16490 17090 16510
rect 17090 16490 17110 16510
rect 17110 16490 17115 16510
rect 17085 16485 17115 16490
rect 17165 16510 17195 16515
rect 17165 16490 17170 16510
rect 17170 16490 17190 16510
rect 17190 16490 17195 16510
rect 17165 16485 17195 16490
rect 17245 16510 17275 16515
rect 17245 16490 17250 16510
rect 17250 16490 17270 16510
rect 17270 16490 17275 16510
rect 17245 16485 17275 16490
rect 17325 16510 17355 16515
rect 17325 16490 17330 16510
rect 17330 16490 17350 16510
rect 17350 16490 17355 16510
rect 17325 16485 17355 16490
rect 17405 16510 17435 16515
rect 17405 16490 17410 16510
rect 17410 16490 17430 16510
rect 17430 16490 17435 16510
rect 17405 16485 17435 16490
rect 17485 16510 17515 16515
rect 17485 16490 17490 16510
rect 17490 16490 17510 16510
rect 17510 16490 17515 16510
rect 17485 16485 17515 16490
rect 17565 16510 17595 16515
rect 17565 16490 17570 16510
rect 17570 16490 17590 16510
rect 17590 16490 17595 16510
rect 17565 16485 17595 16490
rect 17645 16510 17675 16515
rect 17645 16490 17650 16510
rect 17650 16490 17670 16510
rect 17670 16490 17675 16510
rect 17645 16485 17675 16490
rect 17725 16510 17755 16515
rect 17725 16490 17730 16510
rect 17730 16490 17750 16510
rect 17750 16490 17755 16510
rect 17725 16485 17755 16490
rect 17805 16510 17835 16515
rect 17805 16490 17810 16510
rect 17810 16490 17830 16510
rect 17830 16490 17835 16510
rect 17805 16485 17835 16490
rect 17885 16510 17915 16515
rect 17885 16490 17890 16510
rect 17890 16490 17910 16510
rect 17910 16490 17915 16510
rect 17885 16485 17915 16490
rect 17965 16510 17995 16515
rect 17965 16490 17970 16510
rect 17970 16490 17990 16510
rect 17990 16490 17995 16510
rect 17965 16485 17995 16490
rect 18045 16510 18075 16515
rect 18045 16490 18050 16510
rect 18050 16490 18070 16510
rect 18070 16490 18075 16510
rect 18045 16485 18075 16490
rect 18125 16510 18155 16515
rect 18125 16490 18130 16510
rect 18130 16490 18150 16510
rect 18150 16490 18155 16510
rect 18125 16485 18155 16490
rect 18205 16510 18235 16515
rect 18205 16490 18210 16510
rect 18210 16490 18230 16510
rect 18230 16490 18235 16510
rect 18205 16485 18235 16490
rect 18285 16510 18315 16515
rect 18285 16490 18290 16510
rect 18290 16490 18310 16510
rect 18310 16490 18315 16510
rect 18285 16485 18315 16490
rect 18365 16510 18395 16515
rect 18365 16490 18370 16510
rect 18370 16490 18390 16510
rect 18390 16490 18395 16510
rect 18365 16485 18395 16490
rect 18445 16510 18475 16515
rect 18445 16490 18450 16510
rect 18450 16490 18470 16510
rect 18470 16490 18475 16510
rect 18445 16485 18475 16490
rect 18525 16510 18555 16515
rect 18525 16490 18530 16510
rect 18530 16490 18550 16510
rect 18550 16490 18555 16510
rect 18525 16485 18555 16490
rect 18605 16510 18635 16515
rect 18605 16490 18610 16510
rect 18610 16490 18630 16510
rect 18630 16490 18635 16510
rect 18605 16485 18635 16490
rect 18685 16510 18715 16515
rect 18685 16490 18690 16510
rect 18690 16490 18710 16510
rect 18710 16490 18715 16510
rect 18685 16485 18715 16490
rect 18765 16510 18795 16515
rect 18765 16490 18770 16510
rect 18770 16490 18790 16510
rect 18790 16490 18795 16510
rect 18765 16485 18795 16490
rect 18845 16510 18875 16515
rect 18845 16490 18850 16510
rect 18850 16490 18870 16510
rect 18870 16490 18875 16510
rect 18845 16485 18875 16490
rect 18925 16510 18955 16515
rect 18925 16490 18930 16510
rect 18930 16490 18950 16510
rect 18950 16490 18955 16510
rect 18925 16485 18955 16490
rect 19005 16510 19035 16515
rect 19005 16490 19010 16510
rect 19010 16490 19030 16510
rect 19030 16490 19035 16510
rect 19005 16485 19035 16490
rect 19085 16510 19115 16515
rect 19085 16490 19090 16510
rect 19090 16490 19110 16510
rect 19110 16490 19115 16510
rect 19085 16485 19115 16490
rect 19165 16510 19195 16515
rect 19165 16490 19170 16510
rect 19170 16490 19190 16510
rect 19190 16490 19195 16510
rect 19165 16485 19195 16490
rect 19245 16510 19275 16515
rect 19245 16490 19250 16510
rect 19250 16490 19270 16510
rect 19270 16490 19275 16510
rect 19245 16485 19275 16490
rect 19325 16510 19355 16515
rect 19325 16490 19330 16510
rect 19330 16490 19350 16510
rect 19350 16490 19355 16510
rect 19325 16485 19355 16490
rect 19405 16510 19435 16515
rect 19405 16490 19410 16510
rect 19410 16490 19430 16510
rect 19430 16490 19435 16510
rect 19405 16485 19435 16490
rect 19485 16510 19515 16515
rect 19485 16490 19490 16510
rect 19490 16490 19510 16510
rect 19510 16490 19515 16510
rect 19485 16485 19515 16490
rect 19565 16510 19595 16515
rect 19565 16490 19570 16510
rect 19570 16490 19590 16510
rect 19590 16490 19595 16510
rect 19565 16485 19595 16490
rect 19645 16510 19675 16515
rect 19645 16490 19650 16510
rect 19650 16490 19670 16510
rect 19670 16490 19675 16510
rect 19645 16485 19675 16490
rect 19725 16510 19755 16515
rect 19725 16490 19730 16510
rect 19730 16490 19750 16510
rect 19750 16490 19755 16510
rect 19725 16485 19755 16490
rect 19805 16510 19835 16515
rect 19805 16490 19810 16510
rect 19810 16490 19830 16510
rect 19830 16490 19835 16510
rect 19805 16485 19835 16490
rect 19885 16510 19915 16515
rect 19885 16490 19890 16510
rect 19890 16490 19910 16510
rect 19910 16490 19915 16510
rect 19885 16485 19915 16490
rect 19965 16510 19995 16515
rect 19965 16490 19970 16510
rect 19970 16490 19990 16510
rect 19990 16490 19995 16510
rect 19965 16485 19995 16490
rect 20045 16510 20075 16515
rect 20045 16490 20050 16510
rect 20050 16490 20070 16510
rect 20070 16490 20075 16510
rect 20045 16485 20075 16490
rect 20125 16510 20155 16515
rect 20125 16490 20130 16510
rect 20130 16490 20150 16510
rect 20150 16490 20155 16510
rect 20125 16485 20155 16490
rect 20205 16510 20235 16515
rect 20205 16490 20210 16510
rect 20210 16490 20230 16510
rect 20230 16490 20235 16510
rect 20205 16485 20235 16490
rect 20285 16510 20315 16515
rect 20285 16490 20290 16510
rect 20290 16490 20310 16510
rect 20310 16490 20315 16510
rect 20285 16485 20315 16490
rect 20365 16510 20395 16515
rect 20365 16490 20370 16510
rect 20370 16490 20390 16510
rect 20390 16490 20395 16510
rect 20365 16485 20395 16490
rect 20445 16510 20475 16515
rect 20445 16490 20450 16510
rect 20450 16490 20470 16510
rect 20470 16490 20475 16510
rect 20445 16485 20475 16490
rect 20525 16510 20555 16515
rect 20525 16490 20530 16510
rect 20530 16490 20550 16510
rect 20550 16490 20555 16510
rect 20525 16485 20555 16490
rect 20605 16510 20635 16515
rect 20605 16490 20610 16510
rect 20610 16490 20630 16510
rect 20630 16490 20635 16510
rect 20605 16485 20635 16490
rect 20685 16510 20715 16515
rect 20685 16490 20690 16510
rect 20690 16490 20710 16510
rect 20710 16490 20715 16510
rect 20685 16485 20715 16490
rect 20765 16510 20795 16515
rect 20765 16490 20770 16510
rect 20770 16490 20790 16510
rect 20790 16490 20795 16510
rect 20765 16485 20795 16490
rect 20845 16510 20875 16515
rect 20845 16490 20850 16510
rect 20850 16490 20870 16510
rect 20870 16490 20875 16510
rect 20845 16485 20875 16490
rect 20925 16510 20955 16515
rect 20925 16490 20930 16510
rect 20930 16490 20950 16510
rect 20950 16490 20955 16510
rect 20925 16485 20955 16490
rect 5 16430 35 16435
rect 5 16410 10 16430
rect 10 16410 30 16430
rect 30 16410 35 16430
rect 5 16405 35 16410
rect 85 16430 115 16435
rect 85 16410 90 16430
rect 90 16410 110 16430
rect 110 16410 115 16430
rect 85 16405 115 16410
rect 165 16430 195 16435
rect 165 16410 170 16430
rect 170 16410 190 16430
rect 190 16410 195 16430
rect 165 16405 195 16410
rect 245 16430 275 16435
rect 245 16410 250 16430
rect 250 16410 270 16430
rect 270 16410 275 16430
rect 245 16405 275 16410
rect 325 16430 355 16435
rect 325 16410 330 16430
rect 330 16410 350 16430
rect 350 16410 355 16430
rect 325 16405 355 16410
rect 405 16430 435 16435
rect 405 16410 410 16430
rect 410 16410 430 16430
rect 430 16410 435 16430
rect 405 16405 435 16410
rect 485 16430 515 16435
rect 485 16410 490 16430
rect 490 16410 510 16430
rect 510 16410 515 16430
rect 485 16405 515 16410
rect 565 16430 595 16435
rect 565 16410 570 16430
rect 570 16410 590 16430
rect 590 16410 595 16430
rect 565 16405 595 16410
rect 645 16430 675 16435
rect 645 16410 650 16430
rect 650 16410 670 16430
rect 670 16410 675 16430
rect 645 16405 675 16410
rect 725 16430 755 16435
rect 725 16410 730 16430
rect 730 16410 750 16430
rect 750 16410 755 16430
rect 725 16405 755 16410
rect 805 16430 835 16435
rect 805 16410 810 16430
rect 810 16410 830 16430
rect 830 16410 835 16430
rect 805 16405 835 16410
rect 885 16430 915 16435
rect 885 16410 890 16430
rect 890 16410 910 16430
rect 910 16410 915 16430
rect 885 16405 915 16410
rect 965 16430 995 16435
rect 965 16410 970 16430
rect 970 16410 990 16430
rect 990 16410 995 16430
rect 965 16405 995 16410
rect 1045 16430 1075 16435
rect 1045 16410 1050 16430
rect 1050 16410 1070 16430
rect 1070 16410 1075 16430
rect 1045 16405 1075 16410
rect 1125 16430 1155 16435
rect 1125 16410 1130 16430
rect 1130 16410 1150 16430
rect 1150 16410 1155 16430
rect 1125 16405 1155 16410
rect 1205 16430 1235 16435
rect 1205 16410 1210 16430
rect 1210 16410 1230 16430
rect 1230 16410 1235 16430
rect 1205 16405 1235 16410
rect 1285 16430 1315 16435
rect 1285 16410 1290 16430
rect 1290 16410 1310 16430
rect 1310 16410 1315 16430
rect 1285 16405 1315 16410
rect 1365 16430 1395 16435
rect 1365 16410 1370 16430
rect 1370 16410 1390 16430
rect 1390 16410 1395 16430
rect 1365 16405 1395 16410
rect 1445 16430 1475 16435
rect 1445 16410 1450 16430
rect 1450 16410 1470 16430
rect 1470 16410 1475 16430
rect 1445 16405 1475 16410
rect 1525 16430 1555 16435
rect 1525 16410 1530 16430
rect 1530 16410 1550 16430
rect 1550 16410 1555 16430
rect 1525 16405 1555 16410
rect 1605 16430 1635 16435
rect 1605 16410 1610 16430
rect 1610 16410 1630 16430
rect 1630 16410 1635 16430
rect 1605 16405 1635 16410
rect 1685 16430 1715 16435
rect 1685 16410 1690 16430
rect 1690 16410 1710 16430
rect 1710 16410 1715 16430
rect 1685 16405 1715 16410
rect 1765 16430 1795 16435
rect 1765 16410 1770 16430
rect 1770 16410 1790 16430
rect 1790 16410 1795 16430
rect 1765 16405 1795 16410
rect 1845 16430 1875 16435
rect 1845 16410 1850 16430
rect 1850 16410 1870 16430
rect 1870 16410 1875 16430
rect 1845 16405 1875 16410
rect 1925 16430 1955 16435
rect 1925 16410 1930 16430
rect 1930 16410 1950 16430
rect 1950 16410 1955 16430
rect 1925 16405 1955 16410
rect 2005 16430 2035 16435
rect 2005 16410 2010 16430
rect 2010 16410 2030 16430
rect 2030 16410 2035 16430
rect 2005 16405 2035 16410
rect 2085 16430 2115 16435
rect 2085 16410 2090 16430
rect 2090 16410 2110 16430
rect 2110 16410 2115 16430
rect 2085 16405 2115 16410
rect 2165 16430 2195 16435
rect 2165 16410 2170 16430
rect 2170 16410 2190 16430
rect 2190 16410 2195 16430
rect 2165 16405 2195 16410
rect 2245 16430 2275 16435
rect 2245 16410 2250 16430
rect 2250 16410 2270 16430
rect 2270 16410 2275 16430
rect 2245 16405 2275 16410
rect 2325 16430 2355 16435
rect 2325 16410 2330 16430
rect 2330 16410 2350 16430
rect 2350 16410 2355 16430
rect 2325 16405 2355 16410
rect 2405 16430 2435 16435
rect 2405 16410 2410 16430
rect 2410 16410 2430 16430
rect 2430 16410 2435 16430
rect 2405 16405 2435 16410
rect 2485 16430 2515 16435
rect 2485 16410 2490 16430
rect 2490 16410 2510 16430
rect 2510 16410 2515 16430
rect 2485 16405 2515 16410
rect 2565 16430 2595 16435
rect 2565 16410 2570 16430
rect 2570 16410 2590 16430
rect 2590 16410 2595 16430
rect 2565 16405 2595 16410
rect 2645 16430 2675 16435
rect 2645 16410 2650 16430
rect 2650 16410 2670 16430
rect 2670 16410 2675 16430
rect 2645 16405 2675 16410
rect 2725 16430 2755 16435
rect 2725 16410 2730 16430
rect 2730 16410 2750 16430
rect 2750 16410 2755 16430
rect 2725 16405 2755 16410
rect 2805 16430 2835 16435
rect 2805 16410 2810 16430
rect 2810 16410 2830 16430
rect 2830 16410 2835 16430
rect 2805 16405 2835 16410
rect 2885 16430 2915 16435
rect 2885 16410 2890 16430
rect 2890 16410 2910 16430
rect 2910 16410 2915 16430
rect 2885 16405 2915 16410
rect 2965 16430 2995 16435
rect 2965 16410 2970 16430
rect 2970 16410 2990 16430
rect 2990 16410 2995 16430
rect 2965 16405 2995 16410
rect 3045 16430 3075 16435
rect 3045 16410 3050 16430
rect 3050 16410 3070 16430
rect 3070 16410 3075 16430
rect 3045 16405 3075 16410
rect 3125 16430 3155 16435
rect 3125 16410 3130 16430
rect 3130 16410 3150 16430
rect 3150 16410 3155 16430
rect 3125 16405 3155 16410
rect 3205 16430 3235 16435
rect 3205 16410 3210 16430
rect 3210 16410 3230 16430
rect 3230 16410 3235 16430
rect 3205 16405 3235 16410
rect 3285 16430 3315 16435
rect 3285 16410 3290 16430
rect 3290 16410 3310 16430
rect 3310 16410 3315 16430
rect 3285 16405 3315 16410
rect 3365 16430 3395 16435
rect 3365 16410 3370 16430
rect 3370 16410 3390 16430
rect 3390 16410 3395 16430
rect 3365 16405 3395 16410
rect 3445 16430 3475 16435
rect 3445 16410 3450 16430
rect 3450 16410 3470 16430
rect 3470 16410 3475 16430
rect 3445 16405 3475 16410
rect 3525 16430 3555 16435
rect 3525 16410 3530 16430
rect 3530 16410 3550 16430
rect 3550 16410 3555 16430
rect 3525 16405 3555 16410
rect 3605 16430 3635 16435
rect 3605 16410 3610 16430
rect 3610 16410 3630 16430
rect 3630 16410 3635 16430
rect 3605 16405 3635 16410
rect 3685 16430 3715 16435
rect 3685 16410 3690 16430
rect 3690 16410 3710 16430
rect 3710 16410 3715 16430
rect 3685 16405 3715 16410
rect 3765 16430 3795 16435
rect 3765 16410 3770 16430
rect 3770 16410 3790 16430
rect 3790 16410 3795 16430
rect 3765 16405 3795 16410
rect 3845 16430 3875 16435
rect 3845 16410 3850 16430
rect 3850 16410 3870 16430
rect 3870 16410 3875 16430
rect 3845 16405 3875 16410
rect 3925 16430 3955 16435
rect 3925 16410 3930 16430
rect 3930 16410 3950 16430
rect 3950 16410 3955 16430
rect 3925 16405 3955 16410
rect 4005 16430 4035 16435
rect 4005 16410 4010 16430
rect 4010 16410 4030 16430
rect 4030 16410 4035 16430
rect 4005 16405 4035 16410
rect 4085 16430 4115 16435
rect 4085 16410 4090 16430
rect 4090 16410 4110 16430
rect 4110 16410 4115 16430
rect 4085 16405 4115 16410
rect 4165 16430 4195 16435
rect 4165 16410 4170 16430
rect 4170 16410 4190 16430
rect 4190 16410 4195 16430
rect 4165 16405 4195 16410
rect 6245 16430 6275 16435
rect 6245 16410 6250 16430
rect 6250 16410 6270 16430
rect 6270 16410 6275 16430
rect 6245 16405 6275 16410
rect 6325 16430 6355 16435
rect 6325 16410 6330 16430
rect 6330 16410 6350 16430
rect 6350 16410 6355 16430
rect 6325 16405 6355 16410
rect 6405 16430 6435 16435
rect 6405 16410 6410 16430
rect 6410 16410 6430 16430
rect 6430 16410 6435 16430
rect 6405 16405 6435 16410
rect 6485 16430 6515 16435
rect 6485 16410 6490 16430
rect 6490 16410 6510 16430
rect 6510 16410 6515 16430
rect 6485 16405 6515 16410
rect 6565 16430 6595 16435
rect 6565 16410 6570 16430
rect 6570 16410 6590 16430
rect 6590 16410 6595 16430
rect 6565 16405 6595 16410
rect 6645 16430 6675 16435
rect 6645 16410 6650 16430
rect 6650 16410 6670 16430
rect 6670 16410 6675 16430
rect 6645 16405 6675 16410
rect 6725 16430 6755 16435
rect 6725 16410 6730 16430
rect 6730 16410 6750 16430
rect 6750 16410 6755 16430
rect 6725 16405 6755 16410
rect 6805 16430 6835 16435
rect 6805 16410 6810 16430
rect 6810 16410 6830 16430
rect 6830 16410 6835 16430
rect 6805 16405 6835 16410
rect 6885 16430 6915 16435
rect 6885 16410 6890 16430
rect 6890 16410 6910 16430
rect 6910 16410 6915 16430
rect 6885 16405 6915 16410
rect 6965 16430 6995 16435
rect 6965 16410 6970 16430
rect 6970 16410 6990 16430
rect 6990 16410 6995 16430
rect 6965 16405 6995 16410
rect 7045 16430 7075 16435
rect 7045 16410 7050 16430
rect 7050 16410 7070 16430
rect 7070 16410 7075 16430
rect 7045 16405 7075 16410
rect 7125 16430 7155 16435
rect 7125 16410 7130 16430
rect 7130 16410 7150 16430
rect 7150 16410 7155 16430
rect 7125 16405 7155 16410
rect 7205 16430 7235 16435
rect 7205 16410 7210 16430
rect 7210 16410 7230 16430
rect 7230 16410 7235 16430
rect 7205 16405 7235 16410
rect 7285 16430 7315 16435
rect 7285 16410 7290 16430
rect 7290 16410 7310 16430
rect 7310 16410 7315 16430
rect 7285 16405 7315 16410
rect 7365 16430 7395 16435
rect 7365 16410 7370 16430
rect 7370 16410 7390 16430
rect 7390 16410 7395 16430
rect 7365 16405 7395 16410
rect 7445 16430 7475 16435
rect 7445 16410 7450 16430
rect 7450 16410 7470 16430
rect 7470 16410 7475 16430
rect 7445 16405 7475 16410
rect 7525 16430 7555 16435
rect 7525 16410 7530 16430
rect 7530 16410 7550 16430
rect 7550 16410 7555 16430
rect 7525 16405 7555 16410
rect 7605 16430 7635 16435
rect 7605 16410 7610 16430
rect 7610 16410 7630 16430
rect 7630 16410 7635 16430
rect 7605 16405 7635 16410
rect 7685 16430 7715 16435
rect 7685 16410 7690 16430
rect 7690 16410 7710 16430
rect 7710 16410 7715 16430
rect 7685 16405 7715 16410
rect 7765 16430 7795 16435
rect 7765 16410 7770 16430
rect 7770 16410 7790 16430
rect 7790 16410 7795 16430
rect 7765 16405 7795 16410
rect 7845 16430 7875 16435
rect 7845 16410 7850 16430
rect 7850 16410 7870 16430
rect 7870 16410 7875 16430
rect 7845 16405 7875 16410
rect 7925 16430 7955 16435
rect 7925 16410 7930 16430
rect 7930 16410 7950 16430
rect 7950 16410 7955 16430
rect 7925 16405 7955 16410
rect 8005 16430 8035 16435
rect 8005 16410 8010 16430
rect 8010 16410 8030 16430
rect 8030 16410 8035 16430
rect 8005 16405 8035 16410
rect 8085 16430 8115 16435
rect 8085 16410 8090 16430
rect 8090 16410 8110 16430
rect 8110 16410 8115 16430
rect 8085 16405 8115 16410
rect 8165 16430 8195 16435
rect 8165 16410 8170 16430
rect 8170 16410 8190 16430
rect 8190 16410 8195 16430
rect 8165 16405 8195 16410
rect 8245 16430 8275 16435
rect 8245 16410 8250 16430
rect 8250 16410 8270 16430
rect 8270 16410 8275 16430
rect 8245 16405 8275 16410
rect 8325 16430 8355 16435
rect 8325 16410 8330 16430
rect 8330 16410 8350 16430
rect 8350 16410 8355 16430
rect 8325 16405 8355 16410
rect 8405 16430 8435 16435
rect 8405 16410 8410 16430
rect 8410 16410 8430 16430
rect 8430 16410 8435 16430
rect 8405 16405 8435 16410
rect 8485 16430 8515 16435
rect 8485 16410 8490 16430
rect 8490 16410 8510 16430
rect 8510 16410 8515 16430
rect 8485 16405 8515 16410
rect 8565 16430 8595 16435
rect 8565 16410 8570 16430
rect 8570 16410 8590 16430
rect 8590 16410 8595 16430
rect 8565 16405 8595 16410
rect 8645 16430 8675 16435
rect 8645 16410 8650 16430
rect 8650 16410 8670 16430
rect 8670 16410 8675 16430
rect 8645 16405 8675 16410
rect 8725 16430 8755 16435
rect 8725 16410 8730 16430
rect 8730 16410 8750 16430
rect 8750 16410 8755 16430
rect 8725 16405 8755 16410
rect 8805 16430 8835 16435
rect 8805 16410 8810 16430
rect 8810 16410 8830 16430
rect 8830 16410 8835 16430
rect 8805 16405 8835 16410
rect 8885 16430 8915 16435
rect 8885 16410 8890 16430
rect 8890 16410 8910 16430
rect 8910 16410 8915 16430
rect 8885 16405 8915 16410
rect 8965 16430 8995 16435
rect 8965 16410 8970 16430
rect 8970 16410 8990 16430
rect 8990 16410 8995 16430
rect 8965 16405 8995 16410
rect 9045 16430 9075 16435
rect 9045 16410 9050 16430
rect 9050 16410 9070 16430
rect 9070 16410 9075 16430
rect 9045 16405 9075 16410
rect 9125 16430 9155 16435
rect 9125 16410 9130 16430
rect 9130 16410 9150 16430
rect 9150 16410 9155 16430
rect 9125 16405 9155 16410
rect 9205 16430 9235 16435
rect 9205 16410 9210 16430
rect 9210 16410 9230 16430
rect 9230 16410 9235 16430
rect 9205 16405 9235 16410
rect 9285 16430 9315 16435
rect 9285 16410 9290 16430
rect 9290 16410 9310 16430
rect 9310 16410 9315 16430
rect 9285 16405 9315 16410
rect 9365 16430 9395 16435
rect 9365 16410 9370 16430
rect 9370 16410 9390 16430
rect 9390 16410 9395 16430
rect 9365 16405 9395 16410
rect 9445 16430 9475 16435
rect 9445 16410 9450 16430
rect 9450 16410 9470 16430
rect 9470 16410 9475 16430
rect 9445 16405 9475 16410
rect 11565 16430 11595 16435
rect 11565 16410 11570 16430
rect 11570 16410 11590 16430
rect 11590 16410 11595 16430
rect 11565 16405 11595 16410
rect 11645 16430 11675 16435
rect 11645 16410 11650 16430
rect 11650 16410 11670 16430
rect 11670 16410 11675 16430
rect 11645 16405 11675 16410
rect 11725 16430 11755 16435
rect 11725 16410 11730 16430
rect 11730 16410 11750 16430
rect 11750 16410 11755 16430
rect 11725 16405 11755 16410
rect 11805 16430 11835 16435
rect 11805 16410 11810 16430
rect 11810 16410 11830 16430
rect 11830 16410 11835 16430
rect 11805 16405 11835 16410
rect 11885 16430 11915 16435
rect 11885 16410 11890 16430
rect 11890 16410 11910 16430
rect 11910 16410 11915 16430
rect 11885 16405 11915 16410
rect 11965 16430 11995 16435
rect 11965 16410 11970 16430
rect 11970 16410 11990 16430
rect 11990 16410 11995 16430
rect 11965 16405 11995 16410
rect 12045 16430 12075 16435
rect 12045 16410 12050 16430
rect 12050 16410 12070 16430
rect 12070 16410 12075 16430
rect 12045 16405 12075 16410
rect 12125 16430 12155 16435
rect 12125 16410 12130 16430
rect 12130 16410 12150 16430
rect 12150 16410 12155 16430
rect 12125 16405 12155 16410
rect 12205 16430 12235 16435
rect 12205 16410 12210 16430
rect 12210 16410 12230 16430
rect 12230 16410 12235 16430
rect 12205 16405 12235 16410
rect 12285 16430 12315 16435
rect 12285 16410 12290 16430
rect 12290 16410 12310 16430
rect 12310 16410 12315 16430
rect 12285 16405 12315 16410
rect 12365 16430 12395 16435
rect 12365 16410 12370 16430
rect 12370 16410 12390 16430
rect 12390 16410 12395 16430
rect 12365 16405 12395 16410
rect 12445 16430 12475 16435
rect 12445 16410 12450 16430
rect 12450 16410 12470 16430
rect 12470 16410 12475 16430
rect 12445 16405 12475 16410
rect 12525 16430 12555 16435
rect 12525 16410 12530 16430
rect 12530 16410 12550 16430
rect 12550 16410 12555 16430
rect 12525 16405 12555 16410
rect 12605 16430 12635 16435
rect 12605 16410 12610 16430
rect 12610 16410 12630 16430
rect 12630 16410 12635 16430
rect 12605 16405 12635 16410
rect 12685 16430 12715 16435
rect 12685 16410 12690 16430
rect 12690 16410 12710 16430
rect 12710 16410 12715 16430
rect 12685 16405 12715 16410
rect 12765 16430 12795 16435
rect 12765 16410 12770 16430
rect 12770 16410 12790 16430
rect 12790 16410 12795 16430
rect 12765 16405 12795 16410
rect 12845 16430 12875 16435
rect 12845 16410 12850 16430
rect 12850 16410 12870 16430
rect 12870 16410 12875 16430
rect 12845 16405 12875 16410
rect 12925 16430 12955 16435
rect 12925 16410 12930 16430
rect 12930 16410 12950 16430
rect 12950 16410 12955 16430
rect 12925 16405 12955 16410
rect 13005 16430 13035 16435
rect 13005 16410 13010 16430
rect 13010 16410 13030 16430
rect 13030 16410 13035 16430
rect 13005 16405 13035 16410
rect 13085 16430 13115 16435
rect 13085 16410 13090 16430
rect 13090 16410 13110 16430
rect 13110 16410 13115 16430
rect 13085 16405 13115 16410
rect 13165 16430 13195 16435
rect 13165 16410 13170 16430
rect 13170 16410 13190 16430
rect 13190 16410 13195 16430
rect 13165 16405 13195 16410
rect 13245 16430 13275 16435
rect 13245 16410 13250 16430
rect 13250 16410 13270 16430
rect 13270 16410 13275 16430
rect 13245 16405 13275 16410
rect 13325 16430 13355 16435
rect 13325 16410 13330 16430
rect 13330 16410 13350 16430
rect 13350 16410 13355 16430
rect 13325 16405 13355 16410
rect 13405 16430 13435 16435
rect 13405 16410 13410 16430
rect 13410 16410 13430 16430
rect 13430 16410 13435 16430
rect 13405 16405 13435 16410
rect 13485 16430 13515 16435
rect 13485 16410 13490 16430
rect 13490 16410 13510 16430
rect 13510 16410 13515 16430
rect 13485 16405 13515 16410
rect 13565 16430 13595 16435
rect 13565 16410 13570 16430
rect 13570 16410 13590 16430
rect 13590 16410 13595 16430
rect 13565 16405 13595 16410
rect 13645 16430 13675 16435
rect 13645 16410 13650 16430
rect 13650 16410 13670 16430
rect 13670 16410 13675 16430
rect 13645 16405 13675 16410
rect 13725 16430 13755 16435
rect 13725 16410 13730 16430
rect 13730 16410 13750 16430
rect 13750 16410 13755 16430
rect 13725 16405 13755 16410
rect 13805 16430 13835 16435
rect 13805 16410 13810 16430
rect 13810 16410 13830 16430
rect 13830 16410 13835 16430
rect 13805 16405 13835 16410
rect 13885 16430 13915 16435
rect 13885 16410 13890 16430
rect 13890 16410 13910 16430
rect 13910 16410 13915 16430
rect 13885 16405 13915 16410
rect 13965 16430 13995 16435
rect 13965 16410 13970 16430
rect 13970 16410 13990 16430
rect 13990 16410 13995 16430
rect 13965 16405 13995 16410
rect 14045 16430 14075 16435
rect 14045 16410 14050 16430
rect 14050 16410 14070 16430
rect 14070 16410 14075 16430
rect 14045 16405 14075 16410
rect 14125 16430 14155 16435
rect 14125 16410 14130 16430
rect 14130 16410 14150 16430
rect 14150 16410 14155 16430
rect 14125 16405 14155 16410
rect 14205 16430 14235 16435
rect 14205 16410 14210 16430
rect 14210 16410 14230 16430
rect 14230 16410 14235 16430
rect 14205 16405 14235 16410
rect 14285 16430 14315 16435
rect 14285 16410 14290 16430
rect 14290 16410 14310 16430
rect 14310 16410 14315 16430
rect 14285 16405 14315 16410
rect 14365 16430 14395 16435
rect 14365 16410 14370 16430
rect 14370 16410 14390 16430
rect 14390 16410 14395 16430
rect 14365 16405 14395 16410
rect 14445 16430 14475 16435
rect 14445 16410 14450 16430
rect 14450 16410 14470 16430
rect 14470 16410 14475 16430
rect 14445 16405 14475 16410
rect 14525 16430 14555 16435
rect 14525 16410 14530 16430
rect 14530 16410 14550 16430
rect 14550 16410 14555 16430
rect 14525 16405 14555 16410
rect 14605 16430 14635 16435
rect 14605 16410 14610 16430
rect 14610 16410 14630 16430
rect 14630 16410 14635 16430
rect 14605 16405 14635 16410
rect 14685 16430 14715 16435
rect 14685 16410 14690 16430
rect 14690 16410 14710 16430
rect 14710 16410 14715 16430
rect 14685 16405 14715 16410
rect 16765 16430 16795 16435
rect 16765 16410 16770 16430
rect 16770 16410 16790 16430
rect 16790 16410 16795 16430
rect 16765 16405 16795 16410
rect 16845 16430 16875 16435
rect 16845 16410 16850 16430
rect 16850 16410 16870 16430
rect 16870 16410 16875 16430
rect 16845 16405 16875 16410
rect 16925 16430 16955 16435
rect 16925 16410 16930 16430
rect 16930 16410 16950 16430
rect 16950 16410 16955 16430
rect 16925 16405 16955 16410
rect 17005 16430 17035 16435
rect 17005 16410 17010 16430
rect 17010 16410 17030 16430
rect 17030 16410 17035 16430
rect 17005 16405 17035 16410
rect 17085 16430 17115 16435
rect 17085 16410 17090 16430
rect 17090 16410 17110 16430
rect 17110 16410 17115 16430
rect 17085 16405 17115 16410
rect 17165 16430 17195 16435
rect 17165 16410 17170 16430
rect 17170 16410 17190 16430
rect 17190 16410 17195 16430
rect 17165 16405 17195 16410
rect 17245 16430 17275 16435
rect 17245 16410 17250 16430
rect 17250 16410 17270 16430
rect 17270 16410 17275 16430
rect 17245 16405 17275 16410
rect 17325 16430 17355 16435
rect 17325 16410 17330 16430
rect 17330 16410 17350 16430
rect 17350 16410 17355 16430
rect 17325 16405 17355 16410
rect 17405 16430 17435 16435
rect 17405 16410 17410 16430
rect 17410 16410 17430 16430
rect 17430 16410 17435 16430
rect 17405 16405 17435 16410
rect 17485 16430 17515 16435
rect 17485 16410 17490 16430
rect 17490 16410 17510 16430
rect 17510 16410 17515 16430
rect 17485 16405 17515 16410
rect 17565 16430 17595 16435
rect 17565 16410 17570 16430
rect 17570 16410 17590 16430
rect 17590 16410 17595 16430
rect 17565 16405 17595 16410
rect 17645 16430 17675 16435
rect 17645 16410 17650 16430
rect 17650 16410 17670 16430
rect 17670 16410 17675 16430
rect 17645 16405 17675 16410
rect 17725 16430 17755 16435
rect 17725 16410 17730 16430
rect 17730 16410 17750 16430
rect 17750 16410 17755 16430
rect 17725 16405 17755 16410
rect 17805 16430 17835 16435
rect 17805 16410 17810 16430
rect 17810 16410 17830 16430
rect 17830 16410 17835 16430
rect 17805 16405 17835 16410
rect 17885 16430 17915 16435
rect 17885 16410 17890 16430
rect 17890 16410 17910 16430
rect 17910 16410 17915 16430
rect 17885 16405 17915 16410
rect 17965 16430 17995 16435
rect 17965 16410 17970 16430
rect 17970 16410 17990 16430
rect 17990 16410 17995 16430
rect 17965 16405 17995 16410
rect 18045 16430 18075 16435
rect 18045 16410 18050 16430
rect 18050 16410 18070 16430
rect 18070 16410 18075 16430
rect 18045 16405 18075 16410
rect 18125 16430 18155 16435
rect 18125 16410 18130 16430
rect 18130 16410 18150 16430
rect 18150 16410 18155 16430
rect 18125 16405 18155 16410
rect 18205 16430 18235 16435
rect 18205 16410 18210 16430
rect 18210 16410 18230 16430
rect 18230 16410 18235 16430
rect 18205 16405 18235 16410
rect 18285 16430 18315 16435
rect 18285 16410 18290 16430
rect 18290 16410 18310 16430
rect 18310 16410 18315 16430
rect 18285 16405 18315 16410
rect 18365 16430 18395 16435
rect 18365 16410 18370 16430
rect 18370 16410 18390 16430
rect 18390 16410 18395 16430
rect 18365 16405 18395 16410
rect 18445 16430 18475 16435
rect 18445 16410 18450 16430
rect 18450 16410 18470 16430
rect 18470 16410 18475 16430
rect 18445 16405 18475 16410
rect 18525 16430 18555 16435
rect 18525 16410 18530 16430
rect 18530 16410 18550 16430
rect 18550 16410 18555 16430
rect 18525 16405 18555 16410
rect 18605 16430 18635 16435
rect 18605 16410 18610 16430
rect 18610 16410 18630 16430
rect 18630 16410 18635 16430
rect 18605 16405 18635 16410
rect 18685 16430 18715 16435
rect 18685 16410 18690 16430
rect 18690 16410 18710 16430
rect 18710 16410 18715 16430
rect 18685 16405 18715 16410
rect 18765 16430 18795 16435
rect 18765 16410 18770 16430
rect 18770 16410 18790 16430
rect 18790 16410 18795 16430
rect 18765 16405 18795 16410
rect 18845 16430 18875 16435
rect 18845 16410 18850 16430
rect 18850 16410 18870 16430
rect 18870 16410 18875 16430
rect 18845 16405 18875 16410
rect 18925 16430 18955 16435
rect 18925 16410 18930 16430
rect 18930 16410 18950 16430
rect 18950 16410 18955 16430
rect 18925 16405 18955 16410
rect 19005 16430 19035 16435
rect 19005 16410 19010 16430
rect 19010 16410 19030 16430
rect 19030 16410 19035 16430
rect 19005 16405 19035 16410
rect 19085 16430 19115 16435
rect 19085 16410 19090 16430
rect 19090 16410 19110 16430
rect 19110 16410 19115 16430
rect 19085 16405 19115 16410
rect 19165 16430 19195 16435
rect 19165 16410 19170 16430
rect 19170 16410 19190 16430
rect 19190 16410 19195 16430
rect 19165 16405 19195 16410
rect 19245 16430 19275 16435
rect 19245 16410 19250 16430
rect 19250 16410 19270 16430
rect 19270 16410 19275 16430
rect 19245 16405 19275 16410
rect 19325 16430 19355 16435
rect 19325 16410 19330 16430
rect 19330 16410 19350 16430
rect 19350 16410 19355 16430
rect 19325 16405 19355 16410
rect 19405 16430 19435 16435
rect 19405 16410 19410 16430
rect 19410 16410 19430 16430
rect 19430 16410 19435 16430
rect 19405 16405 19435 16410
rect 19485 16430 19515 16435
rect 19485 16410 19490 16430
rect 19490 16410 19510 16430
rect 19510 16410 19515 16430
rect 19485 16405 19515 16410
rect 19565 16430 19595 16435
rect 19565 16410 19570 16430
rect 19570 16410 19590 16430
rect 19590 16410 19595 16430
rect 19565 16405 19595 16410
rect 19645 16430 19675 16435
rect 19645 16410 19650 16430
rect 19650 16410 19670 16430
rect 19670 16410 19675 16430
rect 19645 16405 19675 16410
rect 19725 16430 19755 16435
rect 19725 16410 19730 16430
rect 19730 16410 19750 16430
rect 19750 16410 19755 16430
rect 19725 16405 19755 16410
rect 19805 16430 19835 16435
rect 19805 16410 19810 16430
rect 19810 16410 19830 16430
rect 19830 16410 19835 16430
rect 19805 16405 19835 16410
rect 19885 16430 19915 16435
rect 19885 16410 19890 16430
rect 19890 16410 19910 16430
rect 19910 16410 19915 16430
rect 19885 16405 19915 16410
rect 19965 16430 19995 16435
rect 19965 16410 19970 16430
rect 19970 16410 19990 16430
rect 19990 16410 19995 16430
rect 19965 16405 19995 16410
rect 20045 16430 20075 16435
rect 20045 16410 20050 16430
rect 20050 16410 20070 16430
rect 20070 16410 20075 16430
rect 20045 16405 20075 16410
rect 20125 16430 20155 16435
rect 20125 16410 20130 16430
rect 20130 16410 20150 16430
rect 20150 16410 20155 16430
rect 20125 16405 20155 16410
rect 20205 16430 20235 16435
rect 20205 16410 20210 16430
rect 20210 16410 20230 16430
rect 20230 16410 20235 16430
rect 20205 16405 20235 16410
rect 20285 16430 20315 16435
rect 20285 16410 20290 16430
rect 20290 16410 20310 16430
rect 20310 16410 20315 16430
rect 20285 16405 20315 16410
rect 20365 16430 20395 16435
rect 20365 16410 20370 16430
rect 20370 16410 20390 16430
rect 20390 16410 20395 16430
rect 20365 16405 20395 16410
rect 20445 16430 20475 16435
rect 20445 16410 20450 16430
rect 20450 16410 20470 16430
rect 20470 16410 20475 16430
rect 20445 16405 20475 16410
rect 20525 16430 20555 16435
rect 20525 16410 20530 16430
rect 20530 16410 20550 16430
rect 20550 16410 20555 16430
rect 20525 16405 20555 16410
rect 20605 16430 20635 16435
rect 20605 16410 20610 16430
rect 20610 16410 20630 16430
rect 20630 16410 20635 16430
rect 20605 16405 20635 16410
rect 20685 16430 20715 16435
rect 20685 16410 20690 16430
rect 20690 16410 20710 16430
rect 20710 16410 20715 16430
rect 20685 16405 20715 16410
rect 20765 16430 20795 16435
rect 20765 16410 20770 16430
rect 20770 16410 20790 16430
rect 20790 16410 20795 16430
rect 20765 16405 20795 16410
rect 20845 16430 20875 16435
rect 20845 16410 20850 16430
rect 20850 16410 20870 16430
rect 20870 16410 20875 16430
rect 20845 16405 20875 16410
rect 20925 16430 20955 16435
rect 20925 16410 20930 16430
rect 20930 16410 20950 16430
rect 20950 16410 20955 16430
rect 20925 16405 20955 16410
rect 5 16270 35 16275
rect 5 16250 10 16270
rect 10 16250 30 16270
rect 30 16250 35 16270
rect 5 16245 35 16250
rect 85 16270 115 16275
rect 85 16250 90 16270
rect 90 16250 110 16270
rect 110 16250 115 16270
rect 85 16245 115 16250
rect 165 16270 195 16275
rect 165 16250 170 16270
rect 170 16250 190 16270
rect 190 16250 195 16270
rect 165 16245 195 16250
rect 245 16270 275 16275
rect 245 16250 250 16270
rect 250 16250 270 16270
rect 270 16250 275 16270
rect 245 16245 275 16250
rect 325 16270 355 16275
rect 325 16250 330 16270
rect 330 16250 350 16270
rect 350 16250 355 16270
rect 325 16245 355 16250
rect 405 16270 435 16275
rect 405 16250 410 16270
rect 410 16250 430 16270
rect 430 16250 435 16270
rect 405 16245 435 16250
rect 485 16270 515 16275
rect 485 16250 490 16270
rect 490 16250 510 16270
rect 510 16250 515 16270
rect 485 16245 515 16250
rect 565 16270 595 16275
rect 565 16250 570 16270
rect 570 16250 590 16270
rect 590 16250 595 16270
rect 565 16245 595 16250
rect 645 16270 675 16275
rect 645 16250 650 16270
rect 650 16250 670 16270
rect 670 16250 675 16270
rect 645 16245 675 16250
rect 725 16270 755 16275
rect 725 16250 730 16270
rect 730 16250 750 16270
rect 750 16250 755 16270
rect 725 16245 755 16250
rect 805 16270 835 16275
rect 805 16250 810 16270
rect 810 16250 830 16270
rect 830 16250 835 16270
rect 805 16245 835 16250
rect 885 16270 915 16275
rect 885 16250 890 16270
rect 890 16250 910 16270
rect 910 16250 915 16270
rect 885 16245 915 16250
rect 965 16270 995 16275
rect 965 16250 970 16270
rect 970 16250 990 16270
rect 990 16250 995 16270
rect 965 16245 995 16250
rect 1045 16270 1075 16275
rect 1045 16250 1050 16270
rect 1050 16250 1070 16270
rect 1070 16250 1075 16270
rect 1045 16245 1075 16250
rect 1125 16270 1155 16275
rect 1125 16250 1130 16270
rect 1130 16250 1150 16270
rect 1150 16250 1155 16270
rect 1125 16245 1155 16250
rect 1205 16270 1235 16275
rect 1205 16250 1210 16270
rect 1210 16250 1230 16270
rect 1230 16250 1235 16270
rect 1205 16245 1235 16250
rect 1285 16270 1315 16275
rect 1285 16250 1290 16270
rect 1290 16250 1310 16270
rect 1310 16250 1315 16270
rect 1285 16245 1315 16250
rect 1365 16270 1395 16275
rect 1365 16250 1370 16270
rect 1370 16250 1390 16270
rect 1390 16250 1395 16270
rect 1365 16245 1395 16250
rect 1445 16270 1475 16275
rect 1445 16250 1450 16270
rect 1450 16250 1470 16270
rect 1470 16250 1475 16270
rect 1445 16245 1475 16250
rect 1525 16270 1555 16275
rect 1525 16250 1530 16270
rect 1530 16250 1550 16270
rect 1550 16250 1555 16270
rect 1525 16245 1555 16250
rect 1605 16270 1635 16275
rect 1605 16250 1610 16270
rect 1610 16250 1630 16270
rect 1630 16250 1635 16270
rect 1605 16245 1635 16250
rect 1685 16270 1715 16275
rect 1685 16250 1690 16270
rect 1690 16250 1710 16270
rect 1710 16250 1715 16270
rect 1685 16245 1715 16250
rect 1765 16270 1795 16275
rect 1765 16250 1770 16270
rect 1770 16250 1790 16270
rect 1790 16250 1795 16270
rect 1765 16245 1795 16250
rect 1845 16270 1875 16275
rect 1845 16250 1850 16270
rect 1850 16250 1870 16270
rect 1870 16250 1875 16270
rect 1845 16245 1875 16250
rect 1925 16270 1955 16275
rect 1925 16250 1930 16270
rect 1930 16250 1950 16270
rect 1950 16250 1955 16270
rect 1925 16245 1955 16250
rect 2005 16270 2035 16275
rect 2005 16250 2010 16270
rect 2010 16250 2030 16270
rect 2030 16250 2035 16270
rect 2005 16245 2035 16250
rect 2085 16270 2115 16275
rect 2085 16250 2090 16270
rect 2090 16250 2110 16270
rect 2110 16250 2115 16270
rect 2085 16245 2115 16250
rect 2165 16270 2195 16275
rect 2165 16250 2170 16270
rect 2170 16250 2190 16270
rect 2190 16250 2195 16270
rect 2165 16245 2195 16250
rect 2245 16270 2275 16275
rect 2245 16250 2250 16270
rect 2250 16250 2270 16270
rect 2270 16250 2275 16270
rect 2245 16245 2275 16250
rect 2325 16270 2355 16275
rect 2325 16250 2330 16270
rect 2330 16250 2350 16270
rect 2350 16250 2355 16270
rect 2325 16245 2355 16250
rect 2405 16270 2435 16275
rect 2405 16250 2410 16270
rect 2410 16250 2430 16270
rect 2430 16250 2435 16270
rect 2405 16245 2435 16250
rect 2485 16270 2515 16275
rect 2485 16250 2490 16270
rect 2490 16250 2510 16270
rect 2510 16250 2515 16270
rect 2485 16245 2515 16250
rect 2565 16270 2595 16275
rect 2565 16250 2570 16270
rect 2570 16250 2590 16270
rect 2590 16250 2595 16270
rect 2565 16245 2595 16250
rect 2645 16270 2675 16275
rect 2645 16250 2650 16270
rect 2650 16250 2670 16270
rect 2670 16250 2675 16270
rect 2645 16245 2675 16250
rect 2725 16270 2755 16275
rect 2725 16250 2730 16270
rect 2730 16250 2750 16270
rect 2750 16250 2755 16270
rect 2725 16245 2755 16250
rect 2805 16270 2835 16275
rect 2805 16250 2810 16270
rect 2810 16250 2830 16270
rect 2830 16250 2835 16270
rect 2805 16245 2835 16250
rect 2885 16270 2915 16275
rect 2885 16250 2890 16270
rect 2890 16250 2910 16270
rect 2910 16250 2915 16270
rect 2885 16245 2915 16250
rect 2965 16270 2995 16275
rect 2965 16250 2970 16270
rect 2970 16250 2990 16270
rect 2990 16250 2995 16270
rect 2965 16245 2995 16250
rect 3045 16270 3075 16275
rect 3045 16250 3050 16270
rect 3050 16250 3070 16270
rect 3070 16250 3075 16270
rect 3045 16245 3075 16250
rect 3125 16270 3155 16275
rect 3125 16250 3130 16270
rect 3130 16250 3150 16270
rect 3150 16250 3155 16270
rect 3125 16245 3155 16250
rect 3205 16270 3235 16275
rect 3205 16250 3210 16270
rect 3210 16250 3230 16270
rect 3230 16250 3235 16270
rect 3205 16245 3235 16250
rect 3285 16270 3315 16275
rect 3285 16250 3290 16270
rect 3290 16250 3310 16270
rect 3310 16250 3315 16270
rect 3285 16245 3315 16250
rect 3365 16270 3395 16275
rect 3365 16250 3370 16270
rect 3370 16250 3390 16270
rect 3390 16250 3395 16270
rect 3365 16245 3395 16250
rect 3445 16270 3475 16275
rect 3445 16250 3450 16270
rect 3450 16250 3470 16270
rect 3470 16250 3475 16270
rect 3445 16245 3475 16250
rect 3525 16270 3555 16275
rect 3525 16250 3530 16270
rect 3530 16250 3550 16270
rect 3550 16250 3555 16270
rect 3525 16245 3555 16250
rect 3605 16270 3635 16275
rect 3605 16250 3610 16270
rect 3610 16250 3630 16270
rect 3630 16250 3635 16270
rect 3605 16245 3635 16250
rect 3685 16270 3715 16275
rect 3685 16250 3690 16270
rect 3690 16250 3710 16270
rect 3710 16250 3715 16270
rect 3685 16245 3715 16250
rect 3765 16270 3795 16275
rect 3765 16250 3770 16270
rect 3770 16250 3790 16270
rect 3790 16250 3795 16270
rect 3765 16245 3795 16250
rect 3845 16270 3875 16275
rect 3845 16250 3850 16270
rect 3850 16250 3870 16270
rect 3870 16250 3875 16270
rect 3845 16245 3875 16250
rect 3925 16270 3955 16275
rect 3925 16250 3930 16270
rect 3930 16250 3950 16270
rect 3950 16250 3955 16270
rect 3925 16245 3955 16250
rect 4005 16270 4035 16275
rect 4005 16250 4010 16270
rect 4010 16250 4030 16270
rect 4030 16250 4035 16270
rect 4005 16245 4035 16250
rect 4085 16270 4115 16275
rect 4085 16250 4090 16270
rect 4090 16250 4110 16270
rect 4110 16250 4115 16270
rect 4085 16245 4115 16250
rect 4165 16270 4195 16275
rect 4165 16250 4170 16270
rect 4170 16250 4190 16270
rect 4190 16250 4195 16270
rect 4165 16245 4195 16250
rect 6245 16270 6275 16275
rect 6245 16250 6250 16270
rect 6250 16250 6270 16270
rect 6270 16250 6275 16270
rect 6245 16245 6275 16250
rect 6325 16270 6355 16275
rect 6325 16250 6330 16270
rect 6330 16250 6350 16270
rect 6350 16250 6355 16270
rect 6325 16245 6355 16250
rect 6405 16270 6435 16275
rect 6405 16250 6410 16270
rect 6410 16250 6430 16270
rect 6430 16250 6435 16270
rect 6405 16245 6435 16250
rect 6485 16270 6515 16275
rect 6485 16250 6490 16270
rect 6490 16250 6510 16270
rect 6510 16250 6515 16270
rect 6485 16245 6515 16250
rect 6565 16270 6595 16275
rect 6565 16250 6570 16270
rect 6570 16250 6590 16270
rect 6590 16250 6595 16270
rect 6565 16245 6595 16250
rect 6645 16270 6675 16275
rect 6645 16250 6650 16270
rect 6650 16250 6670 16270
rect 6670 16250 6675 16270
rect 6645 16245 6675 16250
rect 6725 16270 6755 16275
rect 6725 16250 6730 16270
rect 6730 16250 6750 16270
rect 6750 16250 6755 16270
rect 6725 16245 6755 16250
rect 6805 16270 6835 16275
rect 6805 16250 6810 16270
rect 6810 16250 6830 16270
rect 6830 16250 6835 16270
rect 6805 16245 6835 16250
rect 6885 16270 6915 16275
rect 6885 16250 6890 16270
rect 6890 16250 6910 16270
rect 6910 16250 6915 16270
rect 6885 16245 6915 16250
rect 6965 16270 6995 16275
rect 6965 16250 6970 16270
rect 6970 16250 6990 16270
rect 6990 16250 6995 16270
rect 6965 16245 6995 16250
rect 7045 16270 7075 16275
rect 7045 16250 7050 16270
rect 7050 16250 7070 16270
rect 7070 16250 7075 16270
rect 7045 16245 7075 16250
rect 7125 16270 7155 16275
rect 7125 16250 7130 16270
rect 7130 16250 7150 16270
rect 7150 16250 7155 16270
rect 7125 16245 7155 16250
rect 7205 16270 7235 16275
rect 7205 16250 7210 16270
rect 7210 16250 7230 16270
rect 7230 16250 7235 16270
rect 7205 16245 7235 16250
rect 7285 16270 7315 16275
rect 7285 16250 7290 16270
rect 7290 16250 7310 16270
rect 7310 16250 7315 16270
rect 7285 16245 7315 16250
rect 7365 16270 7395 16275
rect 7365 16250 7370 16270
rect 7370 16250 7390 16270
rect 7390 16250 7395 16270
rect 7365 16245 7395 16250
rect 7445 16270 7475 16275
rect 7445 16250 7450 16270
rect 7450 16250 7470 16270
rect 7470 16250 7475 16270
rect 7445 16245 7475 16250
rect 7525 16270 7555 16275
rect 7525 16250 7530 16270
rect 7530 16250 7550 16270
rect 7550 16250 7555 16270
rect 7525 16245 7555 16250
rect 7605 16270 7635 16275
rect 7605 16250 7610 16270
rect 7610 16250 7630 16270
rect 7630 16250 7635 16270
rect 7605 16245 7635 16250
rect 7685 16270 7715 16275
rect 7685 16250 7690 16270
rect 7690 16250 7710 16270
rect 7710 16250 7715 16270
rect 7685 16245 7715 16250
rect 7765 16270 7795 16275
rect 7765 16250 7770 16270
rect 7770 16250 7790 16270
rect 7790 16250 7795 16270
rect 7765 16245 7795 16250
rect 7845 16270 7875 16275
rect 7845 16250 7850 16270
rect 7850 16250 7870 16270
rect 7870 16250 7875 16270
rect 7845 16245 7875 16250
rect 7925 16270 7955 16275
rect 7925 16250 7930 16270
rect 7930 16250 7950 16270
rect 7950 16250 7955 16270
rect 7925 16245 7955 16250
rect 8005 16270 8035 16275
rect 8005 16250 8010 16270
rect 8010 16250 8030 16270
rect 8030 16250 8035 16270
rect 8005 16245 8035 16250
rect 8085 16270 8115 16275
rect 8085 16250 8090 16270
rect 8090 16250 8110 16270
rect 8110 16250 8115 16270
rect 8085 16245 8115 16250
rect 8165 16270 8195 16275
rect 8165 16250 8170 16270
rect 8170 16250 8190 16270
rect 8190 16250 8195 16270
rect 8165 16245 8195 16250
rect 8245 16270 8275 16275
rect 8245 16250 8250 16270
rect 8250 16250 8270 16270
rect 8270 16250 8275 16270
rect 8245 16245 8275 16250
rect 8325 16270 8355 16275
rect 8325 16250 8330 16270
rect 8330 16250 8350 16270
rect 8350 16250 8355 16270
rect 8325 16245 8355 16250
rect 8405 16270 8435 16275
rect 8405 16250 8410 16270
rect 8410 16250 8430 16270
rect 8430 16250 8435 16270
rect 8405 16245 8435 16250
rect 8485 16270 8515 16275
rect 8485 16250 8490 16270
rect 8490 16250 8510 16270
rect 8510 16250 8515 16270
rect 8485 16245 8515 16250
rect 8565 16270 8595 16275
rect 8565 16250 8570 16270
rect 8570 16250 8590 16270
rect 8590 16250 8595 16270
rect 8565 16245 8595 16250
rect 8645 16270 8675 16275
rect 8645 16250 8650 16270
rect 8650 16250 8670 16270
rect 8670 16250 8675 16270
rect 8645 16245 8675 16250
rect 8725 16270 8755 16275
rect 8725 16250 8730 16270
rect 8730 16250 8750 16270
rect 8750 16250 8755 16270
rect 8725 16245 8755 16250
rect 8805 16270 8835 16275
rect 8805 16250 8810 16270
rect 8810 16250 8830 16270
rect 8830 16250 8835 16270
rect 8805 16245 8835 16250
rect 8885 16270 8915 16275
rect 8885 16250 8890 16270
rect 8890 16250 8910 16270
rect 8910 16250 8915 16270
rect 8885 16245 8915 16250
rect 8965 16270 8995 16275
rect 8965 16250 8970 16270
rect 8970 16250 8990 16270
rect 8990 16250 8995 16270
rect 8965 16245 8995 16250
rect 9045 16270 9075 16275
rect 9045 16250 9050 16270
rect 9050 16250 9070 16270
rect 9070 16250 9075 16270
rect 9045 16245 9075 16250
rect 9125 16270 9155 16275
rect 9125 16250 9130 16270
rect 9130 16250 9150 16270
rect 9150 16250 9155 16270
rect 9125 16245 9155 16250
rect 9205 16270 9235 16275
rect 9205 16250 9210 16270
rect 9210 16250 9230 16270
rect 9230 16250 9235 16270
rect 9205 16245 9235 16250
rect 9285 16270 9315 16275
rect 9285 16250 9290 16270
rect 9290 16250 9310 16270
rect 9310 16250 9315 16270
rect 9285 16245 9315 16250
rect 9365 16270 9395 16275
rect 9365 16250 9370 16270
rect 9370 16250 9390 16270
rect 9390 16250 9395 16270
rect 9365 16245 9395 16250
rect 9445 16270 9475 16275
rect 9445 16250 9450 16270
rect 9450 16250 9470 16270
rect 9470 16250 9475 16270
rect 9445 16245 9475 16250
rect 11565 16270 11595 16275
rect 11565 16250 11570 16270
rect 11570 16250 11590 16270
rect 11590 16250 11595 16270
rect 11565 16245 11595 16250
rect 11645 16270 11675 16275
rect 11645 16250 11650 16270
rect 11650 16250 11670 16270
rect 11670 16250 11675 16270
rect 11645 16245 11675 16250
rect 11725 16270 11755 16275
rect 11725 16250 11730 16270
rect 11730 16250 11750 16270
rect 11750 16250 11755 16270
rect 11725 16245 11755 16250
rect 11805 16270 11835 16275
rect 11805 16250 11810 16270
rect 11810 16250 11830 16270
rect 11830 16250 11835 16270
rect 11805 16245 11835 16250
rect 11885 16270 11915 16275
rect 11885 16250 11890 16270
rect 11890 16250 11910 16270
rect 11910 16250 11915 16270
rect 11885 16245 11915 16250
rect 11965 16270 11995 16275
rect 11965 16250 11970 16270
rect 11970 16250 11990 16270
rect 11990 16250 11995 16270
rect 11965 16245 11995 16250
rect 12045 16270 12075 16275
rect 12045 16250 12050 16270
rect 12050 16250 12070 16270
rect 12070 16250 12075 16270
rect 12045 16245 12075 16250
rect 12125 16270 12155 16275
rect 12125 16250 12130 16270
rect 12130 16250 12150 16270
rect 12150 16250 12155 16270
rect 12125 16245 12155 16250
rect 12205 16270 12235 16275
rect 12205 16250 12210 16270
rect 12210 16250 12230 16270
rect 12230 16250 12235 16270
rect 12205 16245 12235 16250
rect 12285 16270 12315 16275
rect 12285 16250 12290 16270
rect 12290 16250 12310 16270
rect 12310 16250 12315 16270
rect 12285 16245 12315 16250
rect 12365 16270 12395 16275
rect 12365 16250 12370 16270
rect 12370 16250 12390 16270
rect 12390 16250 12395 16270
rect 12365 16245 12395 16250
rect 12445 16270 12475 16275
rect 12445 16250 12450 16270
rect 12450 16250 12470 16270
rect 12470 16250 12475 16270
rect 12445 16245 12475 16250
rect 12525 16270 12555 16275
rect 12525 16250 12530 16270
rect 12530 16250 12550 16270
rect 12550 16250 12555 16270
rect 12525 16245 12555 16250
rect 12605 16270 12635 16275
rect 12605 16250 12610 16270
rect 12610 16250 12630 16270
rect 12630 16250 12635 16270
rect 12605 16245 12635 16250
rect 12685 16270 12715 16275
rect 12685 16250 12690 16270
rect 12690 16250 12710 16270
rect 12710 16250 12715 16270
rect 12685 16245 12715 16250
rect 12765 16270 12795 16275
rect 12765 16250 12770 16270
rect 12770 16250 12790 16270
rect 12790 16250 12795 16270
rect 12765 16245 12795 16250
rect 12845 16270 12875 16275
rect 12845 16250 12850 16270
rect 12850 16250 12870 16270
rect 12870 16250 12875 16270
rect 12845 16245 12875 16250
rect 12925 16270 12955 16275
rect 12925 16250 12930 16270
rect 12930 16250 12950 16270
rect 12950 16250 12955 16270
rect 12925 16245 12955 16250
rect 13005 16270 13035 16275
rect 13005 16250 13010 16270
rect 13010 16250 13030 16270
rect 13030 16250 13035 16270
rect 13005 16245 13035 16250
rect 13085 16270 13115 16275
rect 13085 16250 13090 16270
rect 13090 16250 13110 16270
rect 13110 16250 13115 16270
rect 13085 16245 13115 16250
rect 13165 16270 13195 16275
rect 13165 16250 13170 16270
rect 13170 16250 13190 16270
rect 13190 16250 13195 16270
rect 13165 16245 13195 16250
rect 13245 16270 13275 16275
rect 13245 16250 13250 16270
rect 13250 16250 13270 16270
rect 13270 16250 13275 16270
rect 13245 16245 13275 16250
rect 13325 16270 13355 16275
rect 13325 16250 13330 16270
rect 13330 16250 13350 16270
rect 13350 16250 13355 16270
rect 13325 16245 13355 16250
rect 13405 16270 13435 16275
rect 13405 16250 13410 16270
rect 13410 16250 13430 16270
rect 13430 16250 13435 16270
rect 13405 16245 13435 16250
rect 13485 16270 13515 16275
rect 13485 16250 13490 16270
rect 13490 16250 13510 16270
rect 13510 16250 13515 16270
rect 13485 16245 13515 16250
rect 13565 16270 13595 16275
rect 13565 16250 13570 16270
rect 13570 16250 13590 16270
rect 13590 16250 13595 16270
rect 13565 16245 13595 16250
rect 13645 16270 13675 16275
rect 13645 16250 13650 16270
rect 13650 16250 13670 16270
rect 13670 16250 13675 16270
rect 13645 16245 13675 16250
rect 13725 16270 13755 16275
rect 13725 16250 13730 16270
rect 13730 16250 13750 16270
rect 13750 16250 13755 16270
rect 13725 16245 13755 16250
rect 13805 16270 13835 16275
rect 13805 16250 13810 16270
rect 13810 16250 13830 16270
rect 13830 16250 13835 16270
rect 13805 16245 13835 16250
rect 13885 16270 13915 16275
rect 13885 16250 13890 16270
rect 13890 16250 13910 16270
rect 13910 16250 13915 16270
rect 13885 16245 13915 16250
rect 13965 16270 13995 16275
rect 13965 16250 13970 16270
rect 13970 16250 13990 16270
rect 13990 16250 13995 16270
rect 13965 16245 13995 16250
rect 14045 16270 14075 16275
rect 14045 16250 14050 16270
rect 14050 16250 14070 16270
rect 14070 16250 14075 16270
rect 14045 16245 14075 16250
rect 14125 16270 14155 16275
rect 14125 16250 14130 16270
rect 14130 16250 14150 16270
rect 14150 16250 14155 16270
rect 14125 16245 14155 16250
rect 14205 16270 14235 16275
rect 14205 16250 14210 16270
rect 14210 16250 14230 16270
rect 14230 16250 14235 16270
rect 14205 16245 14235 16250
rect 14285 16270 14315 16275
rect 14285 16250 14290 16270
rect 14290 16250 14310 16270
rect 14310 16250 14315 16270
rect 14285 16245 14315 16250
rect 14365 16270 14395 16275
rect 14365 16250 14370 16270
rect 14370 16250 14390 16270
rect 14390 16250 14395 16270
rect 14365 16245 14395 16250
rect 14445 16270 14475 16275
rect 14445 16250 14450 16270
rect 14450 16250 14470 16270
rect 14470 16250 14475 16270
rect 14445 16245 14475 16250
rect 14525 16270 14555 16275
rect 14525 16250 14530 16270
rect 14530 16250 14550 16270
rect 14550 16250 14555 16270
rect 14525 16245 14555 16250
rect 14605 16270 14635 16275
rect 14605 16250 14610 16270
rect 14610 16250 14630 16270
rect 14630 16250 14635 16270
rect 14605 16245 14635 16250
rect 14685 16270 14715 16275
rect 14685 16250 14690 16270
rect 14690 16250 14710 16270
rect 14710 16250 14715 16270
rect 14685 16245 14715 16250
rect 16765 16270 16795 16275
rect 16765 16250 16770 16270
rect 16770 16250 16790 16270
rect 16790 16250 16795 16270
rect 16765 16245 16795 16250
rect 16845 16270 16875 16275
rect 16845 16250 16850 16270
rect 16850 16250 16870 16270
rect 16870 16250 16875 16270
rect 16845 16245 16875 16250
rect 16925 16270 16955 16275
rect 16925 16250 16930 16270
rect 16930 16250 16950 16270
rect 16950 16250 16955 16270
rect 16925 16245 16955 16250
rect 17005 16270 17035 16275
rect 17005 16250 17010 16270
rect 17010 16250 17030 16270
rect 17030 16250 17035 16270
rect 17005 16245 17035 16250
rect 17085 16270 17115 16275
rect 17085 16250 17090 16270
rect 17090 16250 17110 16270
rect 17110 16250 17115 16270
rect 17085 16245 17115 16250
rect 17165 16270 17195 16275
rect 17165 16250 17170 16270
rect 17170 16250 17190 16270
rect 17190 16250 17195 16270
rect 17165 16245 17195 16250
rect 17245 16270 17275 16275
rect 17245 16250 17250 16270
rect 17250 16250 17270 16270
rect 17270 16250 17275 16270
rect 17245 16245 17275 16250
rect 17325 16270 17355 16275
rect 17325 16250 17330 16270
rect 17330 16250 17350 16270
rect 17350 16250 17355 16270
rect 17325 16245 17355 16250
rect 17405 16270 17435 16275
rect 17405 16250 17410 16270
rect 17410 16250 17430 16270
rect 17430 16250 17435 16270
rect 17405 16245 17435 16250
rect 17485 16270 17515 16275
rect 17485 16250 17490 16270
rect 17490 16250 17510 16270
rect 17510 16250 17515 16270
rect 17485 16245 17515 16250
rect 17565 16270 17595 16275
rect 17565 16250 17570 16270
rect 17570 16250 17590 16270
rect 17590 16250 17595 16270
rect 17565 16245 17595 16250
rect 17645 16270 17675 16275
rect 17645 16250 17650 16270
rect 17650 16250 17670 16270
rect 17670 16250 17675 16270
rect 17645 16245 17675 16250
rect 17725 16270 17755 16275
rect 17725 16250 17730 16270
rect 17730 16250 17750 16270
rect 17750 16250 17755 16270
rect 17725 16245 17755 16250
rect 17805 16270 17835 16275
rect 17805 16250 17810 16270
rect 17810 16250 17830 16270
rect 17830 16250 17835 16270
rect 17805 16245 17835 16250
rect 17885 16270 17915 16275
rect 17885 16250 17890 16270
rect 17890 16250 17910 16270
rect 17910 16250 17915 16270
rect 17885 16245 17915 16250
rect 17965 16270 17995 16275
rect 17965 16250 17970 16270
rect 17970 16250 17990 16270
rect 17990 16250 17995 16270
rect 17965 16245 17995 16250
rect 18045 16270 18075 16275
rect 18045 16250 18050 16270
rect 18050 16250 18070 16270
rect 18070 16250 18075 16270
rect 18045 16245 18075 16250
rect 18125 16270 18155 16275
rect 18125 16250 18130 16270
rect 18130 16250 18150 16270
rect 18150 16250 18155 16270
rect 18125 16245 18155 16250
rect 18205 16270 18235 16275
rect 18205 16250 18210 16270
rect 18210 16250 18230 16270
rect 18230 16250 18235 16270
rect 18205 16245 18235 16250
rect 18285 16270 18315 16275
rect 18285 16250 18290 16270
rect 18290 16250 18310 16270
rect 18310 16250 18315 16270
rect 18285 16245 18315 16250
rect 18365 16270 18395 16275
rect 18365 16250 18370 16270
rect 18370 16250 18390 16270
rect 18390 16250 18395 16270
rect 18365 16245 18395 16250
rect 18445 16270 18475 16275
rect 18445 16250 18450 16270
rect 18450 16250 18470 16270
rect 18470 16250 18475 16270
rect 18445 16245 18475 16250
rect 18525 16270 18555 16275
rect 18525 16250 18530 16270
rect 18530 16250 18550 16270
rect 18550 16250 18555 16270
rect 18525 16245 18555 16250
rect 18605 16270 18635 16275
rect 18605 16250 18610 16270
rect 18610 16250 18630 16270
rect 18630 16250 18635 16270
rect 18605 16245 18635 16250
rect 18685 16270 18715 16275
rect 18685 16250 18690 16270
rect 18690 16250 18710 16270
rect 18710 16250 18715 16270
rect 18685 16245 18715 16250
rect 18765 16270 18795 16275
rect 18765 16250 18770 16270
rect 18770 16250 18790 16270
rect 18790 16250 18795 16270
rect 18765 16245 18795 16250
rect 18845 16270 18875 16275
rect 18845 16250 18850 16270
rect 18850 16250 18870 16270
rect 18870 16250 18875 16270
rect 18845 16245 18875 16250
rect 18925 16270 18955 16275
rect 18925 16250 18930 16270
rect 18930 16250 18950 16270
rect 18950 16250 18955 16270
rect 18925 16245 18955 16250
rect 19005 16270 19035 16275
rect 19005 16250 19010 16270
rect 19010 16250 19030 16270
rect 19030 16250 19035 16270
rect 19005 16245 19035 16250
rect 19085 16270 19115 16275
rect 19085 16250 19090 16270
rect 19090 16250 19110 16270
rect 19110 16250 19115 16270
rect 19085 16245 19115 16250
rect 19165 16270 19195 16275
rect 19165 16250 19170 16270
rect 19170 16250 19190 16270
rect 19190 16250 19195 16270
rect 19165 16245 19195 16250
rect 19245 16270 19275 16275
rect 19245 16250 19250 16270
rect 19250 16250 19270 16270
rect 19270 16250 19275 16270
rect 19245 16245 19275 16250
rect 19325 16270 19355 16275
rect 19325 16250 19330 16270
rect 19330 16250 19350 16270
rect 19350 16250 19355 16270
rect 19325 16245 19355 16250
rect 19405 16270 19435 16275
rect 19405 16250 19410 16270
rect 19410 16250 19430 16270
rect 19430 16250 19435 16270
rect 19405 16245 19435 16250
rect 19485 16270 19515 16275
rect 19485 16250 19490 16270
rect 19490 16250 19510 16270
rect 19510 16250 19515 16270
rect 19485 16245 19515 16250
rect 19565 16270 19595 16275
rect 19565 16250 19570 16270
rect 19570 16250 19590 16270
rect 19590 16250 19595 16270
rect 19565 16245 19595 16250
rect 19645 16270 19675 16275
rect 19645 16250 19650 16270
rect 19650 16250 19670 16270
rect 19670 16250 19675 16270
rect 19645 16245 19675 16250
rect 19725 16270 19755 16275
rect 19725 16250 19730 16270
rect 19730 16250 19750 16270
rect 19750 16250 19755 16270
rect 19725 16245 19755 16250
rect 19805 16270 19835 16275
rect 19805 16250 19810 16270
rect 19810 16250 19830 16270
rect 19830 16250 19835 16270
rect 19805 16245 19835 16250
rect 19885 16270 19915 16275
rect 19885 16250 19890 16270
rect 19890 16250 19910 16270
rect 19910 16250 19915 16270
rect 19885 16245 19915 16250
rect 19965 16270 19995 16275
rect 19965 16250 19970 16270
rect 19970 16250 19990 16270
rect 19990 16250 19995 16270
rect 19965 16245 19995 16250
rect 20045 16270 20075 16275
rect 20045 16250 20050 16270
rect 20050 16250 20070 16270
rect 20070 16250 20075 16270
rect 20045 16245 20075 16250
rect 20125 16270 20155 16275
rect 20125 16250 20130 16270
rect 20130 16250 20150 16270
rect 20150 16250 20155 16270
rect 20125 16245 20155 16250
rect 20205 16270 20235 16275
rect 20205 16250 20210 16270
rect 20210 16250 20230 16270
rect 20230 16250 20235 16270
rect 20205 16245 20235 16250
rect 20285 16270 20315 16275
rect 20285 16250 20290 16270
rect 20290 16250 20310 16270
rect 20310 16250 20315 16270
rect 20285 16245 20315 16250
rect 20365 16270 20395 16275
rect 20365 16250 20370 16270
rect 20370 16250 20390 16270
rect 20390 16250 20395 16270
rect 20365 16245 20395 16250
rect 20445 16270 20475 16275
rect 20445 16250 20450 16270
rect 20450 16250 20470 16270
rect 20470 16250 20475 16270
rect 20445 16245 20475 16250
rect 20525 16270 20555 16275
rect 20525 16250 20530 16270
rect 20530 16250 20550 16270
rect 20550 16250 20555 16270
rect 20525 16245 20555 16250
rect 20605 16270 20635 16275
rect 20605 16250 20610 16270
rect 20610 16250 20630 16270
rect 20630 16250 20635 16270
rect 20605 16245 20635 16250
rect 20685 16270 20715 16275
rect 20685 16250 20690 16270
rect 20690 16250 20710 16270
rect 20710 16250 20715 16270
rect 20685 16245 20715 16250
rect 20765 16270 20795 16275
rect 20765 16250 20770 16270
rect 20770 16250 20790 16270
rect 20790 16250 20795 16270
rect 20765 16245 20795 16250
rect 20845 16270 20875 16275
rect 20845 16250 20850 16270
rect 20850 16250 20870 16270
rect 20870 16250 20875 16270
rect 20845 16245 20875 16250
rect 20925 16270 20955 16275
rect 20925 16250 20930 16270
rect 20930 16250 20950 16270
rect 20950 16250 20955 16270
rect 20925 16245 20955 16250
rect 5 16190 35 16195
rect 5 16170 10 16190
rect 10 16170 30 16190
rect 30 16170 35 16190
rect 5 16165 35 16170
rect 85 16190 115 16195
rect 85 16170 90 16190
rect 90 16170 110 16190
rect 110 16170 115 16190
rect 85 16165 115 16170
rect 165 16190 195 16195
rect 165 16170 170 16190
rect 170 16170 190 16190
rect 190 16170 195 16190
rect 165 16165 195 16170
rect 245 16190 275 16195
rect 245 16170 250 16190
rect 250 16170 270 16190
rect 270 16170 275 16190
rect 245 16165 275 16170
rect 325 16190 355 16195
rect 325 16170 330 16190
rect 330 16170 350 16190
rect 350 16170 355 16190
rect 325 16165 355 16170
rect 405 16190 435 16195
rect 405 16170 410 16190
rect 410 16170 430 16190
rect 430 16170 435 16190
rect 405 16165 435 16170
rect 485 16190 515 16195
rect 485 16170 490 16190
rect 490 16170 510 16190
rect 510 16170 515 16190
rect 485 16165 515 16170
rect 565 16190 595 16195
rect 565 16170 570 16190
rect 570 16170 590 16190
rect 590 16170 595 16190
rect 565 16165 595 16170
rect 645 16190 675 16195
rect 645 16170 650 16190
rect 650 16170 670 16190
rect 670 16170 675 16190
rect 645 16165 675 16170
rect 725 16190 755 16195
rect 725 16170 730 16190
rect 730 16170 750 16190
rect 750 16170 755 16190
rect 725 16165 755 16170
rect 805 16190 835 16195
rect 805 16170 810 16190
rect 810 16170 830 16190
rect 830 16170 835 16190
rect 805 16165 835 16170
rect 885 16190 915 16195
rect 885 16170 890 16190
rect 890 16170 910 16190
rect 910 16170 915 16190
rect 885 16165 915 16170
rect 965 16190 995 16195
rect 965 16170 970 16190
rect 970 16170 990 16190
rect 990 16170 995 16190
rect 965 16165 995 16170
rect 1045 16190 1075 16195
rect 1045 16170 1050 16190
rect 1050 16170 1070 16190
rect 1070 16170 1075 16190
rect 1045 16165 1075 16170
rect 1125 16190 1155 16195
rect 1125 16170 1130 16190
rect 1130 16170 1150 16190
rect 1150 16170 1155 16190
rect 1125 16165 1155 16170
rect 1205 16190 1235 16195
rect 1205 16170 1210 16190
rect 1210 16170 1230 16190
rect 1230 16170 1235 16190
rect 1205 16165 1235 16170
rect 1285 16190 1315 16195
rect 1285 16170 1290 16190
rect 1290 16170 1310 16190
rect 1310 16170 1315 16190
rect 1285 16165 1315 16170
rect 1365 16190 1395 16195
rect 1365 16170 1370 16190
rect 1370 16170 1390 16190
rect 1390 16170 1395 16190
rect 1365 16165 1395 16170
rect 1445 16190 1475 16195
rect 1445 16170 1450 16190
rect 1450 16170 1470 16190
rect 1470 16170 1475 16190
rect 1445 16165 1475 16170
rect 1525 16190 1555 16195
rect 1525 16170 1530 16190
rect 1530 16170 1550 16190
rect 1550 16170 1555 16190
rect 1525 16165 1555 16170
rect 1605 16190 1635 16195
rect 1605 16170 1610 16190
rect 1610 16170 1630 16190
rect 1630 16170 1635 16190
rect 1605 16165 1635 16170
rect 1685 16190 1715 16195
rect 1685 16170 1690 16190
rect 1690 16170 1710 16190
rect 1710 16170 1715 16190
rect 1685 16165 1715 16170
rect 1765 16190 1795 16195
rect 1765 16170 1770 16190
rect 1770 16170 1790 16190
rect 1790 16170 1795 16190
rect 1765 16165 1795 16170
rect 1845 16190 1875 16195
rect 1845 16170 1850 16190
rect 1850 16170 1870 16190
rect 1870 16170 1875 16190
rect 1845 16165 1875 16170
rect 1925 16190 1955 16195
rect 1925 16170 1930 16190
rect 1930 16170 1950 16190
rect 1950 16170 1955 16190
rect 1925 16165 1955 16170
rect 2005 16190 2035 16195
rect 2005 16170 2010 16190
rect 2010 16170 2030 16190
rect 2030 16170 2035 16190
rect 2005 16165 2035 16170
rect 2085 16190 2115 16195
rect 2085 16170 2090 16190
rect 2090 16170 2110 16190
rect 2110 16170 2115 16190
rect 2085 16165 2115 16170
rect 2165 16190 2195 16195
rect 2165 16170 2170 16190
rect 2170 16170 2190 16190
rect 2190 16170 2195 16190
rect 2165 16165 2195 16170
rect 2245 16190 2275 16195
rect 2245 16170 2250 16190
rect 2250 16170 2270 16190
rect 2270 16170 2275 16190
rect 2245 16165 2275 16170
rect 2325 16190 2355 16195
rect 2325 16170 2330 16190
rect 2330 16170 2350 16190
rect 2350 16170 2355 16190
rect 2325 16165 2355 16170
rect 2405 16190 2435 16195
rect 2405 16170 2410 16190
rect 2410 16170 2430 16190
rect 2430 16170 2435 16190
rect 2405 16165 2435 16170
rect 2485 16190 2515 16195
rect 2485 16170 2490 16190
rect 2490 16170 2510 16190
rect 2510 16170 2515 16190
rect 2485 16165 2515 16170
rect 2565 16190 2595 16195
rect 2565 16170 2570 16190
rect 2570 16170 2590 16190
rect 2590 16170 2595 16190
rect 2565 16165 2595 16170
rect 2645 16190 2675 16195
rect 2645 16170 2650 16190
rect 2650 16170 2670 16190
rect 2670 16170 2675 16190
rect 2645 16165 2675 16170
rect 2725 16190 2755 16195
rect 2725 16170 2730 16190
rect 2730 16170 2750 16190
rect 2750 16170 2755 16190
rect 2725 16165 2755 16170
rect 2805 16190 2835 16195
rect 2805 16170 2810 16190
rect 2810 16170 2830 16190
rect 2830 16170 2835 16190
rect 2805 16165 2835 16170
rect 2885 16190 2915 16195
rect 2885 16170 2890 16190
rect 2890 16170 2910 16190
rect 2910 16170 2915 16190
rect 2885 16165 2915 16170
rect 2965 16190 2995 16195
rect 2965 16170 2970 16190
rect 2970 16170 2990 16190
rect 2990 16170 2995 16190
rect 2965 16165 2995 16170
rect 3045 16190 3075 16195
rect 3045 16170 3050 16190
rect 3050 16170 3070 16190
rect 3070 16170 3075 16190
rect 3045 16165 3075 16170
rect 3125 16190 3155 16195
rect 3125 16170 3130 16190
rect 3130 16170 3150 16190
rect 3150 16170 3155 16190
rect 3125 16165 3155 16170
rect 3205 16190 3235 16195
rect 3205 16170 3210 16190
rect 3210 16170 3230 16190
rect 3230 16170 3235 16190
rect 3205 16165 3235 16170
rect 3285 16190 3315 16195
rect 3285 16170 3290 16190
rect 3290 16170 3310 16190
rect 3310 16170 3315 16190
rect 3285 16165 3315 16170
rect 3365 16190 3395 16195
rect 3365 16170 3370 16190
rect 3370 16170 3390 16190
rect 3390 16170 3395 16190
rect 3365 16165 3395 16170
rect 3445 16190 3475 16195
rect 3445 16170 3450 16190
rect 3450 16170 3470 16190
rect 3470 16170 3475 16190
rect 3445 16165 3475 16170
rect 3525 16190 3555 16195
rect 3525 16170 3530 16190
rect 3530 16170 3550 16190
rect 3550 16170 3555 16190
rect 3525 16165 3555 16170
rect 3605 16190 3635 16195
rect 3605 16170 3610 16190
rect 3610 16170 3630 16190
rect 3630 16170 3635 16190
rect 3605 16165 3635 16170
rect 3685 16190 3715 16195
rect 3685 16170 3690 16190
rect 3690 16170 3710 16190
rect 3710 16170 3715 16190
rect 3685 16165 3715 16170
rect 3765 16190 3795 16195
rect 3765 16170 3770 16190
rect 3770 16170 3790 16190
rect 3790 16170 3795 16190
rect 3765 16165 3795 16170
rect 3845 16190 3875 16195
rect 3845 16170 3850 16190
rect 3850 16170 3870 16190
rect 3870 16170 3875 16190
rect 3845 16165 3875 16170
rect 3925 16190 3955 16195
rect 3925 16170 3930 16190
rect 3930 16170 3950 16190
rect 3950 16170 3955 16190
rect 3925 16165 3955 16170
rect 4005 16190 4035 16195
rect 4005 16170 4010 16190
rect 4010 16170 4030 16190
rect 4030 16170 4035 16190
rect 4005 16165 4035 16170
rect 4085 16190 4115 16195
rect 4085 16170 4090 16190
rect 4090 16170 4110 16190
rect 4110 16170 4115 16190
rect 4085 16165 4115 16170
rect 4165 16190 4195 16195
rect 4165 16170 4170 16190
rect 4170 16170 4190 16190
rect 4190 16170 4195 16190
rect 4165 16165 4195 16170
rect 6245 16190 6275 16195
rect 6245 16170 6250 16190
rect 6250 16170 6270 16190
rect 6270 16170 6275 16190
rect 6245 16165 6275 16170
rect 6325 16190 6355 16195
rect 6325 16170 6330 16190
rect 6330 16170 6350 16190
rect 6350 16170 6355 16190
rect 6325 16165 6355 16170
rect 6405 16190 6435 16195
rect 6405 16170 6410 16190
rect 6410 16170 6430 16190
rect 6430 16170 6435 16190
rect 6405 16165 6435 16170
rect 6485 16190 6515 16195
rect 6485 16170 6490 16190
rect 6490 16170 6510 16190
rect 6510 16170 6515 16190
rect 6485 16165 6515 16170
rect 6565 16190 6595 16195
rect 6565 16170 6570 16190
rect 6570 16170 6590 16190
rect 6590 16170 6595 16190
rect 6565 16165 6595 16170
rect 6645 16190 6675 16195
rect 6645 16170 6650 16190
rect 6650 16170 6670 16190
rect 6670 16170 6675 16190
rect 6645 16165 6675 16170
rect 6725 16190 6755 16195
rect 6725 16170 6730 16190
rect 6730 16170 6750 16190
rect 6750 16170 6755 16190
rect 6725 16165 6755 16170
rect 6805 16190 6835 16195
rect 6805 16170 6810 16190
rect 6810 16170 6830 16190
rect 6830 16170 6835 16190
rect 6805 16165 6835 16170
rect 6885 16190 6915 16195
rect 6885 16170 6890 16190
rect 6890 16170 6910 16190
rect 6910 16170 6915 16190
rect 6885 16165 6915 16170
rect 6965 16190 6995 16195
rect 6965 16170 6970 16190
rect 6970 16170 6990 16190
rect 6990 16170 6995 16190
rect 6965 16165 6995 16170
rect 7045 16190 7075 16195
rect 7045 16170 7050 16190
rect 7050 16170 7070 16190
rect 7070 16170 7075 16190
rect 7045 16165 7075 16170
rect 7125 16190 7155 16195
rect 7125 16170 7130 16190
rect 7130 16170 7150 16190
rect 7150 16170 7155 16190
rect 7125 16165 7155 16170
rect 7205 16190 7235 16195
rect 7205 16170 7210 16190
rect 7210 16170 7230 16190
rect 7230 16170 7235 16190
rect 7205 16165 7235 16170
rect 7285 16190 7315 16195
rect 7285 16170 7290 16190
rect 7290 16170 7310 16190
rect 7310 16170 7315 16190
rect 7285 16165 7315 16170
rect 7365 16190 7395 16195
rect 7365 16170 7370 16190
rect 7370 16170 7390 16190
rect 7390 16170 7395 16190
rect 7365 16165 7395 16170
rect 7445 16190 7475 16195
rect 7445 16170 7450 16190
rect 7450 16170 7470 16190
rect 7470 16170 7475 16190
rect 7445 16165 7475 16170
rect 7525 16190 7555 16195
rect 7525 16170 7530 16190
rect 7530 16170 7550 16190
rect 7550 16170 7555 16190
rect 7525 16165 7555 16170
rect 7605 16190 7635 16195
rect 7605 16170 7610 16190
rect 7610 16170 7630 16190
rect 7630 16170 7635 16190
rect 7605 16165 7635 16170
rect 7685 16190 7715 16195
rect 7685 16170 7690 16190
rect 7690 16170 7710 16190
rect 7710 16170 7715 16190
rect 7685 16165 7715 16170
rect 7765 16190 7795 16195
rect 7765 16170 7770 16190
rect 7770 16170 7790 16190
rect 7790 16170 7795 16190
rect 7765 16165 7795 16170
rect 7845 16190 7875 16195
rect 7845 16170 7850 16190
rect 7850 16170 7870 16190
rect 7870 16170 7875 16190
rect 7845 16165 7875 16170
rect 7925 16190 7955 16195
rect 7925 16170 7930 16190
rect 7930 16170 7950 16190
rect 7950 16170 7955 16190
rect 7925 16165 7955 16170
rect 8005 16190 8035 16195
rect 8005 16170 8010 16190
rect 8010 16170 8030 16190
rect 8030 16170 8035 16190
rect 8005 16165 8035 16170
rect 8085 16190 8115 16195
rect 8085 16170 8090 16190
rect 8090 16170 8110 16190
rect 8110 16170 8115 16190
rect 8085 16165 8115 16170
rect 8165 16190 8195 16195
rect 8165 16170 8170 16190
rect 8170 16170 8190 16190
rect 8190 16170 8195 16190
rect 8165 16165 8195 16170
rect 8245 16190 8275 16195
rect 8245 16170 8250 16190
rect 8250 16170 8270 16190
rect 8270 16170 8275 16190
rect 8245 16165 8275 16170
rect 8325 16190 8355 16195
rect 8325 16170 8330 16190
rect 8330 16170 8350 16190
rect 8350 16170 8355 16190
rect 8325 16165 8355 16170
rect 8405 16190 8435 16195
rect 8405 16170 8410 16190
rect 8410 16170 8430 16190
rect 8430 16170 8435 16190
rect 8405 16165 8435 16170
rect 8485 16190 8515 16195
rect 8485 16170 8490 16190
rect 8490 16170 8510 16190
rect 8510 16170 8515 16190
rect 8485 16165 8515 16170
rect 8565 16190 8595 16195
rect 8565 16170 8570 16190
rect 8570 16170 8590 16190
rect 8590 16170 8595 16190
rect 8565 16165 8595 16170
rect 8645 16190 8675 16195
rect 8645 16170 8650 16190
rect 8650 16170 8670 16190
rect 8670 16170 8675 16190
rect 8645 16165 8675 16170
rect 8725 16190 8755 16195
rect 8725 16170 8730 16190
rect 8730 16170 8750 16190
rect 8750 16170 8755 16190
rect 8725 16165 8755 16170
rect 8805 16190 8835 16195
rect 8805 16170 8810 16190
rect 8810 16170 8830 16190
rect 8830 16170 8835 16190
rect 8805 16165 8835 16170
rect 8885 16190 8915 16195
rect 8885 16170 8890 16190
rect 8890 16170 8910 16190
rect 8910 16170 8915 16190
rect 8885 16165 8915 16170
rect 8965 16190 8995 16195
rect 8965 16170 8970 16190
rect 8970 16170 8990 16190
rect 8990 16170 8995 16190
rect 8965 16165 8995 16170
rect 9045 16190 9075 16195
rect 9045 16170 9050 16190
rect 9050 16170 9070 16190
rect 9070 16170 9075 16190
rect 9045 16165 9075 16170
rect 9125 16190 9155 16195
rect 9125 16170 9130 16190
rect 9130 16170 9150 16190
rect 9150 16170 9155 16190
rect 9125 16165 9155 16170
rect 9205 16190 9235 16195
rect 9205 16170 9210 16190
rect 9210 16170 9230 16190
rect 9230 16170 9235 16190
rect 9205 16165 9235 16170
rect 9285 16190 9315 16195
rect 9285 16170 9290 16190
rect 9290 16170 9310 16190
rect 9310 16170 9315 16190
rect 9285 16165 9315 16170
rect 9365 16190 9395 16195
rect 9365 16170 9370 16190
rect 9370 16170 9390 16190
rect 9390 16170 9395 16190
rect 9365 16165 9395 16170
rect 9445 16190 9475 16195
rect 9445 16170 9450 16190
rect 9450 16170 9470 16190
rect 9470 16170 9475 16190
rect 9445 16165 9475 16170
rect 11565 16190 11595 16195
rect 11565 16170 11570 16190
rect 11570 16170 11590 16190
rect 11590 16170 11595 16190
rect 11565 16165 11595 16170
rect 11645 16190 11675 16195
rect 11645 16170 11650 16190
rect 11650 16170 11670 16190
rect 11670 16170 11675 16190
rect 11645 16165 11675 16170
rect 11725 16190 11755 16195
rect 11725 16170 11730 16190
rect 11730 16170 11750 16190
rect 11750 16170 11755 16190
rect 11725 16165 11755 16170
rect 11805 16190 11835 16195
rect 11805 16170 11810 16190
rect 11810 16170 11830 16190
rect 11830 16170 11835 16190
rect 11805 16165 11835 16170
rect 11885 16190 11915 16195
rect 11885 16170 11890 16190
rect 11890 16170 11910 16190
rect 11910 16170 11915 16190
rect 11885 16165 11915 16170
rect 11965 16190 11995 16195
rect 11965 16170 11970 16190
rect 11970 16170 11990 16190
rect 11990 16170 11995 16190
rect 11965 16165 11995 16170
rect 12045 16190 12075 16195
rect 12045 16170 12050 16190
rect 12050 16170 12070 16190
rect 12070 16170 12075 16190
rect 12045 16165 12075 16170
rect 12125 16190 12155 16195
rect 12125 16170 12130 16190
rect 12130 16170 12150 16190
rect 12150 16170 12155 16190
rect 12125 16165 12155 16170
rect 12205 16190 12235 16195
rect 12205 16170 12210 16190
rect 12210 16170 12230 16190
rect 12230 16170 12235 16190
rect 12205 16165 12235 16170
rect 12285 16190 12315 16195
rect 12285 16170 12290 16190
rect 12290 16170 12310 16190
rect 12310 16170 12315 16190
rect 12285 16165 12315 16170
rect 12365 16190 12395 16195
rect 12365 16170 12370 16190
rect 12370 16170 12390 16190
rect 12390 16170 12395 16190
rect 12365 16165 12395 16170
rect 12445 16190 12475 16195
rect 12445 16170 12450 16190
rect 12450 16170 12470 16190
rect 12470 16170 12475 16190
rect 12445 16165 12475 16170
rect 12525 16190 12555 16195
rect 12525 16170 12530 16190
rect 12530 16170 12550 16190
rect 12550 16170 12555 16190
rect 12525 16165 12555 16170
rect 12605 16190 12635 16195
rect 12605 16170 12610 16190
rect 12610 16170 12630 16190
rect 12630 16170 12635 16190
rect 12605 16165 12635 16170
rect 12685 16190 12715 16195
rect 12685 16170 12690 16190
rect 12690 16170 12710 16190
rect 12710 16170 12715 16190
rect 12685 16165 12715 16170
rect 12765 16190 12795 16195
rect 12765 16170 12770 16190
rect 12770 16170 12790 16190
rect 12790 16170 12795 16190
rect 12765 16165 12795 16170
rect 12845 16190 12875 16195
rect 12845 16170 12850 16190
rect 12850 16170 12870 16190
rect 12870 16170 12875 16190
rect 12845 16165 12875 16170
rect 12925 16190 12955 16195
rect 12925 16170 12930 16190
rect 12930 16170 12950 16190
rect 12950 16170 12955 16190
rect 12925 16165 12955 16170
rect 13005 16190 13035 16195
rect 13005 16170 13010 16190
rect 13010 16170 13030 16190
rect 13030 16170 13035 16190
rect 13005 16165 13035 16170
rect 13085 16190 13115 16195
rect 13085 16170 13090 16190
rect 13090 16170 13110 16190
rect 13110 16170 13115 16190
rect 13085 16165 13115 16170
rect 13165 16190 13195 16195
rect 13165 16170 13170 16190
rect 13170 16170 13190 16190
rect 13190 16170 13195 16190
rect 13165 16165 13195 16170
rect 13245 16190 13275 16195
rect 13245 16170 13250 16190
rect 13250 16170 13270 16190
rect 13270 16170 13275 16190
rect 13245 16165 13275 16170
rect 13325 16190 13355 16195
rect 13325 16170 13330 16190
rect 13330 16170 13350 16190
rect 13350 16170 13355 16190
rect 13325 16165 13355 16170
rect 13405 16190 13435 16195
rect 13405 16170 13410 16190
rect 13410 16170 13430 16190
rect 13430 16170 13435 16190
rect 13405 16165 13435 16170
rect 13485 16190 13515 16195
rect 13485 16170 13490 16190
rect 13490 16170 13510 16190
rect 13510 16170 13515 16190
rect 13485 16165 13515 16170
rect 13565 16190 13595 16195
rect 13565 16170 13570 16190
rect 13570 16170 13590 16190
rect 13590 16170 13595 16190
rect 13565 16165 13595 16170
rect 13645 16190 13675 16195
rect 13645 16170 13650 16190
rect 13650 16170 13670 16190
rect 13670 16170 13675 16190
rect 13645 16165 13675 16170
rect 13725 16190 13755 16195
rect 13725 16170 13730 16190
rect 13730 16170 13750 16190
rect 13750 16170 13755 16190
rect 13725 16165 13755 16170
rect 13805 16190 13835 16195
rect 13805 16170 13810 16190
rect 13810 16170 13830 16190
rect 13830 16170 13835 16190
rect 13805 16165 13835 16170
rect 13885 16190 13915 16195
rect 13885 16170 13890 16190
rect 13890 16170 13910 16190
rect 13910 16170 13915 16190
rect 13885 16165 13915 16170
rect 13965 16190 13995 16195
rect 13965 16170 13970 16190
rect 13970 16170 13990 16190
rect 13990 16170 13995 16190
rect 13965 16165 13995 16170
rect 14045 16190 14075 16195
rect 14045 16170 14050 16190
rect 14050 16170 14070 16190
rect 14070 16170 14075 16190
rect 14045 16165 14075 16170
rect 14125 16190 14155 16195
rect 14125 16170 14130 16190
rect 14130 16170 14150 16190
rect 14150 16170 14155 16190
rect 14125 16165 14155 16170
rect 14205 16190 14235 16195
rect 14205 16170 14210 16190
rect 14210 16170 14230 16190
rect 14230 16170 14235 16190
rect 14205 16165 14235 16170
rect 14285 16190 14315 16195
rect 14285 16170 14290 16190
rect 14290 16170 14310 16190
rect 14310 16170 14315 16190
rect 14285 16165 14315 16170
rect 14365 16190 14395 16195
rect 14365 16170 14370 16190
rect 14370 16170 14390 16190
rect 14390 16170 14395 16190
rect 14365 16165 14395 16170
rect 14445 16190 14475 16195
rect 14445 16170 14450 16190
rect 14450 16170 14470 16190
rect 14470 16170 14475 16190
rect 14445 16165 14475 16170
rect 14525 16190 14555 16195
rect 14525 16170 14530 16190
rect 14530 16170 14550 16190
rect 14550 16170 14555 16190
rect 14525 16165 14555 16170
rect 14605 16190 14635 16195
rect 14605 16170 14610 16190
rect 14610 16170 14630 16190
rect 14630 16170 14635 16190
rect 14605 16165 14635 16170
rect 14685 16190 14715 16195
rect 14685 16170 14690 16190
rect 14690 16170 14710 16190
rect 14710 16170 14715 16190
rect 14685 16165 14715 16170
rect 16765 16190 16795 16195
rect 16765 16170 16770 16190
rect 16770 16170 16790 16190
rect 16790 16170 16795 16190
rect 16765 16165 16795 16170
rect 16845 16190 16875 16195
rect 16845 16170 16850 16190
rect 16850 16170 16870 16190
rect 16870 16170 16875 16190
rect 16845 16165 16875 16170
rect 16925 16190 16955 16195
rect 16925 16170 16930 16190
rect 16930 16170 16950 16190
rect 16950 16170 16955 16190
rect 16925 16165 16955 16170
rect 17005 16190 17035 16195
rect 17005 16170 17010 16190
rect 17010 16170 17030 16190
rect 17030 16170 17035 16190
rect 17005 16165 17035 16170
rect 17085 16190 17115 16195
rect 17085 16170 17090 16190
rect 17090 16170 17110 16190
rect 17110 16170 17115 16190
rect 17085 16165 17115 16170
rect 17165 16190 17195 16195
rect 17165 16170 17170 16190
rect 17170 16170 17190 16190
rect 17190 16170 17195 16190
rect 17165 16165 17195 16170
rect 17245 16190 17275 16195
rect 17245 16170 17250 16190
rect 17250 16170 17270 16190
rect 17270 16170 17275 16190
rect 17245 16165 17275 16170
rect 17325 16190 17355 16195
rect 17325 16170 17330 16190
rect 17330 16170 17350 16190
rect 17350 16170 17355 16190
rect 17325 16165 17355 16170
rect 17405 16190 17435 16195
rect 17405 16170 17410 16190
rect 17410 16170 17430 16190
rect 17430 16170 17435 16190
rect 17405 16165 17435 16170
rect 17485 16190 17515 16195
rect 17485 16170 17490 16190
rect 17490 16170 17510 16190
rect 17510 16170 17515 16190
rect 17485 16165 17515 16170
rect 17565 16190 17595 16195
rect 17565 16170 17570 16190
rect 17570 16170 17590 16190
rect 17590 16170 17595 16190
rect 17565 16165 17595 16170
rect 17645 16190 17675 16195
rect 17645 16170 17650 16190
rect 17650 16170 17670 16190
rect 17670 16170 17675 16190
rect 17645 16165 17675 16170
rect 17725 16190 17755 16195
rect 17725 16170 17730 16190
rect 17730 16170 17750 16190
rect 17750 16170 17755 16190
rect 17725 16165 17755 16170
rect 17805 16190 17835 16195
rect 17805 16170 17810 16190
rect 17810 16170 17830 16190
rect 17830 16170 17835 16190
rect 17805 16165 17835 16170
rect 17885 16190 17915 16195
rect 17885 16170 17890 16190
rect 17890 16170 17910 16190
rect 17910 16170 17915 16190
rect 17885 16165 17915 16170
rect 17965 16190 17995 16195
rect 17965 16170 17970 16190
rect 17970 16170 17990 16190
rect 17990 16170 17995 16190
rect 17965 16165 17995 16170
rect 18045 16190 18075 16195
rect 18045 16170 18050 16190
rect 18050 16170 18070 16190
rect 18070 16170 18075 16190
rect 18045 16165 18075 16170
rect 18125 16190 18155 16195
rect 18125 16170 18130 16190
rect 18130 16170 18150 16190
rect 18150 16170 18155 16190
rect 18125 16165 18155 16170
rect 18205 16190 18235 16195
rect 18205 16170 18210 16190
rect 18210 16170 18230 16190
rect 18230 16170 18235 16190
rect 18205 16165 18235 16170
rect 18285 16190 18315 16195
rect 18285 16170 18290 16190
rect 18290 16170 18310 16190
rect 18310 16170 18315 16190
rect 18285 16165 18315 16170
rect 18365 16190 18395 16195
rect 18365 16170 18370 16190
rect 18370 16170 18390 16190
rect 18390 16170 18395 16190
rect 18365 16165 18395 16170
rect 18445 16190 18475 16195
rect 18445 16170 18450 16190
rect 18450 16170 18470 16190
rect 18470 16170 18475 16190
rect 18445 16165 18475 16170
rect 18525 16190 18555 16195
rect 18525 16170 18530 16190
rect 18530 16170 18550 16190
rect 18550 16170 18555 16190
rect 18525 16165 18555 16170
rect 18605 16190 18635 16195
rect 18605 16170 18610 16190
rect 18610 16170 18630 16190
rect 18630 16170 18635 16190
rect 18605 16165 18635 16170
rect 18685 16190 18715 16195
rect 18685 16170 18690 16190
rect 18690 16170 18710 16190
rect 18710 16170 18715 16190
rect 18685 16165 18715 16170
rect 18765 16190 18795 16195
rect 18765 16170 18770 16190
rect 18770 16170 18790 16190
rect 18790 16170 18795 16190
rect 18765 16165 18795 16170
rect 18845 16190 18875 16195
rect 18845 16170 18850 16190
rect 18850 16170 18870 16190
rect 18870 16170 18875 16190
rect 18845 16165 18875 16170
rect 18925 16190 18955 16195
rect 18925 16170 18930 16190
rect 18930 16170 18950 16190
rect 18950 16170 18955 16190
rect 18925 16165 18955 16170
rect 19005 16190 19035 16195
rect 19005 16170 19010 16190
rect 19010 16170 19030 16190
rect 19030 16170 19035 16190
rect 19005 16165 19035 16170
rect 19085 16190 19115 16195
rect 19085 16170 19090 16190
rect 19090 16170 19110 16190
rect 19110 16170 19115 16190
rect 19085 16165 19115 16170
rect 19165 16190 19195 16195
rect 19165 16170 19170 16190
rect 19170 16170 19190 16190
rect 19190 16170 19195 16190
rect 19165 16165 19195 16170
rect 19245 16190 19275 16195
rect 19245 16170 19250 16190
rect 19250 16170 19270 16190
rect 19270 16170 19275 16190
rect 19245 16165 19275 16170
rect 19325 16190 19355 16195
rect 19325 16170 19330 16190
rect 19330 16170 19350 16190
rect 19350 16170 19355 16190
rect 19325 16165 19355 16170
rect 19405 16190 19435 16195
rect 19405 16170 19410 16190
rect 19410 16170 19430 16190
rect 19430 16170 19435 16190
rect 19405 16165 19435 16170
rect 19485 16190 19515 16195
rect 19485 16170 19490 16190
rect 19490 16170 19510 16190
rect 19510 16170 19515 16190
rect 19485 16165 19515 16170
rect 19565 16190 19595 16195
rect 19565 16170 19570 16190
rect 19570 16170 19590 16190
rect 19590 16170 19595 16190
rect 19565 16165 19595 16170
rect 19645 16190 19675 16195
rect 19645 16170 19650 16190
rect 19650 16170 19670 16190
rect 19670 16170 19675 16190
rect 19645 16165 19675 16170
rect 19725 16190 19755 16195
rect 19725 16170 19730 16190
rect 19730 16170 19750 16190
rect 19750 16170 19755 16190
rect 19725 16165 19755 16170
rect 19805 16190 19835 16195
rect 19805 16170 19810 16190
rect 19810 16170 19830 16190
rect 19830 16170 19835 16190
rect 19805 16165 19835 16170
rect 19885 16190 19915 16195
rect 19885 16170 19890 16190
rect 19890 16170 19910 16190
rect 19910 16170 19915 16190
rect 19885 16165 19915 16170
rect 19965 16190 19995 16195
rect 19965 16170 19970 16190
rect 19970 16170 19990 16190
rect 19990 16170 19995 16190
rect 19965 16165 19995 16170
rect 20045 16190 20075 16195
rect 20045 16170 20050 16190
rect 20050 16170 20070 16190
rect 20070 16170 20075 16190
rect 20045 16165 20075 16170
rect 20125 16190 20155 16195
rect 20125 16170 20130 16190
rect 20130 16170 20150 16190
rect 20150 16170 20155 16190
rect 20125 16165 20155 16170
rect 20205 16190 20235 16195
rect 20205 16170 20210 16190
rect 20210 16170 20230 16190
rect 20230 16170 20235 16190
rect 20205 16165 20235 16170
rect 20285 16190 20315 16195
rect 20285 16170 20290 16190
rect 20290 16170 20310 16190
rect 20310 16170 20315 16190
rect 20285 16165 20315 16170
rect 20365 16190 20395 16195
rect 20365 16170 20370 16190
rect 20370 16170 20390 16190
rect 20390 16170 20395 16190
rect 20365 16165 20395 16170
rect 20445 16190 20475 16195
rect 20445 16170 20450 16190
rect 20450 16170 20470 16190
rect 20470 16170 20475 16190
rect 20445 16165 20475 16170
rect 20525 16190 20555 16195
rect 20525 16170 20530 16190
rect 20530 16170 20550 16190
rect 20550 16170 20555 16190
rect 20525 16165 20555 16170
rect 20605 16190 20635 16195
rect 20605 16170 20610 16190
rect 20610 16170 20630 16190
rect 20630 16170 20635 16190
rect 20605 16165 20635 16170
rect 20685 16190 20715 16195
rect 20685 16170 20690 16190
rect 20690 16170 20710 16190
rect 20710 16170 20715 16190
rect 20685 16165 20715 16170
rect 20765 16190 20795 16195
rect 20765 16170 20770 16190
rect 20770 16170 20790 16190
rect 20790 16170 20795 16190
rect 20765 16165 20795 16170
rect 20845 16190 20875 16195
rect 20845 16170 20850 16190
rect 20850 16170 20870 16190
rect 20870 16170 20875 16190
rect 20845 16165 20875 16170
rect 20925 16190 20955 16195
rect 20925 16170 20930 16190
rect 20930 16170 20950 16190
rect 20950 16170 20955 16190
rect 20925 16165 20955 16170
rect 5 16030 35 16035
rect 5 16010 10 16030
rect 10 16010 30 16030
rect 30 16010 35 16030
rect 5 16005 35 16010
rect 85 16030 115 16035
rect 85 16010 90 16030
rect 90 16010 110 16030
rect 110 16010 115 16030
rect 85 16005 115 16010
rect 165 16030 195 16035
rect 165 16010 170 16030
rect 170 16010 190 16030
rect 190 16010 195 16030
rect 165 16005 195 16010
rect 245 16030 275 16035
rect 245 16010 250 16030
rect 250 16010 270 16030
rect 270 16010 275 16030
rect 245 16005 275 16010
rect 325 16030 355 16035
rect 325 16010 330 16030
rect 330 16010 350 16030
rect 350 16010 355 16030
rect 325 16005 355 16010
rect 405 16030 435 16035
rect 405 16010 410 16030
rect 410 16010 430 16030
rect 430 16010 435 16030
rect 405 16005 435 16010
rect 485 16030 515 16035
rect 485 16010 490 16030
rect 490 16010 510 16030
rect 510 16010 515 16030
rect 485 16005 515 16010
rect 565 16030 595 16035
rect 565 16010 570 16030
rect 570 16010 590 16030
rect 590 16010 595 16030
rect 565 16005 595 16010
rect 645 16030 675 16035
rect 645 16010 650 16030
rect 650 16010 670 16030
rect 670 16010 675 16030
rect 645 16005 675 16010
rect 725 16030 755 16035
rect 725 16010 730 16030
rect 730 16010 750 16030
rect 750 16010 755 16030
rect 725 16005 755 16010
rect 805 16030 835 16035
rect 805 16010 810 16030
rect 810 16010 830 16030
rect 830 16010 835 16030
rect 805 16005 835 16010
rect 885 16030 915 16035
rect 885 16010 890 16030
rect 890 16010 910 16030
rect 910 16010 915 16030
rect 885 16005 915 16010
rect 965 16030 995 16035
rect 965 16010 970 16030
rect 970 16010 990 16030
rect 990 16010 995 16030
rect 965 16005 995 16010
rect 1045 16030 1075 16035
rect 1045 16010 1050 16030
rect 1050 16010 1070 16030
rect 1070 16010 1075 16030
rect 1045 16005 1075 16010
rect 1125 16030 1155 16035
rect 1125 16010 1130 16030
rect 1130 16010 1150 16030
rect 1150 16010 1155 16030
rect 1125 16005 1155 16010
rect 1205 16030 1235 16035
rect 1205 16010 1210 16030
rect 1210 16010 1230 16030
rect 1230 16010 1235 16030
rect 1205 16005 1235 16010
rect 1285 16030 1315 16035
rect 1285 16010 1290 16030
rect 1290 16010 1310 16030
rect 1310 16010 1315 16030
rect 1285 16005 1315 16010
rect 1365 16030 1395 16035
rect 1365 16010 1370 16030
rect 1370 16010 1390 16030
rect 1390 16010 1395 16030
rect 1365 16005 1395 16010
rect 1445 16030 1475 16035
rect 1445 16010 1450 16030
rect 1450 16010 1470 16030
rect 1470 16010 1475 16030
rect 1445 16005 1475 16010
rect 1525 16030 1555 16035
rect 1525 16010 1530 16030
rect 1530 16010 1550 16030
rect 1550 16010 1555 16030
rect 1525 16005 1555 16010
rect 1605 16030 1635 16035
rect 1605 16010 1610 16030
rect 1610 16010 1630 16030
rect 1630 16010 1635 16030
rect 1605 16005 1635 16010
rect 1685 16030 1715 16035
rect 1685 16010 1690 16030
rect 1690 16010 1710 16030
rect 1710 16010 1715 16030
rect 1685 16005 1715 16010
rect 1765 16030 1795 16035
rect 1765 16010 1770 16030
rect 1770 16010 1790 16030
rect 1790 16010 1795 16030
rect 1765 16005 1795 16010
rect 1845 16030 1875 16035
rect 1845 16010 1850 16030
rect 1850 16010 1870 16030
rect 1870 16010 1875 16030
rect 1845 16005 1875 16010
rect 1925 16030 1955 16035
rect 1925 16010 1930 16030
rect 1930 16010 1950 16030
rect 1950 16010 1955 16030
rect 1925 16005 1955 16010
rect 2005 16030 2035 16035
rect 2005 16010 2010 16030
rect 2010 16010 2030 16030
rect 2030 16010 2035 16030
rect 2005 16005 2035 16010
rect 2085 16030 2115 16035
rect 2085 16010 2090 16030
rect 2090 16010 2110 16030
rect 2110 16010 2115 16030
rect 2085 16005 2115 16010
rect 2165 16030 2195 16035
rect 2165 16010 2170 16030
rect 2170 16010 2190 16030
rect 2190 16010 2195 16030
rect 2165 16005 2195 16010
rect 2245 16030 2275 16035
rect 2245 16010 2250 16030
rect 2250 16010 2270 16030
rect 2270 16010 2275 16030
rect 2245 16005 2275 16010
rect 2325 16030 2355 16035
rect 2325 16010 2330 16030
rect 2330 16010 2350 16030
rect 2350 16010 2355 16030
rect 2325 16005 2355 16010
rect 2405 16030 2435 16035
rect 2405 16010 2410 16030
rect 2410 16010 2430 16030
rect 2430 16010 2435 16030
rect 2405 16005 2435 16010
rect 2485 16030 2515 16035
rect 2485 16010 2490 16030
rect 2490 16010 2510 16030
rect 2510 16010 2515 16030
rect 2485 16005 2515 16010
rect 2565 16030 2595 16035
rect 2565 16010 2570 16030
rect 2570 16010 2590 16030
rect 2590 16010 2595 16030
rect 2565 16005 2595 16010
rect 2645 16030 2675 16035
rect 2645 16010 2650 16030
rect 2650 16010 2670 16030
rect 2670 16010 2675 16030
rect 2645 16005 2675 16010
rect 2725 16030 2755 16035
rect 2725 16010 2730 16030
rect 2730 16010 2750 16030
rect 2750 16010 2755 16030
rect 2725 16005 2755 16010
rect 2805 16030 2835 16035
rect 2805 16010 2810 16030
rect 2810 16010 2830 16030
rect 2830 16010 2835 16030
rect 2805 16005 2835 16010
rect 2885 16030 2915 16035
rect 2885 16010 2890 16030
rect 2890 16010 2910 16030
rect 2910 16010 2915 16030
rect 2885 16005 2915 16010
rect 2965 16030 2995 16035
rect 2965 16010 2970 16030
rect 2970 16010 2990 16030
rect 2990 16010 2995 16030
rect 2965 16005 2995 16010
rect 3045 16030 3075 16035
rect 3045 16010 3050 16030
rect 3050 16010 3070 16030
rect 3070 16010 3075 16030
rect 3045 16005 3075 16010
rect 3125 16030 3155 16035
rect 3125 16010 3130 16030
rect 3130 16010 3150 16030
rect 3150 16010 3155 16030
rect 3125 16005 3155 16010
rect 3205 16030 3235 16035
rect 3205 16010 3210 16030
rect 3210 16010 3230 16030
rect 3230 16010 3235 16030
rect 3205 16005 3235 16010
rect 3285 16030 3315 16035
rect 3285 16010 3290 16030
rect 3290 16010 3310 16030
rect 3310 16010 3315 16030
rect 3285 16005 3315 16010
rect 3365 16030 3395 16035
rect 3365 16010 3370 16030
rect 3370 16010 3390 16030
rect 3390 16010 3395 16030
rect 3365 16005 3395 16010
rect 3445 16030 3475 16035
rect 3445 16010 3450 16030
rect 3450 16010 3470 16030
rect 3470 16010 3475 16030
rect 3445 16005 3475 16010
rect 3525 16030 3555 16035
rect 3525 16010 3530 16030
rect 3530 16010 3550 16030
rect 3550 16010 3555 16030
rect 3525 16005 3555 16010
rect 3605 16030 3635 16035
rect 3605 16010 3610 16030
rect 3610 16010 3630 16030
rect 3630 16010 3635 16030
rect 3605 16005 3635 16010
rect 3685 16030 3715 16035
rect 3685 16010 3690 16030
rect 3690 16010 3710 16030
rect 3710 16010 3715 16030
rect 3685 16005 3715 16010
rect 3765 16030 3795 16035
rect 3765 16010 3770 16030
rect 3770 16010 3790 16030
rect 3790 16010 3795 16030
rect 3765 16005 3795 16010
rect 3845 16030 3875 16035
rect 3845 16010 3850 16030
rect 3850 16010 3870 16030
rect 3870 16010 3875 16030
rect 3845 16005 3875 16010
rect 3925 16030 3955 16035
rect 3925 16010 3930 16030
rect 3930 16010 3950 16030
rect 3950 16010 3955 16030
rect 3925 16005 3955 16010
rect 4005 16030 4035 16035
rect 4005 16010 4010 16030
rect 4010 16010 4030 16030
rect 4030 16010 4035 16030
rect 4005 16005 4035 16010
rect 4085 16030 4115 16035
rect 4085 16010 4090 16030
rect 4090 16010 4110 16030
rect 4110 16010 4115 16030
rect 4085 16005 4115 16010
rect 4165 16030 4195 16035
rect 4165 16010 4170 16030
rect 4170 16010 4190 16030
rect 4190 16010 4195 16030
rect 4165 16005 4195 16010
rect 6245 16030 6275 16035
rect 6245 16010 6250 16030
rect 6250 16010 6270 16030
rect 6270 16010 6275 16030
rect 6245 16005 6275 16010
rect 6325 16030 6355 16035
rect 6325 16010 6330 16030
rect 6330 16010 6350 16030
rect 6350 16010 6355 16030
rect 6325 16005 6355 16010
rect 6405 16030 6435 16035
rect 6405 16010 6410 16030
rect 6410 16010 6430 16030
rect 6430 16010 6435 16030
rect 6405 16005 6435 16010
rect 6485 16030 6515 16035
rect 6485 16010 6490 16030
rect 6490 16010 6510 16030
rect 6510 16010 6515 16030
rect 6485 16005 6515 16010
rect 6565 16030 6595 16035
rect 6565 16010 6570 16030
rect 6570 16010 6590 16030
rect 6590 16010 6595 16030
rect 6565 16005 6595 16010
rect 6645 16030 6675 16035
rect 6645 16010 6650 16030
rect 6650 16010 6670 16030
rect 6670 16010 6675 16030
rect 6645 16005 6675 16010
rect 6725 16030 6755 16035
rect 6725 16010 6730 16030
rect 6730 16010 6750 16030
rect 6750 16010 6755 16030
rect 6725 16005 6755 16010
rect 6805 16030 6835 16035
rect 6805 16010 6810 16030
rect 6810 16010 6830 16030
rect 6830 16010 6835 16030
rect 6805 16005 6835 16010
rect 6885 16030 6915 16035
rect 6885 16010 6890 16030
rect 6890 16010 6910 16030
rect 6910 16010 6915 16030
rect 6885 16005 6915 16010
rect 6965 16030 6995 16035
rect 6965 16010 6970 16030
rect 6970 16010 6990 16030
rect 6990 16010 6995 16030
rect 6965 16005 6995 16010
rect 7045 16030 7075 16035
rect 7045 16010 7050 16030
rect 7050 16010 7070 16030
rect 7070 16010 7075 16030
rect 7045 16005 7075 16010
rect 7125 16030 7155 16035
rect 7125 16010 7130 16030
rect 7130 16010 7150 16030
rect 7150 16010 7155 16030
rect 7125 16005 7155 16010
rect 7205 16030 7235 16035
rect 7205 16010 7210 16030
rect 7210 16010 7230 16030
rect 7230 16010 7235 16030
rect 7205 16005 7235 16010
rect 7285 16030 7315 16035
rect 7285 16010 7290 16030
rect 7290 16010 7310 16030
rect 7310 16010 7315 16030
rect 7285 16005 7315 16010
rect 7365 16030 7395 16035
rect 7365 16010 7370 16030
rect 7370 16010 7390 16030
rect 7390 16010 7395 16030
rect 7365 16005 7395 16010
rect 7445 16030 7475 16035
rect 7445 16010 7450 16030
rect 7450 16010 7470 16030
rect 7470 16010 7475 16030
rect 7445 16005 7475 16010
rect 7525 16030 7555 16035
rect 7525 16010 7530 16030
rect 7530 16010 7550 16030
rect 7550 16010 7555 16030
rect 7525 16005 7555 16010
rect 7605 16030 7635 16035
rect 7605 16010 7610 16030
rect 7610 16010 7630 16030
rect 7630 16010 7635 16030
rect 7605 16005 7635 16010
rect 7685 16030 7715 16035
rect 7685 16010 7690 16030
rect 7690 16010 7710 16030
rect 7710 16010 7715 16030
rect 7685 16005 7715 16010
rect 7765 16030 7795 16035
rect 7765 16010 7770 16030
rect 7770 16010 7790 16030
rect 7790 16010 7795 16030
rect 7765 16005 7795 16010
rect 7845 16030 7875 16035
rect 7845 16010 7850 16030
rect 7850 16010 7870 16030
rect 7870 16010 7875 16030
rect 7845 16005 7875 16010
rect 7925 16030 7955 16035
rect 7925 16010 7930 16030
rect 7930 16010 7950 16030
rect 7950 16010 7955 16030
rect 7925 16005 7955 16010
rect 8005 16030 8035 16035
rect 8005 16010 8010 16030
rect 8010 16010 8030 16030
rect 8030 16010 8035 16030
rect 8005 16005 8035 16010
rect 8085 16030 8115 16035
rect 8085 16010 8090 16030
rect 8090 16010 8110 16030
rect 8110 16010 8115 16030
rect 8085 16005 8115 16010
rect 8165 16030 8195 16035
rect 8165 16010 8170 16030
rect 8170 16010 8190 16030
rect 8190 16010 8195 16030
rect 8165 16005 8195 16010
rect 8245 16030 8275 16035
rect 8245 16010 8250 16030
rect 8250 16010 8270 16030
rect 8270 16010 8275 16030
rect 8245 16005 8275 16010
rect 8325 16030 8355 16035
rect 8325 16010 8330 16030
rect 8330 16010 8350 16030
rect 8350 16010 8355 16030
rect 8325 16005 8355 16010
rect 8405 16030 8435 16035
rect 8405 16010 8410 16030
rect 8410 16010 8430 16030
rect 8430 16010 8435 16030
rect 8405 16005 8435 16010
rect 8485 16030 8515 16035
rect 8485 16010 8490 16030
rect 8490 16010 8510 16030
rect 8510 16010 8515 16030
rect 8485 16005 8515 16010
rect 8565 16030 8595 16035
rect 8565 16010 8570 16030
rect 8570 16010 8590 16030
rect 8590 16010 8595 16030
rect 8565 16005 8595 16010
rect 8645 16030 8675 16035
rect 8645 16010 8650 16030
rect 8650 16010 8670 16030
rect 8670 16010 8675 16030
rect 8645 16005 8675 16010
rect 8725 16030 8755 16035
rect 8725 16010 8730 16030
rect 8730 16010 8750 16030
rect 8750 16010 8755 16030
rect 8725 16005 8755 16010
rect 8805 16030 8835 16035
rect 8805 16010 8810 16030
rect 8810 16010 8830 16030
rect 8830 16010 8835 16030
rect 8805 16005 8835 16010
rect 8885 16030 8915 16035
rect 8885 16010 8890 16030
rect 8890 16010 8910 16030
rect 8910 16010 8915 16030
rect 8885 16005 8915 16010
rect 8965 16030 8995 16035
rect 8965 16010 8970 16030
rect 8970 16010 8990 16030
rect 8990 16010 8995 16030
rect 8965 16005 8995 16010
rect 9045 16030 9075 16035
rect 9045 16010 9050 16030
rect 9050 16010 9070 16030
rect 9070 16010 9075 16030
rect 9045 16005 9075 16010
rect 9125 16030 9155 16035
rect 9125 16010 9130 16030
rect 9130 16010 9150 16030
rect 9150 16010 9155 16030
rect 9125 16005 9155 16010
rect 9205 16030 9235 16035
rect 9205 16010 9210 16030
rect 9210 16010 9230 16030
rect 9230 16010 9235 16030
rect 9205 16005 9235 16010
rect 9285 16030 9315 16035
rect 9285 16010 9290 16030
rect 9290 16010 9310 16030
rect 9310 16010 9315 16030
rect 9285 16005 9315 16010
rect 9365 16030 9395 16035
rect 9365 16010 9370 16030
rect 9370 16010 9390 16030
rect 9390 16010 9395 16030
rect 9365 16005 9395 16010
rect 9445 16030 9475 16035
rect 9445 16010 9450 16030
rect 9450 16010 9470 16030
rect 9470 16010 9475 16030
rect 9445 16005 9475 16010
rect 11565 16030 11595 16035
rect 11565 16010 11570 16030
rect 11570 16010 11590 16030
rect 11590 16010 11595 16030
rect 11565 16005 11595 16010
rect 11645 16030 11675 16035
rect 11645 16010 11650 16030
rect 11650 16010 11670 16030
rect 11670 16010 11675 16030
rect 11645 16005 11675 16010
rect 11725 16030 11755 16035
rect 11725 16010 11730 16030
rect 11730 16010 11750 16030
rect 11750 16010 11755 16030
rect 11725 16005 11755 16010
rect 11805 16030 11835 16035
rect 11805 16010 11810 16030
rect 11810 16010 11830 16030
rect 11830 16010 11835 16030
rect 11805 16005 11835 16010
rect 11885 16030 11915 16035
rect 11885 16010 11890 16030
rect 11890 16010 11910 16030
rect 11910 16010 11915 16030
rect 11885 16005 11915 16010
rect 11965 16030 11995 16035
rect 11965 16010 11970 16030
rect 11970 16010 11990 16030
rect 11990 16010 11995 16030
rect 11965 16005 11995 16010
rect 12045 16030 12075 16035
rect 12045 16010 12050 16030
rect 12050 16010 12070 16030
rect 12070 16010 12075 16030
rect 12045 16005 12075 16010
rect 12125 16030 12155 16035
rect 12125 16010 12130 16030
rect 12130 16010 12150 16030
rect 12150 16010 12155 16030
rect 12125 16005 12155 16010
rect 12205 16030 12235 16035
rect 12205 16010 12210 16030
rect 12210 16010 12230 16030
rect 12230 16010 12235 16030
rect 12205 16005 12235 16010
rect 12285 16030 12315 16035
rect 12285 16010 12290 16030
rect 12290 16010 12310 16030
rect 12310 16010 12315 16030
rect 12285 16005 12315 16010
rect 12365 16030 12395 16035
rect 12365 16010 12370 16030
rect 12370 16010 12390 16030
rect 12390 16010 12395 16030
rect 12365 16005 12395 16010
rect 12445 16030 12475 16035
rect 12445 16010 12450 16030
rect 12450 16010 12470 16030
rect 12470 16010 12475 16030
rect 12445 16005 12475 16010
rect 12525 16030 12555 16035
rect 12525 16010 12530 16030
rect 12530 16010 12550 16030
rect 12550 16010 12555 16030
rect 12525 16005 12555 16010
rect 12605 16030 12635 16035
rect 12605 16010 12610 16030
rect 12610 16010 12630 16030
rect 12630 16010 12635 16030
rect 12605 16005 12635 16010
rect 12685 16030 12715 16035
rect 12685 16010 12690 16030
rect 12690 16010 12710 16030
rect 12710 16010 12715 16030
rect 12685 16005 12715 16010
rect 12765 16030 12795 16035
rect 12765 16010 12770 16030
rect 12770 16010 12790 16030
rect 12790 16010 12795 16030
rect 12765 16005 12795 16010
rect 12845 16030 12875 16035
rect 12845 16010 12850 16030
rect 12850 16010 12870 16030
rect 12870 16010 12875 16030
rect 12845 16005 12875 16010
rect 12925 16030 12955 16035
rect 12925 16010 12930 16030
rect 12930 16010 12950 16030
rect 12950 16010 12955 16030
rect 12925 16005 12955 16010
rect 13005 16030 13035 16035
rect 13005 16010 13010 16030
rect 13010 16010 13030 16030
rect 13030 16010 13035 16030
rect 13005 16005 13035 16010
rect 13085 16030 13115 16035
rect 13085 16010 13090 16030
rect 13090 16010 13110 16030
rect 13110 16010 13115 16030
rect 13085 16005 13115 16010
rect 13165 16030 13195 16035
rect 13165 16010 13170 16030
rect 13170 16010 13190 16030
rect 13190 16010 13195 16030
rect 13165 16005 13195 16010
rect 13245 16030 13275 16035
rect 13245 16010 13250 16030
rect 13250 16010 13270 16030
rect 13270 16010 13275 16030
rect 13245 16005 13275 16010
rect 13325 16030 13355 16035
rect 13325 16010 13330 16030
rect 13330 16010 13350 16030
rect 13350 16010 13355 16030
rect 13325 16005 13355 16010
rect 13405 16030 13435 16035
rect 13405 16010 13410 16030
rect 13410 16010 13430 16030
rect 13430 16010 13435 16030
rect 13405 16005 13435 16010
rect 13485 16030 13515 16035
rect 13485 16010 13490 16030
rect 13490 16010 13510 16030
rect 13510 16010 13515 16030
rect 13485 16005 13515 16010
rect 13565 16030 13595 16035
rect 13565 16010 13570 16030
rect 13570 16010 13590 16030
rect 13590 16010 13595 16030
rect 13565 16005 13595 16010
rect 13645 16030 13675 16035
rect 13645 16010 13650 16030
rect 13650 16010 13670 16030
rect 13670 16010 13675 16030
rect 13645 16005 13675 16010
rect 13725 16030 13755 16035
rect 13725 16010 13730 16030
rect 13730 16010 13750 16030
rect 13750 16010 13755 16030
rect 13725 16005 13755 16010
rect 13805 16030 13835 16035
rect 13805 16010 13810 16030
rect 13810 16010 13830 16030
rect 13830 16010 13835 16030
rect 13805 16005 13835 16010
rect 13885 16030 13915 16035
rect 13885 16010 13890 16030
rect 13890 16010 13910 16030
rect 13910 16010 13915 16030
rect 13885 16005 13915 16010
rect 13965 16030 13995 16035
rect 13965 16010 13970 16030
rect 13970 16010 13990 16030
rect 13990 16010 13995 16030
rect 13965 16005 13995 16010
rect 14045 16030 14075 16035
rect 14045 16010 14050 16030
rect 14050 16010 14070 16030
rect 14070 16010 14075 16030
rect 14045 16005 14075 16010
rect 14125 16030 14155 16035
rect 14125 16010 14130 16030
rect 14130 16010 14150 16030
rect 14150 16010 14155 16030
rect 14125 16005 14155 16010
rect 14205 16030 14235 16035
rect 14205 16010 14210 16030
rect 14210 16010 14230 16030
rect 14230 16010 14235 16030
rect 14205 16005 14235 16010
rect 14285 16030 14315 16035
rect 14285 16010 14290 16030
rect 14290 16010 14310 16030
rect 14310 16010 14315 16030
rect 14285 16005 14315 16010
rect 14365 16030 14395 16035
rect 14365 16010 14370 16030
rect 14370 16010 14390 16030
rect 14390 16010 14395 16030
rect 14365 16005 14395 16010
rect 14445 16030 14475 16035
rect 14445 16010 14450 16030
rect 14450 16010 14470 16030
rect 14470 16010 14475 16030
rect 14445 16005 14475 16010
rect 14525 16030 14555 16035
rect 14525 16010 14530 16030
rect 14530 16010 14550 16030
rect 14550 16010 14555 16030
rect 14525 16005 14555 16010
rect 14605 16030 14635 16035
rect 14605 16010 14610 16030
rect 14610 16010 14630 16030
rect 14630 16010 14635 16030
rect 14605 16005 14635 16010
rect 14685 16030 14715 16035
rect 14685 16010 14690 16030
rect 14690 16010 14710 16030
rect 14710 16010 14715 16030
rect 14685 16005 14715 16010
rect 16765 16030 16795 16035
rect 16765 16010 16770 16030
rect 16770 16010 16790 16030
rect 16790 16010 16795 16030
rect 16765 16005 16795 16010
rect 16845 16030 16875 16035
rect 16845 16010 16850 16030
rect 16850 16010 16870 16030
rect 16870 16010 16875 16030
rect 16845 16005 16875 16010
rect 16925 16030 16955 16035
rect 16925 16010 16930 16030
rect 16930 16010 16950 16030
rect 16950 16010 16955 16030
rect 16925 16005 16955 16010
rect 17005 16030 17035 16035
rect 17005 16010 17010 16030
rect 17010 16010 17030 16030
rect 17030 16010 17035 16030
rect 17005 16005 17035 16010
rect 17085 16030 17115 16035
rect 17085 16010 17090 16030
rect 17090 16010 17110 16030
rect 17110 16010 17115 16030
rect 17085 16005 17115 16010
rect 17165 16030 17195 16035
rect 17165 16010 17170 16030
rect 17170 16010 17190 16030
rect 17190 16010 17195 16030
rect 17165 16005 17195 16010
rect 17245 16030 17275 16035
rect 17245 16010 17250 16030
rect 17250 16010 17270 16030
rect 17270 16010 17275 16030
rect 17245 16005 17275 16010
rect 17325 16030 17355 16035
rect 17325 16010 17330 16030
rect 17330 16010 17350 16030
rect 17350 16010 17355 16030
rect 17325 16005 17355 16010
rect 17405 16030 17435 16035
rect 17405 16010 17410 16030
rect 17410 16010 17430 16030
rect 17430 16010 17435 16030
rect 17405 16005 17435 16010
rect 17485 16030 17515 16035
rect 17485 16010 17490 16030
rect 17490 16010 17510 16030
rect 17510 16010 17515 16030
rect 17485 16005 17515 16010
rect 17565 16030 17595 16035
rect 17565 16010 17570 16030
rect 17570 16010 17590 16030
rect 17590 16010 17595 16030
rect 17565 16005 17595 16010
rect 17645 16030 17675 16035
rect 17645 16010 17650 16030
rect 17650 16010 17670 16030
rect 17670 16010 17675 16030
rect 17645 16005 17675 16010
rect 17725 16030 17755 16035
rect 17725 16010 17730 16030
rect 17730 16010 17750 16030
rect 17750 16010 17755 16030
rect 17725 16005 17755 16010
rect 17805 16030 17835 16035
rect 17805 16010 17810 16030
rect 17810 16010 17830 16030
rect 17830 16010 17835 16030
rect 17805 16005 17835 16010
rect 17885 16030 17915 16035
rect 17885 16010 17890 16030
rect 17890 16010 17910 16030
rect 17910 16010 17915 16030
rect 17885 16005 17915 16010
rect 17965 16030 17995 16035
rect 17965 16010 17970 16030
rect 17970 16010 17990 16030
rect 17990 16010 17995 16030
rect 17965 16005 17995 16010
rect 18045 16030 18075 16035
rect 18045 16010 18050 16030
rect 18050 16010 18070 16030
rect 18070 16010 18075 16030
rect 18045 16005 18075 16010
rect 18125 16030 18155 16035
rect 18125 16010 18130 16030
rect 18130 16010 18150 16030
rect 18150 16010 18155 16030
rect 18125 16005 18155 16010
rect 18205 16030 18235 16035
rect 18205 16010 18210 16030
rect 18210 16010 18230 16030
rect 18230 16010 18235 16030
rect 18205 16005 18235 16010
rect 18285 16030 18315 16035
rect 18285 16010 18290 16030
rect 18290 16010 18310 16030
rect 18310 16010 18315 16030
rect 18285 16005 18315 16010
rect 18365 16030 18395 16035
rect 18365 16010 18370 16030
rect 18370 16010 18390 16030
rect 18390 16010 18395 16030
rect 18365 16005 18395 16010
rect 18445 16030 18475 16035
rect 18445 16010 18450 16030
rect 18450 16010 18470 16030
rect 18470 16010 18475 16030
rect 18445 16005 18475 16010
rect 18525 16030 18555 16035
rect 18525 16010 18530 16030
rect 18530 16010 18550 16030
rect 18550 16010 18555 16030
rect 18525 16005 18555 16010
rect 18605 16030 18635 16035
rect 18605 16010 18610 16030
rect 18610 16010 18630 16030
rect 18630 16010 18635 16030
rect 18605 16005 18635 16010
rect 18685 16030 18715 16035
rect 18685 16010 18690 16030
rect 18690 16010 18710 16030
rect 18710 16010 18715 16030
rect 18685 16005 18715 16010
rect 18765 16030 18795 16035
rect 18765 16010 18770 16030
rect 18770 16010 18790 16030
rect 18790 16010 18795 16030
rect 18765 16005 18795 16010
rect 18845 16030 18875 16035
rect 18845 16010 18850 16030
rect 18850 16010 18870 16030
rect 18870 16010 18875 16030
rect 18845 16005 18875 16010
rect 18925 16030 18955 16035
rect 18925 16010 18930 16030
rect 18930 16010 18950 16030
rect 18950 16010 18955 16030
rect 18925 16005 18955 16010
rect 19005 16030 19035 16035
rect 19005 16010 19010 16030
rect 19010 16010 19030 16030
rect 19030 16010 19035 16030
rect 19005 16005 19035 16010
rect 19085 16030 19115 16035
rect 19085 16010 19090 16030
rect 19090 16010 19110 16030
rect 19110 16010 19115 16030
rect 19085 16005 19115 16010
rect 19165 16030 19195 16035
rect 19165 16010 19170 16030
rect 19170 16010 19190 16030
rect 19190 16010 19195 16030
rect 19165 16005 19195 16010
rect 19245 16030 19275 16035
rect 19245 16010 19250 16030
rect 19250 16010 19270 16030
rect 19270 16010 19275 16030
rect 19245 16005 19275 16010
rect 19325 16030 19355 16035
rect 19325 16010 19330 16030
rect 19330 16010 19350 16030
rect 19350 16010 19355 16030
rect 19325 16005 19355 16010
rect 19405 16030 19435 16035
rect 19405 16010 19410 16030
rect 19410 16010 19430 16030
rect 19430 16010 19435 16030
rect 19405 16005 19435 16010
rect 19485 16030 19515 16035
rect 19485 16010 19490 16030
rect 19490 16010 19510 16030
rect 19510 16010 19515 16030
rect 19485 16005 19515 16010
rect 19565 16030 19595 16035
rect 19565 16010 19570 16030
rect 19570 16010 19590 16030
rect 19590 16010 19595 16030
rect 19565 16005 19595 16010
rect 19645 16030 19675 16035
rect 19645 16010 19650 16030
rect 19650 16010 19670 16030
rect 19670 16010 19675 16030
rect 19645 16005 19675 16010
rect 19725 16030 19755 16035
rect 19725 16010 19730 16030
rect 19730 16010 19750 16030
rect 19750 16010 19755 16030
rect 19725 16005 19755 16010
rect 19805 16030 19835 16035
rect 19805 16010 19810 16030
rect 19810 16010 19830 16030
rect 19830 16010 19835 16030
rect 19805 16005 19835 16010
rect 19885 16030 19915 16035
rect 19885 16010 19890 16030
rect 19890 16010 19910 16030
rect 19910 16010 19915 16030
rect 19885 16005 19915 16010
rect 19965 16030 19995 16035
rect 19965 16010 19970 16030
rect 19970 16010 19990 16030
rect 19990 16010 19995 16030
rect 19965 16005 19995 16010
rect 20045 16030 20075 16035
rect 20045 16010 20050 16030
rect 20050 16010 20070 16030
rect 20070 16010 20075 16030
rect 20045 16005 20075 16010
rect 20125 16030 20155 16035
rect 20125 16010 20130 16030
rect 20130 16010 20150 16030
rect 20150 16010 20155 16030
rect 20125 16005 20155 16010
rect 20205 16030 20235 16035
rect 20205 16010 20210 16030
rect 20210 16010 20230 16030
rect 20230 16010 20235 16030
rect 20205 16005 20235 16010
rect 20285 16030 20315 16035
rect 20285 16010 20290 16030
rect 20290 16010 20310 16030
rect 20310 16010 20315 16030
rect 20285 16005 20315 16010
rect 20365 16030 20395 16035
rect 20365 16010 20370 16030
rect 20370 16010 20390 16030
rect 20390 16010 20395 16030
rect 20365 16005 20395 16010
rect 20445 16030 20475 16035
rect 20445 16010 20450 16030
rect 20450 16010 20470 16030
rect 20470 16010 20475 16030
rect 20445 16005 20475 16010
rect 20525 16030 20555 16035
rect 20525 16010 20530 16030
rect 20530 16010 20550 16030
rect 20550 16010 20555 16030
rect 20525 16005 20555 16010
rect 20605 16030 20635 16035
rect 20605 16010 20610 16030
rect 20610 16010 20630 16030
rect 20630 16010 20635 16030
rect 20605 16005 20635 16010
rect 20685 16030 20715 16035
rect 20685 16010 20690 16030
rect 20690 16010 20710 16030
rect 20710 16010 20715 16030
rect 20685 16005 20715 16010
rect 20765 16030 20795 16035
rect 20765 16010 20770 16030
rect 20770 16010 20790 16030
rect 20790 16010 20795 16030
rect 20765 16005 20795 16010
rect 20845 16030 20875 16035
rect 20845 16010 20850 16030
rect 20850 16010 20870 16030
rect 20870 16010 20875 16030
rect 20845 16005 20875 16010
rect 20925 16030 20955 16035
rect 20925 16010 20930 16030
rect 20930 16010 20950 16030
rect 20950 16010 20955 16030
rect 20925 16005 20955 16010
rect 5 15870 35 15875
rect 5 15850 10 15870
rect 10 15850 30 15870
rect 30 15850 35 15870
rect 5 15845 35 15850
rect 85 15870 115 15875
rect 85 15850 90 15870
rect 90 15850 110 15870
rect 110 15850 115 15870
rect 85 15845 115 15850
rect 165 15870 195 15875
rect 165 15850 170 15870
rect 170 15850 190 15870
rect 190 15850 195 15870
rect 165 15845 195 15850
rect 245 15870 275 15875
rect 245 15850 250 15870
rect 250 15850 270 15870
rect 270 15850 275 15870
rect 245 15845 275 15850
rect 325 15870 355 15875
rect 325 15850 330 15870
rect 330 15850 350 15870
rect 350 15850 355 15870
rect 325 15845 355 15850
rect 405 15870 435 15875
rect 405 15850 410 15870
rect 410 15850 430 15870
rect 430 15850 435 15870
rect 405 15845 435 15850
rect 485 15870 515 15875
rect 485 15850 490 15870
rect 490 15850 510 15870
rect 510 15850 515 15870
rect 485 15845 515 15850
rect 565 15870 595 15875
rect 565 15850 570 15870
rect 570 15850 590 15870
rect 590 15850 595 15870
rect 565 15845 595 15850
rect 645 15870 675 15875
rect 645 15850 650 15870
rect 650 15850 670 15870
rect 670 15850 675 15870
rect 645 15845 675 15850
rect 725 15870 755 15875
rect 725 15850 730 15870
rect 730 15850 750 15870
rect 750 15850 755 15870
rect 725 15845 755 15850
rect 805 15870 835 15875
rect 805 15850 810 15870
rect 810 15850 830 15870
rect 830 15850 835 15870
rect 805 15845 835 15850
rect 885 15870 915 15875
rect 885 15850 890 15870
rect 890 15850 910 15870
rect 910 15850 915 15870
rect 885 15845 915 15850
rect 965 15870 995 15875
rect 965 15850 970 15870
rect 970 15850 990 15870
rect 990 15850 995 15870
rect 965 15845 995 15850
rect 1045 15870 1075 15875
rect 1045 15850 1050 15870
rect 1050 15850 1070 15870
rect 1070 15850 1075 15870
rect 1045 15845 1075 15850
rect 1125 15870 1155 15875
rect 1125 15850 1130 15870
rect 1130 15850 1150 15870
rect 1150 15850 1155 15870
rect 1125 15845 1155 15850
rect 1205 15870 1235 15875
rect 1205 15850 1210 15870
rect 1210 15850 1230 15870
rect 1230 15850 1235 15870
rect 1205 15845 1235 15850
rect 1285 15870 1315 15875
rect 1285 15850 1290 15870
rect 1290 15850 1310 15870
rect 1310 15850 1315 15870
rect 1285 15845 1315 15850
rect 1365 15870 1395 15875
rect 1365 15850 1370 15870
rect 1370 15850 1390 15870
rect 1390 15850 1395 15870
rect 1365 15845 1395 15850
rect 1445 15870 1475 15875
rect 1445 15850 1450 15870
rect 1450 15850 1470 15870
rect 1470 15850 1475 15870
rect 1445 15845 1475 15850
rect 1525 15870 1555 15875
rect 1525 15850 1530 15870
rect 1530 15850 1550 15870
rect 1550 15850 1555 15870
rect 1525 15845 1555 15850
rect 1605 15870 1635 15875
rect 1605 15850 1610 15870
rect 1610 15850 1630 15870
rect 1630 15850 1635 15870
rect 1605 15845 1635 15850
rect 1685 15870 1715 15875
rect 1685 15850 1690 15870
rect 1690 15850 1710 15870
rect 1710 15850 1715 15870
rect 1685 15845 1715 15850
rect 1765 15870 1795 15875
rect 1765 15850 1770 15870
rect 1770 15850 1790 15870
rect 1790 15850 1795 15870
rect 1765 15845 1795 15850
rect 1845 15870 1875 15875
rect 1845 15850 1850 15870
rect 1850 15850 1870 15870
rect 1870 15850 1875 15870
rect 1845 15845 1875 15850
rect 1925 15870 1955 15875
rect 1925 15850 1930 15870
rect 1930 15850 1950 15870
rect 1950 15850 1955 15870
rect 1925 15845 1955 15850
rect 2005 15870 2035 15875
rect 2005 15850 2010 15870
rect 2010 15850 2030 15870
rect 2030 15850 2035 15870
rect 2005 15845 2035 15850
rect 2085 15870 2115 15875
rect 2085 15850 2090 15870
rect 2090 15850 2110 15870
rect 2110 15850 2115 15870
rect 2085 15845 2115 15850
rect 2165 15870 2195 15875
rect 2165 15850 2170 15870
rect 2170 15850 2190 15870
rect 2190 15850 2195 15870
rect 2165 15845 2195 15850
rect 2245 15870 2275 15875
rect 2245 15850 2250 15870
rect 2250 15850 2270 15870
rect 2270 15850 2275 15870
rect 2245 15845 2275 15850
rect 2325 15870 2355 15875
rect 2325 15850 2330 15870
rect 2330 15850 2350 15870
rect 2350 15850 2355 15870
rect 2325 15845 2355 15850
rect 2405 15870 2435 15875
rect 2405 15850 2410 15870
rect 2410 15850 2430 15870
rect 2430 15850 2435 15870
rect 2405 15845 2435 15850
rect 2485 15870 2515 15875
rect 2485 15850 2490 15870
rect 2490 15850 2510 15870
rect 2510 15850 2515 15870
rect 2485 15845 2515 15850
rect 2565 15870 2595 15875
rect 2565 15850 2570 15870
rect 2570 15850 2590 15870
rect 2590 15850 2595 15870
rect 2565 15845 2595 15850
rect 2645 15870 2675 15875
rect 2645 15850 2650 15870
rect 2650 15850 2670 15870
rect 2670 15850 2675 15870
rect 2645 15845 2675 15850
rect 2725 15870 2755 15875
rect 2725 15850 2730 15870
rect 2730 15850 2750 15870
rect 2750 15850 2755 15870
rect 2725 15845 2755 15850
rect 2805 15870 2835 15875
rect 2805 15850 2810 15870
rect 2810 15850 2830 15870
rect 2830 15850 2835 15870
rect 2805 15845 2835 15850
rect 2885 15870 2915 15875
rect 2885 15850 2890 15870
rect 2890 15850 2910 15870
rect 2910 15850 2915 15870
rect 2885 15845 2915 15850
rect 2965 15870 2995 15875
rect 2965 15850 2970 15870
rect 2970 15850 2990 15870
rect 2990 15850 2995 15870
rect 2965 15845 2995 15850
rect 3045 15870 3075 15875
rect 3045 15850 3050 15870
rect 3050 15850 3070 15870
rect 3070 15850 3075 15870
rect 3045 15845 3075 15850
rect 3125 15870 3155 15875
rect 3125 15850 3130 15870
rect 3130 15850 3150 15870
rect 3150 15850 3155 15870
rect 3125 15845 3155 15850
rect 3205 15870 3235 15875
rect 3205 15850 3210 15870
rect 3210 15850 3230 15870
rect 3230 15850 3235 15870
rect 3205 15845 3235 15850
rect 3285 15870 3315 15875
rect 3285 15850 3290 15870
rect 3290 15850 3310 15870
rect 3310 15850 3315 15870
rect 3285 15845 3315 15850
rect 3365 15870 3395 15875
rect 3365 15850 3370 15870
rect 3370 15850 3390 15870
rect 3390 15850 3395 15870
rect 3365 15845 3395 15850
rect 3445 15870 3475 15875
rect 3445 15850 3450 15870
rect 3450 15850 3470 15870
rect 3470 15850 3475 15870
rect 3445 15845 3475 15850
rect 3525 15870 3555 15875
rect 3525 15850 3530 15870
rect 3530 15850 3550 15870
rect 3550 15850 3555 15870
rect 3525 15845 3555 15850
rect 3605 15870 3635 15875
rect 3605 15850 3610 15870
rect 3610 15850 3630 15870
rect 3630 15850 3635 15870
rect 3605 15845 3635 15850
rect 3685 15870 3715 15875
rect 3685 15850 3690 15870
rect 3690 15850 3710 15870
rect 3710 15850 3715 15870
rect 3685 15845 3715 15850
rect 3765 15870 3795 15875
rect 3765 15850 3770 15870
rect 3770 15850 3790 15870
rect 3790 15850 3795 15870
rect 3765 15845 3795 15850
rect 3845 15870 3875 15875
rect 3845 15850 3850 15870
rect 3850 15850 3870 15870
rect 3870 15850 3875 15870
rect 3845 15845 3875 15850
rect 3925 15870 3955 15875
rect 3925 15850 3930 15870
rect 3930 15850 3950 15870
rect 3950 15850 3955 15870
rect 3925 15845 3955 15850
rect 4005 15870 4035 15875
rect 4005 15850 4010 15870
rect 4010 15850 4030 15870
rect 4030 15850 4035 15870
rect 4005 15845 4035 15850
rect 4085 15870 4115 15875
rect 4085 15850 4090 15870
rect 4090 15850 4110 15870
rect 4110 15850 4115 15870
rect 4085 15845 4115 15850
rect 4165 15870 4195 15875
rect 4165 15850 4170 15870
rect 4170 15850 4190 15870
rect 4190 15850 4195 15870
rect 4165 15845 4195 15850
rect 6245 15870 6275 15875
rect 6245 15850 6250 15870
rect 6250 15850 6270 15870
rect 6270 15850 6275 15870
rect 6245 15845 6275 15850
rect 6325 15870 6355 15875
rect 6325 15850 6330 15870
rect 6330 15850 6350 15870
rect 6350 15850 6355 15870
rect 6325 15845 6355 15850
rect 6405 15870 6435 15875
rect 6405 15850 6410 15870
rect 6410 15850 6430 15870
rect 6430 15850 6435 15870
rect 6405 15845 6435 15850
rect 6485 15870 6515 15875
rect 6485 15850 6490 15870
rect 6490 15850 6510 15870
rect 6510 15850 6515 15870
rect 6485 15845 6515 15850
rect 6565 15870 6595 15875
rect 6565 15850 6570 15870
rect 6570 15850 6590 15870
rect 6590 15850 6595 15870
rect 6565 15845 6595 15850
rect 6645 15870 6675 15875
rect 6645 15850 6650 15870
rect 6650 15850 6670 15870
rect 6670 15850 6675 15870
rect 6645 15845 6675 15850
rect 6725 15870 6755 15875
rect 6725 15850 6730 15870
rect 6730 15850 6750 15870
rect 6750 15850 6755 15870
rect 6725 15845 6755 15850
rect 6805 15870 6835 15875
rect 6805 15850 6810 15870
rect 6810 15850 6830 15870
rect 6830 15850 6835 15870
rect 6805 15845 6835 15850
rect 6885 15870 6915 15875
rect 6885 15850 6890 15870
rect 6890 15850 6910 15870
rect 6910 15850 6915 15870
rect 6885 15845 6915 15850
rect 6965 15870 6995 15875
rect 6965 15850 6970 15870
rect 6970 15850 6990 15870
rect 6990 15850 6995 15870
rect 6965 15845 6995 15850
rect 7045 15870 7075 15875
rect 7045 15850 7050 15870
rect 7050 15850 7070 15870
rect 7070 15850 7075 15870
rect 7045 15845 7075 15850
rect 7125 15870 7155 15875
rect 7125 15850 7130 15870
rect 7130 15850 7150 15870
rect 7150 15850 7155 15870
rect 7125 15845 7155 15850
rect 7205 15870 7235 15875
rect 7205 15850 7210 15870
rect 7210 15850 7230 15870
rect 7230 15850 7235 15870
rect 7205 15845 7235 15850
rect 7285 15870 7315 15875
rect 7285 15850 7290 15870
rect 7290 15850 7310 15870
rect 7310 15850 7315 15870
rect 7285 15845 7315 15850
rect 7365 15870 7395 15875
rect 7365 15850 7370 15870
rect 7370 15850 7390 15870
rect 7390 15850 7395 15870
rect 7365 15845 7395 15850
rect 7445 15870 7475 15875
rect 7445 15850 7450 15870
rect 7450 15850 7470 15870
rect 7470 15850 7475 15870
rect 7445 15845 7475 15850
rect 7525 15870 7555 15875
rect 7525 15850 7530 15870
rect 7530 15850 7550 15870
rect 7550 15850 7555 15870
rect 7525 15845 7555 15850
rect 7605 15870 7635 15875
rect 7605 15850 7610 15870
rect 7610 15850 7630 15870
rect 7630 15850 7635 15870
rect 7605 15845 7635 15850
rect 7685 15870 7715 15875
rect 7685 15850 7690 15870
rect 7690 15850 7710 15870
rect 7710 15850 7715 15870
rect 7685 15845 7715 15850
rect 7765 15870 7795 15875
rect 7765 15850 7770 15870
rect 7770 15850 7790 15870
rect 7790 15850 7795 15870
rect 7765 15845 7795 15850
rect 7845 15870 7875 15875
rect 7845 15850 7850 15870
rect 7850 15850 7870 15870
rect 7870 15850 7875 15870
rect 7845 15845 7875 15850
rect 7925 15870 7955 15875
rect 7925 15850 7930 15870
rect 7930 15850 7950 15870
rect 7950 15850 7955 15870
rect 7925 15845 7955 15850
rect 8005 15870 8035 15875
rect 8005 15850 8010 15870
rect 8010 15850 8030 15870
rect 8030 15850 8035 15870
rect 8005 15845 8035 15850
rect 8085 15870 8115 15875
rect 8085 15850 8090 15870
rect 8090 15850 8110 15870
rect 8110 15850 8115 15870
rect 8085 15845 8115 15850
rect 8165 15870 8195 15875
rect 8165 15850 8170 15870
rect 8170 15850 8190 15870
rect 8190 15850 8195 15870
rect 8165 15845 8195 15850
rect 8245 15870 8275 15875
rect 8245 15850 8250 15870
rect 8250 15850 8270 15870
rect 8270 15850 8275 15870
rect 8245 15845 8275 15850
rect 8325 15870 8355 15875
rect 8325 15850 8330 15870
rect 8330 15850 8350 15870
rect 8350 15850 8355 15870
rect 8325 15845 8355 15850
rect 8405 15870 8435 15875
rect 8405 15850 8410 15870
rect 8410 15850 8430 15870
rect 8430 15850 8435 15870
rect 8405 15845 8435 15850
rect 8485 15870 8515 15875
rect 8485 15850 8490 15870
rect 8490 15850 8510 15870
rect 8510 15850 8515 15870
rect 8485 15845 8515 15850
rect 8565 15870 8595 15875
rect 8565 15850 8570 15870
rect 8570 15850 8590 15870
rect 8590 15850 8595 15870
rect 8565 15845 8595 15850
rect 8645 15870 8675 15875
rect 8645 15850 8650 15870
rect 8650 15850 8670 15870
rect 8670 15850 8675 15870
rect 8645 15845 8675 15850
rect 8725 15870 8755 15875
rect 8725 15850 8730 15870
rect 8730 15850 8750 15870
rect 8750 15850 8755 15870
rect 8725 15845 8755 15850
rect 8805 15870 8835 15875
rect 8805 15850 8810 15870
rect 8810 15850 8830 15870
rect 8830 15850 8835 15870
rect 8805 15845 8835 15850
rect 8885 15870 8915 15875
rect 8885 15850 8890 15870
rect 8890 15850 8910 15870
rect 8910 15850 8915 15870
rect 8885 15845 8915 15850
rect 8965 15870 8995 15875
rect 8965 15850 8970 15870
rect 8970 15850 8990 15870
rect 8990 15850 8995 15870
rect 8965 15845 8995 15850
rect 9045 15870 9075 15875
rect 9045 15850 9050 15870
rect 9050 15850 9070 15870
rect 9070 15850 9075 15870
rect 9045 15845 9075 15850
rect 9125 15870 9155 15875
rect 9125 15850 9130 15870
rect 9130 15850 9150 15870
rect 9150 15850 9155 15870
rect 9125 15845 9155 15850
rect 9205 15870 9235 15875
rect 9205 15850 9210 15870
rect 9210 15850 9230 15870
rect 9230 15850 9235 15870
rect 9205 15845 9235 15850
rect 9285 15870 9315 15875
rect 9285 15850 9290 15870
rect 9290 15850 9310 15870
rect 9310 15850 9315 15870
rect 9285 15845 9315 15850
rect 9365 15870 9395 15875
rect 9365 15850 9370 15870
rect 9370 15850 9390 15870
rect 9390 15850 9395 15870
rect 9365 15845 9395 15850
rect 9445 15870 9475 15875
rect 9445 15850 9450 15870
rect 9450 15850 9470 15870
rect 9470 15850 9475 15870
rect 9445 15845 9475 15850
rect 11565 15870 11595 15875
rect 11565 15850 11570 15870
rect 11570 15850 11590 15870
rect 11590 15850 11595 15870
rect 11565 15845 11595 15850
rect 11645 15870 11675 15875
rect 11645 15850 11650 15870
rect 11650 15850 11670 15870
rect 11670 15850 11675 15870
rect 11645 15845 11675 15850
rect 11725 15870 11755 15875
rect 11725 15850 11730 15870
rect 11730 15850 11750 15870
rect 11750 15850 11755 15870
rect 11725 15845 11755 15850
rect 11805 15870 11835 15875
rect 11805 15850 11810 15870
rect 11810 15850 11830 15870
rect 11830 15850 11835 15870
rect 11805 15845 11835 15850
rect 11885 15870 11915 15875
rect 11885 15850 11890 15870
rect 11890 15850 11910 15870
rect 11910 15850 11915 15870
rect 11885 15845 11915 15850
rect 11965 15870 11995 15875
rect 11965 15850 11970 15870
rect 11970 15850 11990 15870
rect 11990 15850 11995 15870
rect 11965 15845 11995 15850
rect 12045 15870 12075 15875
rect 12045 15850 12050 15870
rect 12050 15850 12070 15870
rect 12070 15850 12075 15870
rect 12045 15845 12075 15850
rect 12125 15870 12155 15875
rect 12125 15850 12130 15870
rect 12130 15850 12150 15870
rect 12150 15850 12155 15870
rect 12125 15845 12155 15850
rect 12205 15870 12235 15875
rect 12205 15850 12210 15870
rect 12210 15850 12230 15870
rect 12230 15850 12235 15870
rect 12205 15845 12235 15850
rect 12285 15870 12315 15875
rect 12285 15850 12290 15870
rect 12290 15850 12310 15870
rect 12310 15850 12315 15870
rect 12285 15845 12315 15850
rect 12365 15870 12395 15875
rect 12365 15850 12370 15870
rect 12370 15850 12390 15870
rect 12390 15850 12395 15870
rect 12365 15845 12395 15850
rect 12445 15870 12475 15875
rect 12445 15850 12450 15870
rect 12450 15850 12470 15870
rect 12470 15850 12475 15870
rect 12445 15845 12475 15850
rect 12525 15870 12555 15875
rect 12525 15850 12530 15870
rect 12530 15850 12550 15870
rect 12550 15850 12555 15870
rect 12525 15845 12555 15850
rect 12605 15870 12635 15875
rect 12605 15850 12610 15870
rect 12610 15850 12630 15870
rect 12630 15850 12635 15870
rect 12605 15845 12635 15850
rect 12685 15870 12715 15875
rect 12685 15850 12690 15870
rect 12690 15850 12710 15870
rect 12710 15850 12715 15870
rect 12685 15845 12715 15850
rect 12765 15870 12795 15875
rect 12765 15850 12770 15870
rect 12770 15850 12790 15870
rect 12790 15850 12795 15870
rect 12765 15845 12795 15850
rect 12845 15870 12875 15875
rect 12845 15850 12850 15870
rect 12850 15850 12870 15870
rect 12870 15850 12875 15870
rect 12845 15845 12875 15850
rect 12925 15870 12955 15875
rect 12925 15850 12930 15870
rect 12930 15850 12950 15870
rect 12950 15850 12955 15870
rect 12925 15845 12955 15850
rect 13005 15870 13035 15875
rect 13005 15850 13010 15870
rect 13010 15850 13030 15870
rect 13030 15850 13035 15870
rect 13005 15845 13035 15850
rect 13085 15870 13115 15875
rect 13085 15850 13090 15870
rect 13090 15850 13110 15870
rect 13110 15850 13115 15870
rect 13085 15845 13115 15850
rect 13165 15870 13195 15875
rect 13165 15850 13170 15870
rect 13170 15850 13190 15870
rect 13190 15850 13195 15870
rect 13165 15845 13195 15850
rect 13245 15870 13275 15875
rect 13245 15850 13250 15870
rect 13250 15850 13270 15870
rect 13270 15850 13275 15870
rect 13245 15845 13275 15850
rect 13325 15870 13355 15875
rect 13325 15850 13330 15870
rect 13330 15850 13350 15870
rect 13350 15850 13355 15870
rect 13325 15845 13355 15850
rect 13405 15870 13435 15875
rect 13405 15850 13410 15870
rect 13410 15850 13430 15870
rect 13430 15850 13435 15870
rect 13405 15845 13435 15850
rect 13485 15870 13515 15875
rect 13485 15850 13490 15870
rect 13490 15850 13510 15870
rect 13510 15850 13515 15870
rect 13485 15845 13515 15850
rect 13565 15870 13595 15875
rect 13565 15850 13570 15870
rect 13570 15850 13590 15870
rect 13590 15850 13595 15870
rect 13565 15845 13595 15850
rect 13645 15870 13675 15875
rect 13645 15850 13650 15870
rect 13650 15850 13670 15870
rect 13670 15850 13675 15870
rect 13645 15845 13675 15850
rect 13725 15870 13755 15875
rect 13725 15850 13730 15870
rect 13730 15850 13750 15870
rect 13750 15850 13755 15870
rect 13725 15845 13755 15850
rect 13805 15870 13835 15875
rect 13805 15850 13810 15870
rect 13810 15850 13830 15870
rect 13830 15850 13835 15870
rect 13805 15845 13835 15850
rect 13885 15870 13915 15875
rect 13885 15850 13890 15870
rect 13890 15850 13910 15870
rect 13910 15850 13915 15870
rect 13885 15845 13915 15850
rect 13965 15870 13995 15875
rect 13965 15850 13970 15870
rect 13970 15850 13990 15870
rect 13990 15850 13995 15870
rect 13965 15845 13995 15850
rect 14045 15870 14075 15875
rect 14045 15850 14050 15870
rect 14050 15850 14070 15870
rect 14070 15850 14075 15870
rect 14045 15845 14075 15850
rect 14125 15870 14155 15875
rect 14125 15850 14130 15870
rect 14130 15850 14150 15870
rect 14150 15850 14155 15870
rect 14125 15845 14155 15850
rect 14205 15870 14235 15875
rect 14205 15850 14210 15870
rect 14210 15850 14230 15870
rect 14230 15850 14235 15870
rect 14205 15845 14235 15850
rect 14285 15870 14315 15875
rect 14285 15850 14290 15870
rect 14290 15850 14310 15870
rect 14310 15850 14315 15870
rect 14285 15845 14315 15850
rect 14365 15870 14395 15875
rect 14365 15850 14370 15870
rect 14370 15850 14390 15870
rect 14390 15850 14395 15870
rect 14365 15845 14395 15850
rect 14445 15870 14475 15875
rect 14445 15850 14450 15870
rect 14450 15850 14470 15870
rect 14470 15850 14475 15870
rect 14445 15845 14475 15850
rect 14525 15870 14555 15875
rect 14525 15850 14530 15870
rect 14530 15850 14550 15870
rect 14550 15850 14555 15870
rect 14525 15845 14555 15850
rect 14605 15870 14635 15875
rect 14605 15850 14610 15870
rect 14610 15850 14630 15870
rect 14630 15850 14635 15870
rect 14605 15845 14635 15850
rect 14685 15870 14715 15875
rect 14685 15850 14690 15870
rect 14690 15850 14710 15870
rect 14710 15850 14715 15870
rect 14685 15845 14715 15850
rect 16765 15870 16795 15875
rect 16765 15850 16770 15870
rect 16770 15850 16790 15870
rect 16790 15850 16795 15870
rect 16765 15845 16795 15850
rect 16845 15870 16875 15875
rect 16845 15850 16850 15870
rect 16850 15850 16870 15870
rect 16870 15850 16875 15870
rect 16845 15845 16875 15850
rect 16925 15870 16955 15875
rect 16925 15850 16930 15870
rect 16930 15850 16950 15870
rect 16950 15850 16955 15870
rect 16925 15845 16955 15850
rect 17005 15870 17035 15875
rect 17005 15850 17010 15870
rect 17010 15850 17030 15870
rect 17030 15850 17035 15870
rect 17005 15845 17035 15850
rect 17085 15870 17115 15875
rect 17085 15850 17090 15870
rect 17090 15850 17110 15870
rect 17110 15850 17115 15870
rect 17085 15845 17115 15850
rect 17165 15870 17195 15875
rect 17165 15850 17170 15870
rect 17170 15850 17190 15870
rect 17190 15850 17195 15870
rect 17165 15845 17195 15850
rect 17245 15870 17275 15875
rect 17245 15850 17250 15870
rect 17250 15850 17270 15870
rect 17270 15850 17275 15870
rect 17245 15845 17275 15850
rect 17325 15870 17355 15875
rect 17325 15850 17330 15870
rect 17330 15850 17350 15870
rect 17350 15850 17355 15870
rect 17325 15845 17355 15850
rect 17405 15870 17435 15875
rect 17405 15850 17410 15870
rect 17410 15850 17430 15870
rect 17430 15850 17435 15870
rect 17405 15845 17435 15850
rect 17485 15870 17515 15875
rect 17485 15850 17490 15870
rect 17490 15850 17510 15870
rect 17510 15850 17515 15870
rect 17485 15845 17515 15850
rect 17565 15870 17595 15875
rect 17565 15850 17570 15870
rect 17570 15850 17590 15870
rect 17590 15850 17595 15870
rect 17565 15845 17595 15850
rect 17645 15870 17675 15875
rect 17645 15850 17650 15870
rect 17650 15850 17670 15870
rect 17670 15850 17675 15870
rect 17645 15845 17675 15850
rect 17725 15870 17755 15875
rect 17725 15850 17730 15870
rect 17730 15850 17750 15870
rect 17750 15850 17755 15870
rect 17725 15845 17755 15850
rect 17805 15870 17835 15875
rect 17805 15850 17810 15870
rect 17810 15850 17830 15870
rect 17830 15850 17835 15870
rect 17805 15845 17835 15850
rect 17885 15870 17915 15875
rect 17885 15850 17890 15870
rect 17890 15850 17910 15870
rect 17910 15850 17915 15870
rect 17885 15845 17915 15850
rect 17965 15870 17995 15875
rect 17965 15850 17970 15870
rect 17970 15850 17990 15870
rect 17990 15850 17995 15870
rect 17965 15845 17995 15850
rect 18045 15870 18075 15875
rect 18045 15850 18050 15870
rect 18050 15850 18070 15870
rect 18070 15850 18075 15870
rect 18045 15845 18075 15850
rect 18125 15870 18155 15875
rect 18125 15850 18130 15870
rect 18130 15850 18150 15870
rect 18150 15850 18155 15870
rect 18125 15845 18155 15850
rect 18205 15870 18235 15875
rect 18205 15850 18210 15870
rect 18210 15850 18230 15870
rect 18230 15850 18235 15870
rect 18205 15845 18235 15850
rect 18285 15870 18315 15875
rect 18285 15850 18290 15870
rect 18290 15850 18310 15870
rect 18310 15850 18315 15870
rect 18285 15845 18315 15850
rect 18365 15870 18395 15875
rect 18365 15850 18370 15870
rect 18370 15850 18390 15870
rect 18390 15850 18395 15870
rect 18365 15845 18395 15850
rect 18445 15870 18475 15875
rect 18445 15850 18450 15870
rect 18450 15850 18470 15870
rect 18470 15850 18475 15870
rect 18445 15845 18475 15850
rect 18525 15870 18555 15875
rect 18525 15850 18530 15870
rect 18530 15850 18550 15870
rect 18550 15850 18555 15870
rect 18525 15845 18555 15850
rect 18605 15870 18635 15875
rect 18605 15850 18610 15870
rect 18610 15850 18630 15870
rect 18630 15850 18635 15870
rect 18605 15845 18635 15850
rect 18685 15870 18715 15875
rect 18685 15850 18690 15870
rect 18690 15850 18710 15870
rect 18710 15850 18715 15870
rect 18685 15845 18715 15850
rect 18765 15870 18795 15875
rect 18765 15850 18770 15870
rect 18770 15850 18790 15870
rect 18790 15850 18795 15870
rect 18765 15845 18795 15850
rect 18845 15870 18875 15875
rect 18845 15850 18850 15870
rect 18850 15850 18870 15870
rect 18870 15850 18875 15870
rect 18845 15845 18875 15850
rect 18925 15870 18955 15875
rect 18925 15850 18930 15870
rect 18930 15850 18950 15870
rect 18950 15850 18955 15870
rect 18925 15845 18955 15850
rect 19005 15870 19035 15875
rect 19005 15850 19010 15870
rect 19010 15850 19030 15870
rect 19030 15850 19035 15870
rect 19005 15845 19035 15850
rect 19085 15870 19115 15875
rect 19085 15850 19090 15870
rect 19090 15850 19110 15870
rect 19110 15850 19115 15870
rect 19085 15845 19115 15850
rect 19165 15870 19195 15875
rect 19165 15850 19170 15870
rect 19170 15850 19190 15870
rect 19190 15850 19195 15870
rect 19165 15845 19195 15850
rect 19245 15870 19275 15875
rect 19245 15850 19250 15870
rect 19250 15850 19270 15870
rect 19270 15850 19275 15870
rect 19245 15845 19275 15850
rect 19325 15870 19355 15875
rect 19325 15850 19330 15870
rect 19330 15850 19350 15870
rect 19350 15850 19355 15870
rect 19325 15845 19355 15850
rect 19405 15870 19435 15875
rect 19405 15850 19410 15870
rect 19410 15850 19430 15870
rect 19430 15850 19435 15870
rect 19405 15845 19435 15850
rect 19485 15870 19515 15875
rect 19485 15850 19490 15870
rect 19490 15850 19510 15870
rect 19510 15850 19515 15870
rect 19485 15845 19515 15850
rect 19565 15870 19595 15875
rect 19565 15850 19570 15870
rect 19570 15850 19590 15870
rect 19590 15850 19595 15870
rect 19565 15845 19595 15850
rect 19645 15870 19675 15875
rect 19645 15850 19650 15870
rect 19650 15850 19670 15870
rect 19670 15850 19675 15870
rect 19645 15845 19675 15850
rect 19725 15870 19755 15875
rect 19725 15850 19730 15870
rect 19730 15850 19750 15870
rect 19750 15850 19755 15870
rect 19725 15845 19755 15850
rect 19805 15870 19835 15875
rect 19805 15850 19810 15870
rect 19810 15850 19830 15870
rect 19830 15850 19835 15870
rect 19805 15845 19835 15850
rect 19885 15870 19915 15875
rect 19885 15850 19890 15870
rect 19890 15850 19910 15870
rect 19910 15850 19915 15870
rect 19885 15845 19915 15850
rect 19965 15870 19995 15875
rect 19965 15850 19970 15870
rect 19970 15850 19990 15870
rect 19990 15850 19995 15870
rect 19965 15845 19995 15850
rect 20045 15870 20075 15875
rect 20045 15850 20050 15870
rect 20050 15850 20070 15870
rect 20070 15850 20075 15870
rect 20045 15845 20075 15850
rect 20125 15870 20155 15875
rect 20125 15850 20130 15870
rect 20130 15850 20150 15870
rect 20150 15850 20155 15870
rect 20125 15845 20155 15850
rect 20205 15870 20235 15875
rect 20205 15850 20210 15870
rect 20210 15850 20230 15870
rect 20230 15850 20235 15870
rect 20205 15845 20235 15850
rect 20285 15870 20315 15875
rect 20285 15850 20290 15870
rect 20290 15850 20310 15870
rect 20310 15850 20315 15870
rect 20285 15845 20315 15850
rect 20365 15870 20395 15875
rect 20365 15850 20370 15870
rect 20370 15850 20390 15870
rect 20390 15850 20395 15870
rect 20365 15845 20395 15850
rect 20445 15870 20475 15875
rect 20445 15850 20450 15870
rect 20450 15850 20470 15870
rect 20470 15850 20475 15870
rect 20445 15845 20475 15850
rect 20525 15870 20555 15875
rect 20525 15850 20530 15870
rect 20530 15850 20550 15870
rect 20550 15850 20555 15870
rect 20525 15845 20555 15850
rect 20605 15870 20635 15875
rect 20605 15850 20610 15870
rect 20610 15850 20630 15870
rect 20630 15850 20635 15870
rect 20605 15845 20635 15850
rect 20685 15870 20715 15875
rect 20685 15850 20690 15870
rect 20690 15850 20710 15870
rect 20710 15850 20715 15870
rect 20685 15845 20715 15850
rect 20765 15870 20795 15875
rect 20765 15850 20770 15870
rect 20770 15850 20790 15870
rect 20790 15850 20795 15870
rect 20765 15845 20795 15850
rect 20845 15870 20875 15875
rect 20845 15850 20850 15870
rect 20850 15850 20870 15870
rect 20870 15850 20875 15870
rect 20845 15845 20875 15850
rect 20925 15870 20955 15875
rect 20925 15850 20930 15870
rect 20930 15850 20950 15870
rect 20950 15850 20955 15870
rect 20925 15845 20955 15850
rect 5 15710 35 15715
rect 5 15690 10 15710
rect 10 15690 30 15710
rect 30 15690 35 15710
rect 5 15685 35 15690
rect 85 15710 115 15715
rect 85 15690 90 15710
rect 90 15690 110 15710
rect 110 15690 115 15710
rect 85 15685 115 15690
rect 165 15710 195 15715
rect 165 15690 170 15710
rect 170 15690 190 15710
rect 190 15690 195 15710
rect 165 15685 195 15690
rect 245 15710 275 15715
rect 245 15690 250 15710
rect 250 15690 270 15710
rect 270 15690 275 15710
rect 245 15685 275 15690
rect 325 15710 355 15715
rect 325 15690 330 15710
rect 330 15690 350 15710
rect 350 15690 355 15710
rect 325 15685 355 15690
rect 405 15710 435 15715
rect 405 15690 410 15710
rect 410 15690 430 15710
rect 430 15690 435 15710
rect 405 15685 435 15690
rect 485 15710 515 15715
rect 485 15690 490 15710
rect 490 15690 510 15710
rect 510 15690 515 15710
rect 485 15685 515 15690
rect 565 15710 595 15715
rect 565 15690 570 15710
rect 570 15690 590 15710
rect 590 15690 595 15710
rect 565 15685 595 15690
rect 645 15710 675 15715
rect 645 15690 650 15710
rect 650 15690 670 15710
rect 670 15690 675 15710
rect 645 15685 675 15690
rect 725 15710 755 15715
rect 725 15690 730 15710
rect 730 15690 750 15710
rect 750 15690 755 15710
rect 725 15685 755 15690
rect 805 15710 835 15715
rect 805 15690 810 15710
rect 810 15690 830 15710
rect 830 15690 835 15710
rect 805 15685 835 15690
rect 885 15710 915 15715
rect 885 15690 890 15710
rect 890 15690 910 15710
rect 910 15690 915 15710
rect 885 15685 915 15690
rect 965 15710 995 15715
rect 965 15690 970 15710
rect 970 15690 990 15710
rect 990 15690 995 15710
rect 965 15685 995 15690
rect 1045 15710 1075 15715
rect 1045 15690 1050 15710
rect 1050 15690 1070 15710
rect 1070 15690 1075 15710
rect 1045 15685 1075 15690
rect 1125 15710 1155 15715
rect 1125 15690 1130 15710
rect 1130 15690 1150 15710
rect 1150 15690 1155 15710
rect 1125 15685 1155 15690
rect 1205 15710 1235 15715
rect 1205 15690 1210 15710
rect 1210 15690 1230 15710
rect 1230 15690 1235 15710
rect 1205 15685 1235 15690
rect 1285 15710 1315 15715
rect 1285 15690 1290 15710
rect 1290 15690 1310 15710
rect 1310 15690 1315 15710
rect 1285 15685 1315 15690
rect 1365 15710 1395 15715
rect 1365 15690 1370 15710
rect 1370 15690 1390 15710
rect 1390 15690 1395 15710
rect 1365 15685 1395 15690
rect 1445 15710 1475 15715
rect 1445 15690 1450 15710
rect 1450 15690 1470 15710
rect 1470 15690 1475 15710
rect 1445 15685 1475 15690
rect 1525 15710 1555 15715
rect 1525 15690 1530 15710
rect 1530 15690 1550 15710
rect 1550 15690 1555 15710
rect 1525 15685 1555 15690
rect 1605 15710 1635 15715
rect 1605 15690 1610 15710
rect 1610 15690 1630 15710
rect 1630 15690 1635 15710
rect 1605 15685 1635 15690
rect 1685 15710 1715 15715
rect 1685 15690 1690 15710
rect 1690 15690 1710 15710
rect 1710 15690 1715 15710
rect 1685 15685 1715 15690
rect 1765 15710 1795 15715
rect 1765 15690 1770 15710
rect 1770 15690 1790 15710
rect 1790 15690 1795 15710
rect 1765 15685 1795 15690
rect 1845 15710 1875 15715
rect 1845 15690 1850 15710
rect 1850 15690 1870 15710
rect 1870 15690 1875 15710
rect 1845 15685 1875 15690
rect 1925 15710 1955 15715
rect 1925 15690 1930 15710
rect 1930 15690 1950 15710
rect 1950 15690 1955 15710
rect 1925 15685 1955 15690
rect 2005 15710 2035 15715
rect 2005 15690 2010 15710
rect 2010 15690 2030 15710
rect 2030 15690 2035 15710
rect 2005 15685 2035 15690
rect 2085 15710 2115 15715
rect 2085 15690 2090 15710
rect 2090 15690 2110 15710
rect 2110 15690 2115 15710
rect 2085 15685 2115 15690
rect 2165 15710 2195 15715
rect 2165 15690 2170 15710
rect 2170 15690 2190 15710
rect 2190 15690 2195 15710
rect 2165 15685 2195 15690
rect 2245 15710 2275 15715
rect 2245 15690 2250 15710
rect 2250 15690 2270 15710
rect 2270 15690 2275 15710
rect 2245 15685 2275 15690
rect 2325 15710 2355 15715
rect 2325 15690 2330 15710
rect 2330 15690 2350 15710
rect 2350 15690 2355 15710
rect 2325 15685 2355 15690
rect 2405 15710 2435 15715
rect 2405 15690 2410 15710
rect 2410 15690 2430 15710
rect 2430 15690 2435 15710
rect 2405 15685 2435 15690
rect 2485 15710 2515 15715
rect 2485 15690 2490 15710
rect 2490 15690 2510 15710
rect 2510 15690 2515 15710
rect 2485 15685 2515 15690
rect 2565 15710 2595 15715
rect 2565 15690 2570 15710
rect 2570 15690 2590 15710
rect 2590 15690 2595 15710
rect 2565 15685 2595 15690
rect 2645 15710 2675 15715
rect 2645 15690 2650 15710
rect 2650 15690 2670 15710
rect 2670 15690 2675 15710
rect 2645 15685 2675 15690
rect 2725 15710 2755 15715
rect 2725 15690 2730 15710
rect 2730 15690 2750 15710
rect 2750 15690 2755 15710
rect 2725 15685 2755 15690
rect 2805 15710 2835 15715
rect 2805 15690 2810 15710
rect 2810 15690 2830 15710
rect 2830 15690 2835 15710
rect 2805 15685 2835 15690
rect 2885 15710 2915 15715
rect 2885 15690 2890 15710
rect 2890 15690 2910 15710
rect 2910 15690 2915 15710
rect 2885 15685 2915 15690
rect 2965 15710 2995 15715
rect 2965 15690 2970 15710
rect 2970 15690 2990 15710
rect 2990 15690 2995 15710
rect 2965 15685 2995 15690
rect 3045 15710 3075 15715
rect 3045 15690 3050 15710
rect 3050 15690 3070 15710
rect 3070 15690 3075 15710
rect 3045 15685 3075 15690
rect 3125 15710 3155 15715
rect 3125 15690 3130 15710
rect 3130 15690 3150 15710
rect 3150 15690 3155 15710
rect 3125 15685 3155 15690
rect 3205 15710 3235 15715
rect 3205 15690 3210 15710
rect 3210 15690 3230 15710
rect 3230 15690 3235 15710
rect 3205 15685 3235 15690
rect 3285 15710 3315 15715
rect 3285 15690 3290 15710
rect 3290 15690 3310 15710
rect 3310 15690 3315 15710
rect 3285 15685 3315 15690
rect 3365 15710 3395 15715
rect 3365 15690 3370 15710
rect 3370 15690 3390 15710
rect 3390 15690 3395 15710
rect 3365 15685 3395 15690
rect 3445 15710 3475 15715
rect 3445 15690 3450 15710
rect 3450 15690 3470 15710
rect 3470 15690 3475 15710
rect 3445 15685 3475 15690
rect 3525 15710 3555 15715
rect 3525 15690 3530 15710
rect 3530 15690 3550 15710
rect 3550 15690 3555 15710
rect 3525 15685 3555 15690
rect 3605 15710 3635 15715
rect 3605 15690 3610 15710
rect 3610 15690 3630 15710
rect 3630 15690 3635 15710
rect 3605 15685 3635 15690
rect 3685 15710 3715 15715
rect 3685 15690 3690 15710
rect 3690 15690 3710 15710
rect 3710 15690 3715 15710
rect 3685 15685 3715 15690
rect 3765 15710 3795 15715
rect 3765 15690 3770 15710
rect 3770 15690 3790 15710
rect 3790 15690 3795 15710
rect 3765 15685 3795 15690
rect 3845 15710 3875 15715
rect 3845 15690 3850 15710
rect 3850 15690 3870 15710
rect 3870 15690 3875 15710
rect 3845 15685 3875 15690
rect 3925 15710 3955 15715
rect 3925 15690 3930 15710
rect 3930 15690 3950 15710
rect 3950 15690 3955 15710
rect 3925 15685 3955 15690
rect 4005 15710 4035 15715
rect 4005 15690 4010 15710
rect 4010 15690 4030 15710
rect 4030 15690 4035 15710
rect 4005 15685 4035 15690
rect 4085 15710 4115 15715
rect 4085 15690 4090 15710
rect 4090 15690 4110 15710
rect 4110 15690 4115 15710
rect 4085 15685 4115 15690
rect 4165 15710 4195 15715
rect 4165 15690 4170 15710
rect 4170 15690 4190 15710
rect 4190 15690 4195 15710
rect 4165 15685 4195 15690
rect 6245 15710 6275 15715
rect 6245 15690 6250 15710
rect 6250 15690 6270 15710
rect 6270 15690 6275 15710
rect 6245 15685 6275 15690
rect 6325 15710 6355 15715
rect 6325 15690 6330 15710
rect 6330 15690 6350 15710
rect 6350 15690 6355 15710
rect 6325 15685 6355 15690
rect 6405 15710 6435 15715
rect 6405 15690 6410 15710
rect 6410 15690 6430 15710
rect 6430 15690 6435 15710
rect 6405 15685 6435 15690
rect 6485 15710 6515 15715
rect 6485 15690 6490 15710
rect 6490 15690 6510 15710
rect 6510 15690 6515 15710
rect 6485 15685 6515 15690
rect 6565 15710 6595 15715
rect 6565 15690 6570 15710
rect 6570 15690 6590 15710
rect 6590 15690 6595 15710
rect 6565 15685 6595 15690
rect 6645 15710 6675 15715
rect 6645 15690 6650 15710
rect 6650 15690 6670 15710
rect 6670 15690 6675 15710
rect 6645 15685 6675 15690
rect 6725 15710 6755 15715
rect 6725 15690 6730 15710
rect 6730 15690 6750 15710
rect 6750 15690 6755 15710
rect 6725 15685 6755 15690
rect 6805 15710 6835 15715
rect 6805 15690 6810 15710
rect 6810 15690 6830 15710
rect 6830 15690 6835 15710
rect 6805 15685 6835 15690
rect 6885 15710 6915 15715
rect 6885 15690 6890 15710
rect 6890 15690 6910 15710
rect 6910 15690 6915 15710
rect 6885 15685 6915 15690
rect 6965 15710 6995 15715
rect 6965 15690 6970 15710
rect 6970 15690 6990 15710
rect 6990 15690 6995 15710
rect 6965 15685 6995 15690
rect 7045 15710 7075 15715
rect 7045 15690 7050 15710
rect 7050 15690 7070 15710
rect 7070 15690 7075 15710
rect 7045 15685 7075 15690
rect 7125 15710 7155 15715
rect 7125 15690 7130 15710
rect 7130 15690 7150 15710
rect 7150 15690 7155 15710
rect 7125 15685 7155 15690
rect 7205 15710 7235 15715
rect 7205 15690 7210 15710
rect 7210 15690 7230 15710
rect 7230 15690 7235 15710
rect 7205 15685 7235 15690
rect 7285 15710 7315 15715
rect 7285 15690 7290 15710
rect 7290 15690 7310 15710
rect 7310 15690 7315 15710
rect 7285 15685 7315 15690
rect 7365 15710 7395 15715
rect 7365 15690 7370 15710
rect 7370 15690 7390 15710
rect 7390 15690 7395 15710
rect 7365 15685 7395 15690
rect 7445 15710 7475 15715
rect 7445 15690 7450 15710
rect 7450 15690 7470 15710
rect 7470 15690 7475 15710
rect 7445 15685 7475 15690
rect 7525 15710 7555 15715
rect 7525 15690 7530 15710
rect 7530 15690 7550 15710
rect 7550 15690 7555 15710
rect 7525 15685 7555 15690
rect 7605 15710 7635 15715
rect 7605 15690 7610 15710
rect 7610 15690 7630 15710
rect 7630 15690 7635 15710
rect 7605 15685 7635 15690
rect 7685 15710 7715 15715
rect 7685 15690 7690 15710
rect 7690 15690 7710 15710
rect 7710 15690 7715 15710
rect 7685 15685 7715 15690
rect 7765 15710 7795 15715
rect 7765 15690 7770 15710
rect 7770 15690 7790 15710
rect 7790 15690 7795 15710
rect 7765 15685 7795 15690
rect 7845 15710 7875 15715
rect 7845 15690 7850 15710
rect 7850 15690 7870 15710
rect 7870 15690 7875 15710
rect 7845 15685 7875 15690
rect 7925 15710 7955 15715
rect 7925 15690 7930 15710
rect 7930 15690 7950 15710
rect 7950 15690 7955 15710
rect 7925 15685 7955 15690
rect 8005 15710 8035 15715
rect 8005 15690 8010 15710
rect 8010 15690 8030 15710
rect 8030 15690 8035 15710
rect 8005 15685 8035 15690
rect 8085 15710 8115 15715
rect 8085 15690 8090 15710
rect 8090 15690 8110 15710
rect 8110 15690 8115 15710
rect 8085 15685 8115 15690
rect 8165 15710 8195 15715
rect 8165 15690 8170 15710
rect 8170 15690 8190 15710
rect 8190 15690 8195 15710
rect 8165 15685 8195 15690
rect 8245 15710 8275 15715
rect 8245 15690 8250 15710
rect 8250 15690 8270 15710
rect 8270 15690 8275 15710
rect 8245 15685 8275 15690
rect 8325 15710 8355 15715
rect 8325 15690 8330 15710
rect 8330 15690 8350 15710
rect 8350 15690 8355 15710
rect 8325 15685 8355 15690
rect 8405 15710 8435 15715
rect 8405 15690 8410 15710
rect 8410 15690 8430 15710
rect 8430 15690 8435 15710
rect 8405 15685 8435 15690
rect 8485 15710 8515 15715
rect 8485 15690 8490 15710
rect 8490 15690 8510 15710
rect 8510 15690 8515 15710
rect 8485 15685 8515 15690
rect 8565 15710 8595 15715
rect 8565 15690 8570 15710
rect 8570 15690 8590 15710
rect 8590 15690 8595 15710
rect 8565 15685 8595 15690
rect 8645 15710 8675 15715
rect 8645 15690 8650 15710
rect 8650 15690 8670 15710
rect 8670 15690 8675 15710
rect 8645 15685 8675 15690
rect 8725 15710 8755 15715
rect 8725 15690 8730 15710
rect 8730 15690 8750 15710
rect 8750 15690 8755 15710
rect 8725 15685 8755 15690
rect 8805 15710 8835 15715
rect 8805 15690 8810 15710
rect 8810 15690 8830 15710
rect 8830 15690 8835 15710
rect 8805 15685 8835 15690
rect 8885 15710 8915 15715
rect 8885 15690 8890 15710
rect 8890 15690 8910 15710
rect 8910 15690 8915 15710
rect 8885 15685 8915 15690
rect 8965 15710 8995 15715
rect 8965 15690 8970 15710
rect 8970 15690 8990 15710
rect 8990 15690 8995 15710
rect 8965 15685 8995 15690
rect 9045 15710 9075 15715
rect 9045 15690 9050 15710
rect 9050 15690 9070 15710
rect 9070 15690 9075 15710
rect 9045 15685 9075 15690
rect 9125 15710 9155 15715
rect 9125 15690 9130 15710
rect 9130 15690 9150 15710
rect 9150 15690 9155 15710
rect 9125 15685 9155 15690
rect 9205 15710 9235 15715
rect 9205 15690 9210 15710
rect 9210 15690 9230 15710
rect 9230 15690 9235 15710
rect 9205 15685 9235 15690
rect 9285 15710 9315 15715
rect 9285 15690 9290 15710
rect 9290 15690 9310 15710
rect 9310 15690 9315 15710
rect 9285 15685 9315 15690
rect 9365 15710 9395 15715
rect 9365 15690 9370 15710
rect 9370 15690 9390 15710
rect 9390 15690 9395 15710
rect 9365 15685 9395 15690
rect 9445 15710 9475 15715
rect 9445 15690 9450 15710
rect 9450 15690 9470 15710
rect 9470 15690 9475 15710
rect 9445 15685 9475 15690
rect 11565 15710 11595 15715
rect 11565 15690 11570 15710
rect 11570 15690 11590 15710
rect 11590 15690 11595 15710
rect 11565 15685 11595 15690
rect 11645 15710 11675 15715
rect 11645 15690 11650 15710
rect 11650 15690 11670 15710
rect 11670 15690 11675 15710
rect 11645 15685 11675 15690
rect 11725 15710 11755 15715
rect 11725 15690 11730 15710
rect 11730 15690 11750 15710
rect 11750 15690 11755 15710
rect 11725 15685 11755 15690
rect 11805 15710 11835 15715
rect 11805 15690 11810 15710
rect 11810 15690 11830 15710
rect 11830 15690 11835 15710
rect 11805 15685 11835 15690
rect 11885 15710 11915 15715
rect 11885 15690 11890 15710
rect 11890 15690 11910 15710
rect 11910 15690 11915 15710
rect 11885 15685 11915 15690
rect 11965 15710 11995 15715
rect 11965 15690 11970 15710
rect 11970 15690 11990 15710
rect 11990 15690 11995 15710
rect 11965 15685 11995 15690
rect 12045 15710 12075 15715
rect 12045 15690 12050 15710
rect 12050 15690 12070 15710
rect 12070 15690 12075 15710
rect 12045 15685 12075 15690
rect 12125 15710 12155 15715
rect 12125 15690 12130 15710
rect 12130 15690 12150 15710
rect 12150 15690 12155 15710
rect 12125 15685 12155 15690
rect 12205 15710 12235 15715
rect 12205 15690 12210 15710
rect 12210 15690 12230 15710
rect 12230 15690 12235 15710
rect 12205 15685 12235 15690
rect 12285 15710 12315 15715
rect 12285 15690 12290 15710
rect 12290 15690 12310 15710
rect 12310 15690 12315 15710
rect 12285 15685 12315 15690
rect 12365 15710 12395 15715
rect 12365 15690 12370 15710
rect 12370 15690 12390 15710
rect 12390 15690 12395 15710
rect 12365 15685 12395 15690
rect 12445 15710 12475 15715
rect 12445 15690 12450 15710
rect 12450 15690 12470 15710
rect 12470 15690 12475 15710
rect 12445 15685 12475 15690
rect 12525 15710 12555 15715
rect 12525 15690 12530 15710
rect 12530 15690 12550 15710
rect 12550 15690 12555 15710
rect 12525 15685 12555 15690
rect 12605 15710 12635 15715
rect 12605 15690 12610 15710
rect 12610 15690 12630 15710
rect 12630 15690 12635 15710
rect 12605 15685 12635 15690
rect 12685 15710 12715 15715
rect 12685 15690 12690 15710
rect 12690 15690 12710 15710
rect 12710 15690 12715 15710
rect 12685 15685 12715 15690
rect 12765 15710 12795 15715
rect 12765 15690 12770 15710
rect 12770 15690 12790 15710
rect 12790 15690 12795 15710
rect 12765 15685 12795 15690
rect 12845 15710 12875 15715
rect 12845 15690 12850 15710
rect 12850 15690 12870 15710
rect 12870 15690 12875 15710
rect 12845 15685 12875 15690
rect 12925 15710 12955 15715
rect 12925 15690 12930 15710
rect 12930 15690 12950 15710
rect 12950 15690 12955 15710
rect 12925 15685 12955 15690
rect 13005 15710 13035 15715
rect 13005 15690 13010 15710
rect 13010 15690 13030 15710
rect 13030 15690 13035 15710
rect 13005 15685 13035 15690
rect 13085 15710 13115 15715
rect 13085 15690 13090 15710
rect 13090 15690 13110 15710
rect 13110 15690 13115 15710
rect 13085 15685 13115 15690
rect 13165 15710 13195 15715
rect 13165 15690 13170 15710
rect 13170 15690 13190 15710
rect 13190 15690 13195 15710
rect 13165 15685 13195 15690
rect 13245 15710 13275 15715
rect 13245 15690 13250 15710
rect 13250 15690 13270 15710
rect 13270 15690 13275 15710
rect 13245 15685 13275 15690
rect 13325 15710 13355 15715
rect 13325 15690 13330 15710
rect 13330 15690 13350 15710
rect 13350 15690 13355 15710
rect 13325 15685 13355 15690
rect 13405 15710 13435 15715
rect 13405 15690 13410 15710
rect 13410 15690 13430 15710
rect 13430 15690 13435 15710
rect 13405 15685 13435 15690
rect 13485 15710 13515 15715
rect 13485 15690 13490 15710
rect 13490 15690 13510 15710
rect 13510 15690 13515 15710
rect 13485 15685 13515 15690
rect 13565 15710 13595 15715
rect 13565 15690 13570 15710
rect 13570 15690 13590 15710
rect 13590 15690 13595 15710
rect 13565 15685 13595 15690
rect 13645 15710 13675 15715
rect 13645 15690 13650 15710
rect 13650 15690 13670 15710
rect 13670 15690 13675 15710
rect 13645 15685 13675 15690
rect 13725 15710 13755 15715
rect 13725 15690 13730 15710
rect 13730 15690 13750 15710
rect 13750 15690 13755 15710
rect 13725 15685 13755 15690
rect 13805 15710 13835 15715
rect 13805 15690 13810 15710
rect 13810 15690 13830 15710
rect 13830 15690 13835 15710
rect 13805 15685 13835 15690
rect 13885 15710 13915 15715
rect 13885 15690 13890 15710
rect 13890 15690 13910 15710
rect 13910 15690 13915 15710
rect 13885 15685 13915 15690
rect 13965 15710 13995 15715
rect 13965 15690 13970 15710
rect 13970 15690 13990 15710
rect 13990 15690 13995 15710
rect 13965 15685 13995 15690
rect 14045 15710 14075 15715
rect 14045 15690 14050 15710
rect 14050 15690 14070 15710
rect 14070 15690 14075 15710
rect 14045 15685 14075 15690
rect 14125 15710 14155 15715
rect 14125 15690 14130 15710
rect 14130 15690 14150 15710
rect 14150 15690 14155 15710
rect 14125 15685 14155 15690
rect 14205 15710 14235 15715
rect 14205 15690 14210 15710
rect 14210 15690 14230 15710
rect 14230 15690 14235 15710
rect 14205 15685 14235 15690
rect 14285 15710 14315 15715
rect 14285 15690 14290 15710
rect 14290 15690 14310 15710
rect 14310 15690 14315 15710
rect 14285 15685 14315 15690
rect 14365 15710 14395 15715
rect 14365 15690 14370 15710
rect 14370 15690 14390 15710
rect 14390 15690 14395 15710
rect 14365 15685 14395 15690
rect 14445 15710 14475 15715
rect 14445 15690 14450 15710
rect 14450 15690 14470 15710
rect 14470 15690 14475 15710
rect 14445 15685 14475 15690
rect 14525 15710 14555 15715
rect 14525 15690 14530 15710
rect 14530 15690 14550 15710
rect 14550 15690 14555 15710
rect 14525 15685 14555 15690
rect 14605 15710 14635 15715
rect 14605 15690 14610 15710
rect 14610 15690 14630 15710
rect 14630 15690 14635 15710
rect 14605 15685 14635 15690
rect 14685 15710 14715 15715
rect 14685 15690 14690 15710
rect 14690 15690 14710 15710
rect 14710 15690 14715 15710
rect 14685 15685 14715 15690
rect 16765 15710 16795 15715
rect 16765 15690 16770 15710
rect 16770 15690 16790 15710
rect 16790 15690 16795 15710
rect 16765 15685 16795 15690
rect 16845 15710 16875 15715
rect 16845 15690 16850 15710
rect 16850 15690 16870 15710
rect 16870 15690 16875 15710
rect 16845 15685 16875 15690
rect 16925 15710 16955 15715
rect 16925 15690 16930 15710
rect 16930 15690 16950 15710
rect 16950 15690 16955 15710
rect 16925 15685 16955 15690
rect 17005 15710 17035 15715
rect 17005 15690 17010 15710
rect 17010 15690 17030 15710
rect 17030 15690 17035 15710
rect 17005 15685 17035 15690
rect 17085 15710 17115 15715
rect 17085 15690 17090 15710
rect 17090 15690 17110 15710
rect 17110 15690 17115 15710
rect 17085 15685 17115 15690
rect 17165 15710 17195 15715
rect 17165 15690 17170 15710
rect 17170 15690 17190 15710
rect 17190 15690 17195 15710
rect 17165 15685 17195 15690
rect 17245 15710 17275 15715
rect 17245 15690 17250 15710
rect 17250 15690 17270 15710
rect 17270 15690 17275 15710
rect 17245 15685 17275 15690
rect 17325 15710 17355 15715
rect 17325 15690 17330 15710
rect 17330 15690 17350 15710
rect 17350 15690 17355 15710
rect 17325 15685 17355 15690
rect 17405 15710 17435 15715
rect 17405 15690 17410 15710
rect 17410 15690 17430 15710
rect 17430 15690 17435 15710
rect 17405 15685 17435 15690
rect 17485 15710 17515 15715
rect 17485 15690 17490 15710
rect 17490 15690 17510 15710
rect 17510 15690 17515 15710
rect 17485 15685 17515 15690
rect 17565 15710 17595 15715
rect 17565 15690 17570 15710
rect 17570 15690 17590 15710
rect 17590 15690 17595 15710
rect 17565 15685 17595 15690
rect 17645 15710 17675 15715
rect 17645 15690 17650 15710
rect 17650 15690 17670 15710
rect 17670 15690 17675 15710
rect 17645 15685 17675 15690
rect 17725 15710 17755 15715
rect 17725 15690 17730 15710
rect 17730 15690 17750 15710
rect 17750 15690 17755 15710
rect 17725 15685 17755 15690
rect 17805 15710 17835 15715
rect 17805 15690 17810 15710
rect 17810 15690 17830 15710
rect 17830 15690 17835 15710
rect 17805 15685 17835 15690
rect 17885 15710 17915 15715
rect 17885 15690 17890 15710
rect 17890 15690 17910 15710
rect 17910 15690 17915 15710
rect 17885 15685 17915 15690
rect 17965 15710 17995 15715
rect 17965 15690 17970 15710
rect 17970 15690 17990 15710
rect 17990 15690 17995 15710
rect 17965 15685 17995 15690
rect 18045 15710 18075 15715
rect 18045 15690 18050 15710
rect 18050 15690 18070 15710
rect 18070 15690 18075 15710
rect 18045 15685 18075 15690
rect 18125 15710 18155 15715
rect 18125 15690 18130 15710
rect 18130 15690 18150 15710
rect 18150 15690 18155 15710
rect 18125 15685 18155 15690
rect 18205 15710 18235 15715
rect 18205 15690 18210 15710
rect 18210 15690 18230 15710
rect 18230 15690 18235 15710
rect 18205 15685 18235 15690
rect 18285 15710 18315 15715
rect 18285 15690 18290 15710
rect 18290 15690 18310 15710
rect 18310 15690 18315 15710
rect 18285 15685 18315 15690
rect 18365 15710 18395 15715
rect 18365 15690 18370 15710
rect 18370 15690 18390 15710
rect 18390 15690 18395 15710
rect 18365 15685 18395 15690
rect 18445 15710 18475 15715
rect 18445 15690 18450 15710
rect 18450 15690 18470 15710
rect 18470 15690 18475 15710
rect 18445 15685 18475 15690
rect 18525 15710 18555 15715
rect 18525 15690 18530 15710
rect 18530 15690 18550 15710
rect 18550 15690 18555 15710
rect 18525 15685 18555 15690
rect 18605 15710 18635 15715
rect 18605 15690 18610 15710
rect 18610 15690 18630 15710
rect 18630 15690 18635 15710
rect 18605 15685 18635 15690
rect 18685 15710 18715 15715
rect 18685 15690 18690 15710
rect 18690 15690 18710 15710
rect 18710 15690 18715 15710
rect 18685 15685 18715 15690
rect 18765 15710 18795 15715
rect 18765 15690 18770 15710
rect 18770 15690 18790 15710
rect 18790 15690 18795 15710
rect 18765 15685 18795 15690
rect 18845 15710 18875 15715
rect 18845 15690 18850 15710
rect 18850 15690 18870 15710
rect 18870 15690 18875 15710
rect 18845 15685 18875 15690
rect 18925 15710 18955 15715
rect 18925 15690 18930 15710
rect 18930 15690 18950 15710
rect 18950 15690 18955 15710
rect 18925 15685 18955 15690
rect 19005 15710 19035 15715
rect 19005 15690 19010 15710
rect 19010 15690 19030 15710
rect 19030 15690 19035 15710
rect 19005 15685 19035 15690
rect 19085 15710 19115 15715
rect 19085 15690 19090 15710
rect 19090 15690 19110 15710
rect 19110 15690 19115 15710
rect 19085 15685 19115 15690
rect 19165 15710 19195 15715
rect 19165 15690 19170 15710
rect 19170 15690 19190 15710
rect 19190 15690 19195 15710
rect 19165 15685 19195 15690
rect 19245 15710 19275 15715
rect 19245 15690 19250 15710
rect 19250 15690 19270 15710
rect 19270 15690 19275 15710
rect 19245 15685 19275 15690
rect 19325 15710 19355 15715
rect 19325 15690 19330 15710
rect 19330 15690 19350 15710
rect 19350 15690 19355 15710
rect 19325 15685 19355 15690
rect 19405 15710 19435 15715
rect 19405 15690 19410 15710
rect 19410 15690 19430 15710
rect 19430 15690 19435 15710
rect 19405 15685 19435 15690
rect 19485 15710 19515 15715
rect 19485 15690 19490 15710
rect 19490 15690 19510 15710
rect 19510 15690 19515 15710
rect 19485 15685 19515 15690
rect 19565 15710 19595 15715
rect 19565 15690 19570 15710
rect 19570 15690 19590 15710
rect 19590 15690 19595 15710
rect 19565 15685 19595 15690
rect 19645 15710 19675 15715
rect 19645 15690 19650 15710
rect 19650 15690 19670 15710
rect 19670 15690 19675 15710
rect 19645 15685 19675 15690
rect 19725 15710 19755 15715
rect 19725 15690 19730 15710
rect 19730 15690 19750 15710
rect 19750 15690 19755 15710
rect 19725 15685 19755 15690
rect 19805 15710 19835 15715
rect 19805 15690 19810 15710
rect 19810 15690 19830 15710
rect 19830 15690 19835 15710
rect 19805 15685 19835 15690
rect 19885 15710 19915 15715
rect 19885 15690 19890 15710
rect 19890 15690 19910 15710
rect 19910 15690 19915 15710
rect 19885 15685 19915 15690
rect 19965 15710 19995 15715
rect 19965 15690 19970 15710
rect 19970 15690 19990 15710
rect 19990 15690 19995 15710
rect 19965 15685 19995 15690
rect 20045 15710 20075 15715
rect 20045 15690 20050 15710
rect 20050 15690 20070 15710
rect 20070 15690 20075 15710
rect 20045 15685 20075 15690
rect 20125 15710 20155 15715
rect 20125 15690 20130 15710
rect 20130 15690 20150 15710
rect 20150 15690 20155 15710
rect 20125 15685 20155 15690
rect 20205 15710 20235 15715
rect 20205 15690 20210 15710
rect 20210 15690 20230 15710
rect 20230 15690 20235 15710
rect 20205 15685 20235 15690
rect 20285 15710 20315 15715
rect 20285 15690 20290 15710
rect 20290 15690 20310 15710
rect 20310 15690 20315 15710
rect 20285 15685 20315 15690
rect 20365 15710 20395 15715
rect 20365 15690 20370 15710
rect 20370 15690 20390 15710
rect 20390 15690 20395 15710
rect 20365 15685 20395 15690
rect 20445 15710 20475 15715
rect 20445 15690 20450 15710
rect 20450 15690 20470 15710
rect 20470 15690 20475 15710
rect 20445 15685 20475 15690
rect 20525 15710 20555 15715
rect 20525 15690 20530 15710
rect 20530 15690 20550 15710
rect 20550 15690 20555 15710
rect 20525 15685 20555 15690
rect 20605 15710 20635 15715
rect 20605 15690 20610 15710
rect 20610 15690 20630 15710
rect 20630 15690 20635 15710
rect 20605 15685 20635 15690
rect 20685 15710 20715 15715
rect 20685 15690 20690 15710
rect 20690 15690 20710 15710
rect 20710 15690 20715 15710
rect 20685 15685 20715 15690
rect 20765 15710 20795 15715
rect 20765 15690 20770 15710
rect 20770 15690 20790 15710
rect 20790 15690 20795 15710
rect 20765 15685 20795 15690
rect 20845 15710 20875 15715
rect 20845 15690 20850 15710
rect 20850 15690 20870 15710
rect 20870 15690 20875 15710
rect 20845 15685 20875 15690
rect 20925 15710 20955 15715
rect 20925 15690 20930 15710
rect 20930 15690 20950 15710
rect 20950 15690 20955 15710
rect 20925 15685 20955 15690
rect 5 15550 35 15555
rect 5 15530 10 15550
rect 10 15530 30 15550
rect 30 15530 35 15550
rect 5 15525 35 15530
rect 85 15550 115 15555
rect 85 15530 90 15550
rect 90 15530 110 15550
rect 110 15530 115 15550
rect 85 15525 115 15530
rect 165 15550 195 15555
rect 165 15530 170 15550
rect 170 15530 190 15550
rect 190 15530 195 15550
rect 165 15525 195 15530
rect 245 15550 275 15555
rect 245 15530 250 15550
rect 250 15530 270 15550
rect 270 15530 275 15550
rect 245 15525 275 15530
rect 325 15550 355 15555
rect 325 15530 330 15550
rect 330 15530 350 15550
rect 350 15530 355 15550
rect 325 15525 355 15530
rect 405 15550 435 15555
rect 405 15530 410 15550
rect 410 15530 430 15550
rect 430 15530 435 15550
rect 405 15525 435 15530
rect 485 15550 515 15555
rect 485 15530 490 15550
rect 490 15530 510 15550
rect 510 15530 515 15550
rect 485 15525 515 15530
rect 565 15550 595 15555
rect 565 15530 570 15550
rect 570 15530 590 15550
rect 590 15530 595 15550
rect 565 15525 595 15530
rect 645 15550 675 15555
rect 645 15530 650 15550
rect 650 15530 670 15550
rect 670 15530 675 15550
rect 645 15525 675 15530
rect 725 15550 755 15555
rect 725 15530 730 15550
rect 730 15530 750 15550
rect 750 15530 755 15550
rect 725 15525 755 15530
rect 805 15550 835 15555
rect 805 15530 810 15550
rect 810 15530 830 15550
rect 830 15530 835 15550
rect 805 15525 835 15530
rect 885 15550 915 15555
rect 885 15530 890 15550
rect 890 15530 910 15550
rect 910 15530 915 15550
rect 885 15525 915 15530
rect 965 15550 995 15555
rect 965 15530 970 15550
rect 970 15530 990 15550
rect 990 15530 995 15550
rect 965 15525 995 15530
rect 1045 15550 1075 15555
rect 1045 15530 1050 15550
rect 1050 15530 1070 15550
rect 1070 15530 1075 15550
rect 1045 15525 1075 15530
rect 1125 15550 1155 15555
rect 1125 15530 1130 15550
rect 1130 15530 1150 15550
rect 1150 15530 1155 15550
rect 1125 15525 1155 15530
rect 1205 15550 1235 15555
rect 1205 15530 1210 15550
rect 1210 15530 1230 15550
rect 1230 15530 1235 15550
rect 1205 15525 1235 15530
rect 1285 15550 1315 15555
rect 1285 15530 1290 15550
rect 1290 15530 1310 15550
rect 1310 15530 1315 15550
rect 1285 15525 1315 15530
rect 1365 15550 1395 15555
rect 1365 15530 1370 15550
rect 1370 15530 1390 15550
rect 1390 15530 1395 15550
rect 1365 15525 1395 15530
rect 1445 15550 1475 15555
rect 1445 15530 1450 15550
rect 1450 15530 1470 15550
rect 1470 15530 1475 15550
rect 1445 15525 1475 15530
rect 1525 15550 1555 15555
rect 1525 15530 1530 15550
rect 1530 15530 1550 15550
rect 1550 15530 1555 15550
rect 1525 15525 1555 15530
rect 1605 15550 1635 15555
rect 1605 15530 1610 15550
rect 1610 15530 1630 15550
rect 1630 15530 1635 15550
rect 1605 15525 1635 15530
rect 1685 15550 1715 15555
rect 1685 15530 1690 15550
rect 1690 15530 1710 15550
rect 1710 15530 1715 15550
rect 1685 15525 1715 15530
rect 1765 15550 1795 15555
rect 1765 15530 1770 15550
rect 1770 15530 1790 15550
rect 1790 15530 1795 15550
rect 1765 15525 1795 15530
rect 1845 15550 1875 15555
rect 1845 15530 1850 15550
rect 1850 15530 1870 15550
rect 1870 15530 1875 15550
rect 1845 15525 1875 15530
rect 1925 15550 1955 15555
rect 1925 15530 1930 15550
rect 1930 15530 1950 15550
rect 1950 15530 1955 15550
rect 1925 15525 1955 15530
rect 2005 15550 2035 15555
rect 2005 15530 2010 15550
rect 2010 15530 2030 15550
rect 2030 15530 2035 15550
rect 2005 15525 2035 15530
rect 2085 15550 2115 15555
rect 2085 15530 2090 15550
rect 2090 15530 2110 15550
rect 2110 15530 2115 15550
rect 2085 15525 2115 15530
rect 2165 15550 2195 15555
rect 2165 15530 2170 15550
rect 2170 15530 2190 15550
rect 2190 15530 2195 15550
rect 2165 15525 2195 15530
rect 2245 15550 2275 15555
rect 2245 15530 2250 15550
rect 2250 15530 2270 15550
rect 2270 15530 2275 15550
rect 2245 15525 2275 15530
rect 2325 15550 2355 15555
rect 2325 15530 2330 15550
rect 2330 15530 2350 15550
rect 2350 15530 2355 15550
rect 2325 15525 2355 15530
rect 2405 15550 2435 15555
rect 2405 15530 2410 15550
rect 2410 15530 2430 15550
rect 2430 15530 2435 15550
rect 2405 15525 2435 15530
rect 2485 15550 2515 15555
rect 2485 15530 2490 15550
rect 2490 15530 2510 15550
rect 2510 15530 2515 15550
rect 2485 15525 2515 15530
rect 2565 15550 2595 15555
rect 2565 15530 2570 15550
rect 2570 15530 2590 15550
rect 2590 15530 2595 15550
rect 2565 15525 2595 15530
rect 2645 15550 2675 15555
rect 2645 15530 2650 15550
rect 2650 15530 2670 15550
rect 2670 15530 2675 15550
rect 2645 15525 2675 15530
rect 2725 15550 2755 15555
rect 2725 15530 2730 15550
rect 2730 15530 2750 15550
rect 2750 15530 2755 15550
rect 2725 15525 2755 15530
rect 2805 15550 2835 15555
rect 2805 15530 2810 15550
rect 2810 15530 2830 15550
rect 2830 15530 2835 15550
rect 2805 15525 2835 15530
rect 2885 15550 2915 15555
rect 2885 15530 2890 15550
rect 2890 15530 2910 15550
rect 2910 15530 2915 15550
rect 2885 15525 2915 15530
rect 2965 15550 2995 15555
rect 2965 15530 2970 15550
rect 2970 15530 2990 15550
rect 2990 15530 2995 15550
rect 2965 15525 2995 15530
rect 3045 15550 3075 15555
rect 3045 15530 3050 15550
rect 3050 15530 3070 15550
rect 3070 15530 3075 15550
rect 3045 15525 3075 15530
rect 3125 15550 3155 15555
rect 3125 15530 3130 15550
rect 3130 15530 3150 15550
rect 3150 15530 3155 15550
rect 3125 15525 3155 15530
rect 3205 15550 3235 15555
rect 3205 15530 3210 15550
rect 3210 15530 3230 15550
rect 3230 15530 3235 15550
rect 3205 15525 3235 15530
rect 3285 15550 3315 15555
rect 3285 15530 3290 15550
rect 3290 15530 3310 15550
rect 3310 15530 3315 15550
rect 3285 15525 3315 15530
rect 3365 15550 3395 15555
rect 3365 15530 3370 15550
rect 3370 15530 3390 15550
rect 3390 15530 3395 15550
rect 3365 15525 3395 15530
rect 3445 15550 3475 15555
rect 3445 15530 3450 15550
rect 3450 15530 3470 15550
rect 3470 15530 3475 15550
rect 3445 15525 3475 15530
rect 3525 15550 3555 15555
rect 3525 15530 3530 15550
rect 3530 15530 3550 15550
rect 3550 15530 3555 15550
rect 3525 15525 3555 15530
rect 3605 15550 3635 15555
rect 3605 15530 3610 15550
rect 3610 15530 3630 15550
rect 3630 15530 3635 15550
rect 3605 15525 3635 15530
rect 3685 15550 3715 15555
rect 3685 15530 3690 15550
rect 3690 15530 3710 15550
rect 3710 15530 3715 15550
rect 3685 15525 3715 15530
rect 3765 15550 3795 15555
rect 3765 15530 3770 15550
rect 3770 15530 3790 15550
rect 3790 15530 3795 15550
rect 3765 15525 3795 15530
rect 3845 15550 3875 15555
rect 3845 15530 3850 15550
rect 3850 15530 3870 15550
rect 3870 15530 3875 15550
rect 3845 15525 3875 15530
rect 3925 15550 3955 15555
rect 3925 15530 3930 15550
rect 3930 15530 3950 15550
rect 3950 15530 3955 15550
rect 3925 15525 3955 15530
rect 4005 15550 4035 15555
rect 4005 15530 4010 15550
rect 4010 15530 4030 15550
rect 4030 15530 4035 15550
rect 4005 15525 4035 15530
rect 4085 15550 4115 15555
rect 4085 15530 4090 15550
rect 4090 15530 4110 15550
rect 4110 15530 4115 15550
rect 4085 15525 4115 15530
rect 4165 15550 4195 15555
rect 4165 15530 4170 15550
rect 4170 15530 4190 15550
rect 4190 15530 4195 15550
rect 4165 15525 4195 15530
rect 6245 15550 6275 15555
rect 6245 15530 6250 15550
rect 6250 15530 6270 15550
rect 6270 15530 6275 15550
rect 6245 15525 6275 15530
rect 6325 15550 6355 15555
rect 6325 15530 6330 15550
rect 6330 15530 6350 15550
rect 6350 15530 6355 15550
rect 6325 15525 6355 15530
rect 6405 15550 6435 15555
rect 6405 15530 6410 15550
rect 6410 15530 6430 15550
rect 6430 15530 6435 15550
rect 6405 15525 6435 15530
rect 6485 15550 6515 15555
rect 6485 15530 6490 15550
rect 6490 15530 6510 15550
rect 6510 15530 6515 15550
rect 6485 15525 6515 15530
rect 6565 15550 6595 15555
rect 6565 15530 6570 15550
rect 6570 15530 6590 15550
rect 6590 15530 6595 15550
rect 6565 15525 6595 15530
rect 6645 15550 6675 15555
rect 6645 15530 6650 15550
rect 6650 15530 6670 15550
rect 6670 15530 6675 15550
rect 6645 15525 6675 15530
rect 6725 15550 6755 15555
rect 6725 15530 6730 15550
rect 6730 15530 6750 15550
rect 6750 15530 6755 15550
rect 6725 15525 6755 15530
rect 6805 15550 6835 15555
rect 6805 15530 6810 15550
rect 6810 15530 6830 15550
rect 6830 15530 6835 15550
rect 6805 15525 6835 15530
rect 6885 15550 6915 15555
rect 6885 15530 6890 15550
rect 6890 15530 6910 15550
rect 6910 15530 6915 15550
rect 6885 15525 6915 15530
rect 6965 15550 6995 15555
rect 6965 15530 6970 15550
rect 6970 15530 6990 15550
rect 6990 15530 6995 15550
rect 6965 15525 6995 15530
rect 7045 15550 7075 15555
rect 7045 15530 7050 15550
rect 7050 15530 7070 15550
rect 7070 15530 7075 15550
rect 7045 15525 7075 15530
rect 7125 15550 7155 15555
rect 7125 15530 7130 15550
rect 7130 15530 7150 15550
rect 7150 15530 7155 15550
rect 7125 15525 7155 15530
rect 7205 15550 7235 15555
rect 7205 15530 7210 15550
rect 7210 15530 7230 15550
rect 7230 15530 7235 15550
rect 7205 15525 7235 15530
rect 7285 15550 7315 15555
rect 7285 15530 7290 15550
rect 7290 15530 7310 15550
rect 7310 15530 7315 15550
rect 7285 15525 7315 15530
rect 7365 15550 7395 15555
rect 7365 15530 7370 15550
rect 7370 15530 7390 15550
rect 7390 15530 7395 15550
rect 7365 15525 7395 15530
rect 7445 15550 7475 15555
rect 7445 15530 7450 15550
rect 7450 15530 7470 15550
rect 7470 15530 7475 15550
rect 7445 15525 7475 15530
rect 7525 15550 7555 15555
rect 7525 15530 7530 15550
rect 7530 15530 7550 15550
rect 7550 15530 7555 15550
rect 7525 15525 7555 15530
rect 7605 15550 7635 15555
rect 7605 15530 7610 15550
rect 7610 15530 7630 15550
rect 7630 15530 7635 15550
rect 7605 15525 7635 15530
rect 7685 15550 7715 15555
rect 7685 15530 7690 15550
rect 7690 15530 7710 15550
rect 7710 15530 7715 15550
rect 7685 15525 7715 15530
rect 7765 15550 7795 15555
rect 7765 15530 7770 15550
rect 7770 15530 7790 15550
rect 7790 15530 7795 15550
rect 7765 15525 7795 15530
rect 7845 15550 7875 15555
rect 7845 15530 7850 15550
rect 7850 15530 7870 15550
rect 7870 15530 7875 15550
rect 7845 15525 7875 15530
rect 7925 15550 7955 15555
rect 7925 15530 7930 15550
rect 7930 15530 7950 15550
rect 7950 15530 7955 15550
rect 7925 15525 7955 15530
rect 8005 15550 8035 15555
rect 8005 15530 8010 15550
rect 8010 15530 8030 15550
rect 8030 15530 8035 15550
rect 8005 15525 8035 15530
rect 8085 15550 8115 15555
rect 8085 15530 8090 15550
rect 8090 15530 8110 15550
rect 8110 15530 8115 15550
rect 8085 15525 8115 15530
rect 8165 15550 8195 15555
rect 8165 15530 8170 15550
rect 8170 15530 8190 15550
rect 8190 15530 8195 15550
rect 8165 15525 8195 15530
rect 8245 15550 8275 15555
rect 8245 15530 8250 15550
rect 8250 15530 8270 15550
rect 8270 15530 8275 15550
rect 8245 15525 8275 15530
rect 8325 15550 8355 15555
rect 8325 15530 8330 15550
rect 8330 15530 8350 15550
rect 8350 15530 8355 15550
rect 8325 15525 8355 15530
rect 8405 15550 8435 15555
rect 8405 15530 8410 15550
rect 8410 15530 8430 15550
rect 8430 15530 8435 15550
rect 8405 15525 8435 15530
rect 8485 15550 8515 15555
rect 8485 15530 8490 15550
rect 8490 15530 8510 15550
rect 8510 15530 8515 15550
rect 8485 15525 8515 15530
rect 8565 15550 8595 15555
rect 8565 15530 8570 15550
rect 8570 15530 8590 15550
rect 8590 15530 8595 15550
rect 8565 15525 8595 15530
rect 8645 15550 8675 15555
rect 8645 15530 8650 15550
rect 8650 15530 8670 15550
rect 8670 15530 8675 15550
rect 8645 15525 8675 15530
rect 8725 15550 8755 15555
rect 8725 15530 8730 15550
rect 8730 15530 8750 15550
rect 8750 15530 8755 15550
rect 8725 15525 8755 15530
rect 8805 15550 8835 15555
rect 8805 15530 8810 15550
rect 8810 15530 8830 15550
rect 8830 15530 8835 15550
rect 8805 15525 8835 15530
rect 8885 15550 8915 15555
rect 8885 15530 8890 15550
rect 8890 15530 8910 15550
rect 8910 15530 8915 15550
rect 8885 15525 8915 15530
rect 8965 15550 8995 15555
rect 8965 15530 8970 15550
rect 8970 15530 8990 15550
rect 8990 15530 8995 15550
rect 8965 15525 8995 15530
rect 9045 15550 9075 15555
rect 9045 15530 9050 15550
rect 9050 15530 9070 15550
rect 9070 15530 9075 15550
rect 9045 15525 9075 15530
rect 9125 15550 9155 15555
rect 9125 15530 9130 15550
rect 9130 15530 9150 15550
rect 9150 15530 9155 15550
rect 9125 15525 9155 15530
rect 9205 15550 9235 15555
rect 9205 15530 9210 15550
rect 9210 15530 9230 15550
rect 9230 15530 9235 15550
rect 9205 15525 9235 15530
rect 9285 15550 9315 15555
rect 9285 15530 9290 15550
rect 9290 15530 9310 15550
rect 9310 15530 9315 15550
rect 9285 15525 9315 15530
rect 9365 15550 9395 15555
rect 9365 15530 9370 15550
rect 9370 15530 9390 15550
rect 9390 15530 9395 15550
rect 9365 15525 9395 15530
rect 9445 15550 9475 15555
rect 9445 15530 9450 15550
rect 9450 15530 9470 15550
rect 9470 15530 9475 15550
rect 9445 15525 9475 15530
rect 11565 15550 11595 15555
rect 11565 15530 11570 15550
rect 11570 15530 11590 15550
rect 11590 15530 11595 15550
rect 11565 15525 11595 15530
rect 11645 15550 11675 15555
rect 11645 15530 11650 15550
rect 11650 15530 11670 15550
rect 11670 15530 11675 15550
rect 11645 15525 11675 15530
rect 11725 15550 11755 15555
rect 11725 15530 11730 15550
rect 11730 15530 11750 15550
rect 11750 15530 11755 15550
rect 11725 15525 11755 15530
rect 11805 15550 11835 15555
rect 11805 15530 11810 15550
rect 11810 15530 11830 15550
rect 11830 15530 11835 15550
rect 11805 15525 11835 15530
rect 11885 15550 11915 15555
rect 11885 15530 11890 15550
rect 11890 15530 11910 15550
rect 11910 15530 11915 15550
rect 11885 15525 11915 15530
rect 11965 15550 11995 15555
rect 11965 15530 11970 15550
rect 11970 15530 11990 15550
rect 11990 15530 11995 15550
rect 11965 15525 11995 15530
rect 12045 15550 12075 15555
rect 12045 15530 12050 15550
rect 12050 15530 12070 15550
rect 12070 15530 12075 15550
rect 12045 15525 12075 15530
rect 12125 15550 12155 15555
rect 12125 15530 12130 15550
rect 12130 15530 12150 15550
rect 12150 15530 12155 15550
rect 12125 15525 12155 15530
rect 12205 15550 12235 15555
rect 12205 15530 12210 15550
rect 12210 15530 12230 15550
rect 12230 15530 12235 15550
rect 12205 15525 12235 15530
rect 12285 15550 12315 15555
rect 12285 15530 12290 15550
rect 12290 15530 12310 15550
rect 12310 15530 12315 15550
rect 12285 15525 12315 15530
rect 12365 15550 12395 15555
rect 12365 15530 12370 15550
rect 12370 15530 12390 15550
rect 12390 15530 12395 15550
rect 12365 15525 12395 15530
rect 12445 15550 12475 15555
rect 12445 15530 12450 15550
rect 12450 15530 12470 15550
rect 12470 15530 12475 15550
rect 12445 15525 12475 15530
rect 12525 15550 12555 15555
rect 12525 15530 12530 15550
rect 12530 15530 12550 15550
rect 12550 15530 12555 15550
rect 12525 15525 12555 15530
rect 12605 15550 12635 15555
rect 12605 15530 12610 15550
rect 12610 15530 12630 15550
rect 12630 15530 12635 15550
rect 12605 15525 12635 15530
rect 12685 15550 12715 15555
rect 12685 15530 12690 15550
rect 12690 15530 12710 15550
rect 12710 15530 12715 15550
rect 12685 15525 12715 15530
rect 12765 15550 12795 15555
rect 12765 15530 12770 15550
rect 12770 15530 12790 15550
rect 12790 15530 12795 15550
rect 12765 15525 12795 15530
rect 12845 15550 12875 15555
rect 12845 15530 12850 15550
rect 12850 15530 12870 15550
rect 12870 15530 12875 15550
rect 12845 15525 12875 15530
rect 12925 15550 12955 15555
rect 12925 15530 12930 15550
rect 12930 15530 12950 15550
rect 12950 15530 12955 15550
rect 12925 15525 12955 15530
rect 13005 15550 13035 15555
rect 13005 15530 13010 15550
rect 13010 15530 13030 15550
rect 13030 15530 13035 15550
rect 13005 15525 13035 15530
rect 13085 15550 13115 15555
rect 13085 15530 13090 15550
rect 13090 15530 13110 15550
rect 13110 15530 13115 15550
rect 13085 15525 13115 15530
rect 13165 15550 13195 15555
rect 13165 15530 13170 15550
rect 13170 15530 13190 15550
rect 13190 15530 13195 15550
rect 13165 15525 13195 15530
rect 13245 15550 13275 15555
rect 13245 15530 13250 15550
rect 13250 15530 13270 15550
rect 13270 15530 13275 15550
rect 13245 15525 13275 15530
rect 13325 15550 13355 15555
rect 13325 15530 13330 15550
rect 13330 15530 13350 15550
rect 13350 15530 13355 15550
rect 13325 15525 13355 15530
rect 13405 15550 13435 15555
rect 13405 15530 13410 15550
rect 13410 15530 13430 15550
rect 13430 15530 13435 15550
rect 13405 15525 13435 15530
rect 13485 15550 13515 15555
rect 13485 15530 13490 15550
rect 13490 15530 13510 15550
rect 13510 15530 13515 15550
rect 13485 15525 13515 15530
rect 13565 15550 13595 15555
rect 13565 15530 13570 15550
rect 13570 15530 13590 15550
rect 13590 15530 13595 15550
rect 13565 15525 13595 15530
rect 13645 15550 13675 15555
rect 13645 15530 13650 15550
rect 13650 15530 13670 15550
rect 13670 15530 13675 15550
rect 13645 15525 13675 15530
rect 13725 15550 13755 15555
rect 13725 15530 13730 15550
rect 13730 15530 13750 15550
rect 13750 15530 13755 15550
rect 13725 15525 13755 15530
rect 13805 15550 13835 15555
rect 13805 15530 13810 15550
rect 13810 15530 13830 15550
rect 13830 15530 13835 15550
rect 13805 15525 13835 15530
rect 13885 15550 13915 15555
rect 13885 15530 13890 15550
rect 13890 15530 13910 15550
rect 13910 15530 13915 15550
rect 13885 15525 13915 15530
rect 13965 15550 13995 15555
rect 13965 15530 13970 15550
rect 13970 15530 13990 15550
rect 13990 15530 13995 15550
rect 13965 15525 13995 15530
rect 14045 15550 14075 15555
rect 14045 15530 14050 15550
rect 14050 15530 14070 15550
rect 14070 15530 14075 15550
rect 14045 15525 14075 15530
rect 14125 15550 14155 15555
rect 14125 15530 14130 15550
rect 14130 15530 14150 15550
rect 14150 15530 14155 15550
rect 14125 15525 14155 15530
rect 14205 15550 14235 15555
rect 14205 15530 14210 15550
rect 14210 15530 14230 15550
rect 14230 15530 14235 15550
rect 14205 15525 14235 15530
rect 14285 15550 14315 15555
rect 14285 15530 14290 15550
rect 14290 15530 14310 15550
rect 14310 15530 14315 15550
rect 14285 15525 14315 15530
rect 14365 15550 14395 15555
rect 14365 15530 14370 15550
rect 14370 15530 14390 15550
rect 14390 15530 14395 15550
rect 14365 15525 14395 15530
rect 14445 15550 14475 15555
rect 14445 15530 14450 15550
rect 14450 15530 14470 15550
rect 14470 15530 14475 15550
rect 14445 15525 14475 15530
rect 14525 15550 14555 15555
rect 14525 15530 14530 15550
rect 14530 15530 14550 15550
rect 14550 15530 14555 15550
rect 14525 15525 14555 15530
rect 14605 15550 14635 15555
rect 14605 15530 14610 15550
rect 14610 15530 14630 15550
rect 14630 15530 14635 15550
rect 14605 15525 14635 15530
rect 14685 15550 14715 15555
rect 14685 15530 14690 15550
rect 14690 15530 14710 15550
rect 14710 15530 14715 15550
rect 14685 15525 14715 15530
rect 16765 15550 16795 15555
rect 16765 15530 16770 15550
rect 16770 15530 16790 15550
rect 16790 15530 16795 15550
rect 16765 15525 16795 15530
rect 16845 15550 16875 15555
rect 16845 15530 16850 15550
rect 16850 15530 16870 15550
rect 16870 15530 16875 15550
rect 16845 15525 16875 15530
rect 16925 15550 16955 15555
rect 16925 15530 16930 15550
rect 16930 15530 16950 15550
rect 16950 15530 16955 15550
rect 16925 15525 16955 15530
rect 17005 15550 17035 15555
rect 17005 15530 17010 15550
rect 17010 15530 17030 15550
rect 17030 15530 17035 15550
rect 17005 15525 17035 15530
rect 17085 15550 17115 15555
rect 17085 15530 17090 15550
rect 17090 15530 17110 15550
rect 17110 15530 17115 15550
rect 17085 15525 17115 15530
rect 17165 15550 17195 15555
rect 17165 15530 17170 15550
rect 17170 15530 17190 15550
rect 17190 15530 17195 15550
rect 17165 15525 17195 15530
rect 17245 15550 17275 15555
rect 17245 15530 17250 15550
rect 17250 15530 17270 15550
rect 17270 15530 17275 15550
rect 17245 15525 17275 15530
rect 17325 15550 17355 15555
rect 17325 15530 17330 15550
rect 17330 15530 17350 15550
rect 17350 15530 17355 15550
rect 17325 15525 17355 15530
rect 17405 15550 17435 15555
rect 17405 15530 17410 15550
rect 17410 15530 17430 15550
rect 17430 15530 17435 15550
rect 17405 15525 17435 15530
rect 17485 15550 17515 15555
rect 17485 15530 17490 15550
rect 17490 15530 17510 15550
rect 17510 15530 17515 15550
rect 17485 15525 17515 15530
rect 17565 15550 17595 15555
rect 17565 15530 17570 15550
rect 17570 15530 17590 15550
rect 17590 15530 17595 15550
rect 17565 15525 17595 15530
rect 17645 15550 17675 15555
rect 17645 15530 17650 15550
rect 17650 15530 17670 15550
rect 17670 15530 17675 15550
rect 17645 15525 17675 15530
rect 17725 15550 17755 15555
rect 17725 15530 17730 15550
rect 17730 15530 17750 15550
rect 17750 15530 17755 15550
rect 17725 15525 17755 15530
rect 17805 15550 17835 15555
rect 17805 15530 17810 15550
rect 17810 15530 17830 15550
rect 17830 15530 17835 15550
rect 17805 15525 17835 15530
rect 17885 15550 17915 15555
rect 17885 15530 17890 15550
rect 17890 15530 17910 15550
rect 17910 15530 17915 15550
rect 17885 15525 17915 15530
rect 17965 15550 17995 15555
rect 17965 15530 17970 15550
rect 17970 15530 17990 15550
rect 17990 15530 17995 15550
rect 17965 15525 17995 15530
rect 18045 15550 18075 15555
rect 18045 15530 18050 15550
rect 18050 15530 18070 15550
rect 18070 15530 18075 15550
rect 18045 15525 18075 15530
rect 18125 15550 18155 15555
rect 18125 15530 18130 15550
rect 18130 15530 18150 15550
rect 18150 15530 18155 15550
rect 18125 15525 18155 15530
rect 18205 15550 18235 15555
rect 18205 15530 18210 15550
rect 18210 15530 18230 15550
rect 18230 15530 18235 15550
rect 18205 15525 18235 15530
rect 18285 15550 18315 15555
rect 18285 15530 18290 15550
rect 18290 15530 18310 15550
rect 18310 15530 18315 15550
rect 18285 15525 18315 15530
rect 18365 15550 18395 15555
rect 18365 15530 18370 15550
rect 18370 15530 18390 15550
rect 18390 15530 18395 15550
rect 18365 15525 18395 15530
rect 18445 15550 18475 15555
rect 18445 15530 18450 15550
rect 18450 15530 18470 15550
rect 18470 15530 18475 15550
rect 18445 15525 18475 15530
rect 18525 15550 18555 15555
rect 18525 15530 18530 15550
rect 18530 15530 18550 15550
rect 18550 15530 18555 15550
rect 18525 15525 18555 15530
rect 18605 15550 18635 15555
rect 18605 15530 18610 15550
rect 18610 15530 18630 15550
rect 18630 15530 18635 15550
rect 18605 15525 18635 15530
rect 18685 15550 18715 15555
rect 18685 15530 18690 15550
rect 18690 15530 18710 15550
rect 18710 15530 18715 15550
rect 18685 15525 18715 15530
rect 18765 15550 18795 15555
rect 18765 15530 18770 15550
rect 18770 15530 18790 15550
rect 18790 15530 18795 15550
rect 18765 15525 18795 15530
rect 18845 15550 18875 15555
rect 18845 15530 18850 15550
rect 18850 15530 18870 15550
rect 18870 15530 18875 15550
rect 18845 15525 18875 15530
rect 18925 15550 18955 15555
rect 18925 15530 18930 15550
rect 18930 15530 18950 15550
rect 18950 15530 18955 15550
rect 18925 15525 18955 15530
rect 19005 15550 19035 15555
rect 19005 15530 19010 15550
rect 19010 15530 19030 15550
rect 19030 15530 19035 15550
rect 19005 15525 19035 15530
rect 19085 15550 19115 15555
rect 19085 15530 19090 15550
rect 19090 15530 19110 15550
rect 19110 15530 19115 15550
rect 19085 15525 19115 15530
rect 19165 15550 19195 15555
rect 19165 15530 19170 15550
rect 19170 15530 19190 15550
rect 19190 15530 19195 15550
rect 19165 15525 19195 15530
rect 19245 15550 19275 15555
rect 19245 15530 19250 15550
rect 19250 15530 19270 15550
rect 19270 15530 19275 15550
rect 19245 15525 19275 15530
rect 19325 15550 19355 15555
rect 19325 15530 19330 15550
rect 19330 15530 19350 15550
rect 19350 15530 19355 15550
rect 19325 15525 19355 15530
rect 19405 15550 19435 15555
rect 19405 15530 19410 15550
rect 19410 15530 19430 15550
rect 19430 15530 19435 15550
rect 19405 15525 19435 15530
rect 19485 15550 19515 15555
rect 19485 15530 19490 15550
rect 19490 15530 19510 15550
rect 19510 15530 19515 15550
rect 19485 15525 19515 15530
rect 19565 15550 19595 15555
rect 19565 15530 19570 15550
rect 19570 15530 19590 15550
rect 19590 15530 19595 15550
rect 19565 15525 19595 15530
rect 19645 15550 19675 15555
rect 19645 15530 19650 15550
rect 19650 15530 19670 15550
rect 19670 15530 19675 15550
rect 19645 15525 19675 15530
rect 19725 15550 19755 15555
rect 19725 15530 19730 15550
rect 19730 15530 19750 15550
rect 19750 15530 19755 15550
rect 19725 15525 19755 15530
rect 19805 15550 19835 15555
rect 19805 15530 19810 15550
rect 19810 15530 19830 15550
rect 19830 15530 19835 15550
rect 19805 15525 19835 15530
rect 19885 15550 19915 15555
rect 19885 15530 19890 15550
rect 19890 15530 19910 15550
rect 19910 15530 19915 15550
rect 19885 15525 19915 15530
rect 19965 15550 19995 15555
rect 19965 15530 19970 15550
rect 19970 15530 19990 15550
rect 19990 15530 19995 15550
rect 19965 15525 19995 15530
rect 20045 15550 20075 15555
rect 20045 15530 20050 15550
rect 20050 15530 20070 15550
rect 20070 15530 20075 15550
rect 20045 15525 20075 15530
rect 20125 15550 20155 15555
rect 20125 15530 20130 15550
rect 20130 15530 20150 15550
rect 20150 15530 20155 15550
rect 20125 15525 20155 15530
rect 20205 15550 20235 15555
rect 20205 15530 20210 15550
rect 20210 15530 20230 15550
rect 20230 15530 20235 15550
rect 20205 15525 20235 15530
rect 20285 15550 20315 15555
rect 20285 15530 20290 15550
rect 20290 15530 20310 15550
rect 20310 15530 20315 15550
rect 20285 15525 20315 15530
rect 20365 15550 20395 15555
rect 20365 15530 20370 15550
rect 20370 15530 20390 15550
rect 20390 15530 20395 15550
rect 20365 15525 20395 15530
rect 20445 15550 20475 15555
rect 20445 15530 20450 15550
rect 20450 15530 20470 15550
rect 20470 15530 20475 15550
rect 20445 15525 20475 15530
rect 20525 15550 20555 15555
rect 20525 15530 20530 15550
rect 20530 15530 20550 15550
rect 20550 15530 20555 15550
rect 20525 15525 20555 15530
rect 20605 15550 20635 15555
rect 20605 15530 20610 15550
rect 20610 15530 20630 15550
rect 20630 15530 20635 15550
rect 20605 15525 20635 15530
rect 20685 15550 20715 15555
rect 20685 15530 20690 15550
rect 20690 15530 20710 15550
rect 20710 15530 20715 15550
rect 20685 15525 20715 15530
rect 20765 15550 20795 15555
rect 20765 15530 20770 15550
rect 20770 15530 20790 15550
rect 20790 15530 20795 15550
rect 20765 15525 20795 15530
rect 20845 15550 20875 15555
rect 20845 15530 20850 15550
rect 20850 15530 20870 15550
rect 20870 15530 20875 15550
rect 20845 15525 20875 15530
rect 20925 15550 20955 15555
rect 20925 15530 20930 15550
rect 20930 15530 20950 15550
rect 20950 15530 20955 15550
rect 20925 15525 20955 15530
rect 5 15390 35 15395
rect 5 15370 10 15390
rect 10 15370 30 15390
rect 30 15370 35 15390
rect 5 15365 35 15370
rect 85 15390 115 15395
rect 85 15370 90 15390
rect 90 15370 110 15390
rect 110 15370 115 15390
rect 85 15365 115 15370
rect 165 15390 195 15395
rect 165 15370 170 15390
rect 170 15370 190 15390
rect 190 15370 195 15390
rect 165 15365 195 15370
rect 245 15390 275 15395
rect 245 15370 250 15390
rect 250 15370 270 15390
rect 270 15370 275 15390
rect 245 15365 275 15370
rect 325 15390 355 15395
rect 325 15370 330 15390
rect 330 15370 350 15390
rect 350 15370 355 15390
rect 325 15365 355 15370
rect 405 15390 435 15395
rect 405 15370 410 15390
rect 410 15370 430 15390
rect 430 15370 435 15390
rect 405 15365 435 15370
rect 485 15390 515 15395
rect 485 15370 490 15390
rect 490 15370 510 15390
rect 510 15370 515 15390
rect 485 15365 515 15370
rect 565 15390 595 15395
rect 565 15370 570 15390
rect 570 15370 590 15390
rect 590 15370 595 15390
rect 565 15365 595 15370
rect 645 15390 675 15395
rect 645 15370 650 15390
rect 650 15370 670 15390
rect 670 15370 675 15390
rect 645 15365 675 15370
rect 725 15390 755 15395
rect 725 15370 730 15390
rect 730 15370 750 15390
rect 750 15370 755 15390
rect 725 15365 755 15370
rect 805 15390 835 15395
rect 805 15370 810 15390
rect 810 15370 830 15390
rect 830 15370 835 15390
rect 805 15365 835 15370
rect 885 15390 915 15395
rect 885 15370 890 15390
rect 890 15370 910 15390
rect 910 15370 915 15390
rect 885 15365 915 15370
rect 965 15390 995 15395
rect 965 15370 970 15390
rect 970 15370 990 15390
rect 990 15370 995 15390
rect 965 15365 995 15370
rect 1045 15390 1075 15395
rect 1045 15370 1050 15390
rect 1050 15370 1070 15390
rect 1070 15370 1075 15390
rect 1045 15365 1075 15370
rect 1125 15390 1155 15395
rect 1125 15370 1130 15390
rect 1130 15370 1150 15390
rect 1150 15370 1155 15390
rect 1125 15365 1155 15370
rect 1205 15390 1235 15395
rect 1205 15370 1210 15390
rect 1210 15370 1230 15390
rect 1230 15370 1235 15390
rect 1205 15365 1235 15370
rect 1285 15390 1315 15395
rect 1285 15370 1290 15390
rect 1290 15370 1310 15390
rect 1310 15370 1315 15390
rect 1285 15365 1315 15370
rect 1365 15390 1395 15395
rect 1365 15370 1370 15390
rect 1370 15370 1390 15390
rect 1390 15370 1395 15390
rect 1365 15365 1395 15370
rect 1445 15390 1475 15395
rect 1445 15370 1450 15390
rect 1450 15370 1470 15390
rect 1470 15370 1475 15390
rect 1445 15365 1475 15370
rect 1525 15390 1555 15395
rect 1525 15370 1530 15390
rect 1530 15370 1550 15390
rect 1550 15370 1555 15390
rect 1525 15365 1555 15370
rect 1605 15390 1635 15395
rect 1605 15370 1610 15390
rect 1610 15370 1630 15390
rect 1630 15370 1635 15390
rect 1605 15365 1635 15370
rect 1685 15390 1715 15395
rect 1685 15370 1690 15390
rect 1690 15370 1710 15390
rect 1710 15370 1715 15390
rect 1685 15365 1715 15370
rect 1765 15390 1795 15395
rect 1765 15370 1770 15390
rect 1770 15370 1790 15390
rect 1790 15370 1795 15390
rect 1765 15365 1795 15370
rect 1845 15390 1875 15395
rect 1845 15370 1850 15390
rect 1850 15370 1870 15390
rect 1870 15370 1875 15390
rect 1845 15365 1875 15370
rect 1925 15390 1955 15395
rect 1925 15370 1930 15390
rect 1930 15370 1950 15390
rect 1950 15370 1955 15390
rect 1925 15365 1955 15370
rect 2005 15390 2035 15395
rect 2005 15370 2010 15390
rect 2010 15370 2030 15390
rect 2030 15370 2035 15390
rect 2005 15365 2035 15370
rect 2085 15390 2115 15395
rect 2085 15370 2090 15390
rect 2090 15370 2110 15390
rect 2110 15370 2115 15390
rect 2085 15365 2115 15370
rect 2165 15390 2195 15395
rect 2165 15370 2170 15390
rect 2170 15370 2190 15390
rect 2190 15370 2195 15390
rect 2165 15365 2195 15370
rect 2245 15390 2275 15395
rect 2245 15370 2250 15390
rect 2250 15370 2270 15390
rect 2270 15370 2275 15390
rect 2245 15365 2275 15370
rect 2325 15390 2355 15395
rect 2325 15370 2330 15390
rect 2330 15370 2350 15390
rect 2350 15370 2355 15390
rect 2325 15365 2355 15370
rect 2405 15390 2435 15395
rect 2405 15370 2410 15390
rect 2410 15370 2430 15390
rect 2430 15370 2435 15390
rect 2405 15365 2435 15370
rect 2485 15390 2515 15395
rect 2485 15370 2490 15390
rect 2490 15370 2510 15390
rect 2510 15370 2515 15390
rect 2485 15365 2515 15370
rect 2565 15390 2595 15395
rect 2565 15370 2570 15390
rect 2570 15370 2590 15390
rect 2590 15370 2595 15390
rect 2565 15365 2595 15370
rect 2645 15390 2675 15395
rect 2645 15370 2650 15390
rect 2650 15370 2670 15390
rect 2670 15370 2675 15390
rect 2645 15365 2675 15370
rect 2725 15390 2755 15395
rect 2725 15370 2730 15390
rect 2730 15370 2750 15390
rect 2750 15370 2755 15390
rect 2725 15365 2755 15370
rect 2805 15390 2835 15395
rect 2805 15370 2810 15390
rect 2810 15370 2830 15390
rect 2830 15370 2835 15390
rect 2805 15365 2835 15370
rect 2885 15390 2915 15395
rect 2885 15370 2890 15390
rect 2890 15370 2910 15390
rect 2910 15370 2915 15390
rect 2885 15365 2915 15370
rect 2965 15390 2995 15395
rect 2965 15370 2970 15390
rect 2970 15370 2990 15390
rect 2990 15370 2995 15390
rect 2965 15365 2995 15370
rect 3045 15390 3075 15395
rect 3045 15370 3050 15390
rect 3050 15370 3070 15390
rect 3070 15370 3075 15390
rect 3045 15365 3075 15370
rect 3125 15390 3155 15395
rect 3125 15370 3130 15390
rect 3130 15370 3150 15390
rect 3150 15370 3155 15390
rect 3125 15365 3155 15370
rect 3205 15390 3235 15395
rect 3205 15370 3210 15390
rect 3210 15370 3230 15390
rect 3230 15370 3235 15390
rect 3205 15365 3235 15370
rect 3285 15390 3315 15395
rect 3285 15370 3290 15390
rect 3290 15370 3310 15390
rect 3310 15370 3315 15390
rect 3285 15365 3315 15370
rect 3365 15390 3395 15395
rect 3365 15370 3370 15390
rect 3370 15370 3390 15390
rect 3390 15370 3395 15390
rect 3365 15365 3395 15370
rect 3445 15390 3475 15395
rect 3445 15370 3450 15390
rect 3450 15370 3470 15390
rect 3470 15370 3475 15390
rect 3445 15365 3475 15370
rect 3525 15390 3555 15395
rect 3525 15370 3530 15390
rect 3530 15370 3550 15390
rect 3550 15370 3555 15390
rect 3525 15365 3555 15370
rect 3605 15390 3635 15395
rect 3605 15370 3610 15390
rect 3610 15370 3630 15390
rect 3630 15370 3635 15390
rect 3605 15365 3635 15370
rect 3685 15390 3715 15395
rect 3685 15370 3690 15390
rect 3690 15370 3710 15390
rect 3710 15370 3715 15390
rect 3685 15365 3715 15370
rect 3765 15390 3795 15395
rect 3765 15370 3770 15390
rect 3770 15370 3790 15390
rect 3790 15370 3795 15390
rect 3765 15365 3795 15370
rect 3845 15390 3875 15395
rect 3845 15370 3850 15390
rect 3850 15370 3870 15390
rect 3870 15370 3875 15390
rect 3845 15365 3875 15370
rect 3925 15390 3955 15395
rect 3925 15370 3930 15390
rect 3930 15370 3950 15390
rect 3950 15370 3955 15390
rect 3925 15365 3955 15370
rect 4005 15390 4035 15395
rect 4005 15370 4010 15390
rect 4010 15370 4030 15390
rect 4030 15370 4035 15390
rect 4005 15365 4035 15370
rect 4085 15390 4115 15395
rect 4085 15370 4090 15390
rect 4090 15370 4110 15390
rect 4110 15370 4115 15390
rect 4085 15365 4115 15370
rect 4165 15390 4195 15395
rect 4165 15370 4170 15390
rect 4170 15370 4190 15390
rect 4190 15370 4195 15390
rect 4165 15365 4195 15370
rect 6245 15390 6275 15395
rect 6245 15370 6250 15390
rect 6250 15370 6270 15390
rect 6270 15370 6275 15390
rect 6245 15365 6275 15370
rect 6325 15390 6355 15395
rect 6325 15370 6330 15390
rect 6330 15370 6350 15390
rect 6350 15370 6355 15390
rect 6325 15365 6355 15370
rect 6405 15390 6435 15395
rect 6405 15370 6410 15390
rect 6410 15370 6430 15390
rect 6430 15370 6435 15390
rect 6405 15365 6435 15370
rect 6485 15390 6515 15395
rect 6485 15370 6490 15390
rect 6490 15370 6510 15390
rect 6510 15370 6515 15390
rect 6485 15365 6515 15370
rect 6565 15390 6595 15395
rect 6565 15370 6570 15390
rect 6570 15370 6590 15390
rect 6590 15370 6595 15390
rect 6565 15365 6595 15370
rect 6645 15390 6675 15395
rect 6645 15370 6650 15390
rect 6650 15370 6670 15390
rect 6670 15370 6675 15390
rect 6645 15365 6675 15370
rect 6725 15390 6755 15395
rect 6725 15370 6730 15390
rect 6730 15370 6750 15390
rect 6750 15370 6755 15390
rect 6725 15365 6755 15370
rect 6805 15390 6835 15395
rect 6805 15370 6810 15390
rect 6810 15370 6830 15390
rect 6830 15370 6835 15390
rect 6805 15365 6835 15370
rect 6885 15390 6915 15395
rect 6885 15370 6890 15390
rect 6890 15370 6910 15390
rect 6910 15370 6915 15390
rect 6885 15365 6915 15370
rect 6965 15390 6995 15395
rect 6965 15370 6970 15390
rect 6970 15370 6990 15390
rect 6990 15370 6995 15390
rect 6965 15365 6995 15370
rect 7045 15390 7075 15395
rect 7045 15370 7050 15390
rect 7050 15370 7070 15390
rect 7070 15370 7075 15390
rect 7045 15365 7075 15370
rect 7125 15390 7155 15395
rect 7125 15370 7130 15390
rect 7130 15370 7150 15390
rect 7150 15370 7155 15390
rect 7125 15365 7155 15370
rect 7205 15390 7235 15395
rect 7205 15370 7210 15390
rect 7210 15370 7230 15390
rect 7230 15370 7235 15390
rect 7205 15365 7235 15370
rect 7285 15390 7315 15395
rect 7285 15370 7290 15390
rect 7290 15370 7310 15390
rect 7310 15370 7315 15390
rect 7285 15365 7315 15370
rect 7365 15390 7395 15395
rect 7365 15370 7370 15390
rect 7370 15370 7390 15390
rect 7390 15370 7395 15390
rect 7365 15365 7395 15370
rect 7445 15390 7475 15395
rect 7445 15370 7450 15390
rect 7450 15370 7470 15390
rect 7470 15370 7475 15390
rect 7445 15365 7475 15370
rect 7525 15390 7555 15395
rect 7525 15370 7530 15390
rect 7530 15370 7550 15390
rect 7550 15370 7555 15390
rect 7525 15365 7555 15370
rect 7605 15390 7635 15395
rect 7605 15370 7610 15390
rect 7610 15370 7630 15390
rect 7630 15370 7635 15390
rect 7605 15365 7635 15370
rect 7685 15390 7715 15395
rect 7685 15370 7690 15390
rect 7690 15370 7710 15390
rect 7710 15370 7715 15390
rect 7685 15365 7715 15370
rect 7765 15390 7795 15395
rect 7765 15370 7770 15390
rect 7770 15370 7790 15390
rect 7790 15370 7795 15390
rect 7765 15365 7795 15370
rect 7845 15390 7875 15395
rect 7845 15370 7850 15390
rect 7850 15370 7870 15390
rect 7870 15370 7875 15390
rect 7845 15365 7875 15370
rect 7925 15390 7955 15395
rect 7925 15370 7930 15390
rect 7930 15370 7950 15390
rect 7950 15370 7955 15390
rect 7925 15365 7955 15370
rect 8005 15390 8035 15395
rect 8005 15370 8010 15390
rect 8010 15370 8030 15390
rect 8030 15370 8035 15390
rect 8005 15365 8035 15370
rect 8085 15390 8115 15395
rect 8085 15370 8090 15390
rect 8090 15370 8110 15390
rect 8110 15370 8115 15390
rect 8085 15365 8115 15370
rect 8165 15390 8195 15395
rect 8165 15370 8170 15390
rect 8170 15370 8190 15390
rect 8190 15370 8195 15390
rect 8165 15365 8195 15370
rect 8245 15390 8275 15395
rect 8245 15370 8250 15390
rect 8250 15370 8270 15390
rect 8270 15370 8275 15390
rect 8245 15365 8275 15370
rect 8325 15390 8355 15395
rect 8325 15370 8330 15390
rect 8330 15370 8350 15390
rect 8350 15370 8355 15390
rect 8325 15365 8355 15370
rect 8405 15390 8435 15395
rect 8405 15370 8410 15390
rect 8410 15370 8430 15390
rect 8430 15370 8435 15390
rect 8405 15365 8435 15370
rect 8485 15390 8515 15395
rect 8485 15370 8490 15390
rect 8490 15370 8510 15390
rect 8510 15370 8515 15390
rect 8485 15365 8515 15370
rect 8565 15390 8595 15395
rect 8565 15370 8570 15390
rect 8570 15370 8590 15390
rect 8590 15370 8595 15390
rect 8565 15365 8595 15370
rect 8645 15390 8675 15395
rect 8645 15370 8650 15390
rect 8650 15370 8670 15390
rect 8670 15370 8675 15390
rect 8645 15365 8675 15370
rect 8725 15390 8755 15395
rect 8725 15370 8730 15390
rect 8730 15370 8750 15390
rect 8750 15370 8755 15390
rect 8725 15365 8755 15370
rect 8805 15390 8835 15395
rect 8805 15370 8810 15390
rect 8810 15370 8830 15390
rect 8830 15370 8835 15390
rect 8805 15365 8835 15370
rect 8885 15390 8915 15395
rect 8885 15370 8890 15390
rect 8890 15370 8910 15390
rect 8910 15370 8915 15390
rect 8885 15365 8915 15370
rect 8965 15390 8995 15395
rect 8965 15370 8970 15390
rect 8970 15370 8990 15390
rect 8990 15370 8995 15390
rect 8965 15365 8995 15370
rect 9045 15390 9075 15395
rect 9045 15370 9050 15390
rect 9050 15370 9070 15390
rect 9070 15370 9075 15390
rect 9045 15365 9075 15370
rect 9125 15390 9155 15395
rect 9125 15370 9130 15390
rect 9130 15370 9150 15390
rect 9150 15370 9155 15390
rect 9125 15365 9155 15370
rect 9205 15390 9235 15395
rect 9205 15370 9210 15390
rect 9210 15370 9230 15390
rect 9230 15370 9235 15390
rect 9205 15365 9235 15370
rect 9285 15390 9315 15395
rect 9285 15370 9290 15390
rect 9290 15370 9310 15390
rect 9310 15370 9315 15390
rect 9285 15365 9315 15370
rect 9365 15390 9395 15395
rect 9365 15370 9370 15390
rect 9370 15370 9390 15390
rect 9390 15370 9395 15390
rect 9365 15365 9395 15370
rect 9445 15390 9475 15395
rect 9445 15370 9450 15390
rect 9450 15370 9470 15390
rect 9470 15370 9475 15390
rect 9445 15365 9475 15370
rect 11565 15390 11595 15395
rect 11565 15370 11570 15390
rect 11570 15370 11590 15390
rect 11590 15370 11595 15390
rect 11565 15365 11595 15370
rect 11645 15390 11675 15395
rect 11645 15370 11650 15390
rect 11650 15370 11670 15390
rect 11670 15370 11675 15390
rect 11645 15365 11675 15370
rect 11725 15390 11755 15395
rect 11725 15370 11730 15390
rect 11730 15370 11750 15390
rect 11750 15370 11755 15390
rect 11725 15365 11755 15370
rect 11805 15390 11835 15395
rect 11805 15370 11810 15390
rect 11810 15370 11830 15390
rect 11830 15370 11835 15390
rect 11805 15365 11835 15370
rect 11885 15390 11915 15395
rect 11885 15370 11890 15390
rect 11890 15370 11910 15390
rect 11910 15370 11915 15390
rect 11885 15365 11915 15370
rect 11965 15390 11995 15395
rect 11965 15370 11970 15390
rect 11970 15370 11990 15390
rect 11990 15370 11995 15390
rect 11965 15365 11995 15370
rect 12045 15390 12075 15395
rect 12045 15370 12050 15390
rect 12050 15370 12070 15390
rect 12070 15370 12075 15390
rect 12045 15365 12075 15370
rect 12125 15390 12155 15395
rect 12125 15370 12130 15390
rect 12130 15370 12150 15390
rect 12150 15370 12155 15390
rect 12125 15365 12155 15370
rect 12205 15390 12235 15395
rect 12205 15370 12210 15390
rect 12210 15370 12230 15390
rect 12230 15370 12235 15390
rect 12205 15365 12235 15370
rect 12285 15390 12315 15395
rect 12285 15370 12290 15390
rect 12290 15370 12310 15390
rect 12310 15370 12315 15390
rect 12285 15365 12315 15370
rect 12365 15390 12395 15395
rect 12365 15370 12370 15390
rect 12370 15370 12390 15390
rect 12390 15370 12395 15390
rect 12365 15365 12395 15370
rect 12445 15390 12475 15395
rect 12445 15370 12450 15390
rect 12450 15370 12470 15390
rect 12470 15370 12475 15390
rect 12445 15365 12475 15370
rect 12525 15390 12555 15395
rect 12525 15370 12530 15390
rect 12530 15370 12550 15390
rect 12550 15370 12555 15390
rect 12525 15365 12555 15370
rect 12605 15390 12635 15395
rect 12605 15370 12610 15390
rect 12610 15370 12630 15390
rect 12630 15370 12635 15390
rect 12605 15365 12635 15370
rect 12685 15390 12715 15395
rect 12685 15370 12690 15390
rect 12690 15370 12710 15390
rect 12710 15370 12715 15390
rect 12685 15365 12715 15370
rect 12765 15390 12795 15395
rect 12765 15370 12770 15390
rect 12770 15370 12790 15390
rect 12790 15370 12795 15390
rect 12765 15365 12795 15370
rect 12845 15390 12875 15395
rect 12845 15370 12850 15390
rect 12850 15370 12870 15390
rect 12870 15370 12875 15390
rect 12845 15365 12875 15370
rect 12925 15390 12955 15395
rect 12925 15370 12930 15390
rect 12930 15370 12950 15390
rect 12950 15370 12955 15390
rect 12925 15365 12955 15370
rect 13005 15390 13035 15395
rect 13005 15370 13010 15390
rect 13010 15370 13030 15390
rect 13030 15370 13035 15390
rect 13005 15365 13035 15370
rect 13085 15390 13115 15395
rect 13085 15370 13090 15390
rect 13090 15370 13110 15390
rect 13110 15370 13115 15390
rect 13085 15365 13115 15370
rect 13165 15390 13195 15395
rect 13165 15370 13170 15390
rect 13170 15370 13190 15390
rect 13190 15370 13195 15390
rect 13165 15365 13195 15370
rect 13245 15390 13275 15395
rect 13245 15370 13250 15390
rect 13250 15370 13270 15390
rect 13270 15370 13275 15390
rect 13245 15365 13275 15370
rect 13325 15390 13355 15395
rect 13325 15370 13330 15390
rect 13330 15370 13350 15390
rect 13350 15370 13355 15390
rect 13325 15365 13355 15370
rect 13405 15390 13435 15395
rect 13405 15370 13410 15390
rect 13410 15370 13430 15390
rect 13430 15370 13435 15390
rect 13405 15365 13435 15370
rect 13485 15390 13515 15395
rect 13485 15370 13490 15390
rect 13490 15370 13510 15390
rect 13510 15370 13515 15390
rect 13485 15365 13515 15370
rect 13565 15390 13595 15395
rect 13565 15370 13570 15390
rect 13570 15370 13590 15390
rect 13590 15370 13595 15390
rect 13565 15365 13595 15370
rect 13645 15390 13675 15395
rect 13645 15370 13650 15390
rect 13650 15370 13670 15390
rect 13670 15370 13675 15390
rect 13645 15365 13675 15370
rect 13725 15390 13755 15395
rect 13725 15370 13730 15390
rect 13730 15370 13750 15390
rect 13750 15370 13755 15390
rect 13725 15365 13755 15370
rect 13805 15390 13835 15395
rect 13805 15370 13810 15390
rect 13810 15370 13830 15390
rect 13830 15370 13835 15390
rect 13805 15365 13835 15370
rect 13885 15390 13915 15395
rect 13885 15370 13890 15390
rect 13890 15370 13910 15390
rect 13910 15370 13915 15390
rect 13885 15365 13915 15370
rect 13965 15390 13995 15395
rect 13965 15370 13970 15390
rect 13970 15370 13990 15390
rect 13990 15370 13995 15390
rect 13965 15365 13995 15370
rect 14045 15390 14075 15395
rect 14045 15370 14050 15390
rect 14050 15370 14070 15390
rect 14070 15370 14075 15390
rect 14045 15365 14075 15370
rect 14125 15390 14155 15395
rect 14125 15370 14130 15390
rect 14130 15370 14150 15390
rect 14150 15370 14155 15390
rect 14125 15365 14155 15370
rect 14205 15390 14235 15395
rect 14205 15370 14210 15390
rect 14210 15370 14230 15390
rect 14230 15370 14235 15390
rect 14205 15365 14235 15370
rect 14285 15390 14315 15395
rect 14285 15370 14290 15390
rect 14290 15370 14310 15390
rect 14310 15370 14315 15390
rect 14285 15365 14315 15370
rect 14365 15390 14395 15395
rect 14365 15370 14370 15390
rect 14370 15370 14390 15390
rect 14390 15370 14395 15390
rect 14365 15365 14395 15370
rect 14445 15390 14475 15395
rect 14445 15370 14450 15390
rect 14450 15370 14470 15390
rect 14470 15370 14475 15390
rect 14445 15365 14475 15370
rect 14525 15390 14555 15395
rect 14525 15370 14530 15390
rect 14530 15370 14550 15390
rect 14550 15370 14555 15390
rect 14525 15365 14555 15370
rect 14605 15390 14635 15395
rect 14605 15370 14610 15390
rect 14610 15370 14630 15390
rect 14630 15370 14635 15390
rect 14605 15365 14635 15370
rect 14685 15390 14715 15395
rect 14685 15370 14690 15390
rect 14690 15370 14710 15390
rect 14710 15370 14715 15390
rect 14685 15365 14715 15370
rect 16765 15390 16795 15395
rect 16765 15370 16770 15390
rect 16770 15370 16790 15390
rect 16790 15370 16795 15390
rect 16765 15365 16795 15370
rect 16845 15390 16875 15395
rect 16845 15370 16850 15390
rect 16850 15370 16870 15390
rect 16870 15370 16875 15390
rect 16845 15365 16875 15370
rect 16925 15390 16955 15395
rect 16925 15370 16930 15390
rect 16930 15370 16950 15390
rect 16950 15370 16955 15390
rect 16925 15365 16955 15370
rect 17005 15390 17035 15395
rect 17005 15370 17010 15390
rect 17010 15370 17030 15390
rect 17030 15370 17035 15390
rect 17005 15365 17035 15370
rect 17085 15390 17115 15395
rect 17085 15370 17090 15390
rect 17090 15370 17110 15390
rect 17110 15370 17115 15390
rect 17085 15365 17115 15370
rect 17165 15390 17195 15395
rect 17165 15370 17170 15390
rect 17170 15370 17190 15390
rect 17190 15370 17195 15390
rect 17165 15365 17195 15370
rect 17245 15390 17275 15395
rect 17245 15370 17250 15390
rect 17250 15370 17270 15390
rect 17270 15370 17275 15390
rect 17245 15365 17275 15370
rect 17325 15390 17355 15395
rect 17325 15370 17330 15390
rect 17330 15370 17350 15390
rect 17350 15370 17355 15390
rect 17325 15365 17355 15370
rect 17405 15390 17435 15395
rect 17405 15370 17410 15390
rect 17410 15370 17430 15390
rect 17430 15370 17435 15390
rect 17405 15365 17435 15370
rect 17485 15390 17515 15395
rect 17485 15370 17490 15390
rect 17490 15370 17510 15390
rect 17510 15370 17515 15390
rect 17485 15365 17515 15370
rect 17565 15390 17595 15395
rect 17565 15370 17570 15390
rect 17570 15370 17590 15390
rect 17590 15370 17595 15390
rect 17565 15365 17595 15370
rect 17645 15390 17675 15395
rect 17645 15370 17650 15390
rect 17650 15370 17670 15390
rect 17670 15370 17675 15390
rect 17645 15365 17675 15370
rect 17725 15390 17755 15395
rect 17725 15370 17730 15390
rect 17730 15370 17750 15390
rect 17750 15370 17755 15390
rect 17725 15365 17755 15370
rect 17805 15390 17835 15395
rect 17805 15370 17810 15390
rect 17810 15370 17830 15390
rect 17830 15370 17835 15390
rect 17805 15365 17835 15370
rect 17885 15390 17915 15395
rect 17885 15370 17890 15390
rect 17890 15370 17910 15390
rect 17910 15370 17915 15390
rect 17885 15365 17915 15370
rect 17965 15390 17995 15395
rect 17965 15370 17970 15390
rect 17970 15370 17990 15390
rect 17990 15370 17995 15390
rect 17965 15365 17995 15370
rect 18045 15390 18075 15395
rect 18045 15370 18050 15390
rect 18050 15370 18070 15390
rect 18070 15370 18075 15390
rect 18045 15365 18075 15370
rect 18125 15390 18155 15395
rect 18125 15370 18130 15390
rect 18130 15370 18150 15390
rect 18150 15370 18155 15390
rect 18125 15365 18155 15370
rect 18205 15390 18235 15395
rect 18205 15370 18210 15390
rect 18210 15370 18230 15390
rect 18230 15370 18235 15390
rect 18205 15365 18235 15370
rect 18285 15390 18315 15395
rect 18285 15370 18290 15390
rect 18290 15370 18310 15390
rect 18310 15370 18315 15390
rect 18285 15365 18315 15370
rect 18365 15390 18395 15395
rect 18365 15370 18370 15390
rect 18370 15370 18390 15390
rect 18390 15370 18395 15390
rect 18365 15365 18395 15370
rect 18445 15390 18475 15395
rect 18445 15370 18450 15390
rect 18450 15370 18470 15390
rect 18470 15370 18475 15390
rect 18445 15365 18475 15370
rect 18525 15390 18555 15395
rect 18525 15370 18530 15390
rect 18530 15370 18550 15390
rect 18550 15370 18555 15390
rect 18525 15365 18555 15370
rect 18605 15390 18635 15395
rect 18605 15370 18610 15390
rect 18610 15370 18630 15390
rect 18630 15370 18635 15390
rect 18605 15365 18635 15370
rect 18685 15390 18715 15395
rect 18685 15370 18690 15390
rect 18690 15370 18710 15390
rect 18710 15370 18715 15390
rect 18685 15365 18715 15370
rect 18765 15390 18795 15395
rect 18765 15370 18770 15390
rect 18770 15370 18790 15390
rect 18790 15370 18795 15390
rect 18765 15365 18795 15370
rect 18845 15390 18875 15395
rect 18845 15370 18850 15390
rect 18850 15370 18870 15390
rect 18870 15370 18875 15390
rect 18845 15365 18875 15370
rect 18925 15390 18955 15395
rect 18925 15370 18930 15390
rect 18930 15370 18950 15390
rect 18950 15370 18955 15390
rect 18925 15365 18955 15370
rect 19005 15390 19035 15395
rect 19005 15370 19010 15390
rect 19010 15370 19030 15390
rect 19030 15370 19035 15390
rect 19005 15365 19035 15370
rect 19085 15390 19115 15395
rect 19085 15370 19090 15390
rect 19090 15370 19110 15390
rect 19110 15370 19115 15390
rect 19085 15365 19115 15370
rect 19165 15390 19195 15395
rect 19165 15370 19170 15390
rect 19170 15370 19190 15390
rect 19190 15370 19195 15390
rect 19165 15365 19195 15370
rect 19245 15390 19275 15395
rect 19245 15370 19250 15390
rect 19250 15370 19270 15390
rect 19270 15370 19275 15390
rect 19245 15365 19275 15370
rect 19325 15390 19355 15395
rect 19325 15370 19330 15390
rect 19330 15370 19350 15390
rect 19350 15370 19355 15390
rect 19325 15365 19355 15370
rect 19405 15390 19435 15395
rect 19405 15370 19410 15390
rect 19410 15370 19430 15390
rect 19430 15370 19435 15390
rect 19405 15365 19435 15370
rect 19485 15390 19515 15395
rect 19485 15370 19490 15390
rect 19490 15370 19510 15390
rect 19510 15370 19515 15390
rect 19485 15365 19515 15370
rect 19565 15390 19595 15395
rect 19565 15370 19570 15390
rect 19570 15370 19590 15390
rect 19590 15370 19595 15390
rect 19565 15365 19595 15370
rect 19645 15390 19675 15395
rect 19645 15370 19650 15390
rect 19650 15370 19670 15390
rect 19670 15370 19675 15390
rect 19645 15365 19675 15370
rect 19725 15390 19755 15395
rect 19725 15370 19730 15390
rect 19730 15370 19750 15390
rect 19750 15370 19755 15390
rect 19725 15365 19755 15370
rect 19805 15390 19835 15395
rect 19805 15370 19810 15390
rect 19810 15370 19830 15390
rect 19830 15370 19835 15390
rect 19805 15365 19835 15370
rect 19885 15390 19915 15395
rect 19885 15370 19890 15390
rect 19890 15370 19910 15390
rect 19910 15370 19915 15390
rect 19885 15365 19915 15370
rect 19965 15390 19995 15395
rect 19965 15370 19970 15390
rect 19970 15370 19990 15390
rect 19990 15370 19995 15390
rect 19965 15365 19995 15370
rect 20045 15390 20075 15395
rect 20045 15370 20050 15390
rect 20050 15370 20070 15390
rect 20070 15370 20075 15390
rect 20045 15365 20075 15370
rect 20125 15390 20155 15395
rect 20125 15370 20130 15390
rect 20130 15370 20150 15390
rect 20150 15370 20155 15390
rect 20125 15365 20155 15370
rect 20205 15390 20235 15395
rect 20205 15370 20210 15390
rect 20210 15370 20230 15390
rect 20230 15370 20235 15390
rect 20205 15365 20235 15370
rect 20285 15390 20315 15395
rect 20285 15370 20290 15390
rect 20290 15370 20310 15390
rect 20310 15370 20315 15390
rect 20285 15365 20315 15370
rect 20365 15390 20395 15395
rect 20365 15370 20370 15390
rect 20370 15370 20390 15390
rect 20390 15370 20395 15390
rect 20365 15365 20395 15370
rect 20445 15390 20475 15395
rect 20445 15370 20450 15390
rect 20450 15370 20470 15390
rect 20470 15370 20475 15390
rect 20445 15365 20475 15370
rect 20525 15390 20555 15395
rect 20525 15370 20530 15390
rect 20530 15370 20550 15390
rect 20550 15370 20555 15390
rect 20525 15365 20555 15370
rect 20605 15390 20635 15395
rect 20605 15370 20610 15390
rect 20610 15370 20630 15390
rect 20630 15370 20635 15390
rect 20605 15365 20635 15370
rect 20685 15390 20715 15395
rect 20685 15370 20690 15390
rect 20690 15370 20710 15390
rect 20710 15370 20715 15390
rect 20685 15365 20715 15370
rect 20765 15390 20795 15395
rect 20765 15370 20770 15390
rect 20770 15370 20790 15390
rect 20790 15370 20795 15390
rect 20765 15365 20795 15370
rect 20845 15390 20875 15395
rect 20845 15370 20850 15390
rect 20850 15370 20870 15390
rect 20870 15370 20875 15390
rect 20845 15365 20875 15370
rect 20925 15390 20955 15395
rect 20925 15370 20930 15390
rect 20930 15370 20950 15390
rect 20950 15370 20955 15390
rect 20925 15365 20955 15370
rect 5 15230 35 15235
rect 5 15210 10 15230
rect 10 15210 30 15230
rect 30 15210 35 15230
rect 5 15205 35 15210
rect 85 15230 115 15235
rect 85 15210 90 15230
rect 90 15210 110 15230
rect 110 15210 115 15230
rect 85 15205 115 15210
rect 165 15230 195 15235
rect 165 15210 170 15230
rect 170 15210 190 15230
rect 190 15210 195 15230
rect 165 15205 195 15210
rect 245 15230 275 15235
rect 245 15210 250 15230
rect 250 15210 270 15230
rect 270 15210 275 15230
rect 245 15205 275 15210
rect 325 15230 355 15235
rect 325 15210 330 15230
rect 330 15210 350 15230
rect 350 15210 355 15230
rect 325 15205 355 15210
rect 405 15230 435 15235
rect 405 15210 410 15230
rect 410 15210 430 15230
rect 430 15210 435 15230
rect 405 15205 435 15210
rect 485 15230 515 15235
rect 485 15210 490 15230
rect 490 15210 510 15230
rect 510 15210 515 15230
rect 485 15205 515 15210
rect 565 15230 595 15235
rect 565 15210 570 15230
rect 570 15210 590 15230
rect 590 15210 595 15230
rect 565 15205 595 15210
rect 645 15230 675 15235
rect 645 15210 650 15230
rect 650 15210 670 15230
rect 670 15210 675 15230
rect 645 15205 675 15210
rect 725 15230 755 15235
rect 725 15210 730 15230
rect 730 15210 750 15230
rect 750 15210 755 15230
rect 725 15205 755 15210
rect 805 15230 835 15235
rect 805 15210 810 15230
rect 810 15210 830 15230
rect 830 15210 835 15230
rect 805 15205 835 15210
rect 885 15230 915 15235
rect 885 15210 890 15230
rect 890 15210 910 15230
rect 910 15210 915 15230
rect 885 15205 915 15210
rect 965 15230 995 15235
rect 965 15210 970 15230
rect 970 15210 990 15230
rect 990 15210 995 15230
rect 965 15205 995 15210
rect 1045 15230 1075 15235
rect 1045 15210 1050 15230
rect 1050 15210 1070 15230
rect 1070 15210 1075 15230
rect 1045 15205 1075 15210
rect 1125 15230 1155 15235
rect 1125 15210 1130 15230
rect 1130 15210 1150 15230
rect 1150 15210 1155 15230
rect 1125 15205 1155 15210
rect 1205 15230 1235 15235
rect 1205 15210 1210 15230
rect 1210 15210 1230 15230
rect 1230 15210 1235 15230
rect 1205 15205 1235 15210
rect 1285 15230 1315 15235
rect 1285 15210 1290 15230
rect 1290 15210 1310 15230
rect 1310 15210 1315 15230
rect 1285 15205 1315 15210
rect 1365 15230 1395 15235
rect 1365 15210 1370 15230
rect 1370 15210 1390 15230
rect 1390 15210 1395 15230
rect 1365 15205 1395 15210
rect 1445 15230 1475 15235
rect 1445 15210 1450 15230
rect 1450 15210 1470 15230
rect 1470 15210 1475 15230
rect 1445 15205 1475 15210
rect 1525 15230 1555 15235
rect 1525 15210 1530 15230
rect 1530 15210 1550 15230
rect 1550 15210 1555 15230
rect 1525 15205 1555 15210
rect 1605 15230 1635 15235
rect 1605 15210 1610 15230
rect 1610 15210 1630 15230
rect 1630 15210 1635 15230
rect 1605 15205 1635 15210
rect 1685 15230 1715 15235
rect 1685 15210 1690 15230
rect 1690 15210 1710 15230
rect 1710 15210 1715 15230
rect 1685 15205 1715 15210
rect 1765 15230 1795 15235
rect 1765 15210 1770 15230
rect 1770 15210 1790 15230
rect 1790 15210 1795 15230
rect 1765 15205 1795 15210
rect 1845 15230 1875 15235
rect 1845 15210 1850 15230
rect 1850 15210 1870 15230
rect 1870 15210 1875 15230
rect 1845 15205 1875 15210
rect 1925 15230 1955 15235
rect 1925 15210 1930 15230
rect 1930 15210 1950 15230
rect 1950 15210 1955 15230
rect 1925 15205 1955 15210
rect 2005 15230 2035 15235
rect 2005 15210 2010 15230
rect 2010 15210 2030 15230
rect 2030 15210 2035 15230
rect 2005 15205 2035 15210
rect 2085 15230 2115 15235
rect 2085 15210 2090 15230
rect 2090 15210 2110 15230
rect 2110 15210 2115 15230
rect 2085 15205 2115 15210
rect 2165 15230 2195 15235
rect 2165 15210 2170 15230
rect 2170 15210 2190 15230
rect 2190 15210 2195 15230
rect 2165 15205 2195 15210
rect 2245 15230 2275 15235
rect 2245 15210 2250 15230
rect 2250 15210 2270 15230
rect 2270 15210 2275 15230
rect 2245 15205 2275 15210
rect 2325 15230 2355 15235
rect 2325 15210 2330 15230
rect 2330 15210 2350 15230
rect 2350 15210 2355 15230
rect 2325 15205 2355 15210
rect 2405 15230 2435 15235
rect 2405 15210 2410 15230
rect 2410 15210 2430 15230
rect 2430 15210 2435 15230
rect 2405 15205 2435 15210
rect 2485 15230 2515 15235
rect 2485 15210 2490 15230
rect 2490 15210 2510 15230
rect 2510 15210 2515 15230
rect 2485 15205 2515 15210
rect 2565 15230 2595 15235
rect 2565 15210 2570 15230
rect 2570 15210 2590 15230
rect 2590 15210 2595 15230
rect 2565 15205 2595 15210
rect 2645 15230 2675 15235
rect 2645 15210 2650 15230
rect 2650 15210 2670 15230
rect 2670 15210 2675 15230
rect 2645 15205 2675 15210
rect 2725 15230 2755 15235
rect 2725 15210 2730 15230
rect 2730 15210 2750 15230
rect 2750 15210 2755 15230
rect 2725 15205 2755 15210
rect 2805 15230 2835 15235
rect 2805 15210 2810 15230
rect 2810 15210 2830 15230
rect 2830 15210 2835 15230
rect 2805 15205 2835 15210
rect 2885 15230 2915 15235
rect 2885 15210 2890 15230
rect 2890 15210 2910 15230
rect 2910 15210 2915 15230
rect 2885 15205 2915 15210
rect 2965 15230 2995 15235
rect 2965 15210 2970 15230
rect 2970 15210 2990 15230
rect 2990 15210 2995 15230
rect 2965 15205 2995 15210
rect 3045 15230 3075 15235
rect 3045 15210 3050 15230
rect 3050 15210 3070 15230
rect 3070 15210 3075 15230
rect 3045 15205 3075 15210
rect 3125 15230 3155 15235
rect 3125 15210 3130 15230
rect 3130 15210 3150 15230
rect 3150 15210 3155 15230
rect 3125 15205 3155 15210
rect 3205 15230 3235 15235
rect 3205 15210 3210 15230
rect 3210 15210 3230 15230
rect 3230 15210 3235 15230
rect 3205 15205 3235 15210
rect 3285 15230 3315 15235
rect 3285 15210 3290 15230
rect 3290 15210 3310 15230
rect 3310 15210 3315 15230
rect 3285 15205 3315 15210
rect 3365 15230 3395 15235
rect 3365 15210 3370 15230
rect 3370 15210 3390 15230
rect 3390 15210 3395 15230
rect 3365 15205 3395 15210
rect 3445 15230 3475 15235
rect 3445 15210 3450 15230
rect 3450 15210 3470 15230
rect 3470 15210 3475 15230
rect 3445 15205 3475 15210
rect 3525 15230 3555 15235
rect 3525 15210 3530 15230
rect 3530 15210 3550 15230
rect 3550 15210 3555 15230
rect 3525 15205 3555 15210
rect 3605 15230 3635 15235
rect 3605 15210 3610 15230
rect 3610 15210 3630 15230
rect 3630 15210 3635 15230
rect 3605 15205 3635 15210
rect 3685 15230 3715 15235
rect 3685 15210 3690 15230
rect 3690 15210 3710 15230
rect 3710 15210 3715 15230
rect 3685 15205 3715 15210
rect 3765 15230 3795 15235
rect 3765 15210 3770 15230
rect 3770 15210 3790 15230
rect 3790 15210 3795 15230
rect 3765 15205 3795 15210
rect 3845 15230 3875 15235
rect 3845 15210 3850 15230
rect 3850 15210 3870 15230
rect 3870 15210 3875 15230
rect 3845 15205 3875 15210
rect 3925 15230 3955 15235
rect 3925 15210 3930 15230
rect 3930 15210 3950 15230
rect 3950 15210 3955 15230
rect 3925 15205 3955 15210
rect 4005 15230 4035 15235
rect 4005 15210 4010 15230
rect 4010 15210 4030 15230
rect 4030 15210 4035 15230
rect 4005 15205 4035 15210
rect 4085 15230 4115 15235
rect 4085 15210 4090 15230
rect 4090 15210 4110 15230
rect 4110 15210 4115 15230
rect 4085 15205 4115 15210
rect 4165 15230 4195 15235
rect 4165 15210 4170 15230
rect 4170 15210 4190 15230
rect 4190 15210 4195 15230
rect 4165 15205 4195 15210
rect 6245 15230 6275 15235
rect 6245 15210 6250 15230
rect 6250 15210 6270 15230
rect 6270 15210 6275 15230
rect 6245 15205 6275 15210
rect 6325 15230 6355 15235
rect 6325 15210 6330 15230
rect 6330 15210 6350 15230
rect 6350 15210 6355 15230
rect 6325 15205 6355 15210
rect 6405 15230 6435 15235
rect 6405 15210 6410 15230
rect 6410 15210 6430 15230
rect 6430 15210 6435 15230
rect 6405 15205 6435 15210
rect 6485 15230 6515 15235
rect 6485 15210 6490 15230
rect 6490 15210 6510 15230
rect 6510 15210 6515 15230
rect 6485 15205 6515 15210
rect 6565 15230 6595 15235
rect 6565 15210 6570 15230
rect 6570 15210 6590 15230
rect 6590 15210 6595 15230
rect 6565 15205 6595 15210
rect 6645 15230 6675 15235
rect 6645 15210 6650 15230
rect 6650 15210 6670 15230
rect 6670 15210 6675 15230
rect 6645 15205 6675 15210
rect 6725 15230 6755 15235
rect 6725 15210 6730 15230
rect 6730 15210 6750 15230
rect 6750 15210 6755 15230
rect 6725 15205 6755 15210
rect 6805 15230 6835 15235
rect 6805 15210 6810 15230
rect 6810 15210 6830 15230
rect 6830 15210 6835 15230
rect 6805 15205 6835 15210
rect 6885 15230 6915 15235
rect 6885 15210 6890 15230
rect 6890 15210 6910 15230
rect 6910 15210 6915 15230
rect 6885 15205 6915 15210
rect 6965 15230 6995 15235
rect 6965 15210 6970 15230
rect 6970 15210 6990 15230
rect 6990 15210 6995 15230
rect 6965 15205 6995 15210
rect 7045 15230 7075 15235
rect 7045 15210 7050 15230
rect 7050 15210 7070 15230
rect 7070 15210 7075 15230
rect 7045 15205 7075 15210
rect 7125 15230 7155 15235
rect 7125 15210 7130 15230
rect 7130 15210 7150 15230
rect 7150 15210 7155 15230
rect 7125 15205 7155 15210
rect 7205 15230 7235 15235
rect 7205 15210 7210 15230
rect 7210 15210 7230 15230
rect 7230 15210 7235 15230
rect 7205 15205 7235 15210
rect 7285 15230 7315 15235
rect 7285 15210 7290 15230
rect 7290 15210 7310 15230
rect 7310 15210 7315 15230
rect 7285 15205 7315 15210
rect 7365 15230 7395 15235
rect 7365 15210 7370 15230
rect 7370 15210 7390 15230
rect 7390 15210 7395 15230
rect 7365 15205 7395 15210
rect 7445 15230 7475 15235
rect 7445 15210 7450 15230
rect 7450 15210 7470 15230
rect 7470 15210 7475 15230
rect 7445 15205 7475 15210
rect 7525 15230 7555 15235
rect 7525 15210 7530 15230
rect 7530 15210 7550 15230
rect 7550 15210 7555 15230
rect 7525 15205 7555 15210
rect 7605 15230 7635 15235
rect 7605 15210 7610 15230
rect 7610 15210 7630 15230
rect 7630 15210 7635 15230
rect 7605 15205 7635 15210
rect 7685 15230 7715 15235
rect 7685 15210 7690 15230
rect 7690 15210 7710 15230
rect 7710 15210 7715 15230
rect 7685 15205 7715 15210
rect 7765 15230 7795 15235
rect 7765 15210 7770 15230
rect 7770 15210 7790 15230
rect 7790 15210 7795 15230
rect 7765 15205 7795 15210
rect 7845 15230 7875 15235
rect 7845 15210 7850 15230
rect 7850 15210 7870 15230
rect 7870 15210 7875 15230
rect 7845 15205 7875 15210
rect 7925 15230 7955 15235
rect 7925 15210 7930 15230
rect 7930 15210 7950 15230
rect 7950 15210 7955 15230
rect 7925 15205 7955 15210
rect 8005 15230 8035 15235
rect 8005 15210 8010 15230
rect 8010 15210 8030 15230
rect 8030 15210 8035 15230
rect 8005 15205 8035 15210
rect 8085 15230 8115 15235
rect 8085 15210 8090 15230
rect 8090 15210 8110 15230
rect 8110 15210 8115 15230
rect 8085 15205 8115 15210
rect 8165 15230 8195 15235
rect 8165 15210 8170 15230
rect 8170 15210 8190 15230
rect 8190 15210 8195 15230
rect 8165 15205 8195 15210
rect 8245 15230 8275 15235
rect 8245 15210 8250 15230
rect 8250 15210 8270 15230
rect 8270 15210 8275 15230
rect 8245 15205 8275 15210
rect 8325 15230 8355 15235
rect 8325 15210 8330 15230
rect 8330 15210 8350 15230
rect 8350 15210 8355 15230
rect 8325 15205 8355 15210
rect 8405 15230 8435 15235
rect 8405 15210 8410 15230
rect 8410 15210 8430 15230
rect 8430 15210 8435 15230
rect 8405 15205 8435 15210
rect 8485 15230 8515 15235
rect 8485 15210 8490 15230
rect 8490 15210 8510 15230
rect 8510 15210 8515 15230
rect 8485 15205 8515 15210
rect 8565 15230 8595 15235
rect 8565 15210 8570 15230
rect 8570 15210 8590 15230
rect 8590 15210 8595 15230
rect 8565 15205 8595 15210
rect 8645 15230 8675 15235
rect 8645 15210 8650 15230
rect 8650 15210 8670 15230
rect 8670 15210 8675 15230
rect 8645 15205 8675 15210
rect 8725 15230 8755 15235
rect 8725 15210 8730 15230
rect 8730 15210 8750 15230
rect 8750 15210 8755 15230
rect 8725 15205 8755 15210
rect 8805 15230 8835 15235
rect 8805 15210 8810 15230
rect 8810 15210 8830 15230
rect 8830 15210 8835 15230
rect 8805 15205 8835 15210
rect 8885 15230 8915 15235
rect 8885 15210 8890 15230
rect 8890 15210 8910 15230
rect 8910 15210 8915 15230
rect 8885 15205 8915 15210
rect 8965 15230 8995 15235
rect 8965 15210 8970 15230
rect 8970 15210 8990 15230
rect 8990 15210 8995 15230
rect 8965 15205 8995 15210
rect 9045 15230 9075 15235
rect 9045 15210 9050 15230
rect 9050 15210 9070 15230
rect 9070 15210 9075 15230
rect 9045 15205 9075 15210
rect 9125 15230 9155 15235
rect 9125 15210 9130 15230
rect 9130 15210 9150 15230
rect 9150 15210 9155 15230
rect 9125 15205 9155 15210
rect 9205 15230 9235 15235
rect 9205 15210 9210 15230
rect 9210 15210 9230 15230
rect 9230 15210 9235 15230
rect 9205 15205 9235 15210
rect 9285 15230 9315 15235
rect 9285 15210 9290 15230
rect 9290 15210 9310 15230
rect 9310 15210 9315 15230
rect 9285 15205 9315 15210
rect 9365 15230 9395 15235
rect 9365 15210 9370 15230
rect 9370 15210 9390 15230
rect 9390 15210 9395 15230
rect 9365 15205 9395 15210
rect 9445 15230 9475 15235
rect 9445 15210 9450 15230
rect 9450 15210 9470 15230
rect 9470 15210 9475 15230
rect 9445 15205 9475 15210
rect 11565 15230 11595 15235
rect 11565 15210 11570 15230
rect 11570 15210 11590 15230
rect 11590 15210 11595 15230
rect 11565 15205 11595 15210
rect 11645 15230 11675 15235
rect 11645 15210 11650 15230
rect 11650 15210 11670 15230
rect 11670 15210 11675 15230
rect 11645 15205 11675 15210
rect 11725 15230 11755 15235
rect 11725 15210 11730 15230
rect 11730 15210 11750 15230
rect 11750 15210 11755 15230
rect 11725 15205 11755 15210
rect 11805 15230 11835 15235
rect 11805 15210 11810 15230
rect 11810 15210 11830 15230
rect 11830 15210 11835 15230
rect 11805 15205 11835 15210
rect 11885 15230 11915 15235
rect 11885 15210 11890 15230
rect 11890 15210 11910 15230
rect 11910 15210 11915 15230
rect 11885 15205 11915 15210
rect 11965 15230 11995 15235
rect 11965 15210 11970 15230
rect 11970 15210 11990 15230
rect 11990 15210 11995 15230
rect 11965 15205 11995 15210
rect 12045 15230 12075 15235
rect 12045 15210 12050 15230
rect 12050 15210 12070 15230
rect 12070 15210 12075 15230
rect 12045 15205 12075 15210
rect 12125 15230 12155 15235
rect 12125 15210 12130 15230
rect 12130 15210 12150 15230
rect 12150 15210 12155 15230
rect 12125 15205 12155 15210
rect 12205 15230 12235 15235
rect 12205 15210 12210 15230
rect 12210 15210 12230 15230
rect 12230 15210 12235 15230
rect 12205 15205 12235 15210
rect 12285 15230 12315 15235
rect 12285 15210 12290 15230
rect 12290 15210 12310 15230
rect 12310 15210 12315 15230
rect 12285 15205 12315 15210
rect 12365 15230 12395 15235
rect 12365 15210 12370 15230
rect 12370 15210 12390 15230
rect 12390 15210 12395 15230
rect 12365 15205 12395 15210
rect 12445 15230 12475 15235
rect 12445 15210 12450 15230
rect 12450 15210 12470 15230
rect 12470 15210 12475 15230
rect 12445 15205 12475 15210
rect 12525 15230 12555 15235
rect 12525 15210 12530 15230
rect 12530 15210 12550 15230
rect 12550 15210 12555 15230
rect 12525 15205 12555 15210
rect 12605 15230 12635 15235
rect 12605 15210 12610 15230
rect 12610 15210 12630 15230
rect 12630 15210 12635 15230
rect 12605 15205 12635 15210
rect 12685 15230 12715 15235
rect 12685 15210 12690 15230
rect 12690 15210 12710 15230
rect 12710 15210 12715 15230
rect 12685 15205 12715 15210
rect 12765 15230 12795 15235
rect 12765 15210 12770 15230
rect 12770 15210 12790 15230
rect 12790 15210 12795 15230
rect 12765 15205 12795 15210
rect 12845 15230 12875 15235
rect 12845 15210 12850 15230
rect 12850 15210 12870 15230
rect 12870 15210 12875 15230
rect 12845 15205 12875 15210
rect 12925 15230 12955 15235
rect 12925 15210 12930 15230
rect 12930 15210 12950 15230
rect 12950 15210 12955 15230
rect 12925 15205 12955 15210
rect 13005 15230 13035 15235
rect 13005 15210 13010 15230
rect 13010 15210 13030 15230
rect 13030 15210 13035 15230
rect 13005 15205 13035 15210
rect 13085 15230 13115 15235
rect 13085 15210 13090 15230
rect 13090 15210 13110 15230
rect 13110 15210 13115 15230
rect 13085 15205 13115 15210
rect 13165 15230 13195 15235
rect 13165 15210 13170 15230
rect 13170 15210 13190 15230
rect 13190 15210 13195 15230
rect 13165 15205 13195 15210
rect 13245 15230 13275 15235
rect 13245 15210 13250 15230
rect 13250 15210 13270 15230
rect 13270 15210 13275 15230
rect 13245 15205 13275 15210
rect 13325 15230 13355 15235
rect 13325 15210 13330 15230
rect 13330 15210 13350 15230
rect 13350 15210 13355 15230
rect 13325 15205 13355 15210
rect 13405 15230 13435 15235
rect 13405 15210 13410 15230
rect 13410 15210 13430 15230
rect 13430 15210 13435 15230
rect 13405 15205 13435 15210
rect 13485 15230 13515 15235
rect 13485 15210 13490 15230
rect 13490 15210 13510 15230
rect 13510 15210 13515 15230
rect 13485 15205 13515 15210
rect 13565 15230 13595 15235
rect 13565 15210 13570 15230
rect 13570 15210 13590 15230
rect 13590 15210 13595 15230
rect 13565 15205 13595 15210
rect 13645 15230 13675 15235
rect 13645 15210 13650 15230
rect 13650 15210 13670 15230
rect 13670 15210 13675 15230
rect 13645 15205 13675 15210
rect 13725 15230 13755 15235
rect 13725 15210 13730 15230
rect 13730 15210 13750 15230
rect 13750 15210 13755 15230
rect 13725 15205 13755 15210
rect 13805 15230 13835 15235
rect 13805 15210 13810 15230
rect 13810 15210 13830 15230
rect 13830 15210 13835 15230
rect 13805 15205 13835 15210
rect 13885 15230 13915 15235
rect 13885 15210 13890 15230
rect 13890 15210 13910 15230
rect 13910 15210 13915 15230
rect 13885 15205 13915 15210
rect 13965 15230 13995 15235
rect 13965 15210 13970 15230
rect 13970 15210 13990 15230
rect 13990 15210 13995 15230
rect 13965 15205 13995 15210
rect 14045 15230 14075 15235
rect 14045 15210 14050 15230
rect 14050 15210 14070 15230
rect 14070 15210 14075 15230
rect 14045 15205 14075 15210
rect 14125 15230 14155 15235
rect 14125 15210 14130 15230
rect 14130 15210 14150 15230
rect 14150 15210 14155 15230
rect 14125 15205 14155 15210
rect 14205 15230 14235 15235
rect 14205 15210 14210 15230
rect 14210 15210 14230 15230
rect 14230 15210 14235 15230
rect 14205 15205 14235 15210
rect 14285 15230 14315 15235
rect 14285 15210 14290 15230
rect 14290 15210 14310 15230
rect 14310 15210 14315 15230
rect 14285 15205 14315 15210
rect 14365 15230 14395 15235
rect 14365 15210 14370 15230
rect 14370 15210 14390 15230
rect 14390 15210 14395 15230
rect 14365 15205 14395 15210
rect 14445 15230 14475 15235
rect 14445 15210 14450 15230
rect 14450 15210 14470 15230
rect 14470 15210 14475 15230
rect 14445 15205 14475 15210
rect 14525 15230 14555 15235
rect 14525 15210 14530 15230
rect 14530 15210 14550 15230
rect 14550 15210 14555 15230
rect 14525 15205 14555 15210
rect 14605 15230 14635 15235
rect 14605 15210 14610 15230
rect 14610 15210 14630 15230
rect 14630 15210 14635 15230
rect 14605 15205 14635 15210
rect 14685 15230 14715 15235
rect 14685 15210 14690 15230
rect 14690 15210 14710 15230
rect 14710 15210 14715 15230
rect 14685 15205 14715 15210
rect 16765 15230 16795 15235
rect 16765 15210 16770 15230
rect 16770 15210 16790 15230
rect 16790 15210 16795 15230
rect 16765 15205 16795 15210
rect 16845 15230 16875 15235
rect 16845 15210 16850 15230
rect 16850 15210 16870 15230
rect 16870 15210 16875 15230
rect 16845 15205 16875 15210
rect 16925 15230 16955 15235
rect 16925 15210 16930 15230
rect 16930 15210 16950 15230
rect 16950 15210 16955 15230
rect 16925 15205 16955 15210
rect 17005 15230 17035 15235
rect 17005 15210 17010 15230
rect 17010 15210 17030 15230
rect 17030 15210 17035 15230
rect 17005 15205 17035 15210
rect 17085 15230 17115 15235
rect 17085 15210 17090 15230
rect 17090 15210 17110 15230
rect 17110 15210 17115 15230
rect 17085 15205 17115 15210
rect 17165 15230 17195 15235
rect 17165 15210 17170 15230
rect 17170 15210 17190 15230
rect 17190 15210 17195 15230
rect 17165 15205 17195 15210
rect 17245 15230 17275 15235
rect 17245 15210 17250 15230
rect 17250 15210 17270 15230
rect 17270 15210 17275 15230
rect 17245 15205 17275 15210
rect 17325 15230 17355 15235
rect 17325 15210 17330 15230
rect 17330 15210 17350 15230
rect 17350 15210 17355 15230
rect 17325 15205 17355 15210
rect 17405 15230 17435 15235
rect 17405 15210 17410 15230
rect 17410 15210 17430 15230
rect 17430 15210 17435 15230
rect 17405 15205 17435 15210
rect 17485 15230 17515 15235
rect 17485 15210 17490 15230
rect 17490 15210 17510 15230
rect 17510 15210 17515 15230
rect 17485 15205 17515 15210
rect 17565 15230 17595 15235
rect 17565 15210 17570 15230
rect 17570 15210 17590 15230
rect 17590 15210 17595 15230
rect 17565 15205 17595 15210
rect 17645 15230 17675 15235
rect 17645 15210 17650 15230
rect 17650 15210 17670 15230
rect 17670 15210 17675 15230
rect 17645 15205 17675 15210
rect 17725 15230 17755 15235
rect 17725 15210 17730 15230
rect 17730 15210 17750 15230
rect 17750 15210 17755 15230
rect 17725 15205 17755 15210
rect 17805 15230 17835 15235
rect 17805 15210 17810 15230
rect 17810 15210 17830 15230
rect 17830 15210 17835 15230
rect 17805 15205 17835 15210
rect 17885 15230 17915 15235
rect 17885 15210 17890 15230
rect 17890 15210 17910 15230
rect 17910 15210 17915 15230
rect 17885 15205 17915 15210
rect 17965 15230 17995 15235
rect 17965 15210 17970 15230
rect 17970 15210 17990 15230
rect 17990 15210 17995 15230
rect 17965 15205 17995 15210
rect 18045 15230 18075 15235
rect 18045 15210 18050 15230
rect 18050 15210 18070 15230
rect 18070 15210 18075 15230
rect 18045 15205 18075 15210
rect 18125 15230 18155 15235
rect 18125 15210 18130 15230
rect 18130 15210 18150 15230
rect 18150 15210 18155 15230
rect 18125 15205 18155 15210
rect 18205 15230 18235 15235
rect 18205 15210 18210 15230
rect 18210 15210 18230 15230
rect 18230 15210 18235 15230
rect 18205 15205 18235 15210
rect 18285 15230 18315 15235
rect 18285 15210 18290 15230
rect 18290 15210 18310 15230
rect 18310 15210 18315 15230
rect 18285 15205 18315 15210
rect 18365 15230 18395 15235
rect 18365 15210 18370 15230
rect 18370 15210 18390 15230
rect 18390 15210 18395 15230
rect 18365 15205 18395 15210
rect 18445 15230 18475 15235
rect 18445 15210 18450 15230
rect 18450 15210 18470 15230
rect 18470 15210 18475 15230
rect 18445 15205 18475 15210
rect 18525 15230 18555 15235
rect 18525 15210 18530 15230
rect 18530 15210 18550 15230
rect 18550 15210 18555 15230
rect 18525 15205 18555 15210
rect 18605 15230 18635 15235
rect 18605 15210 18610 15230
rect 18610 15210 18630 15230
rect 18630 15210 18635 15230
rect 18605 15205 18635 15210
rect 18685 15230 18715 15235
rect 18685 15210 18690 15230
rect 18690 15210 18710 15230
rect 18710 15210 18715 15230
rect 18685 15205 18715 15210
rect 18765 15230 18795 15235
rect 18765 15210 18770 15230
rect 18770 15210 18790 15230
rect 18790 15210 18795 15230
rect 18765 15205 18795 15210
rect 18845 15230 18875 15235
rect 18845 15210 18850 15230
rect 18850 15210 18870 15230
rect 18870 15210 18875 15230
rect 18845 15205 18875 15210
rect 18925 15230 18955 15235
rect 18925 15210 18930 15230
rect 18930 15210 18950 15230
rect 18950 15210 18955 15230
rect 18925 15205 18955 15210
rect 19005 15230 19035 15235
rect 19005 15210 19010 15230
rect 19010 15210 19030 15230
rect 19030 15210 19035 15230
rect 19005 15205 19035 15210
rect 19085 15230 19115 15235
rect 19085 15210 19090 15230
rect 19090 15210 19110 15230
rect 19110 15210 19115 15230
rect 19085 15205 19115 15210
rect 19165 15230 19195 15235
rect 19165 15210 19170 15230
rect 19170 15210 19190 15230
rect 19190 15210 19195 15230
rect 19165 15205 19195 15210
rect 19245 15230 19275 15235
rect 19245 15210 19250 15230
rect 19250 15210 19270 15230
rect 19270 15210 19275 15230
rect 19245 15205 19275 15210
rect 19325 15230 19355 15235
rect 19325 15210 19330 15230
rect 19330 15210 19350 15230
rect 19350 15210 19355 15230
rect 19325 15205 19355 15210
rect 19405 15230 19435 15235
rect 19405 15210 19410 15230
rect 19410 15210 19430 15230
rect 19430 15210 19435 15230
rect 19405 15205 19435 15210
rect 19485 15230 19515 15235
rect 19485 15210 19490 15230
rect 19490 15210 19510 15230
rect 19510 15210 19515 15230
rect 19485 15205 19515 15210
rect 19565 15230 19595 15235
rect 19565 15210 19570 15230
rect 19570 15210 19590 15230
rect 19590 15210 19595 15230
rect 19565 15205 19595 15210
rect 19645 15230 19675 15235
rect 19645 15210 19650 15230
rect 19650 15210 19670 15230
rect 19670 15210 19675 15230
rect 19645 15205 19675 15210
rect 19725 15230 19755 15235
rect 19725 15210 19730 15230
rect 19730 15210 19750 15230
rect 19750 15210 19755 15230
rect 19725 15205 19755 15210
rect 19805 15230 19835 15235
rect 19805 15210 19810 15230
rect 19810 15210 19830 15230
rect 19830 15210 19835 15230
rect 19805 15205 19835 15210
rect 19885 15230 19915 15235
rect 19885 15210 19890 15230
rect 19890 15210 19910 15230
rect 19910 15210 19915 15230
rect 19885 15205 19915 15210
rect 19965 15230 19995 15235
rect 19965 15210 19970 15230
rect 19970 15210 19990 15230
rect 19990 15210 19995 15230
rect 19965 15205 19995 15210
rect 20045 15230 20075 15235
rect 20045 15210 20050 15230
rect 20050 15210 20070 15230
rect 20070 15210 20075 15230
rect 20045 15205 20075 15210
rect 20125 15230 20155 15235
rect 20125 15210 20130 15230
rect 20130 15210 20150 15230
rect 20150 15210 20155 15230
rect 20125 15205 20155 15210
rect 20205 15230 20235 15235
rect 20205 15210 20210 15230
rect 20210 15210 20230 15230
rect 20230 15210 20235 15230
rect 20205 15205 20235 15210
rect 20285 15230 20315 15235
rect 20285 15210 20290 15230
rect 20290 15210 20310 15230
rect 20310 15210 20315 15230
rect 20285 15205 20315 15210
rect 20365 15230 20395 15235
rect 20365 15210 20370 15230
rect 20370 15210 20390 15230
rect 20390 15210 20395 15230
rect 20365 15205 20395 15210
rect 20445 15230 20475 15235
rect 20445 15210 20450 15230
rect 20450 15210 20470 15230
rect 20470 15210 20475 15230
rect 20445 15205 20475 15210
rect 20525 15230 20555 15235
rect 20525 15210 20530 15230
rect 20530 15210 20550 15230
rect 20550 15210 20555 15230
rect 20525 15205 20555 15210
rect 20605 15230 20635 15235
rect 20605 15210 20610 15230
rect 20610 15210 20630 15230
rect 20630 15210 20635 15230
rect 20605 15205 20635 15210
rect 20685 15230 20715 15235
rect 20685 15210 20690 15230
rect 20690 15210 20710 15230
rect 20710 15210 20715 15230
rect 20685 15205 20715 15210
rect 20765 15230 20795 15235
rect 20765 15210 20770 15230
rect 20770 15210 20790 15230
rect 20790 15210 20795 15230
rect 20765 15205 20795 15210
rect 20845 15230 20875 15235
rect 20845 15210 20850 15230
rect 20850 15210 20870 15230
rect 20870 15210 20875 15230
rect 20845 15205 20875 15210
rect 20925 15230 20955 15235
rect 20925 15210 20930 15230
rect 20930 15210 20950 15230
rect 20950 15210 20955 15230
rect 20925 15205 20955 15210
rect 5 15150 35 15155
rect 5 15130 10 15150
rect 10 15130 30 15150
rect 30 15130 35 15150
rect 5 15125 35 15130
rect 85 15150 115 15155
rect 85 15130 90 15150
rect 90 15130 110 15150
rect 110 15130 115 15150
rect 85 15125 115 15130
rect 165 15150 195 15155
rect 165 15130 170 15150
rect 170 15130 190 15150
rect 190 15130 195 15150
rect 165 15125 195 15130
rect 245 15150 275 15155
rect 245 15130 250 15150
rect 250 15130 270 15150
rect 270 15130 275 15150
rect 245 15125 275 15130
rect 325 15150 355 15155
rect 325 15130 330 15150
rect 330 15130 350 15150
rect 350 15130 355 15150
rect 325 15125 355 15130
rect 405 15150 435 15155
rect 405 15130 410 15150
rect 410 15130 430 15150
rect 430 15130 435 15150
rect 405 15125 435 15130
rect 485 15150 515 15155
rect 485 15130 490 15150
rect 490 15130 510 15150
rect 510 15130 515 15150
rect 485 15125 515 15130
rect 565 15150 595 15155
rect 565 15130 570 15150
rect 570 15130 590 15150
rect 590 15130 595 15150
rect 565 15125 595 15130
rect 645 15150 675 15155
rect 645 15130 650 15150
rect 650 15130 670 15150
rect 670 15130 675 15150
rect 645 15125 675 15130
rect 725 15150 755 15155
rect 725 15130 730 15150
rect 730 15130 750 15150
rect 750 15130 755 15150
rect 725 15125 755 15130
rect 805 15150 835 15155
rect 805 15130 810 15150
rect 810 15130 830 15150
rect 830 15130 835 15150
rect 805 15125 835 15130
rect 885 15150 915 15155
rect 885 15130 890 15150
rect 890 15130 910 15150
rect 910 15130 915 15150
rect 885 15125 915 15130
rect 965 15150 995 15155
rect 965 15130 970 15150
rect 970 15130 990 15150
rect 990 15130 995 15150
rect 965 15125 995 15130
rect 1045 15150 1075 15155
rect 1045 15130 1050 15150
rect 1050 15130 1070 15150
rect 1070 15130 1075 15150
rect 1045 15125 1075 15130
rect 1125 15150 1155 15155
rect 1125 15130 1130 15150
rect 1130 15130 1150 15150
rect 1150 15130 1155 15150
rect 1125 15125 1155 15130
rect 1205 15150 1235 15155
rect 1205 15130 1210 15150
rect 1210 15130 1230 15150
rect 1230 15130 1235 15150
rect 1205 15125 1235 15130
rect 1285 15150 1315 15155
rect 1285 15130 1290 15150
rect 1290 15130 1310 15150
rect 1310 15130 1315 15150
rect 1285 15125 1315 15130
rect 1365 15150 1395 15155
rect 1365 15130 1370 15150
rect 1370 15130 1390 15150
rect 1390 15130 1395 15150
rect 1365 15125 1395 15130
rect 1445 15150 1475 15155
rect 1445 15130 1450 15150
rect 1450 15130 1470 15150
rect 1470 15130 1475 15150
rect 1445 15125 1475 15130
rect 1525 15150 1555 15155
rect 1525 15130 1530 15150
rect 1530 15130 1550 15150
rect 1550 15130 1555 15150
rect 1525 15125 1555 15130
rect 1605 15150 1635 15155
rect 1605 15130 1610 15150
rect 1610 15130 1630 15150
rect 1630 15130 1635 15150
rect 1605 15125 1635 15130
rect 1685 15150 1715 15155
rect 1685 15130 1690 15150
rect 1690 15130 1710 15150
rect 1710 15130 1715 15150
rect 1685 15125 1715 15130
rect 1765 15150 1795 15155
rect 1765 15130 1770 15150
rect 1770 15130 1790 15150
rect 1790 15130 1795 15150
rect 1765 15125 1795 15130
rect 1845 15150 1875 15155
rect 1845 15130 1850 15150
rect 1850 15130 1870 15150
rect 1870 15130 1875 15150
rect 1845 15125 1875 15130
rect 1925 15150 1955 15155
rect 1925 15130 1930 15150
rect 1930 15130 1950 15150
rect 1950 15130 1955 15150
rect 1925 15125 1955 15130
rect 2005 15150 2035 15155
rect 2005 15130 2010 15150
rect 2010 15130 2030 15150
rect 2030 15130 2035 15150
rect 2005 15125 2035 15130
rect 2085 15150 2115 15155
rect 2085 15130 2090 15150
rect 2090 15130 2110 15150
rect 2110 15130 2115 15150
rect 2085 15125 2115 15130
rect 2165 15150 2195 15155
rect 2165 15130 2170 15150
rect 2170 15130 2190 15150
rect 2190 15130 2195 15150
rect 2165 15125 2195 15130
rect 2245 15150 2275 15155
rect 2245 15130 2250 15150
rect 2250 15130 2270 15150
rect 2270 15130 2275 15150
rect 2245 15125 2275 15130
rect 2325 15150 2355 15155
rect 2325 15130 2330 15150
rect 2330 15130 2350 15150
rect 2350 15130 2355 15150
rect 2325 15125 2355 15130
rect 2405 15150 2435 15155
rect 2405 15130 2410 15150
rect 2410 15130 2430 15150
rect 2430 15130 2435 15150
rect 2405 15125 2435 15130
rect 2485 15150 2515 15155
rect 2485 15130 2490 15150
rect 2490 15130 2510 15150
rect 2510 15130 2515 15150
rect 2485 15125 2515 15130
rect 2565 15150 2595 15155
rect 2565 15130 2570 15150
rect 2570 15130 2590 15150
rect 2590 15130 2595 15150
rect 2565 15125 2595 15130
rect 2645 15150 2675 15155
rect 2645 15130 2650 15150
rect 2650 15130 2670 15150
rect 2670 15130 2675 15150
rect 2645 15125 2675 15130
rect 2725 15150 2755 15155
rect 2725 15130 2730 15150
rect 2730 15130 2750 15150
rect 2750 15130 2755 15150
rect 2725 15125 2755 15130
rect 2805 15150 2835 15155
rect 2805 15130 2810 15150
rect 2810 15130 2830 15150
rect 2830 15130 2835 15150
rect 2805 15125 2835 15130
rect 2885 15150 2915 15155
rect 2885 15130 2890 15150
rect 2890 15130 2910 15150
rect 2910 15130 2915 15150
rect 2885 15125 2915 15130
rect 2965 15150 2995 15155
rect 2965 15130 2970 15150
rect 2970 15130 2990 15150
rect 2990 15130 2995 15150
rect 2965 15125 2995 15130
rect 3045 15150 3075 15155
rect 3045 15130 3050 15150
rect 3050 15130 3070 15150
rect 3070 15130 3075 15150
rect 3045 15125 3075 15130
rect 3125 15150 3155 15155
rect 3125 15130 3130 15150
rect 3130 15130 3150 15150
rect 3150 15130 3155 15150
rect 3125 15125 3155 15130
rect 3205 15150 3235 15155
rect 3205 15130 3210 15150
rect 3210 15130 3230 15150
rect 3230 15130 3235 15150
rect 3205 15125 3235 15130
rect 3285 15150 3315 15155
rect 3285 15130 3290 15150
rect 3290 15130 3310 15150
rect 3310 15130 3315 15150
rect 3285 15125 3315 15130
rect 3365 15150 3395 15155
rect 3365 15130 3370 15150
rect 3370 15130 3390 15150
rect 3390 15130 3395 15150
rect 3365 15125 3395 15130
rect 3445 15150 3475 15155
rect 3445 15130 3450 15150
rect 3450 15130 3470 15150
rect 3470 15130 3475 15150
rect 3445 15125 3475 15130
rect 3525 15150 3555 15155
rect 3525 15130 3530 15150
rect 3530 15130 3550 15150
rect 3550 15130 3555 15150
rect 3525 15125 3555 15130
rect 3605 15150 3635 15155
rect 3605 15130 3610 15150
rect 3610 15130 3630 15150
rect 3630 15130 3635 15150
rect 3605 15125 3635 15130
rect 3685 15150 3715 15155
rect 3685 15130 3690 15150
rect 3690 15130 3710 15150
rect 3710 15130 3715 15150
rect 3685 15125 3715 15130
rect 3765 15150 3795 15155
rect 3765 15130 3770 15150
rect 3770 15130 3790 15150
rect 3790 15130 3795 15150
rect 3765 15125 3795 15130
rect 3845 15150 3875 15155
rect 3845 15130 3850 15150
rect 3850 15130 3870 15150
rect 3870 15130 3875 15150
rect 3845 15125 3875 15130
rect 3925 15150 3955 15155
rect 3925 15130 3930 15150
rect 3930 15130 3950 15150
rect 3950 15130 3955 15150
rect 3925 15125 3955 15130
rect 4005 15150 4035 15155
rect 4005 15130 4010 15150
rect 4010 15130 4030 15150
rect 4030 15130 4035 15150
rect 4005 15125 4035 15130
rect 4085 15150 4115 15155
rect 4085 15130 4090 15150
rect 4090 15130 4110 15150
rect 4110 15130 4115 15150
rect 4085 15125 4115 15130
rect 4165 15150 4195 15155
rect 4165 15130 4170 15150
rect 4170 15130 4190 15150
rect 4190 15130 4195 15150
rect 4165 15125 4195 15130
rect 6245 15150 6275 15155
rect 6245 15130 6250 15150
rect 6250 15130 6270 15150
rect 6270 15130 6275 15150
rect 6245 15125 6275 15130
rect 6325 15150 6355 15155
rect 6325 15130 6330 15150
rect 6330 15130 6350 15150
rect 6350 15130 6355 15150
rect 6325 15125 6355 15130
rect 6405 15150 6435 15155
rect 6405 15130 6410 15150
rect 6410 15130 6430 15150
rect 6430 15130 6435 15150
rect 6405 15125 6435 15130
rect 6485 15150 6515 15155
rect 6485 15130 6490 15150
rect 6490 15130 6510 15150
rect 6510 15130 6515 15150
rect 6485 15125 6515 15130
rect 6565 15150 6595 15155
rect 6565 15130 6570 15150
rect 6570 15130 6590 15150
rect 6590 15130 6595 15150
rect 6565 15125 6595 15130
rect 6645 15150 6675 15155
rect 6645 15130 6650 15150
rect 6650 15130 6670 15150
rect 6670 15130 6675 15150
rect 6645 15125 6675 15130
rect 6725 15150 6755 15155
rect 6725 15130 6730 15150
rect 6730 15130 6750 15150
rect 6750 15130 6755 15150
rect 6725 15125 6755 15130
rect 6805 15150 6835 15155
rect 6805 15130 6810 15150
rect 6810 15130 6830 15150
rect 6830 15130 6835 15150
rect 6805 15125 6835 15130
rect 6885 15150 6915 15155
rect 6885 15130 6890 15150
rect 6890 15130 6910 15150
rect 6910 15130 6915 15150
rect 6885 15125 6915 15130
rect 6965 15150 6995 15155
rect 6965 15130 6970 15150
rect 6970 15130 6990 15150
rect 6990 15130 6995 15150
rect 6965 15125 6995 15130
rect 7045 15150 7075 15155
rect 7045 15130 7050 15150
rect 7050 15130 7070 15150
rect 7070 15130 7075 15150
rect 7045 15125 7075 15130
rect 7125 15150 7155 15155
rect 7125 15130 7130 15150
rect 7130 15130 7150 15150
rect 7150 15130 7155 15150
rect 7125 15125 7155 15130
rect 7205 15150 7235 15155
rect 7205 15130 7210 15150
rect 7210 15130 7230 15150
rect 7230 15130 7235 15150
rect 7205 15125 7235 15130
rect 7285 15150 7315 15155
rect 7285 15130 7290 15150
rect 7290 15130 7310 15150
rect 7310 15130 7315 15150
rect 7285 15125 7315 15130
rect 7365 15150 7395 15155
rect 7365 15130 7370 15150
rect 7370 15130 7390 15150
rect 7390 15130 7395 15150
rect 7365 15125 7395 15130
rect 7445 15150 7475 15155
rect 7445 15130 7450 15150
rect 7450 15130 7470 15150
rect 7470 15130 7475 15150
rect 7445 15125 7475 15130
rect 7525 15150 7555 15155
rect 7525 15130 7530 15150
rect 7530 15130 7550 15150
rect 7550 15130 7555 15150
rect 7525 15125 7555 15130
rect 7605 15150 7635 15155
rect 7605 15130 7610 15150
rect 7610 15130 7630 15150
rect 7630 15130 7635 15150
rect 7605 15125 7635 15130
rect 7685 15150 7715 15155
rect 7685 15130 7690 15150
rect 7690 15130 7710 15150
rect 7710 15130 7715 15150
rect 7685 15125 7715 15130
rect 7765 15150 7795 15155
rect 7765 15130 7770 15150
rect 7770 15130 7790 15150
rect 7790 15130 7795 15150
rect 7765 15125 7795 15130
rect 7845 15150 7875 15155
rect 7845 15130 7850 15150
rect 7850 15130 7870 15150
rect 7870 15130 7875 15150
rect 7845 15125 7875 15130
rect 7925 15150 7955 15155
rect 7925 15130 7930 15150
rect 7930 15130 7950 15150
rect 7950 15130 7955 15150
rect 7925 15125 7955 15130
rect 8005 15150 8035 15155
rect 8005 15130 8010 15150
rect 8010 15130 8030 15150
rect 8030 15130 8035 15150
rect 8005 15125 8035 15130
rect 8085 15150 8115 15155
rect 8085 15130 8090 15150
rect 8090 15130 8110 15150
rect 8110 15130 8115 15150
rect 8085 15125 8115 15130
rect 8165 15150 8195 15155
rect 8165 15130 8170 15150
rect 8170 15130 8190 15150
rect 8190 15130 8195 15150
rect 8165 15125 8195 15130
rect 8245 15150 8275 15155
rect 8245 15130 8250 15150
rect 8250 15130 8270 15150
rect 8270 15130 8275 15150
rect 8245 15125 8275 15130
rect 8325 15150 8355 15155
rect 8325 15130 8330 15150
rect 8330 15130 8350 15150
rect 8350 15130 8355 15150
rect 8325 15125 8355 15130
rect 8405 15150 8435 15155
rect 8405 15130 8410 15150
rect 8410 15130 8430 15150
rect 8430 15130 8435 15150
rect 8405 15125 8435 15130
rect 8485 15150 8515 15155
rect 8485 15130 8490 15150
rect 8490 15130 8510 15150
rect 8510 15130 8515 15150
rect 8485 15125 8515 15130
rect 8565 15150 8595 15155
rect 8565 15130 8570 15150
rect 8570 15130 8590 15150
rect 8590 15130 8595 15150
rect 8565 15125 8595 15130
rect 8645 15150 8675 15155
rect 8645 15130 8650 15150
rect 8650 15130 8670 15150
rect 8670 15130 8675 15150
rect 8645 15125 8675 15130
rect 8725 15150 8755 15155
rect 8725 15130 8730 15150
rect 8730 15130 8750 15150
rect 8750 15130 8755 15150
rect 8725 15125 8755 15130
rect 8805 15150 8835 15155
rect 8805 15130 8810 15150
rect 8810 15130 8830 15150
rect 8830 15130 8835 15150
rect 8805 15125 8835 15130
rect 8885 15150 8915 15155
rect 8885 15130 8890 15150
rect 8890 15130 8910 15150
rect 8910 15130 8915 15150
rect 8885 15125 8915 15130
rect 8965 15150 8995 15155
rect 8965 15130 8970 15150
rect 8970 15130 8990 15150
rect 8990 15130 8995 15150
rect 8965 15125 8995 15130
rect 9045 15150 9075 15155
rect 9045 15130 9050 15150
rect 9050 15130 9070 15150
rect 9070 15130 9075 15150
rect 9045 15125 9075 15130
rect 9125 15150 9155 15155
rect 9125 15130 9130 15150
rect 9130 15130 9150 15150
rect 9150 15130 9155 15150
rect 9125 15125 9155 15130
rect 9205 15150 9235 15155
rect 9205 15130 9210 15150
rect 9210 15130 9230 15150
rect 9230 15130 9235 15150
rect 9205 15125 9235 15130
rect 9285 15150 9315 15155
rect 9285 15130 9290 15150
rect 9290 15130 9310 15150
rect 9310 15130 9315 15150
rect 9285 15125 9315 15130
rect 9365 15150 9395 15155
rect 9365 15130 9370 15150
rect 9370 15130 9390 15150
rect 9390 15130 9395 15150
rect 9365 15125 9395 15130
rect 9445 15150 9475 15155
rect 9445 15130 9450 15150
rect 9450 15130 9470 15150
rect 9470 15130 9475 15150
rect 9445 15125 9475 15130
rect 11565 15150 11595 15155
rect 11565 15130 11570 15150
rect 11570 15130 11590 15150
rect 11590 15130 11595 15150
rect 11565 15125 11595 15130
rect 11645 15150 11675 15155
rect 11645 15130 11650 15150
rect 11650 15130 11670 15150
rect 11670 15130 11675 15150
rect 11645 15125 11675 15130
rect 11725 15150 11755 15155
rect 11725 15130 11730 15150
rect 11730 15130 11750 15150
rect 11750 15130 11755 15150
rect 11725 15125 11755 15130
rect 11805 15150 11835 15155
rect 11805 15130 11810 15150
rect 11810 15130 11830 15150
rect 11830 15130 11835 15150
rect 11805 15125 11835 15130
rect 11885 15150 11915 15155
rect 11885 15130 11890 15150
rect 11890 15130 11910 15150
rect 11910 15130 11915 15150
rect 11885 15125 11915 15130
rect 11965 15150 11995 15155
rect 11965 15130 11970 15150
rect 11970 15130 11990 15150
rect 11990 15130 11995 15150
rect 11965 15125 11995 15130
rect 12045 15150 12075 15155
rect 12045 15130 12050 15150
rect 12050 15130 12070 15150
rect 12070 15130 12075 15150
rect 12045 15125 12075 15130
rect 12125 15150 12155 15155
rect 12125 15130 12130 15150
rect 12130 15130 12150 15150
rect 12150 15130 12155 15150
rect 12125 15125 12155 15130
rect 12205 15150 12235 15155
rect 12205 15130 12210 15150
rect 12210 15130 12230 15150
rect 12230 15130 12235 15150
rect 12205 15125 12235 15130
rect 12285 15150 12315 15155
rect 12285 15130 12290 15150
rect 12290 15130 12310 15150
rect 12310 15130 12315 15150
rect 12285 15125 12315 15130
rect 12365 15150 12395 15155
rect 12365 15130 12370 15150
rect 12370 15130 12390 15150
rect 12390 15130 12395 15150
rect 12365 15125 12395 15130
rect 12445 15150 12475 15155
rect 12445 15130 12450 15150
rect 12450 15130 12470 15150
rect 12470 15130 12475 15150
rect 12445 15125 12475 15130
rect 12525 15150 12555 15155
rect 12525 15130 12530 15150
rect 12530 15130 12550 15150
rect 12550 15130 12555 15150
rect 12525 15125 12555 15130
rect 12605 15150 12635 15155
rect 12605 15130 12610 15150
rect 12610 15130 12630 15150
rect 12630 15130 12635 15150
rect 12605 15125 12635 15130
rect 12685 15150 12715 15155
rect 12685 15130 12690 15150
rect 12690 15130 12710 15150
rect 12710 15130 12715 15150
rect 12685 15125 12715 15130
rect 12765 15150 12795 15155
rect 12765 15130 12770 15150
rect 12770 15130 12790 15150
rect 12790 15130 12795 15150
rect 12765 15125 12795 15130
rect 12845 15150 12875 15155
rect 12845 15130 12850 15150
rect 12850 15130 12870 15150
rect 12870 15130 12875 15150
rect 12845 15125 12875 15130
rect 12925 15150 12955 15155
rect 12925 15130 12930 15150
rect 12930 15130 12950 15150
rect 12950 15130 12955 15150
rect 12925 15125 12955 15130
rect 13005 15150 13035 15155
rect 13005 15130 13010 15150
rect 13010 15130 13030 15150
rect 13030 15130 13035 15150
rect 13005 15125 13035 15130
rect 13085 15150 13115 15155
rect 13085 15130 13090 15150
rect 13090 15130 13110 15150
rect 13110 15130 13115 15150
rect 13085 15125 13115 15130
rect 13165 15150 13195 15155
rect 13165 15130 13170 15150
rect 13170 15130 13190 15150
rect 13190 15130 13195 15150
rect 13165 15125 13195 15130
rect 13245 15150 13275 15155
rect 13245 15130 13250 15150
rect 13250 15130 13270 15150
rect 13270 15130 13275 15150
rect 13245 15125 13275 15130
rect 13325 15150 13355 15155
rect 13325 15130 13330 15150
rect 13330 15130 13350 15150
rect 13350 15130 13355 15150
rect 13325 15125 13355 15130
rect 13405 15150 13435 15155
rect 13405 15130 13410 15150
rect 13410 15130 13430 15150
rect 13430 15130 13435 15150
rect 13405 15125 13435 15130
rect 13485 15150 13515 15155
rect 13485 15130 13490 15150
rect 13490 15130 13510 15150
rect 13510 15130 13515 15150
rect 13485 15125 13515 15130
rect 13565 15150 13595 15155
rect 13565 15130 13570 15150
rect 13570 15130 13590 15150
rect 13590 15130 13595 15150
rect 13565 15125 13595 15130
rect 13645 15150 13675 15155
rect 13645 15130 13650 15150
rect 13650 15130 13670 15150
rect 13670 15130 13675 15150
rect 13645 15125 13675 15130
rect 13725 15150 13755 15155
rect 13725 15130 13730 15150
rect 13730 15130 13750 15150
rect 13750 15130 13755 15150
rect 13725 15125 13755 15130
rect 13805 15150 13835 15155
rect 13805 15130 13810 15150
rect 13810 15130 13830 15150
rect 13830 15130 13835 15150
rect 13805 15125 13835 15130
rect 13885 15150 13915 15155
rect 13885 15130 13890 15150
rect 13890 15130 13910 15150
rect 13910 15130 13915 15150
rect 13885 15125 13915 15130
rect 13965 15150 13995 15155
rect 13965 15130 13970 15150
rect 13970 15130 13990 15150
rect 13990 15130 13995 15150
rect 13965 15125 13995 15130
rect 14045 15150 14075 15155
rect 14045 15130 14050 15150
rect 14050 15130 14070 15150
rect 14070 15130 14075 15150
rect 14045 15125 14075 15130
rect 14125 15150 14155 15155
rect 14125 15130 14130 15150
rect 14130 15130 14150 15150
rect 14150 15130 14155 15150
rect 14125 15125 14155 15130
rect 14205 15150 14235 15155
rect 14205 15130 14210 15150
rect 14210 15130 14230 15150
rect 14230 15130 14235 15150
rect 14205 15125 14235 15130
rect 14285 15150 14315 15155
rect 14285 15130 14290 15150
rect 14290 15130 14310 15150
rect 14310 15130 14315 15150
rect 14285 15125 14315 15130
rect 14365 15150 14395 15155
rect 14365 15130 14370 15150
rect 14370 15130 14390 15150
rect 14390 15130 14395 15150
rect 14365 15125 14395 15130
rect 14445 15150 14475 15155
rect 14445 15130 14450 15150
rect 14450 15130 14470 15150
rect 14470 15130 14475 15150
rect 14445 15125 14475 15130
rect 14525 15150 14555 15155
rect 14525 15130 14530 15150
rect 14530 15130 14550 15150
rect 14550 15130 14555 15150
rect 14525 15125 14555 15130
rect 14605 15150 14635 15155
rect 14605 15130 14610 15150
rect 14610 15130 14630 15150
rect 14630 15130 14635 15150
rect 14605 15125 14635 15130
rect 14685 15150 14715 15155
rect 14685 15130 14690 15150
rect 14690 15130 14710 15150
rect 14710 15130 14715 15150
rect 14685 15125 14715 15130
rect 16765 15150 16795 15155
rect 16765 15130 16770 15150
rect 16770 15130 16790 15150
rect 16790 15130 16795 15150
rect 16765 15125 16795 15130
rect 16845 15150 16875 15155
rect 16845 15130 16850 15150
rect 16850 15130 16870 15150
rect 16870 15130 16875 15150
rect 16845 15125 16875 15130
rect 16925 15150 16955 15155
rect 16925 15130 16930 15150
rect 16930 15130 16950 15150
rect 16950 15130 16955 15150
rect 16925 15125 16955 15130
rect 17005 15150 17035 15155
rect 17005 15130 17010 15150
rect 17010 15130 17030 15150
rect 17030 15130 17035 15150
rect 17005 15125 17035 15130
rect 17085 15150 17115 15155
rect 17085 15130 17090 15150
rect 17090 15130 17110 15150
rect 17110 15130 17115 15150
rect 17085 15125 17115 15130
rect 17165 15150 17195 15155
rect 17165 15130 17170 15150
rect 17170 15130 17190 15150
rect 17190 15130 17195 15150
rect 17165 15125 17195 15130
rect 17245 15150 17275 15155
rect 17245 15130 17250 15150
rect 17250 15130 17270 15150
rect 17270 15130 17275 15150
rect 17245 15125 17275 15130
rect 17325 15150 17355 15155
rect 17325 15130 17330 15150
rect 17330 15130 17350 15150
rect 17350 15130 17355 15150
rect 17325 15125 17355 15130
rect 17405 15150 17435 15155
rect 17405 15130 17410 15150
rect 17410 15130 17430 15150
rect 17430 15130 17435 15150
rect 17405 15125 17435 15130
rect 17485 15150 17515 15155
rect 17485 15130 17490 15150
rect 17490 15130 17510 15150
rect 17510 15130 17515 15150
rect 17485 15125 17515 15130
rect 17565 15150 17595 15155
rect 17565 15130 17570 15150
rect 17570 15130 17590 15150
rect 17590 15130 17595 15150
rect 17565 15125 17595 15130
rect 17645 15150 17675 15155
rect 17645 15130 17650 15150
rect 17650 15130 17670 15150
rect 17670 15130 17675 15150
rect 17645 15125 17675 15130
rect 17725 15150 17755 15155
rect 17725 15130 17730 15150
rect 17730 15130 17750 15150
rect 17750 15130 17755 15150
rect 17725 15125 17755 15130
rect 17805 15150 17835 15155
rect 17805 15130 17810 15150
rect 17810 15130 17830 15150
rect 17830 15130 17835 15150
rect 17805 15125 17835 15130
rect 17885 15150 17915 15155
rect 17885 15130 17890 15150
rect 17890 15130 17910 15150
rect 17910 15130 17915 15150
rect 17885 15125 17915 15130
rect 17965 15150 17995 15155
rect 17965 15130 17970 15150
rect 17970 15130 17990 15150
rect 17990 15130 17995 15150
rect 17965 15125 17995 15130
rect 18045 15150 18075 15155
rect 18045 15130 18050 15150
rect 18050 15130 18070 15150
rect 18070 15130 18075 15150
rect 18045 15125 18075 15130
rect 18125 15150 18155 15155
rect 18125 15130 18130 15150
rect 18130 15130 18150 15150
rect 18150 15130 18155 15150
rect 18125 15125 18155 15130
rect 18205 15150 18235 15155
rect 18205 15130 18210 15150
rect 18210 15130 18230 15150
rect 18230 15130 18235 15150
rect 18205 15125 18235 15130
rect 18285 15150 18315 15155
rect 18285 15130 18290 15150
rect 18290 15130 18310 15150
rect 18310 15130 18315 15150
rect 18285 15125 18315 15130
rect 18365 15150 18395 15155
rect 18365 15130 18370 15150
rect 18370 15130 18390 15150
rect 18390 15130 18395 15150
rect 18365 15125 18395 15130
rect 18445 15150 18475 15155
rect 18445 15130 18450 15150
rect 18450 15130 18470 15150
rect 18470 15130 18475 15150
rect 18445 15125 18475 15130
rect 18525 15150 18555 15155
rect 18525 15130 18530 15150
rect 18530 15130 18550 15150
rect 18550 15130 18555 15150
rect 18525 15125 18555 15130
rect 18605 15150 18635 15155
rect 18605 15130 18610 15150
rect 18610 15130 18630 15150
rect 18630 15130 18635 15150
rect 18605 15125 18635 15130
rect 18685 15150 18715 15155
rect 18685 15130 18690 15150
rect 18690 15130 18710 15150
rect 18710 15130 18715 15150
rect 18685 15125 18715 15130
rect 18765 15150 18795 15155
rect 18765 15130 18770 15150
rect 18770 15130 18790 15150
rect 18790 15130 18795 15150
rect 18765 15125 18795 15130
rect 18845 15150 18875 15155
rect 18845 15130 18850 15150
rect 18850 15130 18870 15150
rect 18870 15130 18875 15150
rect 18845 15125 18875 15130
rect 18925 15150 18955 15155
rect 18925 15130 18930 15150
rect 18930 15130 18950 15150
rect 18950 15130 18955 15150
rect 18925 15125 18955 15130
rect 19005 15150 19035 15155
rect 19005 15130 19010 15150
rect 19010 15130 19030 15150
rect 19030 15130 19035 15150
rect 19005 15125 19035 15130
rect 19085 15150 19115 15155
rect 19085 15130 19090 15150
rect 19090 15130 19110 15150
rect 19110 15130 19115 15150
rect 19085 15125 19115 15130
rect 19165 15150 19195 15155
rect 19165 15130 19170 15150
rect 19170 15130 19190 15150
rect 19190 15130 19195 15150
rect 19165 15125 19195 15130
rect 19245 15150 19275 15155
rect 19245 15130 19250 15150
rect 19250 15130 19270 15150
rect 19270 15130 19275 15150
rect 19245 15125 19275 15130
rect 19325 15150 19355 15155
rect 19325 15130 19330 15150
rect 19330 15130 19350 15150
rect 19350 15130 19355 15150
rect 19325 15125 19355 15130
rect 19405 15150 19435 15155
rect 19405 15130 19410 15150
rect 19410 15130 19430 15150
rect 19430 15130 19435 15150
rect 19405 15125 19435 15130
rect 19485 15150 19515 15155
rect 19485 15130 19490 15150
rect 19490 15130 19510 15150
rect 19510 15130 19515 15150
rect 19485 15125 19515 15130
rect 19565 15150 19595 15155
rect 19565 15130 19570 15150
rect 19570 15130 19590 15150
rect 19590 15130 19595 15150
rect 19565 15125 19595 15130
rect 19645 15150 19675 15155
rect 19645 15130 19650 15150
rect 19650 15130 19670 15150
rect 19670 15130 19675 15150
rect 19645 15125 19675 15130
rect 19725 15150 19755 15155
rect 19725 15130 19730 15150
rect 19730 15130 19750 15150
rect 19750 15130 19755 15150
rect 19725 15125 19755 15130
rect 19805 15150 19835 15155
rect 19805 15130 19810 15150
rect 19810 15130 19830 15150
rect 19830 15130 19835 15150
rect 19805 15125 19835 15130
rect 19885 15150 19915 15155
rect 19885 15130 19890 15150
rect 19890 15130 19910 15150
rect 19910 15130 19915 15150
rect 19885 15125 19915 15130
rect 19965 15150 19995 15155
rect 19965 15130 19970 15150
rect 19970 15130 19990 15150
rect 19990 15130 19995 15150
rect 19965 15125 19995 15130
rect 20045 15150 20075 15155
rect 20045 15130 20050 15150
rect 20050 15130 20070 15150
rect 20070 15130 20075 15150
rect 20045 15125 20075 15130
rect 20125 15150 20155 15155
rect 20125 15130 20130 15150
rect 20130 15130 20150 15150
rect 20150 15130 20155 15150
rect 20125 15125 20155 15130
rect 20205 15150 20235 15155
rect 20205 15130 20210 15150
rect 20210 15130 20230 15150
rect 20230 15130 20235 15150
rect 20205 15125 20235 15130
rect 20285 15150 20315 15155
rect 20285 15130 20290 15150
rect 20290 15130 20310 15150
rect 20310 15130 20315 15150
rect 20285 15125 20315 15130
rect 20365 15150 20395 15155
rect 20365 15130 20370 15150
rect 20370 15130 20390 15150
rect 20390 15130 20395 15150
rect 20365 15125 20395 15130
rect 20445 15150 20475 15155
rect 20445 15130 20450 15150
rect 20450 15130 20470 15150
rect 20470 15130 20475 15150
rect 20445 15125 20475 15130
rect 20525 15150 20555 15155
rect 20525 15130 20530 15150
rect 20530 15130 20550 15150
rect 20550 15130 20555 15150
rect 20525 15125 20555 15130
rect 20605 15150 20635 15155
rect 20605 15130 20610 15150
rect 20610 15130 20630 15150
rect 20630 15130 20635 15150
rect 20605 15125 20635 15130
rect 20685 15150 20715 15155
rect 20685 15130 20690 15150
rect 20690 15130 20710 15150
rect 20710 15130 20715 15150
rect 20685 15125 20715 15130
rect 20765 15150 20795 15155
rect 20765 15130 20770 15150
rect 20770 15130 20790 15150
rect 20790 15130 20795 15150
rect 20765 15125 20795 15130
rect 20845 15150 20875 15155
rect 20845 15130 20850 15150
rect 20850 15130 20870 15150
rect 20870 15130 20875 15150
rect 20845 15125 20875 15130
rect 20925 15150 20955 15155
rect 20925 15130 20930 15150
rect 20930 15130 20950 15150
rect 20950 15130 20955 15150
rect 20925 15125 20955 15130
rect 5 14990 35 14995
rect 5 14970 10 14990
rect 10 14970 30 14990
rect 30 14970 35 14990
rect 5 14965 35 14970
rect 85 14990 115 14995
rect 85 14970 90 14990
rect 90 14970 110 14990
rect 110 14970 115 14990
rect 85 14965 115 14970
rect 165 14990 195 14995
rect 165 14970 170 14990
rect 170 14970 190 14990
rect 190 14970 195 14990
rect 165 14965 195 14970
rect 245 14990 275 14995
rect 245 14970 250 14990
rect 250 14970 270 14990
rect 270 14970 275 14990
rect 245 14965 275 14970
rect 325 14990 355 14995
rect 325 14970 330 14990
rect 330 14970 350 14990
rect 350 14970 355 14990
rect 325 14965 355 14970
rect 405 14990 435 14995
rect 405 14970 410 14990
rect 410 14970 430 14990
rect 430 14970 435 14990
rect 405 14965 435 14970
rect 485 14990 515 14995
rect 485 14970 490 14990
rect 490 14970 510 14990
rect 510 14970 515 14990
rect 485 14965 515 14970
rect 565 14990 595 14995
rect 565 14970 570 14990
rect 570 14970 590 14990
rect 590 14970 595 14990
rect 565 14965 595 14970
rect 645 14990 675 14995
rect 645 14970 650 14990
rect 650 14970 670 14990
rect 670 14970 675 14990
rect 645 14965 675 14970
rect 725 14990 755 14995
rect 725 14970 730 14990
rect 730 14970 750 14990
rect 750 14970 755 14990
rect 725 14965 755 14970
rect 805 14990 835 14995
rect 805 14970 810 14990
rect 810 14970 830 14990
rect 830 14970 835 14990
rect 805 14965 835 14970
rect 885 14990 915 14995
rect 885 14970 890 14990
rect 890 14970 910 14990
rect 910 14970 915 14990
rect 885 14965 915 14970
rect 965 14990 995 14995
rect 965 14970 970 14990
rect 970 14970 990 14990
rect 990 14970 995 14990
rect 965 14965 995 14970
rect 1045 14990 1075 14995
rect 1045 14970 1050 14990
rect 1050 14970 1070 14990
rect 1070 14970 1075 14990
rect 1045 14965 1075 14970
rect 1125 14990 1155 14995
rect 1125 14970 1130 14990
rect 1130 14970 1150 14990
rect 1150 14970 1155 14990
rect 1125 14965 1155 14970
rect 1205 14990 1235 14995
rect 1205 14970 1210 14990
rect 1210 14970 1230 14990
rect 1230 14970 1235 14990
rect 1205 14965 1235 14970
rect 1285 14990 1315 14995
rect 1285 14970 1290 14990
rect 1290 14970 1310 14990
rect 1310 14970 1315 14990
rect 1285 14965 1315 14970
rect 1365 14990 1395 14995
rect 1365 14970 1370 14990
rect 1370 14970 1390 14990
rect 1390 14970 1395 14990
rect 1365 14965 1395 14970
rect 1445 14990 1475 14995
rect 1445 14970 1450 14990
rect 1450 14970 1470 14990
rect 1470 14970 1475 14990
rect 1445 14965 1475 14970
rect 1525 14990 1555 14995
rect 1525 14970 1530 14990
rect 1530 14970 1550 14990
rect 1550 14970 1555 14990
rect 1525 14965 1555 14970
rect 1605 14990 1635 14995
rect 1605 14970 1610 14990
rect 1610 14970 1630 14990
rect 1630 14970 1635 14990
rect 1605 14965 1635 14970
rect 1685 14990 1715 14995
rect 1685 14970 1690 14990
rect 1690 14970 1710 14990
rect 1710 14970 1715 14990
rect 1685 14965 1715 14970
rect 1765 14990 1795 14995
rect 1765 14970 1770 14990
rect 1770 14970 1790 14990
rect 1790 14970 1795 14990
rect 1765 14965 1795 14970
rect 1845 14990 1875 14995
rect 1845 14970 1850 14990
rect 1850 14970 1870 14990
rect 1870 14970 1875 14990
rect 1845 14965 1875 14970
rect 1925 14990 1955 14995
rect 1925 14970 1930 14990
rect 1930 14970 1950 14990
rect 1950 14970 1955 14990
rect 1925 14965 1955 14970
rect 2005 14990 2035 14995
rect 2005 14970 2010 14990
rect 2010 14970 2030 14990
rect 2030 14970 2035 14990
rect 2005 14965 2035 14970
rect 2085 14990 2115 14995
rect 2085 14970 2090 14990
rect 2090 14970 2110 14990
rect 2110 14970 2115 14990
rect 2085 14965 2115 14970
rect 2165 14990 2195 14995
rect 2165 14970 2170 14990
rect 2170 14970 2190 14990
rect 2190 14970 2195 14990
rect 2165 14965 2195 14970
rect 2245 14990 2275 14995
rect 2245 14970 2250 14990
rect 2250 14970 2270 14990
rect 2270 14970 2275 14990
rect 2245 14965 2275 14970
rect 2325 14990 2355 14995
rect 2325 14970 2330 14990
rect 2330 14970 2350 14990
rect 2350 14970 2355 14990
rect 2325 14965 2355 14970
rect 2405 14990 2435 14995
rect 2405 14970 2410 14990
rect 2410 14970 2430 14990
rect 2430 14970 2435 14990
rect 2405 14965 2435 14970
rect 2485 14990 2515 14995
rect 2485 14970 2490 14990
rect 2490 14970 2510 14990
rect 2510 14970 2515 14990
rect 2485 14965 2515 14970
rect 2565 14990 2595 14995
rect 2565 14970 2570 14990
rect 2570 14970 2590 14990
rect 2590 14970 2595 14990
rect 2565 14965 2595 14970
rect 2645 14990 2675 14995
rect 2645 14970 2650 14990
rect 2650 14970 2670 14990
rect 2670 14970 2675 14990
rect 2645 14965 2675 14970
rect 2725 14990 2755 14995
rect 2725 14970 2730 14990
rect 2730 14970 2750 14990
rect 2750 14970 2755 14990
rect 2725 14965 2755 14970
rect 2805 14990 2835 14995
rect 2805 14970 2810 14990
rect 2810 14970 2830 14990
rect 2830 14970 2835 14990
rect 2805 14965 2835 14970
rect 2885 14990 2915 14995
rect 2885 14970 2890 14990
rect 2890 14970 2910 14990
rect 2910 14970 2915 14990
rect 2885 14965 2915 14970
rect 2965 14990 2995 14995
rect 2965 14970 2970 14990
rect 2970 14970 2990 14990
rect 2990 14970 2995 14990
rect 2965 14965 2995 14970
rect 3045 14990 3075 14995
rect 3045 14970 3050 14990
rect 3050 14970 3070 14990
rect 3070 14970 3075 14990
rect 3045 14965 3075 14970
rect 3125 14990 3155 14995
rect 3125 14970 3130 14990
rect 3130 14970 3150 14990
rect 3150 14970 3155 14990
rect 3125 14965 3155 14970
rect 3205 14990 3235 14995
rect 3205 14970 3210 14990
rect 3210 14970 3230 14990
rect 3230 14970 3235 14990
rect 3205 14965 3235 14970
rect 3285 14990 3315 14995
rect 3285 14970 3290 14990
rect 3290 14970 3310 14990
rect 3310 14970 3315 14990
rect 3285 14965 3315 14970
rect 3365 14990 3395 14995
rect 3365 14970 3370 14990
rect 3370 14970 3390 14990
rect 3390 14970 3395 14990
rect 3365 14965 3395 14970
rect 3445 14990 3475 14995
rect 3445 14970 3450 14990
rect 3450 14970 3470 14990
rect 3470 14970 3475 14990
rect 3445 14965 3475 14970
rect 3525 14990 3555 14995
rect 3525 14970 3530 14990
rect 3530 14970 3550 14990
rect 3550 14970 3555 14990
rect 3525 14965 3555 14970
rect 3605 14990 3635 14995
rect 3605 14970 3610 14990
rect 3610 14970 3630 14990
rect 3630 14970 3635 14990
rect 3605 14965 3635 14970
rect 3685 14990 3715 14995
rect 3685 14970 3690 14990
rect 3690 14970 3710 14990
rect 3710 14970 3715 14990
rect 3685 14965 3715 14970
rect 3765 14990 3795 14995
rect 3765 14970 3770 14990
rect 3770 14970 3790 14990
rect 3790 14970 3795 14990
rect 3765 14965 3795 14970
rect 3845 14990 3875 14995
rect 3845 14970 3850 14990
rect 3850 14970 3870 14990
rect 3870 14970 3875 14990
rect 3845 14965 3875 14970
rect 3925 14990 3955 14995
rect 3925 14970 3930 14990
rect 3930 14970 3950 14990
rect 3950 14970 3955 14990
rect 3925 14965 3955 14970
rect 4005 14990 4035 14995
rect 4005 14970 4010 14990
rect 4010 14970 4030 14990
rect 4030 14970 4035 14990
rect 4005 14965 4035 14970
rect 4085 14990 4115 14995
rect 4085 14970 4090 14990
rect 4090 14970 4110 14990
rect 4110 14970 4115 14990
rect 4085 14965 4115 14970
rect 4165 14990 4195 14995
rect 4165 14970 4170 14990
rect 4170 14970 4190 14990
rect 4190 14970 4195 14990
rect 4165 14965 4195 14970
rect 6245 14990 6275 14995
rect 6245 14970 6250 14990
rect 6250 14970 6270 14990
rect 6270 14970 6275 14990
rect 6245 14965 6275 14970
rect 6325 14990 6355 14995
rect 6325 14970 6330 14990
rect 6330 14970 6350 14990
rect 6350 14970 6355 14990
rect 6325 14965 6355 14970
rect 6405 14990 6435 14995
rect 6405 14970 6410 14990
rect 6410 14970 6430 14990
rect 6430 14970 6435 14990
rect 6405 14965 6435 14970
rect 6485 14990 6515 14995
rect 6485 14970 6490 14990
rect 6490 14970 6510 14990
rect 6510 14970 6515 14990
rect 6485 14965 6515 14970
rect 6565 14990 6595 14995
rect 6565 14970 6570 14990
rect 6570 14970 6590 14990
rect 6590 14970 6595 14990
rect 6565 14965 6595 14970
rect 6645 14990 6675 14995
rect 6645 14970 6650 14990
rect 6650 14970 6670 14990
rect 6670 14970 6675 14990
rect 6645 14965 6675 14970
rect 6725 14990 6755 14995
rect 6725 14970 6730 14990
rect 6730 14970 6750 14990
rect 6750 14970 6755 14990
rect 6725 14965 6755 14970
rect 6805 14990 6835 14995
rect 6805 14970 6810 14990
rect 6810 14970 6830 14990
rect 6830 14970 6835 14990
rect 6805 14965 6835 14970
rect 6885 14990 6915 14995
rect 6885 14970 6890 14990
rect 6890 14970 6910 14990
rect 6910 14970 6915 14990
rect 6885 14965 6915 14970
rect 6965 14990 6995 14995
rect 6965 14970 6970 14990
rect 6970 14970 6990 14990
rect 6990 14970 6995 14990
rect 6965 14965 6995 14970
rect 7045 14990 7075 14995
rect 7045 14970 7050 14990
rect 7050 14970 7070 14990
rect 7070 14970 7075 14990
rect 7045 14965 7075 14970
rect 7125 14990 7155 14995
rect 7125 14970 7130 14990
rect 7130 14970 7150 14990
rect 7150 14970 7155 14990
rect 7125 14965 7155 14970
rect 7205 14990 7235 14995
rect 7205 14970 7210 14990
rect 7210 14970 7230 14990
rect 7230 14970 7235 14990
rect 7205 14965 7235 14970
rect 7285 14990 7315 14995
rect 7285 14970 7290 14990
rect 7290 14970 7310 14990
rect 7310 14970 7315 14990
rect 7285 14965 7315 14970
rect 7365 14990 7395 14995
rect 7365 14970 7370 14990
rect 7370 14970 7390 14990
rect 7390 14970 7395 14990
rect 7365 14965 7395 14970
rect 7445 14990 7475 14995
rect 7445 14970 7450 14990
rect 7450 14970 7470 14990
rect 7470 14970 7475 14990
rect 7445 14965 7475 14970
rect 7525 14990 7555 14995
rect 7525 14970 7530 14990
rect 7530 14970 7550 14990
rect 7550 14970 7555 14990
rect 7525 14965 7555 14970
rect 7605 14990 7635 14995
rect 7605 14970 7610 14990
rect 7610 14970 7630 14990
rect 7630 14970 7635 14990
rect 7605 14965 7635 14970
rect 7685 14990 7715 14995
rect 7685 14970 7690 14990
rect 7690 14970 7710 14990
rect 7710 14970 7715 14990
rect 7685 14965 7715 14970
rect 7765 14990 7795 14995
rect 7765 14970 7770 14990
rect 7770 14970 7790 14990
rect 7790 14970 7795 14990
rect 7765 14965 7795 14970
rect 7845 14990 7875 14995
rect 7845 14970 7850 14990
rect 7850 14970 7870 14990
rect 7870 14970 7875 14990
rect 7845 14965 7875 14970
rect 7925 14990 7955 14995
rect 7925 14970 7930 14990
rect 7930 14970 7950 14990
rect 7950 14970 7955 14990
rect 7925 14965 7955 14970
rect 8005 14990 8035 14995
rect 8005 14970 8010 14990
rect 8010 14970 8030 14990
rect 8030 14970 8035 14990
rect 8005 14965 8035 14970
rect 8085 14990 8115 14995
rect 8085 14970 8090 14990
rect 8090 14970 8110 14990
rect 8110 14970 8115 14990
rect 8085 14965 8115 14970
rect 8165 14990 8195 14995
rect 8165 14970 8170 14990
rect 8170 14970 8190 14990
rect 8190 14970 8195 14990
rect 8165 14965 8195 14970
rect 8245 14990 8275 14995
rect 8245 14970 8250 14990
rect 8250 14970 8270 14990
rect 8270 14970 8275 14990
rect 8245 14965 8275 14970
rect 8325 14990 8355 14995
rect 8325 14970 8330 14990
rect 8330 14970 8350 14990
rect 8350 14970 8355 14990
rect 8325 14965 8355 14970
rect 8405 14990 8435 14995
rect 8405 14970 8410 14990
rect 8410 14970 8430 14990
rect 8430 14970 8435 14990
rect 8405 14965 8435 14970
rect 8485 14990 8515 14995
rect 8485 14970 8490 14990
rect 8490 14970 8510 14990
rect 8510 14970 8515 14990
rect 8485 14965 8515 14970
rect 8565 14990 8595 14995
rect 8565 14970 8570 14990
rect 8570 14970 8590 14990
rect 8590 14970 8595 14990
rect 8565 14965 8595 14970
rect 8645 14990 8675 14995
rect 8645 14970 8650 14990
rect 8650 14970 8670 14990
rect 8670 14970 8675 14990
rect 8645 14965 8675 14970
rect 8725 14990 8755 14995
rect 8725 14970 8730 14990
rect 8730 14970 8750 14990
rect 8750 14970 8755 14990
rect 8725 14965 8755 14970
rect 8805 14990 8835 14995
rect 8805 14970 8810 14990
rect 8810 14970 8830 14990
rect 8830 14970 8835 14990
rect 8805 14965 8835 14970
rect 8885 14990 8915 14995
rect 8885 14970 8890 14990
rect 8890 14970 8910 14990
rect 8910 14970 8915 14990
rect 8885 14965 8915 14970
rect 8965 14990 8995 14995
rect 8965 14970 8970 14990
rect 8970 14970 8990 14990
rect 8990 14970 8995 14990
rect 8965 14965 8995 14970
rect 9045 14990 9075 14995
rect 9045 14970 9050 14990
rect 9050 14970 9070 14990
rect 9070 14970 9075 14990
rect 9045 14965 9075 14970
rect 9125 14990 9155 14995
rect 9125 14970 9130 14990
rect 9130 14970 9150 14990
rect 9150 14970 9155 14990
rect 9125 14965 9155 14970
rect 9205 14990 9235 14995
rect 9205 14970 9210 14990
rect 9210 14970 9230 14990
rect 9230 14970 9235 14990
rect 9205 14965 9235 14970
rect 9285 14990 9315 14995
rect 9285 14970 9290 14990
rect 9290 14970 9310 14990
rect 9310 14970 9315 14990
rect 9285 14965 9315 14970
rect 9365 14990 9395 14995
rect 9365 14970 9370 14990
rect 9370 14970 9390 14990
rect 9390 14970 9395 14990
rect 9365 14965 9395 14970
rect 9445 14990 9475 14995
rect 9445 14970 9450 14990
rect 9450 14970 9470 14990
rect 9470 14970 9475 14990
rect 9445 14965 9475 14970
rect 11565 14990 11595 14995
rect 11565 14970 11570 14990
rect 11570 14970 11590 14990
rect 11590 14970 11595 14990
rect 11565 14965 11595 14970
rect 11645 14990 11675 14995
rect 11645 14970 11650 14990
rect 11650 14970 11670 14990
rect 11670 14970 11675 14990
rect 11645 14965 11675 14970
rect 11725 14990 11755 14995
rect 11725 14970 11730 14990
rect 11730 14970 11750 14990
rect 11750 14970 11755 14990
rect 11725 14965 11755 14970
rect 11805 14990 11835 14995
rect 11805 14970 11810 14990
rect 11810 14970 11830 14990
rect 11830 14970 11835 14990
rect 11805 14965 11835 14970
rect 11885 14990 11915 14995
rect 11885 14970 11890 14990
rect 11890 14970 11910 14990
rect 11910 14970 11915 14990
rect 11885 14965 11915 14970
rect 11965 14990 11995 14995
rect 11965 14970 11970 14990
rect 11970 14970 11990 14990
rect 11990 14970 11995 14990
rect 11965 14965 11995 14970
rect 12045 14990 12075 14995
rect 12045 14970 12050 14990
rect 12050 14970 12070 14990
rect 12070 14970 12075 14990
rect 12045 14965 12075 14970
rect 12125 14990 12155 14995
rect 12125 14970 12130 14990
rect 12130 14970 12150 14990
rect 12150 14970 12155 14990
rect 12125 14965 12155 14970
rect 12205 14990 12235 14995
rect 12205 14970 12210 14990
rect 12210 14970 12230 14990
rect 12230 14970 12235 14990
rect 12205 14965 12235 14970
rect 12285 14990 12315 14995
rect 12285 14970 12290 14990
rect 12290 14970 12310 14990
rect 12310 14970 12315 14990
rect 12285 14965 12315 14970
rect 12365 14990 12395 14995
rect 12365 14970 12370 14990
rect 12370 14970 12390 14990
rect 12390 14970 12395 14990
rect 12365 14965 12395 14970
rect 12445 14990 12475 14995
rect 12445 14970 12450 14990
rect 12450 14970 12470 14990
rect 12470 14970 12475 14990
rect 12445 14965 12475 14970
rect 12525 14990 12555 14995
rect 12525 14970 12530 14990
rect 12530 14970 12550 14990
rect 12550 14970 12555 14990
rect 12525 14965 12555 14970
rect 12605 14990 12635 14995
rect 12605 14970 12610 14990
rect 12610 14970 12630 14990
rect 12630 14970 12635 14990
rect 12605 14965 12635 14970
rect 12685 14990 12715 14995
rect 12685 14970 12690 14990
rect 12690 14970 12710 14990
rect 12710 14970 12715 14990
rect 12685 14965 12715 14970
rect 12765 14990 12795 14995
rect 12765 14970 12770 14990
rect 12770 14970 12790 14990
rect 12790 14970 12795 14990
rect 12765 14965 12795 14970
rect 12845 14990 12875 14995
rect 12845 14970 12850 14990
rect 12850 14970 12870 14990
rect 12870 14970 12875 14990
rect 12845 14965 12875 14970
rect 12925 14990 12955 14995
rect 12925 14970 12930 14990
rect 12930 14970 12950 14990
rect 12950 14970 12955 14990
rect 12925 14965 12955 14970
rect 13005 14990 13035 14995
rect 13005 14970 13010 14990
rect 13010 14970 13030 14990
rect 13030 14970 13035 14990
rect 13005 14965 13035 14970
rect 13085 14990 13115 14995
rect 13085 14970 13090 14990
rect 13090 14970 13110 14990
rect 13110 14970 13115 14990
rect 13085 14965 13115 14970
rect 13165 14990 13195 14995
rect 13165 14970 13170 14990
rect 13170 14970 13190 14990
rect 13190 14970 13195 14990
rect 13165 14965 13195 14970
rect 13245 14990 13275 14995
rect 13245 14970 13250 14990
rect 13250 14970 13270 14990
rect 13270 14970 13275 14990
rect 13245 14965 13275 14970
rect 13325 14990 13355 14995
rect 13325 14970 13330 14990
rect 13330 14970 13350 14990
rect 13350 14970 13355 14990
rect 13325 14965 13355 14970
rect 13405 14990 13435 14995
rect 13405 14970 13410 14990
rect 13410 14970 13430 14990
rect 13430 14970 13435 14990
rect 13405 14965 13435 14970
rect 13485 14990 13515 14995
rect 13485 14970 13490 14990
rect 13490 14970 13510 14990
rect 13510 14970 13515 14990
rect 13485 14965 13515 14970
rect 13565 14990 13595 14995
rect 13565 14970 13570 14990
rect 13570 14970 13590 14990
rect 13590 14970 13595 14990
rect 13565 14965 13595 14970
rect 13645 14990 13675 14995
rect 13645 14970 13650 14990
rect 13650 14970 13670 14990
rect 13670 14970 13675 14990
rect 13645 14965 13675 14970
rect 13725 14990 13755 14995
rect 13725 14970 13730 14990
rect 13730 14970 13750 14990
rect 13750 14970 13755 14990
rect 13725 14965 13755 14970
rect 13805 14990 13835 14995
rect 13805 14970 13810 14990
rect 13810 14970 13830 14990
rect 13830 14970 13835 14990
rect 13805 14965 13835 14970
rect 13885 14990 13915 14995
rect 13885 14970 13890 14990
rect 13890 14970 13910 14990
rect 13910 14970 13915 14990
rect 13885 14965 13915 14970
rect 13965 14990 13995 14995
rect 13965 14970 13970 14990
rect 13970 14970 13990 14990
rect 13990 14970 13995 14990
rect 13965 14965 13995 14970
rect 14045 14990 14075 14995
rect 14045 14970 14050 14990
rect 14050 14970 14070 14990
rect 14070 14970 14075 14990
rect 14045 14965 14075 14970
rect 14125 14990 14155 14995
rect 14125 14970 14130 14990
rect 14130 14970 14150 14990
rect 14150 14970 14155 14990
rect 14125 14965 14155 14970
rect 14205 14990 14235 14995
rect 14205 14970 14210 14990
rect 14210 14970 14230 14990
rect 14230 14970 14235 14990
rect 14205 14965 14235 14970
rect 14285 14990 14315 14995
rect 14285 14970 14290 14990
rect 14290 14970 14310 14990
rect 14310 14970 14315 14990
rect 14285 14965 14315 14970
rect 14365 14990 14395 14995
rect 14365 14970 14370 14990
rect 14370 14970 14390 14990
rect 14390 14970 14395 14990
rect 14365 14965 14395 14970
rect 14445 14990 14475 14995
rect 14445 14970 14450 14990
rect 14450 14970 14470 14990
rect 14470 14970 14475 14990
rect 14445 14965 14475 14970
rect 14525 14990 14555 14995
rect 14525 14970 14530 14990
rect 14530 14970 14550 14990
rect 14550 14970 14555 14990
rect 14525 14965 14555 14970
rect 14605 14990 14635 14995
rect 14605 14970 14610 14990
rect 14610 14970 14630 14990
rect 14630 14970 14635 14990
rect 14605 14965 14635 14970
rect 14685 14990 14715 14995
rect 14685 14970 14690 14990
rect 14690 14970 14710 14990
rect 14710 14970 14715 14990
rect 14685 14965 14715 14970
rect 16765 14990 16795 14995
rect 16765 14970 16770 14990
rect 16770 14970 16790 14990
rect 16790 14970 16795 14990
rect 16765 14965 16795 14970
rect 16845 14990 16875 14995
rect 16845 14970 16850 14990
rect 16850 14970 16870 14990
rect 16870 14970 16875 14990
rect 16845 14965 16875 14970
rect 16925 14990 16955 14995
rect 16925 14970 16930 14990
rect 16930 14970 16950 14990
rect 16950 14970 16955 14990
rect 16925 14965 16955 14970
rect 17005 14990 17035 14995
rect 17005 14970 17010 14990
rect 17010 14970 17030 14990
rect 17030 14970 17035 14990
rect 17005 14965 17035 14970
rect 17085 14990 17115 14995
rect 17085 14970 17090 14990
rect 17090 14970 17110 14990
rect 17110 14970 17115 14990
rect 17085 14965 17115 14970
rect 17165 14990 17195 14995
rect 17165 14970 17170 14990
rect 17170 14970 17190 14990
rect 17190 14970 17195 14990
rect 17165 14965 17195 14970
rect 17245 14990 17275 14995
rect 17245 14970 17250 14990
rect 17250 14970 17270 14990
rect 17270 14970 17275 14990
rect 17245 14965 17275 14970
rect 17325 14990 17355 14995
rect 17325 14970 17330 14990
rect 17330 14970 17350 14990
rect 17350 14970 17355 14990
rect 17325 14965 17355 14970
rect 17405 14990 17435 14995
rect 17405 14970 17410 14990
rect 17410 14970 17430 14990
rect 17430 14970 17435 14990
rect 17405 14965 17435 14970
rect 17485 14990 17515 14995
rect 17485 14970 17490 14990
rect 17490 14970 17510 14990
rect 17510 14970 17515 14990
rect 17485 14965 17515 14970
rect 17565 14990 17595 14995
rect 17565 14970 17570 14990
rect 17570 14970 17590 14990
rect 17590 14970 17595 14990
rect 17565 14965 17595 14970
rect 17645 14990 17675 14995
rect 17645 14970 17650 14990
rect 17650 14970 17670 14990
rect 17670 14970 17675 14990
rect 17645 14965 17675 14970
rect 17725 14990 17755 14995
rect 17725 14970 17730 14990
rect 17730 14970 17750 14990
rect 17750 14970 17755 14990
rect 17725 14965 17755 14970
rect 17805 14990 17835 14995
rect 17805 14970 17810 14990
rect 17810 14970 17830 14990
rect 17830 14970 17835 14990
rect 17805 14965 17835 14970
rect 17885 14990 17915 14995
rect 17885 14970 17890 14990
rect 17890 14970 17910 14990
rect 17910 14970 17915 14990
rect 17885 14965 17915 14970
rect 17965 14990 17995 14995
rect 17965 14970 17970 14990
rect 17970 14970 17990 14990
rect 17990 14970 17995 14990
rect 17965 14965 17995 14970
rect 18045 14990 18075 14995
rect 18045 14970 18050 14990
rect 18050 14970 18070 14990
rect 18070 14970 18075 14990
rect 18045 14965 18075 14970
rect 18125 14990 18155 14995
rect 18125 14970 18130 14990
rect 18130 14970 18150 14990
rect 18150 14970 18155 14990
rect 18125 14965 18155 14970
rect 18205 14990 18235 14995
rect 18205 14970 18210 14990
rect 18210 14970 18230 14990
rect 18230 14970 18235 14990
rect 18205 14965 18235 14970
rect 18285 14990 18315 14995
rect 18285 14970 18290 14990
rect 18290 14970 18310 14990
rect 18310 14970 18315 14990
rect 18285 14965 18315 14970
rect 18365 14990 18395 14995
rect 18365 14970 18370 14990
rect 18370 14970 18390 14990
rect 18390 14970 18395 14990
rect 18365 14965 18395 14970
rect 18445 14990 18475 14995
rect 18445 14970 18450 14990
rect 18450 14970 18470 14990
rect 18470 14970 18475 14990
rect 18445 14965 18475 14970
rect 18525 14990 18555 14995
rect 18525 14970 18530 14990
rect 18530 14970 18550 14990
rect 18550 14970 18555 14990
rect 18525 14965 18555 14970
rect 18605 14990 18635 14995
rect 18605 14970 18610 14990
rect 18610 14970 18630 14990
rect 18630 14970 18635 14990
rect 18605 14965 18635 14970
rect 18685 14990 18715 14995
rect 18685 14970 18690 14990
rect 18690 14970 18710 14990
rect 18710 14970 18715 14990
rect 18685 14965 18715 14970
rect 18765 14990 18795 14995
rect 18765 14970 18770 14990
rect 18770 14970 18790 14990
rect 18790 14970 18795 14990
rect 18765 14965 18795 14970
rect 18845 14990 18875 14995
rect 18845 14970 18850 14990
rect 18850 14970 18870 14990
rect 18870 14970 18875 14990
rect 18845 14965 18875 14970
rect 18925 14990 18955 14995
rect 18925 14970 18930 14990
rect 18930 14970 18950 14990
rect 18950 14970 18955 14990
rect 18925 14965 18955 14970
rect 19005 14990 19035 14995
rect 19005 14970 19010 14990
rect 19010 14970 19030 14990
rect 19030 14970 19035 14990
rect 19005 14965 19035 14970
rect 19085 14990 19115 14995
rect 19085 14970 19090 14990
rect 19090 14970 19110 14990
rect 19110 14970 19115 14990
rect 19085 14965 19115 14970
rect 19165 14990 19195 14995
rect 19165 14970 19170 14990
rect 19170 14970 19190 14990
rect 19190 14970 19195 14990
rect 19165 14965 19195 14970
rect 19245 14990 19275 14995
rect 19245 14970 19250 14990
rect 19250 14970 19270 14990
rect 19270 14970 19275 14990
rect 19245 14965 19275 14970
rect 19325 14990 19355 14995
rect 19325 14970 19330 14990
rect 19330 14970 19350 14990
rect 19350 14970 19355 14990
rect 19325 14965 19355 14970
rect 19405 14990 19435 14995
rect 19405 14970 19410 14990
rect 19410 14970 19430 14990
rect 19430 14970 19435 14990
rect 19405 14965 19435 14970
rect 19485 14990 19515 14995
rect 19485 14970 19490 14990
rect 19490 14970 19510 14990
rect 19510 14970 19515 14990
rect 19485 14965 19515 14970
rect 19565 14990 19595 14995
rect 19565 14970 19570 14990
rect 19570 14970 19590 14990
rect 19590 14970 19595 14990
rect 19565 14965 19595 14970
rect 19645 14990 19675 14995
rect 19645 14970 19650 14990
rect 19650 14970 19670 14990
rect 19670 14970 19675 14990
rect 19645 14965 19675 14970
rect 19725 14990 19755 14995
rect 19725 14970 19730 14990
rect 19730 14970 19750 14990
rect 19750 14970 19755 14990
rect 19725 14965 19755 14970
rect 19805 14990 19835 14995
rect 19805 14970 19810 14990
rect 19810 14970 19830 14990
rect 19830 14970 19835 14990
rect 19805 14965 19835 14970
rect 19885 14990 19915 14995
rect 19885 14970 19890 14990
rect 19890 14970 19910 14990
rect 19910 14970 19915 14990
rect 19885 14965 19915 14970
rect 19965 14990 19995 14995
rect 19965 14970 19970 14990
rect 19970 14970 19990 14990
rect 19990 14970 19995 14990
rect 19965 14965 19995 14970
rect 20045 14990 20075 14995
rect 20045 14970 20050 14990
rect 20050 14970 20070 14990
rect 20070 14970 20075 14990
rect 20045 14965 20075 14970
rect 20125 14990 20155 14995
rect 20125 14970 20130 14990
rect 20130 14970 20150 14990
rect 20150 14970 20155 14990
rect 20125 14965 20155 14970
rect 20205 14990 20235 14995
rect 20205 14970 20210 14990
rect 20210 14970 20230 14990
rect 20230 14970 20235 14990
rect 20205 14965 20235 14970
rect 20285 14990 20315 14995
rect 20285 14970 20290 14990
rect 20290 14970 20310 14990
rect 20310 14970 20315 14990
rect 20285 14965 20315 14970
rect 20365 14990 20395 14995
rect 20365 14970 20370 14990
rect 20370 14970 20390 14990
rect 20390 14970 20395 14990
rect 20365 14965 20395 14970
rect 20445 14990 20475 14995
rect 20445 14970 20450 14990
rect 20450 14970 20470 14990
rect 20470 14970 20475 14990
rect 20445 14965 20475 14970
rect 20525 14990 20555 14995
rect 20525 14970 20530 14990
rect 20530 14970 20550 14990
rect 20550 14970 20555 14990
rect 20525 14965 20555 14970
rect 20605 14990 20635 14995
rect 20605 14970 20610 14990
rect 20610 14970 20630 14990
rect 20630 14970 20635 14990
rect 20605 14965 20635 14970
rect 20685 14990 20715 14995
rect 20685 14970 20690 14990
rect 20690 14970 20710 14990
rect 20710 14970 20715 14990
rect 20685 14965 20715 14970
rect 20765 14990 20795 14995
rect 20765 14970 20770 14990
rect 20770 14970 20790 14990
rect 20790 14970 20795 14990
rect 20765 14965 20795 14970
rect 20845 14990 20875 14995
rect 20845 14970 20850 14990
rect 20850 14970 20870 14990
rect 20870 14970 20875 14990
rect 20845 14965 20875 14970
rect 20925 14990 20955 14995
rect 20925 14970 20930 14990
rect 20930 14970 20950 14990
rect 20950 14970 20955 14990
rect 20925 14965 20955 14970
rect 5 14910 35 14915
rect 5 14890 10 14910
rect 10 14890 30 14910
rect 30 14890 35 14910
rect 5 14885 35 14890
rect 85 14910 115 14915
rect 85 14890 90 14910
rect 90 14890 110 14910
rect 110 14890 115 14910
rect 85 14885 115 14890
rect 165 14910 195 14915
rect 165 14890 170 14910
rect 170 14890 190 14910
rect 190 14890 195 14910
rect 165 14885 195 14890
rect 245 14910 275 14915
rect 245 14890 250 14910
rect 250 14890 270 14910
rect 270 14890 275 14910
rect 245 14885 275 14890
rect 325 14910 355 14915
rect 325 14890 330 14910
rect 330 14890 350 14910
rect 350 14890 355 14910
rect 325 14885 355 14890
rect 405 14910 435 14915
rect 405 14890 410 14910
rect 410 14890 430 14910
rect 430 14890 435 14910
rect 405 14885 435 14890
rect 485 14910 515 14915
rect 485 14890 490 14910
rect 490 14890 510 14910
rect 510 14890 515 14910
rect 485 14885 515 14890
rect 565 14910 595 14915
rect 565 14890 570 14910
rect 570 14890 590 14910
rect 590 14890 595 14910
rect 565 14885 595 14890
rect 645 14910 675 14915
rect 645 14890 650 14910
rect 650 14890 670 14910
rect 670 14890 675 14910
rect 645 14885 675 14890
rect 725 14910 755 14915
rect 725 14890 730 14910
rect 730 14890 750 14910
rect 750 14890 755 14910
rect 725 14885 755 14890
rect 805 14910 835 14915
rect 805 14890 810 14910
rect 810 14890 830 14910
rect 830 14890 835 14910
rect 805 14885 835 14890
rect 885 14910 915 14915
rect 885 14890 890 14910
rect 890 14890 910 14910
rect 910 14890 915 14910
rect 885 14885 915 14890
rect 965 14910 995 14915
rect 965 14890 970 14910
rect 970 14890 990 14910
rect 990 14890 995 14910
rect 965 14885 995 14890
rect 1045 14910 1075 14915
rect 1045 14890 1050 14910
rect 1050 14890 1070 14910
rect 1070 14890 1075 14910
rect 1045 14885 1075 14890
rect 1125 14910 1155 14915
rect 1125 14890 1130 14910
rect 1130 14890 1150 14910
rect 1150 14890 1155 14910
rect 1125 14885 1155 14890
rect 1205 14910 1235 14915
rect 1205 14890 1210 14910
rect 1210 14890 1230 14910
rect 1230 14890 1235 14910
rect 1205 14885 1235 14890
rect 1285 14910 1315 14915
rect 1285 14890 1290 14910
rect 1290 14890 1310 14910
rect 1310 14890 1315 14910
rect 1285 14885 1315 14890
rect 1365 14910 1395 14915
rect 1365 14890 1370 14910
rect 1370 14890 1390 14910
rect 1390 14890 1395 14910
rect 1365 14885 1395 14890
rect 1445 14910 1475 14915
rect 1445 14890 1450 14910
rect 1450 14890 1470 14910
rect 1470 14890 1475 14910
rect 1445 14885 1475 14890
rect 1525 14910 1555 14915
rect 1525 14890 1530 14910
rect 1530 14890 1550 14910
rect 1550 14890 1555 14910
rect 1525 14885 1555 14890
rect 1605 14910 1635 14915
rect 1605 14890 1610 14910
rect 1610 14890 1630 14910
rect 1630 14890 1635 14910
rect 1605 14885 1635 14890
rect 1685 14910 1715 14915
rect 1685 14890 1690 14910
rect 1690 14890 1710 14910
rect 1710 14890 1715 14910
rect 1685 14885 1715 14890
rect 1765 14910 1795 14915
rect 1765 14890 1770 14910
rect 1770 14890 1790 14910
rect 1790 14890 1795 14910
rect 1765 14885 1795 14890
rect 1845 14910 1875 14915
rect 1845 14890 1850 14910
rect 1850 14890 1870 14910
rect 1870 14890 1875 14910
rect 1845 14885 1875 14890
rect 1925 14910 1955 14915
rect 1925 14890 1930 14910
rect 1930 14890 1950 14910
rect 1950 14890 1955 14910
rect 1925 14885 1955 14890
rect 2005 14910 2035 14915
rect 2005 14890 2010 14910
rect 2010 14890 2030 14910
rect 2030 14890 2035 14910
rect 2005 14885 2035 14890
rect 2085 14910 2115 14915
rect 2085 14890 2090 14910
rect 2090 14890 2110 14910
rect 2110 14890 2115 14910
rect 2085 14885 2115 14890
rect 2165 14910 2195 14915
rect 2165 14890 2170 14910
rect 2170 14890 2190 14910
rect 2190 14890 2195 14910
rect 2165 14885 2195 14890
rect 2245 14910 2275 14915
rect 2245 14890 2250 14910
rect 2250 14890 2270 14910
rect 2270 14890 2275 14910
rect 2245 14885 2275 14890
rect 2325 14910 2355 14915
rect 2325 14890 2330 14910
rect 2330 14890 2350 14910
rect 2350 14890 2355 14910
rect 2325 14885 2355 14890
rect 2405 14910 2435 14915
rect 2405 14890 2410 14910
rect 2410 14890 2430 14910
rect 2430 14890 2435 14910
rect 2405 14885 2435 14890
rect 2485 14910 2515 14915
rect 2485 14890 2490 14910
rect 2490 14890 2510 14910
rect 2510 14890 2515 14910
rect 2485 14885 2515 14890
rect 2565 14910 2595 14915
rect 2565 14890 2570 14910
rect 2570 14890 2590 14910
rect 2590 14890 2595 14910
rect 2565 14885 2595 14890
rect 2645 14910 2675 14915
rect 2645 14890 2650 14910
rect 2650 14890 2670 14910
rect 2670 14890 2675 14910
rect 2645 14885 2675 14890
rect 2725 14910 2755 14915
rect 2725 14890 2730 14910
rect 2730 14890 2750 14910
rect 2750 14890 2755 14910
rect 2725 14885 2755 14890
rect 2805 14910 2835 14915
rect 2805 14890 2810 14910
rect 2810 14890 2830 14910
rect 2830 14890 2835 14910
rect 2805 14885 2835 14890
rect 2885 14910 2915 14915
rect 2885 14890 2890 14910
rect 2890 14890 2910 14910
rect 2910 14890 2915 14910
rect 2885 14885 2915 14890
rect 2965 14910 2995 14915
rect 2965 14890 2970 14910
rect 2970 14890 2990 14910
rect 2990 14890 2995 14910
rect 2965 14885 2995 14890
rect 3045 14910 3075 14915
rect 3045 14890 3050 14910
rect 3050 14890 3070 14910
rect 3070 14890 3075 14910
rect 3045 14885 3075 14890
rect 3125 14910 3155 14915
rect 3125 14890 3130 14910
rect 3130 14890 3150 14910
rect 3150 14890 3155 14910
rect 3125 14885 3155 14890
rect 3205 14910 3235 14915
rect 3205 14890 3210 14910
rect 3210 14890 3230 14910
rect 3230 14890 3235 14910
rect 3205 14885 3235 14890
rect 3285 14910 3315 14915
rect 3285 14890 3290 14910
rect 3290 14890 3310 14910
rect 3310 14890 3315 14910
rect 3285 14885 3315 14890
rect 3365 14910 3395 14915
rect 3365 14890 3370 14910
rect 3370 14890 3390 14910
rect 3390 14890 3395 14910
rect 3365 14885 3395 14890
rect 3445 14910 3475 14915
rect 3445 14890 3450 14910
rect 3450 14890 3470 14910
rect 3470 14890 3475 14910
rect 3445 14885 3475 14890
rect 3525 14910 3555 14915
rect 3525 14890 3530 14910
rect 3530 14890 3550 14910
rect 3550 14890 3555 14910
rect 3525 14885 3555 14890
rect 3605 14910 3635 14915
rect 3605 14890 3610 14910
rect 3610 14890 3630 14910
rect 3630 14890 3635 14910
rect 3605 14885 3635 14890
rect 3685 14910 3715 14915
rect 3685 14890 3690 14910
rect 3690 14890 3710 14910
rect 3710 14890 3715 14910
rect 3685 14885 3715 14890
rect 3765 14910 3795 14915
rect 3765 14890 3770 14910
rect 3770 14890 3790 14910
rect 3790 14890 3795 14910
rect 3765 14885 3795 14890
rect 3845 14910 3875 14915
rect 3845 14890 3850 14910
rect 3850 14890 3870 14910
rect 3870 14890 3875 14910
rect 3845 14885 3875 14890
rect 3925 14910 3955 14915
rect 3925 14890 3930 14910
rect 3930 14890 3950 14910
rect 3950 14890 3955 14910
rect 3925 14885 3955 14890
rect 4005 14910 4035 14915
rect 4005 14890 4010 14910
rect 4010 14890 4030 14910
rect 4030 14890 4035 14910
rect 4005 14885 4035 14890
rect 4085 14910 4115 14915
rect 4085 14890 4090 14910
rect 4090 14890 4110 14910
rect 4110 14890 4115 14910
rect 4085 14885 4115 14890
rect 4165 14910 4195 14915
rect 4165 14890 4170 14910
rect 4170 14890 4190 14910
rect 4190 14890 4195 14910
rect 4165 14885 4195 14890
rect 6245 14910 6275 14915
rect 6245 14890 6250 14910
rect 6250 14890 6270 14910
rect 6270 14890 6275 14910
rect 6245 14885 6275 14890
rect 6325 14910 6355 14915
rect 6325 14890 6330 14910
rect 6330 14890 6350 14910
rect 6350 14890 6355 14910
rect 6325 14885 6355 14890
rect 6405 14910 6435 14915
rect 6405 14890 6410 14910
rect 6410 14890 6430 14910
rect 6430 14890 6435 14910
rect 6405 14885 6435 14890
rect 6485 14910 6515 14915
rect 6485 14890 6490 14910
rect 6490 14890 6510 14910
rect 6510 14890 6515 14910
rect 6485 14885 6515 14890
rect 6565 14910 6595 14915
rect 6565 14890 6570 14910
rect 6570 14890 6590 14910
rect 6590 14890 6595 14910
rect 6565 14885 6595 14890
rect 6645 14910 6675 14915
rect 6645 14890 6650 14910
rect 6650 14890 6670 14910
rect 6670 14890 6675 14910
rect 6645 14885 6675 14890
rect 6725 14910 6755 14915
rect 6725 14890 6730 14910
rect 6730 14890 6750 14910
rect 6750 14890 6755 14910
rect 6725 14885 6755 14890
rect 6805 14910 6835 14915
rect 6805 14890 6810 14910
rect 6810 14890 6830 14910
rect 6830 14890 6835 14910
rect 6805 14885 6835 14890
rect 6885 14910 6915 14915
rect 6885 14890 6890 14910
rect 6890 14890 6910 14910
rect 6910 14890 6915 14910
rect 6885 14885 6915 14890
rect 6965 14910 6995 14915
rect 6965 14890 6970 14910
rect 6970 14890 6990 14910
rect 6990 14890 6995 14910
rect 6965 14885 6995 14890
rect 7045 14910 7075 14915
rect 7045 14890 7050 14910
rect 7050 14890 7070 14910
rect 7070 14890 7075 14910
rect 7045 14885 7075 14890
rect 7125 14910 7155 14915
rect 7125 14890 7130 14910
rect 7130 14890 7150 14910
rect 7150 14890 7155 14910
rect 7125 14885 7155 14890
rect 7205 14910 7235 14915
rect 7205 14890 7210 14910
rect 7210 14890 7230 14910
rect 7230 14890 7235 14910
rect 7205 14885 7235 14890
rect 7285 14910 7315 14915
rect 7285 14890 7290 14910
rect 7290 14890 7310 14910
rect 7310 14890 7315 14910
rect 7285 14885 7315 14890
rect 7365 14910 7395 14915
rect 7365 14890 7370 14910
rect 7370 14890 7390 14910
rect 7390 14890 7395 14910
rect 7365 14885 7395 14890
rect 7445 14910 7475 14915
rect 7445 14890 7450 14910
rect 7450 14890 7470 14910
rect 7470 14890 7475 14910
rect 7445 14885 7475 14890
rect 7525 14910 7555 14915
rect 7525 14890 7530 14910
rect 7530 14890 7550 14910
rect 7550 14890 7555 14910
rect 7525 14885 7555 14890
rect 7605 14910 7635 14915
rect 7605 14890 7610 14910
rect 7610 14890 7630 14910
rect 7630 14890 7635 14910
rect 7605 14885 7635 14890
rect 7685 14910 7715 14915
rect 7685 14890 7690 14910
rect 7690 14890 7710 14910
rect 7710 14890 7715 14910
rect 7685 14885 7715 14890
rect 7765 14910 7795 14915
rect 7765 14890 7770 14910
rect 7770 14890 7790 14910
rect 7790 14890 7795 14910
rect 7765 14885 7795 14890
rect 7845 14910 7875 14915
rect 7845 14890 7850 14910
rect 7850 14890 7870 14910
rect 7870 14890 7875 14910
rect 7845 14885 7875 14890
rect 7925 14910 7955 14915
rect 7925 14890 7930 14910
rect 7930 14890 7950 14910
rect 7950 14890 7955 14910
rect 7925 14885 7955 14890
rect 8005 14910 8035 14915
rect 8005 14890 8010 14910
rect 8010 14890 8030 14910
rect 8030 14890 8035 14910
rect 8005 14885 8035 14890
rect 8085 14910 8115 14915
rect 8085 14890 8090 14910
rect 8090 14890 8110 14910
rect 8110 14890 8115 14910
rect 8085 14885 8115 14890
rect 8165 14910 8195 14915
rect 8165 14890 8170 14910
rect 8170 14890 8190 14910
rect 8190 14890 8195 14910
rect 8165 14885 8195 14890
rect 8245 14910 8275 14915
rect 8245 14890 8250 14910
rect 8250 14890 8270 14910
rect 8270 14890 8275 14910
rect 8245 14885 8275 14890
rect 8325 14910 8355 14915
rect 8325 14890 8330 14910
rect 8330 14890 8350 14910
rect 8350 14890 8355 14910
rect 8325 14885 8355 14890
rect 8405 14910 8435 14915
rect 8405 14890 8410 14910
rect 8410 14890 8430 14910
rect 8430 14890 8435 14910
rect 8405 14885 8435 14890
rect 8485 14910 8515 14915
rect 8485 14890 8490 14910
rect 8490 14890 8510 14910
rect 8510 14890 8515 14910
rect 8485 14885 8515 14890
rect 8565 14910 8595 14915
rect 8565 14890 8570 14910
rect 8570 14890 8590 14910
rect 8590 14890 8595 14910
rect 8565 14885 8595 14890
rect 8645 14910 8675 14915
rect 8645 14890 8650 14910
rect 8650 14890 8670 14910
rect 8670 14890 8675 14910
rect 8645 14885 8675 14890
rect 8725 14910 8755 14915
rect 8725 14890 8730 14910
rect 8730 14890 8750 14910
rect 8750 14890 8755 14910
rect 8725 14885 8755 14890
rect 8805 14910 8835 14915
rect 8805 14890 8810 14910
rect 8810 14890 8830 14910
rect 8830 14890 8835 14910
rect 8805 14885 8835 14890
rect 8885 14910 8915 14915
rect 8885 14890 8890 14910
rect 8890 14890 8910 14910
rect 8910 14890 8915 14910
rect 8885 14885 8915 14890
rect 8965 14910 8995 14915
rect 8965 14890 8970 14910
rect 8970 14890 8990 14910
rect 8990 14890 8995 14910
rect 8965 14885 8995 14890
rect 9045 14910 9075 14915
rect 9045 14890 9050 14910
rect 9050 14890 9070 14910
rect 9070 14890 9075 14910
rect 9045 14885 9075 14890
rect 9125 14910 9155 14915
rect 9125 14890 9130 14910
rect 9130 14890 9150 14910
rect 9150 14890 9155 14910
rect 9125 14885 9155 14890
rect 9205 14910 9235 14915
rect 9205 14890 9210 14910
rect 9210 14890 9230 14910
rect 9230 14890 9235 14910
rect 9205 14885 9235 14890
rect 9285 14910 9315 14915
rect 9285 14890 9290 14910
rect 9290 14890 9310 14910
rect 9310 14890 9315 14910
rect 9285 14885 9315 14890
rect 9365 14910 9395 14915
rect 9365 14890 9370 14910
rect 9370 14890 9390 14910
rect 9390 14890 9395 14910
rect 9365 14885 9395 14890
rect 9445 14910 9475 14915
rect 9445 14890 9450 14910
rect 9450 14890 9470 14910
rect 9470 14890 9475 14910
rect 9445 14885 9475 14890
rect 11565 14910 11595 14915
rect 11565 14890 11570 14910
rect 11570 14890 11590 14910
rect 11590 14890 11595 14910
rect 11565 14885 11595 14890
rect 11645 14910 11675 14915
rect 11645 14890 11650 14910
rect 11650 14890 11670 14910
rect 11670 14890 11675 14910
rect 11645 14885 11675 14890
rect 11725 14910 11755 14915
rect 11725 14890 11730 14910
rect 11730 14890 11750 14910
rect 11750 14890 11755 14910
rect 11725 14885 11755 14890
rect 11805 14910 11835 14915
rect 11805 14890 11810 14910
rect 11810 14890 11830 14910
rect 11830 14890 11835 14910
rect 11805 14885 11835 14890
rect 11885 14910 11915 14915
rect 11885 14890 11890 14910
rect 11890 14890 11910 14910
rect 11910 14890 11915 14910
rect 11885 14885 11915 14890
rect 11965 14910 11995 14915
rect 11965 14890 11970 14910
rect 11970 14890 11990 14910
rect 11990 14890 11995 14910
rect 11965 14885 11995 14890
rect 12045 14910 12075 14915
rect 12045 14890 12050 14910
rect 12050 14890 12070 14910
rect 12070 14890 12075 14910
rect 12045 14885 12075 14890
rect 12125 14910 12155 14915
rect 12125 14890 12130 14910
rect 12130 14890 12150 14910
rect 12150 14890 12155 14910
rect 12125 14885 12155 14890
rect 12205 14910 12235 14915
rect 12205 14890 12210 14910
rect 12210 14890 12230 14910
rect 12230 14890 12235 14910
rect 12205 14885 12235 14890
rect 12285 14910 12315 14915
rect 12285 14890 12290 14910
rect 12290 14890 12310 14910
rect 12310 14890 12315 14910
rect 12285 14885 12315 14890
rect 12365 14910 12395 14915
rect 12365 14890 12370 14910
rect 12370 14890 12390 14910
rect 12390 14890 12395 14910
rect 12365 14885 12395 14890
rect 12445 14910 12475 14915
rect 12445 14890 12450 14910
rect 12450 14890 12470 14910
rect 12470 14890 12475 14910
rect 12445 14885 12475 14890
rect 12525 14910 12555 14915
rect 12525 14890 12530 14910
rect 12530 14890 12550 14910
rect 12550 14890 12555 14910
rect 12525 14885 12555 14890
rect 12605 14910 12635 14915
rect 12605 14890 12610 14910
rect 12610 14890 12630 14910
rect 12630 14890 12635 14910
rect 12605 14885 12635 14890
rect 12685 14910 12715 14915
rect 12685 14890 12690 14910
rect 12690 14890 12710 14910
rect 12710 14890 12715 14910
rect 12685 14885 12715 14890
rect 12765 14910 12795 14915
rect 12765 14890 12770 14910
rect 12770 14890 12790 14910
rect 12790 14890 12795 14910
rect 12765 14885 12795 14890
rect 12845 14910 12875 14915
rect 12845 14890 12850 14910
rect 12850 14890 12870 14910
rect 12870 14890 12875 14910
rect 12845 14885 12875 14890
rect 12925 14910 12955 14915
rect 12925 14890 12930 14910
rect 12930 14890 12950 14910
rect 12950 14890 12955 14910
rect 12925 14885 12955 14890
rect 13005 14910 13035 14915
rect 13005 14890 13010 14910
rect 13010 14890 13030 14910
rect 13030 14890 13035 14910
rect 13005 14885 13035 14890
rect 13085 14910 13115 14915
rect 13085 14890 13090 14910
rect 13090 14890 13110 14910
rect 13110 14890 13115 14910
rect 13085 14885 13115 14890
rect 13165 14910 13195 14915
rect 13165 14890 13170 14910
rect 13170 14890 13190 14910
rect 13190 14890 13195 14910
rect 13165 14885 13195 14890
rect 13245 14910 13275 14915
rect 13245 14890 13250 14910
rect 13250 14890 13270 14910
rect 13270 14890 13275 14910
rect 13245 14885 13275 14890
rect 13325 14910 13355 14915
rect 13325 14890 13330 14910
rect 13330 14890 13350 14910
rect 13350 14890 13355 14910
rect 13325 14885 13355 14890
rect 13405 14910 13435 14915
rect 13405 14890 13410 14910
rect 13410 14890 13430 14910
rect 13430 14890 13435 14910
rect 13405 14885 13435 14890
rect 13485 14910 13515 14915
rect 13485 14890 13490 14910
rect 13490 14890 13510 14910
rect 13510 14890 13515 14910
rect 13485 14885 13515 14890
rect 13565 14910 13595 14915
rect 13565 14890 13570 14910
rect 13570 14890 13590 14910
rect 13590 14890 13595 14910
rect 13565 14885 13595 14890
rect 13645 14910 13675 14915
rect 13645 14890 13650 14910
rect 13650 14890 13670 14910
rect 13670 14890 13675 14910
rect 13645 14885 13675 14890
rect 13725 14910 13755 14915
rect 13725 14890 13730 14910
rect 13730 14890 13750 14910
rect 13750 14890 13755 14910
rect 13725 14885 13755 14890
rect 13805 14910 13835 14915
rect 13805 14890 13810 14910
rect 13810 14890 13830 14910
rect 13830 14890 13835 14910
rect 13805 14885 13835 14890
rect 13885 14910 13915 14915
rect 13885 14890 13890 14910
rect 13890 14890 13910 14910
rect 13910 14890 13915 14910
rect 13885 14885 13915 14890
rect 13965 14910 13995 14915
rect 13965 14890 13970 14910
rect 13970 14890 13990 14910
rect 13990 14890 13995 14910
rect 13965 14885 13995 14890
rect 14045 14910 14075 14915
rect 14045 14890 14050 14910
rect 14050 14890 14070 14910
rect 14070 14890 14075 14910
rect 14045 14885 14075 14890
rect 14125 14910 14155 14915
rect 14125 14890 14130 14910
rect 14130 14890 14150 14910
rect 14150 14890 14155 14910
rect 14125 14885 14155 14890
rect 14205 14910 14235 14915
rect 14205 14890 14210 14910
rect 14210 14890 14230 14910
rect 14230 14890 14235 14910
rect 14205 14885 14235 14890
rect 14285 14910 14315 14915
rect 14285 14890 14290 14910
rect 14290 14890 14310 14910
rect 14310 14890 14315 14910
rect 14285 14885 14315 14890
rect 14365 14910 14395 14915
rect 14365 14890 14370 14910
rect 14370 14890 14390 14910
rect 14390 14890 14395 14910
rect 14365 14885 14395 14890
rect 14445 14910 14475 14915
rect 14445 14890 14450 14910
rect 14450 14890 14470 14910
rect 14470 14890 14475 14910
rect 14445 14885 14475 14890
rect 14525 14910 14555 14915
rect 14525 14890 14530 14910
rect 14530 14890 14550 14910
rect 14550 14890 14555 14910
rect 14525 14885 14555 14890
rect 14605 14910 14635 14915
rect 14605 14890 14610 14910
rect 14610 14890 14630 14910
rect 14630 14890 14635 14910
rect 14605 14885 14635 14890
rect 14685 14910 14715 14915
rect 14685 14890 14690 14910
rect 14690 14890 14710 14910
rect 14710 14890 14715 14910
rect 14685 14885 14715 14890
rect 16765 14910 16795 14915
rect 16765 14890 16770 14910
rect 16770 14890 16790 14910
rect 16790 14890 16795 14910
rect 16765 14885 16795 14890
rect 16845 14910 16875 14915
rect 16845 14890 16850 14910
rect 16850 14890 16870 14910
rect 16870 14890 16875 14910
rect 16845 14885 16875 14890
rect 16925 14910 16955 14915
rect 16925 14890 16930 14910
rect 16930 14890 16950 14910
rect 16950 14890 16955 14910
rect 16925 14885 16955 14890
rect 17005 14910 17035 14915
rect 17005 14890 17010 14910
rect 17010 14890 17030 14910
rect 17030 14890 17035 14910
rect 17005 14885 17035 14890
rect 17085 14910 17115 14915
rect 17085 14890 17090 14910
rect 17090 14890 17110 14910
rect 17110 14890 17115 14910
rect 17085 14885 17115 14890
rect 17165 14910 17195 14915
rect 17165 14890 17170 14910
rect 17170 14890 17190 14910
rect 17190 14890 17195 14910
rect 17165 14885 17195 14890
rect 17245 14910 17275 14915
rect 17245 14890 17250 14910
rect 17250 14890 17270 14910
rect 17270 14890 17275 14910
rect 17245 14885 17275 14890
rect 17325 14910 17355 14915
rect 17325 14890 17330 14910
rect 17330 14890 17350 14910
rect 17350 14890 17355 14910
rect 17325 14885 17355 14890
rect 17405 14910 17435 14915
rect 17405 14890 17410 14910
rect 17410 14890 17430 14910
rect 17430 14890 17435 14910
rect 17405 14885 17435 14890
rect 17485 14910 17515 14915
rect 17485 14890 17490 14910
rect 17490 14890 17510 14910
rect 17510 14890 17515 14910
rect 17485 14885 17515 14890
rect 17565 14910 17595 14915
rect 17565 14890 17570 14910
rect 17570 14890 17590 14910
rect 17590 14890 17595 14910
rect 17565 14885 17595 14890
rect 17645 14910 17675 14915
rect 17645 14890 17650 14910
rect 17650 14890 17670 14910
rect 17670 14890 17675 14910
rect 17645 14885 17675 14890
rect 17725 14910 17755 14915
rect 17725 14890 17730 14910
rect 17730 14890 17750 14910
rect 17750 14890 17755 14910
rect 17725 14885 17755 14890
rect 17805 14910 17835 14915
rect 17805 14890 17810 14910
rect 17810 14890 17830 14910
rect 17830 14890 17835 14910
rect 17805 14885 17835 14890
rect 17885 14910 17915 14915
rect 17885 14890 17890 14910
rect 17890 14890 17910 14910
rect 17910 14890 17915 14910
rect 17885 14885 17915 14890
rect 17965 14910 17995 14915
rect 17965 14890 17970 14910
rect 17970 14890 17990 14910
rect 17990 14890 17995 14910
rect 17965 14885 17995 14890
rect 18045 14910 18075 14915
rect 18045 14890 18050 14910
rect 18050 14890 18070 14910
rect 18070 14890 18075 14910
rect 18045 14885 18075 14890
rect 18125 14910 18155 14915
rect 18125 14890 18130 14910
rect 18130 14890 18150 14910
rect 18150 14890 18155 14910
rect 18125 14885 18155 14890
rect 18205 14910 18235 14915
rect 18205 14890 18210 14910
rect 18210 14890 18230 14910
rect 18230 14890 18235 14910
rect 18205 14885 18235 14890
rect 18285 14910 18315 14915
rect 18285 14890 18290 14910
rect 18290 14890 18310 14910
rect 18310 14890 18315 14910
rect 18285 14885 18315 14890
rect 18365 14910 18395 14915
rect 18365 14890 18370 14910
rect 18370 14890 18390 14910
rect 18390 14890 18395 14910
rect 18365 14885 18395 14890
rect 18445 14910 18475 14915
rect 18445 14890 18450 14910
rect 18450 14890 18470 14910
rect 18470 14890 18475 14910
rect 18445 14885 18475 14890
rect 18525 14910 18555 14915
rect 18525 14890 18530 14910
rect 18530 14890 18550 14910
rect 18550 14890 18555 14910
rect 18525 14885 18555 14890
rect 18605 14910 18635 14915
rect 18605 14890 18610 14910
rect 18610 14890 18630 14910
rect 18630 14890 18635 14910
rect 18605 14885 18635 14890
rect 18685 14910 18715 14915
rect 18685 14890 18690 14910
rect 18690 14890 18710 14910
rect 18710 14890 18715 14910
rect 18685 14885 18715 14890
rect 18765 14910 18795 14915
rect 18765 14890 18770 14910
rect 18770 14890 18790 14910
rect 18790 14890 18795 14910
rect 18765 14885 18795 14890
rect 18845 14910 18875 14915
rect 18845 14890 18850 14910
rect 18850 14890 18870 14910
rect 18870 14890 18875 14910
rect 18845 14885 18875 14890
rect 18925 14910 18955 14915
rect 18925 14890 18930 14910
rect 18930 14890 18950 14910
rect 18950 14890 18955 14910
rect 18925 14885 18955 14890
rect 19005 14910 19035 14915
rect 19005 14890 19010 14910
rect 19010 14890 19030 14910
rect 19030 14890 19035 14910
rect 19005 14885 19035 14890
rect 19085 14910 19115 14915
rect 19085 14890 19090 14910
rect 19090 14890 19110 14910
rect 19110 14890 19115 14910
rect 19085 14885 19115 14890
rect 19165 14910 19195 14915
rect 19165 14890 19170 14910
rect 19170 14890 19190 14910
rect 19190 14890 19195 14910
rect 19165 14885 19195 14890
rect 19245 14910 19275 14915
rect 19245 14890 19250 14910
rect 19250 14890 19270 14910
rect 19270 14890 19275 14910
rect 19245 14885 19275 14890
rect 19325 14910 19355 14915
rect 19325 14890 19330 14910
rect 19330 14890 19350 14910
rect 19350 14890 19355 14910
rect 19325 14885 19355 14890
rect 19405 14910 19435 14915
rect 19405 14890 19410 14910
rect 19410 14890 19430 14910
rect 19430 14890 19435 14910
rect 19405 14885 19435 14890
rect 19485 14910 19515 14915
rect 19485 14890 19490 14910
rect 19490 14890 19510 14910
rect 19510 14890 19515 14910
rect 19485 14885 19515 14890
rect 19565 14910 19595 14915
rect 19565 14890 19570 14910
rect 19570 14890 19590 14910
rect 19590 14890 19595 14910
rect 19565 14885 19595 14890
rect 19645 14910 19675 14915
rect 19645 14890 19650 14910
rect 19650 14890 19670 14910
rect 19670 14890 19675 14910
rect 19645 14885 19675 14890
rect 19725 14910 19755 14915
rect 19725 14890 19730 14910
rect 19730 14890 19750 14910
rect 19750 14890 19755 14910
rect 19725 14885 19755 14890
rect 19805 14910 19835 14915
rect 19805 14890 19810 14910
rect 19810 14890 19830 14910
rect 19830 14890 19835 14910
rect 19805 14885 19835 14890
rect 19885 14910 19915 14915
rect 19885 14890 19890 14910
rect 19890 14890 19910 14910
rect 19910 14890 19915 14910
rect 19885 14885 19915 14890
rect 19965 14910 19995 14915
rect 19965 14890 19970 14910
rect 19970 14890 19990 14910
rect 19990 14890 19995 14910
rect 19965 14885 19995 14890
rect 20045 14910 20075 14915
rect 20045 14890 20050 14910
rect 20050 14890 20070 14910
rect 20070 14890 20075 14910
rect 20045 14885 20075 14890
rect 20125 14910 20155 14915
rect 20125 14890 20130 14910
rect 20130 14890 20150 14910
rect 20150 14890 20155 14910
rect 20125 14885 20155 14890
rect 20205 14910 20235 14915
rect 20205 14890 20210 14910
rect 20210 14890 20230 14910
rect 20230 14890 20235 14910
rect 20205 14885 20235 14890
rect 20285 14910 20315 14915
rect 20285 14890 20290 14910
rect 20290 14890 20310 14910
rect 20310 14890 20315 14910
rect 20285 14885 20315 14890
rect 20365 14910 20395 14915
rect 20365 14890 20370 14910
rect 20370 14890 20390 14910
rect 20390 14890 20395 14910
rect 20365 14885 20395 14890
rect 20445 14910 20475 14915
rect 20445 14890 20450 14910
rect 20450 14890 20470 14910
rect 20470 14890 20475 14910
rect 20445 14885 20475 14890
rect 20525 14910 20555 14915
rect 20525 14890 20530 14910
rect 20530 14890 20550 14910
rect 20550 14890 20555 14910
rect 20525 14885 20555 14890
rect 20605 14910 20635 14915
rect 20605 14890 20610 14910
rect 20610 14890 20630 14910
rect 20630 14890 20635 14910
rect 20605 14885 20635 14890
rect 20685 14910 20715 14915
rect 20685 14890 20690 14910
rect 20690 14890 20710 14910
rect 20710 14890 20715 14910
rect 20685 14885 20715 14890
rect 20765 14910 20795 14915
rect 20765 14890 20770 14910
rect 20770 14890 20790 14910
rect 20790 14890 20795 14910
rect 20765 14885 20795 14890
rect 20845 14910 20875 14915
rect 20845 14890 20850 14910
rect 20850 14890 20870 14910
rect 20870 14890 20875 14910
rect 20845 14885 20875 14890
rect 20925 14910 20955 14915
rect 20925 14890 20930 14910
rect 20930 14890 20950 14910
rect 20950 14890 20955 14910
rect 20925 14885 20955 14890
rect 5 14750 35 14755
rect 5 14730 10 14750
rect 10 14730 30 14750
rect 30 14730 35 14750
rect 5 14725 35 14730
rect 85 14750 115 14755
rect 85 14730 90 14750
rect 90 14730 110 14750
rect 110 14730 115 14750
rect 85 14725 115 14730
rect 165 14750 195 14755
rect 165 14730 170 14750
rect 170 14730 190 14750
rect 190 14730 195 14750
rect 165 14725 195 14730
rect 245 14750 275 14755
rect 245 14730 250 14750
rect 250 14730 270 14750
rect 270 14730 275 14750
rect 245 14725 275 14730
rect 325 14750 355 14755
rect 325 14730 330 14750
rect 330 14730 350 14750
rect 350 14730 355 14750
rect 325 14725 355 14730
rect 405 14750 435 14755
rect 405 14730 410 14750
rect 410 14730 430 14750
rect 430 14730 435 14750
rect 405 14725 435 14730
rect 485 14750 515 14755
rect 485 14730 490 14750
rect 490 14730 510 14750
rect 510 14730 515 14750
rect 485 14725 515 14730
rect 565 14750 595 14755
rect 565 14730 570 14750
rect 570 14730 590 14750
rect 590 14730 595 14750
rect 565 14725 595 14730
rect 645 14750 675 14755
rect 645 14730 650 14750
rect 650 14730 670 14750
rect 670 14730 675 14750
rect 645 14725 675 14730
rect 725 14750 755 14755
rect 725 14730 730 14750
rect 730 14730 750 14750
rect 750 14730 755 14750
rect 725 14725 755 14730
rect 805 14750 835 14755
rect 805 14730 810 14750
rect 810 14730 830 14750
rect 830 14730 835 14750
rect 805 14725 835 14730
rect 885 14750 915 14755
rect 885 14730 890 14750
rect 890 14730 910 14750
rect 910 14730 915 14750
rect 885 14725 915 14730
rect 965 14750 995 14755
rect 965 14730 970 14750
rect 970 14730 990 14750
rect 990 14730 995 14750
rect 965 14725 995 14730
rect 1045 14750 1075 14755
rect 1045 14730 1050 14750
rect 1050 14730 1070 14750
rect 1070 14730 1075 14750
rect 1045 14725 1075 14730
rect 1125 14750 1155 14755
rect 1125 14730 1130 14750
rect 1130 14730 1150 14750
rect 1150 14730 1155 14750
rect 1125 14725 1155 14730
rect 1205 14750 1235 14755
rect 1205 14730 1210 14750
rect 1210 14730 1230 14750
rect 1230 14730 1235 14750
rect 1205 14725 1235 14730
rect 1285 14750 1315 14755
rect 1285 14730 1290 14750
rect 1290 14730 1310 14750
rect 1310 14730 1315 14750
rect 1285 14725 1315 14730
rect 1365 14750 1395 14755
rect 1365 14730 1370 14750
rect 1370 14730 1390 14750
rect 1390 14730 1395 14750
rect 1365 14725 1395 14730
rect 1445 14750 1475 14755
rect 1445 14730 1450 14750
rect 1450 14730 1470 14750
rect 1470 14730 1475 14750
rect 1445 14725 1475 14730
rect 1525 14750 1555 14755
rect 1525 14730 1530 14750
rect 1530 14730 1550 14750
rect 1550 14730 1555 14750
rect 1525 14725 1555 14730
rect 1605 14750 1635 14755
rect 1605 14730 1610 14750
rect 1610 14730 1630 14750
rect 1630 14730 1635 14750
rect 1605 14725 1635 14730
rect 1685 14750 1715 14755
rect 1685 14730 1690 14750
rect 1690 14730 1710 14750
rect 1710 14730 1715 14750
rect 1685 14725 1715 14730
rect 1765 14750 1795 14755
rect 1765 14730 1770 14750
rect 1770 14730 1790 14750
rect 1790 14730 1795 14750
rect 1765 14725 1795 14730
rect 1845 14750 1875 14755
rect 1845 14730 1850 14750
rect 1850 14730 1870 14750
rect 1870 14730 1875 14750
rect 1845 14725 1875 14730
rect 1925 14750 1955 14755
rect 1925 14730 1930 14750
rect 1930 14730 1950 14750
rect 1950 14730 1955 14750
rect 1925 14725 1955 14730
rect 2005 14750 2035 14755
rect 2005 14730 2010 14750
rect 2010 14730 2030 14750
rect 2030 14730 2035 14750
rect 2005 14725 2035 14730
rect 2085 14750 2115 14755
rect 2085 14730 2090 14750
rect 2090 14730 2110 14750
rect 2110 14730 2115 14750
rect 2085 14725 2115 14730
rect 2165 14750 2195 14755
rect 2165 14730 2170 14750
rect 2170 14730 2190 14750
rect 2190 14730 2195 14750
rect 2165 14725 2195 14730
rect 2245 14750 2275 14755
rect 2245 14730 2250 14750
rect 2250 14730 2270 14750
rect 2270 14730 2275 14750
rect 2245 14725 2275 14730
rect 2325 14750 2355 14755
rect 2325 14730 2330 14750
rect 2330 14730 2350 14750
rect 2350 14730 2355 14750
rect 2325 14725 2355 14730
rect 2405 14750 2435 14755
rect 2405 14730 2410 14750
rect 2410 14730 2430 14750
rect 2430 14730 2435 14750
rect 2405 14725 2435 14730
rect 2485 14750 2515 14755
rect 2485 14730 2490 14750
rect 2490 14730 2510 14750
rect 2510 14730 2515 14750
rect 2485 14725 2515 14730
rect 2565 14750 2595 14755
rect 2565 14730 2570 14750
rect 2570 14730 2590 14750
rect 2590 14730 2595 14750
rect 2565 14725 2595 14730
rect 2645 14750 2675 14755
rect 2645 14730 2650 14750
rect 2650 14730 2670 14750
rect 2670 14730 2675 14750
rect 2645 14725 2675 14730
rect 2725 14750 2755 14755
rect 2725 14730 2730 14750
rect 2730 14730 2750 14750
rect 2750 14730 2755 14750
rect 2725 14725 2755 14730
rect 2805 14750 2835 14755
rect 2805 14730 2810 14750
rect 2810 14730 2830 14750
rect 2830 14730 2835 14750
rect 2805 14725 2835 14730
rect 2885 14750 2915 14755
rect 2885 14730 2890 14750
rect 2890 14730 2910 14750
rect 2910 14730 2915 14750
rect 2885 14725 2915 14730
rect 2965 14750 2995 14755
rect 2965 14730 2970 14750
rect 2970 14730 2990 14750
rect 2990 14730 2995 14750
rect 2965 14725 2995 14730
rect 3045 14750 3075 14755
rect 3045 14730 3050 14750
rect 3050 14730 3070 14750
rect 3070 14730 3075 14750
rect 3045 14725 3075 14730
rect 3125 14750 3155 14755
rect 3125 14730 3130 14750
rect 3130 14730 3150 14750
rect 3150 14730 3155 14750
rect 3125 14725 3155 14730
rect 3205 14750 3235 14755
rect 3205 14730 3210 14750
rect 3210 14730 3230 14750
rect 3230 14730 3235 14750
rect 3205 14725 3235 14730
rect 3285 14750 3315 14755
rect 3285 14730 3290 14750
rect 3290 14730 3310 14750
rect 3310 14730 3315 14750
rect 3285 14725 3315 14730
rect 3365 14750 3395 14755
rect 3365 14730 3370 14750
rect 3370 14730 3390 14750
rect 3390 14730 3395 14750
rect 3365 14725 3395 14730
rect 3445 14750 3475 14755
rect 3445 14730 3450 14750
rect 3450 14730 3470 14750
rect 3470 14730 3475 14750
rect 3445 14725 3475 14730
rect 3525 14750 3555 14755
rect 3525 14730 3530 14750
rect 3530 14730 3550 14750
rect 3550 14730 3555 14750
rect 3525 14725 3555 14730
rect 3605 14750 3635 14755
rect 3605 14730 3610 14750
rect 3610 14730 3630 14750
rect 3630 14730 3635 14750
rect 3605 14725 3635 14730
rect 3685 14750 3715 14755
rect 3685 14730 3690 14750
rect 3690 14730 3710 14750
rect 3710 14730 3715 14750
rect 3685 14725 3715 14730
rect 3765 14750 3795 14755
rect 3765 14730 3770 14750
rect 3770 14730 3790 14750
rect 3790 14730 3795 14750
rect 3765 14725 3795 14730
rect 3845 14750 3875 14755
rect 3845 14730 3850 14750
rect 3850 14730 3870 14750
rect 3870 14730 3875 14750
rect 3845 14725 3875 14730
rect 3925 14750 3955 14755
rect 3925 14730 3930 14750
rect 3930 14730 3950 14750
rect 3950 14730 3955 14750
rect 3925 14725 3955 14730
rect 4005 14750 4035 14755
rect 4005 14730 4010 14750
rect 4010 14730 4030 14750
rect 4030 14730 4035 14750
rect 4005 14725 4035 14730
rect 4085 14750 4115 14755
rect 4085 14730 4090 14750
rect 4090 14730 4110 14750
rect 4110 14730 4115 14750
rect 4085 14725 4115 14730
rect 4165 14750 4195 14755
rect 4165 14730 4170 14750
rect 4170 14730 4190 14750
rect 4190 14730 4195 14750
rect 4165 14725 4195 14730
rect 6245 14750 6275 14755
rect 6245 14730 6250 14750
rect 6250 14730 6270 14750
rect 6270 14730 6275 14750
rect 6245 14725 6275 14730
rect 6325 14750 6355 14755
rect 6325 14730 6330 14750
rect 6330 14730 6350 14750
rect 6350 14730 6355 14750
rect 6325 14725 6355 14730
rect 6405 14750 6435 14755
rect 6405 14730 6410 14750
rect 6410 14730 6430 14750
rect 6430 14730 6435 14750
rect 6405 14725 6435 14730
rect 6485 14750 6515 14755
rect 6485 14730 6490 14750
rect 6490 14730 6510 14750
rect 6510 14730 6515 14750
rect 6485 14725 6515 14730
rect 6565 14750 6595 14755
rect 6565 14730 6570 14750
rect 6570 14730 6590 14750
rect 6590 14730 6595 14750
rect 6565 14725 6595 14730
rect 6645 14750 6675 14755
rect 6645 14730 6650 14750
rect 6650 14730 6670 14750
rect 6670 14730 6675 14750
rect 6645 14725 6675 14730
rect 6725 14750 6755 14755
rect 6725 14730 6730 14750
rect 6730 14730 6750 14750
rect 6750 14730 6755 14750
rect 6725 14725 6755 14730
rect 6805 14750 6835 14755
rect 6805 14730 6810 14750
rect 6810 14730 6830 14750
rect 6830 14730 6835 14750
rect 6805 14725 6835 14730
rect 6885 14750 6915 14755
rect 6885 14730 6890 14750
rect 6890 14730 6910 14750
rect 6910 14730 6915 14750
rect 6885 14725 6915 14730
rect 6965 14750 6995 14755
rect 6965 14730 6970 14750
rect 6970 14730 6990 14750
rect 6990 14730 6995 14750
rect 6965 14725 6995 14730
rect 7045 14750 7075 14755
rect 7045 14730 7050 14750
rect 7050 14730 7070 14750
rect 7070 14730 7075 14750
rect 7045 14725 7075 14730
rect 7125 14750 7155 14755
rect 7125 14730 7130 14750
rect 7130 14730 7150 14750
rect 7150 14730 7155 14750
rect 7125 14725 7155 14730
rect 7205 14750 7235 14755
rect 7205 14730 7210 14750
rect 7210 14730 7230 14750
rect 7230 14730 7235 14750
rect 7205 14725 7235 14730
rect 7285 14750 7315 14755
rect 7285 14730 7290 14750
rect 7290 14730 7310 14750
rect 7310 14730 7315 14750
rect 7285 14725 7315 14730
rect 7365 14750 7395 14755
rect 7365 14730 7370 14750
rect 7370 14730 7390 14750
rect 7390 14730 7395 14750
rect 7365 14725 7395 14730
rect 7445 14750 7475 14755
rect 7445 14730 7450 14750
rect 7450 14730 7470 14750
rect 7470 14730 7475 14750
rect 7445 14725 7475 14730
rect 7525 14750 7555 14755
rect 7525 14730 7530 14750
rect 7530 14730 7550 14750
rect 7550 14730 7555 14750
rect 7525 14725 7555 14730
rect 7605 14750 7635 14755
rect 7605 14730 7610 14750
rect 7610 14730 7630 14750
rect 7630 14730 7635 14750
rect 7605 14725 7635 14730
rect 7685 14750 7715 14755
rect 7685 14730 7690 14750
rect 7690 14730 7710 14750
rect 7710 14730 7715 14750
rect 7685 14725 7715 14730
rect 7765 14750 7795 14755
rect 7765 14730 7770 14750
rect 7770 14730 7790 14750
rect 7790 14730 7795 14750
rect 7765 14725 7795 14730
rect 7845 14750 7875 14755
rect 7845 14730 7850 14750
rect 7850 14730 7870 14750
rect 7870 14730 7875 14750
rect 7845 14725 7875 14730
rect 7925 14750 7955 14755
rect 7925 14730 7930 14750
rect 7930 14730 7950 14750
rect 7950 14730 7955 14750
rect 7925 14725 7955 14730
rect 8005 14750 8035 14755
rect 8005 14730 8010 14750
rect 8010 14730 8030 14750
rect 8030 14730 8035 14750
rect 8005 14725 8035 14730
rect 8085 14750 8115 14755
rect 8085 14730 8090 14750
rect 8090 14730 8110 14750
rect 8110 14730 8115 14750
rect 8085 14725 8115 14730
rect 8165 14750 8195 14755
rect 8165 14730 8170 14750
rect 8170 14730 8190 14750
rect 8190 14730 8195 14750
rect 8165 14725 8195 14730
rect 8245 14750 8275 14755
rect 8245 14730 8250 14750
rect 8250 14730 8270 14750
rect 8270 14730 8275 14750
rect 8245 14725 8275 14730
rect 8325 14750 8355 14755
rect 8325 14730 8330 14750
rect 8330 14730 8350 14750
rect 8350 14730 8355 14750
rect 8325 14725 8355 14730
rect 8405 14750 8435 14755
rect 8405 14730 8410 14750
rect 8410 14730 8430 14750
rect 8430 14730 8435 14750
rect 8405 14725 8435 14730
rect 8485 14750 8515 14755
rect 8485 14730 8490 14750
rect 8490 14730 8510 14750
rect 8510 14730 8515 14750
rect 8485 14725 8515 14730
rect 8565 14750 8595 14755
rect 8565 14730 8570 14750
rect 8570 14730 8590 14750
rect 8590 14730 8595 14750
rect 8565 14725 8595 14730
rect 8645 14750 8675 14755
rect 8645 14730 8650 14750
rect 8650 14730 8670 14750
rect 8670 14730 8675 14750
rect 8645 14725 8675 14730
rect 8725 14750 8755 14755
rect 8725 14730 8730 14750
rect 8730 14730 8750 14750
rect 8750 14730 8755 14750
rect 8725 14725 8755 14730
rect 8805 14750 8835 14755
rect 8805 14730 8810 14750
rect 8810 14730 8830 14750
rect 8830 14730 8835 14750
rect 8805 14725 8835 14730
rect 8885 14750 8915 14755
rect 8885 14730 8890 14750
rect 8890 14730 8910 14750
rect 8910 14730 8915 14750
rect 8885 14725 8915 14730
rect 8965 14750 8995 14755
rect 8965 14730 8970 14750
rect 8970 14730 8990 14750
rect 8990 14730 8995 14750
rect 8965 14725 8995 14730
rect 9045 14750 9075 14755
rect 9045 14730 9050 14750
rect 9050 14730 9070 14750
rect 9070 14730 9075 14750
rect 9045 14725 9075 14730
rect 9125 14750 9155 14755
rect 9125 14730 9130 14750
rect 9130 14730 9150 14750
rect 9150 14730 9155 14750
rect 9125 14725 9155 14730
rect 9205 14750 9235 14755
rect 9205 14730 9210 14750
rect 9210 14730 9230 14750
rect 9230 14730 9235 14750
rect 9205 14725 9235 14730
rect 9285 14750 9315 14755
rect 9285 14730 9290 14750
rect 9290 14730 9310 14750
rect 9310 14730 9315 14750
rect 9285 14725 9315 14730
rect 9365 14750 9395 14755
rect 9365 14730 9370 14750
rect 9370 14730 9390 14750
rect 9390 14730 9395 14750
rect 9365 14725 9395 14730
rect 9445 14750 9475 14755
rect 9445 14730 9450 14750
rect 9450 14730 9470 14750
rect 9470 14730 9475 14750
rect 9445 14725 9475 14730
rect 11565 14750 11595 14755
rect 11565 14730 11570 14750
rect 11570 14730 11590 14750
rect 11590 14730 11595 14750
rect 11565 14725 11595 14730
rect 11645 14750 11675 14755
rect 11645 14730 11650 14750
rect 11650 14730 11670 14750
rect 11670 14730 11675 14750
rect 11645 14725 11675 14730
rect 11725 14750 11755 14755
rect 11725 14730 11730 14750
rect 11730 14730 11750 14750
rect 11750 14730 11755 14750
rect 11725 14725 11755 14730
rect 11805 14750 11835 14755
rect 11805 14730 11810 14750
rect 11810 14730 11830 14750
rect 11830 14730 11835 14750
rect 11805 14725 11835 14730
rect 11885 14750 11915 14755
rect 11885 14730 11890 14750
rect 11890 14730 11910 14750
rect 11910 14730 11915 14750
rect 11885 14725 11915 14730
rect 11965 14750 11995 14755
rect 11965 14730 11970 14750
rect 11970 14730 11990 14750
rect 11990 14730 11995 14750
rect 11965 14725 11995 14730
rect 12045 14750 12075 14755
rect 12045 14730 12050 14750
rect 12050 14730 12070 14750
rect 12070 14730 12075 14750
rect 12045 14725 12075 14730
rect 12125 14750 12155 14755
rect 12125 14730 12130 14750
rect 12130 14730 12150 14750
rect 12150 14730 12155 14750
rect 12125 14725 12155 14730
rect 12205 14750 12235 14755
rect 12205 14730 12210 14750
rect 12210 14730 12230 14750
rect 12230 14730 12235 14750
rect 12205 14725 12235 14730
rect 12285 14750 12315 14755
rect 12285 14730 12290 14750
rect 12290 14730 12310 14750
rect 12310 14730 12315 14750
rect 12285 14725 12315 14730
rect 12365 14750 12395 14755
rect 12365 14730 12370 14750
rect 12370 14730 12390 14750
rect 12390 14730 12395 14750
rect 12365 14725 12395 14730
rect 12445 14750 12475 14755
rect 12445 14730 12450 14750
rect 12450 14730 12470 14750
rect 12470 14730 12475 14750
rect 12445 14725 12475 14730
rect 12525 14750 12555 14755
rect 12525 14730 12530 14750
rect 12530 14730 12550 14750
rect 12550 14730 12555 14750
rect 12525 14725 12555 14730
rect 12605 14750 12635 14755
rect 12605 14730 12610 14750
rect 12610 14730 12630 14750
rect 12630 14730 12635 14750
rect 12605 14725 12635 14730
rect 12685 14750 12715 14755
rect 12685 14730 12690 14750
rect 12690 14730 12710 14750
rect 12710 14730 12715 14750
rect 12685 14725 12715 14730
rect 12765 14750 12795 14755
rect 12765 14730 12770 14750
rect 12770 14730 12790 14750
rect 12790 14730 12795 14750
rect 12765 14725 12795 14730
rect 12845 14750 12875 14755
rect 12845 14730 12850 14750
rect 12850 14730 12870 14750
rect 12870 14730 12875 14750
rect 12845 14725 12875 14730
rect 12925 14750 12955 14755
rect 12925 14730 12930 14750
rect 12930 14730 12950 14750
rect 12950 14730 12955 14750
rect 12925 14725 12955 14730
rect 13005 14750 13035 14755
rect 13005 14730 13010 14750
rect 13010 14730 13030 14750
rect 13030 14730 13035 14750
rect 13005 14725 13035 14730
rect 13085 14750 13115 14755
rect 13085 14730 13090 14750
rect 13090 14730 13110 14750
rect 13110 14730 13115 14750
rect 13085 14725 13115 14730
rect 13165 14750 13195 14755
rect 13165 14730 13170 14750
rect 13170 14730 13190 14750
rect 13190 14730 13195 14750
rect 13165 14725 13195 14730
rect 13245 14750 13275 14755
rect 13245 14730 13250 14750
rect 13250 14730 13270 14750
rect 13270 14730 13275 14750
rect 13245 14725 13275 14730
rect 13325 14750 13355 14755
rect 13325 14730 13330 14750
rect 13330 14730 13350 14750
rect 13350 14730 13355 14750
rect 13325 14725 13355 14730
rect 13405 14750 13435 14755
rect 13405 14730 13410 14750
rect 13410 14730 13430 14750
rect 13430 14730 13435 14750
rect 13405 14725 13435 14730
rect 13485 14750 13515 14755
rect 13485 14730 13490 14750
rect 13490 14730 13510 14750
rect 13510 14730 13515 14750
rect 13485 14725 13515 14730
rect 13565 14750 13595 14755
rect 13565 14730 13570 14750
rect 13570 14730 13590 14750
rect 13590 14730 13595 14750
rect 13565 14725 13595 14730
rect 13645 14750 13675 14755
rect 13645 14730 13650 14750
rect 13650 14730 13670 14750
rect 13670 14730 13675 14750
rect 13645 14725 13675 14730
rect 13725 14750 13755 14755
rect 13725 14730 13730 14750
rect 13730 14730 13750 14750
rect 13750 14730 13755 14750
rect 13725 14725 13755 14730
rect 13805 14750 13835 14755
rect 13805 14730 13810 14750
rect 13810 14730 13830 14750
rect 13830 14730 13835 14750
rect 13805 14725 13835 14730
rect 13885 14750 13915 14755
rect 13885 14730 13890 14750
rect 13890 14730 13910 14750
rect 13910 14730 13915 14750
rect 13885 14725 13915 14730
rect 13965 14750 13995 14755
rect 13965 14730 13970 14750
rect 13970 14730 13990 14750
rect 13990 14730 13995 14750
rect 13965 14725 13995 14730
rect 14045 14750 14075 14755
rect 14045 14730 14050 14750
rect 14050 14730 14070 14750
rect 14070 14730 14075 14750
rect 14045 14725 14075 14730
rect 14125 14750 14155 14755
rect 14125 14730 14130 14750
rect 14130 14730 14150 14750
rect 14150 14730 14155 14750
rect 14125 14725 14155 14730
rect 14205 14750 14235 14755
rect 14205 14730 14210 14750
rect 14210 14730 14230 14750
rect 14230 14730 14235 14750
rect 14205 14725 14235 14730
rect 14285 14750 14315 14755
rect 14285 14730 14290 14750
rect 14290 14730 14310 14750
rect 14310 14730 14315 14750
rect 14285 14725 14315 14730
rect 14365 14750 14395 14755
rect 14365 14730 14370 14750
rect 14370 14730 14390 14750
rect 14390 14730 14395 14750
rect 14365 14725 14395 14730
rect 14445 14750 14475 14755
rect 14445 14730 14450 14750
rect 14450 14730 14470 14750
rect 14470 14730 14475 14750
rect 14445 14725 14475 14730
rect 14525 14750 14555 14755
rect 14525 14730 14530 14750
rect 14530 14730 14550 14750
rect 14550 14730 14555 14750
rect 14525 14725 14555 14730
rect 14605 14750 14635 14755
rect 14605 14730 14610 14750
rect 14610 14730 14630 14750
rect 14630 14730 14635 14750
rect 14605 14725 14635 14730
rect 14685 14750 14715 14755
rect 14685 14730 14690 14750
rect 14690 14730 14710 14750
rect 14710 14730 14715 14750
rect 14685 14725 14715 14730
rect 16765 14750 16795 14755
rect 16765 14730 16770 14750
rect 16770 14730 16790 14750
rect 16790 14730 16795 14750
rect 16765 14725 16795 14730
rect 16845 14750 16875 14755
rect 16845 14730 16850 14750
rect 16850 14730 16870 14750
rect 16870 14730 16875 14750
rect 16845 14725 16875 14730
rect 16925 14750 16955 14755
rect 16925 14730 16930 14750
rect 16930 14730 16950 14750
rect 16950 14730 16955 14750
rect 16925 14725 16955 14730
rect 17005 14750 17035 14755
rect 17005 14730 17010 14750
rect 17010 14730 17030 14750
rect 17030 14730 17035 14750
rect 17005 14725 17035 14730
rect 17085 14750 17115 14755
rect 17085 14730 17090 14750
rect 17090 14730 17110 14750
rect 17110 14730 17115 14750
rect 17085 14725 17115 14730
rect 17165 14750 17195 14755
rect 17165 14730 17170 14750
rect 17170 14730 17190 14750
rect 17190 14730 17195 14750
rect 17165 14725 17195 14730
rect 17245 14750 17275 14755
rect 17245 14730 17250 14750
rect 17250 14730 17270 14750
rect 17270 14730 17275 14750
rect 17245 14725 17275 14730
rect 17325 14750 17355 14755
rect 17325 14730 17330 14750
rect 17330 14730 17350 14750
rect 17350 14730 17355 14750
rect 17325 14725 17355 14730
rect 17405 14750 17435 14755
rect 17405 14730 17410 14750
rect 17410 14730 17430 14750
rect 17430 14730 17435 14750
rect 17405 14725 17435 14730
rect 17485 14750 17515 14755
rect 17485 14730 17490 14750
rect 17490 14730 17510 14750
rect 17510 14730 17515 14750
rect 17485 14725 17515 14730
rect 17565 14750 17595 14755
rect 17565 14730 17570 14750
rect 17570 14730 17590 14750
rect 17590 14730 17595 14750
rect 17565 14725 17595 14730
rect 17645 14750 17675 14755
rect 17645 14730 17650 14750
rect 17650 14730 17670 14750
rect 17670 14730 17675 14750
rect 17645 14725 17675 14730
rect 17725 14750 17755 14755
rect 17725 14730 17730 14750
rect 17730 14730 17750 14750
rect 17750 14730 17755 14750
rect 17725 14725 17755 14730
rect 17805 14750 17835 14755
rect 17805 14730 17810 14750
rect 17810 14730 17830 14750
rect 17830 14730 17835 14750
rect 17805 14725 17835 14730
rect 17885 14750 17915 14755
rect 17885 14730 17890 14750
rect 17890 14730 17910 14750
rect 17910 14730 17915 14750
rect 17885 14725 17915 14730
rect 17965 14750 17995 14755
rect 17965 14730 17970 14750
rect 17970 14730 17990 14750
rect 17990 14730 17995 14750
rect 17965 14725 17995 14730
rect 18045 14750 18075 14755
rect 18045 14730 18050 14750
rect 18050 14730 18070 14750
rect 18070 14730 18075 14750
rect 18045 14725 18075 14730
rect 18125 14750 18155 14755
rect 18125 14730 18130 14750
rect 18130 14730 18150 14750
rect 18150 14730 18155 14750
rect 18125 14725 18155 14730
rect 18205 14750 18235 14755
rect 18205 14730 18210 14750
rect 18210 14730 18230 14750
rect 18230 14730 18235 14750
rect 18205 14725 18235 14730
rect 18285 14750 18315 14755
rect 18285 14730 18290 14750
rect 18290 14730 18310 14750
rect 18310 14730 18315 14750
rect 18285 14725 18315 14730
rect 18365 14750 18395 14755
rect 18365 14730 18370 14750
rect 18370 14730 18390 14750
rect 18390 14730 18395 14750
rect 18365 14725 18395 14730
rect 18445 14750 18475 14755
rect 18445 14730 18450 14750
rect 18450 14730 18470 14750
rect 18470 14730 18475 14750
rect 18445 14725 18475 14730
rect 18525 14750 18555 14755
rect 18525 14730 18530 14750
rect 18530 14730 18550 14750
rect 18550 14730 18555 14750
rect 18525 14725 18555 14730
rect 18605 14750 18635 14755
rect 18605 14730 18610 14750
rect 18610 14730 18630 14750
rect 18630 14730 18635 14750
rect 18605 14725 18635 14730
rect 18685 14750 18715 14755
rect 18685 14730 18690 14750
rect 18690 14730 18710 14750
rect 18710 14730 18715 14750
rect 18685 14725 18715 14730
rect 18765 14750 18795 14755
rect 18765 14730 18770 14750
rect 18770 14730 18790 14750
rect 18790 14730 18795 14750
rect 18765 14725 18795 14730
rect 18845 14750 18875 14755
rect 18845 14730 18850 14750
rect 18850 14730 18870 14750
rect 18870 14730 18875 14750
rect 18845 14725 18875 14730
rect 18925 14750 18955 14755
rect 18925 14730 18930 14750
rect 18930 14730 18950 14750
rect 18950 14730 18955 14750
rect 18925 14725 18955 14730
rect 19005 14750 19035 14755
rect 19005 14730 19010 14750
rect 19010 14730 19030 14750
rect 19030 14730 19035 14750
rect 19005 14725 19035 14730
rect 19085 14750 19115 14755
rect 19085 14730 19090 14750
rect 19090 14730 19110 14750
rect 19110 14730 19115 14750
rect 19085 14725 19115 14730
rect 19165 14750 19195 14755
rect 19165 14730 19170 14750
rect 19170 14730 19190 14750
rect 19190 14730 19195 14750
rect 19165 14725 19195 14730
rect 19245 14750 19275 14755
rect 19245 14730 19250 14750
rect 19250 14730 19270 14750
rect 19270 14730 19275 14750
rect 19245 14725 19275 14730
rect 19325 14750 19355 14755
rect 19325 14730 19330 14750
rect 19330 14730 19350 14750
rect 19350 14730 19355 14750
rect 19325 14725 19355 14730
rect 19405 14750 19435 14755
rect 19405 14730 19410 14750
rect 19410 14730 19430 14750
rect 19430 14730 19435 14750
rect 19405 14725 19435 14730
rect 19485 14750 19515 14755
rect 19485 14730 19490 14750
rect 19490 14730 19510 14750
rect 19510 14730 19515 14750
rect 19485 14725 19515 14730
rect 19565 14750 19595 14755
rect 19565 14730 19570 14750
rect 19570 14730 19590 14750
rect 19590 14730 19595 14750
rect 19565 14725 19595 14730
rect 19645 14750 19675 14755
rect 19645 14730 19650 14750
rect 19650 14730 19670 14750
rect 19670 14730 19675 14750
rect 19645 14725 19675 14730
rect 19725 14750 19755 14755
rect 19725 14730 19730 14750
rect 19730 14730 19750 14750
rect 19750 14730 19755 14750
rect 19725 14725 19755 14730
rect 19805 14750 19835 14755
rect 19805 14730 19810 14750
rect 19810 14730 19830 14750
rect 19830 14730 19835 14750
rect 19805 14725 19835 14730
rect 19885 14750 19915 14755
rect 19885 14730 19890 14750
rect 19890 14730 19910 14750
rect 19910 14730 19915 14750
rect 19885 14725 19915 14730
rect 19965 14750 19995 14755
rect 19965 14730 19970 14750
rect 19970 14730 19990 14750
rect 19990 14730 19995 14750
rect 19965 14725 19995 14730
rect 20045 14750 20075 14755
rect 20045 14730 20050 14750
rect 20050 14730 20070 14750
rect 20070 14730 20075 14750
rect 20045 14725 20075 14730
rect 20125 14750 20155 14755
rect 20125 14730 20130 14750
rect 20130 14730 20150 14750
rect 20150 14730 20155 14750
rect 20125 14725 20155 14730
rect 20205 14750 20235 14755
rect 20205 14730 20210 14750
rect 20210 14730 20230 14750
rect 20230 14730 20235 14750
rect 20205 14725 20235 14730
rect 20285 14750 20315 14755
rect 20285 14730 20290 14750
rect 20290 14730 20310 14750
rect 20310 14730 20315 14750
rect 20285 14725 20315 14730
rect 20365 14750 20395 14755
rect 20365 14730 20370 14750
rect 20370 14730 20390 14750
rect 20390 14730 20395 14750
rect 20365 14725 20395 14730
rect 20445 14750 20475 14755
rect 20445 14730 20450 14750
rect 20450 14730 20470 14750
rect 20470 14730 20475 14750
rect 20445 14725 20475 14730
rect 20525 14750 20555 14755
rect 20525 14730 20530 14750
rect 20530 14730 20550 14750
rect 20550 14730 20555 14750
rect 20525 14725 20555 14730
rect 20605 14750 20635 14755
rect 20605 14730 20610 14750
rect 20610 14730 20630 14750
rect 20630 14730 20635 14750
rect 20605 14725 20635 14730
rect 20685 14750 20715 14755
rect 20685 14730 20690 14750
rect 20690 14730 20710 14750
rect 20710 14730 20715 14750
rect 20685 14725 20715 14730
rect 20765 14750 20795 14755
rect 20765 14730 20770 14750
rect 20770 14730 20790 14750
rect 20790 14730 20795 14750
rect 20765 14725 20795 14730
rect 20845 14750 20875 14755
rect 20845 14730 20850 14750
rect 20850 14730 20870 14750
rect 20870 14730 20875 14750
rect 20845 14725 20875 14730
rect 20925 14750 20955 14755
rect 20925 14730 20930 14750
rect 20930 14730 20950 14750
rect 20950 14730 20955 14750
rect 20925 14725 20955 14730
<< metal2 >>
rect 0 18675 20960 18680
rect 0 18645 5 18675
rect 35 18645 85 18675
rect 115 18645 165 18675
rect 195 18645 245 18675
rect 275 18645 325 18675
rect 355 18645 405 18675
rect 435 18645 485 18675
rect 515 18645 565 18675
rect 595 18645 645 18675
rect 675 18645 725 18675
rect 755 18645 805 18675
rect 835 18645 885 18675
rect 915 18645 965 18675
rect 995 18645 1045 18675
rect 1075 18645 1125 18675
rect 1155 18645 1205 18675
rect 1235 18645 1285 18675
rect 1315 18645 1365 18675
rect 1395 18645 1445 18675
rect 1475 18645 1525 18675
rect 1555 18645 1605 18675
rect 1635 18645 1685 18675
rect 1715 18645 1765 18675
rect 1795 18645 1845 18675
rect 1875 18645 1925 18675
rect 1955 18645 2005 18675
rect 2035 18645 2085 18675
rect 2115 18645 2165 18675
rect 2195 18645 2245 18675
rect 2275 18645 2325 18675
rect 2355 18645 2405 18675
rect 2435 18645 2485 18675
rect 2515 18645 2565 18675
rect 2595 18645 2645 18675
rect 2675 18645 2725 18675
rect 2755 18645 2805 18675
rect 2835 18645 2885 18675
rect 2915 18645 2965 18675
rect 2995 18645 3045 18675
rect 3075 18645 3125 18675
rect 3155 18645 3205 18675
rect 3235 18645 3285 18675
rect 3315 18645 3365 18675
rect 3395 18645 3445 18675
rect 3475 18645 3525 18675
rect 3555 18645 3605 18675
rect 3635 18645 3685 18675
rect 3715 18645 3765 18675
rect 3795 18645 3845 18675
rect 3875 18645 3925 18675
rect 3955 18645 4005 18675
rect 4035 18645 4085 18675
rect 4115 18645 4165 18675
rect 4195 18645 4245 18675
rect 4275 18645 4405 18675
rect 4435 18645 6245 18675
rect 6275 18645 6325 18675
rect 6355 18645 6405 18675
rect 6435 18645 6485 18675
rect 6515 18645 6565 18675
rect 6595 18645 6645 18675
rect 6675 18645 6725 18675
rect 6755 18645 6805 18675
rect 6835 18645 6885 18675
rect 6915 18645 6965 18675
rect 6995 18645 7045 18675
rect 7075 18645 7125 18675
rect 7155 18645 7205 18675
rect 7235 18645 7285 18675
rect 7315 18645 7365 18675
rect 7395 18645 7445 18675
rect 7475 18645 7525 18675
rect 7555 18645 7605 18675
rect 7635 18645 7685 18675
rect 7715 18645 7765 18675
rect 7795 18645 7845 18675
rect 7875 18645 7925 18675
rect 7955 18645 8005 18675
rect 8035 18645 8085 18675
rect 8115 18645 8165 18675
rect 8195 18645 8245 18675
rect 8275 18645 8325 18675
rect 8355 18645 8405 18675
rect 8435 18645 8485 18675
rect 8515 18645 8565 18675
rect 8595 18645 8645 18675
rect 8675 18645 8725 18675
rect 8755 18645 8805 18675
rect 8835 18645 8885 18675
rect 8915 18645 8965 18675
rect 8995 18645 9045 18675
rect 9075 18645 9125 18675
rect 9155 18645 9205 18675
rect 9235 18645 9285 18675
rect 9315 18645 9365 18675
rect 9395 18645 9445 18675
rect 9475 18645 11285 18675
rect 11315 18645 11445 18675
rect 11475 18645 11565 18675
rect 11595 18645 11645 18675
rect 11675 18645 11725 18675
rect 11755 18645 11805 18675
rect 11835 18645 11885 18675
rect 11915 18645 11965 18675
rect 11995 18645 12045 18675
rect 12075 18645 12125 18675
rect 12155 18645 12205 18675
rect 12235 18645 12285 18675
rect 12315 18645 12365 18675
rect 12395 18645 12445 18675
rect 12475 18645 12525 18675
rect 12555 18645 12605 18675
rect 12635 18645 12685 18675
rect 12715 18645 12765 18675
rect 12795 18645 12845 18675
rect 12875 18645 12925 18675
rect 12955 18645 13005 18675
rect 13035 18645 13085 18675
rect 13115 18645 13165 18675
rect 13195 18645 13245 18675
rect 13275 18645 13325 18675
rect 13355 18645 13405 18675
rect 13435 18645 13485 18675
rect 13515 18645 13565 18675
rect 13595 18645 13645 18675
rect 13675 18645 13725 18675
rect 13755 18645 13805 18675
rect 13835 18645 13885 18675
rect 13915 18645 13965 18675
rect 13995 18645 14045 18675
rect 14075 18645 14125 18675
rect 14155 18645 14205 18675
rect 14235 18645 14285 18675
rect 14315 18645 14365 18675
rect 14395 18645 14445 18675
rect 14475 18645 14525 18675
rect 14555 18645 14605 18675
rect 14635 18645 14685 18675
rect 14715 18645 16525 18675
rect 16555 18645 16685 18675
rect 16715 18645 16765 18675
rect 16795 18645 16845 18675
rect 16875 18645 16925 18675
rect 16955 18645 17005 18675
rect 17035 18645 17085 18675
rect 17115 18645 17165 18675
rect 17195 18645 17245 18675
rect 17275 18645 17325 18675
rect 17355 18645 17405 18675
rect 17435 18645 17485 18675
rect 17515 18645 17565 18675
rect 17595 18645 17645 18675
rect 17675 18645 17725 18675
rect 17755 18645 17805 18675
rect 17835 18645 17885 18675
rect 17915 18645 17965 18675
rect 17995 18645 18045 18675
rect 18075 18645 18125 18675
rect 18155 18645 18205 18675
rect 18235 18645 18285 18675
rect 18315 18645 18365 18675
rect 18395 18645 18445 18675
rect 18475 18645 18525 18675
rect 18555 18645 18605 18675
rect 18635 18645 18685 18675
rect 18715 18645 18765 18675
rect 18795 18645 18845 18675
rect 18875 18645 18925 18675
rect 18955 18645 19005 18675
rect 19035 18645 19085 18675
rect 19115 18645 19165 18675
rect 19195 18645 19245 18675
rect 19275 18645 19325 18675
rect 19355 18645 19405 18675
rect 19435 18645 19485 18675
rect 19515 18645 19565 18675
rect 19595 18645 19645 18675
rect 19675 18645 19725 18675
rect 19755 18645 19805 18675
rect 19835 18645 19885 18675
rect 19915 18645 19965 18675
rect 19995 18645 20045 18675
rect 20075 18645 20125 18675
rect 20155 18645 20205 18675
rect 20235 18645 20285 18675
rect 20315 18645 20365 18675
rect 20395 18645 20445 18675
rect 20475 18645 20525 18675
rect 20555 18645 20605 18675
rect 20635 18645 20685 18675
rect 20715 18645 20765 18675
rect 20795 18645 20845 18675
rect 20875 18645 20925 18675
rect 20955 18645 20960 18675
rect 0 18640 20960 18645
rect 0 18595 20960 18600
rect 0 18565 4325 18595
rect 4355 18565 11365 18595
rect 11395 18565 16605 18595
rect 16635 18565 20960 18595
rect 0 18560 20960 18565
rect 0 18515 20960 18520
rect 0 18485 5 18515
rect 35 18485 85 18515
rect 115 18485 165 18515
rect 195 18485 245 18515
rect 275 18485 325 18515
rect 355 18485 405 18515
rect 435 18485 485 18515
rect 515 18485 565 18515
rect 595 18485 645 18515
rect 675 18485 725 18515
rect 755 18485 805 18515
rect 835 18485 885 18515
rect 915 18485 965 18515
rect 995 18485 1045 18515
rect 1075 18485 1125 18515
rect 1155 18485 1205 18515
rect 1235 18485 1285 18515
rect 1315 18485 1365 18515
rect 1395 18485 1445 18515
rect 1475 18485 1525 18515
rect 1555 18485 1605 18515
rect 1635 18485 1685 18515
rect 1715 18485 1765 18515
rect 1795 18485 1845 18515
rect 1875 18485 1925 18515
rect 1955 18485 2005 18515
rect 2035 18485 2085 18515
rect 2115 18485 2165 18515
rect 2195 18485 2245 18515
rect 2275 18485 2325 18515
rect 2355 18485 2405 18515
rect 2435 18485 2485 18515
rect 2515 18485 2565 18515
rect 2595 18485 2645 18515
rect 2675 18485 2725 18515
rect 2755 18485 2805 18515
rect 2835 18485 2885 18515
rect 2915 18485 2965 18515
rect 2995 18485 3045 18515
rect 3075 18485 3125 18515
rect 3155 18485 3205 18515
rect 3235 18485 3285 18515
rect 3315 18485 3365 18515
rect 3395 18485 3445 18515
rect 3475 18485 3525 18515
rect 3555 18485 3605 18515
rect 3635 18485 3685 18515
rect 3715 18485 3765 18515
rect 3795 18485 3845 18515
rect 3875 18485 3925 18515
rect 3955 18485 4005 18515
rect 4035 18485 4085 18515
rect 4115 18485 4165 18515
rect 4195 18485 4245 18515
rect 4275 18485 4405 18515
rect 4435 18485 6245 18515
rect 6275 18485 6325 18515
rect 6355 18485 6405 18515
rect 6435 18485 6485 18515
rect 6515 18485 6565 18515
rect 6595 18485 6645 18515
rect 6675 18485 6725 18515
rect 6755 18485 6805 18515
rect 6835 18485 6885 18515
rect 6915 18485 6965 18515
rect 6995 18485 7045 18515
rect 7075 18485 7125 18515
rect 7155 18485 7205 18515
rect 7235 18485 7285 18515
rect 7315 18485 7365 18515
rect 7395 18485 7445 18515
rect 7475 18485 7525 18515
rect 7555 18485 7605 18515
rect 7635 18485 7685 18515
rect 7715 18485 7765 18515
rect 7795 18485 7845 18515
rect 7875 18485 7925 18515
rect 7955 18485 8005 18515
rect 8035 18485 8085 18515
rect 8115 18485 8165 18515
rect 8195 18485 8245 18515
rect 8275 18485 8325 18515
rect 8355 18485 8405 18515
rect 8435 18485 8485 18515
rect 8515 18485 8565 18515
rect 8595 18485 8645 18515
rect 8675 18485 8725 18515
rect 8755 18485 8805 18515
rect 8835 18485 8885 18515
rect 8915 18485 8965 18515
rect 8995 18485 9045 18515
rect 9075 18485 9125 18515
rect 9155 18485 9205 18515
rect 9235 18485 9285 18515
rect 9315 18485 9365 18515
rect 9395 18485 9445 18515
rect 9475 18485 11285 18515
rect 11315 18485 11445 18515
rect 11475 18485 11565 18515
rect 11595 18485 11645 18515
rect 11675 18485 11725 18515
rect 11755 18485 11805 18515
rect 11835 18485 11885 18515
rect 11915 18485 11965 18515
rect 11995 18485 12045 18515
rect 12075 18485 12125 18515
rect 12155 18485 12205 18515
rect 12235 18485 12285 18515
rect 12315 18485 12365 18515
rect 12395 18485 12445 18515
rect 12475 18485 12525 18515
rect 12555 18485 12605 18515
rect 12635 18485 12685 18515
rect 12715 18485 12765 18515
rect 12795 18485 12845 18515
rect 12875 18485 12925 18515
rect 12955 18485 13005 18515
rect 13035 18485 13085 18515
rect 13115 18485 13165 18515
rect 13195 18485 13245 18515
rect 13275 18485 13325 18515
rect 13355 18485 13405 18515
rect 13435 18485 13485 18515
rect 13515 18485 13565 18515
rect 13595 18485 13645 18515
rect 13675 18485 13725 18515
rect 13755 18485 13805 18515
rect 13835 18485 13885 18515
rect 13915 18485 13965 18515
rect 13995 18485 14045 18515
rect 14075 18485 14125 18515
rect 14155 18485 14205 18515
rect 14235 18485 14285 18515
rect 14315 18485 14365 18515
rect 14395 18485 14445 18515
rect 14475 18485 14525 18515
rect 14555 18485 14605 18515
rect 14635 18485 14685 18515
rect 14715 18485 16525 18515
rect 16555 18485 16685 18515
rect 16715 18485 16765 18515
rect 16795 18485 16845 18515
rect 16875 18485 16925 18515
rect 16955 18485 17005 18515
rect 17035 18485 17085 18515
rect 17115 18485 17165 18515
rect 17195 18485 17245 18515
rect 17275 18485 17325 18515
rect 17355 18485 17405 18515
rect 17435 18485 17485 18515
rect 17515 18485 17565 18515
rect 17595 18485 17645 18515
rect 17675 18485 17725 18515
rect 17755 18485 17805 18515
rect 17835 18485 17885 18515
rect 17915 18485 17965 18515
rect 17995 18485 18045 18515
rect 18075 18485 18125 18515
rect 18155 18485 18205 18515
rect 18235 18485 18285 18515
rect 18315 18485 18365 18515
rect 18395 18485 18445 18515
rect 18475 18485 18525 18515
rect 18555 18485 18605 18515
rect 18635 18485 18685 18515
rect 18715 18485 18765 18515
rect 18795 18485 18845 18515
rect 18875 18485 18925 18515
rect 18955 18485 19005 18515
rect 19035 18485 19085 18515
rect 19115 18485 19165 18515
rect 19195 18485 19245 18515
rect 19275 18485 19325 18515
rect 19355 18485 19405 18515
rect 19435 18485 19485 18515
rect 19515 18485 19565 18515
rect 19595 18485 19645 18515
rect 19675 18485 19725 18515
rect 19755 18485 19805 18515
rect 19835 18485 19885 18515
rect 19915 18485 19965 18515
rect 19995 18485 20045 18515
rect 20075 18485 20125 18515
rect 20155 18485 20205 18515
rect 20235 18485 20285 18515
rect 20315 18485 20365 18515
rect 20395 18485 20445 18515
rect 20475 18485 20525 18515
rect 20555 18485 20605 18515
rect 20635 18485 20685 18515
rect 20715 18485 20765 18515
rect 20795 18485 20845 18515
rect 20875 18485 20925 18515
rect 20955 18485 20960 18515
rect 0 18480 20960 18485
rect 0 18435 20960 18440
rect 0 18405 5 18435
rect 35 18405 85 18435
rect 115 18405 165 18435
rect 195 18405 245 18435
rect 275 18405 325 18435
rect 355 18405 405 18435
rect 435 18405 485 18435
rect 515 18405 565 18435
rect 595 18405 645 18435
rect 675 18405 725 18435
rect 755 18405 805 18435
rect 835 18405 885 18435
rect 915 18405 965 18435
rect 995 18405 1045 18435
rect 1075 18405 1125 18435
rect 1155 18405 1205 18435
rect 1235 18405 1285 18435
rect 1315 18405 1365 18435
rect 1395 18405 1445 18435
rect 1475 18405 1525 18435
rect 1555 18405 1605 18435
rect 1635 18405 1685 18435
rect 1715 18405 1765 18435
rect 1795 18405 1845 18435
rect 1875 18405 1925 18435
rect 1955 18405 2005 18435
rect 2035 18405 2085 18435
rect 2115 18405 2165 18435
rect 2195 18405 2245 18435
rect 2275 18405 2325 18435
rect 2355 18405 2405 18435
rect 2435 18405 2485 18435
rect 2515 18405 2565 18435
rect 2595 18405 2645 18435
rect 2675 18405 2725 18435
rect 2755 18405 2805 18435
rect 2835 18405 2885 18435
rect 2915 18405 2965 18435
rect 2995 18405 3045 18435
rect 3075 18405 3125 18435
rect 3155 18405 3205 18435
rect 3235 18405 3285 18435
rect 3315 18405 3365 18435
rect 3395 18405 3445 18435
rect 3475 18405 3525 18435
rect 3555 18405 3605 18435
rect 3635 18405 3685 18435
rect 3715 18405 3765 18435
rect 3795 18405 3845 18435
rect 3875 18405 3925 18435
rect 3955 18405 4005 18435
rect 4035 18405 4085 18435
rect 4115 18405 4165 18435
rect 4195 18405 4485 18435
rect 4515 18405 4645 18435
rect 4675 18405 6245 18435
rect 6275 18405 6325 18435
rect 6355 18405 6405 18435
rect 6435 18405 6485 18435
rect 6515 18405 6565 18435
rect 6595 18405 6645 18435
rect 6675 18405 6725 18435
rect 6755 18405 6805 18435
rect 6835 18405 6885 18435
rect 6915 18405 6965 18435
rect 6995 18405 7045 18435
rect 7075 18405 7125 18435
rect 7155 18405 7205 18435
rect 7235 18405 7285 18435
rect 7315 18405 7365 18435
rect 7395 18405 7445 18435
rect 7475 18405 7525 18435
rect 7555 18405 7605 18435
rect 7635 18405 7685 18435
rect 7715 18405 7765 18435
rect 7795 18405 7845 18435
rect 7875 18405 7925 18435
rect 7955 18405 8005 18435
rect 8035 18405 8085 18435
rect 8115 18405 8165 18435
rect 8195 18405 8245 18435
rect 8275 18405 8325 18435
rect 8355 18405 8405 18435
rect 8435 18405 8485 18435
rect 8515 18405 8565 18435
rect 8595 18405 8645 18435
rect 8675 18405 8725 18435
rect 8755 18405 8805 18435
rect 8835 18405 8885 18435
rect 8915 18405 8965 18435
rect 8995 18405 9045 18435
rect 9075 18405 9125 18435
rect 9155 18405 9205 18435
rect 9235 18405 9285 18435
rect 9315 18405 9365 18435
rect 9395 18405 9445 18435
rect 9475 18405 11045 18435
rect 11075 18405 11205 18435
rect 11235 18405 11565 18435
rect 11595 18405 11645 18435
rect 11675 18405 11725 18435
rect 11755 18405 11805 18435
rect 11835 18405 11885 18435
rect 11915 18405 11965 18435
rect 11995 18405 12045 18435
rect 12075 18405 12125 18435
rect 12155 18405 12205 18435
rect 12235 18405 12285 18435
rect 12315 18405 12365 18435
rect 12395 18405 12445 18435
rect 12475 18405 12525 18435
rect 12555 18405 12605 18435
rect 12635 18405 12685 18435
rect 12715 18405 12765 18435
rect 12795 18405 12845 18435
rect 12875 18405 12925 18435
rect 12955 18405 13005 18435
rect 13035 18405 13085 18435
rect 13115 18405 13165 18435
rect 13195 18405 13245 18435
rect 13275 18405 13325 18435
rect 13355 18405 13405 18435
rect 13435 18405 13485 18435
rect 13515 18405 13565 18435
rect 13595 18405 13645 18435
rect 13675 18405 13725 18435
rect 13755 18405 13805 18435
rect 13835 18405 13885 18435
rect 13915 18405 13965 18435
rect 13995 18405 14045 18435
rect 14075 18405 14125 18435
rect 14155 18405 14205 18435
rect 14235 18405 14285 18435
rect 14315 18405 14365 18435
rect 14395 18405 14445 18435
rect 14475 18405 14525 18435
rect 14555 18405 14605 18435
rect 14635 18405 14685 18435
rect 14715 18405 16285 18435
rect 16315 18405 16445 18435
rect 16475 18405 16765 18435
rect 16795 18405 16845 18435
rect 16875 18405 16925 18435
rect 16955 18405 17005 18435
rect 17035 18405 17085 18435
rect 17115 18405 17165 18435
rect 17195 18405 17245 18435
rect 17275 18405 17325 18435
rect 17355 18405 17405 18435
rect 17435 18405 17485 18435
rect 17515 18405 17565 18435
rect 17595 18405 17645 18435
rect 17675 18405 17725 18435
rect 17755 18405 17805 18435
rect 17835 18405 17885 18435
rect 17915 18405 17965 18435
rect 17995 18405 18045 18435
rect 18075 18405 18125 18435
rect 18155 18405 18205 18435
rect 18235 18405 18285 18435
rect 18315 18405 18365 18435
rect 18395 18405 18445 18435
rect 18475 18405 18525 18435
rect 18555 18405 18605 18435
rect 18635 18405 18685 18435
rect 18715 18405 18765 18435
rect 18795 18405 18845 18435
rect 18875 18405 18925 18435
rect 18955 18405 19005 18435
rect 19035 18405 19085 18435
rect 19115 18405 19165 18435
rect 19195 18405 19245 18435
rect 19275 18405 19325 18435
rect 19355 18405 19405 18435
rect 19435 18405 19485 18435
rect 19515 18405 19565 18435
rect 19595 18405 19645 18435
rect 19675 18405 19725 18435
rect 19755 18405 19805 18435
rect 19835 18405 19885 18435
rect 19915 18405 19965 18435
rect 19995 18405 20045 18435
rect 20075 18405 20125 18435
rect 20155 18405 20205 18435
rect 20235 18405 20285 18435
rect 20315 18405 20365 18435
rect 20395 18405 20445 18435
rect 20475 18405 20525 18435
rect 20555 18405 20605 18435
rect 20635 18405 20685 18435
rect 20715 18405 20765 18435
rect 20795 18405 20845 18435
rect 20875 18405 20925 18435
rect 20955 18405 20960 18435
rect 0 18400 20960 18405
rect 0 18355 20960 18360
rect 0 18325 4565 18355
rect 4595 18325 11125 18355
rect 11155 18325 16365 18355
rect 16395 18325 20960 18355
rect 0 18320 20960 18325
rect 0 18275 20960 18280
rect 0 18245 5 18275
rect 35 18245 85 18275
rect 115 18245 165 18275
rect 195 18245 245 18275
rect 275 18245 325 18275
rect 355 18245 405 18275
rect 435 18245 485 18275
rect 515 18245 565 18275
rect 595 18245 645 18275
rect 675 18245 725 18275
rect 755 18245 805 18275
rect 835 18245 885 18275
rect 915 18245 965 18275
rect 995 18245 1045 18275
rect 1075 18245 1125 18275
rect 1155 18245 1205 18275
rect 1235 18245 1285 18275
rect 1315 18245 1365 18275
rect 1395 18245 1445 18275
rect 1475 18245 1525 18275
rect 1555 18245 1605 18275
rect 1635 18245 1685 18275
rect 1715 18245 1765 18275
rect 1795 18245 1845 18275
rect 1875 18245 1925 18275
rect 1955 18245 2005 18275
rect 2035 18245 2085 18275
rect 2115 18245 2165 18275
rect 2195 18245 2245 18275
rect 2275 18245 2325 18275
rect 2355 18245 2405 18275
rect 2435 18245 2485 18275
rect 2515 18245 2565 18275
rect 2595 18245 2645 18275
rect 2675 18245 2725 18275
rect 2755 18245 2805 18275
rect 2835 18245 2885 18275
rect 2915 18245 2965 18275
rect 2995 18245 3045 18275
rect 3075 18245 3125 18275
rect 3155 18245 3205 18275
rect 3235 18245 3285 18275
rect 3315 18245 3365 18275
rect 3395 18245 3445 18275
rect 3475 18245 3525 18275
rect 3555 18245 3605 18275
rect 3635 18245 3685 18275
rect 3715 18245 3765 18275
rect 3795 18245 3845 18275
rect 3875 18245 3925 18275
rect 3955 18245 4005 18275
rect 4035 18245 4085 18275
rect 4115 18245 4165 18275
rect 4195 18245 4485 18275
rect 4515 18245 4645 18275
rect 4675 18245 6245 18275
rect 6275 18245 6325 18275
rect 6355 18245 6405 18275
rect 6435 18245 6485 18275
rect 6515 18245 6565 18275
rect 6595 18245 6645 18275
rect 6675 18245 6725 18275
rect 6755 18245 6805 18275
rect 6835 18245 6885 18275
rect 6915 18245 6965 18275
rect 6995 18245 7045 18275
rect 7075 18245 7125 18275
rect 7155 18245 7205 18275
rect 7235 18245 7285 18275
rect 7315 18245 7365 18275
rect 7395 18245 7445 18275
rect 7475 18245 7525 18275
rect 7555 18245 7605 18275
rect 7635 18245 7685 18275
rect 7715 18245 7765 18275
rect 7795 18245 7845 18275
rect 7875 18245 7925 18275
rect 7955 18245 8005 18275
rect 8035 18245 8085 18275
rect 8115 18245 8165 18275
rect 8195 18245 8245 18275
rect 8275 18245 8325 18275
rect 8355 18245 8405 18275
rect 8435 18245 8485 18275
rect 8515 18245 8565 18275
rect 8595 18245 8645 18275
rect 8675 18245 8725 18275
rect 8755 18245 8805 18275
rect 8835 18245 8885 18275
rect 8915 18245 8965 18275
rect 8995 18245 9045 18275
rect 9075 18245 9125 18275
rect 9155 18245 9205 18275
rect 9235 18245 9285 18275
rect 9315 18245 9365 18275
rect 9395 18245 9445 18275
rect 9475 18245 11045 18275
rect 11075 18245 11205 18275
rect 11235 18245 11565 18275
rect 11595 18245 11645 18275
rect 11675 18245 11725 18275
rect 11755 18245 11805 18275
rect 11835 18245 11885 18275
rect 11915 18245 11965 18275
rect 11995 18245 12045 18275
rect 12075 18245 12125 18275
rect 12155 18245 12205 18275
rect 12235 18245 12285 18275
rect 12315 18245 12365 18275
rect 12395 18245 12445 18275
rect 12475 18245 12525 18275
rect 12555 18245 12605 18275
rect 12635 18245 12685 18275
rect 12715 18245 12765 18275
rect 12795 18245 12845 18275
rect 12875 18245 12925 18275
rect 12955 18245 13005 18275
rect 13035 18245 13085 18275
rect 13115 18245 13165 18275
rect 13195 18245 13245 18275
rect 13275 18245 13325 18275
rect 13355 18245 13405 18275
rect 13435 18245 13485 18275
rect 13515 18245 13565 18275
rect 13595 18245 13645 18275
rect 13675 18245 13725 18275
rect 13755 18245 13805 18275
rect 13835 18245 13885 18275
rect 13915 18245 13965 18275
rect 13995 18245 14045 18275
rect 14075 18245 14125 18275
rect 14155 18245 14205 18275
rect 14235 18245 14285 18275
rect 14315 18245 14365 18275
rect 14395 18245 14445 18275
rect 14475 18245 14525 18275
rect 14555 18245 14605 18275
rect 14635 18245 14685 18275
rect 14715 18245 16285 18275
rect 16315 18245 16445 18275
rect 16475 18245 16765 18275
rect 16795 18245 16845 18275
rect 16875 18245 16925 18275
rect 16955 18245 17005 18275
rect 17035 18245 17085 18275
rect 17115 18245 17165 18275
rect 17195 18245 17245 18275
rect 17275 18245 17325 18275
rect 17355 18245 17405 18275
rect 17435 18245 17485 18275
rect 17515 18245 17565 18275
rect 17595 18245 17645 18275
rect 17675 18245 17725 18275
rect 17755 18245 17805 18275
rect 17835 18245 17885 18275
rect 17915 18245 17965 18275
rect 17995 18245 18045 18275
rect 18075 18245 18125 18275
rect 18155 18245 18205 18275
rect 18235 18245 18285 18275
rect 18315 18245 18365 18275
rect 18395 18245 18445 18275
rect 18475 18245 18525 18275
rect 18555 18245 18605 18275
rect 18635 18245 18685 18275
rect 18715 18245 18765 18275
rect 18795 18245 18845 18275
rect 18875 18245 18925 18275
rect 18955 18245 19005 18275
rect 19035 18245 19085 18275
rect 19115 18245 19165 18275
rect 19195 18245 19245 18275
rect 19275 18245 19325 18275
rect 19355 18245 19405 18275
rect 19435 18245 19485 18275
rect 19515 18245 19565 18275
rect 19595 18245 19645 18275
rect 19675 18245 19725 18275
rect 19755 18245 19805 18275
rect 19835 18245 19885 18275
rect 19915 18245 19965 18275
rect 19995 18245 20045 18275
rect 20075 18245 20125 18275
rect 20155 18245 20205 18275
rect 20235 18245 20285 18275
rect 20315 18245 20365 18275
rect 20395 18245 20445 18275
rect 20475 18245 20525 18275
rect 20555 18245 20605 18275
rect 20635 18245 20685 18275
rect 20715 18245 20765 18275
rect 20795 18245 20845 18275
rect 20875 18245 20925 18275
rect 20955 18245 20960 18275
rect 0 18240 20960 18245
rect 0 18195 20960 18200
rect 0 18165 5 18195
rect 35 18165 85 18195
rect 115 18165 165 18195
rect 195 18165 245 18195
rect 275 18165 325 18195
rect 355 18165 405 18195
rect 435 18165 485 18195
rect 515 18165 565 18195
rect 595 18165 645 18195
rect 675 18165 725 18195
rect 755 18165 805 18195
rect 835 18165 885 18195
rect 915 18165 965 18195
rect 995 18165 1045 18195
rect 1075 18165 1125 18195
rect 1155 18165 1205 18195
rect 1235 18165 1285 18195
rect 1315 18165 1365 18195
rect 1395 18165 1445 18195
rect 1475 18165 1525 18195
rect 1555 18165 1605 18195
rect 1635 18165 1685 18195
rect 1715 18165 1765 18195
rect 1795 18165 1845 18195
rect 1875 18165 1925 18195
rect 1955 18165 2005 18195
rect 2035 18165 2085 18195
rect 2115 18165 2165 18195
rect 2195 18165 2245 18195
rect 2275 18165 2325 18195
rect 2355 18165 2405 18195
rect 2435 18165 2485 18195
rect 2515 18165 2565 18195
rect 2595 18165 2645 18195
rect 2675 18165 2725 18195
rect 2755 18165 2805 18195
rect 2835 18165 2885 18195
rect 2915 18165 2965 18195
rect 2995 18165 3045 18195
rect 3075 18165 3125 18195
rect 3155 18165 3205 18195
rect 3235 18165 3285 18195
rect 3315 18165 3365 18195
rect 3395 18165 3445 18195
rect 3475 18165 3525 18195
rect 3555 18165 3605 18195
rect 3635 18165 3685 18195
rect 3715 18165 3765 18195
rect 3795 18165 3845 18195
rect 3875 18165 3925 18195
rect 3955 18165 4005 18195
rect 4035 18165 4085 18195
rect 4115 18165 4165 18195
rect 4195 18165 4725 18195
rect 4755 18165 4885 18195
rect 4915 18165 5045 18195
rect 5075 18165 5205 18195
rect 5235 18165 5365 18195
rect 5395 18165 5525 18195
rect 5555 18165 5685 18195
rect 5715 18165 6245 18195
rect 6275 18165 6325 18195
rect 6355 18165 6405 18195
rect 6435 18165 6485 18195
rect 6515 18165 6565 18195
rect 6595 18165 6645 18195
rect 6675 18165 6725 18195
rect 6755 18165 6805 18195
rect 6835 18165 6885 18195
rect 6915 18165 6965 18195
rect 6995 18165 7045 18195
rect 7075 18165 7125 18195
rect 7155 18165 7205 18195
rect 7235 18165 7285 18195
rect 7315 18165 7365 18195
rect 7395 18165 7445 18195
rect 7475 18165 7525 18195
rect 7555 18165 7605 18195
rect 7635 18165 7685 18195
rect 7715 18165 7765 18195
rect 7795 18165 7845 18195
rect 7875 18165 7925 18195
rect 7955 18165 8005 18195
rect 8035 18165 8085 18195
rect 8115 18165 8165 18195
rect 8195 18165 8245 18195
rect 8275 18165 8325 18195
rect 8355 18165 8405 18195
rect 8435 18165 8485 18195
rect 8515 18165 8565 18195
rect 8595 18165 8645 18195
rect 8675 18165 8725 18195
rect 8755 18165 8805 18195
rect 8835 18165 8885 18195
rect 8915 18165 8965 18195
rect 8995 18165 9045 18195
rect 9075 18165 9125 18195
rect 9155 18165 9205 18195
rect 9235 18165 9285 18195
rect 9315 18165 9365 18195
rect 9395 18165 9445 18195
rect 9475 18165 10005 18195
rect 10035 18165 10165 18195
rect 10195 18165 10325 18195
rect 10355 18165 10485 18195
rect 10515 18165 10645 18195
rect 10675 18165 10805 18195
rect 10835 18165 10965 18195
rect 10995 18165 11565 18195
rect 11595 18165 11645 18195
rect 11675 18165 11725 18195
rect 11755 18165 11805 18195
rect 11835 18165 11885 18195
rect 11915 18165 11965 18195
rect 11995 18165 12045 18195
rect 12075 18165 12125 18195
rect 12155 18165 12205 18195
rect 12235 18165 12285 18195
rect 12315 18165 12365 18195
rect 12395 18165 12445 18195
rect 12475 18165 12525 18195
rect 12555 18165 12605 18195
rect 12635 18165 12685 18195
rect 12715 18165 12765 18195
rect 12795 18165 12845 18195
rect 12875 18165 12925 18195
rect 12955 18165 13005 18195
rect 13035 18165 13085 18195
rect 13115 18165 13165 18195
rect 13195 18165 13245 18195
rect 13275 18165 13325 18195
rect 13355 18165 13405 18195
rect 13435 18165 13485 18195
rect 13515 18165 13565 18195
rect 13595 18165 13645 18195
rect 13675 18165 13725 18195
rect 13755 18165 13805 18195
rect 13835 18165 13885 18195
rect 13915 18165 13965 18195
rect 13995 18165 14045 18195
rect 14075 18165 14125 18195
rect 14155 18165 14205 18195
rect 14235 18165 14285 18195
rect 14315 18165 14365 18195
rect 14395 18165 14445 18195
rect 14475 18165 14525 18195
rect 14555 18165 14605 18195
rect 14635 18165 14685 18195
rect 14715 18165 15245 18195
rect 15275 18165 15405 18195
rect 15435 18165 15565 18195
rect 15595 18165 15725 18195
rect 15755 18165 15885 18195
rect 15915 18165 16045 18195
rect 16075 18165 16205 18195
rect 16235 18165 16765 18195
rect 16795 18165 16845 18195
rect 16875 18165 16925 18195
rect 16955 18165 17005 18195
rect 17035 18165 17085 18195
rect 17115 18165 17165 18195
rect 17195 18165 17245 18195
rect 17275 18165 17325 18195
rect 17355 18165 17405 18195
rect 17435 18165 17485 18195
rect 17515 18165 17565 18195
rect 17595 18165 17645 18195
rect 17675 18165 17725 18195
rect 17755 18165 17805 18195
rect 17835 18165 17885 18195
rect 17915 18165 17965 18195
rect 17995 18165 18045 18195
rect 18075 18165 18125 18195
rect 18155 18165 18205 18195
rect 18235 18165 18285 18195
rect 18315 18165 18365 18195
rect 18395 18165 18445 18195
rect 18475 18165 18525 18195
rect 18555 18165 18605 18195
rect 18635 18165 18685 18195
rect 18715 18165 18765 18195
rect 18795 18165 18845 18195
rect 18875 18165 18925 18195
rect 18955 18165 19005 18195
rect 19035 18165 19085 18195
rect 19115 18165 19165 18195
rect 19195 18165 19245 18195
rect 19275 18165 19325 18195
rect 19355 18165 19405 18195
rect 19435 18165 19485 18195
rect 19515 18165 19565 18195
rect 19595 18165 19645 18195
rect 19675 18165 19725 18195
rect 19755 18165 19805 18195
rect 19835 18165 19885 18195
rect 19915 18165 19965 18195
rect 19995 18165 20045 18195
rect 20075 18165 20125 18195
rect 20155 18165 20205 18195
rect 20235 18165 20285 18195
rect 20315 18165 20365 18195
rect 20395 18165 20445 18195
rect 20475 18165 20525 18195
rect 20555 18165 20605 18195
rect 20635 18165 20685 18195
rect 20715 18165 20765 18195
rect 20795 18165 20845 18195
rect 20875 18165 20925 18195
rect 20955 18165 20960 18195
rect 0 18160 20960 18165
rect 0 18115 20960 18120
rect 0 18085 4805 18115
rect 4835 18085 10885 18115
rect 10915 18085 16125 18115
rect 16155 18085 20960 18115
rect 0 18080 20960 18085
rect 0 18035 20960 18040
rect 0 18005 5 18035
rect 35 18005 85 18035
rect 115 18005 165 18035
rect 195 18005 245 18035
rect 275 18005 325 18035
rect 355 18005 405 18035
rect 435 18005 485 18035
rect 515 18005 565 18035
rect 595 18005 645 18035
rect 675 18005 725 18035
rect 755 18005 805 18035
rect 835 18005 885 18035
rect 915 18005 965 18035
rect 995 18005 1045 18035
rect 1075 18005 1125 18035
rect 1155 18005 1205 18035
rect 1235 18005 1285 18035
rect 1315 18005 1365 18035
rect 1395 18005 1445 18035
rect 1475 18005 1525 18035
rect 1555 18005 1605 18035
rect 1635 18005 1685 18035
rect 1715 18005 1765 18035
rect 1795 18005 1845 18035
rect 1875 18005 1925 18035
rect 1955 18005 2005 18035
rect 2035 18005 2085 18035
rect 2115 18005 2165 18035
rect 2195 18005 2245 18035
rect 2275 18005 2325 18035
rect 2355 18005 2405 18035
rect 2435 18005 2485 18035
rect 2515 18005 2565 18035
rect 2595 18005 2645 18035
rect 2675 18005 2725 18035
rect 2755 18005 2805 18035
rect 2835 18005 2885 18035
rect 2915 18005 2965 18035
rect 2995 18005 3045 18035
rect 3075 18005 3125 18035
rect 3155 18005 3205 18035
rect 3235 18005 3285 18035
rect 3315 18005 3365 18035
rect 3395 18005 3445 18035
rect 3475 18005 3525 18035
rect 3555 18005 3605 18035
rect 3635 18005 3685 18035
rect 3715 18005 3765 18035
rect 3795 18005 3845 18035
rect 3875 18005 3925 18035
rect 3955 18005 4005 18035
rect 4035 18005 4085 18035
rect 4115 18005 4165 18035
rect 4195 18005 4725 18035
rect 4755 18005 4885 18035
rect 4915 18005 5045 18035
rect 5075 18005 5205 18035
rect 5235 18005 5365 18035
rect 5395 18005 5525 18035
rect 5555 18005 5685 18035
rect 5715 18005 6245 18035
rect 6275 18005 6325 18035
rect 6355 18005 6405 18035
rect 6435 18005 6485 18035
rect 6515 18005 6565 18035
rect 6595 18005 6645 18035
rect 6675 18005 6725 18035
rect 6755 18005 6805 18035
rect 6835 18005 6885 18035
rect 6915 18005 6965 18035
rect 6995 18005 7045 18035
rect 7075 18005 7125 18035
rect 7155 18005 7205 18035
rect 7235 18005 7285 18035
rect 7315 18005 7365 18035
rect 7395 18005 7445 18035
rect 7475 18005 7525 18035
rect 7555 18005 7605 18035
rect 7635 18005 7685 18035
rect 7715 18005 7765 18035
rect 7795 18005 7845 18035
rect 7875 18005 7925 18035
rect 7955 18005 8005 18035
rect 8035 18005 8085 18035
rect 8115 18005 8165 18035
rect 8195 18005 8245 18035
rect 8275 18005 8325 18035
rect 8355 18005 8405 18035
rect 8435 18005 8485 18035
rect 8515 18005 8565 18035
rect 8595 18005 8645 18035
rect 8675 18005 8725 18035
rect 8755 18005 8805 18035
rect 8835 18005 8885 18035
rect 8915 18005 8965 18035
rect 8995 18005 9045 18035
rect 9075 18005 9125 18035
rect 9155 18005 9205 18035
rect 9235 18005 9285 18035
rect 9315 18005 9365 18035
rect 9395 18005 9445 18035
rect 9475 18005 10005 18035
rect 10035 18005 10165 18035
rect 10195 18005 10325 18035
rect 10355 18005 10485 18035
rect 10515 18005 10645 18035
rect 10675 18005 10805 18035
rect 10835 18005 10965 18035
rect 10995 18005 11565 18035
rect 11595 18005 11645 18035
rect 11675 18005 11725 18035
rect 11755 18005 11805 18035
rect 11835 18005 11885 18035
rect 11915 18005 11965 18035
rect 11995 18005 12045 18035
rect 12075 18005 12125 18035
rect 12155 18005 12205 18035
rect 12235 18005 12285 18035
rect 12315 18005 12365 18035
rect 12395 18005 12445 18035
rect 12475 18005 12525 18035
rect 12555 18005 12605 18035
rect 12635 18005 12685 18035
rect 12715 18005 12765 18035
rect 12795 18005 12845 18035
rect 12875 18005 12925 18035
rect 12955 18005 13005 18035
rect 13035 18005 13085 18035
rect 13115 18005 13165 18035
rect 13195 18005 13245 18035
rect 13275 18005 13325 18035
rect 13355 18005 13405 18035
rect 13435 18005 13485 18035
rect 13515 18005 13565 18035
rect 13595 18005 13645 18035
rect 13675 18005 13725 18035
rect 13755 18005 13805 18035
rect 13835 18005 13885 18035
rect 13915 18005 13965 18035
rect 13995 18005 14045 18035
rect 14075 18005 14125 18035
rect 14155 18005 14205 18035
rect 14235 18005 14285 18035
rect 14315 18005 14365 18035
rect 14395 18005 14445 18035
rect 14475 18005 14525 18035
rect 14555 18005 14605 18035
rect 14635 18005 14685 18035
rect 14715 18005 15245 18035
rect 15275 18005 15405 18035
rect 15435 18005 15565 18035
rect 15595 18005 15725 18035
rect 15755 18005 15885 18035
rect 15915 18005 16045 18035
rect 16075 18005 16205 18035
rect 16235 18005 16765 18035
rect 16795 18005 16845 18035
rect 16875 18005 16925 18035
rect 16955 18005 17005 18035
rect 17035 18005 17085 18035
rect 17115 18005 17165 18035
rect 17195 18005 17245 18035
rect 17275 18005 17325 18035
rect 17355 18005 17405 18035
rect 17435 18005 17485 18035
rect 17515 18005 17565 18035
rect 17595 18005 17645 18035
rect 17675 18005 17725 18035
rect 17755 18005 17805 18035
rect 17835 18005 17885 18035
rect 17915 18005 17965 18035
rect 17995 18005 18045 18035
rect 18075 18005 18125 18035
rect 18155 18005 18205 18035
rect 18235 18005 18285 18035
rect 18315 18005 18365 18035
rect 18395 18005 18445 18035
rect 18475 18005 18525 18035
rect 18555 18005 18605 18035
rect 18635 18005 18685 18035
rect 18715 18005 18765 18035
rect 18795 18005 18845 18035
rect 18875 18005 18925 18035
rect 18955 18005 19005 18035
rect 19035 18005 19085 18035
rect 19115 18005 19165 18035
rect 19195 18005 19245 18035
rect 19275 18005 19325 18035
rect 19355 18005 19405 18035
rect 19435 18005 19485 18035
rect 19515 18005 19565 18035
rect 19595 18005 19645 18035
rect 19675 18005 19725 18035
rect 19755 18005 19805 18035
rect 19835 18005 19885 18035
rect 19915 18005 19965 18035
rect 19995 18005 20045 18035
rect 20075 18005 20125 18035
rect 20155 18005 20205 18035
rect 20235 18005 20285 18035
rect 20315 18005 20365 18035
rect 20395 18005 20445 18035
rect 20475 18005 20525 18035
rect 20555 18005 20605 18035
rect 20635 18005 20685 18035
rect 20715 18005 20765 18035
rect 20795 18005 20845 18035
rect 20875 18005 20925 18035
rect 20955 18005 20960 18035
rect 0 18000 20960 18005
rect 0 17955 20960 17960
rect 0 17925 4965 17955
rect 4995 17925 10725 17955
rect 10755 17925 15965 17955
rect 15995 17925 20960 17955
rect 0 17920 20960 17925
rect 0 17875 20960 17880
rect 0 17845 5 17875
rect 35 17845 85 17875
rect 115 17845 165 17875
rect 195 17845 245 17875
rect 275 17845 325 17875
rect 355 17845 405 17875
rect 435 17845 485 17875
rect 515 17845 565 17875
rect 595 17845 645 17875
rect 675 17845 725 17875
rect 755 17845 805 17875
rect 835 17845 885 17875
rect 915 17845 965 17875
rect 995 17845 1045 17875
rect 1075 17845 1125 17875
rect 1155 17845 1205 17875
rect 1235 17845 1285 17875
rect 1315 17845 1365 17875
rect 1395 17845 1445 17875
rect 1475 17845 1525 17875
rect 1555 17845 1605 17875
rect 1635 17845 1685 17875
rect 1715 17845 1765 17875
rect 1795 17845 1845 17875
rect 1875 17845 1925 17875
rect 1955 17845 2005 17875
rect 2035 17845 2085 17875
rect 2115 17845 2165 17875
rect 2195 17845 2245 17875
rect 2275 17845 2325 17875
rect 2355 17845 2405 17875
rect 2435 17845 2485 17875
rect 2515 17845 2565 17875
rect 2595 17845 2645 17875
rect 2675 17845 2725 17875
rect 2755 17845 2805 17875
rect 2835 17845 2885 17875
rect 2915 17845 2965 17875
rect 2995 17845 3045 17875
rect 3075 17845 3125 17875
rect 3155 17845 3205 17875
rect 3235 17845 3285 17875
rect 3315 17845 3365 17875
rect 3395 17845 3445 17875
rect 3475 17845 3525 17875
rect 3555 17845 3605 17875
rect 3635 17845 3685 17875
rect 3715 17845 3765 17875
rect 3795 17845 3845 17875
rect 3875 17845 3925 17875
rect 3955 17845 4005 17875
rect 4035 17845 4085 17875
rect 4115 17845 4165 17875
rect 4195 17845 4725 17875
rect 4755 17845 4885 17875
rect 4915 17845 5045 17875
rect 5075 17845 5205 17875
rect 5235 17845 5365 17875
rect 5395 17845 5525 17875
rect 5555 17845 5685 17875
rect 5715 17845 6245 17875
rect 6275 17845 6325 17875
rect 6355 17845 6405 17875
rect 6435 17845 6485 17875
rect 6515 17845 6565 17875
rect 6595 17845 6645 17875
rect 6675 17845 6725 17875
rect 6755 17845 6805 17875
rect 6835 17845 6885 17875
rect 6915 17845 6965 17875
rect 6995 17845 7045 17875
rect 7075 17845 7125 17875
rect 7155 17845 7205 17875
rect 7235 17845 7285 17875
rect 7315 17845 7365 17875
rect 7395 17845 7445 17875
rect 7475 17845 7525 17875
rect 7555 17845 7605 17875
rect 7635 17845 7685 17875
rect 7715 17845 7765 17875
rect 7795 17845 7845 17875
rect 7875 17845 7925 17875
rect 7955 17845 8005 17875
rect 8035 17845 8085 17875
rect 8115 17845 8165 17875
rect 8195 17845 8245 17875
rect 8275 17845 8325 17875
rect 8355 17845 8405 17875
rect 8435 17845 8485 17875
rect 8515 17845 8565 17875
rect 8595 17845 8645 17875
rect 8675 17845 8725 17875
rect 8755 17845 8805 17875
rect 8835 17845 8885 17875
rect 8915 17845 8965 17875
rect 8995 17845 9045 17875
rect 9075 17845 9125 17875
rect 9155 17845 9205 17875
rect 9235 17845 9285 17875
rect 9315 17845 9365 17875
rect 9395 17845 9445 17875
rect 9475 17845 10005 17875
rect 10035 17845 10165 17875
rect 10195 17845 10325 17875
rect 10355 17845 10485 17875
rect 10515 17845 10645 17875
rect 10675 17845 10805 17875
rect 10835 17845 10965 17875
rect 10995 17845 11565 17875
rect 11595 17845 11645 17875
rect 11675 17845 11725 17875
rect 11755 17845 11805 17875
rect 11835 17845 11885 17875
rect 11915 17845 11965 17875
rect 11995 17845 12045 17875
rect 12075 17845 12125 17875
rect 12155 17845 12205 17875
rect 12235 17845 12285 17875
rect 12315 17845 12365 17875
rect 12395 17845 12445 17875
rect 12475 17845 12525 17875
rect 12555 17845 12605 17875
rect 12635 17845 12685 17875
rect 12715 17845 12765 17875
rect 12795 17845 12845 17875
rect 12875 17845 12925 17875
rect 12955 17845 13005 17875
rect 13035 17845 13085 17875
rect 13115 17845 13165 17875
rect 13195 17845 13245 17875
rect 13275 17845 13325 17875
rect 13355 17845 13405 17875
rect 13435 17845 13485 17875
rect 13515 17845 13565 17875
rect 13595 17845 13645 17875
rect 13675 17845 13725 17875
rect 13755 17845 13805 17875
rect 13835 17845 13885 17875
rect 13915 17845 13965 17875
rect 13995 17845 14045 17875
rect 14075 17845 14125 17875
rect 14155 17845 14205 17875
rect 14235 17845 14285 17875
rect 14315 17845 14365 17875
rect 14395 17845 14445 17875
rect 14475 17845 14525 17875
rect 14555 17845 14605 17875
rect 14635 17845 14685 17875
rect 14715 17845 15245 17875
rect 15275 17845 15405 17875
rect 15435 17845 15565 17875
rect 15595 17845 15725 17875
rect 15755 17845 15885 17875
rect 15915 17845 16045 17875
rect 16075 17845 16205 17875
rect 16235 17845 16765 17875
rect 16795 17845 16845 17875
rect 16875 17845 16925 17875
rect 16955 17845 17005 17875
rect 17035 17845 17085 17875
rect 17115 17845 17165 17875
rect 17195 17845 17245 17875
rect 17275 17845 17325 17875
rect 17355 17845 17405 17875
rect 17435 17845 17485 17875
rect 17515 17845 17565 17875
rect 17595 17845 17645 17875
rect 17675 17845 17725 17875
rect 17755 17845 17805 17875
rect 17835 17845 17885 17875
rect 17915 17845 17965 17875
rect 17995 17845 18045 17875
rect 18075 17845 18125 17875
rect 18155 17845 18205 17875
rect 18235 17845 18285 17875
rect 18315 17845 18365 17875
rect 18395 17845 18445 17875
rect 18475 17845 18525 17875
rect 18555 17845 18605 17875
rect 18635 17845 18685 17875
rect 18715 17845 18765 17875
rect 18795 17845 18845 17875
rect 18875 17845 18925 17875
rect 18955 17845 19005 17875
rect 19035 17845 19085 17875
rect 19115 17845 19165 17875
rect 19195 17845 19245 17875
rect 19275 17845 19325 17875
rect 19355 17845 19405 17875
rect 19435 17845 19485 17875
rect 19515 17845 19565 17875
rect 19595 17845 19645 17875
rect 19675 17845 19725 17875
rect 19755 17845 19805 17875
rect 19835 17845 19885 17875
rect 19915 17845 19965 17875
rect 19995 17845 20045 17875
rect 20075 17845 20125 17875
rect 20155 17845 20205 17875
rect 20235 17845 20285 17875
rect 20315 17845 20365 17875
rect 20395 17845 20445 17875
rect 20475 17845 20525 17875
rect 20555 17845 20605 17875
rect 20635 17845 20685 17875
rect 20715 17845 20765 17875
rect 20795 17845 20845 17875
rect 20875 17845 20925 17875
rect 20955 17845 20960 17875
rect 0 17840 20960 17845
rect 0 17795 20960 17800
rect 0 17765 5125 17795
rect 5155 17765 10565 17795
rect 10595 17765 15805 17795
rect 15835 17765 20960 17795
rect 0 17760 20960 17765
rect 0 17715 20960 17720
rect 0 17685 5 17715
rect 35 17685 85 17715
rect 115 17685 165 17715
rect 195 17685 245 17715
rect 275 17685 325 17715
rect 355 17685 405 17715
rect 435 17685 485 17715
rect 515 17685 565 17715
rect 595 17685 645 17715
rect 675 17685 725 17715
rect 755 17685 805 17715
rect 835 17685 885 17715
rect 915 17685 965 17715
rect 995 17685 1045 17715
rect 1075 17685 1125 17715
rect 1155 17685 1205 17715
rect 1235 17685 1285 17715
rect 1315 17685 1365 17715
rect 1395 17685 1445 17715
rect 1475 17685 1525 17715
rect 1555 17685 1605 17715
rect 1635 17685 1685 17715
rect 1715 17685 1765 17715
rect 1795 17685 1845 17715
rect 1875 17685 1925 17715
rect 1955 17685 2005 17715
rect 2035 17685 2085 17715
rect 2115 17685 2165 17715
rect 2195 17685 2245 17715
rect 2275 17685 2325 17715
rect 2355 17685 2405 17715
rect 2435 17685 2485 17715
rect 2515 17685 2565 17715
rect 2595 17685 2645 17715
rect 2675 17685 2725 17715
rect 2755 17685 2805 17715
rect 2835 17685 2885 17715
rect 2915 17685 2965 17715
rect 2995 17685 3045 17715
rect 3075 17685 3125 17715
rect 3155 17685 3205 17715
rect 3235 17685 3285 17715
rect 3315 17685 3365 17715
rect 3395 17685 3445 17715
rect 3475 17685 3525 17715
rect 3555 17685 3605 17715
rect 3635 17685 3685 17715
rect 3715 17685 3765 17715
rect 3795 17685 3845 17715
rect 3875 17685 3925 17715
rect 3955 17685 4005 17715
rect 4035 17685 4085 17715
rect 4115 17685 4165 17715
rect 4195 17685 4725 17715
rect 4755 17685 4885 17715
rect 4915 17685 5045 17715
rect 5075 17685 5205 17715
rect 5235 17685 5365 17715
rect 5395 17685 5525 17715
rect 5555 17685 5685 17715
rect 5715 17685 6245 17715
rect 6275 17685 6325 17715
rect 6355 17685 6405 17715
rect 6435 17685 6485 17715
rect 6515 17685 6565 17715
rect 6595 17685 6645 17715
rect 6675 17685 6725 17715
rect 6755 17685 6805 17715
rect 6835 17685 6885 17715
rect 6915 17685 6965 17715
rect 6995 17685 7045 17715
rect 7075 17685 7125 17715
rect 7155 17685 7205 17715
rect 7235 17685 7285 17715
rect 7315 17685 7365 17715
rect 7395 17685 7445 17715
rect 7475 17685 7525 17715
rect 7555 17685 7605 17715
rect 7635 17685 7685 17715
rect 7715 17685 7765 17715
rect 7795 17685 7845 17715
rect 7875 17685 7925 17715
rect 7955 17685 8005 17715
rect 8035 17685 8085 17715
rect 8115 17685 8165 17715
rect 8195 17685 8245 17715
rect 8275 17685 8325 17715
rect 8355 17685 8405 17715
rect 8435 17685 8485 17715
rect 8515 17685 8565 17715
rect 8595 17685 8645 17715
rect 8675 17685 8725 17715
rect 8755 17685 8805 17715
rect 8835 17685 8885 17715
rect 8915 17685 8965 17715
rect 8995 17685 9045 17715
rect 9075 17685 9125 17715
rect 9155 17685 9205 17715
rect 9235 17685 9285 17715
rect 9315 17685 9365 17715
rect 9395 17685 9445 17715
rect 9475 17685 10005 17715
rect 10035 17685 10165 17715
rect 10195 17685 10325 17715
rect 10355 17685 10485 17715
rect 10515 17685 10645 17715
rect 10675 17685 10805 17715
rect 10835 17685 10965 17715
rect 10995 17685 11565 17715
rect 11595 17685 11645 17715
rect 11675 17685 11725 17715
rect 11755 17685 11805 17715
rect 11835 17685 11885 17715
rect 11915 17685 11965 17715
rect 11995 17685 12045 17715
rect 12075 17685 12125 17715
rect 12155 17685 12205 17715
rect 12235 17685 12285 17715
rect 12315 17685 12365 17715
rect 12395 17685 12445 17715
rect 12475 17685 12525 17715
rect 12555 17685 12605 17715
rect 12635 17685 12685 17715
rect 12715 17685 12765 17715
rect 12795 17685 12845 17715
rect 12875 17685 12925 17715
rect 12955 17685 13005 17715
rect 13035 17685 13085 17715
rect 13115 17685 13165 17715
rect 13195 17685 13245 17715
rect 13275 17685 13325 17715
rect 13355 17685 13405 17715
rect 13435 17685 13485 17715
rect 13515 17685 13565 17715
rect 13595 17685 13645 17715
rect 13675 17685 13725 17715
rect 13755 17685 13805 17715
rect 13835 17685 13885 17715
rect 13915 17685 13965 17715
rect 13995 17685 14045 17715
rect 14075 17685 14125 17715
rect 14155 17685 14205 17715
rect 14235 17685 14285 17715
rect 14315 17685 14365 17715
rect 14395 17685 14445 17715
rect 14475 17685 14525 17715
rect 14555 17685 14605 17715
rect 14635 17685 14685 17715
rect 14715 17685 15245 17715
rect 15275 17685 15405 17715
rect 15435 17685 15565 17715
rect 15595 17685 15725 17715
rect 15755 17685 15885 17715
rect 15915 17685 16045 17715
rect 16075 17685 16205 17715
rect 16235 17685 16765 17715
rect 16795 17685 16845 17715
rect 16875 17685 16925 17715
rect 16955 17685 17005 17715
rect 17035 17685 17085 17715
rect 17115 17685 17165 17715
rect 17195 17685 17245 17715
rect 17275 17685 17325 17715
rect 17355 17685 17405 17715
rect 17435 17685 17485 17715
rect 17515 17685 17565 17715
rect 17595 17685 17645 17715
rect 17675 17685 17725 17715
rect 17755 17685 17805 17715
rect 17835 17685 17885 17715
rect 17915 17685 17965 17715
rect 17995 17685 18045 17715
rect 18075 17685 18125 17715
rect 18155 17685 18205 17715
rect 18235 17685 18285 17715
rect 18315 17685 18365 17715
rect 18395 17685 18445 17715
rect 18475 17685 18525 17715
rect 18555 17685 18605 17715
rect 18635 17685 18685 17715
rect 18715 17685 18765 17715
rect 18795 17685 18845 17715
rect 18875 17685 18925 17715
rect 18955 17685 19005 17715
rect 19035 17685 19085 17715
rect 19115 17685 19165 17715
rect 19195 17685 19245 17715
rect 19275 17685 19325 17715
rect 19355 17685 19405 17715
rect 19435 17685 19485 17715
rect 19515 17685 19565 17715
rect 19595 17685 19645 17715
rect 19675 17685 19725 17715
rect 19755 17685 19805 17715
rect 19835 17685 19885 17715
rect 19915 17685 19965 17715
rect 19995 17685 20045 17715
rect 20075 17685 20125 17715
rect 20155 17685 20205 17715
rect 20235 17685 20285 17715
rect 20315 17685 20365 17715
rect 20395 17685 20445 17715
rect 20475 17685 20525 17715
rect 20555 17685 20605 17715
rect 20635 17685 20685 17715
rect 20715 17685 20765 17715
rect 20795 17685 20845 17715
rect 20875 17685 20925 17715
rect 20955 17685 20960 17715
rect 0 17680 20960 17685
rect 0 17635 20960 17640
rect 0 17605 5285 17635
rect 5315 17605 10405 17635
rect 10435 17605 15645 17635
rect 15675 17605 20960 17635
rect 0 17600 20960 17605
rect 0 17555 20960 17560
rect 0 17525 5 17555
rect 35 17525 85 17555
rect 115 17525 165 17555
rect 195 17525 245 17555
rect 275 17525 325 17555
rect 355 17525 405 17555
rect 435 17525 485 17555
rect 515 17525 565 17555
rect 595 17525 645 17555
rect 675 17525 725 17555
rect 755 17525 805 17555
rect 835 17525 885 17555
rect 915 17525 965 17555
rect 995 17525 1045 17555
rect 1075 17525 1125 17555
rect 1155 17525 1205 17555
rect 1235 17525 1285 17555
rect 1315 17525 1365 17555
rect 1395 17525 1445 17555
rect 1475 17525 1525 17555
rect 1555 17525 1605 17555
rect 1635 17525 1685 17555
rect 1715 17525 1765 17555
rect 1795 17525 1845 17555
rect 1875 17525 1925 17555
rect 1955 17525 2005 17555
rect 2035 17525 2085 17555
rect 2115 17525 2165 17555
rect 2195 17525 2245 17555
rect 2275 17525 2325 17555
rect 2355 17525 2405 17555
rect 2435 17525 2485 17555
rect 2515 17525 2565 17555
rect 2595 17525 2645 17555
rect 2675 17525 2725 17555
rect 2755 17525 2805 17555
rect 2835 17525 2885 17555
rect 2915 17525 2965 17555
rect 2995 17525 3045 17555
rect 3075 17525 3125 17555
rect 3155 17525 3205 17555
rect 3235 17525 3285 17555
rect 3315 17525 3365 17555
rect 3395 17525 3445 17555
rect 3475 17525 3525 17555
rect 3555 17525 3605 17555
rect 3635 17525 3685 17555
rect 3715 17525 3765 17555
rect 3795 17525 3845 17555
rect 3875 17525 3925 17555
rect 3955 17525 4005 17555
rect 4035 17525 4085 17555
rect 4115 17525 4165 17555
rect 4195 17525 4725 17555
rect 4755 17525 4885 17555
rect 4915 17525 5045 17555
rect 5075 17525 5205 17555
rect 5235 17525 5365 17555
rect 5395 17525 5525 17555
rect 5555 17525 5685 17555
rect 5715 17525 6245 17555
rect 6275 17525 6325 17555
rect 6355 17525 6405 17555
rect 6435 17525 6485 17555
rect 6515 17525 6565 17555
rect 6595 17525 6645 17555
rect 6675 17525 6725 17555
rect 6755 17525 6805 17555
rect 6835 17525 6885 17555
rect 6915 17525 6965 17555
rect 6995 17525 7045 17555
rect 7075 17525 7125 17555
rect 7155 17525 7205 17555
rect 7235 17525 7285 17555
rect 7315 17525 7365 17555
rect 7395 17525 7445 17555
rect 7475 17525 7525 17555
rect 7555 17525 7605 17555
rect 7635 17525 7685 17555
rect 7715 17525 7765 17555
rect 7795 17525 7845 17555
rect 7875 17525 7925 17555
rect 7955 17525 8005 17555
rect 8035 17525 8085 17555
rect 8115 17525 8165 17555
rect 8195 17525 8245 17555
rect 8275 17525 8325 17555
rect 8355 17525 8405 17555
rect 8435 17525 8485 17555
rect 8515 17525 8565 17555
rect 8595 17525 8645 17555
rect 8675 17525 8725 17555
rect 8755 17525 8805 17555
rect 8835 17525 8885 17555
rect 8915 17525 8965 17555
rect 8995 17525 9045 17555
rect 9075 17525 9125 17555
rect 9155 17525 9205 17555
rect 9235 17525 9285 17555
rect 9315 17525 9365 17555
rect 9395 17525 9445 17555
rect 9475 17525 10005 17555
rect 10035 17525 10165 17555
rect 10195 17525 10325 17555
rect 10355 17525 10485 17555
rect 10515 17525 10645 17555
rect 10675 17525 10805 17555
rect 10835 17525 10965 17555
rect 10995 17525 11565 17555
rect 11595 17525 11645 17555
rect 11675 17525 11725 17555
rect 11755 17525 11805 17555
rect 11835 17525 11885 17555
rect 11915 17525 11965 17555
rect 11995 17525 12045 17555
rect 12075 17525 12125 17555
rect 12155 17525 12205 17555
rect 12235 17525 12285 17555
rect 12315 17525 12365 17555
rect 12395 17525 12445 17555
rect 12475 17525 12525 17555
rect 12555 17525 12605 17555
rect 12635 17525 12685 17555
rect 12715 17525 12765 17555
rect 12795 17525 12845 17555
rect 12875 17525 12925 17555
rect 12955 17525 13005 17555
rect 13035 17525 13085 17555
rect 13115 17525 13165 17555
rect 13195 17525 13245 17555
rect 13275 17525 13325 17555
rect 13355 17525 13405 17555
rect 13435 17525 13485 17555
rect 13515 17525 13565 17555
rect 13595 17525 13645 17555
rect 13675 17525 13725 17555
rect 13755 17525 13805 17555
rect 13835 17525 13885 17555
rect 13915 17525 13965 17555
rect 13995 17525 14045 17555
rect 14075 17525 14125 17555
rect 14155 17525 14205 17555
rect 14235 17525 14285 17555
rect 14315 17525 14365 17555
rect 14395 17525 14445 17555
rect 14475 17525 14525 17555
rect 14555 17525 14605 17555
rect 14635 17525 14685 17555
rect 14715 17525 15245 17555
rect 15275 17525 15405 17555
rect 15435 17525 15565 17555
rect 15595 17525 15725 17555
rect 15755 17525 15885 17555
rect 15915 17525 16045 17555
rect 16075 17525 16205 17555
rect 16235 17525 16765 17555
rect 16795 17525 16845 17555
rect 16875 17525 16925 17555
rect 16955 17525 17005 17555
rect 17035 17525 17085 17555
rect 17115 17525 17165 17555
rect 17195 17525 17245 17555
rect 17275 17525 17325 17555
rect 17355 17525 17405 17555
rect 17435 17525 17485 17555
rect 17515 17525 17565 17555
rect 17595 17525 17645 17555
rect 17675 17525 17725 17555
rect 17755 17525 17805 17555
rect 17835 17525 17885 17555
rect 17915 17525 17965 17555
rect 17995 17525 18045 17555
rect 18075 17525 18125 17555
rect 18155 17525 18205 17555
rect 18235 17525 18285 17555
rect 18315 17525 18365 17555
rect 18395 17525 18445 17555
rect 18475 17525 18525 17555
rect 18555 17525 18605 17555
rect 18635 17525 18685 17555
rect 18715 17525 18765 17555
rect 18795 17525 18845 17555
rect 18875 17525 18925 17555
rect 18955 17525 19005 17555
rect 19035 17525 19085 17555
rect 19115 17525 19165 17555
rect 19195 17525 19245 17555
rect 19275 17525 19325 17555
rect 19355 17525 19405 17555
rect 19435 17525 19485 17555
rect 19515 17525 19565 17555
rect 19595 17525 19645 17555
rect 19675 17525 19725 17555
rect 19755 17525 19805 17555
rect 19835 17525 19885 17555
rect 19915 17525 19965 17555
rect 19995 17525 20045 17555
rect 20075 17525 20125 17555
rect 20155 17525 20205 17555
rect 20235 17525 20285 17555
rect 20315 17525 20365 17555
rect 20395 17525 20445 17555
rect 20475 17525 20525 17555
rect 20555 17525 20605 17555
rect 20635 17525 20685 17555
rect 20715 17525 20765 17555
rect 20795 17525 20845 17555
rect 20875 17525 20925 17555
rect 20955 17525 20960 17555
rect 0 17520 20960 17525
rect 0 17475 20960 17480
rect 0 17445 5445 17475
rect 5475 17445 10245 17475
rect 10275 17445 15485 17475
rect 15515 17445 20960 17475
rect 0 17440 20960 17445
rect 0 17395 20960 17400
rect 0 17365 5 17395
rect 35 17365 85 17395
rect 115 17365 165 17395
rect 195 17365 245 17395
rect 275 17365 325 17395
rect 355 17365 405 17395
rect 435 17365 485 17395
rect 515 17365 565 17395
rect 595 17365 645 17395
rect 675 17365 725 17395
rect 755 17365 805 17395
rect 835 17365 885 17395
rect 915 17365 965 17395
rect 995 17365 1045 17395
rect 1075 17365 1125 17395
rect 1155 17365 1205 17395
rect 1235 17365 1285 17395
rect 1315 17365 1365 17395
rect 1395 17365 1445 17395
rect 1475 17365 1525 17395
rect 1555 17365 1605 17395
rect 1635 17365 1685 17395
rect 1715 17365 1765 17395
rect 1795 17365 1845 17395
rect 1875 17365 1925 17395
rect 1955 17365 2005 17395
rect 2035 17365 2085 17395
rect 2115 17365 2165 17395
rect 2195 17365 2245 17395
rect 2275 17365 2325 17395
rect 2355 17365 2405 17395
rect 2435 17365 2485 17395
rect 2515 17365 2565 17395
rect 2595 17365 2645 17395
rect 2675 17365 2725 17395
rect 2755 17365 2805 17395
rect 2835 17365 2885 17395
rect 2915 17365 2965 17395
rect 2995 17365 3045 17395
rect 3075 17365 3125 17395
rect 3155 17365 3205 17395
rect 3235 17365 3285 17395
rect 3315 17365 3365 17395
rect 3395 17365 3445 17395
rect 3475 17365 3525 17395
rect 3555 17365 3605 17395
rect 3635 17365 3685 17395
rect 3715 17365 3765 17395
rect 3795 17365 3845 17395
rect 3875 17365 3925 17395
rect 3955 17365 4005 17395
rect 4035 17365 4085 17395
rect 4115 17365 4165 17395
rect 4195 17365 4725 17395
rect 4755 17365 4885 17395
rect 4915 17365 5045 17395
rect 5075 17365 5205 17395
rect 5235 17365 5365 17395
rect 5395 17365 5525 17395
rect 5555 17365 5685 17395
rect 5715 17365 6245 17395
rect 6275 17365 6325 17395
rect 6355 17365 6405 17395
rect 6435 17365 6485 17395
rect 6515 17365 6565 17395
rect 6595 17365 6645 17395
rect 6675 17365 6725 17395
rect 6755 17365 6805 17395
rect 6835 17365 6885 17395
rect 6915 17365 6965 17395
rect 6995 17365 7045 17395
rect 7075 17365 7125 17395
rect 7155 17365 7205 17395
rect 7235 17365 7285 17395
rect 7315 17365 7365 17395
rect 7395 17365 7445 17395
rect 7475 17365 7525 17395
rect 7555 17365 7605 17395
rect 7635 17365 7685 17395
rect 7715 17365 7765 17395
rect 7795 17365 7845 17395
rect 7875 17365 7925 17395
rect 7955 17365 8005 17395
rect 8035 17365 8085 17395
rect 8115 17365 8165 17395
rect 8195 17365 8245 17395
rect 8275 17365 8325 17395
rect 8355 17365 8405 17395
rect 8435 17365 8485 17395
rect 8515 17365 8565 17395
rect 8595 17365 8645 17395
rect 8675 17365 8725 17395
rect 8755 17365 8805 17395
rect 8835 17365 8885 17395
rect 8915 17365 8965 17395
rect 8995 17365 9045 17395
rect 9075 17365 9125 17395
rect 9155 17365 9205 17395
rect 9235 17365 9285 17395
rect 9315 17365 9365 17395
rect 9395 17365 9445 17395
rect 9475 17365 10005 17395
rect 10035 17365 10165 17395
rect 10195 17365 10325 17395
rect 10355 17365 10485 17395
rect 10515 17365 10645 17395
rect 10675 17365 10805 17395
rect 10835 17365 10965 17395
rect 10995 17365 11565 17395
rect 11595 17365 11645 17395
rect 11675 17365 11725 17395
rect 11755 17365 11805 17395
rect 11835 17365 11885 17395
rect 11915 17365 11965 17395
rect 11995 17365 12045 17395
rect 12075 17365 12125 17395
rect 12155 17365 12205 17395
rect 12235 17365 12285 17395
rect 12315 17365 12365 17395
rect 12395 17365 12445 17395
rect 12475 17365 12525 17395
rect 12555 17365 12605 17395
rect 12635 17365 12685 17395
rect 12715 17365 12765 17395
rect 12795 17365 12845 17395
rect 12875 17365 12925 17395
rect 12955 17365 13005 17395
rect 13035 17365 13085 17395
rect 13115 17365 13165 17395
rect 13195 17365 13245 17395
rect 13275 17365 13325 17395
rect 13355 17365 13405 17395
rect 13435 17365 13485 17395
rect 13515 17365 13565 17395
rect 13595 17365 13645 17395
rect 13675 17365 13725 17395
rect 13755 17365 13805 17395
rect 13835 17365 13885 17395
rect 13915 17365 13965 17395
rect 13995 17365 14045 17395
rect 14075 17365 14125 17395
rect 14155 17365 14205 17395
rect 14235 17365 14285 17395
rect 14315 17365 14365 17395
rect 14395 17365 14445 17395
rect 14475 17365 14525 17395
rect 14555 17365 14605 17395
rect 14635 17365 14685 17395
rect 14715 17365 15245 17395
rect 15275 17365 15405 17395
rect 15435 17365 15565 17395
rect 15595 17365 15725 17395
rect 15755 17365 15885 17395
rect 15915 17365 16045 17395
rect 16075 17365 16205 17395
rect 16235 17365 16765 17395
rect 16795 17365 16845 17395
rect 16875 17365 16925 17395
rect 16955 17365 17005 17395
rect 17035 17365 17085 17395
rect 17115 17365 17165 17395
rect 17195 17365 17245 17395
rect 17275 17365 17325 17395
rect 17355 17365 17405 17395
rect 17435 17365 17485 17395
rect 17515 17365 17565 17395
rect 17595 17365 17645 17395
rect 17675 17365 17725 17395
rect 17755 17365 17805 17395
rect 17835 17365 17885 17395
rect 17915 17365 17965 17395
rect 17995 17365 18045 17395
rect 18075 17365 18125 17395
rect 18155 17365 18205 17395
rect 18235 17365 18285 17395
rect 18315 17365 18365 17395
rect 18395 17365 18445 17395
rect 18475 17365 18525 17395
rect 18555 17365 18605 17395
rect 18635 17365 18685 17395
rect 18715 17365 18765 17395
rect 18795 17365 18845 17395
rect 18875 17365 18925 17395
rect 18955 17365 19005 17395
rect 19035 17365 19085 17395
rect 19115 17365 19165 17395
rect 19195 17365 19245 17395
rect 19275 17365 19325 17395
rect 19355 17365 19405 17395
rect 19435 17365 19485 17395
rect 19515 17365 19565 17395
rect 19595 17365 19645 17395
rect 19675 17365 19725 17395
rect 19755 17365 19805 17395
rect 19835 17365 19885 17395
rect 19915 17365 19965 17395
rect 19995 17365 20045 17395
rect 20075 17365 20125 17395
rect 20155 17365 20205 17395
rect 20235 17365 20285 17395
rect 20315 17365 20365 17395
rect 20395 17365 20445 17395
rect 20475 17365 20525 17395
rect 20555 17365 20605 17395
rect 20635 17365 20685 17395
rect 20715 17365 20765 17395
rect 20795 17365 20845 17395
rect 20875 17365 20925 17395
rect 20955 17365 20960 17395
rect 0 17360 20960 17365
rect 0 17315 20960 17320
rect 0 17285 5605 17315
rect 5635 17285 10085 17315
rect 10115 17285 15325 17315
rect 15355 17285 20960 17315
rect 0 17280 20960 17285
rect 0 17235 20960 17240
rect 0 17205 5 17235
rect 35 17205 85 17235
rect 115 17205 165 17235
rect 195 17205 245 17235
rect 275 17205 325 17235
rect 355 17205 405 17235
rect 435 17205 485 17235
rect 515 17205 565 17235
rect 595 17205 645 17235
rect 675 17205 725 17235
rect 755 17205 805 17235
rect 835 17205 885 17235
rect 915 17205 965 17235
rect 995 17205 1045 17235
rect 1075 17205 1125 17235
rect 1155 17205 1205 17235
rect 1235 17205 1285 17235
rect 1315 17205 1365 17235
rect 1395 17205 1445 17235
rect 1475 17205 1525 17235
rect 1555 17205 1605 17235
rect 1635 17205 1685 17235
rect 1715 17205 1765 17235
rect 1795 17205 1845 17235
rect 1875 17205 1925 17235
rect 1955 17205 2005 17235
rect 2035 17205 2085 17235
rect 2115 17205 2165 17235
rect 2195 17205 2245 17235
rect 2275 17205 2325 17235
rect 2355 17205 2405 17235
rect 2435 17205 2485 17235
rect 2515 17205 2565 17235
rect 2595 17205 2645 17235
rect 2675 17205 2725 17235
rect 2755 17205 2805 17235
rect 2835 17205 2885 17235
rect 2915 17205 2965 17235
rect 2995 17205 3045 17235
rect 3075 17205 3125 17235
rect 3155 17205 3205 17235
rect 3235 17205 3285 17235
rect 3315 17205 3365 17235
rect 3395 17205 3445 17235
rect 3475 17205 3525 17235
rect 3555 17205 3605 17235
rect 3635 17205 3685 17235
rect 3715 17205 3765 17235
rect 3795 17205 3845 17235
rect 3875 17205 3925 17235
rect 3955 17205 4005 17235
rect 4035 17205 4085 17235
rect 4115 17205 4165 17235
rect 4195 17205 4725 17235
rect 4755 17205 4885 17235
rect 4915 17205 5045 17235
rect 5075 17205 5205 17235
rect 5235 17205 5365 17235
rect 5395 17205 5525 17235
rect 5555 17205 5685 17235
rect 5715 17205 6245 17235
rect 6275 17205 6325 17235
rect 6355 17205 6405 17235
rect 6435 17205 6485 17235
rect 6515 17205 6565 17235
rect 6595 17205 6645 17235
rect 6675 17205 6725 17235
rect 6755 17205 6805 17235
rect 6835 17205 6885 17235
rect 6915 17205 6965 17235
rect 6995 17205 7045 17235
rect 7075 17205 7125 17235
rect 7155 17205 7205 17235
rect 7235 17205 7285 17235
rect 7315 17205 7365 17235
rect 7395 17205 7445 17235
rect 7475 17205 7525 17235
rect 7555 17205 7605 17235
rect 7635 17205 7685 17235
rect 7715 17205 7765 17235
rect 7795 17205 7845 17235
rect 7875 17205 7925 17235
rect 7955 17205 8005 17235
rect 8035 17205 8085 17235
rect 8115 17205 8165 17235
rect 8195 17205 8245 17235
rect 8275 17205 8325 17235
rect 8355 17205 8405 17235
rect 8435 17205 8485 17235
rect 8515 17205 8565 17235
rect 8595 17205 8645 17235
rect 8675 17205 8725 17235
rect 8755 17205 8805 17235
rect 8835 17205 8885 17235
rect 8915 17205 8965 17235
rect 8995 17205 9045 17235
rect 9075 17205 9125 17235
rect 9155 17205 9205 17235
rect 9235 17205 9285 17235
rect 9315 17205 9365 17235
rect 9395 17205 9445 17235
rect 9475 17205 10005 17235
rect 10035 17205 10165 17235
rect 10195 17205 10325 17235
rect 10355 17205 10485 17235
rect 10515 17205 10645 17235
rect 10675 17205 10805 17235
rect 10835 17205 10965 17235
rect 10995 17205 11565 17235
rect 11595 17205 11645 17235
rect 11675 17205 11725 17235
rect 11755 17205 11805 17235
rect 11835 17205 11885 17235
rect 11915 17205 11965 17235
rect 11995 17205 12045 17235
rect 12075 17205 12125 17235
rect 12155 17205 12205 17235
rect 12235 17205 12285 17235
rect 12315 17205 12365 17235
rect 12395 17205 12445 17235
rect 12475 17205 12525 17235
rect 12555 17205 12605 17235
rect 12635 17205 12685 17235
rect 12715 17205 12765 17235
rect 12795 17205 12845 17235
rect 12875 17205 12925 17235
rect 12955 17205 13005 17235
rect 13035 17205 13085 17235
rect 13115 17205 13165 17235
rect 13195 17205 13245 17235
rect 13275 17205 13325 17235
rect 13355 17205 13405 17235
rect 13435 17205 13485 17235
rect 13515 17205 13565 17235
rect 13595 17205 13645 17235
rect 13675 17205 13725 17235
rect 13755 17205 13805 17235
rect 13835 17205 13885 17235
rect 13915 17205 13965 17235
rect 13995 17205 14045 17235
rect 14075 17205 14125 17235
rect 14155 17205 14205 17235
rect 14235 17205 14285 17235
rect 14315 17205 14365 17235
rect 14395 17205 14445 17235
rect 14475 17205 14525 17235
rect 14555 17205 14605 17235
rect 14635 17205 14685 17235
rect 14715 17205 15245 17235
rect 15275 17205 15405 17235
rect 15435 17205 15565 17235
rect 15595 17205 15725 17235
rect 15755 17205 15885 17235
rect 15915 17205 16045 17235
rect 16075 17205 16205 17235
rect 16235 17205 16765 17235
rect 16795 17205 16845 17235
rect 16875 17205 16925 17235
rect 16955 17205 17005 17235
rect 17035 17205 17085 17235
rect 17115 17205 17165 17235
rect 17195 17205 17245 17235
rect 17275 17205 17325 17235
rect 17355 17205 17405 17235
rect 17435 17205 17485 17235
rect 17515 17205 17565 17235
rect 17595 17205 17645 17235
rect 17675 17205 17725 17235
rect 17755 17205 17805 17235
rect 17835 17205 17885 17235
rect 17915 17205 17965 17235
rect 17995 17205 18045 17235
rect 18075 17205 18125 17235
rect 18155 17205 18205 17235
rect 18235 17205 18285 17235
rect 18315 17205 18365 17235
rect 18395 17205 18445 17235
rect 18475 17205 18525 17235
rect 18555 17205 18605 17235
rect 18635 17205 18685 17235
rect 18715 17205 18765 17235
rect 18795 17205 18845 17235
rect 18875 17205 18925 17235
rect 18955 17205 19005 17235
rect 19035 17205 19085 17235
rect 19115 17205 19165 17235
rect 19195 17205 19245 17235
rect 19275 17205 19325 17235
rect 19355 17205 19405 17235
rect 19435 17205 19485 17235
rect 19515 17205 19565 17235
rect 19595 17205 19645 17235
rect 19675 17205 19725 17235
rect 19755 17205 19805 17235
rect 19835 17205 19885 17235
rect 19915 17205 19965 17235
rect 19995 17205 20045 17235
rect 20075 17205 20125 17235
rect 20155 17205 20205 17235
rect 20235 17205 20285 17235
rect 20315 17205 20365 17235
rect 20395 17205 20445 17235
rect 20475 17205 20525 17235
rect 20555 17205 20605 17235
rect 20635 17205 20685 17235
rect 20715 17205 20765 17235
rect 20795 17205 20845 17235
rect 20875 17205 20925 17235
rect 20955 17205 20960 17235
rect 0 17200 20960 17205
rect 0 17155 20960 17160
rect 0 17125 5 17155
rect 35 17125 85 17155
rect 115 17125 165 17155
rect 195 17125 245 17155
rect 275 17125 325 17155
rect 355 17125 405 17155
rect 435 17125 485 17155
rect 515 17125 565 17155
rect 595 17125 645 17155
rect 675 17125 725 17155
rect 755 17125 805 17155
rect 835 17125 885 17155
rect 915 17125 965 17155
rect 995 17125 1045 17155
rect 1075 17125 1125 17155
rect 1155 17125 1205 17155
rect 1235 17125 1285 17155
rect 1315 17125 1365 17155
rect 1395 17125 1445 17155
rect 1475 17125 1525 17155
rect 1555 17125 1605 17155
rect 1635 17125 1685 17155
rect 1715 17125 1765 17155
rect 1795 17125 1845 17155
rect 1875 17125 1925 17155
rect 1955 17125 2005 17155
rect 2035 17125 2085 17155
rect 2115 17125 2165 17155
rect 2195 17125 2245 17155
rect 2275 17125 2325 17155
rect 2355 17125 2405 17155
rect 2435 17125 2485 17155
rect 2515 17125 2565 17155
rect 2595 17125 2645 17155
rect 2675 17125 2725 17155
rect 2755 17125 2805 17155
rect 2835 17125 2885 17155
rect 2915 17125 2965 17155
rect 2995 17125 3045 17155
rect 3075 17125 3125 17155
rect 3155 17125 3205 17155
rect 3235 17125 3285 17155
rect 3315 17125 3365 17155
rect 3395 17125 3445 17155
rect 3475 17125 3525 17155
rect 3555 17125 3605 17155
rect 3635 17125 3685 17155
rect 3715 17125 3765 17155
rect 3795 17125 3845 17155
rect 3875 17125 3925 17155
rect 3955 17125 4005 17155
rect 4035 17125 4085 17155
rect 4115 17125 4165 17155
rect 4195 17125 5765 17155
rect 5795 17125 5925 17155
rect 5955 17125 6245 17155
rect 6275 17125 6325 17155
rect 6355 17125 6405 17155
rect 6435 17125 6485 17155
rect 6515 17125 6565 17155
rect 6595 17125 6645 17155
rect 6675 17125 6725 17155
rect 6755 17125 6805 17155
rect 6835 17125 6885 17155
rect 6915 17125 6965 17155
rect 6995 17125 7045 17155
rect 7075 17125 7125 17155
rect 7155 17125 7205 17155
rect 7235 17125 7285 17155
rect 7315 17125 7365 17155
rect 7395 17125 7445 17155
rect 7475 17125 7525 17155
rect 7555 17125 7605 17155
rect 7635 17125 7685 17155
rect 7715 17125 7765 17155
rect 7795 17125 7845 17155
rect 7875 17125 7925 17155
rect 7955 17125 8005 17155
rect 8035 17125 8085 17155
rect 8115 17125 8165 17155
rect 8195 17125 8245 17155
rect 8275 17125 8325 17155
rect 8355 17125 8405 17155
rect 8435 17125 8485 17155
rect 8515 17125 8565 17155
rect 8595 17125 8645 17155
rect 8675 17125 8725 17155
rect 8755 17125 8805 17155
rect 8835 17125 8885 17155
rect 8915 17125 8965 17155
rect 8995 17125 9045 17155
rect 9075 17125 9125 17155
rect 9155 17125 9205 17155
rect 9235 17125 9285 17155
rect 9315 17125 9365 17155
rect 9395 17125 9445 17155
rect 9475 17125 9765 17155
rect 9795 17125 9925 17155
rect 9955 17125 11565 17155
rect 11595 17125 11645 17155
rect 11675 17125 11725 17155
rect 11755 17125 11805 17155
rect 11835 17125 11885 17155
rect 11915 17125 11965 17155
rect 11995 17125 12045 17155
rect 12075 17125 12125 17155
rect 12155 17125 12205 17155
rect 12235 17125 12285 17155
rect 12315 17125 12365 17155
rect 12395 17125 12445 17155
rect 12475 17125 12525 17155
rect 12555 17125 12605 17155
rect 12635 17125 12685 17155
rect 12715 17125 12765 17155
rect 12795 17125 12845 17155
rect 12875 17125 12925 17155
rect 12955 17125 13005 17155
rect 13035 17125 13085 17155
rect 13115 17125 13165 17155
rect 13195 17125 13245 17155
rect 13275 17125 13325 17155
rect 13355 17125 13405 17155
rect 13435 17125 13485 17155
rect 13515 17125 13565 17155
rect 13595 17125 13645 17155
rect 13675 17125 13725 17155
rect 13755 17125 13805 17155
rect 13835 17125 13885 17155
rect 13915 17125 13965 17155
rect 13995 17125 14045 17155
rect 14075 17125 14125 17155
rect 14155 17125 14205 17155
rect 14235 17125 14285 17155
rect 14315 17125 14365 17155
rect 14395 17125 14445 17155
rect 14475 17125 14525 17155
rect 14555 17125 14605 17155
rect 14635 17125 14685 17155
rect 14715 17125 15005 17155
rect 15035 17125 15165 17155
rect 15195 17125 16765 17155
rect 16795 17125 16845 17155
rect 16875 17125 16925 17155
rect 16955 17125 17005 17155
rect 17035 17125 17085 17155
rect 17115 17125 17165 17155
rect 17195 17125 17245 17155
rect 17275 17125 17325 17155
rect 17355 17125 17405 17155
rect 17435 17125 17485 17155
rect 17515 17125 17565 17155
rect 17595 17125 17645 17155
rect 17675 17125 17725 17155
rect 17755 17125 17805 17155
rect 17835 17125 17885 17155
rect 17915 17125 17965 17155
rect 17995 17125 18045 17155
rect 18075 17125 18125 17155
rect 18155 17125 18205 17155
rect 18235 17125 18285 17155
rect 18315 17125 18365 17155
rect 18395 17125 18445 17155
rect 18475 17125 18525 17155
rect 18555 17125 18605 17155
rect 18635 17125 18685 17155
rect 18715 17125 18765 17155
rect 18795 17125 18845 17155
rect 18875 17125 18925 17155
rect 18955 17125 19005 17155
rect 19035 17125 19085 17155
rect 19115 17125 19165 17155
rect 19195 17125 19245 17155
rect 19275 17125 19325 17155
rect 19355 17125 19405 17155
rect 19435 17125 19485 17155
rect 19515 17125 19565 17155
rect 19595 17125 19645 17155
rect 19675 17125 19725 17155
rect 19755 17125 19805 17155
rect 19835 17125 19885 17155
rect 19915 17125 19965 17155
rect 19995 17125 20045 17155
rect 20075 17125 20125 17155
rect 20155 17125 20205 17155
rect 20235 17125 20285 17155
rect 20315 17125 20365 17155
rect 20395 17125 20445 17155
rect 20475 17125 20525 17155
rect 20555 17125 20605 17155
rect 20635 17125 20685 17155
rect 20715 17125 20765 17155
rect 20795 17125 20845 17155
rect 20875 17125 20925 17155
rect 20955 17125 20960 17155
rect 0 17120 20960 17125
rect 0 17075 20960 17080
rect 0 17045 5845 17075
rect 5875 17045 9845 17075
rect 9875 17045 15085 17075
rect 15115 17045 20960 17075
rect 0 17040 20960 17045
rect 0 16995 20960 17000
rect 0 16965 5 16995
rect 35 16965 85 16995
rect 115 16965 165 16995
rect 195 16965 245 16995
rect 275 16965 325 16995
rect 355 16965 405 16995
rect 435 16965 485 16995
rect 515 16965 565 16995
rect 595 16965 645 16995
rect 675 16965 725 16995
rect 755 16965 805 16995
rect 835 16965 885 16995
rect 915 16965 965 16995
rect 995 16965 1045 16995
rect 1075 16965 1125 16995
rect 1155 16965 1205 16995
rect 1235 16965 1285 16995
rect 1315 16965 1365 16995
rect 1395 16965 1445 16995
rect 1475 16965 1525 16995
rect 1555 16965 1605 16995
rect 1635 16965 1685 16995
rect 1715 16965 1765 16995
rect 1795 16965 1845 16995
rect 1875 16965 1925 16995
rect 1955 16965 2005 16995
rect 2035 16965 2085 16995
rect 2115 16965 2165 16995
rect 2195 16965 2245 16995
rect 2275 16965 2325 16995
rect 2355 16965 2405 16995
rect 2435 16965 2485 16995
rect 2515 16965 2565 16995
rect 2595 16965 2645 16995
rect 2675 16965 2725 16995
rect 2755 16965 2805 16995
rect 2835 16965 2885 16995
rect 2915 16965 2965 16995
rect 2995 16965 3045 16995
rect 3075 16965 3125 16995
rect 3155 16965 3205 16995
rect 3235 16965 3285 16995
rect 3315 16965 3365 16995
rect 3395 16965 3445 16995
rect 3475 16965 3525 16995
rect 3555 16965 3605 16995
rect 3635 16965 3685 16995
rect 3715 16965 3765 16995
rect 3795 16965 3845 16995
rect 3875 16965 3925 16995
rect 3955 16965 4005 16995
rect 4035 16965 4085 16995
rect 4115 16965 4165 16995
rect 4195 16965 5765 16995
rect 5795 16965 5925 16995
rect 5955 16965 6245 16995
rect 6275 16965 6325 16995
rect 6355 16965 6405 16995
rect 6435 16965 6485 16995
rect 6515 16965 6565 16995
rect 6595 16965 6645 16995
rect 6675 16965 6725 16995
rect 6755 16965 6805 16995
rect 6835 16965 6885 16995
rect 6915 16965 6965 16995
rect 6995 16965 7045 16995
rect 7075 16965 7125 16995
rect 7155 16965 7205 16995
rect 7235 16965 7285 16995
rect 7315 16965 7365 16995
rect 7395 16965 7445 16995
rect 7475 16965 7525 16995
rect 7555 16965 7605 16995
rect 7635 16965 7685 16995
rect 7715 16965 7765 16995
rect 7795 16965 7845 16995
rect 7875 16965 7925 16995
rect 7955 16965 8005 16995
rect 8035 16965 8085 16995
rect 8115 16965 8165 16995
rect 8195 16965 8245 16995
rect 8275 16965 8325 16995
rect 8355 16965 8405 16995
rect 8435 16965 8485 16995
rect 8515 16965 8565 16995
rect 8595 16965 8645 16995
rect 8675 16965 8725 16995
rect 8755 16965 8805 16995
rect 8835 16965 8885 16995
rect 8915 16965 8965 16995
rect 8995 16965 9045 16995
rect 9075 16965 9125 16995
rect 9155 16965 9205 16995
rect 9235 16965 9285 16995
rect 9315 16965 9365 16995
rect 9395 16965 9445 16995
rect 9475 16965 9765 16995
rect 9795 16965 9925 16995
rect 9955 16965 11565 16995
rect 11595 16965 11645 16995
rect 11675 16965 11725 16995
rect 11755 16965 11805 16995
rect 11835 16965 11885 16995
rect 11915 16965 11965 16995
rect 11995 16965 12045 16995
rect 12075 16965 12125 16995
rect 12155 16965 12205 16995
rect 12235 16965 12285 16995
rect 12315 16965 12365 16995
rect 12395 16965 12445 16995
rect 12475 16965 12525 16995
rect 12555 16965 12605 16995
rect 12635 16965 12685 16995
rect 12715 16965 12765 16995
rect 12795 16965 12845 16995
rect 12875 16965 12925 16995
rect 12955 16965 13005 16995
rect 13035 16965 13085 16995
rect 13115 16965 13165 16995
rect 13195 16965 13245 16995
rect 13275 16965 13325 16995
rect 13355 16965 13405 16995
rect 13435 16965 13485 16995
rect 13515 16965 13565 16995
rect 13595 16965 13645 16995
rect 13675 16965 13725 16995
rect 13755 16965 13805 16995
rect 13835 16965 13885 16995
rect 13915 16965 13965 16995
rect 13995 16965 14045 16995
rect 14075 16965 14125 16995
rect 14155 16965 14205 16995
rect 14235 16965 14285 16995
rect 14315 16965 14365 16995
rect 14395 16965 14445 16995
rect 14475 16965 14525 16995
rect 14555 16965 14605 16995
rect 14635 16965 14685 16995
rect 14715 16965 15005 16995
rect 15035 16965 15165 16995
rect 15195 16965 16765 16995
rect 16795 16965 16845 16995
rect 16875 16965 16925 16995
rect 16955 16965 17005 16995
rect 17035 16965 17085 16995
rect 17115 16965 17165 16995
rect 17195 16965 17245 16995
rect 17275 16965 17325 16995
rect 17355 16965 17405 16995
rect 17435 16965 17485 16995
rect 17515 16965 17565 16995
rect 17595 16965 17645 16995
rect 17675 16965 17725 16995
rect 17755 16965 17805 16995
rect 17835 16965 17885 16995
rect 17915 16965 17965 16995
rect 17995 16965 18045 16995
rect 18075 16965 18125 16995
rect 18155 16965 18205 16995
rect 18235 16965 18285 16995
rect 18315 16965 18365 16995
rect 18395 16965 18445 16995
rect 18475 16965 18525 16995
rect 18555 16965 18605 16995
rect 18635 16965 18685 16995
rect 18715 16965 18765 16995
rect 18795 16965 18845 16995
rect 18875 16965 18925 16995
rect 18955 16965 19005 16995
rect 19035 16965 19085 16995
rect 19115 16965 19165 16995
rect 19195 16965 19245 16995
rect 19275 16965 19325 16995
rect 19355 16965 19405 16995
rect 19435 16965 19485 16995
rect 19515 16965 19565 16995
rect 19595 16965 19645 16995
rect 19675 16965 19725 16995
rect 19755 16965 19805 16995
rect 19835 16965 19885 16995
rect 19915 16965 19965 16995
rect 19995 16965 20045 16995
rect 20075 16965 20125 16995
rect 20155 16965 20205 16995
rect 20235 16965 20285 16995
rect 20315 16965 20365 16995
rect 20395 16965 20445 16995
rect 20475 16965 20525 16995
rect 20555 16965 20605 16995
rect 20635 16965 20685 16995
rect 20715 16965 20765 16995
rect 20795 16965 20845 16995
rect 20875 16965 20925 16995
rect 20955 16965 20960 16995
rect 0 16960 20960 16965
rect 0 16915 20960 16920
rect 0 16885 5 16915
rect 35 16885 85 16915
rect 115 16885 165 16915
rect 195 16885 245 16915
rect 275 16885 325 16915
rect 355 16885 405 16915
rect 435 16885 485 16915
rect 515 16885 565 16915
rect 595 16885 645 16915
rect 675 16885 725 16915
rect 755 16885 805 16915
rect 835 16885 885 16915
rect 915 16885 965 16915
rect 995 16885 1045 16915
rect 1075 16885 1125 16915
rect 1155 16885 1205 16915
rect 1235 16885 1285 16915
rect 1315 16885 1365 16915
rect 1395 16885 1445 16915
rect 1475 16885 1525 16915
rect 1555 16885 1605 16915
rect 1635 16885 1685 16915
rect 1715 16885 1765 16915
rect 1795 16885 1845 16915
rect 1875 16885 1925 16915
rect 1955 16885 2005 16915
rect 2035 16885 2085 16915
rect 2115 16885 2165 16915
rect 2195 16885 2245 16915
rect 2275 16885 2325 16915
rect 2355 16885 2405 16915
rect 2435 16885 2485 16915
rect 2515 16885 2565 16915
rect 2595 16885 2645 16915
rect 2675 16885 2725 16915
rect 2755 16885 2805 16915
rect 2835 16885 2885 16915
rect 2915 16885 2965 16915
rect 2995 16885 3045 16915
rect 3075 16885 3125 16915
rect 3155 16885 3205 16915
rect 3235 16885 3285 16915
rect 3315 16885 3365 16915
rect 3395 16885 3445 16915
rect 3475 16885 3525 16915
rect 3555 16885 3605 16915
rect 3635 16885 3685 16915
rect 3715 16885 3765 16915
rect 3795 16885 3845 16915
rect 3875 16885 3925 16915
rect 3955 16885 4005 16915
rect 4035 16885 4085 16915
rect 4115 16885 4165 16915
rect 4195 16885 6005 16915
rect 6035 16885 6165 16915
rect 6195 16885 6245 16915
rect 6275 16885 6325 16915
rect 6355 16885 6405 16915
rect 6435 16885 6485 16915
rect 6515 16885 6565 16915
rect 6595 16885 6645 16915
rect 6675 16885 6725 16915
rect 6755 16885 6805 16915
rect 6835 16885 6885 16915
rect 6915 16885 6965 16915
rect 6995 16885 7045 16915
rect 7075 16885 7125 16915
rect 7155 16885 7205 16915
rect 7235 16885 7285 16915
rect 7315 16885 7365 16915
rect 7395 16885 7445 16915
rect 7475 16885 7525 16915
rect 7555 16885 7605 16915
rect 7635 16885 7685 16915
rect 7715 16885 7765 16915
rect 7795 16885 7845 16915
rect 7875 16885 7925 16915
rect 7955 16885 8005 16915
rect 8035 16885 8085 16915
rect 8115 16885 8165 16915
rect 8195 16885 8245 16915
rect 8275 16885 8325 16915
rect 8355 16885 8405 16915
rect 8435 16885 8485 16915
rect 8515 16885 8565 16915
rect 8595 16885 8645 16915
rect 8675 16885 8725 16915
rect 8755 16885 8805 16915
rect 8835 16885 8885 16915
rect 8915 16885 8965 16915
rect 8995 16885 9045 16915
rect 9075 16885 9125 16915
rect 9155 16885 9205 16915
rect 9235 16885 9285 16915
rect 9315 16885 9365 16915
rect 9395 16885 9445 16915
rect 9475 16885 9525 16915
rect 9555 16885 9685 16915
rect 9715 16885 11565 16915
rect 11595 16885 11645 16915
rect 11675 16885 11725 16915
rect 11755 16885 11805 16915
rect 11835 16885 11885 16915
rect 11915 16885 11965 16915
rect 11995 16885 12045 16915
rect 12075 16885 12125 16915
rect 12155 16885 12205 16915
rect 12235 16885 12285 16915
rect 12315 16885 12365 16915
rect 12395 16885 12445 16915
rect 12475 16885 12525 16915
rect 12555 16885 12605 16915
rect 12635 16885 12685 16915
rect 12715 16885 12765 16915
rect 12795 16885 12845 16915
rect 12875 16885 12925 16915
rect 12955 16885 13005 16915
rect 13035 16885 13085 16915
rect 13115 16885 13165 16915
rect 13195 16885 13245 16915
rect 13275 16885 13325 16915
rect 13355 16885 13405 16915
rect 13435 16885 13485 16915
rect 13515 16885 13565 16915
rect 13595 16885 13645 16915
rect 13675 16885 13725 16915
rect 13755 16885 13805 16915
rect 13835 16885 13885 16915
rect 13915 16885 13965 16915
rect 13995 16885 14045 16915
rect 14075 16885 14125 16915
rect 14155 16885 14205 16915
rect 14235 16885 14285 16915
rect 14315 16885 14365 16915
rect 14395 16885 14445 16915
rect 14475 16885 14525 16915
rect 14555 16885 14605 16915
rect 14635 16885 14685 16915
rect 14715 16885 14765 16915
rect 14795 16885 14925 16915
rect 14955 16885 16765 16915
rect 16795 16885 16845 16915
rect 16875 16885 16925 16915
rect 16955 16885 17005 16915
rect 17035 16885 17085 16915
rect 17115 16885 17165 16915
rect 17195 16885 17245 16915
rect 17275 16885 17325 16915
rect 17355 16885 17405 16915
rect 17435 16885 17485 16915
rect 17515 16885 17565 16915
rect 17595 16885 17645 16915
rect 17675 16885 17725 16915
rect 17755 16885 17805 16915
rect 17835 16885 17885 16915
rect 17915 16885 17965 16915
rect 17995 16885 18045 16915
rect 18075 16885 18125 16915
rect 18155 16885 18205 16915
rect 18235 16885 18285 16915
rect 18315 16885 18365 16915
rect 18395 16885 18445 16915
rect 18475 16885 18525 16915
rect 18555 16885 18605 16915
rect 18635 16885 18685 16915
rect 18715 16885 18765 16915
rect 18795 16885 18845 16915
rect 18875 16885 18925 16915
rect 18955 16885 19005 16915
rect 19035 16885 19085 16915
rect 19115 16885 19165 16915
rect 19195 16885 19245 16915
rect 19275 16885 19325 16915
rect 19355 16885 19405 16915
rect 19435 16885 19485 16915
rect 19515 16885 19565 16915
rect 19595 16885 19645 16915
rect 19675 16885 19725 16915
rect 19755 16885 19805 16915
rect 19835 16885 19885 16915
rect 19915 16885 19965 16915
rect 19995 16885 20045 16915
rect 20075 16885 20125 16915
rect 20155 16885 20205 16915
rect 20235 16885 20285 16915
rect 20315 16885 20365 16915
rect 20395 16885 20445 16915
rect 20475 16885 20525 16915
rect 20555 16885 20605 16915
rect 20635 16885 20685 16915
rect 20715 16885 20765 16915
rect 20795 16885 20845 16915
rect 20875 16885 20925 16915
rect 20955 16885 20960 16915
rect 0 16880 20960 16885
rect 0 16835 20960 16840
rect 0 16805 6085 16835
rect 6115 16805 9605 16835
rect 9635 16805 14845 16835
rect 14875 16805 20960 16835
rect 0 16800 20960 16805
rect 0 16755 20960 16760
rect 0 16725 5 16755
rect 35 16725 85 16755
rect 115 16725 165 16755
rect 195 16725 245 16755
rect 275 16725 325 16755
rect 355 16725 405 16755
rect 435 16725 485 16755
rect 515 16725 565 16755
rect 595 16725 645 16755
rect 675 16725 725 16755
rect 755 16725 805 16755
rect 835 16725 885 16755
rect 915 16725 965 16755
rect 995 16725 1045 16755
rect 1075 16725 1125 16755
rect 1155 16725 1205 16755
rect 1235 16725 1285 16755
rect 1315 16725 1365 16755
rect 1395 16725 1445 16755
rect 1475 16725 1525 16755
rect 1555 16725 1605 16755
rect 1635 16725 1685 16755
rect 1715 16725 1765 16755
rect 1795 16725 1845 16755
rect 1875 16725 1925 16755
rect 1955 16725 2005 16755
rect 2035 16725 2085 16755
rect 2115 16725 2165 16755
rect 2195 16725 2245 16755
rect 2275 16725 2325 16755
rect 2355 16725 2405 16755
rect 2435 16725 2485 16755
rect 2515 16725 2565 16755
rect 2595 16725 2645 16755
rect 2675 16725 2725 16755
rect 2755 16725 2805 16755
rect 2835 16725 2885 16755
rect 2915 16725 2965 16755
rect 2995 16725 3045 16755
rect 3075 16725 3125 16755
rect 3155 16725 3205 16755
rect 3235 16725 3285 16755
rect 3315 16725 3365 16755
rect 3395 16725 3445 16755
rect 3475 16725 3525 16755
rect 3555 16725 3605 16755
rect 3635 16725 3685 16755
rect 3715 16725 3765 16755
rect 3795 16725 3845 16755
rect 3875 16725 3925 16755
rect 3955 16725 4005 16755
rect 4035 16725 4085 16755
rect 4115 16725 4165 16755
rect 4195 16725 6005 16755
rect 6035 16725 6165 16755
rect 6195 16725 6245 16755
rect 6275 16725 6325 16755
rect 6355 16725 6405 16755
rect 6435 16725 6485 16755
rect 6515 16725 6565 16755
rect 6595 16725 6645 16755
rect 6675 16725 6725 16755
rect 6755 16725 6805 16755
rect 6835 16725 6885 16755
rect 6915 16725 6965 16755
rect 6995 16725 7045 16755
rect 7075 16725 7125 16755
rect 7155 16725 7205 16755
rect 7235 16725 7285 16755
rect 7315 16725 7365 16755
rect 7395 16725 7445 16755
rect 7475 16725 7525 16755
rect 7555 16725 7605 16755
rect 7635 16725 7685 16755
rect 7715 16725 7765 16755
rect 7795 16725 7845 16755
rect 7875 16725 7925 16755
rect 7955 16725 8005 16755
rect 8035 16725 8085 16755
rect 8115 16725 8165 16755
rect 8195 16725 8245 16755
rect 8275 16725 8325 16755
rect 8355 16725 8405 16755
rect 8435 16725 8485 16755
rect 8515 16725 8565 16755
rect 8595 16725 8645 16755
rect 8675 16725 8725 16755
rect 8755 16725 8805 16755
rect 8835 16725 8885 16755
rect 8915 16725 8965 16755
rect 8995 16725 9045 16755
rect 9075 16725 9125 16755
rect 9155 16725 9205 16755
rect 9235 16725 9285 16755
rect 9315 16725 9365 16755
rect 9395 16725 9445 16755
rect 9475 16725 9525 16755
rect 9555 16725 9685 16755
rect 9715 16725 11565 16755
rect 11595 16725 11645 16755
rect 11675 16725 11725 16755
rect 11755 16725 11805 16755
rect 11835 16725 11885 16755
rect 11915 16725 11965 16755
rect 11995 16725 12045 16755
rect 12075 16725 12125 16755
rect 12155 16725 12205 16755
rect 12235 16725 12285 16755
rect 12315 16725 12365 16755
rect 12395 16725 12445 16755
rect 12475 16725 12525 16755
rect 12555 16725 12605 16755
rect 12635 16725 12685 16755
rect 12715 16725 12765 16755
rect 12795 16725 12845 16755
rect 12875 16725 12925 16755
rect 12955 16725 13005 16755
rect 13035 16725 13085 16755
rect 13115 16725 13165 16755
rect 13195 16725 13245 16755
rect 13275 16725 13325 16755
rect 13355 16725 13405 16755
rect 13435 16725 13485 16755
rect 13515 16725 13565 16755
rect 13595 16725 13645 16755
rect 13675 16725 13725 16755
rect 13755 16725 13805 16755
rect 13835 16725 13885 16755
rect 13915 16725 13965 16755
rect 13995 16725 14045 16755
rect 14075 16725 14125 16755
rect 14155 16725 14205 16755
rect 14235 16725 14285 16755
rect 14315 16725 14365 16755
rect 14395 16725 14445 16755
rect 14475 16725 14525 16755
rect 14555 16725 14605 16755
rect 14635 16725 14685 16755
rect 14715 16725 14765 16755
rect 14795 16725 14925 16755
rect 14955 16725 16765 16755
rect 16795 16725 16845 16755
rect 16875 16725 16925 16755
rect 16955 16725 17005 16755
rect 17035 16725 17085 16755
rect 17115 16725 17165 16755
rect 17195 16725 17245 16755
rect 17275 16725 17325 16755
rect 17355 16725 17405 16755
rect 17435 16725 17485 16755
rect 17515 16725 17565 16755
rect 17595 16725 17645 16755
rect 17675 16725 17725 16755
rect 17755 16725 17805 16755
rect 17835 16725 17885 16755
rect 17915 16725 17965 16755
rect 17995 16725 18045 16755
rect 18075 16725 18125 16755
rect 18155 16725 18205 16755
rect 18235 16725 18285 16755
rect 18315 16725 18365 16755
rect 18395 16725 18445 16755
rect 18475 16725 18525 16755
rect 18555 16725 18605 16755
rect 18635 16725 18685 16755
rect 18715 16725 18765 16755
rect 18795 16725 18845 16755
rect 18875 16725 18925 16755
rect 18955 16725 19005 16755
rect 19035 16725 19085 16755
rect 19115 16725 19165 16755
rect 19195 16725 19245 16755
rect 19275 16725 19325 16755
rect 19355 16725 19405 16755
rect 19435 16725 19485 16755
rect 19515 16725 19565 16755
rect 19595 16725 19645 16755
rect 19675 16725 19725 16755
rect 19755 16725 19805 16755
rect 19835 16725 19885 16755
rect 19915 16725 19965 16755
rect 19995 16725 20045 16755
rect 20075 16725 20125 16755
rect 20155 16725 20205 16755
rect 20235 16725 20285 16755
rect 20315 16725 20365 16755
rect 20395 16725 20445 16755
rect 20475 16725 20525 16755
rect 20555 16725 20605 16755
rect 20635 16725 20685 16755
rect 20715 16725 20765 16755
rect 20795 16725 20845 16755
rect 20875 16725 20925 16755
rect 20955 16725 20960 16755
rect 0 16720 20960 16725
rect 0 16675 20960 16680
rect 0 16645 5 16675
rect 35 16645 85 16675
rect 115 16645 165 16675
rect 195 16645 245 16675
rect 275 16645 325 16675
rect 355 16645 405 16675
rect 435 16645 485 16675
rect 515 16645 565 16675
rect 595 16645 645 16675
rect 675 16645 725 16675
rect 755 16645 805 16675
rect 835 16645 885 16675
rect 915 16645 965 16675
rect 995 16645 1045 16675
rect 1075 16645 1125 16675
rect 1155 16645 1205 16675
rect 1235 16645 1285 16675
rect 1315 16645 1365 16675
rect 1395 16645 1445 16675
rect 1475 16645 1525 16675
rect 1555 16645 1605 16675
rect 1635 16645 1685 16675
rect 1715 16645 1765 16675
rect 1795 16645 1845 16675
rect 1875 16645 1925 16675
rect 1955 16645 2005 16675
rect 2035 16645 2085 16675
rect 2115 16645 2165 16675
rect 2195 16645 2245 16675
rect 2275 16645 2325 16675
rect 2355 16645 2405 16675
rect 2435 16645 2485 16675
rect 2515 16645 2565 16675
rect 2595 16645 2645 16675
rect 2675 16645 2725 16675
rect 2755 16645 2805 16675
rect 2835 16645 2885 16675
rect 2915 16645 2965 16675
rect 2995 16645 3045 16675
rect 3075 16645 3125 16675
rect 3155 16645 3205 16675
rect 3235 16645 3285 16675
rect 3315 16645 3365 16675
rect 3395 16645 3445 16675
rect 3475 16645 3525 16675
rect 3555 16645 3605 16675
rect 3635 16645 3685 16675
rect 3715 16645 3765 16675
rect 3795 16645 3845 16675
rect 3875 16645 3925 16675
rect 3955 16645 4005 16675
rect 4035 16645 4085 16675
rect 4115 16645 4165 16675
rect 4195 16645 4245 16675
rect 4275 16645 4405 16675
rect 4435 16645 6245 16675
rect 6275 16645 6325 16675
rect 6355 16645 6405 16675
rect 6435 16645 6485 16675
rect 6515 16645 6565 16675
rect 6595 16645 6645 16675
rect 6675 16645 6725 16675
rect 6755 16645 6805 16675
rect 6835 16645 6885 16675
rect 6915 16645 6965 16675
rect 6995 16645 7045 16675
rect 7075 16645 7125 16675
rect 7155 16645 7205 16675
rect 7235 16645 7285 16675
rect 7315 16645 7365 16675
rect 7395 16645 7445 16675
rect 7475 16645 7525 16675
rect 7555 16645 7605 16675
rect 7635 16645 7685 16675
rect 7715 16645 7765 16675
rect 7795 16645 7845 16675
rect 7875 16645 7925 16675
rect 7955 16645 8005 16675
rect 8035 16645 8085 16675
rect 8115 16645 8165 16675
rect 8195 16645 8245 16675
rect 8275 16645 8325 16675
rect 8355 16645 8405 16675
rect 8435 16645 8485 16675
rect 8515 16645 8565 16675
rect 8595 16645 8645 16675
rect 8675 16645 8725 16675
rect 8755 16645 8805 16675
rect 8835 16645 8885 16675
rect 8915 16645 8965 16675
rect 8995 16645 9045 16675
rect 9075 16645 9125 16675
rect 9155 16645 9205 16675
rect 9235 16645 9285 16675
rect 9315 16645 9365 16675
rect 9395 16645 9445 16675
rect 9475 16645 9525 16675
rect 9555 16645 9685 16675
rect 9715 16645 11565 16675
rect 11595 16645 11645 16675
rect 11675 16645 11725 16675
rect 11755 16645 11805 16675
rect 11835 16645 11885 16675
rect 11915 16645 11965 16675
rect 11995 16645 12045 16675
rect 12075 16645 12125 16675
rect 12155 16645 12205 16675
rect 12235 16645 12285 16675
rect 12315 16645 12365 16675
rect 12395 16645 12445 16675
rect 12475 16645 12525 16675
rect 12555 16645 12605 16675
rect 12635 16645 12685 16675
rect 12715 16645 12765 16675
rect 12795 16645 12845 16675
rect 12875 16645 12925 16675
rect 12955 16645 13005 16675
rect 13035 16645 13085 16675
rect 13115 16645 13165 16675
rect 13195 16645 13245 16675
rect 13275 16645 13325 16675
rect 13355 16645 13405 16675
rect 13435 16645 13485 16675
rect 13515 16645 13565 16675
rect 13595 16645 13645 16675
rect 13675 16645 13725 16675
rect 13755 16645 13805 16675
rect 13835 16645 13885 16675
rect 13915 16645 13965 16675
rect 13995 16645 14045 16675
rect 14075 16645 14125 16675
rect 14155 16645 14205 16675
rect 14235 16645 14285 16675
rect 14315 16645 14365 16675
rect 14395 16645 14445 16675
rect 14475 16645 14525 16675
rect 14555 16645 14605 16675
rect 14635 16645 14685 16675
rect 14715 16645 16525 16675
rect 16555 16645 16685 16675
rect 16715 16645 16765 16675
rect 16795 16645 16845 16675
rect 16875 16645 16925 16675
rect 16955 16645 17005 16675
rect 17035 16645 17085 16675
rect 17115 16645 17165 16675
rect 17195 16645 17245 16675
rect 17275 16645 17325 16675
rect 17355 16645 17405 16675
rect 17435 16645 17485 16675
rect 17515 16645 17565 16675
rect 17595 16645 17645 16675
rect 17675 16645 17725 16675
rect 17755 16645 17805 16675
rect 17835 16645 17885 16675
rect 17915 16645 17965 16675
rect 17995 16645 18045 16675
rect 18075 16645 18125 16675
rect 18155 16645 18205 16675
rect 18235 16645 18285 16675
rect 18315 16645 18365 16675
rect 18395 16645 18445 16675
rect 18475 16645 18525 16675
rect 18555 16645 18605 16675
rect 18635 16645 18685 16675
rect 18715 16645 18765 16675
rect 18795 16645 18845 16675
rect 18875 16645 18925 16675
rect 18955 16645 19005 16675
rect 19035 16645 19085 16675
rect 19115 16645 19165 16675
rect 19195 16645 19245 16675
rect 19275 16645 19325 16675
rect 19355 16645 19405 16675
rect 19435 16645 19485 16675
rect 19515 16645 19565 16675
rect 19595 16645 19645 16675
rect 19675 16645 19725 16675
rect 19755 16645 19805 16675
rect 19835 16645 19885 16675
rect 19915 16645 19965 16675
rect 19995 16645 20045 16675
rect 20075 16645 20125 16675
rect 20155 16645 20205 16675
rect 20235 16645 20285 16675
rect 20315 16645 20365 16675
rect 20395 16645 20445 16675
rect 20475 16645 20525 16675
rect 20555 16645 20605 16675
rect 20635 16645 20685 16675
rect 20715 16645 20765 16675
rect 20795 16645 20845 16675
rect 20875 16645 20925 16675
rect 20955 16645 20960 16675
rect 0 16640 20960 16645
rect 0 16595 20960 16600
rect 0 16565 4325 16595
rect 4355 16565 9605 16595
rect 9635 16565 16605 16595
rect 16635 16565 20960 16595
rect 0 16560 20960 16565
rect 0 16515 20960 16520
rect 0 16485 5 16515
rect 35 16485 85 16515
rect 115 16485 165 16515
rect 195 16485 245 16515
rect 275 16485 325 16515
rect 355 16485 405 16515
rect 435 16485 485 16515
rect 515 16485 565 16515
rect 595 16485 645 16515
rect 675 16485 725 16515
rect 755 16485 805 16515
rect 835 16485 885 16515
rect 915 16485 965 16515
rect 995 16485 1045 16515
rect 1075 16485 1125 16515
rect 1155 16485 1205 16515
rect 1235 16485 1285 16515
rect 1315 16485 1365 16515
rect 1395 16485 1445 16515
rect 1475 16485 1525 16515
rect 1555 16485 1605 16515
rect 1635 16485 1685 16515
rect 1715 16485 1765 16515
rect 1795 16485 1845 16515
rect 1875 16485 1925 16515
rect 1955 16485 2005 16515
rect 2035 16485 2085 16515
rect 2115 16485 2165 16515
rect 2195 16485 2245 16515
rect 2275 16485 2325 16515
rect 2355 16485 2405 16515
rect 2435 16485 2485 16515
rect 2515 16485 2565 16515
rect 2595 16485 2645 16515
rect 2675 16485 2725 16515
rect 2755 16485 2805 16515
rect 2835 16485 2885 16515
rect 2915 16485 2965 16515
rect 2995 16485 3045 16515
rect 3075 16485 3125 16515
rect 3155 16485 3205 16515
rect 3235 16485 3285 16515
rect 3315 16485 3365 16515
rect 3395 16485 3445 16515
rect 3475 16485 3525 16515
rect 3555 16485 3605 16515
rect 3635 16485 3685 16515
rect 3715 16485 3765 16515
rect 3795 16485 3845 16515
rect 3875 16485 3925 16515
rect 3955 16485 4005 16515
rect 4035 16485 4085 16515
rect 4115 16485 4165 16515
rect 4195 16485 4245 16515
rect 4275 16485 4405 16515
rect 4435 16485 6245 16515
rect 6275 16485 6325 16515
rect 6355 16485 6405 16515
rect 6435 16485 6485 16515
rect 6515 16485 6565 16515
rect 6595 16485 6645 16515
rect 6675 16485 6725 16515
rect 6755 16485 6805 16515
rect 6835 16485 6885 16515
rect 6915 16485 6965 16515
rect 6995 16485 7045 16515
rect 7075 16485 7125 16515
rect 7155 16485 7205 16515
rect 7235 16485 7285 16515
rect 7315 16485 7365 16515
rect 7395 16485 7445 16515
rect 7475 16485 7525 16515
rect 7555 16485 7605 16515
rect 7635 16485 7685 16515
rect 7715 16485 7765 16515
rect 7795 16485 7845 16515
rect 7875 16485 7925 16515
rect 7955 16485 8005 16515
rect 8035 16485 8085 16515
rect 8115 16485 8165 16515
rect 8195 16485 8245 16515
rect 8275 16485 8325 16515
rect 8355 16485 8405 16515
rect 8435 16485 8485 16515
rect 8515 16485 8565 16515
rect 8595 16485 8645 16515
rect 8675 16485 8725 16515
rect 8755 16485 8805 16515
rect 8835 16485 8885 16515
rect 8915 16485 8965 16515
rect 8995 16485 9045 16515
rect 9075 16485 9125 16515
rect 9155 16485 9205 16515
rect 9235 16485 9285 16515
rect 9315 16485 9365 16515
rect 9395 16485 9445 16515
rect 9475 16485 9525 16515
rect 9555 16485 9685 16515
rect 9715 16485 11565 16515
rect 11595 16485 11645 16515
rect 11675 16485 11725 16515
rect 11755 16485 11805 16515
rect 11835 16485 11885 16515
rect 11915 16485 11965 16515
rect 11995 16485 12045 16515
rect 12075 16485 12125 16515
rect 12155 16485 12205 16515
rect 12235 16485 12285 16515
rect 12315 16485 12365 16515
rect 12395 16485 12445 16515
rect 12475 16485 12525 16515
rect 12555 16485 12605 16515
rect 12635 16485 12685 16515
rect 12715 16485 12765 16515
rect 12795 16485 12845 16515
rect 12875 16485 12925 16515
rect 12955 16485 13005 16515
rect 13035 16485 13085 16515
rect 13115 16485 13165 16515
rect 13195 16485 13245 16515
rect 13275 16485 13325 16515
rect 13355 16485 13405 16515
rect 13435 16485 13485 16515
rect 13515 16485 13565 16515
rect 13595 16485 13645 16515
rect 13675 16485 13725 16515
rect 13755 16485 13805 16515
rect 13835 16485 13885 16515
rect 13915 16485 13965 16515
rect 13995 16485 14045 16515
rect 14075 16485 14125 16515
rect 14155 16485 14205 16515
rect 14235 16485 14285 16515
rect 14315 16485 14365 16515
rect 14395 16485 14445 16515
rect 14475 16485 14525 16515
rect 14555 16485 14605 16515
rect 14635 16485 14685 16515
rect 14715 16485 16525 16515
rect 16555 16485 16685 16515
rect 16715 16485 16765 16515
rect 16795 16485 16845 16515
rect 16875 16485 16925 16515
rect 16955 16485 17005 16515
rect 17035 16485 17085 16515
rect 17115 16485 17165 16515
rect 17195 16485 17245 16515
rect 17275 16485 17325 16515
rect 17355 16485 17405 16515
rect 17435 16485 17485 16515
rect 17515 16485 17565 16515
rect 17595 16485 17645 16515
rect 17675 16485 17725 16515
rect 17755 16485 17805 16515
rect 17835 16485 17885 16515
rect 17915 16485 17965 16515
rect 17995 16485 18045 16515
rect 18075 16485 18125 16515
rect 18155 16485 18205 16515
rect 18235 16485 18285 16515
rect 18315 16485 18365 16515
rect 18395 16485 18445 16515
rect 18475 16485 18525 16515
rect 18555 16485 18605 16515
rect 18635 16485 18685 16515
rect 18715 16485 18765 16515
rect 18795 16485 18845 16515
rect 18875 16485 18925 16515
rect 18955 16485 19005 16515
rect 19035 16485 19085 16515
rect 19115 16485 19165 16515
rect 19195 16485 19245 16515
rect 19275 16485 19325 16515
rect 19355 16485 19405 16515
rect 19435 16485 19485 16515
rect 19515 16485 19565 16515
rect 19595 16485 19645 16515
rect 19675 16485 19725 16515
rect 19755 16485 19805 16515
rect 19835 16485 19885 16515
rect 19915 16485 19965 16515
rect 19995 16485 20045 16515
rect 20075 16485 20125 16515
rect 20155 16485 20205 16515
rect 20235 16485 20285 16515
rect 20315 16485 20365 16515
rect 20395 16485 20445 16515
rect 20475 16485 20525 16515
rect 20555 16485 20605 16515
rect 20635 16485 20685 16515
rect 20715 16485 20765 16515
rect 20795 16485 20845 16515
rect 20875 16485 20925 16515
rect 20955 16485 20960 16515
rect 0 16480 20960 16485
rect 0 16435 20960 16440
rect 0 16405 5 16435
rect 35 16405 85 16435
rect 115 16405 165 16435
rect 195 16405 245 16435
rect 275 16405 325 16435
rect 355 16405 405 16435
rect 435 16405 485 16435
rect 515 16405 565 16435
rect 595 16405 645 16435
rect 675 16405 725 16435
rect 755 16405 805 16435
rect 835 16405 885 16435
rect 915 16405 965 16435
rect 995 16405 1045 16435
rect 1075 16405 1125 16435
rect 1155 16405 1205 16435
rect 1235 16405 1285 16435
rect 1315 16405 1365 16435
rect 1395 16405 1445 16435
rect 1475 16405 1525 16435
rect 1555 16405 1605 16435
rect 1635 16405 1685 16435
rect 1715 16405 1765 16435
rect 1795 16405 1845 16435
rect 1875 16405 1925 16435
rect 1955 16405 2005 16435
rect 2035 16405 2085 16435
rect 2115 16405 2165 16435
rect 2195 16405 2245 16435
rect 2275 16405 2325 16435
rect 2355 16405 2405 16435
rect 2435 16405 2485 16435
rect 2515 16405 2565 16435
rect 2595 16405 2645 16435
rect 2675 16405 2725 16435
rect 2755 16405 2805 16435
rect 2835 16405 2885 16435
rect 2915 16405 2965 16435
rect 2995 16405 3045 16435
rect 3075 16405 3125 16435
rect 3155 16405 3205 16435
rect 3235 16405 3285 16435
rect 3315 16405 3365 16435
rect 3395 16405 3445 16435
rect 3475 16405 3525 16435
rect 3555 16405 3605 16435
rect 3635 16405 3685 16435
rect 3715 16405 3765 16435
rect 3795 16405 3845 16435
rect 3875 16405 3925 16435
rect 3955 16405 4005 16435
rect 4035 16405 4085 16435
rect 4115 16405 4165 16435
rect 4195 16405 4485 16435
rect 4515 16405 4645 16435
rect 4675 16405 6245 16435
rect 6275 16405 6325 16435
rect 6355 16405 6405 16435
rect 6435 16405 6485 16435
rect 6515 16405 6565 16435
rect 6595 16405 6645 16435
rect 6675 16405 6725 16435
rect 6755 16405 6805 16435
rect 6835 16405 6885 16435
rect 6915 16405 6965 16435
rect 6995 16405 7045 16435
rect 7075 16405 7125 16435
rect 7155 16405 7205 16435
rect 7235 16405 7285 16435
rect 7315 16405 7365 16435
rect 7395 16405 7445 16435
rect 7475 16405 7525 16435
rect 7555 16405 7605 16435
rect 7635 16405 7685 16435
rect 7715 16405 7765 16435
rect 7795 16405 7845 16435
rect 7875 16405 7925 16435
rect 7955 16405 8005 16435
rect 8035 16405 8085 16435
rect 8115 16405 8165 16435
rect 8195 16405 8245 16435
rect 8275 16405 8325 16435
rect 8355 16405 8405 16435
rect 8435 16405 8485 16435
rect 8515 16405 8565 16435
rect 8595 16405 8645 16435
rect 8675 16405 8725 16435
rect 8755 16405 8805 16435
rect 8835 16405 8885 16435
rect 8915 16405 8965 16435
rect 8995 16405 9045 16435
rect 9075 16405 9125 16435
rect 9155 16405 9205 16435
rect 9235 16405 9285 16435
rect 9315 16405 9365 16435
rect 9395 16405 9445 16435
rect 9475 16405 9765 16435
rect 9795 16405 9925 16435
rect 9955 16405 11565 16435
rect 11595 16405 11645 16435
rect 11675 16405 11725 16435
rect 11755 16405 11805 16435
rect 11835 16405 11885 16435
rect 11915 16405 11965 16435
rect 11995 16405 12045 16435
rect 12075 16405 12125 16435
rect 12155 16405 12205 16435
rect 12235 16405 12285 16435
rect 12315 16405 12365 16435
rect 12395 16405 12445 16435
rect 12475 16405 12525 16435
rect 12555 16405 12605 16435
rect 12635 16405 12685 16435
rect 12715 16405 12765 16435
rect 12795 16405 12845 16435
rect 12875 16405 12925 16435
rect 12955 16405 13005 16435
rect 13035 16405 13085 16435
rect 13115 16405 13165 16435
rect 13195 16405 13245 16435
rect 13275 16405 13325 16435
rect 13355 16405 13405 16435
rect 13435 16405 13485 16435
rect 13515 16405 13565 16435
rect 13595 16405 13645 16435
rect 13675 16405 13725 16435
rect 13755 16405 13805 16435
rect 13835 16405 13885 16435
rect 13915 16405 13965 16435
rect 13995 16405 14045 16435
rect 14075 16405 14125 16435
rect 14155 16405 14205 16435
rect 14235 16405 14285 16435
rect 14315 16405 14365 16435
rect 14395 16405 14445 16435
rect 14475 16405 14525 16435
rect 14555 16405 14605 16435
rect 14635 16405 14685 16435
rect 14715 16405 16285 16435
rect 16315 16405 16445 16435
rect 16475 16405 16765 16435
rect 16795 16405 16845 16435
rect 16875 16405 16925 16435
rect 16955 16405 17005 16435
rect 17035 16405 17085 16435
rect 17115 16405 17165 16435
rect 17195 16405 17245 16435
rect 17275 16405 17325 16435
rect 17355 16405 17405 16435
rect 17435 16405 17485 16435
rect 17515 16405 17565 16435
rect 17595 16405 17645 16435
rect 17675 16405 17725 16435
rect 17755 16405 17805 16435
rect 17835 16405 17885 16435
rect 17915 16405 17965 16435
rect 17995 16405 18045 16435
rect 18075 16405 18125 16435
rect 18155 16405 18205 16435
rect 18235 16405 18285 16435
rect 18315 16405 18365 16435
rect 18395 16405 18445 16435
rect 18475 16405 18525 16435
rect 18555 16405 18605 16435
rect 18635 16405 18685 16435
rect 18715 16405 18765 16435
rect 18795 16405 18845 16435
rect 18875 16405 18925 16435
rect 18955 16405 19005 16435
rect 19035 16405 19085 16435
rect 19115 16405 19165 16435
rect 19195 16405 19245 16435
rect 19275 16405 19325 16435
rect 19355 16405 19405 16435
rect 19435 16405 19485 16435
rect 19515 16405 19565 16435
rect 19595 16405 19645 16435
rect 19675 16405 19725 16435
rect 19755 16405 19805 16435
rect 19835 16405 19885 16435
rect 19915 16405 19965 16435
rect 19995 16405 20045 16435
rect 20075 16405 20125 16435
rect 20155 16405 20205 16435
rect 20235 16405 20285 16435
rect 20315 16405 20365 16435
rect 20395 16405 20445 16435
rect 20475 16405 20525 16435
rect 20555 16405 20605 16435
rect 20635 16405 20685 16435
rect 20715 16405 20765 16435
rect 20795 16405 20845 16435
rect 20875 16405 20925 16435
rect 20955 16405 20960 16435
rect 0 16400 20960 16405
rect 0 16355 20960 16360
rect 0 16325 4565 16355
rect 4595 16325 9845 16355
rect 9875 16325 16365 16355
rect 16395 16325 20960 16355
rect 0 16320 20960 16325
rect 0 16275 20960 16280
rect 0 16245 5 16275
rect 35 16245 85 16275
rect 115 16245 165 16275
rect 195 16245 245 16275
rect 275 16245 325 16275
rect 355 16245 405 16275
rect 435 16245 485 16275
rect 515 16245 565 16275
rect 595 16245 645 16275
rect 675 16245 725 16275
rect 755 16245 805 16275
rect 835 16245 885 16275
rect 915 16245 965 16275
rect 995 16245 1045 16275
rect 1075 16245 1125 16275
rect 1155 16245 1205 16275
rect 1235 16245 1285 16275
rect 1315 16245 1365 16275
rect 1395 16245 1445 16275
rect 1475 16245 1525 16275
rect 1555 16245 1605 16275
rect 1635 16245 1685 16275
rect 1715 16245 1765 16275
rect 1795 16245 1845 16275
rect 1875 16245 1925 16275
rect 1955 16245 2005 16275
rect 2035 16245 2085 16275
rect 2115 16245 2165 16275
rect 2195 16245 2245 16275
rect 2275 16245 2325 16275
rect 2355 16245 2405 16275
rect 2435 16245 2485 16275
rect 2515 16245 2565 16275
rect 2595 16245 2645 16275
rect 2675 16245 2725 16275
rect 2755 16245 2805 16275
rect 2835 16245 2885 16275
rect 2915 16245 2965 16275
rect 2995 16245 3045 16275
rect 3075 16245 3125 16275
rect 3155 16245 3205 16275
rect 3235 16245 3285 16275
rect 3315 16245 3365 16275
rect 3395 16245 3445 16275
rect 3475 16245 3525 16275
rect 3555 16245 3605 16275
rect 3635 16245 3685 16275
rect 3715 16245 3765 16275
rect 3795 16245 3845 16275
rect 3875 16245 3925 16275
rect 3955 16245 4005 16275
rect 4035 16245 4085 16275
rect 4115 16245 4165 16275
rect 4195 16245 4485 16275
rect 4515 16245 4645 16275
rect 4675 16245 6245 16275
rect 6275 16245 6325 16275
rect 6355 16245 6405 16275
rect 6435 16245 6485 16275
rect 6515 16245 6565 16275
rect 6595 16245 6645 16275
rect 6675 16245 6725 16275
rect 6755 16245 6805 16275
rect 6835 16245 6885 16275
rect 6915 16245 6965 16275
rect 6995 16245 7045 16275
rect 7075 16245 7125 16275
rect 7155 16245 7205 16275
rect 7235 16245 7285 16275
rect 7315 16245 7365 16275
rect 7395 16245 7445 16275
rect 7475 16245 7525 16275
rect 7555 16245 7605 16275
rect 7635 16245 7685 16275
rect 7715 16245 7765 16275
rect 7795 16245 7845 16275
rect 7875 16245 7925 16275
rect 7955 16245 8005 16275
rect 8035 16245 8085 16275
rect 8115 16245 8165 16275
rect 8195 16245 8245 16275
rect 8275 16245 8325 16275
rect 8355 16245 8405 16275
rect 8435 16245 8485 16275
rect 8515 16245 8565 16275
rect 8595 16245 8645 16275
rect 8675 16245 8725 16275
rect 8755 16245 8805 16275
rect 8835 16245 8885 16275
rect 8915 16245 8965 16275
rect 8995 16245 9045 16275
rect 9075 16245 9125 16275
rect 9155 16245 9205 16275
rect 9235 16245 9285 16275
rect 9315 16245 9365 16275
rect 9395 16245 9445 16275
rect 9475 16245 9765 16275
rect 9795 16245 9925 16275
rect 9955 16245 11565 16275
rect 11595 16245 11645 16275
rect 11675 16245 11725 16275
rect 11755 16245 11805 16275
rect 11835 16245 11885 16275
rect 11915 16245 11965 16275
rect 11995 16245 12045 16275
rect 12075 16245 12125 16275
rect 12155 16245 12205 16275
rect 12235 16245 12285 16275
rect 12315 16245 12365 16275
rect 12395 16245 12445 16275
rect 12475 16245 12525 16275
rect 12555 16245 12605 16275
rect 12635 16245 12685 16275
rect 12715 16245 12765 16275
rect 12795 16245 12845 16275
rect 12875 16245 12925 16275
rect 12955 16245 13005 16275
rect 13035 16245 13085 16275
rect 13115 16245 13165 16275
rect 13195 16245 13245 16275
rect 13275 16245 13325 16275
rect 13355 16245 13405 16275
rect 13435 16245 13485 16275
rect 13515 16245 13565 16275
rect 13595 16245 13645 16275
rect 13675 16245 13725 16275
rect 13755 16245 13805 16275
rect 13835 16245 13885 16275
rect 13915 16245 13965 16275
rect 13995 16245 14045 16275
rect 14075 16245 14125 16275
rect 14155 16245 14205 16275
rect 14235 16245 14285 16275
rect 14315 16245 14365 16275
rect 14395 16245 14445 16275
rect 14475 16245 14525 16275
rect 14555 16245 14605 16275
rect 14635 16245 14685 16275
rect 14715 16245 16285 16275
rect 16315 16245 16445 16275
rect 16475 16245 16765 16275
rect 16795 16245 16845 16275
rect 16875 16245 16925 16275
rect 16955 16245 17005 16275
rect 17035 16245 17085 16275
rect 17115 16245 17165 16275
rect 17195 16245 17245 16275
rect 17275 16245 17325 16275
rect 17355 16245 17405 16275
rect 17435 16245 17485 16275
rect 17515 16245 17565 16275
rect 17595 16245 17645 16275
rect 17675 16245 17725 16275
rect 17755 16245 17805 16275
rect 17835 16245 17885 16275
rect 17915 16245 17965 16275
rect 17995 16245 18045 16275
rect 18075 16245 18125 16275
rect 18155 16245 18205 16275
rect 18235 16245 18285 16275
rect 18315 16245 18365 16275
rect 18395 16245 18445 16275
rect 18475 16245 18525 16275
rect 18555 16245 18605 16275
rect 18635 16245 18685 16275
rect 18715 16245 18765 16275
rect 18795 16245 18845 16275
rect 18875 16245 18925 16275
rect 18955 16245 19005 16275
rect 19035 16245 19085 16275
rect 19115 16245 19165 16275
rect 19195 16245 19245 16275
rect 19275 16245 19325 16275
rect 19355 16245 19405 16275
rect 19435 16245 19485 16275
rect 19515 16245 19565 16275
rect 19595 16245 19645 16275
rect 19675 16245 19725 16275
rect 19755 16245 19805 16275
rect 19835 16245 19885 16275
rect 19915 16245 19965 16275
rect 19995 16245 20045 16275
rect 20075 16245 20125 16275
rect 20155 16245 20205 16275
rect 20235 16245 20285 16275
rect 20315 16245 20365 16275
rect 20395 16245 20445 16275
rect 20475 16245 20525 16275
rect 20555 16245 20605 16275
rect 20635 16245 20685 16275
rect 20715 16245 20765 16275
rect 20795 16245 20845 16275
rect 20875 16245 20925 16275
rect 20955 16245 20960 16275
rect 0 16240 20960 16245
rect 0 16195 20960 16200
rect 0 16165 5 16195
rect 35 16165 85 16195
rect 115 16165 165 16195
rect 195 16165 245 16195
rect 275 16165 325 16195
rect 355 16165 405 16195
rect 435 16165 485 16195
rect 515 16165 565 16195
rect 595 16165 645 16195
rect 675 16165 725 16195
rect 755 16165 805 16195
rect 835 16165 885 16195
rect 915 16165 965 16195
rect 995 16165 1045 16195
rect 1075 16165 1125 16195
rect 1155 16165 1205 16195
rect 1235 16165 1285 16195
rect 1315 16165 1365 16195
rect 1395 16165 1445 16195
rect 1475 16165 1525 16195
rect 1555 16165 1605 16195
rect 1635 16165 1685 16195
rect 1715 16165 1765 16195
rect 1795 16165 1845 16195
rect 1875 16165 1925 16195
rect 1955 16165 2005 16195
rect 2035 16165 2085 16195
rect 2115 16165 2165 16195
rect 2195 16165 2245 16195
rect 2275 16165 2325 16195
rect 2355 16165 2405 16195
rect 2435 16165 2485 16195
rect 2515 16165 2565 16195
rect 2595 16165 2645 16195
rect 2675 16165 2725 16195
rect 2755 16165 2805 16195
rect 2835 16165 2885 16195
rect 2915 16165 2965 16195
rect 2995 16165 3045 16195
rect 3075 16165 3125 16195
rect 3155 16165 3205 16195
rect 3235 16165 3285 16195
rect 3315 16165 3365 16195
rect 3395 16165 3445 16195
rect 3475 16165 3525 16195
rect 3555 16165 3605 16195
rect 3635 16165 3685 16195
rect 3715 16165 3765 16195
rect 3795 16165 3845 16195
rect 3875 16165 3925 16195
rect 3955 16165 4005 16195
rect 4035 16165 4085 16195
rect 4115 16165 4165 16195
rect 4195 16165 4725 16195
rect 4755 16165 4885 16195
rect 4915 16165 5045 16195
rect 5075 16165 5205 16195
rect 5235 16165 5365 16195
rect 5395 16165 5525 16195
rect 5555 16165 5685 16195
rect 5715 16165 6245 16195
rect 6275 16165 6325 16195
rect 6355 16165 6405 16195
rect 6435 16165 6485 16195
rect 6515 16165 6565 16195
rect 6595 16165 6645 16195
rect 6675 16165 6725 16195
rect 6755 16165 6805 16195
rect 6835 16165 6885 16195
rect 6915 16165 6965 16195
rect 6995 16165 7045 16195
rect 7075 16165 7125 16195
rect 7155 16165 7205 16195
rect 7235 16165 7285 16195
rect 7315 16165 7365 16195
rect 7395 16165 7445 16195
rect 7475 16165 7525 16195
rect 7555 16165 7605 16195
rect 7635 16165 7685 16195
rect 7715 16165 7765 16195
rect 7795 16165 7845 16195
rect 7875 16165 7925 16195
rect 7955 16165 8005 16195
rect 8035 16165 8085 16195
rect 8115 16165 8165 16195
rect 8195 16165 8245 16195
rect 8275 16165 8325 16195
rect 8355 16165 8405 16195
rect 8435 16165 8485 16195
rect 8515 16165 8565 16195
rect 8595 16165 8645 16195
rect 8675 16165 8725 16195
rect 8755 16165 8805 16195
rect 8835 16165 8885 16195
rect 8915 16165 8965 16195
rect 8995 16165 9045 16195
rect 9075 16165 9125 16195
rect 9155 16165 9205 16195
rect 9235 16165 9285 16195
rect 9315 16165 9365 16195
rect 9395 16165 9445 16195
rect 9475 16165 10005 16195
rect 10035 16165 10165 16195
rect 10195 16165 10325 16195
rect 10355 16165 10485 16195
rect 10515 16165 10645 16195
rect 10675 16165 10805 16195
rect 10835 16165 10965 16195
rect 10995 16165 11565 16195
rect 11595 16165 11645 16195
rect 11675 16165 11725 16195
rect 11755 16165 11805 16195
rect 11835 16165 11885 16195
rect 11915 16165 11965 16195
rect 11995 16165 12045 16195
rect 12075 16165 12125 16195
rect 12155 16165 12205 16195
rect 12235 16165 12285 16195
rect 12315 16165 12365 16195
rect 12395 16165 12445 16195
rect 12475 16165 12525 16195
rect 12555 16165 12605 16195
rect 12635 16165 12685 16195
rect 12715 16165 12765 16195
rect 12795 16165 12845 16195
rect 12875 16165 12925 16195
rect 12955 16165 13005 16195
rect 13035 16165 13085 16195
rect 13115 16165 13165 16195
rect 13195 16165 13245 16195
rect 13275 16165 13325 16195
rect 13355 16165 13405 16195
rect 13435 16165 13485 16195
rect 13515 16165 13565 16195
rect 13595 16165 13645 16195
rect 13675 16165 13725 16195
rect 13755 16165 13805 16195
rect 13835 16165 13885 16195
rect 13915 16165 13965 16195
rect 13995 16165 14045 16195
rect 14075 16165 14125 16195
rect 14155 16165 14205 16195
rect 14235 16165 14285 16195
rect 14315 16165 14365 16195
rect 14395 16165 14445 16195
rect 14475 16165 14525 16195
rect 14555 16165 14605 16195
rect 14635 16165 14685 16195
rect 14715 16165 15245 16195
rect 15275 16165 15405 16195
rect 15435 16165 15565 16195
rect 15595 16165 15725 16195
rect 15755 16165 15885 16195
rect 15915 16165 16045 16195
rect 16075 16165 16205 16195
rect 16235 16165 16765 16195
rect 16795 16165 16845 16195
rect 16875 16165 16925 16195
rect 16955 16165 17005 16195
rect 17035 16165 17085 16195
rect 17115 16165 17165 16195
rect 17195 16165 17245 16195
rect 17275 16165 17325 16195
rect 17355 16165 17405 16195
rect 17435 16165 17485 16195
rect 17515 16165 17565 16195
rect 17595 16165 17645 16195
rect 17675 16165 17725 16195
rect 17755 16165 17805 16195
rect 17835 16165 17885 16195
rect 17915 16165 17965 16195
rect 17995 16165 18045 16195
rect 18075 16165 18125 16195
rect 18155 16165 18205 16195
rect 18235 16165 18285 16195
rect 18315 16165 18365 16195
rect 18395 16165 18445 16195
rect 18475 16165 18525 16195
rect 18555 16165 18605 16195
rect 18635 16165 18685 16195
rect 18715 16165 18765 16195
rect 18795 16165 18845 16195
rect 18875 16165 18925 16195
rect 18955 16165 19005 16195
rect 19035 16165 19085 16195
rect 19115 16165 19165 16195
rect 19195 16165 19245 16195
rect 19275 16165 19325 16195
rect 19355 16165 19405 16195
rect 19435 16165 19485 16195
rect 19515 16165 19565 16195
rect 19595 16165 19645 16195
rect 19675 16165 19725 16195
rect 19755 16165 19805 16195
rect 19835 16165 19885 16195
rect 19915 16165 19965 16195
rect 19995 16165 20045 16195
rect 20075 16165 20125 16195
rect 20155 16165 20205 16195
rect 20235 16165 20285 16195
rect 20315 16165 20365 16195
rect 20395 16165 20445 16195
rect 20475 16165 20525 16195
rect 20555 16165 20605 16195
rect 20635 16165 20685 16195
rect 20715 16165 20765 16195
rect 20795 16165 20845 16195
rect 20875 16165 20925 16195
rect 20955 16165 20960 16195
rect 0 16160 20960 16165
rect 0 16115 20960 16120
rect 0 16085 4805 16115
rect 4835 16085 10085 16115
rect 10115 16085 16125 16115
rect 16155 16085 20960 16115
rect 0 16080 20960 16085
rect 0 16035 20960 16040
rect 0 16005 5 16035
rect 35 16005 85 16035
rect 115 16005 165 16035
rect 195 16005 245 16035
rect 275 16005 325 16035
rect 355 16005 405 16035
rect 435 16005 485 16035
rect 515 16005 565 16035
rect 595 16005 645 16035
rect 675 16005 725 16035
rect 755 16005 805 16035
rect 835 16005 885 16035
rect 915 16005 965 16035
rect 995 16005 1045 16035
rect 1075 16005 1125 16035
rect 1155 16005 1205 16035
rect 1235 16005 1285 16035
rect 1315 16005 1365 16035
rect 1395 16005 1445 16035
rect 1475 16005 1525 16035
rect 1555 16005 1605 16035
rect 1635 16005 1685 16035
rect 1715 16005 1765 16035
rect 1795 16005 1845 16035
rect 1875 16005 1925 16035
rect 1955 16005 2005 16035
rect 2035 16005 2085 16035
rect 2115 16005 2165 16035
rect 2195 16005 2245 16035
rect 2275 16005 2325 16035
rect 2355 16005 2405 16035
rect 2435 16005 2485 16035
rect 2515 16005 2565 16035
rect 2595 16005 2645 16035
rect 2675 16005 2725 16035
rect 2755 16005 2805 16035
rect 2835 16005 2885 16035
rect 2915 16005 2965 16035
rect 2995 16005 3045 16035
rect 3075 16005 3125 16035
rect 3155 16005 3205 16035
rect 3235 16005 3285 16035
rect 3315 16005 3365 16035
rect 3395 16005 3445 16035
rect 3475 16005 3525 16035
rect 3555 16005 3605 16035
rect 3635 16005 3685 16035
rect 3715 16005 3765 16035
rect 3795 16005 3845 16035
rect 3875 16005 3925 16035
rect 3955 16005 4005 16035
rect 4035 16005 4085 16035
rect 4115 16005 4165 16035
rect 4195 16005 4725 16035
rect 4755 16005 4885 16035
rect 4915 16005 5045 16035
rect 5075 16005 5205 16035
rect 5235 16005 5365 16035
rect 5395 16005 5525 16035
rect 5555 16005 5685 16035
rect 5715 16005 6245 16035
rect 6275 16005 6325 16035
rect 6355 16005 6405 16035
rect 6435 16005 6485 16035
rect 6515 16005 6565 16035
rect 6595 16005 6645 16035
rect 6675 16005 6725 16035
rect 6755 16005 6805 16035
rect 6835 16005 6885 16035
rect 6915 16005 6965 16035
rect 6995 16005 7045 16035
rect 7075 16005 7125 16035
rect 7155 16005 7205 16035
rect 7235 16005 7285 16035
rect 7315 16005 7365 16035
rect 7395 16005 7445 16035
rect 7475 16005 7525 16035
rect 7555 16005 7605 16035
rect 7635 16005 7685 16035
rect 7715 16005 7765 16035
rect 7795 16005 7845 16035
rect 7875 16005 7925 16035
rect 7955 16005 8005 16035
rect 8035 16005 8085 16035
rect 8115 16005 8165 16035
rect 8195 16005 8245 16035
rect 8275 16005 8325 16035
rect 8355 16005 8405 16035
rect 8435 16005 8485 16035
rect 8515 16005 8565 16035
rect 8595 16005 8645 16035
rect 8675 16005 8725 16035
rect 8755 16005 8805 16035
rect 8835 16005 8885 16035
rect 8915 16005 8965 16035
rect 8995 16005 9045 16035
rect 9075 16005 9125 16035
rect 9155 16005 9205 16035
rect 9235 16005 9285 16035
rect 9315 16005 9365 16035
rect 9395 16005 9445 16035
rect 9475 16005 10005 16035
rect 10035 16005 10165 16035
rect 10195 16005 10325 16035
rect 10355 16005 10485 16035
rect 10515 16005 10645 16035
rect 10675 16005 10805 16035
rect 10835 16005 10965 16035
rect 10995 16005 11565 16035
rect 11595 16005 11645 16035
rect 11675 16005 11725 16035
rect 11755 16005 11805 16035
rect 11835 16005 11885 16035
rect 11915 16005 11965 16035
rect 11995 16005 12045 16035
rect 12075 16005 12125 16035
rect 12155 16005 12205 16035
rect 12235 16005 12285 16035
rect 12315 16005 12365 16035
rect 12395 16005 12445 16035
rect 12475 16005 12525 16035
rect 12555 16005 12605 16035
rect 12635 16005 12685 16035
rect 12715 16005 12765 16035
rect 12795 16005 12845 16035
rect 12875 16005 12925 16035
rect 12955 16005 13005 16035
rect 13035 16005 13085 16035
rect 13115 16005 13165 16035
rect 13195 16005 13245 16035
rect 13275 16005 13325 16035
rect 13355 16005 13405 16035
rect 13435 16005 13485 16035
rect 13515 16005 13565 16035
rect 13595 16005 13645 16035
rect 13675 16005 13725 16035
rect 13755 16005 13805 16035
rect 13835 16005 13885 16035
rect 13915 16005 13965 16035
rect 13995 16005 14045 16035
rect 14075 16005 14125 16035
rect 14155 16005 14205 16035
rect 14235 16005 14285 16035
rect 14315 16005 14365 16035
rect 14395 16005 14445 16035
rect 14475 16005 14525 16035
rect 14555 16005 14605 16035
rect 14635 16005 14685 16035
rect 14715 16005 15245 16035
rect 15275 16005 15405 16035
rect 15435 16005 15565 16035
rect 15595 16005 15725 16035
rect 15755 16005 15885 16035
rect 15915 16005 16045 16035
rect 16075 16005 16205 16035
rect 16235 16005 16765 16035
rect 16795 16005 16845 16035
rect 16875 16005 16925 16035
rect 16955 16005 17005 16035
rect 17035 16005 17085 16035
rect 17115 16005 17165 16035
rect 17195 16005 17245 16035
rect 17275 16005 17325 16035
rect 17355 16005 17405 16035
rect 17435 16005 17485 16035
rect 17515 16005 17565 16035
rect 17595 16005 17645 16035
rect 17675 16005 17725 16035
rect 17755 16005 17805 16035
rect 17835 16005 17885 16035
rect 17915 16005 17965 16035
rect 17995 16005 18045 16035
rect 18075 16005 18125 16035
rect 18155 16005 18205 16035
rect 18235 16005 18285 16035
rect 18315 16005 18365 16035
rect 18395 16005 18445 16035
rect 18475 16005 18525 16035
rect 18555 16005 18605 16035
rect 18635 16005 18685 16035
rect 18715 16005 18765 16035
rect 18795 16005 18845 16035
rect 18875 16005 18925 16035
rect 18955 16005 19005 16035
rect 19035 16005 19085 16035
rect 19115 16005 19165 16035
rect 19195 16005 19245 16035
rect 19275 16005 19325 16035
rect 19355 16005 19405 16035
rect 19435 16005 19485 16035
rect 19515 16005 19565 16035
rect 19595 16005 19645 16035
rect 19675 16005 19725 16035
rect 19755 16005 19805 16035
rect 19835 16005 19885 16035
rect 19915 16005 19965 16035
rect 19995 16005 20045 16035
rect 20075 16005 20125 16035
rect 20155 16005 20205 16035
rect 20235 16005 20285 16035
rect 20315 16005 20365 16035
rect 20395 16005 20445 16035
rect 20475 16005 20525 16035
rect 20555 16005 20605 16035
rect 20635 16005 20685 16035
rect 20715 16005 20765 16035
rect 20795 16005 20845 16035
rect 20875 16005 20925 16035
rect 20955 16005 20960 16035
rect 0 16000 20960 16005
rect 0 15955 20960 15960
rect 0 15925 4965 15955
rect 4995 15925 10245 15955
rect 10275 15925 15965 15955
rect 15995 15925 20960 15955
rect 0 15920 20960 15925
rect 0 15875 20960 15880
rect 0 15845 5 15875
rect 35 15845 85 15875
rect 115 15845 165 15875
rect 195 15845 245 15875
rect 275 15845 325 15875
rect 355 15845 405 15875
rect 435 15845 485 15875
rect 515 15845 565 15875
rect 595 15845 645 15875
rect 675 15845 725 15875
rect 755 15845 805 15875
rect 835 15845 885 15875
rect 915 15845 965 15875
rect 995 15845 1045 15875
rect 1075 15845 1125 15875
rect 1155 15845 1205 15875
rect 1235 15845 1285 15875
rect 1315 15845 1365 15875
rect 1395 15845 1445 15875
rect 1475 15845 1525 15875
rect 1555 15845 1605 15875
rect 1635 15845 1685 15875
rect 1715 15845 1765 15875
rect 1795 15845 1845 15875
rect 1875 15845 1925 15875
rect 1955 15845 2005 15875
rect 2035 15845 2085 15875
rect 2115 15845 2165 15875
rect 2195 15845 2245 15875
rect 2275 15845 2325 15875
rect 2355 15845 2405 15875
rect 2435 15845 2485 15875
rect 2515 15845 2565 15875
rect 2595 15845 2645 15875
rect 2675 15845 2725 15875
rect 2755 15845 2805 15875
rect 2835 15845 2885 15875
rect 2915 15845 2965 15875
rect 2995 15845 3045 15875
rect 3075 15845 3125 15875
rect 3155 15845 3205 15875
rect 3235 15845 3285 15875
rect 3315 15845 3365 15875
rect 3395 15845 3445 15875
rect 3475 15845 3525 15875
rect 3555 15845 3605 15875
rect 3635 15845 3685 15875
rect 3715 15845 3765 15875
rect 3795 15845 3845 15875
rect 3875 15845 3925 15875
rect 3955 15845 4005 15875
rect 4035 15845 4085 15875
rect 4115 15845 4165 15875
rect 4195 15845 4725 15875
rect 4755 15845 4885 15875
rect 4915 15845 5045 15875
rect 5075 15845 5205 15875
rect 5235 15845 5365 15875
rect 5395 15845 5525 15875
rect 5555 15845 5685 15875
rect 5715 15845 6245 15875
rect 6275 15845 6325 15875
rect 6355 15845 6405 15875
rect 6435 15845 6485 15875
rect 6515 15845 6565 15875
rect 6595 15845 6645 15875
rect 6675 15845 6725 15875
rect 6755 15845 6805 15875
rect 6835 15845 6885 15875
rect 6915 15845 6965 15875
rect 6995 15845 7045 15875
rect 7075 15845 7125 15875
rect 7155 15845 7205 15875
rect 7235 15845 7285 15875
rect 7315 15845 7365 15875
rect 7395 15845 7445 15875
rect 7475 15845 7525 15875
rect 7555 15845 7605 15875
rect 7635 15845 7685 15875
rect 7715 15845 7765 15875
rect 7795 15845 7845 15875
rect 7875 15845 7925 15875
rect 7955 15845 8005 15875
rect 8035 15845 8085 15875
rect 8115 15845 8165 15875
rect 8195 15845 8245 15875
rect 8275 15845 8325 15875
rect 8355 15845 8405 15875
rect 8435 15845 8485 15875
rect 8515 15845 8565 15875
rect 8595 15845 8645 15875
rect 8675 15845 8725 15875
rect 8755 15845 8805 15875
rect 8835 15845 8885 15875
rect 8915 15845 8965 15875
rect 8995 15845 9045 15875
rect 9075 15845 9125 15875
rect 9155 15845 9205 15875
rect 9235 15845 9285 15875
rect 9315 15845 9365 15875
rect 9395 15845 9445 15875
rect 9475 15845 10005 15875
rect 10035 15845 10165 15875
rect 10195 15845 10325 15875
rect 10355 15845 10485 15875
rect 10515 15845 10645 15875
rect 10675 15845 10805 15875
rect 10835 15845 10965 15875
rect 10995 15845 11565 15875
rect 11595 15845 11645 15875
rect 11675 15845 11725 15875
rect 11755 15845 11805 15875
rect 11835 15845 11885 15875
rect 11915 15845 11965 15875
rect 11995 15845 12045 15875
rect 12075 15845 12125 15875
rect 12155 15845 12205 15875
rect 12235 15845 12285 15875
rect 12315 15845 12365 15875
rect 12395 15845 12445 15875
rect 12475 15845 12525 15875
rect 12555 15845 12605 15875
rect 12635 15845 12685 15875
rect 12715 15845 12765 15875
rect 12795 15845 12845 15875
rect 12875 15845 12925 15875
rect 12955 15845 13005 15875
rect 13035 15845 13085 15875
rect 13115 15845 13165 15875
rect 13195 15845 13245 15875
rect 13275 15845 13325 15875
rect 13355 15845 13405 15875
rect 13435 15845 13485 15875
rect 13515 15845 13565 15875
rect 13595 15845 13645 15875
rect 13675 15845 13725 15875
rect 13755 15845 13805 15875
rect 13835 15845 13885 15875
rect 13915 15845 13965 15875
rect 13995 15845 14045 15875
rect 14075 15845 14125 15875
rect 14155 15845 14205 15875
rect 14235 15845 14285 15875
rect 14315 15845 14365 15875
rect 14395 15845 14445 15875
rect 14475 15845 14525 15875
rect 14555 15845 14605 15875
rect 14635 15845 14685 15875
rect 14715 15845 15245 15875
rect 15275 15845 15405 15875
rect 15435 15845 15565 15875
rect 15595 15845 15725 15875
rect 15755 15845 15885 15875
rect 15915 15845 16045 15875
rect 16075 15845 16205 15875
rect 16235 15845 16765 15875
rect 16795 15845 16845 15875
rect 16875 15845 16925 15875
rect 16955 15845 17005 15875
rect 17035 15845 17085 15875
rect 17115 15845 17165 15875
rect 17195 15845 17245 15875
rect 17275 15845 17325 15875
rect 17355 15845 17405 15875
rect 17435 15845 17485 15875
rect 17515 15845 17565 15875
rect 17595 15845 17645 15875
rect 17675 15845 17725 15875
rect 17755 15845 17805 15875
rect 17835 15845 17885 15875
rect 17915 15845 17965 15875
rect 17995 15845 18045 15875
rect 18075 15845 18125 15875
rect 18155 15845 18205 15875
rect 18235 15845 18285 15875
rect 18315 15845 18365 15875
rect 18395 15845 18445 15875
rect 18475 15845 18525 15875
rect 18555 15845 18605 15875
rect 18635 15845 18685 15875
rect 18715 15845 18765 15875
rect 18795 15845 18845 15875
rect 18875 15845 18925 15875
rect 18955 15845 19005 15875
rect 19035 15845 19085 15875
rect 19115 15845 19165 15875
rect 19195 15845 19245 15875
rect 19275 15845 19325 15875
rect 19355 15845 19405 15875
rect 19435 15845 19485 15875
rect 19515 15845 19565 15875
rect 19595 15845 19645 15875
rect 19675 15845 19725 15875
rect 19755 15845 19805 15875
rect 19835 15845 19885 15875
rect 19915 15845 19965 15875
rect 19995 15845 20045 15875
rect 20075 15845 20125 15875
rect 20155 15845 20205 15875
rect 20235 15845 20285 15875
rect 20315 15845 20365 15875
rect 20395 15845 20445 15875
rect 20475 15845 20525 15875
rect 20555 15845 20605 15875
rect 20635 15845 20685 15875
rect 20715 15845 20765 15875
rect 20795 15845 20845 15875
rect 20875 15845 20925 15875
rect 20955 15845 20960 15875
rect 0 15840 20960 15845
rect 0 15795 20960 15800
rect 0 15765 5125 15795
rect 5155 15765 10405 15795
rect 10435 15765 15805 15795
rect 15835 15765 20960 15795
rect 0 15760 20960 15765
rect 0 15715 20960 15720
rect 0 15685 5 15715
rect 35 15685 85 15715
rect 115 15685 165 15715
rect 195 15685 245 15715
rect 275 15685 325 15715
rect 355 15685 405 15715
rect 435 15685 485 15715
rect 515 15685 565 15715
rect 595 15685 645 15715
rect 675 15685 725 15715
rect 755 15685 805 15715
rect 835 15685 885 15715
rect 915 15685 965 15715
rect 995 15685 1045 15715
rect 1075 15685 1125 15715
rect 1155 15685 1205 15715
rect 1235 15685 1285 15715
rect 1315 15685 1365 15715
rect 1395 15685 1445 15715
rect 1475 15685 1525 15715
rect 1555 15685 1605 15715
rect 1635 15685 1685 15715
rect 1715 15685 1765 15715
rect 1795 15685 1845 15715
rect 1875 15685 1925 15715
rect 1955 15685 2005 15715
rect 2035 15685 2085 15715
rect 2115 15685 2165 15715
rect 2195 15685 2245 15715
rect 2275 15685 2325 15715
rect 2355 15685 2405 15715
rect 2435 15685 2485 15715
rect 2515 15685 2565 15715
rect 2595 15685 2645 15715
rect 2675 15685 2725 15715
rect 2755 15685 2805 15715
rect 2835 15685 2885 15715
rect 2915 15685 2965 15715
rect 2995 15685 3045 15715
rect 3075 15685 3125 15715
rect 3155 15685 3205 15715
rect 3235 15685 3285 15715
rect 3315 15685 3365 15715
rect 3395 15685 3445 15715
rect 3475 15685 3525 15715
rect 3555 15685 3605 15715
rect 3635 15685 3685 15715
rect 3715 15685 3765 15715
rect 3795 15685 3845 15715
rect 3875 15685 3925 15715
rect 3955 15685 4005 15715
rect 4035 15685 4085 15715
rect 4115 15685 4165 15715
rect 4195 15685 4725 15715
rect 4755 15685 4885 15715
rect 4915 15685 5045 15715
rect 5075 15685 5205 15715
rect 5235 15685 5365 15715
rect 5395 15685 5525 15715
rect 5555 15685 5685 15715
rect 5715 15685 6245 15715
rect 6275 15685 6325 15715
rect 6355 15685 6405 15715
rect 6435 15685 6485 15715
rect 6515 15685 6565 15715
rect 6595 15685 6645 15715
rect 6675 15685 6725 15715
rect 6755 15685 6805 15715
rect 6835 15685 6885 15715
rect 6915 15685 6965 15715
rect 6995 15685 7045 15715
rect 7075 15685 7125 15715
rect 7155 15685 7205 15715
rect 7235 15685 7285 15715
rect 7315 15685 7365 15715
rect 7395 15685 7445 15715
rect 7475 15685 7525 15715
rect 7555 15685 7605 15715
rect 7635 15685 7685 15715
rect 7715 15685 7765 15715
rect 7795 15685 7845 15715
rect 7875 15685 7925 15715
rect 7955 15685 8005 15715
rect 8035 15685 8085 15715
rect 8115 15685 8165 15715
rect 8195 15685 8245 15715
rect 8275 15685 8325 15715
rect 8355 15685 8405 15715
rect 8435 15685 8485 15715
rect 8515 15685 8565 15715
rect 8595 15685 8645 15715
rect 8675 15685 8725 15715
rect 8755 15685 8805 15715
rect 8835 15685 8885 15715
rect 8915 15685 8965 15715
rect 8995 15685 9045 15715
rect 9075 15685 9125 15715
rect 9155 15685 9205 15715
rect 9235 15685 9285 15715
rect 9315 15685 9365 15715
rect 9395 15685 9445 15715
rect 9475 15685 10005 15715
rect 10035 15685 10165 15715
rect 10195 15685 10325 15715
rect 10355 15685 10485 15715
rect 10515 15685 10645 15715
rect 10675 15685 10805 15715
rect 10835 15685 10965 15715
rect 10995 15685 11565 15715
rect 11595 15685 11645 15715
rect 11675 15685 11725 15715
rect 11755 15685 11805 15715
rect 11835 15685 11885 15715
rect 11915 15685 11965 15715
rect 11995 15685 12045 15715
rect 12075 15685 12125 15715
rect 12155 15685 12205 15715
rect 12235 15685 12285 15715
rect 12315 15685 12365 15715
rect 12395 15685 12445 15715
rect 12475 15685 12525 15715
rect 12555 15685 12605 15715
rect 12635 15685 12685 15715
rect 12715 15685 12765 15715
rect 12795 15685 12845 15715
rect 12875 15685 12925 15715
rect 12955 15685 13005 15715
rect 13035 15685 13085 15715
rect 13115 15685 13165 15715
rect 13195 15685 13245 15715
rect 13275 15685 13325 15715
rect 13355 15685 13405 15715
rect 13435 15685 13485 15715
rect 13515 15685 13565 15715
rect 13595 15685 13645 15715
rect 13675 15685 13725 15715
rect 13755 15685 13805 15715
rect 13835 15685 13885 15715
rect 13915 15685 13965 15715
rect 13995 15685 14045 15715
rect 14075 15685 14125 15715
rect 14155 15685 14205 15715
rect 14235 15685 14285 15715
rect 14315 15685 14365 15715
rect 14395 15685 14445 15715
rect 14475 15685 14525 15715
rect 14555 15685 14605 15715
rect 14635 15685 14685 15715
rect 14715 15685 15245 15715
rect 15275 15685 15405 15715
rect 15435 15685 15565 15715
rect 15595 15685 15725 15715
rect 15755 15685 15885 15715
rect 15915 15685 16045 15715
rect 16075 15685 16205 15715
rect 16235 15685 16765 15715
rect 16795 15685 16845 15715
rect 16875 15685 16925 15715
rect 16955 15685 17005 15715
rect 17035 15685 17085 15715
rect 17115 15685 17165 15715
rect 17195 15685 17245 15715
rect 17275 15685 17325 15715
rect 17355 15685 17405 15715
rect 17435 15685 17485 15715
rect 17515 15685 17565 15715
rect 17595 15685 17645 15715
rect 17675 15685 17725 15715
rect 17755 15685 17805 15715
rect 17835 15685 17885 15715
rect 17915 15685 17965 15715
rect 17995 15685 18045 15715
rect 18075 15685 18125 15715
rect 18155 15685 18205 15715
rect 18235 15685 18285 15715
rect 18315 15685 18365 15715
rect 18395 15685 18445 15715
rect 18475 15685 18525 15715
rect 18555 15685 18605 15715
rect 18635 15685 18685 15715
rect 18715 15685 18765 15715
rect 18795 15685 18845 15715
rect 18875 15685 18925 15715
rect 18955 15685 19005 15715
rect 19035 15685 19085 15715
rect 19115 15685 19165 15715
rect 19195 15685 19245 15715
rect 19275 15685 19325 15715
rect 19355 15685 19405 15715
rect 19435 15685 19485 15715
rect 19515 15685 19565 15715
rect 19595 15685 19645 15715
rect 19675 15685 19725 15715
rect 19755 15685 19805 15715
rect 19835 15685 19885 15715
rect 19915 15685 19965 15715
rect 19995 15685 20045 15715
rect 20075 15685 20125 15715
rect 20155 15685 20205 15715
rect 20235 15685 20285 15715
rect 20315 15685 20365 15715
rect 20395 15685 20445 15715
rect 20475 15685 20525 15715
rect 20555 15685 20605 15715
rect 20635 15685 20685 15715
rect 20715 15685 20765 15715
rect 20795 15685 20845 15715
rect 20875 15685 20925 15715
rect 20955 15685 20960 15715
rect 0 15680 20960 15685
rect 0 15635 20960 15640
rect 0 15605 5285 15635
rect 5315 15605 10565 15635
rect 10595 15605 15645 15635
rect 15675 15605 20960 15635
rect 0 15600 20960 15605
rect 0 15555 20960 15560
rect 0 15525 5 15555
rect 35 15525 85 15555
rect 115 15525 165 15555
rect 195 15525 245 15555
rect 275 15525 325 15555
rect 355 15525 405 15555
rect 435 15525 485 15555
rect 515 15525 565 15555
rect 595 15525 645 15555
rect 675 15525 725 15555
rect 755 15525 805 15555
rect 835 15525 885 15555
rect 915 15525 965 15555
rect 995 15525 1045 15555
rect 1075 15525 1125 15555
rect 1155 15525 1205 15555
rect 1235 15525 1285 15555
rect 1315 15525 1365 15555
rect 1395 15525 1445 15555
rect 1475 15525 1525 15555
rect 1555 15525 1605 15555
rect 1635 15525 1685 15555
rect 1715 15525 1765 15555
rect 1795 15525 1845 15555
rect 1875 15525 1925 15555
rect 1955 15525 2005 15555
rect 2035 15525 2085 15555
rect 2115 15525 2165 15555
rect 2195 15525 2245 15555
rect 2275 15525 2325 15555
rect 2355 15525 2405 15555
rect 2435 15525 2485 15555
rect 2515 15525 2565 15555
rect 2595 15525 2645 15555
rect 2675 15525 2725 15555
rect 2755 15525 2805 15555
rect 2835 15525 2885 15555
rect 2915 15525 2965 15555
rect 2995 15525 3045 15555
rect 3075 15525 3125 15555
rect 3155 15525 3205 15555
rect 3235 15525 3285 15555
rect 3315 15525 3365 15555
rect 3395 15525 3445 15555
rect 3475 15525 3525 15555
rect 3555 15525 3605 15555
rect 3635 15525 3685 15555
rect 3715 15525 3765 15555
rect 3795 15525 3845 15555
rect 3875 15525 3925 15555
rect 3955 15525 4005 15555
rect 4035 15525 4085 15555
rect 4115 15525 4165 15555
rect 4195 15525 4725 15555
rect 4755 15525 4885 15555
rect 4915 15525 5045 15555
rect 5075 15525 5205 15555
rect 5235 15525 5365 15555
rect 5395 15525 5525 15555
rect 5555 15525 5685 15555
rect 5715 15525 6245 15555
rect 6275 15525 6325 15555
rect 6355 15525 6405 15555
rect 6435 15525 6485 15555
rect 6515 15525 6565 15555
rect 6595 15525 6645 15555
rect 6675 15525 6725 15555
rect 6755 15525 6805 15555
rect 6835 15525 6885 15555
rect 6915 15525 6965 15555
rect 6995 15525 7045 15555
rect 7075 15525 7125 15555
rect 7155 15525 7205 15555
rect 7235 15525 7285 15555
rect 7315 15525 7365 15555
rect 7395 15525 7445 15555
rect 7475 15525 7525 15555
rect 7555 15525 7605 15555
rect 7635 15525 7685 15555
rect 7715 15525 7765 15555
rect 7795 15525 7845 15555
rect 7875 15525 7925 15555
rect 7955 15525 8005 15555
rect 8035 15525 8085 15555
rect 8115 15525 8165 15555
rect 8195 15525 8245 15555
rect 8275 15525 8325 15555
rect 8355 15525 8405 15555
rect 8435 15525 8485 15555
rect 8515 15525 8565 15555
rect 8595 15525 8645 15555
rect 8675 15525 8725 15555
rect 8755 15525 8805 15555
rect 8835 15525 8885 15555
rect 8915 15525 8965 15555
rect 8995 15525 9045 15555
rect 9075 15525 9125 15555
rect 9155 15525 9205 15555
rect 9235 15525 9285 15555
rect 9315 15525 9365 15555
rect 9395 15525 9445 15555
rect 9475 15525 10005 15555
rect 10035 15525 10165 15555
rect 10195 15525 10325 15555
rect 10355 15525 10485 15555
rect 10515 15525 10645 15555
rect 10675 15525 10805 15555
rect 10835 15525 10965 15555
rect 10995 15525 11565 15555
rect 11595 15525 11645 15555
rect 11675 15525 11725 15555
rect 11755 15525 11805 15555
rect 11835 15525 11885 15555
rect 11915 15525 11965 15555
rect 11995 15525 12045 15555
rect 12075 15525 12125 15555
rect 12155 15525 12205 15555
rect 12235 15525 12285 15555
rect 12315 15525 12365 15555
rect 12395 15525 12445 15555
rect 12475 15525 12525 15555
rect 12555 15525 12605 15555
rect 12635 15525 12685 15555
rect 12715 15525 12765 15555
rect 12795 15525 12845 15555
rect 12875 15525 12925 15555
rect 12955 15525 13005 15555
rect 13035 15525 13085 15555
rect 13115 15525 13165 15555
rect 13195 15525 13245 15555
rect 13275 15525 13325 15555
rect 13355 15525 13405 15555
rect 13435 15525 13485 15555
rect 13515 15525 13565 15555
rect 13595 15525 13645 15555
rect 13675 15525 13725 15555
rect 13755 15525 13805 15555
rect 13835 15525 13885 15555
rect 13915 15525 13965 15555
rect 13995 15525 14045 15555
rect 14075 15525 14125 15555
rect 14155 15525 14205 15555
rect 14235 15525 14285 15555
rect 14315 15525 14365 15555
rect 14395 15525 14445 15555
rect 14475 15525 14525 15555
rect 14555 15525 14605 15555
rect 14635 15525 14685 15555
rect 14715 15525 15245 15555
rect 15275 15525 15405 15555
rect 15435 15525 15565 15555
rect 15595 15525 15725 15555
rect 15755 15525 15885 15555
rect 15915 15525 16045 15555
rect 16075 15525 16205 15555
rect 16235 15525 16765 15555
rect 16795 15525 16845 15555
rect 16875 15525 16925 15555
rect 16955 15525 17005 15555
rect 17035 15525 17085 15555
rect 17115 15525 17165 15555
rect 17195 15525 17245 15555
rect 17275 15525 17325 15555
rect 17355 15525 17405 15555
rect 17435 15525 17485 15555
rect 17515 15525 17565 15555
rect 17595 15525 17645 15555
rect 17675 15525 17725 15555
rect 17755 15525 17805 15555
rect 17835 15525 17885 15555
rect 17915 15525 17965 15555
rect 17995 15525 18045 15555
rect 18075 15525 18125 15555
rect 18155 15525 18205 15555
rect 18235 15525 18285 15555
rect 18315 15525 18365 15555
rect 18395 15525 18445 15555
rect 18475 15525 18525 15555
rect 18555 15525 18605 15555
rect 18635 15525 18685 15555
rect 18715 15525 18765 15555
rect 18795 15525 18845 15555
rect 18875 15525 18925 15555
rect 18955 15525 19005 15555
rect 19035 15525 19085 15555
rect 19115 15525 19165 15555
rect 19195 15525 19245 15555
rect 19275 15525 19325 15555
rect 19355 15525 19405 15555
rect 19435 15525 19485 15555
rect 19515 15525 19565 15555
rect 19595 15525 19645 15555
rect 19675 15525 19725 15555
rect 19755 15525 19805 15555
rect 19835 15525 19885 15555
rect 19915 15525 19965 15555
rect 19995 15525 20045 15555
rect 20075 15525 20125 15555
rect 20155 15525 20205 15555
rect 20235 15525 20285 15555
rect 20315 15525 20365 15555
rect 20395 15525 20445 15555
rect 20475 15525 20525 15555
rect 20555 15525 20605 15555
rect 20635 15525 20685 15555
rect 20715 15525 20765 15555
rect 20795 15525 20845 15555
rect 20875 15525 20925 15555
rect 20955 15525 20960 15555
rect 0 15520 20960 15525
rect 0 15475 20960 15480
rect 0 15445 5445 15475
rect 5475 15445 10725 15475
rect 10755 15445 15485 15475
rect 15515 15445 20960 15475
rect 0 15440 20960 15445
rect 0 15395 20960 15400
rect 0 15365 5 15395
rect 35 15365 85 15395
rect 115 15365 165 15395
rect 195 15365 245 15395
rect 275 15365 325 15395
rect 355 15365 405 15395
rect 435 15365 485 15395
rect 515 15365 565 15395
rect 595 15365 645 15395
rect 675 15365 725 15395
rect 755 15365 805 15395
rect 835 15365 885 15395
rect 915 15365 965 15395
rect 995 15365 1045 15395
rect 1075 15365 1125 15395
rect 1155 15365 1205 15395
rect 1235 15365 1285 15395
rect 1315 15365 1365 15395
rect 1395 15365 1445 15395
rect 1475 15365 1525 15395
rect 1555 15365 1605 15395
rect 1635 15365 1685 15395
rect 1715 15365 1765 15395
rect 1795 15365 1845 15395
rect 1875 15365 1925 15395
rect 1955 15365 2005 15395
rect 2035 15365 2085 15395
rect 2115 15365 2165 15395
rect 2195 15365 2245 15395
rect 2275 15365 2325 15395
rect 2355 15365 2405 15395
rect 2435 15365 2485 15395
rect 2515 15365 2565 15395
rect 2595 15365 2645 15395
rect 2675 15365 2725 15395
rect 2755 15365 2805 15395
rect 2835 15365 2885 15395
rect 2915 15365 2965 15395
rect 2995 15365 3045 15395
rect 3075 15365 3125 15395
rect 3155 15365 3205 15395
rect 3235 15365 3285 15395
rect 3315 15365 3365 15395
rect 3395 15365 3445 15395
rect 3475 15365 3525 15395
rect 3555 15365 3605 15395
rect 3635 15365 3685 15395
rect 3715 15365 3765 15395
rect 3795 15365 3845 15395
rect 3875 15365 3925 15395
rect 3955 15365 4005 15395
rect 4035 15365 4085 15395
rect 4115 15365 4165 15395
rect 4195 15365 4725 15395
rect 4755 15365 4885 15395
rect 4915 15365 5045 15395
rect 5075 15365 5205 15395
rect 5235 15365 5365 15395
rect 5395 15365 5525 15395
rect 5555 15365 5685 15395
rect 5715 15365 6245 15395
rect 6275 15365 6325 15395
rect 6355 15365 6405 15395
rect 6435 15365 6485 15395
rect 6515 15365 6565 15395
rect 6595 15365 6645 15395
rect 6675 15365 6725 15395
rect 6755 15365 6805 15395
rect 6835 15365 6885 15395
rect 6915 15365 6965 15395
rect 6995 15365 7045 15395
rect 7075 15365 7125 15395
rect 7155 15365 7205 15395
rect 7235 15365 7285 15395
rect 7315 15365 7365 15395
rect 7395 15365 7445 15395
rect 7475 15365 7525 15395
rect 7555 15365 7605 15395
rect 7635 15365 7685 15395
rect 7715 15365 7765 15395
rect 7795 15365 7845 15395
rect 7875 15365 7925 15395
rect 7955 15365 8005 15395
rect 8035 15365 8085 15395
rect 8115 15365 8165 15395
rect 8195 15365 8245 15395
rect 8275 15365 8325 15395
rect 8355 15365 8405 15395
rect 8435 15365 8485 15395
rect 8515 15365 8565 15395
rect 8595 15365 8645 15395
rect 8675 15365 8725 15395
rect 8755 15365 8805 15395
rect 8835 15365 8885 15395
rect 8915 15365 8965 15395
rect 8995 15365 9045 15395
rect 9075 15365 9125 15395
rect 9155 15365 9205 15395
rect 9235 15365 9285 15395
rect 9315 15365 9365 15395
rect 9395 15365 9445 15395
rect 9475 15365 10005 15395
rect 10035 15365 10165 15395
rect 10195 15365 10325 15395
rect 10355 15365 10485 15395
rect 10515 15365 10645 15395
rect 10675 15365 10805 15395
rect 10835 15365 10965 15395
rect 10995 15365 11565 15395
rect 11595 15365 11645 15395
rect 11675 15365 11725 15395
rect 11755 15365 11805 15395
rect 11835 15365 11885 15395
rect 11915 15365 11965 15395
rect 11995 15365 12045 15395
rect 12075 15365 12125 15395
rect 12155 15365 12205 15395
rect 12235 15365 12285 15395
rect 12315 15365 12365 15395
rect 12395 15365 12445 15395
rect 12475 15365 12525 15395
rect 12555 15365 12605 15395
rect 12635 15365 12685 15395
rect 12715 15365 12765 15395
rect 12795 15365 12845 15395
rect 12875 15365 12925 15395
rect 12955 15365 13005 15395
rect 13035 15365 13085 15395
rect 13115 15365 13165 15395
rect 13195 15365 13245 15395
rect 13275 15365 13325 15395
rect 13355 15365 13405 15395
rect 13435 15365 13485 15395
rect 13515 15365 13565 15395
rect 13595 15365 13645 15395
rect 13675 15365 13725 15395
rect 13755 15365 13805 15395
rect 13835 15365 13885 15395
rect 13915 15365 13965 15395
rect 13995 15365 14045 15395
rect 14075 15365 14125 15395
rect 14155 15365 14205 15395
rect 14235 15365 14285 15395
rect 14315 15365 14365 15395
rect 14395 15365 14445 15395
rect 14475 15365 14525 15395
rect 14555 15365 14605 15395
rect 14635 15365 14685 15395
rect 14715 15365 15245 15395
rect 15275 15365 15405 15395
rect 15435 15365 15565 15395
rect 15595 15365 15725 15395
rect 15755 15365 15885 15395
rect 15915 15365 16045 15395
rect 16075 15365 16205 15395
rect 16235 15365 16765 15395
rect 16795 15365 16845 15395
rect 16875 15365 16925 15395
rect 16955 15365 17005 15395
rect 17035 15365 17085 15395
rect 17115 15365 17165 15395
rect 17195 15365 17245 15395
rect 17275 15365 17325 15395
rect 17355 15365 17405 15395
rect 17435 15365 17485 15395
rect 17515 15365 17565 15395
rect 17595 15365 17645 15395
rect 17675 15365 17725 15395
rect 17755 15365 17805 15395
rect 17835 15365 17885 15395
rect 17915 15365 17965 15395
rect 17995 15365 18045 15395
rect 18075 15365 18125 15395
rect 18155 15365 18205 15395
rect 18235 15365 18285 15395
rect 18315 15365 18365 15395
rect 18395 15365 18445 15395
rect 18475 15365 18525 15395
rect 18555 15365 18605 15395
rect 18635 15365 18685 15395
rect 18715 15365 18765 15395
rect 18795 15365 18845 15395
rect 18875 15365 18925 15395
rect 18955 15365 19005 15395
rect 19035 15365 19085 15395
rect 19115 15365 19165 15395
rect 19195 15365 19245 15395
rect 19275 15365 19325 15395
rect 19355 15365 19405 15395
rect 19435 15365 19485 15395
rect 19515 15365 19565 15395
rect 19595 15365 19645 15395
rect 19675 15365 19725 15395
rect 19755 15365 19805 15395
rect 19835 15365 19885 15395
rect 19915 15365 19965 15395
rect 19995 15365 20045 15395
rect 20075 15365 20125 15395
rect 20155 15365 20205 15395
rect 20235 15365 20285 15395
rect 20315 15365 20365 15395
rect 20395 15365 20445 15395
rect 20475 15365 20525 15395
rect 20555 15365 20605 15395
rect 20635 15365 20685 15395
rect 20715 15365 20765 15395
rect 20795 15365 20845 15395
rect 20875 15365 20925 15395
rect 20955 15365 20960 15395
rect 0 15360 20960 15365
rect 0 15315 20960 15320
rect 0 15285 5605 15315
rect 5635 15285 10885 15315
rect 10915 15285 15325 15315
rect 15355 15285 20960 15315
rect 0 15280 20960 15285
rect 0 15235 20960 15240
rect 0 15205 5 15235
rect 35 15205 85 15235
rect 115 15205 165 15235
rect 195 15205 245 15235
rect 275 15205 325 15235
rect 355 15205 405 15235
rect 435 15205 485 15235
rect 515 15205 565 15235
rect 595 15205 645 15235
rect 675 15205 725 15235
rect 755 15205 805 15235
rect 835 15205 885 15235
rect 915 15205 965 15235
rect 995 15205 1045 15235
rect 1075 15205 1125 15235
rect 1155 15205 1205 15235
rect 1235 15205 1285 15235
rect 1315 15205 1365 15235
rect 1395 15205 1445 15235
rect 1475 15205 1525 15235
rect 1555 15205 1605 15235
rect 1635 15205 1685 15235
rect 1715 15205 1765 15235
rect 1795 15205 1845 15235
rect 1875 15205 1925 15235
rect 1955 15205 2005 15235
rect 2035 15205 2085 15235
rect 2115 15205 2165 15235
rect 2195 15205 2245 15235
rect 2275 15205 2325 15235
rect 2355 15205 2405 15235
rect 2435 15205 2485 15235
rect 2515 15205 2565 15235
rect 2595 15205 2645 15235
rect 2675 15205 2725 15235
rect 2755 15205 2805 15235
rect 2835 15205 2885 15235
rect 2915 15205 2965 15235
rect 2995 15205 3045 15235
rect 3075 15205 3125 15235
rect 3155 15205 3205 15235
rect 3235 15205 3285 15235
rect 3315 15205 3365 15235
rect 3395 15205 3445 15235
rect 3475 15205 3525 15235
rect 3555 15205 3605 15235
rect 3635 15205 3685 15235
rect 3715 15205 3765 15235
rect 3795 15205 3845 15235
rect 3875 15205 3925 15235
rect 3955 15205 4005 15235
rect 4035 15205 4085 15235
rect 4115 15205 4165 15235
rect 4195 15205 4725 15235
rect 4755 15205 4885 15235
rect 4915 15205 5045 15235
rect 5075 15205 5205 15235
rect 5235 15205 5365 15235
rect 5395 15205 5525 15235
rect 5555 15205 5685 15235
rect 5715 15205 6245 15235
rect 6275 15205 6325 15235
rect 6355 15205 6405 15235
rect 6435 15205 6485 15235
rect 6515 15205 6565 15235
rect 6595 15205 6645 15235
rect 6675 15205 6725 15235
rect 6755 15205 6805 15235
rect 6835 15205 6885 15235
rect 6915 15205 6965 15235
rect 6995 15205 7045 15235
rect 7075 15205 7125 15235
rect 7155 15205 7205 15235
rect 7235 15205 7285 15235
rect 7315 15205 7365 15235
rect 7395 15205 7445 15235
rect 7475 15205 7525 15235
rect 7555 15205 7605 15235
rect 7635 15205 7685 15235
rect 7715 15205 7765 15235
rect 7795 15205 7845 15235
rect 7875 15205 7925 15235
rect 7955 15205 8005 15235
rect 8035 15205 8085 15235
rect 8115 15205 8165 15235
rect 8195 15205 8245 15235
rect 8275 15205 8325 15235
rect 8355 15205 8405 15235
rect 8435 15205 8485 15235
rect 8515 15205 8565 15235
rect 8595 15205 8645 15235
rect 8675 15205 8725 15235
rect 8755 15205 8805 15235
rect 8835 15205 8885 15235
rect 8915 15205 8965 15235
rect 8995 15205 9045 15235
rect 9075 15205 9125 15235
rect 9155 15205 9205 15235
rect 9235 15205 9285 15235
rect 9315 15205 9365 15235
rect 9395 15205 9445 15235
rect 9475 15205 10005 15235
rect 10035 15205 10165 15235
rect 10195 15205 10325 15235
rect 10355 15205 10485 15235
rect 10515 15205 10645 15235
rect 10675 15205 10805 15235
rect 10835 15205 10965 15235
rect 10995 15205 11565 15235
rect 11595 15205 11645 15235
rect 11675 15205 11725 15235
rect 11755 15205 11805 15235
rect 11835 15205 11885 15235
rect 11915 15205 11965 15235
rect 11995 15205 12045 15235
rect 12075 15205 12125 15235
rect 12155 15205 12205 15235
rect 12235 15205 12285 15235
rect 12315 15205 12365 15235
rect 12395 15205 12445 15235
rect 12475 15205 12525 15235
rect 12555 15205 12605 15235
rect 12635 15205 12685 15235
rect 12715 15205 12765 15235
rect 12795 15205 12845 15235
rect 12875 15205 12925 15235
rect 12955 15205 13005 15235
rect 13035 15205 13085 15235
rect 13115 15205 13165 15235
rect 13195 15205 13245 15235
rect 13275 15205 13325 15235
rect 13355 15205 13405 15235
rect 13435 15205 13485 15235
rect 13515 15205 13565 15235
rect 13595 15205 13645 15235
rect 13675 15205 13725 15235
rect 13755 15205 13805 15235
rect 13835 15205 13885 15235
rect 13915 15205 13965 15235
rect 13995 15205 14045 15235
rect 14075 15205 14125 15235
rect 14155 15205 14205 15235
rect 14235 15205 14285 15235
rect 14315 15205 14365 15235
rect 14395 15205 14445 15235
rect 14475 15205 14525 15235
rect 14555 15205 14605 15235
rect 14635 15205 14685 15235
rect 14715 15205 15245 15235
rect 15275 15205 15405 15235
rect 15435 15205 15565 15235
rect 15595 15205 15725 15235
rect 15755 15205 15885 15235
rect 15915 15205 16045 15235
rect 16075 15205 16205 15235
rect 16235 15205 16765 15235
rect 16795 15205 16845 15235
rect 16875 15205 16925 15235
rect 16955 15205 17005 15235
rect 17035 15205 17085 15235
rect 17115 15205 17165 15235
rect 17195 15205 17245 15235
rect 17275 15205 17325 15235
rect 17355 15205 17405 15235
rect 17435 15205 17485 15235
rect 17515 15205 17565 15235
rect 17595 15205 17645 15235
rect 17675 15205 17725 15235
rect 17755 15205 17805 15235
rect 17835 15205 17885 15235
rect 17915 15205 17965 15235
rect 17995 15205 18045 15235
rect 18075 15205 18125 15235
rect 18155 15205 18205 15235
rect 18235 15205 18285 15235
rect 18315 15205 18365 15235
rect 18395 15205 18445 15235
rect 18475 15205 18525 15235
rect 18555 15205 18605 15235
rect 18635 15205 18685 15235
rect 18715 15205 18765 15235
rect 18795 15205 18845 15235
rect 18875 15205 18925 15235
rect 18955 15205 19005 15235
rect 19035 15205 19085 15235
rect 19115 15205 19165 15235
rect 19195 15205 19245 15235
rect 19275 15205 19325 15235
rect 19355 15205 19405 15235
rect 19435 15205 19485 15235
rect 19515 15205 19565 15235
rect 19595 15205 19645 15235
rect 19675 15205 19725 15235
rect 19755 15205 19805 15235
rect 19835 15205 19885 15235
rect 19915 15205 19965 15235
rect 19995 15205 20045 15235
rect 20075 15205 20125 15235
rect 20155 15205 20205 15235
rect 20235 15205 20285 15235
rect 20315 15205 20365 15235
rect 20395 15205 20445 15235
rect 20475 15205 20525 15235
rect 20555 15205 20605 15235
rect 20635 15205 20685 15235
rect 20715 15205 20765 15235
rect 20795 15205 20845 15235
rect 20875 15205 20925 15235
rect 20955 15205 20960 15235
rect 0 15200 20960 15205
rect 0 15155 20960 15160
rect 0 15125 5 15155
rect 35 15125 85 15155
rect 115 15125 165 15155
rect 195 15125 245 15155
rect 275 15125 325 15155
rect 355 15125 405 15155
rect 435 15125 485 15155
rect 515 15125 565 15155
rect 595 15125 645 15155
rect 675 15125 725 15155
rect 755 15125 805 15155
rect 835 15125 885 15155
rect 915 15125 965 15155
rect 995 15125 1045 15155
rect 1075 15125 1125 15155
rect 1155 15125 1205 15155
rect 1235 15125 1285 15155
rect 1315 15125 1365 15155
rect 1395 15125 1445 15155
rect 1475 15125 1525 15155
rect 1555 15125 1605 15155
rect 1635 15125 1685 15155
rect 1715 15125 1765 15155
rect 1795 15125 1845 15155
rect 1875 15125 1925 15155
rect 1955 15125 2005 15155
rect 2035 15125 2085 15155
rect 2115 15125 2165 15155
rect 2195 15125 2245 15155
rect 2275 15125 2325 15155
rect 2355 15125 2405 15155
rect 2435 15125 2485 15155
rect 2515 15125 2565 15155
rect 2595 15125 2645 15155
rect 2675 15125 2725 15155
rect 2755 15125 2805 15155
rect 2835 15125 2885 15155
rect 2915 15125 2965 15155
rect 2995 15125 3045 15155
rect 3075 15125 3125 15155
rect 3155 15125 3205 15155
rect 3235 15125 3285 15155
rect 3315 15125 3365 15155
rect 3395 15125 3445 15155
rect 3475 15125 3525 15155
rect 3555 15125 3605 15155
rect 3635 15125 3685 15155
rect 3715 15125 3765 15155
rect 3795 15125 3845 15155
rect 3875 15125 3925 15155
rect 3955 15125 4005 15155
rect 4035 15125 4085 15155
rect 4115 15125 4165 15155
rect 4195 15125 5765 15155
rect 5795 15125 5925 15155
rect 5955 15125 6245 15155
rect 6275 15125 6325 15155
rect 6355 15125 6405 15155
rect 6435 15125 6485 15155
rect 6515 15125 6565 15155
rect 6595 15125 6645 15155
rect 6675 15125 6725 15155
rect 6755 15125 6805 15155
rect 6835 15125 6885 15155
rect 6915 15125 6965 15155
rect 6995 15125 7045 15155
rect 7075 15125 7125 15155
rect 7155 15125 7205 15155
rect 7235 15125 7285 15155
rect 7315 15125 7365 15155
rect 7395 15125 7445 15155
rect 7475 15125 7525 15155
rect 7555 15125 7605 15155
rect 7635 15125 7685 15155
rect 7715 15125 7765 15155
rect 7795 15125 7845 15155
rect 7875 15125 7925 15155
rect 7955 15125 8005 15155
rect 8035 15125 8085 15155
rect 8115 15125 8165 15155
rect 8195 15125 8245 15155
rect 8275 15125 8325 15155
rect 8355 15125 8405 15155
rect 8435 15125 8485 15155
rect 8515 15125 8565 15155
rect 8595 15125 8645 15155
rect 8675 15125 8725 15155
rect 8755 15125 8805 15155
rect 8835 15125 8885 15155
rect 8915 15125 8965 15155
rect 8995 15125 9045 15155
rect 9075 15125 9125 15155
rect 9155 15125 9205 15155
rect 9235 15125 9285 15155
rect 9315 15125 9365 15155
rect 9395 15125 9445 15155
rect 9475 15125 11045 15155
rect 11075 15125 11205 15155
rect 11235 15125 11565 15155
rect 11595 15125 11645 15155
rect 11675 15125 11725 15155
rect 11755 15125 11805 15155
rect 11835 15125 11885 15155
rect 11915 15125 11965 15155
rect 11995 15125 12045 15155
rect 12075 15125 12125 15155
rect 12155 15125 12205 15155
rect 12235 15125 12285 15155
rect 12315 15125 12365 15155
rect 12395 15125 12445 15155
rect 12475 15125 12525 15155
rect 12555 15125 12605 15155
rect 12635 15125 12685 15155
rect 12715 15125 12765 15155
rect 12795 15125 12845 15155
rect 12875 15125 12925 15155
rect 12955 15125 13005 15155
rect 13035 15125 13085 15155
rect 13115 15125 13165 15155
rect 13195 15125 13245 15155
rect 13275 15125 13325 15155
rect 13355 15125 13405 15155
rect 13435 15125 13485 15155
rect 13515 15125 13565 15155
rect 13595 15125 13645 15155
rect 13675 15125 13725 15155
rect 13755 15125 13805 15155
rect 13835 15125 13885 15155
rect 13915 15125 13965 15155
rect 13995 15125 14045 15155
rect 14075 15125 14125 15155
rect 14155 15125 14205 15155
rect 14235 15125 14285 15155
rect 14315 15125 14365 15155
rect 14395 15125 14445 15155
rect 14475 15125 14525 15155
rect 14555 15125 14605 15155
rect 14635 15125 14685 15155
rect 14715 15125 15005 15155
rect 15035 15125 15165 15155
rect 15195 15125 16765 15155
rect 16795 15125 16845 15155
rect 16875 15125 16925 15155
rect 16955 15125 17005 15155
rect 17035 15125 17085 15155
rect 17115 15125 17165 15155
rect 17195 15125 17245 15155
rect 17275 15125 17325 15155
rect 17355 15125 17405 15155
rect 17435 15125 17485 15155
rect 17515 15125 17565 15155
rect 17595 15125 17645 15155
rect 17675 15125 17725 15155
rect 17755 15125 17805 15155
rect 17835 15125 17885 15155
rect 17915 15125 17965 15155
rect 17995 15125 18045 15155
rect 18075 15125 18125 15155
rect 18155 15125 18205 15155
rect 18235 15125 18285 15155
rect 18315 15125 18365 15155
rect 18395 15125 18445 15155
rect 18475 15125 18525 15155
rect 18555 15125 18605 15155
rect 18635 15125 18685 15155
rect 18715 15125 18765 15155
rect 18795 15125 18845 15155
rect 18875 15125 18925 15155
rect 18955 15125 19005 15155
rect 19035 15125 19085 15155
rect 19115 15125 19165 15155
rect 19195 15125 19245 15155
rect 19275 15125 19325 15155
rect 19355 15125 19405 15155
rect 19435 15125 19485 15155
rect 19515 15125 19565 15155
rect 19595 15125 19645 15155
rect 19675 15125 19725 15155
rect 19755 15125 19805 15155
rect 19835 15125 19885 15155
rect 19915 15125 19965 15155
rect 19995 15125 20045 15155
rect 20075 15125 20125 15155
rect 20155 15125 20205 15155
rect 20235 15125 20285 15155
rect 20315 15125 20365 15155
rect 20395 15125 20445 15155
rect 20475 15125 20525 15155
rect 20555 15125 20605 15155
rect 20635 15125 20685 15155
rect 20715 15125 20765 15155
rect 20795 15125 20845 15155
rect 20875 15125 20925 15155
rect 20955 15125 20960 15155
rect 0 15120 20960 15125
rect 0 15075 20960 15080
rect 0 15045 5845 15075
rect 5875 15045 11125 15075
rect 11155 15045 15085 15075
rect 15115 15045 20960 15075
rect 0 15040 20960 15045
rect 0 14995 20960 15000
rect 0 14965 5 14995
rect 35 14965 85 14995
rect 115 14965 165 14995
rect 195 14965 245 14995
rect 275 14965 325 14995
rect 355 14965 405 14995
rect 435 14965 485 14995
rect 515 14965 565 14995
rect 595 14965 645 14995
rect 675 14965 725 14995
rect 755 14965 805 14995
rect 835 14965 885 14995
rect 915 14965 965 14995
rect 995 14965 1045 14995
rect 1075 14965 1125 14995
rect 1155 14965 1205 14995
rect 1235 14965 1285 14995
rect 1315 14965 1365 14995
rect 1395 14965 1445 14995
rect 1475 14965 1525 14995
rect 1555 14965 1605 14995
rect 1635 14965 1685 14995
rect 1715 14965 1765 14995
rect 1795 14965 1845 14995
rect 1875 14965 1925 14995
rect 1955 14965 2005 14995
rect 2035 14965 2085 14995
rect 2115 14965 2165 14995
rect 2195 14965 2245 14995
rect 2275 14965 2325 14995
rect 2355 14965 2405 14995
rect 2435 14965 2485 14995
rect 2515 14965 2565 14995
rect 2595 14965 2645 14995
rect 2675 14965 2725 14995
rect 2755 14965 2805 14995
rect 2835 14965 2885 14995
rect 2915 14965 2965 14995
rect 2995 14965 3045 14995
rect 3075 14965 3125 14995
rect 3155 14965 3205 14995
rect 3235 14965 3285 14995
rect 3315 14965 3365 14995
rect 3395 14965 3445 14995
rect 3475 14965 3525 14995
rect 3555 14965 3605 14995
rect 3635 14965 3685 14995
rect 3715 14965 3765 14995
rect 3795 14965 3845 14995
rect 3875 14965 3925 14995
rect 3955 14965 4005 14995
rect 4035 14965 4085 14995
rect 4115 14965 4165 14995
rect 4195 14965 5765 14995
rect 5795 14965 5925 14995
rect 5955 14965 6245 14995
rect 6275 14965 6325 14995
rect 6355 14965 6405 14995
rect 6435 14965 6485 14995
rect 6515 14965 6565 14995
rect 6595 14965 6645 14995
rect 6675 14965 6725 14995
rect 6755 14965 6805 14995
rect 6835 14965 6885 14995
rect 6915 14965 6965 14995
rect 6995 14965 7045 14995
rect 7075 14965 7125 14995
rect 7155 14965 7205 14995
rect 7235 14965 7285 14995
rect 7315 14965 7365 14995
rect 7395 14965 7445 14995
rect 7475 14965 7525 14995
rect 7555 14965 7605 14995
rect 7635 14965 7685 14995
rect 7715 14965 7765 14995
rect 7795 14965 7845 14995
rect 7875 14965 7925 14995
rect 7955 14965 8005 14995
rect 8035 14965 8085 14995
rect 8115 14965 8165 14995
rect 8195 14965 8245 14995
rect 8275 14965 8325 14995
rect 8355 14965 8405 14995
rect 8435 14965 8485 14995
rect 8515 14965 8565 14995
rect 8595 14965 8645 14995
rect 8675 14965 8725 14995
rect 8755 14965 8805 14995
rect 8835 14965 8885 14995
rect 8915 14965 8965 14995
rect 8995 14965 9045 14995
rect 9075 14965 9125 14995
rect 9155 14965 9205 14995
rect 9235 14965 9285 14995
rect 9315 14965 9365 14995
rect 9395 14965 9445 14995
rect 9475 14965 11045 14995
rect 11075 14965 11205 14995
rect 11235 14965 11565 14995
rect 11595 14965 11645 14995
rect 11675 14965 11725 14995
rect 11755 14965 11805 14995
rect 11835 14965 11885 14995
rect 11915 14965 11965 14995
rect 11995 14965 12045 14995
rect 12075 14965 12125 14995
rect 12155 14965 12205 14995
rect 12235 14965 12285 14995
rect 12315 14965 12365 14995
rect 12395 14965 12445 14995
rect 12475 14965 12525 14995
rect 12555 14965 12605 14995
rect 12635 14965 12685 14995
rect 12715 14965 12765 14995
rect 12795 14965 12845 14995
rect 12875 14965 12925 14995
rect 12955 14965 13005 14995
rect 13035 14965 13085 14995
rect 13115 14965 13165 14995
rect 13195 14965 13245 14995
rect 13275 14965 13325 14995
rect 13355 14965 13405 14995
rect 13435 14965 13485 14995
rect 13515 14965 13565 14995
rect 13595 14965 13645 14995
rect 13675 14965 13725 14995
rect 13755 14965 13805 14995
rect 13835 14965 13885 14995
rect 13915 14965 13965 14995
rect 13995 14965 14045 14995
rect 14075 14965 14125 14995
rect 14155 14965 14205 14995
rect 14235 14965 14285 14995
rect 14315 14965 14365 14995
rect 14395 14965 14445 14995
rect 14475 14965 14525 14995
rect 14555 14965 14605 14995
rect 14635 14965 14685 14995
rect 14715 14965 15005 14995
rect 15035 14965 15165 14995
rect 15195 14965 16765 14995
rect 16795 14965 16845 14995
rect 16875 14965 16925 14995
rect 16955 14965 17005 14995
rect 17035 14965 17085 14995
rect 17115 14965 17165 14995
rect 17195 14965 17245 14995
rect 17275 14965 17325 14995
rect 17355 14965 17405 14995
rect 17435 14965 17485 14995
rect 17515 14965 17565 14995
rect 17595 14965 17645 14995
rect 17675 14965 17725 14995
rect 17755 14965 17805 14995
rect 17835 14965 17885 14995
rect 17915 14965 17965 14995
rect 17995 14965 18045 14995
rect 18075 14965 18125 14995
rect 18155 14965 18205 14995
rect 18235 14965 18285 14995
rect 18315 14965 18365 14995
rect 18395 14965 18445 14995
rect 18475 14965 18525 14995
rect 18555 14965 18605 14995
rect 18635 14965 18685 14995
rect 18715 14965 18765 14995
rect 18795 14965 18845 14995
rect 18875 14965 18925 14995
rect 18955 14965 19005 14995
rect 19035 14965 19085 14995
rect 19115 14965 19165 14995
rect 19195 14965 19245 14995
rect 19275 14965 19325 14995
rect 19355 14965 19405 14995
rect 19435 14965 19485 14995
rect 19515 14965 19565 14995
rect 19595 14965 19645 14995
rect 19675 14965 19725 14995
rect 19755 14965 19805 14995
rect 19835 14965 19885 14995
rect 19915 14965 19965 14995
rect 19995 14965 20045 14995
rect 20075 14965 20125 14995
rect 20155 14965 20205 14995
rect 20235 14965 20285 14995
rect 20315 14965 20365 14995
rect 20395 14965 20445 14995
rect 20475 14965 20525 14995
rect 20555 14965 20605 14995
rect 20635 14965 20685 14995
rect 20715 14965 20765 14995
rect 20795 14965 20845 14995
rect 20875 14965 20925 14995
rect 20955 14965 20960 14995
rect 0 14960 20960 14965
rect 0 14915 20960 14920
rect 0 14885 5 14915
rect 35 14885 85 14915
rect 115 14885 165 14915
rect 195 14885 245 14915
rect 275 14885 325 14915
rect 355 14885 405 14915
rect 435 14885 485 14915
rect 515 14885 565 14915
rect 595 14885 645 14915
rect 675 14885 725 14915
rect 755 14885 805 14915
rect 835 14885 885 14915
rect 915 14885 965 14915
rect 995 14885 1045 14915
rect 1075 14885 1125 14915
rect 1155 14885 1205 14915
rect 1235 14885 1285 14915
rect 1315 14885 1365 14915
rect 1395 14885 1445 14915
rect 1475 14885 1525 14915
rect 1555 14885 1605 14915
rect 1635 14885 1685 14915
rect 1715 14885 1765 14915
rect 1795 14885 1845 14915
rect 1875 14885 1925 14915
rect 1955 14885 2005 14915
rect 2035 14885 2085 14915
rect 2115 14885 2165 14915
rect 2195 14885 2245 14915
rect 2275 14885 2325 14915
rect 2355 14885 2405 14915
rect 2435 14885 2485 14915
rect 2515 14885 2565 14915
rect 2595 14885 2645 14915
rect 2675 14885 2725 14915
rect 2755 14885 2805 14915
rect 2835 14885 2885 14915
rect 2915 14885 2965 14915
rect 2995 14885 3045 14915
rect 3075 14885 3125 14915
rect 3155 14885 3205 14915
rect 3235 14885 3285 14915
rect 3315 14885 3365 14915
rect 3395 14885 3445 14915
rect 3475 14885 3525 14915
rect 3555 14885 3605 14915
rect 3635 14885 3685 14915
rect 3715 14885 3765 14915
rect 3795 14885 3845 14915
rect 3875 14885 3925 14915
rect 3955 14885 4005 14915
rect 4035 14885 4085 14915
rect 4115 14885 4165 14915
rect 4195 14885 6005 14915
rect 6035 14885 6165 14915
rect 6195 14885 6245 14915
rect 6275 14885 6325 14915
rect 6355 14885 6405 14915
rect 6435 14885 6485 14915
rect 6515 14885 6565 14915
rect 6595 14885 6645 14915
rect 6675 14885 6725 14915
rect 6755 14885 6805 14915
rect 6835 14885 6885 14915
rect 6915 14885 6965 14915
rect 6995 14885 7045 14915
rect 7075 14885 7125 14915
rect 7155 14885 7205 14915
rect 7235 14885 7285 14915
rect 7315 14885 7365 14915
rect 7395 14885 7445 14915
rect 7475 14885 7525 14915
rect 7555 14885 7605 14915
rect 7635 14885 7685 14915
rect 7715 14885 7765 14915
rect 7795 14885 7845 14915
rect 7875 14885 7925 14915
rect 7955 14885 8005 14915
rect 8035 14885 8085 14915
rect 8115 14885 8165 14915
rect 8195 14885 8245 14915
rect 8275 14885 8325 14915
rect 8355 14885 8405 14915
rect 8435 14885 8485 14915
rect 8515 14885 8565 14915
rect 8595 14885 8645 14915
rect 8675 14885 8725 14915
rect 8755 14885 8805 14915
rect 8835 14885 8885 14915
rect 8915 14885 8965 14915
rect 8995 14885 9045 14915
rect 9075 14885 9125 14915
rect 9155 14885 9205 14915
rect 9235 14885 9285 14915
rect 9315 14885 9365 14915
rect 9395 14885 9445 14915
rect 9475 14885 11285 14915
rect 11315 14885 11445 14915
rect 11475 14885 11565 14915
rect 11595 14885 11645 14915
rect 11675 14885 11725 14915
rect 11755 14885 11805 14915
rect 11835 14885 11885 14915
rect 11915 14885 11965 14915
rect 11995 14885 12045 14915
rect 12075 14885 12125 14915
rect 12155 14885 12205 14915
rect 12235 14885 12285 14915
rect 12315 14885 12365 14915
rect 12395 14885 12445 14915
rect 12475 14885 12525 14915
rect 12555 14885 12605 14915
rect 12635 14885 12685 14915
rect 12715 14885 12765 14915
rect 12795 14885 12845 14915
rect 12875 14885 12925 14915
rect 12955 14885 13005 14915
rect 13035 14885 13085 14915
rect 13115 14885 13165 14915
rect 13195 14885 13245 14915
rect 13275 14885 13325 14915
rect 13355 14885 13405 14915
rect 13435 14885 13485 14915
rect 13515 14885 13565 14915
rect 13595 14885 13645 14915
rect 13675 14885 13725 14915
rect 13755 14885 13805 14915
rect 13835 14885 13885 14915
rect 13915 14885 13965 14915
rect 13995 14885 14045 14915
rect 14075 14885 14125 14915
rect 14155 14885 14205 14915
rect 14235 14885 14285 14915
rect 14315 14885 14365 14915
rect 14395 14885 14445 14915
rect 14475 14885 14525 14915
rect 14555 14885 14605 14915
rect 14635 14885 14685 14915
rect 14715 14885 14765 14915
rect 14795 14885 14925 14915
rect 14955 14885 16765 14915
rect 16795 14885 16845 14915
rect 16875 14885 16925 14915
rect 16955 14885 17005 14915
rect 17035 14885 17085 14915
rect 17115 14885 17165 14915
rect 17195 14885 17245 14915
rect 17275 14885 17325 14915
rect 17355 14885 17405 14915
rect 17435 14885 17485 14915
rect 17515 14885 17565 14915
rect 17595 14885 17645 14915
rect 17675 14885 17725 14915
rect 17755 14885 17805 14915
rect 17835 14885 17885 14915
rect 17915 14885 17965 14915
rect 17995 14885 18045 14915
rect 18075 14885 18125 14915
rect 18155 14885 18205 14915
rect 18235 14885 18285 14915
rect 18315 14885 18365 14915
rect 18395 14885 18445 14915
rect 18475 14885 18525 14915
rect 18555 14885 18605 14915
rect 18635 14885 18685 14915
rect 18715 14885 18765 14915
rect 18795 14885 18845 14915
rect 18875 14885 18925 14915
rect 18955 14885 19005 14915
rect 19035 14885 19085 14915
rect 19115 14885 19165 14915
rect 19195 14885 19245 14915
rect 19275 14885 19325 14915
rect 19355 14885 19405 14915
rect 19435 14885 19485 14915
rect 19515 14885 19565 14915
rect 19595 14885 19645 14915
rect 19675 14885 19725 14915
rect 19755 14885 19805 14915
rect 19835 14885 19885 14915
rect 19915 14885 19965 14915
rect 19995 14885 20045 14915
rect 20075 14885 20125 14915
rect 20155 14885 20205 14915
rect 20235 14885 20285 14915
rect 20315 14885 20365 14915
rect 20395 14885 20445 14915
rect 20475 14885 20525 14915
rect 20555 14885 20605 14915
rect 20635 14885 20685 14915
rect 20715 14885 20765 14915
rect 20795 14885 20845 14915
rect 20875 14885 20925 14915
rect 20955 14885 20960 14915
rect 0 14880 20960 14885
rect 0 14835 20960 14840
rect 0 14805 6085 14835
rect 6115 14805 11365 14835
rect 11395 14805 14845 14835
rect 14875 14805 20960 14835
rect 0 14800 20960 14805
rect 0 14755 20960 14760
rect 0 14725 5 14755
rect 35 14725 85 14755
rect 115 14725 165 14755
rect 195 14725 245 14755
rect 275 14725 325 14755
rect 355 14725 405 14755
rect 435 14725 485 14755
rect 515 14725 565 14755
rect 595 14725 645 14755
rect 675 14725 725 14755
rect 755 14725 805 14755
rect 835 14725 885 14755
rect 915 14725 965 14755
rect 995 14725 1045 14755
rect 1075 14725 1125 14755
rect 1155 14725 1205 14755
rect 1235 14725 1285 14755
rect 1315 14725 1365 14755
rect 1395 14725 1445 14755
rect 1475 14725 1525 14755
rect 1555 14725 1605 14755
rect 1635 14725 1685 14755
rect 1715 14725 1765 14755
rect 1795 14725 1845 14755
rect 1875 14725 1925 14755
rect 1955 14725 2005 14755
rect 2035 14725 2085 14755
rect 2115 14725 2165 14755
rect 2195 14725 2245 14755
rect 2275 14725 2325 14755
rect 2355 14725 2405 14755
rect 2435 14725 2485 14755
rect 2515 14725 2565 14755
rect 2595 14725 2645 14755
rect 2675 14725 2725 14755
rect 2755 14725 2805 14755
rect 2835 14725 2885 14755
rect 2915 14725 2965 14755
rect 2995 14725 3045 14755
rect 3075 14725 3125 14755
rect 3155 14725 3205 14755
rect 3235 14725 3285 14755
rect 3315 14725 3365 14755
rect 3395 14725 3445 14755
rect 3475 14725 3525 14755
rect 3555 14725 3605 14755
rect 3635 14725 3685 14755
rect 3715 14725 3765 14755
rect 3795 14725 3845 14755
rect 3875 14725 3925 14755
rect 3955 14725 4005 14755
rect 4035 14725 4085 14755
rect 4115 14725 4165 14755
rect 4195 14725 6005 14755
rect 6035 14725 6165 14755
rect 6195 14725 6245 14755
rect 6275 14725 6325 14755
rect 6355 14725 6405 14755
rect 6435 14725 6485 14755
rect 6515 14725 6565 14755
rect 6595 14725 6645 14755
rect 6675 14725 6725 14755
rect 6755 14725 6805 14755
rect 6835 14725 6885 14755
rect 6915 14725 6965 14755
rect 6995 14725 7045 14755
rect 7075 14725 7125 14755
rect 7155 14725 7205 14755
rect 7235 14725 7285 14755
rect 7315 14725 7365 14755
rect 7395 14725 7445 14755
rect 7475 14725 7525 14755
rect 7555 14725 7605 14755
rect 7635 14725 7685 14755
rect 7715 14725 7765 14755
rect 7795 14725 7845 14755
rect 7875 14725 7925 14755
rect 7955 14725 8005 14755
rect 8035 14725 8085 14755
rect 8115 14725 8165 14755
rect 8195 14725 8245 14755
rect 8275 14725 8325 14755
rect 8355 14725 8405 14755
rect 8435 14725 8485 14755
rect 8515 14725 8565 14755
rect 8595 14725 8645 14755
rect 8675 14725 8725 14755
rect 8755 14725 8805 14755
rect 8835 14725 8885 14755
rect 8915 14725 8965 14755
rect 8995 14725 9045 14755
rect 9075 14725 9125 14755
rect 9155 14725 9205 14755
rect 9235 14725 9285 14755
rect 9315 14725 9365 14755
rect 9395 14725 9445 14755
rect 9475 14725 11285 14755
rect 11315 14725 11445 14755
rect 11475 14725 11565 14755
rect 11595 14725 11645 14755
rect 11675 14725 11725 14755
rect 11755 14725 11805 14755
rect 11835 14725 11885 14755
rect 11915 14725 11965 14755
rect 11995 14725 12045 14755
rect 12075 14725 12125 14755
rect 12155 14725 12205 14755
rect 12235 14725 12285 14755
rect 12315 14725 12365 14755
rect 12395 14725 12445 14755
rect 12475 14725 12525 14755
rect 12555 14725 12605 14755
rect 12635 14725 12685 14755
rect 12715 14725 12765 14755
rect 12795 14725 12845 14755
rect 12875 14725 12925 14755
rect 12955 14725 13005 14755
rect 13035 14725 13085 14755
rect 13115 14725 13165 14755
rect 13195 14725 13245 14755
rect 13275 14725 13325 14755
rect 13355 14725 13405 14755
rect 13435 14725 13485 14755
rect 13515 14725 13565 14755
rect 13595 14725 13645 14755
rect 13675 14725 13725 14755
rect 13755 14725 13805 14755
rect 13835 14725 13885 14755
rect 13915 14725 13965 14755
rect 13995 14725 14045 14755
rect 14075 14725 14125 14755
rect 14155 14725 14205 14755
rect 14235 14725 14285 14755
rect 14315 14725 14365 14755
rect 14395 14725 14445 14755
rect 14475 14725 14525 14755
rect 14555 14725 14605 14755
rect 14635 14725 14685 14755
rect 14715 14725 14765 14755
rect 14795 14725 14925 14755
rect 14955 14725 16765 14755
rect 16795 14725 16845 14755
rect 16875 14725 16925 14755
rect 16955 14725 17005 14755
rect 17035 14725 17085 14755
rect 17115 14725 17165 14755
rect 17195 14725 17245 14755
rect 17275 14725 17325 14755
rect 17355 14725 17405 14755
rect 17435 14725 17485 14755
rect 17515 14725 17565 14755
rect 17595 14725 17645 14755
rect 17675 14725 17725 14755
rect 17755 14725 17805 14755
rect 17835 14725 17885 14755
rect 17915 14725 17965 14755
rect 17995 14725 18045 14755
rect 18075 14725 18125 14755
rect 18155 14725 18205 14755
rect 18235 14725 18285 14755
rect 18315 14725 18365 14755
rect 18395 14725 18445 14755
rect 18475 14725 18525 14755
rect 18555 14725 18605 14755
rect 18635 14725 18685 14755
rect 18715 14725 18765 14755
rect 18795 14725 18845 14755
rect 18875 14725 18925 14755
rect 18955 14725 19005 14755
rect 19035 14725 19085 14755
rect 19115 14725 19165 14755
rect 19195 14725 19245 14755
rect 19275 14725 19325 14755
rect 19355 14725 19405 14755
rect 19435 14725 19485 14755
rect 19515 14725 19565 14755
rect 19595 14725 19645 14755
rect 19675 14725 19725 14755
rect 19755 14725 19805 14755
rect 19835 14725 19885 14755
rect 19915 14725 19965 14755
rect 19995 14725 20045 14755
rect 20075 14725 20125 14755
rect 20155 14725 20205 14755
rect 20235 14725 20285 14755
rect 20315 14725 20365 14755
rect 20395 14725 20445 14755
rect 20475 14725 20525 14755
rect 20555 14725 20605 14755
rect 20635 14725 20685 14755
rect 20715 14725 20765 14755
rect 20795 14725 20845 14755
rect 20875 14725 20925 14755
rect 20955 14725 20960 14755
rect 0 14720 20960 14725
<< via2 >>
rect 5 18645 35 18675
rect 85 18645 115 18675
rect 165 18645 195 18675
rect 245 18645 275 18675
rect 325 18645 355 18675
rect 405 18645 435 18675
rect 485 18645 515 18675
rect 565 18645 595 18675
rect 645 18645 675 18675
rect 725 18645 755 18675
rect 805 18645 835 18675
rect 885 18645 915 18675
rect 965 18645 995 18675
rect 1045 18645 1075 18675
rect 1125 18645 1155 18675
rect 1205 18645 1235 18675
rect 1285 18645 1315 18675
rect 1365 18645 1395 18675
rect 1445 18645 1475 18675
rect 1525 18645 1555 18675
rect 1605 18645 1635 18675
rect 1685 18645 1715 18675
rect 1765 18645 1795 18675
rect 1845 18645 1875 18675
rect 1925 18645 1955 18675
rect 2005 18645 2035 18675
rect 2085 18645 2115 18675
rect 2165 18645 2195 18675
rect 2245 18645 2275 18675
rect 2325 18645 2355 18675
rect 2405 18645 2435 18675
rect 2485 18645 2515 18675
rect 2565 18645 2595 18675
rect 2645 18645 2675 18675
rect 2725 18645 2755 18675
rect 2805 18645 2835 18675
rect 2885 18645 2915 18675
rect 2965 18645 2995 18675
rect 3045 18645 3075 18675
rect 3125 18645 3155 18675
rect 3205 18645 3235 18675
rect 3285 18645 3315 18675
rect 3365 18645 3395 18675
rect 3445 18645 3475 18675
rect 3525 18645 3555 18675
rect 3605 18645 3635 18675
rect 3685 18645 3715 18675
rect 3765 18645 3795 18675
rect 3845 18645 3875 18675
rect 3925 18645 3955 18675
rect 4005 18645 4035 18675
rect 4085 18645 4115 18675
rect 4165 18645 4195 18675
rect 4245 18645 4275 18675
rect 4405 18645 4435 18675
rect 6245 18645 6275 18675
rect 6325 18645 6355 18675
rect 6405 18645 6435 18675
rect 6485 18645 6515 18675
rect 6565 18645 6595 18675
rect 6645 18645 6675 18675
rect 6725 18645 6755 18675
rect 6805 18645 6835 18675
rect 6885 18645 6915 18675
rect 6965 18645 6995 18675
rect 7045 18645 7075 18675
rect 7125 18645 7155 18675
rect 7205 18645 7235 18675
rect 7285 18645 7315 18675
rect 7365 18645 7395 18675
rect 7445 18645 7475 18675
rect 7525 18645 7555 18675
rect 7605 18645 7635 18675
rect 7685 18645 7715 18675
rect 7765 18645 7795 18675
rect 7845 18645 7875 18675
rect 7925 18645 7955 18675
rect 8005 18645 8035 18675
rect 8085 18645 8115 18675
rect 8165 18645 8195 18675
rect 8245 18645 8275 18675
rect 8325 18645 8355 18675
rect 8405 18645 8435 18675
rect 8485 18645 8515 18675
rect 8565 18645 8595 18675
rect 8645 18645 8675 18675
rect 8725 18645 8755 18675
rect 8805 18645 8835 18675
rect 8885 18645 8915 18675
rect 8965 18645 8995 18675
rect 9045 18645 9075 18675
rect 9125 18645 9155 18675
rect 9205 18645 9235 18675
rect 9285 18645 9315 18675
rect 9365 18645 9395 18675
rect 9445 18645 9475 18675
rect 11285 18645 11315 18675
rect 11445 18645 11475 18675
rect 11565 18645 11595 18675
rect 11645 18645 11675 18675
rect 11725 18645 11755 18675
rect 11805 18645 11835 18675
rect 11885 18645 11915 18675
rect 11965 18645 11995 18675
rect 12045 18645 12075 18675
rect 12125 18645 12155 18675
rect 12205 18645 12235 18675
rect 12285 18645 12315 18675
rect 12365 18645 12395 18675
rect 12445 18645 12475 18675
rect 12525 18645 12555 18675
rect 12605 18645 12635 18675
rect 12685 18645 12715 18675
rect 12765 18645 12795 18675
rect 12845 18645 12875 18675
rect 12925 18645 12955 18675
rect 13005 18645 13035 18675
rect 13085 18645 13115 18675
rect 13165 18645 13195 18675
rect 13245 18645 13275 18675
rect 13325 18645 13355 18675
rect 13405 18645 13435 18675
rect 13485 18645 13515 18675
rect 13565 18645 13595 18675
rect 13645 18645 13675 18675
rect 13725 18645 13755 18675
rect 13805 18645 13835 18675
rect 13885 18645 13915 18675
rect 13965 18645 13995 18675
rect 14045 18645 14075 18675
rect 14125 18645 14155 18675
rect 14205 18645 14235 18675
rect 14285 18645 14315 18675
rect 14365 18645 14395 18675
rect 14445 18645 14475 18675
rect 14525 18645 14555 18675
rect 14605 18645 14635 18675
rect 14685 18645 14715 18675
rect 16525 18645 16555 18675
rect 16685 18645 16715 18675
rect 16765 18645 16795 18675
rect 16845 18645 16875 18675
rect 16925 18645 16955 18675
rect 17005 18645 17035 18675
rect 17085 18645 17115 18675
rect 17165 18645 17195 18675
rect 17245 18645 17275 18675
rect 17325 18645 17355 18675
rect 17405 18645 17435 18675
rect 17485 18645 17515 18675
rect 17565 18645 17595 18675
rect 17645 18645 17675 18675
rect 17725 18645 17755 18675
rect 17805 18645 17835 18675
rect 17885 18645 17915 18675
rect 17965 18645 17995 18675
rect 18045 18645 18075 18675
rect 18125 18645 18155 18675
rect 18205 18645 18235 18675
rect 18285 18645 18315 18675
rect 18365 18645 18395 18675
rect 18445 18645 18475 18675
rect 18525 18645 18555 18675
rect 18605 18645 18635 18675
rect 18685 18645 18715 18675
rect 18765 18645 18795 18675
rect 18845 18645 18875 18675
rect 18925 18645 18955 18675
rect 19005 18645 19035 18675
rect 19085 18645 19115 18675
rect 19165 18645 19195 18675
rect 19245 18645 19275 18675
rect 19325 18645 19355 18675
rect 19405 18645 19435 18675
rect 19485 18645 19515 18675
rect 19565 18645 19595 18675
rect 19645 18645 19675 18675
rect 19725 18645 19755 18675
rect 19805 18645 19835 18675
rect 19885 18645 19915 18675
rect 19965 18645 19995 18675
rect 20045 18645 20075 18675
rect 20125 18645 20155 18675
rect 20205 18645 20235 18675
rect 20285 18645 20315 18675
rect 20365 18645 20395 18675
rect 20445 18645 20475 18675
rect 20525 18645 20555 18675
rect 20605 18645 20635 18675
rect 20685 18645 20715 18675
rect 20765 18645 20795 18675
rect 20845 18645 20875 18675
rect 20925 18645 20955 18675
rect 4325 18565 4355 18595
rect 11365 18565 11395 18595
rect 16605 18565 16635 18595
rect 5 18485 35 18515
rect 85 18485 115 18515
rect 165 18485 195 18515
rect 245 18485 275 18515
rect 325 18485 355 18515
rect 405 18485 435 18515
rect 485 18485 515 18515
rect 565 18485 595 18515
rect 645 18485 675 18515
rect 725 18485 755 18515
rect 805 18485 835 18515
rect 885 18485 915 18515
rect 965 18485 995 18515
rect 1045 18485 1075 18515
rect 1125 18485 1155 18515
rect 1205 18485 1235 18515
rect 1285 18485 1315 18515
rect 1365 18485 1395 18515
rect 1445 18485 1475 18515
rect 1525 18485 1555 18515
rect 1605 18485 1635 18515
rect 1685 18485 1715 18515
rect 1765 18485 1795 18515
rect 1845 18485 1875 18515
rect 1925 18485 1955 18515
rect 2005 18485 2035 18515
rect 2085 18485 2115 18515
rect 2165 18485 2195 18515
rect 2245 18485 2275 18515
rect 2325 18485 2355 18515
rect 2405 18485 2435 18515
rect 2485 18485 2515 18515
rect 2565 18485 2595 18515
rect 2645 18485 2675 18515
rect 2725 18485 2755 18515
rect 2805 18485 2835 18515
rect 2885 18485 2915 18515
rect 2965 18485 2995 18515
rect 3045 18485 3075 18515
rect 3125 18485 3155 18515
rect 3205 18485 3235 18515
rect 3285 18485 3315 18515
rect 3365 18485 3395 18515
rect 3445 18485 3475 18515
rect 3525 18485 3555 18515
rect 3605 18485 3635 18515
rect 3685 18485 3715 18515
rect 3765 18485 3795 18515
rect 3845 18485 3875 18515
rect 3925 18485 3955 18515
rect 4005 18485 4035 18515
rect 4085 18485 4115 18515
rect 4165 18485 4195 18515
rect 4245 18485 4275 18515
rect 4405 18485 4435 18515
rect 6245 18485 6275 18515
rect 6325 18485 6355 18515
rect 6405 18485 6435 18515
rect 6485 18485 6515 18515
rect 6565 18485 6595 18515
rect 6645 18485 6675 18515
rect 6725 18485 6755 18515
rect 6805 18485 6835 18515
rect 6885 18485 6915 18515
rect 6965 18485 6995 18515
rect 7045 18485 7075 18515
rect 7125 18485 7155 18515
rect 7205 18485 7235 18515
rect 7285 18485 7315 18515
rect 7365 18485 7395 18515
rect 7445 18485 7475 18515
rect 7525 18485 7555 18515
rect 7605 18485 7635 18515
rect 7685 18485 7715 18515
rect 7765 18485 7795 18515
rect 7845 18485 7875 18515
rect 7925 18485 7955 18515
rect 8005 18485 8035 18515
rect 8085 18485 8115 18515
rect 8165 18485 8195 18515
rect 8245 18485 8275 18515
rect 8325 18485 8355 18515
rect 8405 18485 8435 18515
rect 8485 18485 8515 18515
rect 8565 18485 8595 18515
rect 8645 18485 8675 18515
rect 8725 18485 8755 18515
rect 8805 18485 8835 18515
rect 8885 18485 8915 18515
rect 8965 18485 8995 18515
rect 9045 18485 9075 18515
rect 9125 18485 9155 18515
rect 9205 18485 9235 18515
rect 9285 18485 9315 18515
rect 9365 18485 9395 18515
rect 9445 18485 9475 18515
rect 11285 18485 11315 18515
rect 11445 18485 11475 18515
rect 11565 18485 11595 18515
rect 11645 18485 11675 18515
rect 11725 18485 11755 18515
rect 11805 18485 11835 18515
rect 11885 18485 11915 18515
rect 11965 18485 11995 18515
rect 12045 18485 12075 18515
rect 12125 18485 12155 18515
rect 12205 18485 12235 18515
rect 12285 18485 12315 18515
rect 12365 18485 12395 18515
rect 12445 18485 12475 18515
rect 12525 18485 12555 18515
rect 12605 18485 12635 18515
rect 12685 18485 12715 18515
rect 12765 18485 12795 18515
rect 12845 18485 12875 18515
rect 12925 18485 12955 18515
rect 13005 18485 13035 18515
rect 13085 18485 13115 18515
rect 13165 18485 13195 18515
rect 13245 18485 13275 18515
rect 13325 18485 13355 18515
rect 13405 18485 13435 18515
rect 13485 18485 13515 18515
rect 13565 18485 13595 18515
rect 13645 18485 13675 18515
rect 13725 18485 13755 18515
rect 13805 18485 13835 18515
rect 13885 18485 13915 18515
rect 13965 18485 13995 18515
rect 14045 18485 14075 18515
rect 14125 18485 14155 18515
rect 14205 18485 14235 18515
rect 14285 18485 14315 18515
rect 14365 18485 14395 18515
rect 14445 18485 14475 18515
rect 14525 18485 14555 18515
rect 14605 18485 14635 18515
rect 14685 18485 14715 18515
rect 16525 18485 16555 18515
rect 16685 18485 16715 18515
rect 16765 18485 16795 18515
rect 16845 18485 16875 18515
rect 16925 18485 16955 18515
rect 17005 18485 17035 18515
rect 17085 18485 17115 18515
rect 17165 18485 17195 18515
rect 17245 18485 17275 18515
rect 17325 18485 17355 18515
rect 17405 18485 17435 18515
rect 17485 18485 17515 18515
rect 17565 18485 17595 18515
rect 17645 18485 17675 18515
rect 17725 18485 17755 18515
rect 17805 18485 17835 18515
rect 17885 18485 17915 18515
rect 17965 18485 17995 18515
rect 18045 18485 18075 18515
rect 18125 18485 18155 18515
rect 18205 18485 18235 18515
rect 18285 18485 18315 18515
rect 18365 18485 18395 18515
rect 18445 18485 18475 18515
rect 18525 18485 18555 18515
rect 18605 18485 18635 18515
rect 18685 18485 18715 18515
rect 18765 18485 18795 18515
rect 18845 18485 18875 18515
rect 18925 18485 18955 18515
rect 19005 18485 19035 18515
rect 19085 18485 19115 18515
rect 19165 18485 19195 18515
rect 19245 18485 19275 18515
rect 19325 18485 19355 18515
rect 19405 18485 19435 18515
rect 19485 18485 19515 18515
rect 19565 18485 19595 18515
rect 19645 18485 19675 18515
rect 19725 18485 19755 18515
rect 19805 18485 19835 18515
rect 19885 18485 19915 18515
rect 19965 18485 19995 18515
rect 20045 18485 20075 18515
rect 20125 18485 20155 18515
rect 20205 18485 20235 18515
rect 20285 18485 20315 18515
rect 20365 18485 20395 18515
rect 20445 18485 20475 18515
rect 20525 18485 20555 18515
rect 20605 18485 20635 18515
rect 20685 18485 20715 18515
rect 20765 18485 20795 18515
rect 20845 18485 20875 18515
rect 20925 18485 20955 18515
rect 5 18405 35 18435
rect 85 18405 115 18435
rect 165 18405 195 18435
rect 245 18405 275 18435
rect 325 18405 355 18435
rect 405 18405 435 18435
rect 485 18405 515 18435
rect 565 18405 595 18435
rect 645 18405 675 18435
rect 725 18405 755 18435
rect 805 18405 835 18435
rect 885 18405 915 18435
rect 965 18405 995 18435
rect 1045 18405 1075 18435
rect 1125 18405 1155 18435
rect 1205 18405 1235 18435
rect 1285 18405 1315 18435
rect 1365 18405 1395 18435
rect 1445 18405 1475 18435
rect 1525 18405 1555 18435
rect 1605 18405 1635 18435
rect 1685 18405 1715 18435
rect 1765 18405 1795 18435
rect 1845 18405 1875 18435
rect 1925 18405 1955 18435
rect 2005 18405 2035 18435
rect 2085 18405 2115 18435
rect 2165 18405 2195 18435
rect 2245 18405 2275 18435
rect 2325 18405 2355 18435
rect 2405 18405 2435 18435
rect 2485 18405 2515 18435
rect 2565 18405 2595 18435
rect 2645 18405 2675 18435
rect 2725 18405 2755 18435
rect 2805 18405 2835 18435
rect 2885 18405 2915 18435
rect 2965 18405 2995 18435
rect 3045 18405 3075 18435
rect 3125 18405 3155 18435
rect 3205 18405 3235 18435
rect 3285 18405 3315 18435
rect 3365 18405 3395 18435
rect 3445 18405 3475 18435
rect 3525 18405 3555 18435
rect 3605 18405 3635 18435
rect 3685 18405 3715 18435
rect 3765 18405 3795 18435
rect 3845 18405 3875 18435
rect 3925 18405 3955 18435
rect 4005 18405 4035 18435
rect 4085 18405 4115 18435
rect 4165 18405 4195 18435
rect 4485 18405 4515 18435
rect 4645 18405 4675 18435
rect 6245 18405 6275 18435
rect 6325 18405 6355 18435
rect 6405 18405 6435 18435
rect 6485 18405 6515 18435
rect 6565 18405 6595 18435
rect 6645 18405 6675 18435
rect 6725 18405 6755 18435
rect 6805 18405 6835 18435
rect 6885 18405 6915 18435
rect 6965 18405 6995 18435
rect 7045 18405 7075 18435
rect 7125 18405 7155 18435
rect 7205 18405 7235 18435
rect 7285 18405 7315 18435
rect 7365 18405 7395 18435
rect 7445 18405 7475 18435
rect 7525 18405 7555 18435
rect 7605 18405 7635 18435
rect 7685 18405 7715 18435
rect 7765 18405 7795 18435
rect 7845 18405 7875 18435
rect 7925 18405 7955 18435
rect 8005 18405 8035 18435
rect 8085 18405 8115 18435
rect 8165 18405 8195 18435
rect 8245 18405 8275 18435
rect 8325 18405 8355 18435
rect 8405 18405 8435 18435
rect 8485 18405 8515 18435
rect 8565 18405 8595 18435
rect 8645 18405 8675 18435
rect 8725 18405 8755 18435
rect 8805 18405 8835 18435
rect 8885 18405 8915 18435
rect 8965 18405 8995 18435
rect 9045 18405 9075 18435
rect 9125 18405 9155 18435
rect 9205 18405 9235 18435
rect 9285 18405 9315 18435
rect 9365 18405 9395 18435
rect 9445 18405 9475 18435
rect 11045 18405 11075 18435
rect 11205 18405 11235 18435
rect 11565 18405 11595 18435
rect 11645 18405 11675 18435
rect 11725 18405 11755 18435
rect 11805 18405 11835 18435
rect 11885 18405 11915 18435
rect 11965 18405 11995 18435
rect 12045 18405 12075 18435
rect 12125 18405 12155 18435
rect 12205 18405 12235 18435
rect 12285 18405 12315 18435
rect 12365 18405 12395 18435
rect 12445 18405 12475 18435
rect 12525 18405 12555 18435
rect 12605 18405 12635 18435
rect 12685 18405 12715 18435
rect 12765 18405 12795 18435
rect 12845 18405 12875 18435
rect 12925 18405 12955 18435
rect 13005 18405 13035 18435
rect 13085 18405 13115 18435
rect 13165 18405 13195 18435
rect 13245 18405 13275 18435
rect 13325 18405 13355 18435
rect 13405 18405 13435 18435
rect 13485 18405 13515 18435
rect 13565 18405 13595 18435
rect 13645 18405 13675 18435
rect 13725 18405 13755 18435
rect 13805 18405 13835 18435
rect 13885 18405 13915 18435
rect 13965 18405 13995 18435
rect 14045 18405 14075 18435
rect 14125 18405 14155 18435
rect 14205 18405 14235 18435
rect 14285 18405 14315 18435
rect 14365 18405 14395 18435
rect 14445 18405 14475 18435
rect 14525 18405 14555 18435
rect 14605 18405 14635 18435
rect 14685 18405 14715 18435
rect 16285 18405 16315 18435
rect 16445 18405 16475 18435
rect 16765 18405 16795 18435
rect 16845 18405 16875 18435
rect 16925 18405 16955 18435
rect 17005 18405 17035 18435
rect 17085 18405 17115 18435
rect 17165 18405 17195 18435
rect 17245 18405 17275 18435
rect 17325 18405 17355 18435
rect 17405 18405 17435 18435
rect 17485 18405 17515 18435
rect 17565 18405 17595 18435
rect 17645 18405 17675 18435
rect 17725 18405 17755 18435
rect 17805 18405 17835 18435
rect 17885 18405 17915 18435
rect 17965 18405 17995 18435
rect 18045 18405 18075 18435
rect 18125 18405 18155 18435
rect 18205 18405 18235 18435
rect 18285 18405 18315 18435
rect 18365 18405 18395 18435
rect 18445 18405 18475 18435
rect 18525 18405 18555 18435
rect 18605 18405 18635 18435
rect 18685 18405 18715 18435
rect 18765 18405 18795 18435
rect 18845 18405 18875 18435
rect 18925 18405 18955 18435
rect 19005 18405 19035 18435
rect 19085 18405 19115 18435
rect 19165 18405 19195 18435
rect 19245 18405 19275 18435
rect 19325 18405 19355 18435
rect 19405 18405 19435 18435
rect 19485 18405 19515 18435
rect 19565 18405 19595 18435
rect 19645 18405 19675 18435
rect 19725 18405 19755 18435
rect 19805 18405 19835 18435
rect 19885 18405 19915 18435
rect 19965 18405 19995 18435
rect 20045 18405 20075 18435
rect 20125 18405 20155 18435
rect 20205 18405 20235 18435
rect 20285 18405 20315 18435
rect 20365 18405 20395 18435
rect 20445 18405 20475 18435
rect 20525 18405 20555 18435
rect 20605 18405 20635 18435
rect 20685 18405 20715 18435
rect 20765 18405 20795 18435
rect 20845 18405 20875 18435
rect 20925 18405 20955 18435
rect 4565 18325 4595 18355
rect 11125 18325 11155 18355
rect 16365 18325 16395 18355
rect 5 18245 35 18275
rect 85 18245 115 18275
rect 165 18245 195 18275
rect 245 18245 275 18275
rect 325 18245 355 18275
rect 405 18245 435 18275
rect 485 18245 515 18275
rect 565 18245 595 18275
rect 645 18245 675 18275
rect 725 18245 755 18275
rect 805 18245 835 18275
rect 885 18245 915 18275
rect 965 18245 995 18275
rect 1045 18245 1075 18275
rect 1125 18245 1155 18275
rect 1205 18245 1235 18275
rect 1285 18245 1315 18275
rect 1365 18245 1395 18275
rect 1445 18245 1475 18275
rect 1525 18245 1555 18275
rect 1605 18245 1635 18275
rect 1685 18245 1715 18275
rect 1765 18245 1795 18275
rect 1845 18245 1875 18275
rect 1925 18245 1955 18275
rect 2005 18245 2035 18275
rect 2085 18245 2115 18275
rect 2165 18245 2195 18275
rect 2245 18245 2275 18275
rect 2325 18245 2355 18275
rect 2405 18245 2435 18275
rect 2485 18245 2515 18275
rect 2565 18245 2595 18275
rect 2645 18245 2675 18275
rect 2725 18245 2755 18275
rect 2805 18245 2835 18275
rect 2885 18245 2915 18275
rect 2965 18245 2995 18275
rect 3045 18245 3075 18275
rect 3125 18245 3155 18275
rect 3205 18245 3235 18275
rect 3285 18245 3315 18275
rect 3365 18245 3395 18275
rect 3445 18245 3475 18275
rect 3525 18245 3555 18275
rect 3605 18245 3635 18275
rect 3685 18245 3715 18275
rect 3765 18245 3795 18275
rect 3845 18245 3875 18275
rect 3925 18245 3955 18275
rect 4005 18245 4035 18275
rect 4085 18245 4115 18275
rect 4165 18245 4195 18275
rect 4485 18245 4515 18275
rect 4645 18245 4675 18275
rect 6245 18245 6275 18275
rect 6325 18245 6355 18275
rect 6405 18245 6435 18275
rect 6485 18245 6515 18275
rect 6565 18245 6595 18275
rect 6645 18245 6675 18275
rect 6725 18245 6755 18275
rect 6805 18245 6835 18275
rect 6885 18245 6915 18275
rect 6965 18245 6995 18275
rect 7045 18245 7075 18275
rect 7125 18245 7155 18275
rect 7205 18245 7235 18275
rect 7285 18245 7315 18275
rect 7365 18245 7395 18275
rect 7445 18245 7475 18275
rect 7525 18245 7555 18275
rect 7605 18245 7635 18275
rect 7685 18245 7715 18275
rect 7765 18245 7795 18275
rect 7845 18245 7875 18275
rect 7925 18245 7955 18275
rect 8005 18245 8035 18275
rect 8085 18245 8115 18275
rect 8165 18245 8195 18275
rect 8245 18245 8275 18275
rect 8325 18245 8355 18275
rect 8405 18245 8435 18275
rect 8485 18245 8515 18275
rect 8565 18245 8595 18275
rect 8645 18245 8675 18275
rect 8725 18245 8755 18275
rect 8805 18245 8835 18275
rect 8885 18245 8915 18275
rect 8965 18245 8995 18275
rect 9045 18245 9075 18275
rect 9125 18245 9155 18275
rect 9205 18245 9235 18275
rect 9285 18245 9315 18275
rect 9365 18245 9395 18275
rect 9445 18245 9475 18275
rect 11045 18245 11075 18275
rect 11205 18245 11235 18275
rect 11565 18245 11595 18275
rect 11645 18245 11675 18275
rect 11725 18245 11755 18275
rect 11805 18245 11835 18275
rect 11885 18245 11915 18275
rect 11965 18245 11995 18275
rect 12045 18245 12075 18275
rect 12125 18245 12155 18275
rect 12205 18245 12235 18275
rect 12285 18245 12315 18275
rect 12365 18245 12395 18275
rect 12445 18245 12475 18275
rect 12525 18245 12555 18275
rect 12605 18245 12635 18275
rect 12685 18245 12715 18275
rect 12765 18245 12795 18275
rect 12845 18245 12875 18275
rect 12925 18245 12955 18275
rect 13005 18245 13035 18275
rect 13085 18245 13115 18275
rect 13165 18245 13195 18275
rect 13245 18245 13275 18275
rect 13325 18245 13355 18275
rect 13405 18245 13435 18275
rect 13485 18245 13515 18275
rect 13565 18245 13595 18275
rect 13645 18245 13675 18275
rect 13725 18245 13755 18275
rect 13805 18245 13835 18275
rect 13885 18245 13915 18275
rect 13965 18245 13995 18275
rect 14045 18245 14075 18275
rect 14125 18245 14155 18275
rect 14205 18245 14235 18275
rect 14285 18245 14315 18275
rect 14365 18245 14395 18275
rect 14445 18245 14475 18275
rect 14525 18245 14555 18275
rect 14605 18245 14635 18275
rect 14685 18245 14715 18275
rect 16285 18245 16315 18275
rect 16445 18245 16475 18275
rect 16765 18245 16795 18275
rect 16845 18245 16875 18275
rect 16925 18245 16955 18275
rect 17005 18245 17035 18275
rect 17085 18245 17115 18275
rect 17165 18245 17195 18275
rect 17245 18245 17275 18275
rect 17325 18245 17355 18275
rect 17405 18245 17435 18275
rect 17485 18245 17515 18275
rect 17565 18245 17595 18275
rect 17645 18245 17675 18275
rect 17725 18245 17755 18275
rect 17805 18245 17835 18275
rect 17885 18245 17915 18275
rect 17965 18245 17995 18275
rect 18045 18245 18075 18275
rect 18125 18245 18155 18275
rect 18205 18245 18235 18275
rect 18285 18245 18315 18275
rect 18365 18245 18395 18275
rect 18445 18245 18475 18275
rect 18525 18245 18555 18275
rect 18605 18245 18635 18275
rect 18685 18245 18715 18275
rect 18765 18245 18795 18275
rect 18845 18245 18875 18275
rect 18925 18245 18955 18275
rect 19005 18245 19035 18275
rect 19085 18245 19115 18275
rect 19165 18245 19195 18275
rect 19245 18245 19275 18275
rect 19325 18245 19355 18275
rect 19405 18245 19435 18275
rect 19485 18245 19515 18275
rect 19565 18245 19595 18275
rect 19645 18245 19675 18275
rect 19725 18245 19755 18275
rect 19805 18245 19835 18275
rect 19885 18245 19915 18275
rect 19965 18245 19995 18275
rect 20045 18245 20075 18275
rect 20125 18245 20155 18275
rect 20205 18245 20235 18275
rect 20285 18245 20315 18275
rect 20365 18245 20395 18275
rect 20445 18245 20475 18275
rect 20525 18245 20555 18275
rect 20605 18245 20635 18275
rect 20685 18245 20715 18275
rect 20765 18245 20795 18275
rect 20845 18245 20875 18275
rect 20925 18245 20955 18275
rect 5 18165 35 18195
rect 85 18165 115 18195
rect 165 18165 195 18195
rect 245 18165 275 18195
rect 325 18165 355 18195
rect 405 18165 435 18195
rect 485 18165 515 18195
rect 565 18165 595 18195
rect 645 18165 675 18195
rect 725 18165 755 18195
rect 805 18165 835 18195
rect 885 18165 915 18195
rect 965 18165 995 18195
rect 1045 18165 1075 18195
rect 1125 18165 1155 18195
rect 1205 18165 1235 18195
rect 1285 18165 1315 18195
rect 1365 18165 1395 18195
rect 1445 18165 1475 18195
rect 1525 18165 1555 18195
rect 1605 18165 1635 18195
rect 1685 18165 1715 18195
rect 1765 18165 1795 18195
rect 1845 18165 1875 18195
rect 1925 18165 1955 18195
rect 2005 18165 2035 18195
rect 2085 18165 2115 18195
rect 2165 18165 2195 18195
rect 2245 18165 2275 18195
rect 2325 18165 2355 18195
rect 2405 18165 2435 18195
rect 2485 18165 2515 18195
rect 2565 18165 2595 18195
rect 2645 18165 2675 18195
rect 2725 18165 2755 18195
rect 2805 18165 2835 18195
rect 2885 18165 2915 18195
rect 2965 18165 2995 18195
rect 3045 18165 3075 18195
rect 3125 18165 3155 18195
rect 3205 18165 3235 18195
rect 3285 18165 3315 18195
rect 3365 18165 3395 18195
rect 3445 18165 3475 18195
rect 3525 18165 3555 18195
rect 3605 18165 3635 18195
rect 3685 18165 3715 18195
rect 3765 18165 3795 18195
rect 3845 18165 3875 18195
rect 3925 18165 3955 18195
rect 4005 18165 4035 18195
rect 4085 18165 4115 18195
rect 4165 18165 4195 18195
rect 4725 18165 4755 18195
rect 4885 18165 4915 18195
rect 5045 18165 5075 18195
rect 5205 18165 5235 18195
rect 5365 18165 5395 18195
rect 5525 18165 5555 18195
rect 5685 18165 5715 18195
rect 6245 18165 6275 18195
rect 6325 18165 6355 18195
rect 6405 18165 6435 18195
rect 6485 18165 6515 18195
rect 6565 18165 6595 18195
rect 6645 18165 6675 18195
rect 6725 18165 6755 18195
rect 6805 18165 6835 18195
rect 6885 18165 6915 18195
rect 6965 18165 6995 18195
rect 7045 18165 7075 18195
rect 7125 18165 7155 18195
rect 7205 18165 7235 18195
rect 7285 18165 7315 18195
rect 7365 18165 7395 18195
rect 7445 18165 7475 18195
rect 7525 18165 7555 18195
rect 7605 18165 7635 18195
rect 7685 18165 7715 18195
rect 7765 18165 7795 18195
rect 7845 18165 7875 18195
rect 7925 18165 7955 18195
rect 8005 18165 8035 18195
rect 8085 18165 8115 18195
rect 8165 18165 8195 18195
rect 8245 18165 8275 18195
rect 8325 18165 8355 18195
rect 8405 18165 8435 18195
rect 8485 18165 8515 18195
rect 8565 18165 8595 18195
rect 8645 18165 8675 18195
rect 8725 18165 8755 18195
rect 8805 18165 8835 18195
rect 8885 18165 8915 18195
rect 8965 18165 8995 18195
rect 9045 18165 9075 18195
rect 9125 18165 9155 18195
rect 9205 18165 9235 18195
rect 9285 18165 9315 18195
rect 9365 18165 9395 18195
rect 9445 18165 9475 18195
rect 10005 18165 10035 18195
rect 10165 18165 10195 18195
rect 10325 18165 10355 18195
rect 10485 18165 10515 18195
rect 10645 18165 10675 18195
rect 10805 18165 10835 18195
rect 10965 18165 10995 18195
rect 11565 18165 11595 18195
rect 11645 18165 11675 18195
rect 11725 18165 11755 18195
rect 11805 18165 11835 18195
rect 11885 18165 11915 18195
rect 11965 18165 11995 18195
rect 12045 18165 12075 18195
rect 12125 18165 12155 18195
rect 12205 18165 12235 18195
rect 12285 18165 12315 18195
rect 12365 18165 12395 18195
rect 12445 18165 12475 18195
rect 12525 18165 12555 18195
rect 12605 18165 12635 18195
rect 12685 18165 12715 18195
rect 12765 18165 12795 18195
rect 12845 18165 12875 18195
rect 12925 18165 12955 18195
rect 13005 18165 13035 18195
rect 13085 18165 13115 18195
rect 13165 18165 13195 18195
rect 13245 18165 13275 18195
rect 13325 18165 13355 18195
rect 13405 18165 13435 18195
rect 13485 18165 13515 18195
rect 13565 18165 13595 18195
rect 13645 18165 13675 18195
rect 13725 18165 13755 18195
rect 13805 18165 13835 18195
rect 13885 18165 13915 18195
rect 13965 18165 13995 18195
rect 14045 18165 14075 18195
rect 14125 18165 14155 18195
rect 14205 18165 14235 18195
rect 14285 18165 14315 18195
rect 14365 18165 14395 18195
rect 14445 18165 14475 18195
rect 14525 18165 14555 18195
rect 14605 18165 14635 18195
rect 14685 18165 14715 18195
rect 15245 18165 15275 18195
rect 15405 18165 15435 18195
rect 15565 18165 15595 18195
rect 15725 18165 15755 18195
rect 15885 18165 15915 18195
rect 16045 18165 16075 18195
rect 16205 18165 16235 18195
rect 16765 18165 16795 18195
rect 16845 18165 16875 18195
rect 16925 18165 16955 18195
rect 17005 18165 17035 18195
rect 17085 18165 17115 18195
rect 17165 18165 17195 18195
rect 17245 18165 17275 18195
rect 17325 18165 17355 18195
rect 17405 18165 17435 18195
rect 17485 18165 17515 18195
rect 17565 18165 17595 18195
rect 17645 18165 17675 18195
rect 17725 18165 17755 18195
rect 17805 18165 17835 18195
rect 17885 18165 17915 18195
rect 17965 18165 17995 18195
rect 18045 18165 18075 18195
rect 18125 18165 18155 18195
rect 18205 18165 18235 18195
rect 18285 18165 18315 18195
rect 18365 18165 18395 18195
rect 18445 18165 18475 18195
rect 18525 18165 18555 18195
rect 18605 18165 18635 18195
rect 18685 18165 18715 18195
rect 18765 18165 18795 18195
rect 18845 18165 18875 18195
rect 18925 18165 18955 18195
rect 19005 18165 19035 18195
rect 19085 18165 19115 18195
rect 19165 18165 19195 18195
rect 19245 18165 19275 18195
rect 19325 18165 19355 18195
rect 19405 18165 19435 18195
rect 19485 18165 19515 18195
rect 19565 18165 19595 18195
rect 19645 18165 19675 18195
rect 19725 18165 19755 18195
rect 19805 18165 19835 18195
rect 19885 18165 19915 18195
rect 19965 18165 19995 18195
rect 20045 18165 20075 18195
rect 20125 18165 20155 18195
rect 20205 18165 20235 18195
rect 20285 18165 20315 18195
rect 20365 18165 20395 18195
rect 20445 18165 20475 18195
rect 20525 18165 20555 18195
rect 20605 18165 20635 18195
rect 20685 18165 20715 18195
rect 20765 18165 20795 18195
rect 20845 18165 20875 18195
rect 20925 18165 20955 18195
rect 4805 18085 4835 18115
rect 10885 18085 10915 18115
rect 16125 18085 16155 18115
rect 5 18005 35 18035
rect 85 18005 115 18035
rect 165 18005 195 18035
rect 245 18005 275 18035
rect 325 18005 355 18035
rect 405 18005 435 18035
rect 485 18005 515 18035
rect 565 18005 595 18035
rect 645 18005 675 18035
rect 725 18005 755 18035
rect 805 18005 835 18035
rect 885 18005 915 18035
rect 965 18005 995 18035
rect 1045 18005 1075 18035
rect 1125 18005 1155 18035
rect 1205 18005 1235 18035
rect 1285 18005 1315 18035
rect 1365 18005 1395 18035
rect 1445 18005 1475 18035
rect 1525 18005 1555 18035
rect 1605 18005 1635 18035
rect 1685 18005 1715 18035
rect 1765 18005 1795 18035
rect 1845 18005 1875 18035
rect 1925 18005 1955 18035
rect 2005 18005 2035 18035
rect 2085 18005 2115 18035
rect 2165 18005 2195 18035
rect 2245 18005 2275 18035
rect 2325 18005 2355 18035
rect 2405 18005 2435 18035
rect 2485 18005 2515 18035
rect 2565 18005 2595 18035
rect 2645 18005 2675 18035
rect 2725 18005 2755 18035
rect 2805 18005 2835 18035
rect 2885 18005 2915 18035
rect 2965 18005 2995 18035
rect 3045 18005 3075 18035
rect 3125 18005 3155 18035
rect 3205 18005 3235 18035
rect 3285 18005 3315 18035
rect 3365 18005 3395 18035
rect 3445 18005 3475 18035
rect 3525 18005 3555 18035
rect 3605 18005 3635 18035
rect 3685 18005 3715 18035
rect 3765 18005 3795 18035
rect 3845 18005 3875 18035
rect 3925 18005 3955 18035
rect 4005 18005 4035 18035
rect 4085 18005 4115 18035
rect 4165 18005 4195 18035
rect 4725 18005 4755 18035
rect 4885 18005 4915 18035
rect 5045 18005 5075 18035
rect 5205 18005 5235 18035
rect 5365 18005 5395 18035
rect 5525 18005 5555 18035
rect 5685 18005 5715 18035
rect 6245 18005 6275 18035
rect 6325 18005 6355 18035
rect 6405 18005 6435 18035
rect 6485 18005 6515 18035
rect 6565 18005 6595 18035
rect 6645 18005 6675 18035
rect 6725 18005 6755 18035
rect 6805 18005 6835 18035
rect 6885 18005 6915 18035
rect 6965 18005 6995 18035
rect 7045 18005 7075 18035
rect 7125 18005 7155 18035
rect 7205 18005 7235 18035
rect 7285 18005 7315 18035
rect 7365 18005 7395 18035
rect 7445 18005 7475 18035
rect 7525 18005 7555 18035
rect 7605 18005 7635 18035
rect 7685 18005 7715 18035
rect 7765 18005 7795 18035
rect 7845 18005 7875 18035
rect 7925 18005 7955 18035
rect 8005 18005 8035 18035
rect 8085 18005 8115 18035
rect 8165 18005 8195 18035
rect 8245 18005 8275 18035
rect 8325 18005 8355 18035
rect 8405 18005 8435 18035
rect 8485 18005 8515 18035
rect 8565 18005 8595 18035
rect 8645 18005 8675 18035
rect 8725 18005 8755 18035
rect 8805 18005 8835 18035
rect 8885 18005 8915 18035
rect 8965 18005 8995 18035
rect 9045 18005 9075 18035
rect 9125 18005 9155 18035
rect 9205 18005 9235 18035
rect 9285 18005 9315 18035
rect 9365 18005 9395 18035
rect 9445 18005 9475 18035
rect 10005 18005 10035 18035
rect 10165 18005 10195 18035
rect 10325 18005 10355 18035
rect 10485 18005 10515 18035
rect 10645 18005 10675 18035
rect 10805 18005 10835 18035
rect 10965 18005 10995 18035
rect 11565 18005 11595 18035
rect 11645 18005 11675 18035
rect 11725 18005 11755 18035
rect 11805 18005 11835 18035
rect 11885 18005 11915 18035
rect 11965 18005 11995 18035
rect 12045 18005 12075 18035
rect 12125 18005 12155 18035
rect 12205 18005 12235 18035
rect 12285 18005 12315 18035
rect 12365 18005 12395 18035
rect 12445 18005 12475 18035
rect 12525 18005 12555 18035
rect 12605 18005 12635 18035
rect 12685 18005 12715 18035
rect 12765 18005 12795 18035
rect 12845 18005 12875 18035
rect 12925 18005 12955 18035
rect 13005 18005 13035 18035
rect 13085 18005 13115 18035
rect 13165 18005 13195 18035
rect 13245 18005 13275 18035
rect 13325 18005 13355 18035
rect 13405 18005 13435 18035
rect 13485 18005 13515 18035
rect 13565 18005 13595 18035
rect 13645 18005 13675 18035
rect 13725 18005 13755 18035
rect 13805 18005 13835 18035
rect 13885 18005 13915 18035
rect 13965 18005 13995 18035
rect 14045 18005 14075 18035
rect 14125 18005 14155 18035
rect 14205 18005 14235 18035
rect 14285 18005 14315 18035
rect 14365 18005 14395 18035
rect 14445 18005 14475 18035
rect 14525 18005 14555 18035
rect 14605 18005 14635 18035
rect 14685 18005 14715 18035
rect 15245 18005 15275 18035
rect 15405 18005 15435 18035
rect 15565 18005 15595 18035
rect 15725 18005 15755 18035
rect 15885 18005 15915 18035
rect 16045 18005 16075 18035
rect 16205 18005 16235 18035
rect 16765 18005 16795 18035
rect 16845 18005 16875 18035
rect 16925 18005 16955 18035
rect 17005 18005 17035 18035
rect 17085 18005 17115 18035
rect 17165 18005 17195 18035
rect 17245 18005 17275 18035
rect 17325 18005 17355 18035
rect 17405 18005 17435 18035
rect 17485 18005 17515 18035
rect 17565 18005 17595 18035
rect 17645 18005 17675 18035
rect 17725 18005 17755 18035
rect 17805 18005 17835 18035
rect 17885 18005 17915 18035
rect 17965 18005 17995 18035
rect 18045 18005 18075 18035
rect 18125 18005 18155 18035
rect 18205 18005 18235 18035
rect 18285 18005 18315 18035
rect 18365 18005 18395 18035
rect 18445 18005 18475 18035
rect 18525 18005 18555 18035
rect 18605 18005 18635 18035
rect 18685 18005 18715 18035
rect 18765 18005 18795 18035
rect 18845 18005 18875 18035
rect 18925 18005 18955 18035
rect 19005 18005 19035 18035
rect 19085 18005 19115 18035
rect 19165 18005 19195 18035
rect 19245 18005 19275 18035
rect 19325 18005 19355 18035
rect 19405 18005 19435 18035
rect 19485 18005 19515 18035
rect 19565 18005 19595 18035
rect 19645 18005 19675 18035
rect 19725 18005 19755 18035
rect 19805 18005 19835 18035
rect 19885 18005 19915 18035
rect 19965 18005 19995 18035
rect 20045 18005 20075 18035
rect 20125 18005 20155 18035
rect 20205 18005 20235 18035
rect 20285 18005 20315 18035
rect 20365 18005 20395 18035
rect 20445 18005 20475 18035
rect 20525 18005 20555 18035
rect 20605 18005 20635 18035
rect 20685 18005 20715 18035
rect 20765 18005 20795 18035
rect 20845 18005 20875 18035
rect 20925 18005 20955 18035
rect 4965 17925 4995 17955
rect 10725 17925 10755 17955
rect 15965 17925 15995 17955
rect 5 17845 35 17875
rect 85 17845 115 17875
rect 165 17845 195 17875
rect 245 17845 275 17875
rect 325 17845 355 17875
rect 405 17845 435 17875
rect 485 17845 515 17875
rect 565 17845 595 17875
rect 645 17845 675 17875
rect 725 17845 755 17875
rect 805 17845 835 17875
rect 885 17845 915 17875
rect 965 17845 995 17875
rect 1045 17845 1075 17875
rect 1125 17845 1155 17875
rect 1205 17845 1235 17875
rect 1285 17845 1315 17875
rect 1365 17845 1395 17875
rect 1445 17845 1475 17875
rect 1525 17845 1555 17875
rect 1605 17845 1635 17875
rect 1685 17845 1715 17875
rect 1765 17845 1795 17875
rect 1845 17845 1875 17875
rect 1925 17845 1955 17875
rect 2005 17845 2035 17875
rect 2085 17845 2115 17875
rect 2165 17845 2195 17875
rect 2245 17845 2275 17875
rect 2325 17845 2355 17875
rect 2405 17845 2435 17875
rect 2485 17845 2515 17875
rect 2565 17845 2595 17875
rect 2645 17845 2675 17875
rect 2725 17845 2755 17875
rect 2805 17845 2835 17875
rect 2885 17845 2915 17875
rect 2965 17845 2995 17875
rect 3045 17845 3075 17875
rect 3125 17845 3155 17875
rect 3205 17845 3235 17875
rect 3285 17845 3315 17875
rect 3365 17845 3395 17875
rect 3445 17845 3475 17875
rect 3525 17845 3555 17875
rect 3605 17845 3635 17875
rect 3685 17845 3715 17875
rect 3765 17845 3795 17875
rect 3845 17845 3875 17875
rect 3925 17845 3955 17875
rect 4005 17845 4035 17875
rect 4085 17845 4115 17875
rect 4165 17845 4195 17875
rect 4725 17845 4755 17875
rect 4885 17845 4915 17875
rect 5045 17845 5075 17875
rect 5205 17845 5235 17875
rect 5365 17845 5395 17875
rect 5525 17845 5555 17875
rect 5685 17845 5715 17875
rect 6245 17845 6275 17875
rect 6325 17845 6355 17875
rect 6405 17845 6435 17875
rect 6485 17845 6515 17875
rect 6565 17845 6595 17875
rect 6645 17845 6675 17875
rect 6725 17845 6755 17875
rect 6805 17845 6835 17875
rect 6885 17845 6915 17875
rect 6965 17845 6995 17875
rect 7045 17845 7075 17875
rect 7125 17845 7155 17875
rect 7205 17845 7235 17875
rect 7285 17845 7315 17875
rect 7365 17845 7395 17875
rect 7445 17845 7475 17875
rect 7525 17845 7555 17875
rect 7605 17845 7635 17875
rect 7685 17845 7715 17875
rect 7765 17845 7795 17875
rect 7845 17845 7875 17875
rect 7925 17845 7955 17875
rect 8005 17845 8035 17875
rect 8085 17845 8115 17875
rect 8165 17845 8195 17875
rect 8245 17845 8275 17875
rect 8325 17845 8355 17875
rect 8405 17845 8435 17875
rect 8485 17845 8515 17875
rect 8565 17845 8595 17875
rect 8645 17845 8675 17875
rect 8725 17845 8755 17875
rect 8805 17845 8835 17875
rect 8885 17845 8915 17875
rect 8965 17845 8995 17875
rect 9045 17845 9075 17875
rect 9125 17845 9155 17875
rect 9205 17845 9235 17875
rect 9285 17845 9315 17875
rect 9365 17845 9395 17875
rect 9445 17845 9475 17875
rect 10005 17845 10035 17875
rect 10165 17845 10195 17875
rect 10325 17845 10355 17875
rect 10485 17845 10515 17875
rect 10645 17845 10675 17875
rect 10805 17845 10835 17875
rect 10965 17845 10995 17875
rect 11565 17845 11595 17875
rect 11645 17845 11675 17875
rect 11725 17845 11755 17875
rect 11805 17845 11835 17875
rect 11885 17845 11915 17875
rect 11965 17845 11995 17875
rect 12045 17845 12075 17875
rect 12125 17845 12155 17875
rect 12205 17845 12235 17875
rect 12285 17845 12315 17875
rect 12365 17845 12395 17875
rect 12445 17845 12475 17875
rect 12525 17845 12555 17875
rect 12605 17845 12635 17875
rect 12685 17845 12715 17875
rect 12765 17845 12795 17875
rect 12845 17845 12875 17875
rect 12925 17845 12955 17875
rect 13005 17845 13035 17875
rect 13085 17845 13115 17875
rect 13165 17845 13195 17875
rect 13245 17845 13275 17875
rect 13325 17845 13355 17875
rect 13405 17845 13435 17875
rect 13485 17845 13515 17875
rect 13565 17845 13595 17875
rect 13645 17845 13675 17875
rect 13725 17845 13755 17875
rect 13805 17845 13835 17875
rect 13885 17845 13915 17875
rect 13965 17845 13995 17875
rect 14045 17845 14075 17875
rect 14125 17845 14155 17875
rect 14205 17845 14235 17875
rect 14285 17845 14315 17875
rect 14365 17845 14395 17875
rect 14445 17845 14475 17875
rect 14525 17845 14555 17875
rect 14605 17845 14635 17875
rect 14685 17845 14715 17875
rect 15245 17845 15275 17875
rect 15405 17845 15435 17875
rect 15565 17845 15595 17875
rect 15725 17845 15755 17875
rect 15885 17845 15915 17875
rect 16045 17845 16075 17875
rect 16205 17845 16235 17875
rect 16765 17845 16795 17875
rect 16845 17845 16875 17875
rect 16925 17845 16955 17875
rect 17005 17845 17035 17875
rect 17085 17845 17115 17875
rect 17165 17845 17195 17875
rect 17245 17845 17275 17875
rect 17325 17845 17355 17875
rect 17405 17845 17435 17875
rect 17485 17845 17515 17875
rect 17565 17845 17595 17875
rect 17645 17845 17675 17875
rect 17725 17845 17755 17875
rect 17805 17845 17835 17875
rect 17885 17845 17915 17875
rect 17965 17845 17995 17875
rect 18045 17845 18075 17875
rect 18125 17845 18155 17875
rect 18205 17845 18235 17875
rect 18285 17845 18315 17875
rect 18365 17845 18395 17875
rect 18445 17845 18475 17875
rect 18525 17845 18555 17875
rect 18605 17845 18635 17875
rect 18685 17845 18715 17875
rect 18765 17845 18795 17875
rect 18845 17845 18875 17875
rect 18925 17845 18955 17875
rect 19005 17845 19035 17875
rect 19085 17845 19115 17875
rect 19165 17845 19195 17875
rect 19245 17845 19275 17875
rect 19325 17845 19355 17875
rect 19405 17845 19435 17875
rect 19485 17845 19515 17875
rect 19565 17845 19595 17875
rect 19645 17845 19675 17875
rect 19725 17845 19755 17875
rect 19805 17845 19835 17875
rect 19885 17845 19915 17875
rect 19965 17845 19995 17875
rect 20045 17845 20075 17875
rect 20125 17845 20155 17875
rect 20205 17845 20235 17875
rect 20285 17845 20315 17875
rect 20365 17845 20395 17875
rect 20445 17845 20475 17875
rect 20525 17845 20555 17875
rect 20605 17845 20635 17875
rect 20685 17845 20715 17875
rect 20765 17845 20795 17875
rect 20845 17845 20875 17875
rect 20925 17845 20955 17875
rect 5125 17765 5155 17795
rect 10565 17765 10595 17795
rect 15805 17765 15835 17795
rect 5 17685 35 17715
rect 85 17685 115 17715
rect 165 17685 195 17715
rect 245 17685 275 17715
rect 325 17685 355 17715
rect 405 17685 435 17715
rect 485 17685 515 17715
rect 565 17685 595 17715
rect 645 17685 675 17715
rect 725 17685 755 17715
rect 805 17685 835 17715
rect 885 17685 915 17715
rect 965 17685 995 17715
rect 1045 17685 1075 17715
rect 1125 17685 1155 17715
rect 1205 17685 1235 17715
rect 1285 17685 1315 17715
rect 1365 17685 1395 17715
rect 1445 17685 1475 17715
rect 1525 17685 1555 17715
rect 1605 17685 1635 17715
rect 1685 17685 1715 17715
rect 1765 17685 1795 17715
rect 1845 17685 1875 17715
rect 1925 17685 1955 17715
rect 2005 17685 2035 17715
rect 2085 17685 2115 17715
rect 2165 17685 2195 17715
rect 2245 17685 2275 17715
rect 2325 17685 2355 17715
rect 2405 17685 2435 17715
rect 2485 17685 2515 17715
rect 2565 17685 2595 17715
rect 2645 17685 2675 17715
rect 2725 17685 2755 17715
rect 2805 17685 2835 17715
rect 2885 17685 2915 17715
rect 2965 17685 2995 17715
rect 3045 17685 3075 17715
rect 3125 17685 3155 17715
rect 3205 17685 3235 17715
rect 3285 17685 3315 17715
rect 3365 17685 3395 17715
rect 3445 17685 3475 17715
rect 3525 17685 3555 17715
rect 3605 17685 3635 17715
rect 3685 17685 3715 17715
rect 3765 17685 3795 17715
rect 3845 17685 3875 17715
rect 3925 17685 3955 17715
rect 4005 17685 4035 17715
rect 4085 17685 4115 17715
rect 4165 17685 4195 17715
rect 4725 17685 4755 17715
rect 4885 17685 4915 17715
rect 5045 17685 5075 17715
rect 5205 17685 5235 17715
rect 5365 17685 5395 17715
rect 5525 17685 5555 17715
rect 5685 17685 5715 17715
rect 6245 17685 6275 17715
rect 6325 17685 6355 17715
rect 6405 17685 6435 17715
rect 6485 17685 6515 17715
rect 6565 17685 6595 17715
rect 6645 17685 6675 17715
rect 6725 17685 6755 17715
rect 6805 17685 6835 17715
rect 6885 17685 6915 17715
rect 6965 17685 6995 17715
rect 7045 17685 7075 17715
rect 7125 17685 7155 17715
rect 7205 17685 7235 17715
rect 7285 17685 7315 17715
rect 7365 17685 7395 17715
rect 7445 17685 7475 17715
rect 7525 17685 7555 17715
rect 7605 17685 7635 17715
rect 7685 17685 7715 17715
rect 7765 17685 7795 17715
rect 7845 17685 7875 17715
rect 7925 17685 7955 17715
rect 8005 17685 8035 17715
rect 8085 17685 8115 17715
rect 8165 17685 8195 17715
rect 8245 17685 8275 17715
rect 8325 17685 8355 17715
rect 8405 17685 8435 17715
rect 8485 17685 8515 17715
rect 8565 17685 8595 17715
rect 8645 17685 8675 17715
rect 8725 17685 8755 17715
rect 8805 17685 8835 17715
rect 8885 17685 8915 17715
rect 8965 17685 8995 17715
rect 9045 17685 9075 17715
rect 9125 17685 9155 17715
rect 9205 17685 9235 17715
rect 9285 17685 9315 17715
rect 9365 17685 9395 17715
rect 9445 17685 9475 17715
rect 10005 17685 10035 17715
rect 10165 17685 10195 17715
rect 10325 17685 10355 17715
rect 10485 17685 10515 17715
rect 10645 17685 10675 17715
rect 10805 17685 10835 17715
rect 10965 17685 10995 17715
rect 11565 17685 11595 17715
rect 11645 17685 11675 17715
rect 11725 17685 11755 17715
rect 11805 17685 11835 17715
rect 11885 17685 11915 17715
rect 11965 17685 11995 17715
rect 12045 17685 12075 17715
rect 12125 17685 12155 17715
rect 12205 17685 12235 17715
rect 12285 17685 12315 17715
rect 12365 17685 12395 17715
rect 12445 17685 12475 17715
rect 12525 17685 12555 17715
rect 12605 17685 12635 17715
rect 12685 17685 12715 17715
rect 12765 17685 12795 17715
rect 12845 17685 12875 17715
rect 12925 17685 12955 17715
rect 13005 17685 13035 17715
rect 13085 17685 13115 17715
rect 13165 17685 13195 17715
rect 13245 17685 13275 17715
rect 13325 17685 13355 17715
rect 13405 17685 13435 17715
rect 13485 17685 13515 17715
rect 13565 17685 13595 17715
rect 13645 17685 13675 17715
rect 13725 17685 13755 17715
rect 13805 17685 13835 17715
rect 13885 17685 13915 17715
rect 13965 17685 13995 17715
rect 14045 17685 14075 17715
rect 14125 17685 14155 17715
rect 14205 17685 14235 17715
rect 14285 17685 14315 17715
rect 14365 17685 14395 17715
rect 14445 17685 14475 17715
rect 14525 17685 14555 17715
rect 14605 17685 14635 17715
rect 14685 17685 14715 17715
rect 15245 17685 15275 17715
rect 15405 17685 15435 17715
rect 15565 17685 15595 17715
rect 15725 17685 15755 17715
rect 15885 17685 15915 17715
rect 16045 17685 16075 17715
rect 16205 17685 16235 17715
rect 16765 17685 16795 17715
rect 16845 17685 16875 17715
rect 16925 17685 16955 17715
rect 17005 17685 17035 17715
rect 17085 17685 17115 17715
rect 17165 17685 17195 17715
rect 17245 17685 17275 17715
rect 17325 17685 17355 17715
rect 17405 17685 17435 17715
rect 17485 17685 17515 17715
rect 17565 17685 17595 17715
rect 17645 17685 17675 17715
rect 17725 17685 17755 17715
rect 17805 17685 17835 17715
rect 17885 17685 17915 17715
rect 17965 17685 17995 17715
rect 18045 17685 18075 17715
rect 18125 17685 18155 17715
rect 18205 17685 18235 17715
rect 18285 17685 18315 17715
rect 18365 17685 18395 17715
rect 18445 17685 18475 17715
rect 18525 17685 18555 17715
rect 18605 17685 18635 17715
rect 18685 17685 18715 17715
rect 18765 17685 18795 17715
rect 18845 17685 18875 17715
rect 18925 17685 18955 17715
rect 19005 17685 19035 17715
rect 19085 17685 19115 17715
rect 19165 17685 19195 17715
rect 19245 17685 19275 17715
rect 19325 17685 19355 17715
rect 19405 17685 19435 17715
rect 19485 17685 19515 17715
rect 19565 17685 19595 17715
rect 19645 17685 19675 17715
rect 19725 17685 19755 17715
rect 19805 17685 19835 17715
rect 19885 17685 19915 17715
rect 19965 17685 19995 17715
rect 20045 17685 20075 17715
rect 20125 17685 20155 17715
rect 20205 17685 20235 17715
rect 20285 17685 20315 17715
rect 20365 17685 20395 17715
rect 20445 17685 20475 17715
rect 20525 17685 20555 17715
rect 20605 17685 20635 17715
rect 20685 17685 20715 17715
rect 20765 17685 20795 17715
rect 20845 17685 20875 17715
rect 20925 17685 20955 17715
rect 5285 17605 5315 17635
rect 10405 17605 10435 17635
rect 15645 17605 15675 17635
rect 5 17525 35 17555
rect 85 17525 115 17555
rect 165 17525 195 17555
rect 245 17525 275 17555
rect 325 17525 355 17555
rect 405 17525 435 17555
rect 485 17525 515 17555
rect 565 17525 595 17555
rect 645 17525 675 17555
rect 725 17525 755 17555
rect 805 17525 835 17555
rect 885 17525 915 17555
rect 965 17525 995 17555
rect 1045 17525 1075 17555
rect 1125 17525 1155 17555
rect 1205 17525 1235 17555
rect 1285 17525 1315 17555
rect 1365 17525 1395 17555
rect 1445 17525 1475 17555
rect 1525 17525 1555 17555
rect 1605 17525 1635 17555
rect 1685 17525 1715 17555
rect 1765 17525 1795 17555
rect 1845 17525 1875 17555
rect 1925 17525 1955 17555
rect 2005 17525 2035 17555
rect 2085 17525 2115 17555
rect 2165 17525 2195 17555
rect 2245 17525 2275 17555
rect 2325 17525 2355 17555
rect 2405 17525 2435 17555
rect 2485 17525 2515 17555
rect 2565 17525 2595 17555
rect 2645 17525 2675 17555
rect 2725 17525 2755 17555
rect 2805 17525 2835 17555
rect 2885 17525 2915 17555
rect 2965 17525 2995 17555
rect 3045 17525 3075 17555
rect 3125 17525 3155 17555
rect 3205 17525 3235 17555
rect 3285 17525 3315 17555
rect 3365 17525 3395 17555
rect 3445 17525 3475 17555
rect 3525 17525 3555 17555
rect 3605 17525 3635 17555
rect 3685 17525 3715 17555
rect 3765 17525 3795 17555
rect 3845 17525 3875 17555
rect 3925 17525 3955 17555
rect 4005 17525 4035 17555
rect 4085 17525 4115 17555
rect 4165 17525 4195 17555
rect 4725 17525 4755 17555
rect 4885 17525 4915 17555
rect 5045 17525 5075 17555
rect 5205 17525 5235 17555
rect 5365 17525 5395 17555
rect 5525 17525 5555 17555
rect 5685 17525 5715 17555
rect 6245 17525 6275 17555
rect 6325 17525 6355 17555
rect 6405 17525 6435 17555
rect 6485 17525 6515 17555
rect 6565 17525 6595 17555
rect 6645 17525 6675 17555
rect 6725 17525 6755 17555
rect 6805 17525 6835 17555
rect 6885 17525 6915 17555
rect 6965 17525 6995 17555
rect 7045 17525 7075 17555
rect 7125 17525 7155 17555
rect 7205 17525 7235 17555
rect 7285 17525 7315 17555
rect 7365 17525 7395 17555
rect 7445 17525 7475 17555
rect 7525 17525 7555 17555
rect 7605 17525 7635 17555
rect 7685 17525 7715 17555
rect 7765 17525 7795 17555
rect 7845 17525 7875 17555
rect 7925 17525 7955 17555
rect 8005 17525 8035 17555
rect 8085 17525 8115 17555
rect 8165 17525 8195 17555
rect 8245 17525 8275 17555
rect 8325 17525 8355 17555
rect 8405 17525 8435 17555
rect 8485 17525 8515 17555
rect 8565 17525 8595 17555
rect 8645 17525 8675 17555
rect 8725 17525 8755 17555
rect 8805 17525 8835 17555
rect 8885 17525 8915 17555
rect 8965 17525 8995 17555
rect 9045 17525 9075 17555
rect 9125 17525 9155 17555
rect 9205 17525 9235 17555
rect 9285 17525 9315 17555
rect 9365 17525 9395 17555
rect 9445 17525 9475 17555
rect 10005 17525 10035 17555
rect 10165 17525 10195 17555
rect 10325 17525 10355 17555
rect 10485 17525 10515 17555
rect 10645 17525 10675 17555
rect 10805 17525 10835 17555
rect 10965 17525 10995 17555
rect 11565 17525 11595 17555
rect 11645 17525 11675 17555
rect 11725 17525 11755 17555
rect 11805 17525 11835 17555
rect 11885 17525 11915 17555
rect 11965 17525 11995 17555
rect 12045 17525 12075 17555
rect 12125 17525 12155 17555
rect 12205 17525 12235 17555
rect 12285 17525 12315 17555
rect 12365 17525 12395 17555
rect 12445 17525 12475 17555
rect 12525 17525 12555 17555
rect 12605 17525 12635 17555
rect 12685 17525 12715 17555
rect 12765 17525 12795 17555
rect 12845 17525 12875 17555
rect 12925 17525 12955 17555
rect 13005 17525 13035 17555
rect 13085 17525 13115 17555
rect 13165 17525 13195 17555
rect 13245 17525 13275 17555
rect 13325 17525 13355 17555
rect 13405 17525 13435 17555
rect 13485 17525 13515 17555
rect 13565 17525 13595 17555
rect 13645 17525 13675 17555
rect 13725 17525 13755 17555
rect 13805 17525 13835 17555
rect 13885 17525 13915 17555
rect 13965 17525 13995 17555
rect 14045 17525 14075 17555
rect 14125 17525 14155 17555
rect 14205 17525 14235 17555
rect 14285 17525 14315 17555
rect 14365 17525 14395 17555
rect 14445 17525 14475 17555
rect 14525 17525 14555 17555
rect 14605 17525 14635 17555
rect 14685 17525 14715 17555
rect 15245 17525 15275 17555
rect 15405 17525 15435 17555
rect 15565 17525 15595 17555
rect 15725 17525 15755 17555
rect 15885 17525 15915 17555
rect 16045 17525 16075 17555
rect 16205 17525 16235 17555
rect 16765 17525 16795 17555
rect 16845 17525 16875 17555
rect 16925 17525 16955 17555
rect 17005 17525 17035 17555
rect 17085 17525 17115 17555
rect 17165 17525 17195 17555
rect 17245 17525 17275 17555
rect 17325 17525 17355 17555
rect 17405 17525 17435 17555
rect 17485 17525 17515 17555
rect 17565 17525 17595 17555
rect 17645 17525 17675 17555
rect 17725 17525 17755 17555
rect 17805 17525 17835 17555
rect 17885 17525 17915 17555
rect 17965 17525 17995 17555
rect 18045 17525 18075 17555
rect 18125 17525 18155 17555
rect 18205 17525 18235 17555
rect 18285 17525 18315 17555
rect 18365 17525 18395 17555
rect 18445 17525 18475 17555
rect 18525 17525 18555 17555
rect 18605 17525 18635 17555
rect 18685 17525 18715 17555
rect 18765 17525 18795 17555
rect 18845 17525 18875 17555
rect 18925 17525 18955 17555
rect 19005 17525 19035 17555
rect 19085 17525 19115 17555
rect 19165 17525 19195 17555
rect 19245 17525 19275 17555
rect 19325 17525 19355 17555
rect 19405 17525 19435 17555
rect 19485 17525 19515 17555
rect 19565 17525 19595 17555
rect 19645 17525 19675 17555
rect 19725 17525 19755 17555
rect 19805 17525 19835 17555
rect 19885 17525 19915 17555
rect 19965 17525 19995 17555
rect 20045 17525 20075 17555
rect 20125 17525 20155 17555
rect 20205 17525 20235 17555
rect 20285 17525 20315 17555
rect 20365 17525 20395 17555
rect 20445 17525 20475 17555
rect 20525 17525 20555 17555
rect 20605 17525 20635 17555
rect 20685 17525 20715 17555
rect 20765 17525 20795 17555
rect 20845 17525 20875 17555
rect 20925 17525 20955 17555
rect 5445 17445 5475 17475
rect 10245 17445 10275 17475
rect 15485 17445 15515 17475
rect 5 17365 35 17395
rect 85 17365 115 17395
rect 165 17365 195 17395
rect 245 17365 275 17395
rect 325 17365 355 17395
rect 405 17365 435 17395
rect 485 17365 515 17395
rect 565 17365 595 17395
rect 645 17365 675 17395
rect 725 17365 755 17395
rect 805 17365 835 17395
rect 885 17365 915 17395
rect 965 17365 995 17395
rect 1045 17365 1075 17395
rect 1125 17365 1155 17395
rect 1205 17365 1235 17395
rect 1285 17365 1315 17395
rect 1365 17365 1395 17395
rect 1445 17365 1475 17395
rect 1525 17365 1555 17395
rect 1605 17365 1635 17395
rect 1685 17365 1715 17395
rect 1765 17365 1795 17395
rect 1845 17365 1875 17395
rect 1925 17365 1955 17395
rect 2005 17365 2035 17395
rect 2085 17365 2115 17395
rect 2165 17365 2195 17395
rect 2245 17365 2275 17395
rect 2325 17365 2355 17395
rect 2405 17365 2435 17395
rect 2485 17365 2515 17395
rect 2565 17365 2595 17395
rect 2645 17365 2675 17395
rect 2725 17365 2755 17395
rect 2805 17365 2835 17395
rect 2885 17365 2915 17395
rect 2965 17365 2995 17395
rect 3045 17365 3075 17395
rect 3125 17365 3155 17395
rect 3205 17365 3235 17395
rect 3285 17365 3315 17395
rect 3365 17365 3395 17395
rect 3445 17365 3475 17395
rect 3525 17365 3555 17395
rect 3605 17365 3635 17395
rect 3685 17365 3715 17395
rect 3765 17365 3795 17395
rect 3845 17365 3875 17395
rect 3925 17365 3955 17395
rect 4005 17365 4035 17395
rect 4085 17365 4115 17395
rect 4165 17365 4195 17395
rect 4725 17365 4755 17395
rect 4885 17365 4915 17395
rect 5045 17365 5075 17395
rect 5205 17365 5235 17395
rect 5365 17365 5395 17395
rect 5525 17365 5555 17395
rect 5685 17365 5715 17395
rect 6245 17365 6275 17395
rect 6325 17365 6355 17395
rect 6405 17365 6435 17395
rect 6485 17365 6515 17395
rect 6565 17365 6595 17395
rect 6645 17365 6675 17395
rect 6725 17365 6755 17395
rect 6805 17365 6835 17395
rect 6885 17365 6915 17395
rect 6965 17365 6995 17395
rect 7045 17365 7075 17395
rect 7125 17365 7155 17395
rect 7205 17365 7235 17395
rect 7285 17365 7315 17395
rect 7365 17365 7395 17395
rect 7445 17365 7475 17395
rect 7525 17365 7555 17395
rect 7605 17365 7635 17395
rect 7685 17365 7715 17395
rect 7765 17365 7795 17395
rect 7845 17365 7875 17395
rect 7925 17365 7955 17395
rect 8005 17365 8035 17395
rect 8085 17365 8115 17395
rect 8165 17365 8195 17395
rect 8245 17365 8275 17395
rect 8325 17365 8355 17395
rect 8405 17365 8435 17395
rect 8485 17365 8515 17395
rect 8565 17365 8595 17395
rect 8645 17365 8675 17395
rect 8725 17365 8755 17395
rect 8805 17365 8835 17395
rect 8885 17365 8915 17395
rect 8965 17365 8995 17395
rect 9045 17365 9075 17395
rect 9125 17365 9155 17395
rect 9205 17365 9235 17395
rect 9285 17365 9315 17395
rect 9365 17365 9395 17395
rect 9445 17365 9475 17395
rect 10005 17365 10035 17395
rect 10165 17365 10195 17395
rect 10325 17365 10355 17395
rect 10485 17365 10515 17395
rect 10645 17365 10675 17395
rect 10805 17365 10835 17395
rect 10965 17365 10995 17395
rect 11565 17365 11595 17395
rect 11645 17365 11675 17395
rect 11725 17365 11755 17395
rect 11805 17365 11835 17395
rect 11885 17365 11915 17395
rect 11965 17365 11995 17395
rect 12045 17365 12075 17395
rect 12125 17365 12155 17395
rect 12205 17365 12235 17395
rect 12285 17365 12315 17395
rect 12365 17365 12395 17395
rect 12445 17365 12475 17395
rect 12525 17365 12555 17395
rect 12605 17365 12635 17395
rect 12685 17365 12715 17395
rect 12765 17365 12795 17395
rect 12845 17365 12875 17395
rect 12925 17365 12955 17395
rect 13005 17365 13035 17395
rect 13085 17365 13115 17395
rect 13165 17365 13195 17395
rect 13245 17365 13275 17395
rect 13325 17365 13355 17395
rect 13405 17365 13435 17395
rect 13485 17365 13515 17395
rect 13565 17365 13595 17395
rect 13645 17365 13675 17395
rect 13725 17365 13755 17395
rect 13805 17365 13835 17395
rect 13885 17365 13915 17395
rect 13965 17365 13995 17395
rect 14045 17365 14075 17395
rect 14125 17365 14155 17395
rect 14205 17365 14235 17395
rect 14285 17365 14315 17395
rect 14365 17365 14395 17395
rect 14445 17365 14475 17395
rect 14525 17365 14555 17395
rect 14605 17365 14635 17395
rect 14685 17365 14715 17395
rect 15245 17365 15275 17395
rect 15405 17365 15435 17395
rect 15565 17365 15595 17395
rect 15725 17365 15755 17395
rect 15885 17365 15915 17395
rect 16045 17365 16075 17395
rect 16205 17365 16235 17395
rect 16765 17365 16795 17395
rect 16845 17365 16875 17395
rect 16925 17365 16955 17395
rect 17005 17365 17035 17395
rect 17085 17365 17115 17395
rect 17165 17365 17195 17395
rect 17245 17365 17275 17395
rect 17325 17365 17355 17395
rect 17405 17365 17435 17395
rect 17485 17365 17515 17395
rect 17565 17365 17595 17395
rect 17645 17365 17675 17395
rect 17725 17365 17755 17395
rect 17805 17365 17835 17395
rect 17885 17365 17915 17395
rect 17965 17365 17995 17395
rect 18045 17365 18075 17395
rect 18125 17365 18155 17395
rect 18205 17365 18235 17395
rect 18285 17365 18315 17395
rect 18365 17365 18395 17395
rect 18445 17365 18475 17395
rect 18525 17365 18555 17395
rect 18605 17365 18635 17395
rect 18685 17365 18715 17395
rect 18765 17365 18795 17395
rect 18845 17365 18875 17395
rect 18925 17365 18955 17395
rect 19005 17365 19035 17395
rect 19085 17365 19115 17395
rect 19165 17365 19195 17395
rect 19245 17365 19275 17395
rect 19325 17365 19355 17395
rect 19405 17365 19435 17395
rect 19485 17365 19515 17395
rect 19565 17365 19595 17395
rect 19645 17365 19675 17395
rect 19725 17365 19755 17395
rect 19805 17365 19835 17395
rect 19885 17365 19915 17395
rect 19965 17365 19995 17395
rect 20045 17365 20075 17395
rect 20125 17365 20155 17395
rect 20205 17365 20235 17395
rect 20285 17365 20315 17395
rect 20365 17365 20395 17395
rect 20445 17365 20475 17395
rect 20525 17365 20555 17395
rect 20605 17365 20635 17395
rect 20685 17365 20715 17395
rect 20765 17365 20795 17395
rect 20845 17365 20875 17395
rect 20925 17365 20955 17395
rect 5605 17285 5635 17315
rect 10085 17285 10115 17315
rect 15325 17285 15355 17315
rect 5 17205 35 17235
rect 85 17205 115 17235
rect 165 17205 195 17235
rect 245 17205 275 17235
rect 325 17205 355 17235
rect 405 17205 435 17235
rect 485 17205 515 17235
rect 565 17205 595 17235
rect 645 17205 675 17235
rect 725 17205 755 17235
rect 805 17205 835 17235
rect 885 17205 915 17235
rect 965 17205 995 17235
rect 1045 17205 1075 17235
rect 1125 17205 1155 17235
rect 1205 17205 1235 17235
rect 1285 17205 1315 17235
rect 1365 17205 1395 17235
rect 1445 17205 1475 17235
rect 1525 17205 1555 17235
rect 1605 17205 1635 17235
rect 1685 17205 1715 17235
rect 1765 17205 1795 17235
rect 1845 17205 1875 17235
rect 1925 17205 1955 17235
rect 2005 17205 2035 17235
rect 2085 17205 2115 17235
rect 2165 17205 2195 17235
rect 2245 17205 2275 17235
rect 2325 17205 2355 17235
rect 2405 17205 2435 17235
rect 2485 17205 2515 17235
rect 2565 17205 2595 17235
rect 2645 17205 2675 17235
rect 2725 17205 2755 17235
rect 2805 17205 2835 17235
rect 2885 17205 2915 17235
rect 2965 17205 2995 17235
rect 3045 17205 3075 17235
rect 3125 17205 3155 17235
rect 3205 17205 3235 17235
rect 3285 17205 3315 17235
rect 3365 17205 3395 17235
rect 3445 17205 3475 17235
rect 3525 17205 3555 17235
rect 3605 17205 3635 17235
rect 3685 17205 3715 17235
rect 3765 17205 3795 17235
rect 3845 17205 3875 17235
rect 3925 17205 3955 17235
rect 4005 17205 4035 17235
rect 4085 17205 4115 17235
rect 4165 17205 4195 17235
rect 4725 17205 4755 17235
rect 4885 17205 4915 17235
rect 5045 17205 5075 17235
rect 5205 17205 5235 17235
rect 5365 17205 5395 17235
rect 5525 17205 5555 17235
rect 5685 17205 5715 17235
rect 6245 17205 6275 17235
rect 6325 17205 6355 17235
rect 6405 17205 6435 17235
rect 6485 17205 6515 17235
rect 6565 17205 6595 17235
rect 6645 17205 6675 17235
rect 6725 17205 6755 17235
rect 6805 17205 6835 17235
rect 6885 17205 6915 17235
rect 6965 17205 6995 17235
rect 7045 17205 7075 17235
rect 7125 17205 7155 17235
rect 7205 17205 7235 17235
rect 7285 17205 7315 17235
rect 7365 17205 7395 17235
rect 7445 17205 7475 17235
rect 7525 17205 7555 17235
rect 7605 17205 7635 17235
rect 7685 17205 7715 17235
rect 7765 17205 7795 17235
rect 7845 17205 7875 17235
rect 7925 17205 7955 17235
rect 8005 17205 8035 17235
rect 8085 17205 8115 17235
rect 8165 17205 8195 17235
rect 8245 17205 8275 17235
rect 8325 17205 8355 17235
rect 8405 17205 8435 17235
rect 8485 17205 8515 17235
rect 8565 17205 8595 17235
rect 8645 17205 8675 17235
rect 8725 17205 8755 17235
rect 8805 17205 8835 17235
rect 8885 17205 8915 17235
rect 8965 17205 8995 17235
rect 9045 17205 9075 17235
rect 9125 17205 9155 17235
rect 9205 17205 9235 17235
rect 9285 17205 9315 17235
rect 9365 17205 9395 17235
rect 9445 17205 9475 17235
rect 10005 17205 10035 17235
rect 10165 17205 10195 17235
rect 10325 17205 10355 17235
rect 10485 17205 10515 17235
rect 10645 17205 10675 17235
rect 10805 17205 10835 17235
rect 10965 17205 10995 17235
rect 11565 17205 11595 17235
rect 11645 17205 11675 17235
rect 11725 17205 11755 17235
rect 11805 17205 11835 17235
rect 11885 17205 11915 17235
rect 11965 17205 11995 17235
rect 12045 17205 12075 17235
rect 12125 17205 12155 17235
rect 12205 17205 12235 17235
rect 12285 17205 12315 17235
rect 12365 17205 12395 17235
rect 12445 17205 12475 17235
rect 12525 17205 12555 17235
rect 12605 17205 12635 17235
rect 12685 17205 12715 17235
rect 12765 17205 12795 17235
rect 12845 17205 12875 17235
rect 12925 17205 12955 17235
rect 13005 17205 13035 17235
rect 13085 17205 13115 17235
rect 13165 17205 13195 17235
rect 13245 17205 13275 17235
rect 13325 17205 13355 17235
rect 13405 17205 13435 17235
rect 13485 17205 13515 17235
rect 13565 17205 13595 17235
rect 13645 17205 13675 17235
rect 13725 17205 13755 17235
rect 13805 17205 13835 17235
rect 13885 17205 13915 17235
rect 13965 17205 13995 17235
rect 14045 17205 14075 17235
rect 14125 17205 14155 17235
rect 14205 17205 14235 17235
rect 14285 17205 14315 17235
rect 14365 17205 14395 17235
rect 14445 17205 14475 17235
rect 14525 17205 14555 17235
rect 14605 17205 14635 17235
rect 14685 17205 14715 17235
rect 15245 17205 15275 17235
rect 15405 17205 15435 17235
rect 15565 17205 15595 17235
rect 15725 17205 15755 17235
rect 15885 17205 15915 17235
rect 16045 17205 16075 17235
rect 16205 17205 16235 17235
rect 16765 17205 16795 17235
rect 16845 17205 16875 17235
rect 16925 17205 16955 17235
rect 17005 17205 17035 17235
rect 17085 17205 17115 17235
rect 17165 17205 17195 17235
rect 17245 17205 17275 17235
rect 17325 17205 17355 17235
rect 17405 17205 17435 17235
rect 17485 17205 17515 17235
rect 17565 17205 17595 17235
rect 17645 17205 17675 17235
rect 17725 17205 17755 17235
rect 17805 17205 17835 17235
rect 17885 17205 17915 17235
rect 17965 17205 17995 17235
rect 18045 17205 18075 17235
rect 18125 17205 18155 17235
rect 18205 17205 18235 17235
rect 18285 17205 18315 17235
rect 18365 17205 18395 17235
rect 18445 17205 18475 17235
rect 18525 17205 18555 17235
rect 18605 17205 18635 17235
rect 18685 17205 18715 17235
rect 18765 17205 18795 17235
rect 18845 17205 18875 17235
rect 18925 17205 18955 17235
rect 19005 17205 19035 17235
rect 19085 17205 19115 17235
rect 19165 17205 19195 17235
rect 19245 17205 19275 17235
rect 19325 17205 19355 17235
rect 19405 17205 19435 17235
rect 19485 17205 19515 17235
rect 19565 17205 19595 17235
rect 19645 17205 19675 17235
rect 19725 17205 19755 17235
rect 19805 17205 19835 17235
rect 19885 17205 19915 17235
rect 19965 17205 19995 17235
rect 20045 17205 20075 17235
rect 20125 17205 20155 17235
rect 20205 17205 20235 17235
rect 20285 17205 20315 17235
rect 20365 17205 20395 17235
rect 20445 17205 20475 17235
rect 20525 17205 20555 17235
rect 20605 17205 20635 17235
rect 20685 17205 20715 17235
rect 20765 17205 20795 17235
rect 20845 17205 20875 17235
rect 20925 17205 20955 17235
rect 5 17125 35 17155
rect 85 17125 115 17155
rect 165 17125 195 17155
rect 245 17125 275 17155
rect 325 17125 355 17155
rect 405 17125 435 17155
rect 485 17125 515 17155
rect 565 17125 595 17155
rect 645 17125 675 17155
rect 725 17125 755 17155
rect 805 17125 835 17155
rect 885 17125 915 17155
rect 965 17125 995 17155
rect 1045 17125 1075 17155
rect 1125 17125 1155 17155
rect 1205 17125 1235 17155
rect 1285 17125 1315 17155
rect 1365 17125 1395 17155
rect 1445 17125 1475 17155
rect 1525 17125 1555 17155
rect 1605 17125 1635 17155
rect 1685 17125 1715 17155
rect 1765 17125 1795 17155
rect 1845 17125 1875 17155
rect 1925 17125 1955 17155
rect 2005 17125 2035 17155
rect 2085 17125 2115 17155
rect 2165 17125 2195 17155
rect 2245 17125 2275 17155
rect 2325 17125 2355 17155
rect 2405 17125 2435 17155
rect 2485 17125 2515 17155
rect 2565 17125 2595 17155
rect 2645 17125 2675 17155
rect 2725 17125 2755 17155
rect 2805 17125 2835 17155
rect 2885 17125 2915 17155
rect 2965 17125 2995 17155
rect 3045 17125 3075 17155
rect 3125 17125 3155 17155
rect 3205 17125 3235 17155
rect 3285 17125 3315 17155
rect 3365 17125 3395 17155
rect 3445 17125 3475 17155
rect 3525 17125 3555 17155
rect 3605 17125 3635 17155
rect 3685 17125 3715 17155
rect 3765 17125 3795 17155
rect 3845 17125 3875 17155
rect 3925 17125 3955 17155
rect 4005 17125 4035 17155
rect 4085 17125 4115 17155
rect 4165 17125 4195 17155
rect 5765 17125 5795 17155
rect 5925 17125 5955 17155
rect 6245 17125 6275 17155
rect 6325 17125 6355 17155
rect 6405 17125 6435 17155
rect 6485 17125 6515 17155
rect 6565 17125 6595 17155
rect 6645 17125 6675 17155
rect 6725 17125 6755 17155
rect 6805 17125 6835 17155
rect 6885 17125 6915 17155
rect 6965 17125 6995 17155
rect 7045 17125 7075 17155
rect 7125 17125 7155 17155
rect 7205 17125 7235 17155
rect 7285 17125 7315 17155
rect 7365 17125 7395 17155
rect 7445 17125 7475 17155
rect 7525 17125 7555 17155
rect 7605 17125 7635 17155
rect 7685 17125 7715 17155
rect 7765 17125 7795 17155
rect 7845 17125 7875 17155
rect 7925 17125 7955 17155
rect 8005 17125 8035 17155
rect 8085 17125 8115 17155
rect 8165 17125 8195 17155
rect 8245 17125 8275 17155
rect 8325 17125 8355 17155
rect 8405 17125 8435 17155
rect 8485 17125 8515 17155
rect 8565 17125 8595 17155
rect 8645 17125 8675 17155
rect 8725 17125 8755 17155
rect 8805 17125 8835 17155
rect 8885 17125 8915 17155
rect 8965 17125 8995 17155
rect 9045 17125 9075 17155
rect 9125 17125 9155 17155
rect 9205 17125 9235 17155
rect 9285 17125 9315 17155
rect 9365 17125 9395 17155
rect 9445 17125 9475 17155
rect 9765 17125 9795 17155
rect 9925 17125 9955 17155
rect 11565 17125 11595 17155
rect 11645 17125 11675 17155
rect 11725 17125 11755 17155
rect 11805 17125 11835 17155
rect 11885 17125 11915 17155
rect 11965 17125 11995 17155
rect 12045 17125 12075 17155
rect 12125 17125 12155 17155
rect 12205 17125 12235 17155
rect 12285 17125 12315 17155
rect 12365 17125 12395 17155
rect 12445 17125 12475 17155
rect 12525 17125 12555 17155
rect 12605 17125 12635 17155
rect 12685 17125 12715 17155
rect 12765 17125 12795 17155
rect 12845 17125 12875 17155
rect 12925 17125 12955 17155
rect 13005 17125 13035 17155
rect 13085 17125 13115 17155
rect 13165 17125 13195 17155
rect 13245 17125 13275 17155
rect 13325 17125 13355 17155
rect 13405 17125 13435 17155
rect 13485 17125 13515 17155
rect 13565 17125 13595 17155
rect 13645 17125 13675 17155
rect 13725 17125 13755 17155
rect 13805 17125 13835 17155
rect 13885 17125 13915 17155
rect 13965 17125 13995 17155
rect 14045 17125 14075 17155
rect 14125 17125 14155 17155
rect 14205 17125 14235 17155
rect 14285 17125 14315 17155
rect 14365 17125 14395 17155
rect 14445 17125 14475 17155
rect 14525 17125 14555 17155
rect 14605 17125 14635 17155
rect 14685 17125 14715 17155
rect 15005 17125 15035 17155
rect 15165 17125 15195 17155
rect 16765 17125 16795 17155
rect 16845 17125 16875 17155
rect 16925 17125 16955 17155
rect 17005 17125 17035 17155
rect 17085 17125 17115 17155
rect 17165 17125 17195 17155
rect 17245 17125 17275 17155
rect 17325 17125 17355 17155
rect 17405 17125 17435 17155
rect 17485 17125 17515 17155
rect 17565 17125 17595 17155
rect 17645 17125 17675 17155
rect 17725 17125 17755 17155
rect 17805 17125 17835 17155
rect 17885 17125 17915 17155
rect 17965 17125 17995 17155
rect 18045 17125 18075 17155
rect 18125 17125 18155 17155
rect 18205 17125 18235 17155
rect 18285 17125 18315 17155
rect 18365 17125 18395 17155
rect 18445 17125 18475 17155
rect 18525 17125 18555 17155
rect 18605 17125 18635 17155
rect 18685 17125 18715 17155
rect 18765 17125 18795 17155
rect 18845 17125 18875 17155
rect 18925 17125 18955 17155
rect 19005 17125 19035 17155
rect 19085 17125 19115 17155
rect 19165 17125 19195 17155
rect 19245 17125 19275 17155
rect 19325 17125 19355 17155
rect 19405 17125 19435 17155
rect 19485 17125 19515 17155
rect 19565 17125 19595 17155
rect 19645 17125 19675 17155
rect 19725 17125 19755 17155
rect 19805 17125 19835 17155
rect 19885 17125 19915 17155
rect 19965 17125 19995 17155
rect 20045 17125 20075 17155
rect 20125 17125 20155 17155
rect 20205 17125 20235 17155
rect 20285 17125 20315 17155
rect 20365 17125 20395 17155
rect 20445 17125 20475 17155
rect 20525 17125 20555 17155
rect 20605 17125 20635 17155
rect 20685 17125 20715 17155
rect 20765 17125 20795 17155
rect 20845 17125 20875 17155
rect 20925 17125 20955 17155
rect 5845 17045 5875 17075
rect 9845 17045 9875 17075
rect 15085 17045 15115 17075
rect 5 16965 35 16995
rect 85 16965 115 16995
rect 165 16965 195 16995
rect 245 16965 275 16995
rect 325 16965 355 16995
rect 405 16965 435 16995
rect 485 16965 515 16995
rect 565 16965 595 16995
rect 645 16965 675 16995
rect 725 16965 755 16995
rect 805 16965 835 16995
rect 885 16965 915 16995
rect 965 16965 995 16995
rect 1045 16965 1075 16995
rect 1125 16965 1155 16995
rect 1205 16965 1235 16995
rect 1285 16965 1315 16995
rect 1365 16965 1395 16995
rect 1445 16965 1475 16995
rect 1525 16965 1555 16995
rect 1605 16965 1635 16995
rect 1685 16965 1715 16995
rect 1765 16965 1795 16995
rect 1845 16965 1875 16995
rect 1925 16965 1955 16995
rect 2005 16965 2035 16995
rect 2085 16965 2115 16995
rect 2165 16965 2195 16995
rect 2245 16965 2275 16995
rect 2325 16965 2355 16995
rect 2405 16965 2435 16995
rect 2485 16965 2515 16995
rect 2565 16965 2595 16995
rect 2645 16965 2675 16995
rect 2725 16965 2755 16995
rect 2805 16965 2835 16995
rect 2885 16965 2915 16995
rect 2965 16965 2995 16995
rect 3045 16965 3075 16995
rect 3125 16965 3155 16995
rect 3205 16965 3235 16995
rect 3285 16965 3315 16995
rect 3365 16965 3395 16995
rect 3445 16965 3475 16995
rect 3525 16965 3555 16995
rect 3605 16965 3635 16995
rect 3685 16965 3715 16995
rect 3765 16965 3795 16995
rect 3845 16965 3875 16995
rect 3925 16965 3955 16995
rect 4005 16965 4035 16995
rect 4085 16965 4115 16995
rect 4165 16965 4195 16995
rect 5765 16965 5795 16995
rect 5925 16965 5955 16995
rect 6245 16965 6275 16995
rect 6325 16965 6355 16995
rect 6405 16965 6435 16995
rect 6485 16965 6515 16995
rect 6565 16965 6595 16995
rect 6645 16965 6675 16995
rect 6725 16965 6755 16995
rect 6805 16965 6835 16995
rect 6885 16965 6915 16995
rect 6965 16965 6995 16995
rect 7045 16965 7075 16995
rect 7125 16965 7155 16995
rect 7205 16965 7235 16995
rect 7285 16965 7315 16995
rect 7365 16965 7395 16995
rect 7445 16965 7475 16995
rect 7525 16965 7555 16995
rect 7605 16965 7635 16995
rect 7685 16965 7715 16995
rect 7765 16965 7795 16995
rect 7845 16965 7875 16995
rect 7925 16965 7955 16995
rect 8005 16965 8035 16995
rect 8085 16965 8115 16995
rect 8165 16965 8195 16995
rect 8245 16965 8275 16995
rect 8325 16965 8355 16995
rect 8405 16965 8435 16995
rect 8485 16965 8515 16995
rect 8565 16965 8595 16995
rect 8645 16965 8675 16995
rect 8725 16965 8755 16995
rect 8805 16965 8835 16995
rect 8885 16965 8915 16995
rect 8965 16965 8995 16995
rect 9045 16965 9075 16995
rect 9125 16965 9155 16995
rect 9205 16965 9235 16995
rect 9285 16965 9315 16995
rect 9365 16965 9395 16995
rect 9445 16965 9475 16995
rect 9765 16965 9795 16995
rect 9925 16965 9955 16995
rect 11565 16965 11595 16995
rect 11645 16965 11675 16995
rect 11725 16965 11755 16995
rect 11805 16965 11835 16995
rect 11885 16965 11915 16995
rect 11965 16965 11995 16995
rect 12045 16965 12075 16995
rect 12125 16965 12155 16995
rect 12205 16965 12235 16995
rect 12285 16965 12315 16995
rect 12365 16965 12395 16995
rect 12445 16965 12475 16995
rect 12525 16965 12555 16995
rect 12605 16965 12635 16995
rect 12685 16965 12715 16995
rect 12765 16965 12795 16995
rect 12845 16965 12875 16995
rect 12925 16965 12955 16995
rect 13005 16965 13035 16995
rect 13085 16965 13115 16995
rect 13165 16965 13195 16995
rect 13245 16965 13275 16995
rect 13325 16965 13355 16995
rect 13405 16965 13435 16995
rect 13485 16965 13515 16995
rect 13565 16965 13595 16995
rect 13645 16965 13675 16995
rect 13725 16965 13755 16995
rect 13805 16965 13835 16995
rect 13885 16965 13915 16995
rect 13965 16965 13995 16995
rect 14045 16965 14075 16995
rect 14125 16965 14155 16995
rect 14205 16965 14235 16995
rect 14285 16965 14315 16995
rect 14365 16965 14395 16995
rect 14445 16965 14475 16995
rect 14525 16965 14555 16995
rect 14605 16965 14635 16995
rect 14685 16965 14715 16995
rect 15005 16965 15035 16995
rect 15165 16965 15195 16995
rect 16765 16965 16795 16995
rect 16845 16965 16875 16995
rect 16925 16965 16955 16995
rect 17005 16965 17035 16995
rect 17085 16965 17115 16995
rect 17165 16965 17195 16995
rect 17245 16965 17275 16995
rect 17325 16965 17355 16995
rect 17405 16965 17435 16995
rect 17485 16965 17515 16995
rect 17565 16965 17595 16995
rect 17645 16965 17675 16995
rect 17725 16965 17755 16995
rect 17805 16965 17835 16995
rect 17885 16965 17915 16995
rect 17965 16965 17995 16995
rect 18045 16965 18075 16995
rect 18125 16965 18155 16995
rect 18205 16965 18235 16995
rect 18285 16965 18315 16995
rect 18365 16965 18395 16995
rect 18445 16965 18475 16995
rect 18525 16965 18555 16995
rect 18605 16965 18635 16995
rect 18685 16965 18715 16995
rect 18765 16965 18795 16995
rect 18845 16965 18875 16995
rect 18925 16965 18955 16995
rect 19005 16965 19035 16995
rect 19085 16965 19115 16995
rect 19165 16965 19195 16995
rect 19245 16965 19275 16995
rect 19325 16965 19355 16995
rect 19405 16965 19435 16995
rect 19485 16965 19515 16995
rect 19565 16965 19595 16995
rect 19645 16965 19675 16995
rect 19725 16965 19755 16995
rect 19805 16965 19835 16995
rect 19885 16965 19915 16995
rect 19965 16965 19995 16995
rect 20045 16965 20075 16995
rect 20125 16965 20155 16995
rect 20205 16965 20235 16995
rect 20285 16965 20315 16995
rect 20365 16965 20395 16995
rect 20445 16965 20475 16995
rect 20525 16965 20555 16995
rect 20605 16965 20635 16995
rect 20685 16965 20715 16995
rect 20765 16965 20795 16995
rect 20845 16965 20875 16995
rect 20925 16965 20955 16995
rect 5 16885 35 16915
rect 85 16885 115 16915
rect 165 16885 195 16915
rect 245 16885 275 16915
rect 325 16885 355 16915
rect 405 16885 435 16915
rect 485 16885 515 16915
rect 565 16885 595 16915
rect 645 16885 675 16915
rect 725 16885 755 16915
rect 805 16885 835 16915
rect 885 16885 915 16915
rect 965 16885 995 16915
rect 1045 16885 1075 16915
rect 1125 16885 1155 16915
rect 1205 16885 1235 16915
rect 1285 16885 1315 16915
rect 1365 16885 1395 16915
rect 1445 16885 1475 16915
rect 1525 16885 1555 16915
rect 1605 16885 1635 16915
rect 1685 16885 1715 16915
rect 1765 16885 1795 16915
rect 1845 16885 1875 16915
rect 1925 16885 1955 16915
rect 2005 16885 2035 16915
rect 2085 16885 2115 16915
rect 2165 16885 2195 16915
rect 2245 16885 2275 16915
rect 2325 16885 2355 16915
rect 2405 16885 2435 16915
rect 2485 16885 2515 16915
rect 2565 16885 2595 16915
rect 2645 16885 2675 16915
rect 2725 16885 2755 16915
rect 2805 16885 2835 16915
rect 2885 16885 2915 16915
rect 2965 16885 2995 16915
rect 3045 16885 3075 16915
rect 3125 16885 3155 16915
rect 3205 16885 3235 16915
rect 3285 16885 3315 16915
rect 3365 16885 3395 16915
rect 3445 16885 3475 16915
rect 3525 16885 3555 16915
rect 3605 16885 3635 16915
rect 3685 16885 3715 16915
rect 3765 16885 3795 16915
rect 3845 16885 3875 16915
rect 3925 16885 3955 16915
rect 4005 16885 4035 16915
rect 4085 16885 4115 16915
rect 4165 16885 4195 16915
rect 6005 16885 6035 16915
rect 6165 16885 6195 16915
rect 6245 16885 6275 16915
rect 6325 16885 6355 16915
rect 6405 16885 6435 16915
rect 6485 16885 6515 16915
rect 6565 16885 6595 16915
rect 6645 16885 6675 16915
rect 6725 16885 6755 16915
rect 6805 16885 6835 16915
rect 6885 16885 6915 16915
rect 6965 16885 6995 16915
rect 7045 16885 7075 16915
rect 7125 16885 7155 16915
rect 7205 16885 7235 16915
rect 7285 16885 7315 16915
rect 7365 16885 7395 16915
rect 7445 16885 7475 16915
rect 7525 16885 7555 16915
rect 7605 16885 7635 16915
rect 7685 16885 7715 16915
rect 7765 16885 7795 16915
rect 7845 16885 7875 16915
rect 7925 16885 7955 16915
rect 8005 16885 8035 16915
rect 8085 16885 8115 16915
rect 8165 16885 8195 16915
rect 8245 16885 8275 16915
rect 8325 16885 8355 16915
rect 8405 16885 8435 16915
rect 8485 16885 8515 16915
rect 8565 16885 8595 16915
rect 8645 16885 8675 16915
rect 8725 16885 8755 16915
rect 8805 16885 8835 16915
rect 8885 16885 8915 16915
rect 8965 16885 8995 16915
rect 9045 16885 9075 16915
rect 9125 16885 9155 16915
rect 9205 16885 9235 16915
rect 9285 16885 9315 16915
rect 9365 16885 9395 16915
rect 9445 16885 9475 16915
rect 9525 16885 9555 16915
rect 9685 16885 9715 16915
rect 11565 16885 11595 16915
rect 11645 16885 11675 16915
rect 11725 16885 11755 16915
rect 11805 16885 11835 16915
rect 11885 16885 11915 16915
rect 11965 16885 11995 16915
rect 12045 16885 12075 16915
rect 12125 16885 12155 16915
rect 12205 16885 12235 16915
rect 12285 16885 12315 16915
rect 12365 16885 12395 16915
rect 12445 16885 12475 16915
rect 12525 16885 12555 16915
rect 12605 16885 12635 16915
rect 12685 16885 12715 16915
rect 12765 16885 12795 16915
rect 12845 16885 12875 16915
rect 12925 16885 12955 16915
rect 13005 16885 13035 16915
rect 13085 16885 13115 16915
rect 13165 16885 13195 16915
rect 13245 16885 13275 16915
rect 13325 16885 13355 16915
rect 13405 16885 13435 16915
rect 13485 16885 13515 16915
rect 13565 16885 13595 16915
rect 13645 16885 13675 16915
rect 13725 16885 13755 16915
rect 13805 16885 13835 16915
rect 13885 16885 13915 16915
rect 13965 16885 13995 16915
rect 14045 16885 14075 16915
rect 14125 16885 14155 16915
rect 14205 16885 14235 16915
rect 14285 16885 14315 16915
rect 14365 16885 14395 16915
rect 14445 16885 14475 16915
rect 14525 16885 14555 16915
rect 14605 16885 14635 16915
rect 14685 16885 14715 16915
rect 14765 16885 14795 16915
rect 14925 16885 14955 16915
rect 16765 16885 16795 16915
rect 16845 16885 16875 16915
rect 16925 16885 16955 16915
rect 17005 16885 17035 16915
rect 17085 16885 17115 16915
rect 17165 16885 17195 16915
rect 17245 16885 17275 16915
rect 17325 16885 17355 16915
rect 17405 16885 17435 16915
rect 17485 16885 17515 16915
rect 17565 16885 17595 16915
rect 17645 16885 17675 16915
rect 17725 16885 17755 16915
rect 17805 16885 17835 16915
rect 17885 16885 17915 16915
rect 17965 16885 17995 16915
rect 18045 16885 18075 16915
rect 18125 16885 18155 16915
rect 18205 16885 18235 16915
rect 18285 16885 18315 16915
rect 18365 16885 18395 16915
rect 18445 16885 18475 16915
rect 18525 16885 18555 16915
rect 18605 16885 18635 16915
rect 18685 16885 18715 16915
rect 18765 16885 18795 16915
rect 18845 16885 18875 16915
rect 18925 16885 18955 16915
rect 19005 16885 19035 16915
rect 19085 16885 19115 16915
rect 19165 16885 19195 16915
rect 19245 16885 19275 16915
rect 19325 16885 19355 16915
rect 19405 16885 19435 16915
rect 19485 16885 19515 16915
rect 19565 16885 19595 16915
rect 19645 16885 19675 16915
rect 19725 16885 19755 16915
rect 19805 16885 19835 16915
rect 19885 16885 19915 16915
rect 19965 16885 19995 16915
rect 20045 16885 20075 16915
rect 20125 16885 20155 16915
rect 20205 16885 20235 16915
rect 20285 16885 20315 16915
rect 20365 16885 20395 16915
rect 20445 16885 20475 16915
rect 20525 16885 20555 16915
rect 20605 16885 20635 16915
rect 20685 16885 20715 16915
rect 20765 16885 20795 16915
rect 20845 16885 20875 16915
rect 20925 16885 20955 16915
rect 6085 16805 6115 16835
rect 9605 16805 9635 16835
rect 14845 16805 14875 16835
rect 5 16725 35 16755
rect 85 16725 115 16755
rect 165 16725 195 16755
rect 245 16725 275 16755
rect 325 16725 355 16755
rect 405 16725 435 16755
rect 485 16725 515 16755
rect 565 16725 595 16755
rect 645 16725 675 16755
rect 725 16725 755 16755
rect 805 16725 835 16755
rect 885 16725 915 16755
rect 965 16725 995 16755
rect 1045 16725 1075 16755
rect 1125 16725 1155 16755
rect 1205 16725 1235 16755
rect 1285 16725 1315 16755
rect 1365 16725 1395 16755
rect 1445 16725 1475 16755
rect 1525 16725 1555 16755
rect 1605 16725 1635 16755
rect 1685 16725 1715 16755
rect 1765 16725 1795 16755
rect 1845 16725 1875 16755
rect 1925 16725 1955 16755
rect 2005 16725 2035 16755
rect 2085 16725 2115 16755
rect 2165 16725 2195 16755
rect 2245 16725 2275 16755
rect 2325 16725 2355 16755
rect 2405 16725 2435 16755
rect 2485 16725 2515 16755
rect 2565 16725 2595 16755
rect 2645 16725 2675 16755
rect 2725 16725 2755 16755
rect 2805 16725 2835 16755
rect 2885 16725 2915 16755
rect 2965 16725 2995 16755
rect 3045 16725 3075 16755
rect 3125 16725 3155 16755
rect 3205 16725 3235 16755
rect 3285 16725 3315 16755
rect 3365 16725 3395 16755
rect 3445 16725 3475 16755
rect 3525 16725 3555 16755
rect 3605 16725 3635 16755
rect 3685 16725 3715 16755
rect 3765 16725 3795 16755
rect 3845 16725 3875 16755
rect 3925 16725 3955 16755
rect 4005 16725 4035 16755
rect 4085 16725 4115 16755
rect 4165 16725 4195 16755
rect 6005 16725 6035 16755
rect 6165 16725 6195 16755
rect 6245 16725 6275 16755
rect 6325 16725 6355 16755
rect 6405 16725 6435 16755
rect 6485 16725 6515 16755
rect 6565 16725 6595 16755
rect 6645 16725 6675 16755
rect 6725 16725 6755 16755
rect 6805 16725 6835 16755
rect 6885 16725 6915 16755
rect 6965 16725 6995 16755
rect 7045 16725 7075 16755
rect 7125 16725 7155 16755
rect 7205 16725 7235 16755
rect 7285 16725 7315 16755
rect 7365 16725 7395 16755
rect 7445 16725 7475 16755
rect 7525 16725 7555 16755
rect 7605 16725 7635 16755
rect 7685 16725 7715 16755
rect 7765 16725 7795 16755
rect 7845 16725 7875 16755
rect 7925 16725 7955 16755
rect 8005 16725 8035 16755
rect 8085 16725 8115 16755
rect 8165 16725 8195 16755
rect 8245 16725 8275 16755
rect 8325 16725 8355 16755
rect 8405 16725 8435 16755
rect 8485 16725 8515 16755
rect 8565 16725 8595 16755
rect 8645 16725 8675 16755
rect 8725 16725 8755 16755
rect 8805 16725 8835 16755
rect 8885 16725 8915 16755
rect 8965 16725 8995 16755
rect 9045 16725 9075 16755
rect 9125 16725 9155 16755
rect 9205 16725 9235 16755
rect 9285 16725 9315 16755
rect 9365 16725 9395 16755
rect 9445 16725 9475 16755
rect 9525 16725 9555 16755
rect 9685 16725 9715 16755
rect 11565 16725 11595 16755
rect 11645 16725 11675 16755
rect 11725 16725 11755 16755
rect 11805 16725 11835 16755
rect 11885 16725 11915 16755
rect 11965 16725 11995 16755
rect 12045 16725 12075 16755
rect 12125 16725 12155 16755
rect 12205 16725 12235 16755
rect 12285 16725 12315 16755
rect 12365 16725 12395 16755
rect 12445 16725 12475 16755
rect 12525 16725 12555 16755
rect 12605 16725 12635 16755
rect 12685 16725 12715 16755
rect 12765 16725 12795 16755
rect 12845 16725 12875 16755
rect 12925 16725 12955 16755
rect 13005 16725 13035 16755
rect 13085 16725 13115 16755
rect 13165 16725 13195 16755
rect 13245 16725 13275 16755
rect 13325 16725 13355 16755
rect 13405 16725 13435 16755
rect 13485 16725 13515 16755
rect 13565 16725 13595 16755
rect 13645 16725 13675 16755
rect 13725 16725 13755 16755
rect 13805 16725 13835 16755
rect 13885 16725 13915 16755
rect 13965 16725 13995 16755
rect 14045 16725 14075 16755
rect 14125 16725 14155 16755
rect 14205 16725 14235 16755
rect 14285 16725 14315 16755
rect 14365 16725 14395 16755
rect 14445 16725 14475 16755
rect 14525 16725 14555 16755
rect 14605 16725 14635 16755
rect 14685 16725 14715 16755
rect 14765 16725 14795 16755
rect 14925 16725 14955 16755
rect 16765 16725 16795 16755
rect 16845 16725 16875 16755
rect 16925 16725 16955 16755
rect 17005 16725 17035 16755
rect 17085 16725 17115 16755
rect 17165 16725 17195 16755
rect 17245 16725 17275 16755
rect 17325 16725 17355 16755
rect 17405 16725 17435 16755
rect 17485 16725 17515 16755
rect 17565 16725 17595 16755
rect 17645 16725 17675 16755
rect 17725 16725 17755 16755
rect 17805 16725 17835 16755
rect 17885 16725 17915 16755
rect 17965 16725 17995 16755
rect 18045 16725 18075 16755
rect 18125 16725 18155 16755
rect 18205 16725 18235 16755
rect 18285 16725 18315 16755
rect 18365 16725 18395 16755
rect 18445 16725 18475 16755
rect 18525 16725 18555 16755
rect 18605 16725 18635 16755
rect 18685 16725 18715 16755
rect 18765 16725 18795 16755
rect 18845 16725 18875 16755
rect 18925 16725 18955 16755
rect 19005 16725 19035 16755
rect 19085 16725 19115 16755
rect 19165 16725 19195 16755
rect 19245 16725 19275 16755
rect 19325 16725 19355 16755
rect 19405 16725 19435 16755
rect 19485 16725 19515 16755
rect 19565 16725 19595 16755
rect 19645 16725 19675 16755
rect 19725 16725 19755 16755
rect 19805 16725 19835 16755
rect 19885 16725 19915 16755
rect 19965 16725 19995 16755
rect 20045 16725 20075 16755
rect 20125 16725 20155 16755
rect 20205 16725 20235 16755
rect 20285 16725 20315 16755
rect 20365 16725 20395 16755
rect 20445 16725 20475 16755
rect 20525 16725 20555 16755
rect 20605 16725 20635 16755
rect 20685 16725 20715 16755
rect 20765 16725 20795 16755
rect 20845 16725 20875 16755
rect 20925 16725 20955 16755
rect 5 16645 35 16675
rect 85 16645 115 16675
rect 165 16645 195 16675
rect 245 16645 275 16675
rect 325 16645 355 16675
rect 405 16645 435 16675
rect 485 16645 515 16675
rect 565 16645 595 16675
rect 645 16645 675 16675
rect 725 16645 755 16675
rect 805 16645 835 16675
rect 885 16645 915 16675
rect 965 16645 995 16675
rect 1045 16645 1075 16675
rect 1125 16645 1155 16675
rect 1205 16645 1235 16675
rect 1285 16645 1315 16675
rect 1365 16645 1395 16675
rect 1445 16645 1475 16675
rect 1525 16645 1555 16675
rect 1605 16645 1635 16675
rect 1685 16645 1715 16675
rect 1765 16645 1795 16675
rect 1845 16645 1875 16675
rect 1925 16645 1955 16675
rect 2005 16645 2035 16675
rect 2085 16645 2115 16675
rect 2165 16645 2195 16675
rect 2245 16645 2275 16675
rect 2325 16645 2355 16675
rect 2405 16645 2435 16675
rect 2485 16645 2515 16675
rect 2565 16645 2595 16675
rect 2645 16645 2675 16675
rect 2725 16645 2755 16675
rect 2805 16645 2835 16675
rect 2885 16645 2915 16675
rect 2965 16645 2995 16675
rect 3045 16645 3075 16675
rect 3125 16645 3155 16675
rect 3205 16645 3235 16675
rect 3285 16645 3315 16675
rect 3365 16645 3395 16675
rect 3445 16645 3475 16675
rect 3525 16645 3555 16675
rect 3605 16645 3635 16675
rect 3685 16645 3715 16675
rect 3765 16645 3795 16675
rect 3845 16645 3875 16675
rect 3925 16645 3955 16675
rect 4005 16645 4035 16675
rect 4085 16645 4115 16675
rect 4165 16645 4195 16675
rect 4245 16645 4275 16675
rect 4405 16645 4435 16675
rect 6245 16645 6275 16675
rect 6325 16645 6355 16675
rect 6405 16645 6435 16675
rect 6485 16645 6515 16675
rect 6565 16645 6595 16675
rect 6645 16645 6675 16675
rect 6725 16645 6755 16675
rect 6805 16645 6835 16675
rect 6885 16645 6915 16675
rect 6965 16645 6995 16675
rect 7045 16645 7075 16675
rect 7125 16645 7155 16675
rect 7205 16645 7235 16675
rect 7285 16645 7315 16675
rect 7365 16645 7395 16675
rect 7445 16645 7475 16675
rect 7525 16645 7555 16675
rect 7605 16645 7635 16675
rect 7685 16645 7715 16675
rect 7765 16645 7795 16675
rect 7845 16645 7875 16675
rect 7925 16645 7955 16675
rect 8005 16645 8035 16675
rect 8085 16645 8115 16675
rect 8165 16645 8195 16675
rect 8245 16645 8275 16675
rect 8325 16645 8355 16675
rect 8405 16645 8435 16675
rect 8485 16645 8515 16675
rect 8565 16645 8595 16675
rect 8645 16645 8675 16675
rect 8725 16645 8755 16675
rect 8805 16645 8835 16675
rect 8885 16645 8915 16675
rect 8965 16645 8995 16675
rect 9045 16645 9075 16675
rect 9125 16645 9155 16675
rect 9205 16645 9235 16675
rect 9285 16645 9315 16675
rect 9365 16645 9395 16675
rect 9445 16645 9475 16675
rect 9525 16645 9555 16675
rect 9685 16645 9715 16675
rect 11565 16645 11595 16675
rect 11645 16645 11675 16675
rect 11725 16645 11755 16675
rect 11805 16645 11835 16675
rect 11885 16645 11915 16675
rect 11965 16645 11995 16675
rect 12045 16645 12075 16675
rect 12125 16645 12155 16675
rect 12205 16645 12235 16675
rect 12285 16645 12315 16675
rect 12365 16645 12395 16675
rect 12445 16645 12475 16675
rect 12525 16645 12555 16675
rect 12605 16645 12635 16675
rect 12685 16645 12715 16675
rect 12765 16645 12795 16675
rect 12845 16645 12875 16675
rect 12925 16645 12955 16675
rect 13005 16645 13035 16675
rect 13085 16645 13115 16675
rect 13165 16645 13195 16675
rect 13245 16645 13275 16675
rect 13325 16645 13355 16675
rect 13405 16645 13435 16675
rect 13485 16645 13515 16675
rect 13565 16645 13595 16675
rect 13645 16645 13675 16675
rect 13725 16645 13755 16675
rect 13805 16645 13835 16675
rect 13885 16645 13915 16675
rect 13965 16645 13995 16675
rect 14045 16645 14075 16675
rect 14125 16645 14155 16675
rect 14205 16645 14235 16675
rect 14285 16645 14315 16675
rect 14365 16645 14395 16675
rect 14445 16645 14475 16675
rect 14525 16645 14555 16675
rect 14605 16645 14635 16675
rect 14685 16645 14715 16675
rect 16525 16645 16555 16675
rect 16685 16645 16715 16675
rect 16765 16645 16795 16675
rect 16845 16645 16875 16675
rect 16925 16645 16955 16675
rect 17005 16645 17035 16675
rect 17085 16645 17115 16675
rect 17165 16645 17195 16675
rect 17245 16645 17275 16675
rect 17325 16645 17355 16675
rect 17405 16645 17435 16675
rect 17485 16645 17515 16675
rect 17565 16645 17595 16675
rect 17645 16645 17675 16675
rect 17725 16645 17755 16675
rect 17805 16645 17835 16675
rect 17885 16645 17915 16675
rect 17965 16645 17995 16675
rect 18045 16645 18075 16675
rect 18125 16645 18155 16675
rect 18205 16645 18235 16675
rect 18285 16645 18315 16675
rect 18365 16645 18395 16675
rect 18445 16645 18475 16675
rect 18525 16645 18555 16675
rect 18605 16645 18635 16675
rect 18685 16645 18715 16675
rect 18765 16645 18795 16675
rect 18845 16645 18875 16675
rect 18925 16645 18955 16675
rect 19005 16645 19035 16675
rect 19085 16645 19115 16675
rect 19165 16645 19195 16675
rect 19245 16645 19275 16675
rect 19325 16645 19355 16675
rect 19405 16645 19435 16675
rect 19485 16645 19515 16675
rect 19565 16645 19595 16675
rect 19645 16645 19675 16675
rect 19725 16645 19755 16675
rect 19805 16645 19835 16675
rect 19885 16645 19915 16675
rect 19965 16645 19995 16675
rect 20045 16645 20075 16675
rect 20125 16645 20155 16675
rect 20205 16645 20235 16675
rect 20285 16645 20315 16675
rect 20365 16645 20395 16675
rect 20445 16645 20475 16675
rect 20525 16645 20555 16675
rect 20605 16645 20635 16675
rect 20685 16645 20715 16675
rect 20765 16645 20795 16675
rect 20845 16645 20875 16675
rect 20925 16645 20955 16675
rect 4325 16565 4355 16595
rect 9605 16565 9635 16595
rect 16605 16565 16635 16595
rect 5 16485 35 16515
rect 85 16485 115 16515
rect 165 16485 195 16515
rect 245 16485 275 16515
rect 325 16485 355 16515
rect 405 16485 435 16515
rect 485 16485 515 16515
rect 565 16485 595 16515
rect 645 16485 675 16515
rect 725 16485 755 16515
rect 805 16485 835 16515
rect 885 16485 915 16515
rect 965 16485 995 16515
rect 1045 16485 1075 16515
rect 1125 16485 1155 16515
rect 1205 16485 1235 16515
rect 1285 16485 1315 16515
rect 1365 16485 1395 16515
rect 1445 16485 1475 16515
rect 1525 16485 1555 16515
rect 1605 16485 1635 16515
rect 1685 16485 1715 16515
rect 1765 16485 1795 16515
rect 1845 16485 1875 16515
rect 1925 16485 1955 16515
rect 2005 16485 2035 16515
rect 2085 16485 2115 16515
rect 2165 16485 2195 16515
rect 2245 16485 2275 16515
rect 2325 16485 2355 16515
rect 2405 16485 2435 16515
rect 2485 16485 2515 16515
rect 2565 16485 2595 16515
rect 2645 16485 2675 16515
rect 2725 16485 2755 16515
rect 2805 16485 2835 16515
rect 2885 16485 2915 16515
rect 2965 16485 2995 16515
rect 3045 16485 3075 16515
rect 3125 16485 3155 16515
rect 3205 16485 3235 16515
rect 3285 16485 3315 16515
rect 3365 16485 3395 16515
rect 3445 16485 3475 16515
rect 3525 16485 3555 16515
rect 3605 16485 3635 16515
rect 3685 16485 3715 16515
rect 3765 16485 3795 16515
rect 3845 16485 3875 16515
rect 3925 16485 3955 16515
rect 4005 16485 4035 16515
rect 4085 16485 4115 16515
rect 4165 16485 4195 16515
rect 4245 16485 4275 16515
rect 4405 16485 4435 16515
rect 6245 16485 6275 16515
rect 6325 16485 6355 16515
rect 6405 16485 6435 16515
rect 6485 16485 6515 16515
rect 6565 16485 6595 16515
rect 6645 16485 6675 16515
rect 6725 16485 6755 16515
rect 6805 16485 6835 16515
rect 6885 16485 6915 16515
rect 6965 16485 6995 16515
rect 7045 16485 7075 16515
rect 7125 16485 7155 16515
rect 7205 16485 7235 16515
rect 7285 16485 7315 16515
rect 7365 16485 7395 16515
rect 7445 16485 7475 16515
rect 7525 16485 7555 16515
rect 7605 16485 7635 16515
rect 7685 16485 7715 16515
rect 7765 16485 7795 16515
rect 7845 16485 7875 16515
rect 7925 16485 7955 16515
rect 8005 16485 8035 16515
rect 8085 16485 8115 16515
rect 8165 16485 8195 16515
rect 8245 16485 8275 16515
rect 8325 16485 8355 16515
rect 8405 16485 8435 16515
rect 8485 16485 8515 16515
rect 8565 16485 8595 16515
rect 8645 16485 8675 16515
rect 8725 16485 8755 16515
rect 8805 16485 8835 16515
rect 8885 16485 8915 16515
rect 8965 16485 8995 16515
rect 9045 16485 9075 16515
rect 9125 16485 9155 16515
rect 9205 16485 9235 16515
rect 9285 16485 9315 16515
rect 9365 16485 9395 16515
rect 9445 16485 9475 16515
rect 9525 16485 9555 16515
rect 9685 16485 9715 16515
rect 11565 16485 11595 16515
rect 11645 16485 11675 16515
rect 11725 16485 11755 16515
rect 11805 16485 11835 16515
rect 11885 16485 11915 16515
rect 11965 16485 11995 16515
rect 12045 16485 12075 16515
rect 12125 16485 12155 16515
rect 12205 16485 12235 16515
rect 12285 16485 12315 16515
rect 12365 16485 12395 16515
rect 12445 16485 12475 16515
rect 12525 16485 12555 16515
rect 12605 16485 12635 16515
rect 12685 16485 12715 16515
rect 12765 16485 12795 16515
rect 12845 16485 12875 16515
rect 12925 16485 12955 16515
rect 13005 16485 13035 16515
rect 13085 16485 13115 16515
rect 13165 16485 13195 16515
rect 13245 16485 13275 16515
rect 13325 16485 13355 16515
rect 13405 16485 13435 16515
rect 13485 16485 13515 16515
rect 13565 16485 13595 16515
rect 13645 16485 13675 16515
rect 13725 16485 13755 16515
rect 13805 16485 13835 16515
rect 13885 16485 13915 16515
rect 13965 16485 13995 16515
rect 14045 16485 14075 16515
rect 14125 16485 14155 16515
rect 14205 16485 14235 16515
rect 14285 16485 14315 16515
rect 14365 16485 14395 16515
rect 14445 16485 14475 16515
rect 14525 16485 14555 16515
rect 14605 16485 14635 16515
rect 14685 16485 14715 16515
rect 16525 16485 16555 16515
rect 16685 16485 16715 16515
rect 16765 16485 16795 16515
rect 16845 16485 16875 16515
rect 16925 16485 16955 16515
rect 17005 16485 17035 16515
rect 17085 16485 17115 16515
rect 17165 16485 17195 16515
rect 17245 16485 17275 16515
rect 17325 16485 17355 16515
rect 17405 16485 17435 16515
rect 17485 16485 17515 16515
rect 17565 16485 17595 16515
rect 17645 16485 17675 16515
rect 17725 16485 17755 16515
rect 17805 16485 17835 16515
rect 17885 16485 17915 16515
rect 17965 16485 17995 16515
rect 18045 16485 18075 16515
rect 18125 16485 18155 16515
rect 18205 16485 18235 16515
rect 18285 16485 18315 16515
rect 18365 16485 18395 16515
rect 18445 16485 18475 16515
rect 18525 16485 18555 16515
rect 18605 16485 18635 16515
rect 18685 16485 18715 16515
rect 18765 16485 18795 16515
rect 18845 16485 18875 16515
rect 18925 16485 18955 16515
rect 19005 16485 19035 16515
rect 19085 16485 19115 16515
rect 19165 16485 19195 16515
rect 19245 16485 19275 16515
rect 19325 16485 19355 16515
rect 19405 16485 19435 16515
rect 19485 16485 19515 16515
rect 19565 16485 19595 16515
rect 19645 16485 19675 16515
rect 19725 16485 19755 16515
rect 19805 16485 19835 16515
rect 19885 16485 19915 16515
rect 19965 16485 19995 16515
rect 20045 16485 20075 16515
rect 20125 16485 20155 16515
rect 20205 16485 20235 16515
rect 20285 16485 20315 16515
rect 20365 16485 20395 16515
rect 20445 16485 20475 16515
rect 20525 16485 20555 16515
rect 20605 16485 20635 16515
rect 20685 16485 20715 16515
rect 20765 16485 20795 16515
rect 20845 16485 20875 16515
rect 20925 16485 20955 16515
rect 5 16405 35 16435
rect 85 16405 115 16435
rect 165 16405 195 16435
rect 245 16405 275 16435
rect 325 16405 355 16435
rect 405 16405 435 16435
rect 485 16405 515 16435
rect 565 16405 595 16435
rect 645 16405 675 16435
rect 725 16405 755 16435
rect 805 16405 835 16435
rect 885 16405 915 16435
rect 965 16405 995 16435
rect 1045 16405 1075 16435
rect 1125 16405 1155 16435
rect 1205 16405 1235 16435
rect 1285 16405 1315 16435
rect 1365 16405 1395 16435
rect 1445 16405 1475 16435
rect 1525 16405 1555 16435
rect 1605 16405 1635 16435
rect 1685 16405 1715 16435
rect 1765 16405 1795 16435
rect 1845 16405 1875 16435
rect 1925 16405 1955 16435
rect 2005 16405 2035 16435
rect 2085 16405 2115 16435
rect 2165 16405 2195 16435
rect 2245 16405 2275 16435
rect 2325 16405 2355 16435
rect 2405 16405 2435 16435
rect 2485 16405 2515 16435
rect 2565 16405 2595 16435
rect 2645 16405 2675 16435
rect 2725 16405 2755 16435
rect 2805 16405 2835 16435
rect 2885 16405 2915 16435
rect 2965 16405 2995 16435
rect 3045 16405 3075 16435
rect 3125 16405 3155 16435
rect 3205 16405 3235 16435
rect 3285 16405 3315 16435
rect 3365 16405 3395 16435
rect 3445 16405 3475 16435
rect 3525 16405 3555 16435
rect 3605 16405 3635 16435
rect 3685 16405 3715 16435
rect 3765 16405 3795 16435
rect 3845 16405 3875 16435
rect 3925 16405 3955 16435
rect 4005 16405 4035 16435
rect 4085 16405 4115 16435
rect 4165 16405 4195 16435
rect 4485 16405 4515 16435
rect 4645 16405 4675 16435
rect 6245 16405 6275 16435
rect 6325 16405 6355 16435
rect 6405 16405 6435 16435
rect 6485 16405 6515 16435
rect 6565 16405 6595 16435
rect 6645 16405 6675 16435
rect 6725 16405 6755 16435
rect 6805 16405 6835 16435
rect 6885 16405 6915 16435
rect 6965 16405 6995 16435
rect 7045 16405 7075 16435
rect 7125 16405 7155 16435
rect 7205 16405 7235 16435
rect 7285 16405 7315 16435
rect 7365 16405 7395 16435
rect 7445 16405 7475 16435
rect 7525 16405 7555 16435
rect 7605 16405 7635 16435
rect 7685 16405 7715 16435
rect 7765 16405 7795 16435
rect 7845 16405 7875 16435
rect 7925 16405 7955 16435
rect 8005 16405 8035 16435
rect 8085 16405 8115 16435
rect 8165 16405 8195 16435
rect 8245 16405 8275 16435
rect 8325 16405 8355 16435
rect 8405 16405 8435 16435
rect 8485 16405 8515 16435
rect 8565 16405 8595 16435
rect 8645 16405 8675 16435
rect 8725 16405 8755 16435
rect 8805 16405 8835 16435
rect 8885 16405 8915 16435
rect 8965 16405 8995 16435
rect 9045 16405 9075 16435
rect 9125 16405 9155 16435
rect 9205 16405 9235 16435
rect 9285 16405 9315 16435
rect 9365 16405 9395 16435
rect 9445 16405 9475 16435
rect 9765 16405 9795 16435
rect 9925 16405 9955 16435
rect 11565 16405 11595 16435
rect 11645 16405 11675 16435
rect 11725 16405 11755 16435
rect 11805 16405 11835 16435
rect 11885 16405 11915 16435
rect 11965 16405 11995 16435
rect 12045 16405 12075 16435
rect 12125 16405 12155 16435
rect 12205 16405 12235 16435
rect 12285 16405 12315 16435
rect 12365 16405 12395 16435
rect 12445 16405 12475 16435
rect 12525 16405 12555 16435
rect 12605 16405 12635 16435
rect 12685 16405 12715 16435
rect 12765 16405 12795 16435
rect 12845 16405 12875 16435
rect 12925 16405 12955 16435
rect 13005 16405 13035 16435
rect 13085 16405 13115 16435
rect 13165 16405 13195 16435
rect 13245 16405 13275 16435
rect 13325 16405 13355 16435
rect 13405 16405 13435 16435
rect 13485 16405 13515 16435
rect 13565 16405 13595 16435
rect 13645 16405 13675 16435
rect 13725 16405 13755 16435
rect 13805 16405 13835 16435
rect 13885 16405 13915 16435
rect 13965 16405 13995 16435
rect 14045 16405 14075 16435
rect 14125 16405 14155 16435
rect 14205 16405 14235 16435
rect 14285 16405 14315 16435
rect 14365 16405 14395 16435
rect 14445 16405 14475 16435
rect 14525 16405 14555 16435
rect 14605 16405 14635 16435
rect 14685 16405 14715 16435
rect 16285 16405 16315 16435
rect 16445 16405 16475 16435
rect 16765 16405 16795 16435
rect 16845 16405 16875 16435
rect 16925 16405 16955 16435
rect 17005 16405 17035 16435
rect 17085 16405 17115 16435
rect 17165 16405 17195 16435
rect 17245 16405 17275 16435
rect 17325 16405 17355 16435
rect 17405 16405 17435 16435
rect 17485 16405 17515 16435
rect 17565 16405 17595 16435
rect 17645 16405 17675 16435
rect 17725 16405 17755 16435
rect 17805 16405 17835 16435
rect 17885 16405 17915 16435
rect 17965 16405 17995 16435
rect 18045 16405 18075 16435
rect 18125 16405 18155 16435
rect 18205 16405 18235 16435
rect 18285 16405 18315 16435
rect 18365 16405 18395 16435
rect 18445 16405 18475 16435
rect 18525 16405 18555 16435
rect 18605 16405 18635 16435
rect 18685 16405 18715 16435
rect 18765 16405 18795 16435
rect 18845 16405 18875 16435
rect 18925 16405 18955 16435
rect 19005 16405 19035 16435
rect 19085 16405 19115 16435
rect 19165 16405 19195 16435
rect 19245 16405 19275 16435
rect 19325 16405 19355 16435
rect 19405 16405 19435 16435
rect 19485 16405 19515 16435
rect 19565 16405 19595 16435
rect 19645 16405 19675 16435
rect 19725 16405 19755 16435
rect 19805 16405 19835 16435
rect 19885 16405 19915 16435
rect 19965 16405 19995 16435
rect 20045 16405 20075 16435
rect 20125 16405 20155 16435
rect 20205 16405 20235 16435
rect 20285 16405 20315 16435
rect 20365 16405 20395 16435
rect 20445 16405 20475 16435
rect 20525 16405 20555 16435
rect 20605 16405 20635 16435
rect 20685 16405 20715 16435
rect 20765 16405 20795 16435
rect 20845 16405 20875 16435
rect 20925 16405 20955 16435
rect 4565 16325 4595 16355
rect 9845 16325 9875 16355
rect 16365 16325 16395 16355
rect 5 16245 35 16275
rect 85 16245 115 16275
rect 165 16245 195 16275
rect 245 16245 275 16275
rect 325 16245 355 16275
rect 405 16245 435 16275
rect 485 16245 515 16275
rect 565 16245 595 16275
rect 645 16245 675 16275
rect 725 16245 755 16275
rect 805 16245 835 16275
rect 885 16245 915 16275
rect 965 16245 995 16275
rect 1045 16245 1075 16275
rect 1125 16245 1155 16275
rect 1205 16245 1235 16275
rect 1285 16245 1315 16275
rect 1365 16245 1395 16275
rect 1445 16245 1475 16275
rect 1525 16245 1555 16275
rect 1605 16245 1635 16275
rect 1685 16245 1715 16275
rect 1765 16245 1795 16275
rect 1845 16245 1875 16275
rect 1925 16245 1955 16275
rect 2005 16245 2035 16275
rect 2085 16245 2115 16275
rect 2165 16245 2195 16275
rect 2245 16245 2275 16275
rect 2325 16245 2355 16275
rect 2405 16245 2435 16275
rect 2485 16245 2515 16275
rect 2565 16245 2595 16275
rect 2645 16245 2675 16275
rect 2725 16245 2755 16275
rect 2805 16245 2835 16275
rect 2885 16245 2915 16275
rect 2965 16245 2995 16275
rect 3045 16245 3075 16275
rect 3125 16245 3155 16275
rect 3205 16245 3235 16275
rect 3285 16245 3315 16275
rect 3365 16245 3395 16275
rect 3445 16245 3475 16275
rect 3525 16245 3555 16275
rect 3605 16245 3635 16275
rect 3685 16245 3715 16275
rect 3765 16245 3795 16275
rect 3845 16245 3875 16275
rect 3925 16245 3955 16275
rect 4005 16245 4035 16275
rect 4085 16245 4115 16275
rect 4165 16245 4195 16275
rect 4485 16245 4515 16275
rect 4645 16245 4675 16275
rect 6245 16245 6275 16275
rect 6325 16245 6355 16275
rect 6405 16245 6435 16275
rect 6485 16245 6515 16275
rect 6565 16245 6595 16275
rect 6645 16245 6675 16275
rect 6725 16245 6755 16275
rect 6805 16245 6835 16275
rect 6885 16245 6915 16275
rect 6965 16245 6995 16275
rect 7045 16245 7075 16275
rect 7125 16245 7155 16275
rect 7205 16245 7235 16275
rect 7285 16245 7315 16275
rect 7365 16245 7395 16275
rect 7445 16245 7475 16275
rect 7525 16245 7555 16275
rect 7605 16245 7635 16275
rect 7685 16245 7715 16275
rect 7765 16245 7795 16275
rect 7845 16245 7875 16275
rect 7925 16245 7955 16275
rect 8005 16245 8035 16275
rect 8085 16245 8115 16275
rect 8165 16245 8195 16275
rect 8245 16245 8275 16275
rect 8325 16245 8355 16275
rect 8405 16245 8435 16275
rect 8485 16245 8515 16275
rect 8565 16245 8595 16275
rect 8645 16245 8675 16275
rect 8725 16245 8755 16275
rect 8805 16245 8835 16275
rect 8885 16245 8915 16275
rect 8965 16245 8995 16275
rect 9045 16245 9075 16275
rect 9125 16245 9155 16275
rect 9205 16245 9235 16275
rect 9285 16245 9315 16275
rect 9365 16245 9395 16275
rect 9445 16245 9475 16275
rect 9765 16245 9795 16275
rect 9925 16245 9955 16275
rect 11565 16245 11595 16275
rect 11645 16245 11675 16275
rect 11725 16245 11755 16275
rect 11805 16245 11835 16275
rect 11885 16245 11915 16275
rect 11965 16245 11995 16275
rect 12045 16245 12075 16275
rect 12125 16245 12155 16275
rect 12205 16245 12235 16275
rect 12285 16245 12315 16275
rect 12365 16245 12395 16275
rect 12445 16245 12475 16275
rect 12525 16245 12555 16275
rect 12605 16245 12635 16275
rect 12685 16245 12715 16275
rect 12765 16245 12795 16275
rect 12845 16245 12875 16275
rect 12925 16245 12955 16275
rect 13005 16245 13035 16275
rect 13085 16245 13115 16275
rect 13165 16245 13195 16275
rect 13245 16245 13275 16275
rect 13325 16245 13355 16275
rect 13405 16245 13435 16275
rect 13485 16245 13515 16275
rect 13565 16245 13595 16275
rect 13645 16245 13675 16275
rect 13725 16245 13755 16275
rect 13805 16245 13835 16275
rect 13885 16245 13915 16275
rect 13965 16245 13995 16275
rect 14045 16245 14075 16275
rect 14125 16245 14155 16275
rect 14205 16245 14235 16275
rect 14285 16245 14315 16275
rect 14365 16245 14395 16275
rect 14445 16245 14475 16275
rect 14525 16245 14555 16275
rect 14605 16245 14635 16275
rect 14685 16245 14715 16275
rect 16285 16245 16315 16275
rect 16445 16245 16475 16275
rect 16765 16245 16795 16275
rect 16845 16245 16875 16275
rect 16925 16245 16955 16275
rect 17005 16245 17035 16275
rect 17085 16245 17115 16275
rect 17165 16245 17195 16275
rect 17245 16245 17275 16275
rect 17325 16245 17355 16275
rect 17405 16245 17435 16275
rect 17485 16245 17515 16275
rect 17565 16245 17595 16275
rect 17645 16245 17675 16275
rect 17725 16245 17755 16275
rect 17805 16245 17835 16275
rect 17885 16245 17915 16275
rect 17965 16245 17995 16275
rect 18045 16245 18075 16275
rect 18125 16245 18155 16275
rect 18205 16245 18235 16275
rect 18285 16245 18315 16275
rect 18365 16245 18395 16275
rect 18445 16245 18475 16275
rect 18525 16245 18555 16275
rect 18605 16245 18635 16275
rect 18685 16245 18715 16275
rect 18765 16245 18795 16275
rect 18845 16245 18875 16275
rect 18925 16245 18955 16275
rect 19005 16245 19035 16275
rect 19085 16245 19115 16275
rect 19165 16245 19195 16275
rect 19245 16245 19275 16275
rect 19325 16245 19355 16275
rect 19405 16245 19435 16275
rect 19485 16245 19515 16275
rect 19565 16245 19595 16275
rect 19645 16245 19675 16275
rect 19725 16245 19755 16275
rect 19805 16245 19835 16275
rect 19885 16245 19915 16275
rect 19965 16245 19995 16275
rect 20045 16245 20075 16275
rect 20125 16245 20155 16275
rect 20205 16245 20235 16275
rect 20285 16245 20315 16275
rect 20365 16245 20395 16275
rect 20445 16245 20475 16275
rect 20525 16245 20555 16275
rect 20605 16245 20635 16275
rect 20685 16245 20715 16275
rect 20765 16245 20795 16275
rect 20845 16245 20875 16275
rect 20925 16245 20955 16275
rect 5 16165 35 16195
rect 85 16165 115 16195
rect 165 16165 195 16195
rect 245 16165 275 16195
rect 325 16165 355 16195
rect 405 16165 435 16195
rect 485 16165 515 16195
rect 565 16165 595 16195
rect 645 16165 675 16195
rect 725 16165 755 16195
rect 805 16165 835 16195
rect 885 16165 915 16195
rect 965 16165 995 16195
rect 1045 16165 1075 16195
rect 1125 16165 1155 16195
rect 1205 16165 1235 16195
rect 1285 16165 1315 16195
rect 1365 16165 1395 16195
rect 1445 16165 1475 16195
rect 1525 16165 1555 16195
rect 1605 16165 1635 16195
rect 1685 16165 1715 16195
rect 1765 16165 1795 16195
rect 1845 16165 1875 16195
rect 1925 16165 1955 16195
rect 2005 16165 2035 16195
rect 2085 16165 2115 16195
rect 2165 16165 2195 16195
rect 2245 16165 2275 16195
rect 2325 16165 2355 16195
rect 2405 16165 2435 16195
rect 2485 16165 2515 16195
rect 2565 16165 2595 16195
rect 2645 16165 2675 16195
rect 2725 16165 2755 16195
rect 2805 16165 2835 16195
rect 2885 16165 2915 16195
rect 2965 16165 2995 16195
rect 3045 16165 3075 16195
rect 3125 16165 3155 16195
rect 3205 16165 3235 16195
rect 3285 16165 3315 16195
rect 3365 16165 3395 16195
rect 3445 16165 3475 16195
rect 3525 16165 3555 16195
rect 3605 16165 3635 16195
rect 3685 16165 3715 16195
rect 3765 16165 3795 16195
rect 3845 16165 3875 16195
rect 3925 16165 3955 16195
rect 4005 16165 4035 16195
rect 4085 16165 4115 16195
rect 4165 16165 4195 16195
rect 4725 16165 4755 16195
rect 4885 16165 4915 16195
rect 5045 16165 5075 16195
rect 5205 16165 5235 16195
rect 5365 16165 5395 16195
rect 5525 16165 5555 16195
rect 5685 16165 5715 16195
rect 6245 16165 6275 16195
rect 6325 16165 6355 16195
rect 6405 16165 6435 16195
rect 6485 16165 6515 16195
rect 6565 16165 6595 16195
rect 6645 16165 6675 16195
rect 6725 16165 6755 16195
rect 6805 16165 6835 16195
rect 6885 16165 6915 16195
rect 6965 16165 6995 16195
rect 7045 16165 7075 16195
rect 7125 16165 7155 16195
rect 7205 16165 7235 16195
rect 7285 16165 7315 16195
rect 7365 16165 7395 16195
rect 7445 16165 7475 16195
rect 7525 16165 7555 16195
rect 7605 16165 7635 16195
rect 7685 16165 7715 16195
rect 7765 16165 7795 16195
rect 7845 16165 7875 16195
rect 7925 16165 7955 16195
rect 8005 16165 8035 16195
rect 8085 16165 8115 16195
rect 8165 16165 8195 16195
rect 8245 16165 8275 16195
rect 8325 16165 8355 16195
rect 8405 16165 8435 16195
rect 8485 16165 8515 16195
rect 8565 16165 8595 16195
rect 8645 16165 8675 16195
rect 8725 16165 8755 16195
rect 8805 16165 8835 16195
rect 8885 16165 8915 16195
rect 8965 16165 8995 16195
rect 9045 16165 9075 16195
rect 9125 16165 9155 16195
rect 9205 16165 9235 16195
rect 9285 16165 9315 16195
rect 9365 16165 9395 16195
rect 9445 16165 9475 16195
rect 10005 16165 10035 16195
rect 10165 16165 10195 16195
rect 10325 16165 10355 16195
rect 10485 16165 10515 16195
rect 10645 16165 10675 16195
rect 10805 16165 10835 16195
rect 10965 16165 10995 16195
rect 11565 16165 11595 16195
rect 11645 16165 11675 16195
rect 11725 16165 11755 16195
rect 11805 16165 11835 16195
rect 11885 16165 11915 16195
rect 11965 16165 11995 16195
rect 12045 16165 12075 16195
rect 12125 16165 12155 16195
rect 12205 16165 12235 16195
rect 12285 16165 12315 16195
rect 12365 16165 12395 16195
rect 12445 16165 12475 16195
rect 12525 16165 12555 16195
rect 12605 16165 12635 16195
rect 12685 16165 12715 16195
rect 12765 16165 12795 16195
rect 12845 16165 12875 16195
rect 12925 16165 12955 16195
rect 13005 16165 13035 16195
rect 13085 16165 13115 16195
rect 13165 16165 13195 16195
rect 13245 16165 13275 16195
rect 13325 16165 13355 16195
rect 13405 16165 13435 16195
rect 13485 16165 13515 16195
rect 13565 16165 13595 16195
rect 13645 16165 13675 16195
rect 13725 16165 13755 16195
rect 13805 16165 13835 16195
rect 13885 16165 13915 16195
rect 13965 16165 13995 16195
rect 14045 16165 14075 16195
rect 14125 16165 14155 16195
rect 14205 16165 14235 16195
rect 14285 16165 14315 16195
rect 14365 16165 14395 16195
rect 14445 16165 14475 16195
rect 14525 16165 14555 16195
rect 14605 16165 14635 16195
rect 14685 16165 14715 16195
rect 15245 16165 15275 16195
rect 15405 16165 15435 16195
rect 15565 16165 15595 16195
rect 15725 16165 15755 16195
rect 15885 16165 15915 16195
rect 16045 16165 16075 16195
rect 16205 16165 16235 16195
rect 16765 16165 16795 16195
rect 16845 16165 16875 16195
rect 16925 16165 16955 16195
rect 17005 16165 17035 16195
rect 17085 16165 17115 16195
rect 17165 16165 17195 16195
rect 17245 16165 17275 16195
rect 17325 16165 17355 16195
rect 17405 16165 17435 16195
rect 17485 16165 17515 16195
rect 17565 16165 17595 16195
rect 17645 16165 17675 16195
rect 17725 16165 17755 16195
rect 17805 16165 17835 16195
rect 17885 16165 17915 16195
rect 17965 16165 17995 16195
rect 18045 16165 18075 16195
rect 18125 16165 18155 16195
rect 18205 16165 18235 16195
rect 18285 16165 18315 16195
rect 18365 16165 18395 16195
rect 18445 16165 18475 16195
rect 18525 16165 18555 16195
rect 18605 16165 18635 16195
rect 18685 16165 18715 16195
rect 18765 16165 18795 16195
rect 18845 16165 18875 16195
rect 18925 16165 18955 16195
rect 19005 16165 19035 16195
rect 19085 16165 19115 16195
rect 19165 16165 19195 16195
rect 19245 16165 19275 16195
rect 19325 16165 19355 16195
rect 19405 16165 19435 16195
rect 19485 16165 19515 16195
rect 19565 16165 19595 16195
rect 19645 16165 19675 16195
rect 19725 16165 19755 16195
rect 19805 16165 19835 16195
rect 19885 16165 19915 16195
rect 19965 16165 19995 16195
rect 20045 16165 20075 16195
rect 20125 16165 20155 16195
rect 20205 16165 20235 16195
rect 20285 16165 20315 16195
rect 20365 16165 20395 16195
rect 20445 16165 20475 16195
rect 20525 16165 20555 16195
rect 20605 16165 20635 16195
rect 20685 16165 20715 16195
rect 20765 16165 20795 16195
rect 20845 16165 20875 16195
rect 20925 16165 20955 16195
rect 4805 16085 4835 16115
rect 10085 16085 10115 16115
rect 16125 16085 16155 16115
rect 5 16005 35 16035
rect 85 16005 115 16035
rect 165 16005 195 16035
rect 245 16005 275 16035
rect 325 16005 355 16035
rect 405 16005 435 16035
rect 485 16005 515 16035
rect 565 16005 595 16035
rect 645 16005 675 16035
rect 725 16005 755 16035
rect 805 16005 835 16035
rect 885 16005 915 16035
rect 965 16005 995 16035
rect 1045 16005 1075 16035
rect 1125 16005 1155 16035
rect 1205 16005 1235 16035
rect 1285 16005 1315 16035
rect 1365 16005 1395 16035
rect 1445 16005 1475 16035
rect 1525 16005 1555 16035
rect 1605 16005 1635 16035
rect 1685 16005 1715 16035
rect 1765 16005 1795 16035
rect 1845 16005 1875 16035
rect 1925 16005 1955 16035
rect 2005 16005 2035 16035
rect 2085 16005 2115 16035
rect 2165 16005 2195 16035
rect 2245 16005 2275 16035
rect 2325 16005 2355 16035
rect 2405 16005 2435 16035
rect 2485 16005 2515 16035
rect 2565 16005 2595 16035
rect 2645 16005 2675 16035
rect 2725 16005 2755 16035
rect 2805 16005 2835 16035
rect 2885 16005 2915 16035
rect 2965 16005 2995 16035
rect 3045 16005 3075 16035
rect 3125 16005 3155 16035
rect 3205 16005 3235 16035
rect 3285 16005 3315 16035
rect 3365 16005 3395 16035
rect 3445 16005 3475 16035
rect 3525 16005 3555 16035
rect 3605 16005 3635 16035
rect 3685 16005 3715 16035
rect 3765 16005 3795 16035
rect 3845 16005 3875 16035
rect 3925 16005 3955 16035
rect 4005 16005 4035 16035
rect 4085 16005 4115 16035
rect 4165 16005 4195 16035
rect 4725 16005 4755 16035
rect 4885 16005 4915 16035
rect 5045 16005 5075 16035
rect 5205 16005 5235 16035
rect 5365 16005 5395 16035
rect 5525 16005 5555 16035
rect 5685 16005 5715 16035
rect 6245 16005 6275 16035
rect 6325 16005 6355 16035
rect 6405 16005 6435 16035
rect 6485 16005 6515 16035
rect 6565 16005 6595 16035
rect 6645 16005 6675 16035
rect 6725 16005 6755 16035
rect 6805 16005 6835 16035
rect 6885 16005 6915 16035
rect 6965 16005 6995 16035
rect 7045 16005 7075 16035
rect 7125 16005 7155 16035
rect 7205 16005 7235 16035
rect 7285 16005 7315 16035
rect 7365 16005 7395 16035
rect 7445 16005 7475 16035
rect 7525 16005 7555 16035
rect 7605 16005 7635 16035
rect 7685 16005 7715 16035
rect 7765 16005 7795 16035
rect 7845 16005 7875 16035
rect 7925 16005 7955 16035
rect 8005 16005 8035 16035
rect 8085 16005 8115 16035
rect 8165 16005 8195 16035
rect 8245 16005 8275 16035
rect 8325 16005 8355 16035
rect 8405 16005 8435 16035
rect 8485 16005 8515 16035
rect 8565 16005 8595 16035
rect 8645 16005 8675 16035
rect 8725 16005 8755 16035
rect 8805 16005 8835 16035
rect 8885 16005 8915 16035
rect 8965 16005 8995 16035
rect 9045 16005 9075 16035
rect 9125 16005 9155 16035
rect 9205 16005 9235 16035
rect 9285 16005 9315 16035
rect 9365 16005 9395 16035
rect 9445 16005 9475 16035
rect 10005 16005 10035 16035
rect 10165 16005 10195 16035
rect 10325 16005 10355 16035
rect 10485 16005 10515 16035
rect 10645 16005 10675 16035
rect 10805 16005 10835 16035
rect 10965 16005 10995 16035
rect 11565 16005 11595 16035
rect 11645 16005 11675 16035
rect 11725 16005 11755 16035
rect 11805 16005 11835 16035
rect 11885 16005 11915 16035
rect 11965 16005 11995 16035
rect 12045 16005 12075 16035
rect 12125 16005 12155 16035
rect 12205 16005 12235 16035
rect 12285 16005 12315 16035
rect 12365 16005 12395 16035
rect 12445 16005 12475 16035
rect 12525 16005 12555 16035
rect 12605 16005 12635 16035
rect 12685 16005 12715 16035
rect 12765 16005 12795 16035
rect 12845 16005 12875 16035
rect 12925 16005 12955 16035
rect 13005 16005 13035 16035
rect 13085 16005 13115 16035
rect 13165 16005 13195 16035
rect 13245 16005 13275 16035
rect 13325 16005 13355 16035
rect 13405 16005 13435 16035
rect 13485 16005 13515 16035
rect 13565 16005 13595 16035
rect 13645 16005 13675 16035
rect 13725 16005 13755 16035
rect 13805 16005 13835 16035
rect 13885 16005 13915 16035
rect 13965 16005 13995 16035
rect 14045 16005 14075 16035
rect 14125 16005 14155 16035
rect 14205 16005 14235 16035
rect 14285 16005 14315 16035
rect 14365 16005 14395 16035
rect 14445 16005 14475 16035
rect 14525 16005 14555 16035
rect 14605 16005 14635 16035
rect 14685 16005 14715 16035
rect 15245 16005 15275 16035
rect 15405 16005 15435 16035
rect 15565 16005 15595 16035
rect 15725 16005 15755 16035
rect 15885 16005 15915 16035
rect 16045 16005 16075 16035
rect 16205 16005 16235 16035
rect 16765 16005 16795 16035
rect 16845 16005 16875 16035
rect 16925 16005 16955 16035
rect 17005 16005 17035 16035
rect 17085 16005 17115 16035
rect 17165 16005 17195 16035
rect 17245 16005 17275 16035
rect 17325 16005 17355 16035
rect 17405 16005 17435 16035
rect 17485 16005 17515 16035
rect 17565 16005 17595 16035
rect 17645 16005 17675 16035
rect 17725 16005 17755 16035
rect 17805 16005 17835 16035
rect 17885 16005 17915 16035
rect 17965 16005 17995 16035
rect 18045 16005 18075 16035
rect 18125 16005 18155 16035
rect 18205 16005 18235 16035
rect 18285 16005 18315 16035
rect 18365 16005 18395 16035
rect 18445 16005 18475 16035
rect 18525 16005 18555 16035
rect 18605 16005 18635 16035
rect 18685 16005 18715 16035
rect 18765 16005 18795 16035
rect 18845 16005 18875 16035
rect 18925 16005 18955 16035
rect 19005 16005 19035 16035
rect 19085 16005 19115 16035
rect 19165 16005 19195 16035
rect 19245 16005 19275 16035
rect 19325 16005 19355 16035
rect 19405 16005 19435 16035
rect 19485 16005 19515 16035
rect 19565 16005 19595 16035
rect 19645 16005 19675 16035
rect 19725 16005 19755 16035
rect 19805 16005 19835 16035
rect 19885 16005 19915 16035
rect 19965 16005 19995 16035
rect 20045 16005 20075 16035
rect 20125 16005 20155 16035
rect 20205 16005 20235 16035
rect 20285 16005 20315 16035
rect 20365 16005 20395 16035
rect 20445 16005 20475 16035
rect 20525 16005 20555 16035
rect 20605 16005 20635 16035
rect 20685 16005 20715 16035
rect 20765 16005 20795 16035
rect 20845 16005 20875 16035
rect 20925 16005 20955 16035
rect 4965 15925 4995 15955
rect 10245 15925 10275 15955
rect 15965 15925 15995 15955
rect 5 15845 35 15875
rect 85 15845 115 15875
rect 165 15845 195 15875
rect 245 15845 275 15875
rect 325 15845 355 15875
rect 405 15845 435 15875
rect 485 15845 515 15875
rect 565 15845 595 15875
rect 645 15845 675 15875
rect 725 15845 755 15875
rect 805 15845 835 15875
rect 885 15845 915 15875
rect 965 15845 995 15875
rect 1045 15845 1075 15875
rect 1125 15845 1155 15875
rect 1205 15845 1235 15875
rect 1285 15845 1315 15875
rect 1365 15845 1395 15875
rect 1445 15845 1475 15875
rect 1525 15845 1555 15875
rect 1605 15845 1635 15875
rect 1685 15845 1715 15875
rect 1765 15845 1795 15875
rect 1845 15845 1875 15875
rect 1925 15845 1955 15875
rect 2005 15845 2035 15875
rect 2085 15845 2115 15875
rect 2165 15845 2195 15875
rect 2245 15845 2275 15875
rect 2325 15845 2355 15875
rect 2405 15845 2435 15875
rect 2485 15845 2515 15875
rect 2565 15845 2595 15875
rect 2645 15845 2675 15875
rect 2725 15845 2755 15875
rect 2805 15845 2835 15875
rect 2885 15845 2915 15875
rect 2965 15845 2995 15875
rect 3045 15845 3075 15875
rect 3125 15845 3155 15875
rect 3205 15845 3235 15875
rect 3285 15845 3315 15875
rect 3365 15845 3395 15875
rect 3445 15845 3475 15875
rect 3525 15845 3555 15875
rect 3605 15845 3635 15875
rect 3685 15845 3715 15875
rect 3765 15845 3795 15875
rect 3845 15845 3875 15875
rect 3925 15845 3955 15875
rect 4005 15845 4035 15875
rect 4085 15845 4115 15875
rect 4165 15845 4195 15875
rect 4725 15845 4755 15875
rect 4885 15845 4915 15875
rect 5045 15845 5075 15875
rect 5205 15845 5235 15875
rect 5365 15845 5395 15875
rect 5525 15845 5555 15875
rect 5685 15845 5715 15875
rect 6245 15845 6275 15875
rect 6325 15845 6355 15875
rect 6405 15845 6435 15875
rect 6485 15845 6515 15875
rect 6565 15845 6595 15875
rect 6645 15845 6675 15875
rect 6725 15845 6755 15875
rect 6805 15845 6835 15875
rect 6885 15845 6915 15875
rect 6965 15845 6995 15875
rect 7045 15845 7075 15875
rect 7125 15845 7155 15875
rect 7205 15845 7235 15875
rect 7285 15845 7315 15875
rect 7365 15845 7395 15875
rect 7445 15845 7475 15875
rect 7525 15845 7555 15875
rect 7605 15845 7635 15875
rect 7685 15845 7715 15875
rect 7765 15845 7795 15875
rect 7845 15845 7875 15875
rect 7925 15845 7955 15875
rect 8005 15845 8035 15875
rect 8085 15845 8115 15875
rect 8165 15845 8195 15875
rect 8245 15845 8275 15875
rect 8325 15845 8355 15875
rect 8405 15845 8435 15875
rect 8485 15845 8515 15875
rect 8565 15845 8595 15875
rect 8645 15845 8675 15875
rect 8725 15845 8755 15875
rect 8805 15845 8835 15875
rect 8885 15845 8915 15875
rect 8965 15845 8995 15875
rect 9045 15845 9075 15875
rect 9125 15845 9155 15875
rect 9205 15845 9235 15875
rect 9285 15845 9315 15875
rect 9365 15845 9395 15875
rect 9445 15845 9475 15875
rect 10005 15845 10035 15875
rect 10165 15845 10195 15875
rect 10325 15845 10355 15875
rect 10485 15845 10515 15875
rect 10645 15845 10675 15875
rect 10805 15845 10835 15875
rect 10965 15845 10995 15875
rect 11565 15845 11595 15875
rect 11645 15845 11675 15875
rect 11725 15845 11755 15875
rect 11805 15845 11835 15875
rect 11885 15845 11915 15875
rect 11965 15845 11995 15875
rect 12045 15845 12075 15875
rect 12125 15845 12155 15875
rect 12205 15845 12235 15875
rect 12285 15845 12315 15875
rect 12365 15845 12395 15875
rect 12445 15845 12475 15875
rect 12525 15845 12555 15875
rect 12605 15845 12635 15875
rect 12685 15845 12715 15875
rect 12765 15845 12795 15875
rect 12845 15845 12875 15875
rect 12925 15845 12955 15875
rect 13005 15845 13035 15875
rect 13085 15845 13115 15875
rect 13165 15845 13195 15875
rect 13245 15845 13275 15875
rect 13325 15845 13355 15875
rect 13405 15845 13435 15875
rect 13485 15845 13515 15875
rect 13565 15845 13595 15875
rect 13645 15845 13675 15875
rect 13725 15845 13755 15875
rect 13805 15845 13835 15875
rect 13885 15845 13915 15875
rect 13965 15845 13995 15875
rect 14045 15845 14075 15875
rect 14125 15845 14155 15875
rect 14205 15845 14235 15875
rect 14285 15845 14315 15875
rect 14365 15845 14395 15875
rect 14445 15845 14475 15875
rect 14525 15845 14555 15875
rect 14605 15845 14635 15875
rect 14685 15845 14715 15875
rect 15245 15845 15275 15875
rect 15405 15845 15435 15875
rect 15565 15845 15595 15875
rect 15725 15845 15755 15875
rect 15885 15845 15915 15875
rect 16045 15845 16075 15875
rect 16205 15845 16235 15875
rect 16765 15845 16795 15875
rect 16845 15845 16875 15875
rect 16925 15845 16955 15875
rect 17005 15845 17035 15875
rect 17085 15845 17115 15875
rect 17165 15845 17195 15875
rect 17245 15845 17275 15875
rect 17325 15845 17355 15875
rect 17405 15845 17435 15875
rect 17485 15845 17515 15875
rect 17565 15845 17595 15875
rect 17645 15845 17675 15875
rect 17725 15845 17755 15875
rect 17805 15845 17835 15875
rect 17885 15845 17915 15875
rect 17965 15845 17995 15875
rect 18045 15845 18075 15875
rect 18125 15845 18155 15875
rect 18205 15845 18235 15875
rect 18285 15845 18315 15875
rect 18365 15845 18395 15875
rect 18445 15845 18475 15875
rect 18525 15845 18555 15875
rect 18605 15845 18635 15875
rect 18685 15845 18715 15875
rect 18765 15845 18795 15875
rect 18845 15845 18875 15875
rect 18925 15845 18955 15875
rect 19005 15845 19035 15875
rect 19085 15845 19115 15875
rect 19165 15845 19195 15875
rect 19245 15845 19275 15875
rect 19325 15845 19355 15875
rect 19405 15845 19435 15875
rect 19485 15845 19515 15875
rect 19565 15845 19595 15875
rect 19645 15845 19675 15875
rect 19725 15845 19755 15875
rect 19805 15845 19835 15875
rect 19885 15845 19915 15875
rect 19965 15845 19995 15875
rect 20045 15845 20075 15875
rect 20125 15845 20155 15875
rect 20205 15845 20235 15875
rect 20285 15845 20315 15875
rect 20365 15845 20395 15875
rect 20445 15845 20475 15875
rect 20525 15845 20555 15875
rect 20605 15845 20635 15875
rect 20685 15845 20715 15875
rect 20765 15845 20795 15875
rect 20845 15845 20875 15875
rect 20925 15845 20955 15875
rect 5125 15765 5155 15795
rect 10405 15765 10435 15795
rect 15805 15765 15835 15795
rect 5 15685 35 15715
rect 85 15685 115 15715
rect 165 15685 195 15715
rect 245 15685 275 15715
rect 325 15685 355 15715
rect 405 15685 435 15715
rect 485 15685 515 15715
rect 565 15685 595 15715
rect 645 15685 675 15715
rect 725 15685 755 15715
rect 805 15685 835 15715
rect 885 15685 915 15715
rect 965 15685 995 15715
rect 1045 15685 1075 15715
rect 1125 15685 1155 15715
rect 1205 15685 1235 15715
rect 1285 15685 1315 15715
rect 1365 15685 1395 15715
rect 1445 15685 1475 15715
rect 1525 15685 1555 15715
rect 1605 15685 1635 15715
rect 1685 15685 1715 15715
rect 1765 15685 1795 15715
rect 1845 15685 1875 15715
rect 1925 15685 1955 15715
rect 2005 15685 2035 15715
rect 2085 15685 2115 15715
rect 2165 15685 2195 15715
rect 2245 15685 2275 15715
rect 2325 15685 2355 15715
rect 2405 15685 2435 15715
rect 2485 15685 2515 15715
rect 2565 15685 2595 15715
rect 2645 15685 2675 15715
rect 2725 15685 2755 15715
rect 2805 15685 2835 15715
rect 2885 15685 2915 15715
rect 2965 15685 2995 15715
rect 3045 15685 3075 15715
rect 3125 15685 3155 15715
rect 3205 15685 3235 15715
rect 3285 15685 3315 15715
rect 3365 15685 3395 15715
rect 3445 15685 3475 15715
rect 3525 15685 3555 15715
rect 3605 15685 3635 15715
rect 3685 15685 3715 15715
rect 3765 15685 3795 15715
rect 3845 15685 3875 15715
rect 3925 15685 3955 15715
rect 4005 15685 4035 15715
rect 4085 15685 4115 15715
rect 4165 15685 4195 15715
rect 4725 15685 4755 15715
rect 4885 15685 4915 15715
rect 5045 15685 5075 15715
rect 5205 15685 5235 15715
rect 5365 15685 5395 15715
rect 5525 15685 5555 15715
rect 5685 15685 5715 15715
rect 6245 15685 6275 15715
rect 6325 15685 6355 15715
rect 6405 15685 6435 15715
rect 6485 15685 6515 15715
rect 6565 15685 6595 15715
rect 6645 15685 6675 15715
rect 6725 15685 6755 15715
rect 6805 15685 6835 15715
rect 6885 15685 6915 15715
rect 6965 15685 6995 15715
rect 7045 15685 7075 15715
rect 7125 15685 7155 15715
rect 7205 15685 7235 15715
rect 7285 15685 7315 15715
rect 7365 15685 7395 15715
rect 7445 15685 7475 15715
rect 7525 15685 7555 15715
rect 7605 15685 7635 15715
rect 7685 15685 7715 15715
rect 7765 15685 7795 15715
rect 7845 15685 7875 15715
rect 7925 15685 7955 15715
rect 8005 15685 8035 15715
rect 8085 15685 8115 15715
rect 8165 15685 8195 15715
rect 8245 15685 8275 15715
rect 8325 15685 8355 15715
rect 8405 15685 8435 15715
rect 8485 15685 8515 15715
rect 8565 15685 8595 15715
rect 8645 15685 8675 15715
rect 8725 15685 8755 15715
rect 8805 15685 8835 15715
rect 8885 15685 8915 15715
rect 8965 15685 8995 15715
rect 9045 15685 9075 15715
rect 9125 15685 9155 15715
rect 9205 15685 9235 15715
rect 9285 15685 9315 15715
rect 9365 15685 9395 15715
rect 9445 15685 9475 15715
rect 10005 15685 10035 15715
rect 10165 15685 10195 15715
rect 10325 15685 10355 15715
rect 10485 15685 10515 15715
rect 10645 15685 10675 15715
rect 10805 15685 10835 15715
rect 10965 15685 10995 15715
rect 11565 15685 11595 15715
rect 11645 15685 11675 15715
rect 11725 15685 11755 15715
rect 11805 15685 11835 15715
rect 11885 15685 11915 15715
rect 11965 15685 11995 15715
rect 12045 15685 12075 15715
rect 12125 15685 12155 15715
rect 12205 15685 12235 15715
rect 12285 15685 12315 15715
rect 12365 15685 12395 15715
rect 12445 15685 12475 15715
rect 12525 15685 12555 15715
rect 12605 15685 12635 15715
rect 12685 15685 12715 15715
rect 12765 15685 12795 15715
rect 12845 15685 12875 15715
rect 12925 15685 12955 15715
rect 13005 15685 13035 15715
rect 13085 15685 13115 15715
rect 13165 15685 13195 15715
rect 13245 15685 13275 15715
rect 13325 15685 13355 15715
rect 13405 15685 13435 15715
rect 13485 15685 13515 15715
rect 13565 15685 13595 15715
rect 13645 15685 13675 15715
rect 13725 15685 13755 15715
rect 13805 15685 13835 15715
rect 13885 15685 13915 15715
rect 13965 15685 13995 15715
rect 14045 15685 14075 15715
rect 14125 15685 14155 15715
rect 14205 15685 14235 15715
rect 14285 15685 14315 15715
rect 14365 15685 14395 15715
rect 14445 15685 14475 15715
rect 14525 15685 14555 15715
rect 14605 15685 14635 15715
rect 14685 15685 14715 15715
rect 15245 15685 15275 15715
rect 15405 15685 15435 15715
rect 15565 15685 15595 15715
rect 15725 15685 15755 15715
rect 15885 15685 15915 15715
rect 16045 15685 16075 15715
rect 16205 15685 16235 15715
rect 16765 15685 16795 15715
rect 16845 15685 16875 15715
rect 16925 15685 16955 15715
rect 17005 15685 17035 15715
rect 17085 15685 17115 15715
rect 17165 15685 17195 15715
rect 17245 15685 17275 15715
rect 17325 15685 17355 15715
rect 17405 15685 17435 15715
rect 17485 15685 17515 15715
rect 17565 15685 17595 15715
rect 17645 15685 17675 15715
rect 17725 15685 17755 15715
rect 17805 15685 17835 15715
rect 17885 15685 17915 15715
rect 17965 15685 17995 15715
rect 18045 15685 18075 15715
rect 18125 15685 18155 15715
rect 18205 15685 18235 15715
rect 18285 15685 18315 15715
rect 18365 15685 18395 15715
rect 18445 15685 18475 15715
rect 18525 15685 18555 15715
rect 18605 15685 18635 15715
rect 18685 15685 18715 15715
rect 18765 15685 18795 15715
rect 18845 15685 18875 15715
rect 18925 15685 18955 15715
rect 19005 15685 19035 15715
rect 19085 15685 19115 15715
rect 19165 15685 19195 15715
rect 19245 15685 19275 15715
rect 19325 15685 19355 15715
rect 19405 15685 19435 15715
rect 19485 15685 19515 15715
rect 19565 15685 19595 15715
rect 19645 15685 19675 15715
rect 19725 15685 19755 15715
rect 19805 15685 19835 15715
rect 19885 15685 19915 15715
rect 19965 15685 19995 15715
rect 20045 15685 20075 15715
rect 20125 15685 20155 15715
rect 20205 15685 20235 15715
rect 20285 15685 20315 15715
rect 20365 15685 20395 15715
rect 20445 15685 20475 15715
rect 20525 15685 20555 15715
rect 20605 15685 20635 15715
rect 20685 15685 20715 15715
rect 20765 15685 20795 15715
rect 20845 15685 20875 15715
rect 20925 15685 20955 15715
rect 5285 15605 5315 15635
rect 10565 15605 10595 15635
rect 15645 15605 15675 15635
rect 5 15525 35 15555
rect 85 15525 115 15555
rect 165 15525 195 15555
rect 245 15525 275 15555
rect 325 15525 355 15555
rect 405 15525 435 15555
rect 485 15525 515 15555
rect 565 15525 595 15555
rect 645 15525 675 15555
rect 725 15525 755 15555
rect 805 15525 835 15555
rect 885 15525 915 15555
rect 965 15525 995 15555
rect 1045 15525 1075 15555
rect 1125 15525 1155 15555
rect 1205 15525 1235 15555
rect 1285 15525 1315 15555
rect 1365 15525 1395 15555
rect 1445 15525 1475 15555
rect 1525 15525 1555 15555
rect 1605 15525 1635 15555
rect 1685 15525 1715 15555
rect 1765 15525 1795 15555
rect 1845 15525 1875 15555
rect 1925 15525 1955 15555
rect 2005 15525 2035 15555
rect 2085 15525 2115 15555
rect 2165 15525 2195 15555
rect 2245 15525 2275 15555
rect 2325 15525 2355 15555
rect 2405 15525 2435 15555
rect 2485 15525 2515 15555
rect 2565 15525 2595 15555
rect 2645 15525 2675 15555
rect 2725 15525 2755 15555
rect 2805 15525 2835 15555
rect 2885 15525 2915 15555
rect 2965 15525 2995 15555
rect 3045 15525 3075 15555
rect 3125 15525 3155 15555
rect 3205 15525 3235 15555
rect 3285 15525 3315 15555
rect 3365 15525 3395 15555
rect 3445 15525 3475 15555
rect 3525 15525 3555 15555
rect 3605 15525 3635 15555
rect 3685 15525 3715 15555
rect 3765 15525 3795 15555
rect 3845 15525 3875 15555
rect 3925 15525 3955 15555
rect 4005 15525 4035 15555
rect 4085 15525 4115 15555
rect 4165 15525 4195 15555
rect 4725 15525 4755 15555
rect 4885 15525 4915 15555
rect 5045 15525 5075 15555
rect 5205 15525 5235 15555
rect 5365 15525 5395 15555
rect 5525 15525 5555 15555
rect 5685 15525 5715 15555
rect 6245 15525 6275 15555
rect 6325 15525 6355 15555
rect 6405 15525 6435 15555
rect 6485 15525 6515 15555
rect 6565 15525 6595 15555
rect 6645 15525 6675 15555
rect 6725 15525 6755 15555
rect 6805 15525 6835 15555
rect 6885 15525 6915 15555
rect 6965 15525 6995 15555
rect 7045 15525 7075 15555
rect 7125 15525 7155 15555
rect 7205 15525 7235 15555
rect 7285 15525 7315 15555
rect 7365 15525 7395 15555
rect 7445 15525 7475 15555
rect 7525 15525 7555 15555
rect 7605 15525 7635 15555
rect 7685 15525 7715 15555
rect 7765 15525 7795 15555
rect 7845 15525 7875 15555
rect 7925 15525 7955 15555
rect 8005 15525 8035 15555
rect 8085 15525 8115 15555
rect 8165 15525 8195 15555
rect 8245 15525 8275 15555
rect 8325 15525 8355 15555
rect 8405 15525 8435 15555
rect 8485 15525 8515 15555
rect 8565 15525 8595 15555
rect 8645 15525 8675 15555
rect 8725 15525 8755 15555
rect 8805 15525 8835 15555
rect 8885 15525 8915 15555
rect 8965 15525 8995 15555
rect 9045 15525 9075 15555
rect 9125 15525 9155 15555
rect 9205 15525 9235 15555
rect 9285 15525 9315 15555
rect 9365 15525 9395 15555
rect 9445 15525 9475 15555
rect 10005 15525 10035 15555
rect 10165 15525 10195 15555
rect 10325 15525 10355 15555
rect 10485 15525 10515 15555
rect 10645 15525 10675 15555
rect 10805 15525 10835 15555
rect 10965 15525 10995 15555
rect 11565 15525 11595 15555
rect 11645 15525 11675 15555
rect 11725 15525 11755 15555
rect 11805 15525 11835 15555
rect 11885 15525 11915 15555
rect 11965 15525 11995 15555
rect 12045 15525 12075 15555
rect 12125 15525 12155 15555
rect 12205 15525 12235 15555
rect 12285 15525 12315 15555
rect 12365 15525 12395 15555
rect 12445 15525 12475 15555
rect 12525 15525 12555 15555
rect 12605 15525 12635 15555
rect 12685 15525 12715 15555
rect 12765 15525 12795 15555
rect 12845 15525 12875 15555
rect 12925 15525 12955 15555
rect 13005 15525 13035 15555
rect 13085 15525 13115 15555
rect 13165 15525 13195 15555
rect 13245 15525 13275 15555
rect 13325 15525 13355 15555
rect 13405 15525 13435 15555
rect 13485 15525 13515 15555
rect 13565 15525 13595 15555
rect 13645 15525 13675 15555
rect 13725 15525 13755 15555
rect 13805 15525 13835 15555
rect 13885 15525 13915 15555
rect 13965 15525 13995 15555
rect 14045 15525 14075 15555
rect 14125 15525 14155 15555
rect 14205 15525 14235 15555
rect 14285 15525 14315 15555
rect 14365 15525 14395 15555
rect 14445 15525 14475 15555
rect 14525 15525 14555 15555
rect 14605 15525 14635 15555
rect 14685 15525 14715 15555
rect 15245 15525 15275 15555
rect 15405 15525 15435 15555
rect 15565 15525 15595 15555
rect 15725 15525 15755 15555
rect 15885 15525 15915 15555
rect 16045 15525 16075 15555
rect 16205 15525 16235 15555
rect 16765 15525 16795 15555
rect 16845 15525 16875 15555
rect 16925 15525 16955 15555
rect 17005 15525 17035 15555
rect 17085 15525 17115 15555
rect 17165 15525 17195 15555
rect 17245 15525 17275 15555
rect 17325 15525 17355 15555
rect 17405 15525 17435 15555
rect 17485 15525 17515 15555
rect 17565 15525 17595 15555
rect 17645 15525 17675 15555
rect 17725 15525 17755 15555
rect 17805 15525 17835 15555
rect 17885 15525 17915 15555
rect 17965 15525 17995 15555
rect 18045 15525 18075 15555
rect 18125 15525 18155 15555
rect 18205 15525 18235 15555
rect 18285 15525 18315 15555
rect 18365 15525 18395 15555
rect 18445 15525 18475 15555
rect 18525 15525 18555 15555
rect 18605 15525 18635 15555
rect 18685 15525 18715 15555
rect 18765 15525 18795 15555
rect 18845 15525 18875 15555
rect 18925 15525 18955 15555
rect 19005 15525 19035 15555
rect 19085 15525 19115 15555
rect 19165 15525 19195 15555
rect 19245 15525 19275 15555
rect 19325 15525 19355 15555
rect 19405 15525 19435 15555
rect 19485 15525 19515 15555
rect 19565 15525 19595 15555
rect 19645 15525 19675 15555
rect 19725 15525 19755 15555
rect 19805 15525 19835 15555
rect 19885 15525 19915 15555
rect 19965 15525 19995 15555
rect 20045 15525 20075 15555
rect 20125 15525 20155 15555
rect 20205 15525 20235 15555
rect 20285 15525 20315 15555
rect 20365 15525 20395 15555
rect 20445 15525 20475 15555
rect 20525 15525 20555 15555
rect 20605 15525 20635 15555
rect 20685 15525 20715 15555
rect 20765 15525 20795 15555
rect 20845 15525 20875 15555
rect 20925 15525 20955 15555
rect 5445 15445 5475 15475
rect 10725 15445 10755 15475
rect 15485 15445 15515 15475
rect 5 15365 35 15395
rect 85 15365 115 15395
rect 165 15365 195 15395
rect 245 15365 275 15395
rect 325 15365 355 15395
rect 405 15365 435 15395
rect 485 15365 515 15395
rect 565 15365 595 15395
rect 645 15365 675 15395
rect 725 15365 755 15395
rect 805 15365 835 15395
rect 885 15365 915 15395
rect 965 15365 995 15395
rect 1045 15365 1075 15395
rect 1125 15365 1155 15395
rect 1205 15365 1235 15395
rect 1285 15365 1315 15395
rect 1365 15365 1395 15395
rect 1445 15365 1475 15395
rect 1525 15365 1555 15395
rect 1605 15365 1635 15395
rect 1685 15365 1715 15395
rect 1765 15365 1795 15395
rect 1845 15365 1875 15395
rect 1925 15365 1955 15395
rect 2005 15365 2035 15395
rect 2085 15365 2115 15395
rect 2165 15365 2195 15395
rect 2245 15365 2275 15395
rect 2325 15365 2355 15395
rect 2405 15365 2435 15395
rect 2485 15365 2515 15395
rect 2565 15365 2595 15395
rect 2645 15365 2675 15395
rect 2725 15365 2755 15395
rect 2805 15365 2835 15395
rect 2885 15365 2915 15395
rect 2965 15365 2995 15395
rect 3045 15365 3075 15395
rect 3125 15365 3155 15395
rect 3205 15365 3235 15395
rect 3285 15365 3315 15395
rect 3365 15365 3395 15395
rect 3445 15365 3475 15395
rect 3525 15365 3555 15395
rect 3605 15365 3635 15395
rect 3685 15365 3715 15395
rect 3765 15365 3795 15395
rect 3845 15365 3875 15395
rect 3925 15365 3955 15395
rect 4005 15365 4035 15395
rect 4085 15365 4115 15395
rect 4165 15365 4195 15395
rect 4725 15365 4755 15395
rect 4885 15365 4915 15395
rect 5045 15365 5075 15395
rect 5205 15365 5235 15395
rect 5365 15365 5395 15395
rect 5525 15365 5555 15395
rect 5685 15365 5715 15395
rect 6245 15365 6275 15395
rect 6325 15365 6355 15395
rect 6405 15365 6435 15395
rect 6485 15365 6515 15395
rect 6565 15365 6595 15395
rect 6645 15365 6675 15395
rect 6725 15365 6755 15395
rect 6805 15365 6835 15395
rect 6885 15365 6915 15395
rect 6965 15365 6995 15395
rect 7045 15365 7075 15395
rect 7125 15365 7155 15395
rect 7205 15365 7235 15395
rect 7285 15365 7315 15395
rect 7365 15365 7395 15395
rect 7445 15365 7475 15395
rect 7525 15365 7555 15395
rect 7605 15365 7635 15395
rect 7685 15365 7715 15395
rect 7765 15365 7795 15395
rect 7845 15365 7875 15395
rect 7925 15365 7955 15395
rect 8005 15365 8035 15395
rect 8085 15365 8115 15395
rect 8165 15365 8195 15395
rect 8245 15365 8275 15395
rect 8325 15365 8355 15395
rect 8405 15365 8435 15395
rect 8485 15365 8515 15395
rect 8565 15365 8595 15395
rect 8645 15365 8675 15395
rect 8725 15365 8755 15395
rect 8805 15365 8835 15395
rect 8885 15365 8915 15395
rect 8965 15365 8995 15395
rect 9045 15365 9075 15395
rect 9125 15365 9155 15395
rect 9205 15365 9235 15395
rect 9285 15365 9315 15395
rect 9365 15365 9395 15395
rect 9445 15365 9475 15395
rect 10005 15365 10035 15395
rect 10165 15365 10195 15395
rect 10325 15365 10355 15395
rect 10485 15365 10515 15395
rect 10645 15365 10675 15395
rect 10805 15365 10835 15395
rect 10965 15365 10995 15395
rect 11565 15365 11595 15395
rect 11645 15365 11675 15395
rect 11725 15365 11755 15395
rect 11805 15365 11835 15395
rect 11885 15365 11915 15395
rect 11965 15365 11995 15395
rect 12045 15365 12075 15395
rect 12125 15365 12155 15395
rect 12205 15365 12235 15395
rect 12285 15365 12315 15395
rect 12365 15365 12395 15395
rect 12445 15365 12475 15395
rect 12525 15365 12555 15395
rect 12605 15365 12635 15395
rect 12685 15365 12715 15395
rect 12765 15365 12795 15395
rect 12845 15365 12875 15395
rect 12925 15365 12955 15395
rect 13005 15365 13035 15395
rect 13085 15365 13115 15395
rect 13165 15365 13195 15395
rect 13245 15365 13275 15395
rect 13325 15365 13355 15395
rect 13405 15365 13435 15395
rect 13485 15365 13515 15395
rect 13565 15365 13595 15395
rect 13645 15365 13675 15395
rect 13725 15365 13755 15395
rect 13805 15365 13835 15395
rect 13885 15365 13915 15395
rect 13965 15365 13995 15395
rect 14045 15365 14075 15395
rect 14125 15365 14155 15395
rect 14205 15365 14235 15395
rect 14285 15365 14315 15395
rect 14365 15365 14395 15395
rect 14445 15365 14475 15395
rect 14525 15365 14555 15395
rect 14605 15365 14635 15395
rect 14685 15365 14715 15395
rect 15245 15365 15275 15395
rect 15405 15365 15435 15395
rect 15565 15365 15595 15395
rect 15725 15365 15755 15395
rect 15885 15365 15915 15395
rect 16045 15365 16075 15395
rect 16205 15365 16235 15395
rect 16765 15365 16795 15395
rect 16845 15365 16875 15395
rect 16925 15365 16955 15395
rect 17005 15365 17035 15395
rect 17085 15365 17115 15395
rect 17165 15365 17195 15395
rect 17245 15365 17275 15395
rect 17325 15365 17355 15395
rect 17405 15365 17435 15395
rect 17485 15365 17515 15395
rect 17565 15365 17595 15395
rect 17645 15365 17675 15395
rect 17725 15365 17755 15395
rect 17805 15365 17835 15395
rect 17885 15365 17915 15395
rect 17965 15365 17995 15395
rect 18045 15365 18075 15395
rect 18125 15365 18155 15395
rect 18205 15365 18235 15395
rect 18285 15365 18315 15395
rect 18365 15365 18395 15395
rect 18445 15365 18475 15395
rect 18525 15365 18555 15395
rect 18605 15365 18635 15395
rect 18685 15365 18715 15395
rect 18765 15365 18795 15395
rect 18845 15365 18875 15395
rect 18925 15365 18955 15395
rect 19005 15365 19035 15395
rect 19085 15365 19115 15395
rect 19165 15365 19195 15395
rect 19245 15365 19275 15395
rect 19325 15365 19355 15395
rect 19405 15365 19435 15395
rect 19485 15365 19515 15395
rect 19565 15365 19595 15395
rect 19645 15365 19675 15395
rect 19725 15365 19755 15395
rect 19805 15365 19835 15395
rect 19885 15365 19915 15395
rect 19965 15365 19995 15395
rect 20045 15365 20075 15395
rect 20125 15365 20155 15395
rect 20205 15365 20235 15395
rect 20285 15365 20315 15395
rect 20365 15365 20395 15395
rect 20445 15365 20475 15395
rect 20525 15365 20555 15395
rect 20605 15365 20635 15395
rect 20685 15365 20715 15395
rect 20765 15365 20795 15395
rect 20845 15365 20875 15395
rect 20925 15365 20955 15395
rect 5605 15285 5635 15315
rect 10885 15285 10915 15315
rect 15325 15285 15355 15315
rect 5 15205 35 15235
rect 85 15205 115 15235
rect 165 15205 195 15235
rect 245 15205 275 15235
rect 325 15205 355 15235
rect 405 15205 435 15235
rect 485 15205 515 15235
rect 565 15205 595 15235
rect 645 15205 675 15235
rect 725 15205 755 15235
rect 805 15205 835 15235
rect 885 15205 915 15235
rect 965 15205 995 15235
rect 1045 15205 1075 15235
rect 1125 15205 1155 15235
rect 1205 15205 1235 15235
rect 1285 15205 1315 15235
rect 1365 15205 1395 15235
rect 1445 15205 1475 15235
rect 1525 15205 1555 15235
rect 1605 15205 1635 15235
rect 1685 15205 1715 15235
rect 1765 15205 1795 15235
rect 1845 15205 1875 15235
rect 1925 15205 1955 15235
rect 2005 15205 2035 15235
rect 2085 15205 2115 15235
rect 2165 15205 2195 15235
rect 2245 15205 2275 15235
rect 2325 15205 2355 15235
rect 2405 15205 2435 15235
rect 2485 15205 2515 15235
rect 2565 15205 2595 15235
rect 2645 15205 2675 15235
rect 2725 15205 2755 15235
rect 2805 15205 2835 15235
rect 2885 15205 2915 15235
rect 2965 15205 2995 15235
rect 3045 15205 3075 15235
rect 3125 15205 3155 15235
rect 3205 15205 3235 15235
rect 3285 15205 3315 15235
rect 3365 15205 3395 15235
rect 3445 15205 3475 15235
rect 3525 15205 3555 15235
rect 3605 15205 3635 15235
rect 3685 15205 3715 15235
rect 3765 15205 3795 15235
rect 3845 15205 3875 15235
rect 3925 15205 3955 15235
rect 4005 15205 4035 15235
rect 4085 15205 4115 15235
rect 4165 15205 4195 15235
rect 4725 15205 4755 15235
rect 4885 15205 4915 15235
rect 5045 15205 5075 15235
rect 5205 15205 5235 15235
rect 5365 15205 5395 15235
rect 5525 15205 5555 15235
rect 5685 15205 5715 15235
rect 6245 15205 6275 15235
rect 6325 15205 6355 15235
rect 6405 15205 6435 15235
rect 6485 15205 6515 15235
rect 6565 15205 6595 15235
rect 6645 15205 6675 15235
rect 6725 15205 6755 15235
rect 6805 15205 6835 15235
rect 6885 15205 6915 15235
rect 6965 15205 6995 15235
rect 7045 15205 7075 15235
rect 7125 15205 7155 15235
rect 7205 15205 7235 15235
rect 7285 15205 7315 15235
rect 7365 15205 7395 15235
rect 7445 15205 7475 15235
rect 7525 15205 7555 15235
rect 7605 15205 7635 15235
rect 7685 15205 7715 15235
rect 7765 15205 7795 15235
rect 7845 15205 7875 15235
rect 7925 15205 7955 15235
rect 8005 15205 8035 15235
rect 8085 15205 8115 15235
rect 8165 15205 8195 15235
rect 8245 15205 8275 15235
rect 8325 15205 8355 15235
rect 8405 15205 8435 15235
rect 8485 15205 8515 15235
rect 8565 15205 8595 15235
rect 8645 15205 8675 15235
rect 8725 15205 8755 15235
rect 8805 15205 8835 15235
rect 8885 15205 8915 15235
rect 8965 15205 8995 15235
rect 9045 15205 9075 15235
rect 9125 15205 9155 15235
rect 9205 15205 9235 15235
rect 9285 15205 9315 15235
rect 9365 15205 9395 15235
rect 9445 15205 9475 15235
rect 10005 15205 10035 15235
rect 10165 15205 10195 15235
rect 10325 15205 10355 15235
rect 10485 15205 10515 15235
rect 10645 15205 10675 15235
rect 10805 15205 10835 15235
rect 10965 15205 10995 15235
rect 11565 15205 11595 15235
rect 11645 15205 11675 15235
rect 11725 15205 11755 15235
rect 11805 15205 11835 15235
rect 11885 15205 11915 15235
rect 11965 15205 11995 15235
rect 12045 15205 12075 15235
rect 12125 15205 12155 15235
rect 12205 15205 12235 15235
rect 12285 15205 12315 15235
rect 12365 15205 12395 15235
rect 12445 15205 12475 15235
rect 12525 15205 12555 15235
rect 12605 15205 12635 15235
rect 12685 15205 12715 15235
rect 12765 15205 12795 15235
rect 12845 15205 12875 15235
rect 12925 15205 12955 15235
rect 13005 15205 13035 15235
rect 13085 15205 13115 15235
rect 13165 15205 13195 15235
rect 13245 15205 13275 15235
rect 13325 15205 13355 15235
rect 13405 15205 13435 15235
rect 13485 15205 13515 15235
rect 13565 15205 13595 15235
rect 13645 15205 13675 15235
rect 13725 15205 13755 15235
rect 13805 15205 13835 15235
rect 13885 15205 13915 15235
rect 13965 15205 13995 15235
rect 14045 15205 14075 15235
rect 14125 15205 14155 15235
rect 14205 15205 14235 15235
rect 14285 15205 14315 15235
rect 14365 15205 14395 15235
rect 14445 15205 14475 15235
rect 14525 15205 14555 15235
rect 14605 15205 14635 15235
rect 14685 15205 14715 15235
rect 15245 15205 15275 15235
rect 15405 15205 15435 15235
rect 15565 15205 15595 15235
rect 15725 15205 15755 15235
rect 15885 15205 15915 15235
rect 16045 15205 16075 15235
rect 16205 15205 16235 15235
rect 16765 15205 16795 15235
rect 16845 15205 16875 15235
rect 16925 15205 16955 15235
rect 17005 15205 17035 15235
rect 17085 15205 17115 15235
rect 17165 15205 17195 15235
rect 17245 15205 17275 15235
rect 17325 15205 17355 15235
rect 17405 15205 17435 15235
rect 17485 15205 17515 15235
rect 17565 15205 17595 15235
rect 17645 15205 17675 15235
rect 17725 15205 17755 15235
rect 17805 15205 17835 15235
rect 17885 15205 17915 15235
rect 17965 15205 17995 15235
rect 18045 15205 18075 15235
rect 18125 15205 18155 15235
rect 18205 15205 18235 15235
rect 18285 15205 18315 15235
rect 18365 15205 18395 15235
rect 18445 15205 18475 15235
rect 18525 15205 18555 15235
rect 18605 15205 18635 15235
rect 18685 15205 18715 15235
rect 18765 15205 18795 15235
rect 18845 15205 18875 15235
rect 18925 15205 18955 15235
rect 19005 15205 19035 15235
rect 19085 15205 19115 15235
rect 19165 15205 19195 15235
rect 19245 15205 19275 15235
rect 19325 15205 19355 15235
rect 19405 15205 19435 15235
rect 19485 15205 19515 15235
rect 19565 15205 19595 15235
rect 19645 15205 19675 15235
rect 19725 15205 19755 15235
rect 19805 15205 19835 15235
rect 19885 15205 19915 15235
rect 19965 15205 19995 15235
rect 20045 15205 20075 15235
rect 20125 15205 20155 15235
rect 20205 15205 20235 15235
rect 20285 15205 20315 15235
rect 20365 15205 20395 15235
rect 20445 15205 20475 15235
rect 20525 15205 20555 15235
rect 20605 15205 20635 15235
rect 20685 15205 20715 15235
rect 20765 15205 20795 15235
rect 20845 15205 20875 15235
rect 20925 15205 20955 15235
rect 5 15125 35 15155
rect 85 15125 115 15155
rect 165 15125 195 15155
rect 245 15125 275 15155
rect 325 15125 355 15155
rect 405 15125 435 15155
rect 485 15125 515 15155
rect 565 15125 595 15155
rect 645 15125 675 15155
rect 725 15125 755 15155
rect 805 15125 835 15155
rect 885 15125 915 15155
rect 965 15125 995 15155
rect 1045 15125 1075 15155
rect 1125 15125 1155 15155
rect 1205 15125 1235 15155
rect 1285 15125 1315 15155
rect 1365 15125 1395 15155
rect 1445 15125 1475 15155
rect 1525 15125 1555 15155
rect 1605 15125 1635 15155
rect 1685 15125 1715 15155
rect 1765 15125 1795 15155
rect 1845 15125 1875 15155
rect 1925 15125 1955 15155
rect 2005 15125 2035 15155
rect 2085 15125 2115 15155
rect 2165 15125 2195 15155
rect 2245 15125 2275 15155
rect 2325 15125 2355 15155
rect 2405 15125 2435 15155
rect 2485 15125 2515 15155
rect 2565 15125 2595 15155
rect 2645 15125 2675 15155
rect 2725 15125 2755 15155
rect 2805 15125 2835 15155
rect 2885 15125 2915 15155
rect 2965 15125 2995 15155
rect 3045 15125 3075 15155
rect 3125 15125 3155 15155
rect 3205 15125 3235 15155
rect 3285 15125 3315 15155
rect 3365 15125 3395 15155
rect 3445 15125 3475 15155
rect 3525 15125 3555 15155
rect 3605 15125 3635 15155
rect 3685 15125 3715 15155
rect 3765 15125 3795 15155
rect 3845 15125 3875 15155
rect 3925 15125 3955 15155
rect 4005 15125 4035 15155
rect 4085 15125 4115 15155
rect 4165 15125 4195 15155
rect 5765 15125 5795 15155
rect 5925 15125 5955 15155
rect 6245 15125 6275 15155
rect 6325 15125 6355 15155
rect 6405 15125 6435 15155
rect 6485 15125 6515 15155
rect 6565 15125 6595 15155
rect 6645 15125 6675 15155
rect 6725 15125 6755 15155
rect 6805 15125 6835 15155
rect 6885 15125 6915 15155
rect 6965 15125 6995 15155
rect 7045 15125 7075 15155
rect 7125 15125 7155 15155
rect 7205 15125 7235 15155
rect 7285 15125 7315 15155
rect 7365 15125 7395 15155
rect 7445 15125 7475 15155
rect 7525 15125 7555 15155
rect 7605 15125 7635 15155
rect 7685 15125 7715 15155
rect 7765 15125 7795 15155
rect 7845 15125 7875 15155
rect 7925 15125 7955 15155
rect 8005 15125 8035 15155
rect 8085 15125 8115 15155
rect 8165 15125 8195 15155
rect 8245 15125 8275 15155
rect 8325 15125 8355 15155
rect 8405 15125 8435 15155
rect 8485 15125 8515 15155
rect 8565 15125 8595 15155
rect 8645 15125 8675 15155
rect 8725 15125 8755 15155
rect 8805 15125 8835 15155
rect 8885 15125 8915 15155
rect 8965 15125 8995 15155
rect 9045 15125 9075 15155
rect 9125 15125 9155 15155
rect 9205 15125 9235 15155
rect 9285 15125 9315 15155
rect 9365 15125 9395 15155
rect 9445 15125 9475 15155
rect 11045 15125 11075 15155
rect 11205 15125 11235 15155
rect 11565 15125 11595 15155
rect 11645 15125 11675 15155
rect 11725 15125 11755 15155
rect 11805 15125 11835 15155
rect 11885 15125 11915 15155
rect 11965 15125 11995 15155
rect 12045 15125 12075 15155
rect 12125 15125 12155 15155
rect 12205 15125 12235 15155
rect 12285 15125 12315 15155
rect 12365 15125 12395 15155
rect 12445 15125 12475 15155
rect 12525 15125 12555 15155
rect 12605 15125 12635 15155
rect 12685 15125 12715 15155
rect 12765 15125 12795 15155
rect 12845 15125 12875 15155
rect 12925 15125 12955 15155
rect 13005 15125 13035 15155
rect 13085 15125 13115 15155
rect 13165 15125 13195 15155
rect 13245 15125 13275 15155
rect 13325 15125 13355 15155
rect 13405 15125 13435 15155
rect 13485 15125 13515 15155
rect 13565 15125 13595 15155
rect 13645 15125 13675 15155
rect 13725 15125 13755 15155
rect 13805 15125 13835 15155
rect 13885 15125 13915 15155
rect 13965 15125 13995 15155
rect 14045 15125 14075 15155
rect 14125 15125 14155 15155
rect 14205 15125 14235 15155
rect 14285 15125 14315 15155
rect 14365 15125 14395 15155
rect 14445 15125 14475 15155
rect 14525 15125 14555 15155
rect 14605 15125 14635 15155
rect 14685 15125 14715 15155
rect 15005 15125 15035 15155
rect 15165 15125 15195 15155
rect 16765 15125 16795 15155
rect 16845 15125 16875 15155
rect 16925 15125 16955 15155
rect 17005 15125 17035 15155
rect 17085 15125 17115 15155
rect 17165 15125 17195 15155
rect 17245 15125 17275 15155
rect 17325 15125 17355 15155
rect 17405 15125 17435 15155
rect 17485 15125 17515 15155
rect 17565 15125 17595 15155
rect 17645 15125 17675 15155
rect 17725 15125 17755 15155
rect 17805 15125 17835 15155
rect 17885 15125 17915 15155
rect 17965 15125 17995 15155
rect 18045 15125 18075 15155
rect 18125 15125 18155 15155
rect 18205 15125 18235 15155
rect 18285 15125 18315 15155
rect 18365 15125 18395 15155
rect 18445 15125 18475 15155
rect 18525 15125 18555 15155
rect 18605 15125 18635 15155
rect 18685 15125 18715 15155
rect 18765 15125 18795 15155
rect 18845 15125 18875 15155
rect 18925 15125 18955 15155
rect 19005 15125 19035 15155
rect 19085 15125 19115 15155
rect 19165 15125 19195 15155
rect 19245 15125 19275 15155
rect 19325 15125 19355 15155
rect 19405 15125 19435 15155
rect 19485 15125 19515 15155
rect 19565 15125 19595 15155
rect 19645 15125 19675 15155
rect 19725 15125 19755 15155
rect 19805 15125 19835 15155
rect 19885 15125 19915 15155
rect 19965 15125 19995 15155
rect 20045 15125 20075 15155
rect 20125 15125 20155 15155
rect 20205 15125 20235 15155
rect 20285 15125 20315 15155
rect 20365 15125 20395 15155
rect 20445 15125 20475 15155
rect 20525 15125 20555 15155
rect 20605 15125 20635 15155
rect 20685 15125 20715 15155
rect 20765 15125 20795 15155
rect 20845 15125 20875 15155
rect 20925 15125 20955 15155
rect 5845 15045 5875 15075
rect 11125 15045 11155 15075
rect 15085 15045 15115 15075
rect 5 14965 35 14995
rect 85 14965 115 14995
rect 165 14965 195 14995
rect 245 14965 275 14995
rect 325 14965 355 14995
rect 405 14965 435 14995
rect 485 14965 515 14995
rect 565 14965 595 14995
rect 645 14965 675 14995
rect 725 14965 755 14995
rect 805 14965 835 14995
rect 885 14965 915 14995
rect 965 14965 995 14995
rect 1045 14965 1075 14995
rect 1125 14965 1155 14995
rect 1205 14965 1235 14995
rect 1285 14965 1315 14995
rect 1365 14965 1395 14995
rect 1445 14965 1475 14995
rect 1525 14965 1555 14995
rect 1605 14965 1635 14995
rect 1685 14965 1715 14995
rect 1765 14965 1795 14995
rect 1845 14965 1875 14995
rect 1925 14965 1955 14995
rect 2005 14965 2035 14995
rect 2085 14965 2115 14995
rect 2165 14965 2195 14995
rect 2245 14965 2275 14995
rect 2325 14965 2355 14995
rect 2405 14965 2435 14995
rect 2485 14965 2515 14995
rect 2565 14965 2595 14995
rect 2645 14965 2675 14995
rect 2725 14965 2755 14995
rect 2805 14965 2835 14995
rect 2885 14965 2915 14995
rect 2965 14965 2995 14995
rect 3045 14965 3075 14995
rect 3125 14965 3155 14995
rect 3205 14965 3235 14995
rect 3285 14965 3315 14995
rect 3365 14965 3395 14995
rect 3445 14965 3475 14995
rect 3525 14965 3555 14995
rect 3605 14965 3635 14995
rect 3685 14965 3715 14995
rect 3765 14965 3795 14995
rect 3845 14965 3875 14995
rect 3925 14965 3955 14995
rect 4005 14965 4035 14995
rect 4085 14965 4115 14995
rect 4165 14965 4195 14995
rect 5765 14965 5795 14995
rect 5925 14965 5955 14995
rect 6245 14965 6275 14995
rect 6325 14965 6355 14995
rect 6405 14965 6435 14995
rect 6485 14965 6515 14995
rect 6565 14965 6595 14995
rect 6645 14965 6675 14995
rect 6725 14965 6755 14995
rect 6805 14965 6835 14995
rect 6885 14965 6915 14995
rect 6965 14965 6995 14995
rect 7045 14965 7075 14995
rect 7125 14965 7155 14995
rect 7205 14965 7235 14995
rect 7285 14965 7315 14995
rect 7365 14965 7395 14995
rect 7445 14965 7475 14995
rect 7525 14965 7555 14995
rect 7605 14965 7635 14995
rect 7685 14965 7715 14995
rect 7765 14965 7795 14995
rect 7845 14965 7875 14995
rect 7925 14965 7955 14995
rect 8005 14965 8035 14995
rect 8085 14965 8115 14995
rect 8165 14965 8195 14995
rect 8245 14965 8275 14995
rect 8325 14965 8355 14995
rect 8405 14965 8435 14995
rect 8485 14965 8515 14995
rect 8565 14965 8595 14995
rect 8645 14965 8675 14995
rect 8725 14965 8755 14995
rect 8805 14965 8835 14995
rect 8885 14965 8915 14995
rect 8965 14965 8995 14995
rect 9045 14965 9075 14995
rect 9125 14965 9155 14995
rect 9205 14965 9235 14995
rect 9285 14965 9315 14995
rect 9365 14965 9395 14995
rect 9445 14965 9475 14995
rect 11045 14965 11075 14995
rect 11205 14965 11235 14995
rect 11565 14965 11595 14995
rect 11645 14965 11675 14995
rect 11725 14965 11755 14995
rect 11805 14965 11835 14995
rect 11885 14965 11915 14995
rect 11965 14965 11995 14995
rect 12045 14965 12075 14995
rect 12125 14965 12155 14995
rect 12205 14965 12235 14995
rect 12285 14965 12315 14995
rect 12365 14965 12395 14995
rect 12445 14965 12475 14995
rect 12525 14965 12555 14995
rect 12605 14965 12635 14995
rect 12685 14965 12715 14995
rect 12765 14965 12795 14995
rect 12845 14965 12875 14995
rect 12925 14965 12955 14995
rect 13005 14965 13035 14995
rect 13085 14965 13115 14995
rect 13165 14965 13195 14995
rect 13245 14965 13275 14995
rect 13325 14965 13355 14995
rect 13405 14965 13435 14995
rect 13485 14965 13515 14995
rect 13565 14965 13595 14995
rect 13645 14965 13675 14995
rect 13725 14965 13755 14995
rect 13805 14965 13835 14995
rect 13885 14965 13915 14995
rect 13965 14965 13995 14995
rect 14045 14965 14075 14995
rect 14125 14965 14155 14995
rect 14205 14965 14235 14995
rect 14285 14965 14315 14995
rect 14365 14965 14395 14995
rect 14445 14965 14475 14995
rect 14525 14965 14555 14995
rect 14605 14965 14635 14995
rect 14685 14965 14715 14995
rect 15005 14965 15035 14995
rect 15165 14965 15195 14995
rect 16765 14965 16795 14995
rect 16845 14965 16875 14995
rect 16925 14965 16955 14995
rect 17005 14965 17035 14995
rect 17085 14965 17115 14995
rect 17165 14965 17195 14995
rect 17245 14965 17275 14995
rect 17325 14965 17355 14995
rect 17405 14965 17435 14995
rect 17485 14965 17515 14995
rect 17565 14965 17595 14995
rect 17645 14965 17675 14995
rect 17725 14965 17755 14995
rect 17805 14965 17835 14995
rect 17885 14965 17915 14995
rect 17965 14965 17995 14995
rect 18045 14965 18075 14995
rect 18125 14965 18155 14995
rect 18205 14965 18235 14995
rect 18285 14965 18315 14995
rect 18365 14965 18395 14995
rect 18445 14965 18475 14995
rect 18525 14965 18555 14995
rect 18605 14965 18635 14995
rect 18685 14965 18715 14995
rect 18765 14965 18795 14995
rect 18845 14965 18875 14995
rect 18925 14965 18955 14995
rect 19005 14965 19035 14995
rect 19085 14965 19115 14995
rect 19165 14965 19195 14995
rect 19245 14965 19275 14995
rect 19325 14965 19355 14995
rect 19405 14965 19435 14995
rect 19485 14965 19515 14995
rect 19565 14965 19595 14995
rect 19645 14965 19675 14995
rect 19725 14965 19755 14995
rect 19805 14965 19835 14995
rect 19885 14965 19915 14995
rect 19965 14965 19995 14995
rect 20045 14965 20075 14995
rect 20125 14965 20155 14995
rect 20205 14965 20235 14995
rect 20285 14965 20315 14995
rect 20365 14965 20395 14995
rect 20445 14965 20475 14995
rect 20525 14965 20555 14995
rect 20605 14965 20635 14995
rect 20685 14965 20715 14995
rect 20765 14965 20795 14995
rect 20845 14965 20875 14995
rect 20925 14965 20955 14995
rect 5 14885 35 14915
rect 85 14885 115 14915
rect 165 14885 195 14915
rect 245 14885 275 14915
rect 325 14885 355 14915
rect 405 14885 435 14915
rect 485 14885 515 14915
rect 565 14885 595 14915
rect 645 14885 675 14915
rect 725 14885 755 14915
rect 805 14885 835 14915
rect 885 14885 915 14915
rect 965 14885 995 14915
rect 1045 14885 1075 14915
rect 1125 14885 1155 14915
rect 1205 14885 1235 14915
rect 1285 14885 1315 14915
rect 1365 14885 1395 14915
rect 1445 14885 1475 14915
rect 1525 14885 1555 14915
rect 1605 14885 1635 14915
rect 1685 14885 1715 14915
rect 1765 14885 1795 14915
rect 1845 14885 1875 14915
rect 1925 14885 1955 14915
rect 2005 14885 2035 14915
rect 2085 14885 2115 14915
rect 2165 14885 2195 14915
rect 2245 14885 2275 14915
rect 2325 14885 2355 14915
rect 2405 14885 2435 14915
rect 2485 14885 2515 14915
rect 2565 14885 2595 14915
rect 2645 14885 2675 14915
rect 2725 14885 2755 14915
rect 2805 14885 2835 14915
rect 2885 14885 2915 14915
rect 2965 14885 2995 14915
rect 3045 14885 3075 14915
rect 3125 14885 3155 14915
rect 3205 14885 3235 14915
rect 3285 14885 3315 14915
rect 3365 14885 3395 14915
rect 3445 14885 3475 14915
rect 3525 14885 3555 14915
rect 3605 14885 3635 14915
rect 3685 14885 3715 14915
rect 3765 14885 3795 14915
rect 3845 14885 3875 14915
rect 3925 14885 3955 14915
rect 4005 14885 4035 14915
rect 4085 14885 4115 14915
rect 4165 14885 4195 14915
rect 6005 14885 6035 14915
rect 6165 14885 6195 14915
rect 6245 14885 6275 14915
rect 6325 14885 6355 14915
rect 6405 14885 6435 14915
rect 6485 14885 6515 14915
rect 6565 14885 6595 14915
rect 6645 14885 6675 14915
rect 6725 14885 6755 14915
rect 6805 14885 6835 14915
rect 6885 14885 6915 14915
rect 6965 14885 6995 14915
rect 7045 14885 7075 14915
rect 7125 14885 7155 14915
rect 7205 14885 7235 14915
rect 7285 14885 7315 14915
rect 7365 14885 7395 14915
rect 7445 14885 7475 14915
rect 7525 14885 7555 14915
rect 7605 14885 7635 14915
rect 7685 14885 7715 14915
rect 7765 14885 7795 14915
rect 7845 14885 7875 14915
rect 7925 14885 7955 14915
rect 8005 14885 8035 14915
rect 8085 14885 8115 14915
rect 8165 14885 8195 14915
rect 8245 14885 8275 14915
rect 8325 14885 8355 14915
rect 8405 14885 8435 14915
rect 8485 14885 8515 14915
rect 8565 14885 8595 14915
rect 8645 14885 8675 14915
rect 8725 14885 8755 14915
rect 8805 14885 8835 14915
rect 8885 14885 8915 14915
rect 8965 14885 8995 14915
rect 9045 14885 9075 14915
rect 9125 14885 9155 14915
rect 9205 14885 9235 14915
rect 9285 14885 9315 14915
rect 9365 14885 9395 14915
rect 9445 14885 9475 14915
rect 11285 14885 11315 14915
rect 11445 14885 11475 14915
rect 11565 14885 11595 14915
rect 11645 14885 11675 14915
rect 11725 14885 11755 14915
rect 11805 14885 11835 14915
rect 11885 14885 11915 14915
rect 11965 14885 11995 14915
rect 12045 14885 12075 14915
rect 12125 14885 12155 14915
rect 12205 14885 12235 14915
rect 12285 14885 12315 14915
rect 12365 14885 12395 14915
rect 12445 14885 12475 14915
rect 12525 14885 12555 14915
rect 12605 14885 12635 14915
rect 12685 14885 12715 14915
rect 12765 14885 12795 14915
rect 12845 14885 12875 14915
rect 12925 14885 12955 14915
rect 13005 14885 13035 14915
rect 13085 14885 13115 14915
rect 13165 14885 13195 14915
rect 13245 14885 13275 14915
rect 13325 14885 13355 14915
rect 13405 14885 13435 14915
rect 13485 14885 13515 14915
rect 13565 14885 13595 14915
rect 13645 14885 13675 14915
rect 13725 14885 13755 14915
rect 13805 14885 13835 14915
rect 13885 14885 13915 14915
rect 13965 14885 13995 14915
rect 14045 14885 14075 14915
rect 14125 14885 14155 14915
rect 14205 14885 14235 14915
rect 14285 14885 14315 14915
rect 14365 14885 14395 14915
rect 14445 14885 14475 14915
rect 14525 14885 14555 14915
rect 14605 14885 14635 14915
rect 14685 14885 14715 14915
rect 14765 14885 14795 14915
rect 14925 14885 14955 14915
rect 16765 14885 16795 14915
rect 16845 14885 16875 14915
rect 16925 14885 16955 14915
rect 17005 14885 17035 14915
rect 17085 14885 17115 14915
rect 17165 14885 17195 14915
rect 17245 14885 17275 14915
rect 17325 14885 17355 14915
rect 17405 14885 17435 14915
rect 17485 14885 17515 14915
rect 17565 14885 17595 14915
rect 17645 14885 17675 14915
rect 17725 14885 17755 14915
rect 17805 14885 17835 14915
rect 17885 14885 17915 14915
rect 17965 14885 17995 14915
rect 18045 14885 18075 14915
rect 18125 14885 18155 14915
rect 18205 14885 18235 14915
rect 18285 14885 18315 14915
rect 18365 14885 18395 14915
rect 18445 14885 18475 14915
rect 18525 14885 18555 14915
rect 18605 14885 18635 14915
rect 18685 14885 18715 14915
rect 18765 14885 18795 14915
rect 18845 14885 18875 14915
rect 18925 14885 18955 14915
rect 19005 14885 19035 14915
rect 19085 14885 19115 14915
rect 19165 14885 19195 14915
rect 19245 14885 19275 14915
rect 19325 14885 19355 14915
rect 19405 14885 19435 14915
rect 19485 14885 19515 14915
rect 19565 14885 19595 14915
rect 19645 14885 19675 14915
rect 19725 14885 19755 14915
rect 19805 14885 19835 14915
rect 19885 14885 19915 14915
rect 19965 14885 19995 14915
rect 20045 14885 20075 14915
rect 20125 14885 20155 14915
rect 20205 14885 20235 14915
rect 20285 14885 20315 14915
rect 20365 14885 20395 14915
rect 20445 14885 20475 14915
rect 20525 14885 20555 14915
rect 20605 14885 20635 14915
rect 20685 14885 20715 14915
rect 20765 14885 20795 14915
rect 20845 14885 20875 14915
rect 20925 14885 20955 14915
rect 6085 14805 6115 14835
rect 11365 14805 11395 14835
rect 14845 14805 14875 14835
rect 5 14725 35 14755
rect 85 14725 115 14755
rect 165 14725 195 14755
rect 245 14725 275 14755
rect 325 14725 355 14755
rect 405 14725 435 14755
rect 485 14725 515 14755
rect 565 14725 595 14755
rect 645 14725 675 14755
rect 725 14725 755 14755
rect 805 14725 835 14755
rect 885 14725 915 14755
rect 965 14725 995 14755
rect 1045 14725 1075 14755
rect 1125 14725 1155 14755
rect 1205 14725 1235 14755
rect 1285 14725 1315 14755
rect 1365 14725 1395 14755
rect 1445 14725 1475 14755
rect 1525 14725 1555 14755
rect 1605 14725 1635 14755
rect 1685 14725 1715 14755
rect 1765 14725 1795 14755
rect 1845 14725 1875 14755
rect 1925 14725 1955 14755
rect 2005 14725 2035 14755
rect 2085 14725 2115 14755
rect 2165 14725 2195 14755
rect 2245 14725 2275 14755
rect 2325 14725 2355 14755
rect 2405 14725 2435 14755
rect 2485 14725 2515 14755
rect 2565 14725 2595 14755
rect 2645 14725 2675 14755
rect 2725 14725 2755 14755
rect 2805 14725 2835 14755
rect 2885 14725 2915 14755
rect 2965 14725 2995 14755
rect 3045 14725 3075 14755
rect 3125 14725 3155 14755
rect 3205 14725 3235 14755
rect 3285 14725 3315 14755
rect 3365 14725 3395 14755
rect 3445 14725 3475 14755
rect 3525 14725 3555 14755
rect 3605 14725 3635 14755
rect 3685 14725 3715 14755
rect 3765 14725 3795 14755
rect 3845 14725 3875 14755
rect 3925 14725 3955 14755
rect 4005 14725 4035 14755
rect 4085 14725 4115 14755
rect 4165 14725 4195 14755
rect 6005 14725 6035 14755
rect 6165 14725 6195 14755
rect 6245 14725 6275 14755
rect 6325 14725 6355 14755
rect 6405 14725 6435 14755
rect 6485 14725 6515 14755
rect 6565 14725 6595 14755
rect 6645 14725 6675 14755
rect 6725 14725 6755 14755
rect 6805 14725 6835 14755
rect 6885 14725 6915 14755
rect 6965 14725 6995 14755
rect 7045 14725 7075 14755
rect 7125 14725 7155 14755
rect 7205 14725 7235 14755
rect 7285 14725 7315 14755
rect 7365 14725 7395 14755
rect 7445 14725 7475 14755
rect 7525 14725 7555 14755
rect 7605 14725 7635 14755
rect 7685 14725 7715 14755
rect 7765 14725 7795 14755
rect 7845 14725 7875 14755
rect 7925 14725 7955 14755
rect 8005 14725 8035 14755
rect 8085 14725 8115 14755
rect 8165 14725 8195 14755
rect 8245 14725 8275 14755
rect 8325 14725 8355 14755
rect 8405 14725 8435 14755
rect 8485 14725 8515 14755
rect 8565 14725 8595 14755
rect 8645 14725 8675 14755
rect 8725 14725 8755 14755
rect 8805 14725 8835 14755
rect 8885 14725 8915 14755
rect 8965 14725 8995 14755
rect 9045 14725 9075 14755
rect 9125 14725 9155 14755
rect 9205 14725 9235 14755
rect 9285 14725 9315 14755
rect 9365 14725 9395 14755
rect 9445 14725 9475 14755
rect 11285 14725 11315 14755
rect 11445 14725 11475 14755
rect 11565 14725 11595 14755
rect 11645 14725 11675 14755
rect 11725 14725 11755 14755
rect 11805 14725 11835 14755
rect 11885 14725 11915 14755
rect 11965 14725 11995 14755
rect 12045 14725 12075 14755
rect 12125 14725 12155 14755
rect 12205 14725 12235 14755
rect 12285 14725 12315 14755
rect 12365 14725 12395 14755
rect 12445 14725 12475 14755
rect 12525 14725 12555 14755
rect 12605 14725 12635 14755
rect 12685 14725 12715 14755
rect 12765 14725 12795 14755
rect 12845 14725 12875 14755
rect 12925 14725 12955 14755
rect 13005 14725 13035 14755
rect 13085 14725 13115 14755
rect 13165 14725 13195 14755
rect 13245 14725 13275 14755
rect 13325 14725 13355 14755
rect 13405 14725 13435 14755
rect 13485 14725 13515 14755
rect 13565 14725 13595 14755
rect 13645 14725 13675 14755
rect 13725 14725 13755 14755
rect 13805 14725 13835 14755
rect 13885 14725 13915 14755
rect 13965 14725 13995 14755
rect 14045 14725 14075 14755
rect 14125 14725 14155 14755
rect 14205 14725 14235 14755
rect 14285 14725 14315 14755
rect 14365 14725 14395 14755
rect 14445 14725 14475 14755
rect 14525 14725 14555 14755
rect 14605 14725 14635 14755
rect 14685 14725 14715 14755
rect 14765 14725 14795 14755
rect 14925 14725 14955 14755
rect 16765 14725 16795 14755
rect 16845 14725 16875 14755
rect 16925 14725 16955 14755
rect 17005 14725 17035 14755
rect 17085 14725 17115 14755
rect 17165 14725 17195 14755
rect 17245 14725 17275 14755
rect 17325 14725 17355 14755
rect 17405 14725 17435 14755
rect 17485 14725 17515 14755
rect 17565 14725 17595 14755
rect 17645 14725 17675 14755
rect 17725 14725 17755 14755
rect 17805 14725 17835 14755
rect 17885 14725 17915 14755
rect 17965 14725 17995 14755
rect 18045 14725 18075 14755
rect 18125 14725 18155 14755
rect 18205 14725 18235 14755
rect 18285 14725 18315 14755
rect 18365 14725 18395 14755
rect 18445 14725 18475 14755
rect 18525 14725 18555 14755
rect 18605 14725 18635 14755
rect 18685 14725 18715 14755
rect 18765 14725 18795 14755
rect 18845 14725 18875 14755
rect 18925 14725 18955 14755
rect 19005 14725 19035 14755
rect 19085 14725 19115 14755
rect 19165 14725 19195 14755
rect 19245 14725 19275 14755
rect 19325 14725 19355 14755
rect 19405 14725 19435 14755
rect 19485 14725 19515 14755
rect 19565 14725 19595 14755
rect 19645 14725 19675 14755
rect 19725 14725 19755 14755
rect 19805 14725 19835 14755
rect 19885 14725 19915 14755
rect 19965 14725 19995 14755
rect 20045 14725 20075 14755
rect 20125 14725 20155 14755
rect 20205 14725 20235 14755
rect 20285 14725 20315 14755
rect 20365 14725 20395 14755
rect 20445 14725 20475 14755
rect 20525 14725 20555 14755
rect 20605 14725 20635 14755
rect 20685 14725 20715 14755
rect 20765 14725 20795 14755
rect 20845 14725 20875 14755
rect 20925 14725 20955 14755
<< metal3 >>
rect 0 18675 40 18680
rect 0 18645 5 18675
rect 35 18645 40 18675
rect 0 18515 40 18645
rect 0 18485 5 18515
rect 35 18485 40 18515
rect 0 18480 40 18485
rect 80 18675 120 18680
rect 80 18645 85 18675
rect 115 18645 120 18675
rect 80 18515 120 18645
rect 80 18485 85 18515
rect 115 18485 120 18515
rect 80 18480 120 18485
rect 160 18675 200 18680
rect 160 18645 165 18675
rect 195 18645 200 18675
rect 160 18515 200 18645
rect 160 18485 165 18515
rect 195 18485 200 18515
rect 160 18480 200 18485
rect 240 18675 280 18680
rect 240 18645 245 18675
rect 275 18645 280 18675
rect 240 18515 280 18645
rect 240 18485 245 18515
rect 275 18485 280 18515
rect 240 18480 280 18485
rect 320 18675 360 18680
rect 320 18645 325 18675
rect 355 18645 360 18675
rect 320 18515 360 18645
rect 320 18485 325 18515
rect 355 18485 360 18515
rect 320 18480 360 18485
rect 400 18675 440 18680
rect 400 18645 405 18675
rect 435 18645 440 18675
rect 400 18515 440 18645
rect 400 18485 405 18515
rect 435 18485 440 18515
rect 400 18480 440 18485
rect 480 18675 520 18680
rect 480 18645 485 18675
rect 515 18645 520 18675
rect 480 18515 520 18645
rect 480 18485 485 18515
rect 515 18485 520 18515
rect 480 18480 520 18485
rect 560 18675 600 18680
rect 560 18645 565 18675
rect 595 18645 600 18675
rect 560 18515 600 18645
rect 560 18485 565 18515
rect 595 18485 600 18515
rect 560 18480 600 18485
rect 640 18675 680 18680
rect 640 18645 645 18675
rect 675 18645 680 18675
rect 640 18515 680 18645
rect 640 18485 645 18515
rect 675 18485 680 18515
rect 640 18480 680 18485
rect 720 18675 760 18680
rect 720 18645 725 18675
rect 755 18645 760 18675
rect 720 18515 760 18645
rect 720 18485 725 18515
rect 755 18485 760 18515
rect 720 18480 760 18485
rect 800 18675 840 18680
rect 800 18645 805 18675
rect 835 18645 840 18675
rect 800 18515 840 18645
rect 800 18485 805 18515
rect 835 18485 840 18515
rect 800 18480 840 18485
rect 880 18675 920 18680
rect 880 18645 885 18675
rect 915 18645 920 18675
rect 880 18515 920 18645
rect 880 18485 885 18515
rect 915 18485 920 18515
rect 880 18480 920 18485
rect 960 18675 1000 18680
rect 960 18645 965 18675
rect 995 18645 1000 18675
rect 960 18515 1000 18645
rect 960 18485 965 18515
rect 995 18485 1000 18515
rect 960 18480 1000 18485
rect 1040 18675 1080 18680
rect 1040 18645 1045 18675
rect 1075 18645 1080 18675
rect 1040 18515 1080 18645
rect 1040 18485 1045 18515
rect 1075 18485 1080 18515
rect 1040 18480 1080 18485
rect 1120 18675 1160 18680
rect 1120 18645 1125 18675
rect 1155 18645 1160 18675
rect 1120 18515 1160 18645
rect 1120 18485 1125 18515
rect 1155 18485 1160 18515
rect 1120 18480 1160 18485
rect 1200 18675 1240 18680
rect 1200 18645 1205 18675
rect 1235 18645 1240 18675
rect 1200 18515 1240 18645
rect 1200 18485 1205 18515
rect 1235 18485 1240 18515
rect 1200 18480 1240 18485
rect 1280 18675 1320 18680
rect 1280 18645 1285 18675
rect 1315 18645 1320 18675
rect 1280 18515 1320 18645
rect 1280 18485 1285 18515
rect 1315 18485 1320 18515
rect 1280 18480 1320 18485
rect 1360 18675 1400 18680
rect 1360 18645 1365 18675
rect 1395 18645 1400 18675
rect 1360 18515 1400 18645
rect 1360 18485 1365 18515
rect 1395 18485 1400 18515
rect 1360 18480 1400 18485
rect 1440 18675 1480 18680
rect 1440 18645 1445 18675
rect 1475 18645 1480 18675
rect 1440 18515 1480 18645
rect 1440 18485 1445 18515
rect 1475 18485 1480 18515
rect 1440 18480 1480 18485
rect 1520 18675 1560 18680
rect 1520 18645 1525 18675
rect 1555 18645 1560 18675
rect 1520 18515 1560 18645
rect 1520 18485 1525 18515
rect 1555 18485 1560 18515
rect 1520 18480 1560 18485
rect 1600 18675 1640 18680
rect 1600 18645 1605 18675
rect 1635 18645 1640 18675
rect 1600 18515 1640 18645
rect 1600 18485 1605 18515
rect 1635 18485 1640 18515
rect 1600 18480 1640 18485
rect 1680 18675 1720 18680
rect 1680 18645 1685 18675
rect 1715 18645 1720 18675
rect 1680 18515 1720 18645
rect 1680 18485 1685 18515
rect 1715 18485 1720 18515
rect 1680 18480 1720 18485
rect 1760 18675 1800 18680
rect 1760 18645 1765 18675
rect 1795 18645 1800 18675
rect 1760 18515 1800 18645
rect 1760 18485 1765 18515
rect 1795 18485 1800 18515
rect 1760 18480 1800 18485
rect 1840 18675 1880 18680
rect 1840 18645 1845 18675
rect 1875 18645 1880 18675
rect 1840 18515 1880 18645
rect 1840 18485 1845 18515
rect 1875 18485 1880 18515
rect 1840 18480 1880 18485
rect 1920 18675 1960 18680
rect 1920 18645 1925 18675
rect 1955 18645 1960 18675
rect 1920 18515 1960 18645
rect 1920 18485 1925 18515
rect 1955 18485 1960 18515
rect 1920 18480 1960 18485
rect 2000 18675 2040 18680
rect 2000 18645 2005 18675
rect 2035 18645 2040 18675
rect 2000 18515 2040 18645
rect 2000 18485 2005 18515
rect 2035 18485 2040 18515
rect 2000 18480 2040 18485
rect 2080 18675 2120 18680
rect 2080 18645 2085 18675
rect 2115 18645 2120 18675
rect 2080 18515 2120 18645
rect 2080 18485 2085 18515
rect 2115 18485 2120 18515
rect 2080 18480 2120 18485
rect 2160 18675 2200 18680
rect 2160 18645 2165 18675
rect 2195 18645 2200 18675
rect 2160 18515 2200 18645
rect 2160 18485 2165 18515
rect 2195 18485 2200 18515
rect 2160 18480 2200 18485
rect 2240 18675 2280 18680
rect 2240 18645 2245 18675
rect 2275 18645 2280 18675
rect 2240 18515 2280 18645
rect 2240 18485 2245 18515
rect 2275 18485 2280 18515
rect 2240 18480 2280 18485
rect 2320 18675 2360 18680
rect 2320 18645 2325 18675
rect 2355 18645 2360 18675
rect 2320 18515 2360 18645
rect 2320 18485 2325 18515
rect 2355 18485 2360 18515
rect 2320 18480 2360 18485
rect 2400 18675 2440 18680
rect 2400 18645 2405 18675
rect 2435 18645 2440 18675
rect 2400 18515 2440 18645
rect 2400 18485 2405 18515
rect 2435 18485 2440 18515
rect 2400 18480 2440 18485
rect 2480 18675 2520 18680
rect 2480 18645 2485 18675
rect 2515 18645 2520 18675
rect 2480 18515 2520 18645
rect 2480 18485 2485 18515
rect 2515 18485 2520 18515
rect 2480 18480 2520 18485
rect 2560 18675 2600 18680
rect 2560 18645 2565 18675
rect 2595 18645 2600 18675
rect 2560 18515 2600 18645
rect 2560 18485 2565 18515
rect 2595 18485 2600 18515
rect 2560 18480 2600 18485
rect 2640 18675 2680 18680
rect 2640 18645 2645 18675
rect 2675 18645 2680 18675
rect 2640 18515 2680 18645
rect 2640 18485 2645 18515
rect 2675 18485 2680 18515
rect 2640 18480 2680 18485
rect 2720 18675 2760 18680
rect 2720 18645 2725 18675
rect 2755 18645 2760 18675
rect 2720 18515 2760 18645
rect 2720 18485 2725 18515
rect 2755 18485 2760 18515
rect 2720 18480 2760 18485
rect 2800 18675 2840 18680
rect 2800 18645 2805 18675
rect 2835 18645 2840 18675
rect 2800 18515 2840 18645
rect 2800 18485 2805 18515
rect 2835 18485 2840 18515
rect 2800 18480 2840 18485
rect 2880 18675 2920 18680
rect 2880 18645 2885 18675
rect 2915 18645 2920 18675
rect 2880 18515 2920 18645
rect 2880 18485 2885 18515
rect 2915 18485 2920 18515
rect 2880 18480 2920 18485
rect 2960 18675 3000 18680
rect 2960 18645 2965 18675
rect 2995 18645 3000 18675
rect 2960 18515 3000 18645
rect 2960 18485 2965 18515
rect 2995 18485 3000 18515
rect 2960 18480 3000 18485
rect 3040 18675 3080 18680
rect 3040 18645 3045 18675
rect 3075 18645 3080 18675
rect 3040 18515 3080 18645
rect 3040 18485 3045 18515
rect 3075 18485 3080 18515
rect 3040 18480 3080 18485
rect 3120 18675 3160 18680
rect 3120 18645 3125 18675
rect 3155 18645 3160 18675
rect 3120 18515 3160 18645
rect 3120 18485 3125 18515
rect 3155 18485 3160 18515
rect 3120 18480 3160 18485
rect 3200 18675 3240 18680
rect 3200 18645 3205 18675
rect 3235 18645 3240 18675
rect 3200 18515 3240 18645
rect 3200 18485 3205 18515
rect 3235 18485 3240 18515
rect 3200 18480 3240 18485
rect 3280 18675 3320 18680
rect 3280 18645 3285 18675
rect 3315 18645 3320 18675
rect 3280 18515 3320 18645
rect 3280 18485 3285 18515
rect 3315 18485 3320 18515
rect 3280 18480 3320 18485
rect 3360 18675 3400 18680
rect 3360 18645 3365 18675
rect 3395 18645 3400 18675
rect 3360 18515 3400 18645
rect 3360 18485 3365 18515
rect 3395 18485 3400 18515
rect 3360 18480 3400 18485
rect 3440 18675 3480 18680
rect 3440 18645 3445 18675
rect 3475 18645 3480 18675
rect 3440 18515 3480 18645
rect 3440 18485 3445 18515
rect 3475 18485 3480 18515
rect 3440 18480 3480 18485
rect 3520 18675 3560 18680
rect 3520 18645 3525 18675
rect 3555 18645 3560 18675
rect 3520 18515 3560 18645
rect 3520 18485 3525 18515
rect 3555 18485 3560 18515
rect 3520 18480 3560 18485
rect 3600 18675 3640 18680
rect 3600 18645 3605 18675
rect 3635 18645 3640 18675
rect 3600 18515 3640 18645
rect 3600 18485 3605 18515
rect 3635 18485 3640 18515
rect 3600 18480 3640 18485
rect 3680 18675 3720 18680
rect 3680 18645 3685 18675
rect 3715 18645 3720 18675
rect 3680 18515 3720 18645
rect 3680 18485 3685 18515
rect 3715 18485 3720 18515
rect 3680 18480 3720 18485
rect 3760 18675 3800 18680
rect 3760 18645 3765 18675
rect 3795 18645 3800 18675
rect 3760 18515 3800 18645
rect 3760 18485 3765 18515
rect 3795 18485 3800 18515
rect 3760 18480 3800 18485
rect 3840 18675 3880 18680
rect 3840 18645 3845 18675
rect 3875 18645 3880 18675
rect 3840 18515 3880 18645
rect 3840 18485 3845 18515
rect 3875 18485 3880 18515
rect 3840 18480 3880 18485
rect 3920 18675 3960 18680
rect 3920 18645 3925 18675
rect 3955 18645 3960 18675
rect 3920 18515 3960 18645
rect 3920 18485 3925 18515
rect 3955 18485 3960 18515
rect 3920 18480 3960 18485
rect 4000 18675 4040 18680
rect 4000 18645 4005 18675
rect 4035 18645 4040 18675
rect 4000 18515 4040 18645
rect 4000 18485 4005 18515
rect 4035 18485 4040 18515
rect 4000 18480 4040 18485
rect 4080 18675 4120 18680
rect 4080 18645 4085 18675
rect 4115 18645 4120 18675
rect 4080 18515 4120 18645
rect 4080 18485 4085 18515
rect 4115 18485 4120 18515
rect 4080 18480 4120 18485
rect 4160 18675 4200 18680
rect 4160 18645 4165 18675
rect 4195 18645 4200 18675
rect 4160 18515 4200 18645
rect 4160 18485 4165 18515
rect 4195 18485 4200 18515
rect 4160 18480 4200 18485
rect 4240 18675 4280 18720
rect 4240 18645 4245 18675
rect 4275 18645 4280 18675
rect 4240 18515 4280 18645
rect 4240 18485 4245 18515
rect 4275 18485 4280 18515
rect 0 18435 40 18440
rect 0 18405 5 18435
rect 35 18405 40 18435
rect 0 18275 40 18405
rect 0 18245 5 18275
rect 35 18245 40 18275
rect 0 18240 40 18245
rect 80 18435 120 18440
rect 80 18405 85 18435
rect 115 18405 120 18435
rect 80 18275 120 18405
rect 80 18245 85 18275
rect 115 18245 120 18275
rect 80 18240 120 18245
rect 160 18435 200 18440
rect 160 18405 165 18435
rect 195 18405 200 18435
rect 160 18275 200 18405
rect 160 18245 165 18275
rect 195 18245 200 18275
rect 160 18240 200 18245
rect 240 18435 280 18440
rect 240 18405 245 18435
rect 275 18405 280 18435
rect 240 18275 280 18405
rect 240 18245 245 18275
rect 275 18245 280 18275
rect 240 18240 280 18245
rect 320 18435 360 18440
rect 320 18405 325 18435
rect 355 18405 360 18435
rect 320 18275 360 18405
rect 320 18245 325 18275
rect 355 18245 360 18275
rect 320 18240 360 18245
rect 400 18435 440 18440
rect 400 18405 405 18435
rect 435 18405 440 18435
rect 400 18275 440 18405
rect 400 18245 405 18275
rect 435 18245 440 18275
rect 400 18240 440 18245
rect 480 18435 520 18440
rect 480 18405 485 18435
rect 515 18405 520 18435
rect 480 18275 520 18405
rect 480 18245 485 18275
rect 515 18245 520 18275
rect 480 18240 520 18245
rect 560 18435 600 18440
rect 560 18405 565 18435
rect 595 18405 600 18435
rect 560 18275 600 18405
rect 560 18245 565 18275
rect 595 18245 600 18275
rect 560 18240 600 18245
rect 640 18435 680 18440
rect 640 18405 645 18435
rect 675 18405 680 18435
rect 640 18275 680 18405
rect 640 18245 645 18275
rect 675 18245 680 18275
rect 640 18240 680 18245
rect 720 18435 760 18440
rect 720 18405 725 18435
rect 755 18405 760 18435
rect 720 18275 760 18405
rect 720 18245 725 18275
rect 755 18245 760 18275
rect 720 18240 760 18245
rect 800 18435 840 18440
rect 800 18405 805 18435
rect 835 18405 840 18435
rect 800 18275 840 18405
rect 800 18245 805 18275
rect 835 18245 840 18275
rect 800 18240 840 18245
rect 880 18435 920 18440
rect 880 18405 885 18435
rect 915 18405 920 18435
rect 880 18275 920 18405
rect 880 18245 885 18275
rect 915 18245 920 18275
rect 880 18240 920 18245
rect 960 18435 1000 18440
rect 960 18405 965 18435
rect 995 18405 1000 18435
rect 960 18275 1000 18405
rect 960 18245 965 18275
rect 995 18245 1000 18275
rect 960 18240 1000 18245
rect 1040 18435 1080 18440
rect 1040 18405 1045 18435
rect 1075 18405 1080 18435
rect 1040 18275 1080 18405
rect 1040 18245 1045 18275
rect 1075 18245 1080 18275
rect 1040 18240 1080 18245
rect 1120 18435 1160 18440
rect 1120 18405 1125 18435
rect 1155 18405 1160 18435
rect 1120 18275 1160 18405
rect 1120 18245 1125 18275
rect 1155 18245 1160 18275
rect 1120 18240 1160 18245
rect 1200 18435 1240 18440
rect 1200 18405 1205 18435
rect 1235 18405 1240 18435
rect 1200 18275 1240 18405
rect 1200 18245 1205 18275
rect 1235 18245 1240 18275
rect 1200 18240 1240 18245
rect 1280 18435 1320 18440
rect 1280 18405 1285 18435
rect 1315 18405 1320 18435
rect 1280 18275 1320 18405
rect 1280 18245 1285 18275
rect 1315 18245 1320 18275
rect 1280 18240 1320 18245
rect 1360 18435 1400 18440
rect 1360 18405 1365 18435
rect 1395 18405 1400 18435
rect 1360 18275 1400 18405
rect 1360 18245 1365 18275
rect 1395 18245 1400 18275
rect 1360 18240 1400 18245
rect 1440 18435 1480 18440
rect 1440 18405 1445 18435
rect 1475 18405 1480 18435
rect 1440 18275 1480 18405
rect 1440 18245 1445 18275
rect 1475 18245 1480 18275
rect 1440 18240 1480 18245
rect 1520 18435 1560 18440
rect 1520 18405 1525 18435
rect 1555 18405 1560 18435
rect 1520 18275 1560 18405
rect 1520 18245 1525 18275
rect 1555 18245 1560 18275
rect 1520 18240 1560 18245
rect 1600 18435 1640 18440
rect 1600 18405 1605 18435
rect 1635 18405 1640 18435
rect 1600 18275 1640 18405
rect 1600 18245 1605 18275
rect 1635 18245 1640 18275
rect 1600 18240 1640 18245
rect 1680 18435 1720 18440
rect 1680 18405 1685 18435
rect 1715 18405 1720 18435
rect 1680 18275 1720 18405
rect 1680 18245 1685 18275
rect 1715 18245 1720 18275
rect 1680 18240 1720 18245
rect 1760 18435 1800 18440
rect 1760 18405 1765 18435
rect 1795 18405 1800 18435
rect 1760 18275 1800 18405
rect 1760 18245 1765 18275
rect 1795 18245 1800 18275
rect 1760 18240 1800 18245
rect 1840 18435 1880 18440
rect 1840 18405 1845 18435
rect 1875 18405 1880 18435
rect 1840 18275 1880 18405
rect 1840 18245 1845 18275
rect 1875 18245 1880 18275
rect 1840 18240 1880 18245
rect 1920 18435 1960 18440
rect 1920 18405 1925 18435
rect 1955 18405 1960 18435
rect 1920 18275 1960 18405
rect 1920 18245 1925 18275
rect 1955 18245 1960 18275
rect 1920 18240 1960 18245
rect 2000 18435 2040 18440
rect 2000 18405 2005 18435
rect 2035 18405 2040 18435
rect 2000 18275 2040 18405
rect 2000 18245 2005 18275
rect 2035 18245 2040 18275
rect 2000 18240 2040 18245
rect 2080 18435 2120 18440
rect 2080 18405 2085 18435
rect 2115 18405 2120 18435
rect 2080 18275 2120 18405
rect 2080 18245 2085 18275
rect 2115 18245 2120 18275
rect 2080 18240 2120 18245
rect 2160 18435 2200 18440
rect 2160 18405 2165 18435
rect 2195 18405 2200 18435
rect 2160 18275 2200 18405
rect 2160 18245 2165 18275
rect 2195 18245 2200 18275
rect 2160 18240 2200 18245
rect 2240 18435 2280 18440
rect 2240 18405 2245 18435
rect 2275 18405 2280 18435
rect 2240 18275 2280 18405
rect 2240 18245 2245 18275
rect 2275 18245 2280 18275
rect 2240 18240 2280 18245
rect 2320 18435 2360 18440
rect 2320 18405 2325 18435
rect 2355 18405 2360 18435
rect 2320 18275 2360 18405
rect 2320 18245 2325 18275
rect 2355 18245 2360 18275
rect 2320 18240 2360 18245
rect 2400 18435 2440 18440
rect 2400 18405 2405 18435
rect 2435 18405 2440 18435
rect 2400 18275 2440 18405
rect 2400 18245 2405 18275
rect 2435 18245 2440 18275
rect 2400 18240 2440 18245
rect 2480 18435 2520 18440
rect 2480 18405 2485 18435
rect 2515 18405 2520 18435
rect 2480 18275 2520 18405
rect 2480 18245 2485 18275
rect 2515 18245 2520 18275
rect 2480 18240 2520 18245
rect 2560 18435 2600 18440
rect 2560 18405 2565 18435
rect 2595 18405 2600 18435
rect 2560 18275 2600 18405
rect 2560 18245 2565 18275
rect 2595 18245 2600 18275
rect 2560 18240 2600 18245
rect 2640 18435 2680 18440
rect 2640 18405 2645 18435
rect 2675 18405 2680 18435
rect 2640 18275 2680 18405
rect 2640 18245 2645 18275
rect 2675 18245 2680 18275
rect 2640 18240 2680 18245
rect 2720 18435 2760 18440
rect 2720 18405 2725 18435
rect 2755 18405 2760 18435
rect 2720 18275 2760 18405
rect 2720 18245 2725 18275
rect 2755 18245 2760 18275
rect 2720 18240 2760 18245
rect 2800 18435 2840 18440
rect 2800 18405 2805 18435
rect 2835 18405 2840 18435
rect 2800 18275 2840 18405
rect 2800 18245 2805 18275
rect 2835 18245 2840 18275
rect 2800 18240 2840 18245
rect 2880 18435 2920 18440
rect 2880 18405 2885 18435
rect 2915 18405 2920 18435
rect 2880 18275 2920 18405
rect 2880 18245 2885 18275
rect 2915 18245 2920 18275
rect 2880 18240 2920 18245
rect 2960 18435 3000 18440
rect 2960 18405 2965 18435
rect 2995 18405 3000 18435
rect 2960 18275 3000 18405
rect 2960 18245 2965 18275
rect 2995 18245 3000 18275
rect 2960 18240 3000 18245
rect 3040 18435 3080 18440
rect 3040 18405 3045 18435
rect 3075 18405 3080 18435
rect 3040 18275 3080 18405
rect 3040 18245 3045 18275
rect 3075 18245 3080 18275
rect 3040 18240 3080 18245
rect 3120 18435 3160 18440
rect 3120 18405 3125 18435
rect 3155 18405 3160 18435
rect 3120 18275 3160 18405
rect 3120 18245 3125 18275
rect 3155 18245 3160 18275
rect 3120 18240 3160 18245
rect 3200 18435 3240 18440
rect 3200 18405 3205 18435
rect 3235 18405 3240 18435
rect 3200 18275 3240 18405
rect 3200 18245 3205 18275
rect 3235 18245 3240 18275
rect 3200 18240 3240 18245
rect 3280 18435 3320 18440
rect 3280 18405 3285 18435
rect 3315 18405 3320 18435
rect 3280 18275 3320 18405
rect 3280 18245 3285 18275
rect 3315 18245 3320 18275
rect 3280 18240 3320 18245
rect 3360 18435 3400 18440
rect 3360 18405 3365 18435
rect 3395 18405 3400 18435
rect 3360 18275 3400 18405
rect 3360 18245 3365 18275
rect 3395 18245 3400 18275
rect 3360 18240 3400 18245
rect 3440 18435 3480 18440
rect 3440 18405 3445 18435
rect 3475 18405 3480 18435
rect 3440 18275 3480 18405
rect 3440 18245 3445 18275
rect 3475 18245 3480 18275
rect 3440 18240 3480 18245
rect 3520 18435 3560 18440
rect 3520 18405 3525 18435
rect 3555 18405 3560 18435
rect 3520 18275 3560 18405
rect 3520 18245 3525 18275
rect 3555 18245 3560 18275
rect 3520 18240 3560 18245
rect 3600 18435 3640 18440
rect 3600 18405 3605 18435
rect 3635 18405 3640 18435
rect 3600 18275 3640 18405
rect 3600 18245 3605 18275
rect 3635 18245 3640 18275
rect 3600 18240 3640 18245
rect 3680 18435 3720 18440
rect 3680 18405 3685 18435
rect 3715 18405 3720 18435
rect 3680 18275 3720 18405
rect 3680 18245 3685 18275
rect 3715 18245 3720 18275
rect 3680 18240 3720 18245
rect 3760 18435 3800 18440
rect 3760 18405 3765 18435
rect 3795 18405 3800 18435
rect 3760 18275 3800 18405
rect 3760 18245 3765 18275
rect 3795 18245 3800 18275
rect 3760 18240 3800 18245
rect 3840 18435 3880 18440
rect 3840 18405 3845 18435
rect 3875 18405 3880 18435
rect 3840 18275 3880 18405
rect 3840 18245 3845 18275
rect 3875 18245 3880 18275
rect 3840 18240 3880 18245
rect 3920 18435 3960 18440
rect 3920 18405 3925 18435
rect 3955 18405 3960 18435
rect 3920 18275 3960 18405
rect 3920 18245 3925 18275
rect 3955 18245 3960 18275
rect 3920 18240 3960 18245
rect 4000 18435 4040 18440
rect 4000 18405 4005 18435
rect 4035 18405 4040 18435
rect 4000 18275 4040 18405
rect 4000 18245 4005 18275
rect 4035 18245 4040 18275
rect 4000 18240 4040 18245
rect 4080 18435 4120 18440
rect 4080 18405 4085 18435
rect 4115 18405 4120 18435
rect 4080 18275 4120 18405
rect 4080 18245 4085 18275
rect 4115 18245 4120 18275
rect 4080 18240 4120 18245
rect 4160 18435 4200 18440
rect 4160 18405 4165 18435
rect 4195 18405 4200 18435
rect 4160 18275 4200 18405
rect 4160 18245 4165 18275
rect 4195 18245 4200 18275
rect 4160 18240 4200 18245
rect 0 18195 40 18200
rect 0 18165 5 18195
rect 35 18165 40 18195
rect 0 18035 40 18165
rect 0 18005 5 18035
rect 35 18005 40 18035
rect 0 17875 40 18005
rect 0 17845 5 17875
rect 35 17845 40 17875
rect 0 17715 40 17845
rect 0 17685 5 17715
rect 35 17685 40 17715
rect 0 17555 40 17685
rect 0 17525 5 17555
rect 35 17525 40 17555
rect 0 17395 40 17525
rect 0 17365 5 17395
rect 35 17365 40 17395
rect 0 17235 40 17365
rect 0 17205 5 17235
rect 35 17205 40 17235
rect 0 17200 40 17205
rect 80 18195 120 18200
rect 80 18165 85 18195
rect 115 18165 120 18195
rect 80 18035 120 18165
rect 80 18005 85 18035
rect 115 18005 120 18035
rect 80 17875 120 18005
rect 80 17845 85 17875
rect 115 17845 120 17875
rect 80 17715 120 17845
rect 80 17685 85 17715
rect 115 17685 120 17715
rect 80 17555 120 17685
rect 80 17525 85 17555
rect 115 17525 120 17555
rect 80 17395 120 17525
rect 80 17365 85 17395
rect 115 17365 120 17395
rect 80 17235 120 17365
rect 80 17205 85 17235
rect 115 17205 120 17235
rect 80 17200 120 17205
rect 160 18195 200 18200
rect 160 18165 165 18195
rect 195 18165 200 18195
rect 160 18035 200 18165
rect 160 18005 165 18035
rect 195 18005 200 18035
rect 160 17875 200 18005
rect 160 17845 165 17875
rect 195 17845 200 17875
rect 160 17715 200 17845
rect 160 17685 165 17715
rect 195 17685 200 17715
rect 160 17555 200 17685
rect 160 17525 165 17555
rect 195 17525 200 17555
rect 160 17395 200 17525
rect 160 17365 165 17395
rect 195 17365 200 17395
rect 160 17235 200 17365
rect 160 17205 165 17235
rect 195 17205 200 17235
rect 160 17200 200 17205
rect 240 18195 280 18200
rect 240 18165 245 18195
rect 275 18165 280 18195
rect 240 18035 280 18165
rect 240 18005 245 18035
rect 275 18005 280 18035
rect 240 17875 280 18005
rect 240 17845 245 17875
rect 275 17845 280 17875
rect 240 17715 280 17845
rect 240 17685 245 17715
rect 275 17685 280 17715
rect 240 17555 280 17685
rect 240 17525 245 17555
rect 275 17525 280 17555
rect 240 17395 280 17525
rect 240 17365 245 17395
rect 275 17365 280 17395
rect 240 17235 280 17365
rect 240 17205 245 17235
rect 275 17205 280 17235
rect 240 17200 280 17205
rect 320 18195 360 18200
rect 320 18165 325 18195
rect 355 18165 360 18195
rect 320 18035 360 18165
rect 320 18005 325 18035
rect 355 18005 360 18035
rect 320 17875 360 18005
rect 320 17845 325 17875
rect 355 17845 360 17875
rect 320 17715 360 17845
rect 320 17685 325 17715
rect 355 17685 360 17715
rect 320 17555 360 17685
rect 320 17525 325 17555
rect 355 17525 360 17555
rect 320 17395 360 17525
rect 320 17365 325 17395
rect 355 17365 360 17395
rect 320 17235 360 17365
rect 320 17205 325 17235
rect 355 17205 360 17235
rect 320 17200 360 17205
rect 400 18195 440 18200
rect 400 18165 405 18195
rect 435 18165 440 18195
rect 400 18035 440 18165
rect 400 18005 405 18035
rect 435 18005 440 18035
rect 400 17875 440 18005
rect 400 17845 405 17875
rect 435 17845 440 17875
rect 400 17715 440 17845
rect 400 17685 405 17715
rect 435 17685 440 17715
rect 400 17555 440 17685
rect 400 17525 405 17555
rect 435 17525 440 17555
rect 400 17395 440 17525
rect 400 17365 405 17395
rect 435 17365 440 17395
rect 400 17235 440 17365
rect 400 17205 405 17235
rect 435 17205 440 17235
rect 400 17200 440 17205
rect 480 18195 520 18200
rect 480 18165 485 18195
rect 515 18165 520 18195
rect 480 18035 520 18165
rect 480 18005 485 18035
rect 515 18005 520 18035
rect 480 17875 520 18005
rect 480 17845 485 17875
rect 515 17845 520 17875
rect 480 17715 520 17845
rect 480 17685 485 17715
rect 515 17685 520 17715
rect 480 17555 520 17685
rect 480 17525 485 17555
rect 515 17525 520 17555
rect 480 17395 520 17525
rect 480 17365 485 17395
rect 515 17365 520 17395
rect 480 17235 520 17365
rect 480 17205 485 17235
rect 515 17205 520 17235
rect 480 17200 520 17205
rect 560 18195 600 18200
rect 560 18165 565 18195
rect 595 18165 600 18195
rect 560 18035 600 18165
rect 560 18005 565 18035
rect 595 18005 600 18035
rect 560 17875 600 18005
rect 560 17845 565 17875
rect 595 17845 600 17875
rect 560 17715 600 17845
rect 560 17685 565 17715
rect 595 17685 600 17715
rect 560 17555 600 17685
rect 560 17525 565 17555
rect 595 17525 600 17555
rect 560 17395 600 17525
rect 560 17365 565 17395
rect 595 17365 600 17395
rect 560 17235 600 17365
rect 560 17205 565 17235
rect 595 17205 600 17235
rect 560 17200 600 17205
rect 640 18195 680 18200
rect 640 18165 645 18195
rect 675 18165 680 18195
rect 640 18035 680 18165
rect 640 18005 645 18035
rect 675 18005 680 18035
rect 640 17875 680 18005
rect 640 17845 645 17875
rect 675 17845 680 17875
rect 640 17715 680 17845
rect 640 17685 645 17715
rect 675 17685 680 17715
rect 640 17555 680 17685
rect 640 17525 645 17555
rect 675 17525 680 17555
rect 640 17395 680 17525
rect 640 17365 645 17395
rect 675 17365 680 17395
rect 640 17235 680 17365
rect 640 17205 645 17235
rect 675 17205 680 17235
rect 640 17200 680 17205
rect 720 18195 760 18200
rect 720 18165 725 18195
rect 755 18165 760 18195
rect 720 18035 760 18165
rect 720 18005 725 18035
rect 755 18005 760 18035
rect 720 17875 760 18005
rect 720 17845 725 17875
rect 755 17845 760 17875
rect 720 17715 760 17845
rect 720 17685 725 17715
rect 755 17685 760 17715
rect 720 17555 760 17685
rect 720 17525 725 17555
rect 755 17525 760 17555
rect 720 17395 760 17525
rect 720 17365 725 17395
rect 755 17365 760 17395
rect 720 17235 760 17365
rect 720 17205 725 17235
rect 755 17205 760 17235
rect 720 17200 760 17205
rect 800 18195 840 18200
rect 800 18165 805 18195
rect 835 18165 840 18195
rect 800 18035 840 18165
rect 800 18005 805 18035
rect 835 18005 840 18035
rect 800 17875 840 18005
rect 800 17845 805 17875
rect 835 17845 840 17875
rect 800 17715 840 17845
rect 800 17685 805 17715
rect 835 17685 840 17715
rect 800 17555 840 17685
rect 800 17525 805 17555
rect 835 17525 840 17555
rect 800 17395 840 17525
rect 800 17365 805 17395
rect 835 17365 840 17395
rect 800 17235 840 17365
rect 800 17205 805 17235
rect 835 17205 840 17235
rect 800 17200 840 17205
rect 880 18195 920 18200
rect 880 18165 885 18195
rect 915 18165 920 18195
rect 880 18035 920 18165
rect 880 18005 885 18035
rect 915 18005 920 18035
rect 880 17875 920 18005
rect 880 17845 885 17875
rect 915 17845 920 17875
rect 880 17715 920 17845
rect 880 17685 885 17715
rect 915 17685 920 17715
rect 880 17555 920 17685
rect 880 17525 885 17555
rect 915 17525 920 17555
rect 880 17395 920 17525
rect 880 17365 885 17395
rect 915 17365 920 17395
rect 880 17235 920 17365
rect 880 17205 885 17235
rect 915 17205 920 17235
rect 880 17200 920 17205
rect 960 18195 1000 18200
rect 960 18165 965 18195
rect 995 18165 1000 18195
rect 960 18035 1000 18165
rect 960 18005 965 18035
rect 995 18005 1000 18035
rect 960 17875 1000 18005
rect 960 17845 965 17875
rect 995 17845 1000 17875
rect 960 17715 1000 17845
rect 960 17685 965 17715
rect 995 17685 1000 17715
rect 960 17555 1000 17685
rect 960 17525 965 17555
rect 995 17525 1000 17555
rect 960 17395 1000 17525
rect 960 17365 965 17395
rect 995 17365 1000 17395
rect 960 17235 1000 17365
rect 960 17205 965 17235
rect 995 17205 1000 17235
rect 960 17200 1000 17205
rect 1040 18195 1080 18200
rect 1040 18165 1045 18195
rect 1075 18165 1080 18195
rect 1040 18035 1080 18165
rect 1040 18005 1045 18035
rect 1075 18005 1080 18035
rect 1040 17875 1080 18005
rect 1040 17845 1045 17875
rect 1075 17845 1080 17875
rect 1040 17715 1080 17845
rect 1040 17685 1045 17715
rect 1075 17685 1080 17715
rect 1040 17555 1080 17685
rect 1040 17525 1045 17555
rect 1075 17525 1080 17555
rect 1040 17395 1080 17525
rect 1040 17365 1045 17395
rect 1075 17365 1080 17395
rect 1040 17235 1080 17365
rect 1040 17205 1045 17235
rect 1075 17205 1080 17235
rect 1040 17200 1080 17205
rect 1120 18195 1160 18200
rect 1120 18165 1125 18195
rect 1155 18165 1160 18195
rect 1120 18035 1160 18165
rect 1120 18005 1125 18035
rect 1155 18005 1160 18035
rect 1120 17875 1160 18005
rect 1120 17845 1125 17875
rect 1155 17845 1160 17875
rect 1120 17715 1160 17845
rect 1120 17685 1125 17715
rect 1155 17685 1160 17715
rect 1120 17555 1160 17685
rect 1120 17525 1125 17555
rect 1155 17525 1160 17555
rect 1120 17395 1160 17525
rect 1120 17365 1125 17395
rect 1155 17365 1160 17395
rect 1120 17235 1160 17365
rect 1120 17205 1125 17235
rect 1155 17205 1160 17235
rect 1120 17200 1160 17205
rect 1200 18195 1240 18200
rect 1200 18165 1205 18195
rect 1235 18165 1240 18195
rect 1200 18035 1240 18165
rect 1200 18005 1205 18035
rect 1235 18005 1240 18035
rect 1200 17875 1240 18005
rect 1200 17845 1205 17875
rect 1235 17845 1240 17875
rect 1200 17715 1240 17845
rect 1200 17685 1205 17715
rect 1235 17685 1240 17715
rect 1200 17555 1240 17685
rect 1200 17525 1205 17555
rect 1235 17525 1240 17555
rect 1200 17395 1240 17525
rect 1200 17365 1205 17395
rect 1235 17365 1240 17395
rect 1200 17235 1240 17365
rect 1200 17205 1205 17235
rect 1235 17205 1240 17235
rect 1200 17200 1240 17205
rect 1280 18195 1320 18200
rect 1280 18165 1285 18195
rect 1315 18165 1320 18195
rect 1280 18035 1320 18165
rect 1280 18005 1285 18035
rect 1315 18005 1320 18035
rect 1280 17875 1320 18005
rect 1280 17845 1285 17875
rect 1315 17845 1320 17875
rect 1280 17715 1320 17845
rect 1280 17685 1285 17715
rect 1315 17685 1320 17715
rect 1280 17555 1320 17685
rect 1280 17525 1285 17555
rect 1315 17525 1320 17555
rect 1280 17395 1320 17525
rect 1280 17365 1285 17395
rect 1315 17365 1320 17395
rect 1280 17235 1320 17365
rect 1280 17205 1285 17235
rect 1315 17205 1320 17235
rect 1280 17200 1320 17205
rect 1360 18195 1400 18200
rect 1360 18165 1365 18195
rect 1395 18165 1400 18195
rect 1360 18035 1400 18165
rect 1360 18005 1365 18035
rect 1395 18005 1400 18035
rect 1360 17875 1400 18005
rect 1360 17845 1365 17875
rect 1395 17845 1400 17875
rect 1360 17715 1400 17845
rect 1360 17685 1365 17715
rect 1395 17685 1400 17715
rect 1360 17555 1400 17685
rect 1360 17525 1365 17555
rect 1395 17525 1400 17555
rect 1360 17395 1400 17525
rect 1360 17365 1365 17395
rect 1395 17365 1400 17395
rect 1360 17235 1400 17365
rect 1360 17205 1365 17235
rect 1395 17205 1400 17235
rect 1360 17200 1400 17205
rect 1440 18195 1480 18200
rect 1440 18165 1445 18195
rect 1475 18165 1480 18195
rect 1440 18035 1480 18165
rect 1440 18005 1445 18035
rect 1475 18005 1480 18035
rect 1440 17875 1480 18005
rect 1440 17845 1445 17875
rect 1475 17845 1480 17875
rect 1440 17715 1480 17845
rect 1440 17685 1445 17715
rect 1475 17685 1480 17715
rect 1440 17555 1480 17685
rect 1440 17525 1445 17555
rect 1475 17525 1480 17555
rect 1440 17395 1480 17525
rect 1440 17365 1445 17395
rect 1475 17365 1480 17395
rect 1440 17235 1480 17365
rect 1440 17205 1445 17235
rect 1475 17205 1480 17235
rect 1440 17200 1480 17205
rect 1520 18195 1560 18200
rect 1520 18165 1525 18195
rect 1555 18165 1560 18195
rect 1520 18035 1560 18165
rect 1520 18005 1525 18035
rect 1555 18005 1560 18035
rect 1520 17875 1560 18005
rect 1520 17845 1525 17875
rect 1555 17845 1560 17875
rect 1520 17715 1560 17845
rect 1520 17685 1525 17715
rect 1555 17685 1560 17715
rect 1520 17555 1560 17685
rect 1520 17525 1525 17555
rect 1555 17525 1560 17555
rect 1520 17395 1560 17525
rect 1520 17365 1525 17395
rect 1555 17365 1560 17395
rect 1520 17235 1560 17365
rect 1520 17205 1525 17235
rect 1555 17205 1560 17235
rect 1520 17200 1560 17205
rect 1600 18195 1640 18200
rect 1600 18165 1605 18195
rect 1635 18165 1640 18195
rect 1600 18035 1640 18165
rect 1600 18005 1605 18035
rect 1635 18005 1640 18035
rect 1600 17875 1640 18005
rect 1600 17845 1605 17875
rect 1635 17845 1640 17875
rect 1600 17715 1640 17845
rect 1600 17685 1605 17715
rect 1635 17685 1640 17715
rect 1600 17555 1640 17685
rect 1600 17525 1605 17555
rect 1635 17525 1640 17555
rect 1600 17395 1640 17525
rect 1600 17365 1605 17395
rect 1635 17365 1640 17395
rect 1600 17235 1640 17365
rect 1600 17205 1605 17235
rect 1635 17205 1640 17235
rect 1600 17200 1640 17205
rect 1680 18195 1720 18200
rect 1680 18165 1685 18195
rect 1715 18165 1720 18195
rect 1680 18035 1720 18165
rect 1680 18005 1685 18035
rect 1715 18005 1720 18035
rect 1680 17875 1720 18005
rect 1680 17845 1685 17875
rect 1715 17845 1720 17875
rect 1680 17715 1720 17845
rect 1680 17685 1685 17715
rect 1715 17685 1720 17715
rect 1680 17555 1720 17685
rect 1680 17525 1685 17555
rect 1715 17525 1720 17555
rect 1680 17395 1720 17525
rect 1680 17365 1685 17395
rect 1715 17365 1720 17395
rect 1680 17235 1720 17365
rect 1680 17205 1685 17235
rect 1715 17205 1720 17235
rect 1680 17200 1720 17205
rect 1760 18195 1800 18200
rect 1760 18165 1765 18195
rect 1795 18165 1800 18195
rect 1760 18035 1800 18165
rect 1760 18005 1765 18035
rect 1795 18005 1800 18035
rect 1760 17875 1800 18005
rect 1760 17845 1765 17875
rect 1795 17845 1800 17875
rect 1760 17715 1800 17845
rect 1760 17685 1765 17715
rect 1795 17685 1800 17715
rect 1760 17555 1800 17685
rect 1760 17525 1765 17555
rect 1795 17525 1800 17555
rect 1760 17395 1800 17525
rect 1760 17365 1765 17395
rect 1795 17365 1800 17395
rect 1760 17235 1800 17365
rect 1760 17205 1765 17235
rect 1795 17205 1800 17235
rect 1760 17200 1800 17205
rect 1840 18195 1880 18200
rect 1840 18165 1845 18195
rect 1875 18165 1880 18195
rect 1840 18035 1880 18165
rect 1840 18005 1845 18035
rect 1875 18005 1880 18035
rect 1840 17875 1880 18005
rect 1840 17845 1845 17875
rect 1875 17845 1880 17875
rect 1840 17715 1880 17845
rect 1840 17685 1845 17715
rect 1875 17685 1880 17715
rect 1840 17555 1880 17685
rect 1840 17525 1845 17555
rect 1875 17525 1880 17555
rect 1840 17395 1880 17525
rect 1840 17365 1845 17395
rect 1875 17365 1880 17395
rect 1840 17235 1880 17365
rect 1840 17205 1845 17235
rect 1875 17205 1880 17235
rect 1840 17200 1880 17205
rect 1920 18195 1960 18200
rect 1920 18165 1925 18195
rect 1955 18165 1960 18195
rect 1920 18035 1960 18165
rect 1920 18005 1925 18035
rect 1955 18005 1960 18035
rect 1920 17875 1960 18005
rect 1920 17845 1925 17875
rect 1955 17845 1960 17875
rect 1920 17715 1960 17845
rect 1920 17685 1925 17715
rect 1955 17685 1960 17715
rect 1920 17555 1960 17685
rect 1920 17525 1925 17555
rect 1955 17525 1960 17555
rect 1920 17395 1960 17525
rect 1920 17365 1925 17395
rect 1955 17365 1960 17395
rect 1920 17235 1960 17365
rect 1920 17205 1925 17235
rect 1955 17205 1960 17235
rect 1920 17200 1960 17205
rect 2000 18195 2040 18200
rect 2000 18165 2005 18195
rect 2035 18165 2040 18195
rect 2000 18035 2040 18165
rect 2000 18005 2005 18035
rect 2035 18005 2040 18035
rect 2000 17875 2040 18005
rect 2000 17845 2005 17875
rect 2035 17845 2040 17875
rect 2000 17715 2040 17845
rect 2000 17685 2005 17715
rect 2035 17685 2040 17715
rect 2000 17555 2040 17685
rect 2000 17525 2005 17555
rect 2035 17525 2040 17555
rect 2000 17395 2040 17525
rect 2000 17365 2005 17395
rect 2035 17365 2040 17395
rect 2000 17235 2040 17365
rect 2000 17205 2005 17235
rect 2035 17205 2040 17235
rect 2000 17200 2040 17205
rect 2080 18195 2120 18200
rect 2080 18165 2085 18195
rect 2115 18165 2120 18195
rect 2080 18035 2120 18165
rect 2080 18005 2085 18035
rect 2115 18005 2120 18035
rect 2080 17875 2120 18005
rect 2080 17845 2085 17875
rect 2115 17845 2120 17875
rect 2080 17715 2120 17845
rect 2080 17685 2085 17715
rect 2115 17685 2120 17715
rect 2080 17555 2120 17685
rect 2080 17525 2085 17555
rect 2115 17525 2120 17555
rect 2080 17395 2120 17525
rect 2080 17365 2085 17395
rect 2115 17365 2120 17395
rect 2080 17235 2120 17365
rect 2080 17205 2085 17235
rect 2115 17205 2120 17235
rect 2080 17200 2120 17205
rect 2160 18195 2200 18200
rect 2160 18165 2165 18195
rect 2195 18165 2200 18195
rect 2160 18035 2200 18165
rect 2160 18005 2165 18035
rect 2195 18005 2200 18035
rect 2160 17875 2200 18005
rect 2160 17845 2165 17875
rect 2195 17845 2200 17875
rect 2160 17715 2200 17845
rect 2160 17685 2165 17715
rect 2195 17685 2200 17715
rect 2160 17555 2200 17685
rect 2160 17525 2165 17555
rect 2195 17525 2200 17555
rect 2160 17395 2200 17525
rect 2160 17365 2165 17395
rect 2195 17365 2200 17395
rect 2160 17235 2200 17365
rect 2160 17205 2165 17235
rect 2195 17205 2200 17235
rect 2160 17200 2200 17205
rect 2240 18195 2280 18200
rect 2240 18165 2245 18195
rect 2275 18165 2280 18195
rect 2240 18035 2280 18165
rect 2240 18005 2245 18035
rect 2275 18005 2280 18035
rect 2240 17875 2280 18005
rect 2240 17845 2245 17875
rect 2275 17845 2280 17875
rect 2240 17715 2280 17845
rect 2240 17685 2245 17715
rect 2275 17685 2280 17715
rect 2240 17555 2280 17685
rect 2240 17525 2245 17555
rect 2275 17525 2280 17555
rect 2240 17395 2280 17525
rect 2240 17365 2245 17395
rect 2275 17365 2280 17395
rect 2240 17235 2280 17365
rect 2240 17205 2245 17235
rect 2275 17205 2280 17235
rect 2240 17200 2280 17205
rect 2320 18195 2360 18200
rect 2320 18165 2325 18195
rect 2355 18165 2360 18195
rect 2320 18035 2360 18165
rect 2320 18005 2325 18035
rect 2355 18005 2360 18035
rect 2320 17875 2360 18005
rect 2320 17845 2325 17875
rect 2355 17845 2360 17875
rect 2320 17715 2360 17845
rect 2320 17685 2325 17715
rect 2355 17685 2360 17715
rect 2320 17555 2360 17685
rect 2320 17525 2325 17555
rect 2355 17525 2360 17555
rect 2320 17395 2360 17525
rect 2320 17365 2325 17395
rect 2355 17365 2360 17395
rect 2320 17235 2360 17365
rect 2320 17205 2325 17235
rect 2355 17205 2360 17235
rect 2320 17200 2360 17205
rect 2400 18195 2440 18200
rect 2400 18165 2405 18195
rect 2435 18165 2440 18195
rect 2400 18035 2440 18165
rect 2400 18005 2405 18035
rect 2435 18005 2440 18035
rect 2400 17875 2440 18005
rect 2400 17845 2405 17875
rect 2435 17845 2440 17875
rect 2400 17715 2440 17845
rect 2400 17685 2405 17715
rect 2435 17685 2440 17715
rect 2400 17555 2440 17685
rect 2400 17525 2405 17555
rect 2435 17525 2440 17555
rect 2400 17395 2440 17525
rect 2400 17365 2405 17395
rect 2435 17365 2440 17395
rect 2400 17235 2440 17365
rect 2400 17205 2405 17235
rect 2435 17205 2440 17235
rect 2400 17200 2440 17205
rect 2480 18195 2520 18200
rect 2480 18165 2485 18195
rect 2515 18165 2520 18195
rect 2480 18035 2520 18165
rect 2480 18005 2485 18035
rect 2515 18005 2520 18035
rect 2480 17875 2520 18005
rect 2480 17845 2485 17875
rect 2515 17845 2520 17875
rect 2480 17715 2520 17845
rect 2480 17685 2485 17715
rect 2515 17685 2520 17715
rect 2480 17555 2520 17685
rect 2480 17525 2485 17555
rect 2515 17525 2520 17555
rect 2480 17395 2520 17525
rect 2480 17365 2485 17395
rect 2515 17365 2520 17395
rect 2480 17235 2520 17365
rect 2480 17205 2485 17235
rect 2515 17205 2520 17235
rect 2480 17200 2520 17205
rect 2560 18195 2600 18200
rect 2560 18165 2565 18195
rect 2595 18165 2600 18195
rect 2560 18035 2600 18165
rect 2560 18005 2565 18035
rect 2595 18005 2600 18035
rect 2560 17875 2600 18005
rect 2560 17845 2565 17875
rect 2595 17845 2600 17875
rect 2560 17715 2600 17845
rect 2560 17685 2565 17715
rect 2595 17685 2600 17715
rect 2560 17555 2600 17685
rect 2560 17525 2565 17555
rect 2595 17525 2600 17555
rect 2560 17395 2600 17525
rect 2560 17365 2565 17395
rect 2595 17365 2600 17395
rect 2560 17235 2600 17365
rect 2560 17205 2565 17235
rect 2595 17205 2600 17235
rect 2560 17200 2600 17205
rect 2640 18195 2680 18200
rect 2640 18165 2645 18195
rect 2675 18165 2680 18195
rect 2640 18035 2680 18165
rect 2640 18005 2645 18035
rect 2675 18005 2680 18035
rect 2640 17875 2680 18005
rect 2640 17845 2645 17875
rect 2675 17845 2680 17875
rect 2640 17715 2680 17845
rect 2640 17685 2645 17715
rect 2675 17685 2680 17715
rect 2640 17555 2680 17685
rect 2640 17525 2645 17555
rect 2675 17525 2680 17555
rect 2640 17395 2680 17525
rect 2640 17365 2645 17395
rect 2675 17365 2680 17395
rect 2640 17235 2680 17365
rect 2640 17205 2645 17235
rect 2675 17205 2680 17235
rect 2640 17200 2680 17205
rect 2720 18195 2760 18200
rect 2720 18165 2725 18195
rect 2755 18165 2760 18195
rect 2720 18035 2760 18165
rect 2720 18005 2725 18035
rect 2755 18005 2760 18035
rect 2720 17875 2760 18005
rect 2720 17845 2725 17875
rect 2755 17845 2760 17875
rect 2720 17715 2760 17845
rect 2720 17685 2725 17715
rect 2755 17685 2760 17715
rect 2720 17555 2760 17685
rect 2720 17525 2725 17555
rect 2755 17525 2760 17555
rect 2720 17395 2760 17525
rect 2720 17365 2725 17395
rect 2755 17365 2760 17395
rect 2720 17235 2760 17365
rect 2720 17205 2725 17235
rect 2755 17205 2760 17235
rect 2720 17200 2760 17205
rect 2800 18195 2840 18200
rect 2800 18165 2805 18195
rect 2835 18165 2840 18195
rect 2800 18035 2840 18165
rect 2800 18005 2805 18035
rect 2835 18005 2840 18035
rect 2800 17875 2840 18005
rect 2800 17845 2805 17875
rect 2835 17845 2840 17875
rect 2800 17715 2840 17845
rect 2800 17685 2805 17715
rect 2835 17685 2840 17715
rect 2800 17555 2840 17685
rect 2800 17525 2805 17555
rect 2835 17525 2840 17555
rect 2800 17395 2840 17525
rect 2800 17365 2805 17395
rect 2835 17365 2840 17395
rect 2800 17235 2840 17365
rect 2800 17205 2805 17235
rect 2835 17205 2840 17235
rect 2800 17200 2840 17205
rect 2880 18195 2920 18200
rect 2880 18165 2885 18195
rect 2915 18165 2920 18195
rect 2880 18035 2920 18165
rect 2880 18005 2885 18035
rect 2915 18005 2920 18035
rect 2880 17875 2920 18005
rect 2880 17845 2885 17875
rect 2915 17845 2920 17875
rect 2880 17715 2920 17845
rect 2880 17685 2885 17715
rect 2915 17685 2920 17715
rect 2880 17555 2920 17685
rect 2880 17525 2885 17555
rect 2915 17525 2920 17555
rect 2880 17395 2920 17525
rect 2880 17365 2885 17395
rect 2915 17365 2920 17395
rect 2880 17235 2920 17365
rect 2880 17205 2885 17235
rect 2915 17205 2920 17235
rect 2880 17200 2920 17205
rect 2960 18195 3000 18200
rect 2960 18165 2965 18195
rect 2995 18165 3000 18195
rect 2960 18035 3000 18165
rect 2960 18005 2965 18035
rect 2995 18005 3000 18035
rect 2960 17875 3000 18005
rect 2960 17845 2965 17875
rect 2995 17845 3000 17875
rect 2960 17715 3000 17845
rect 2960 17685 2965 17715
rect 2995 17685 3000 17715
rect 2960 17555 3000 17685
rect 2960 17525 2965 17555
rect 2995 17525 3000 17555
rect 2960 17395 3000 17525
rect 2960 17365 2965 17395
rect 2995 17365 3000 17395
rect 2960 17235 3000 17365
rect 2960 17205 2965 17235
rect 2995 17205 3000 17235
rect 2960 17200 3000 17205
rect 3040 18195 3080 18200
rect 3040 18165 3045 18195
rect 3075 18165 3080 18195
rect 3040 18035 3080 18165
rect 3040 18005 3045 18035
rect 3075 18005 3080 18035
rect 3040 17875 3080 18005
rect 3040 17845 3045 17875
rect 3075 17845 3080 17875
rect 3040 17715 3080 17845
rect 3040 17685 3045 17715
rect 3075 17685 3080 17715
rect 3040 17555 3080 17685
rect 3040 17525 3045 17555
rect 3075 17525 3080 17555
rect 3040 17395 3080 17525
rect 3040 17365 3045 17395
rect 3075 17365 3080 17395
rect 3040 17235 3080 17365
rect 3040 17205 3045 17235
rect 3075 17205 3080 17235
rect 3040 17200 3080 17205
rect 3120 18195 3160 18200
rect 3120 18165 3125 18195
rect 3155 18165 3160 18195
rect 3120 18035 3160 18165
rect 3120 18005 3125 18035
rect 3155 18005 3160 18035
rect 3120 17875 3160 18005
rect 3120 17845 3125 17875
rect 3155 17845 3160 17875
rect 3120 17715 3160 17845
rect 3120 17685 3125 17715
rect 3155 17685 3160 17715
rect 3120 17555 3160 17685
rect 3120 17525 3125 17555
rect 3155 17525 3160 17555
rect 3120 17395 3160 17525
rect 3120 17365 3125 17395
rect 3155 17365 3160 17395
rect 3120 17235 3160 17365
rect 3120 17205 3125 17235
rect 3155 17205 3160 17235
rect 3120 17200 3160 17205
rect 3200 18195 3240 18200
rect 3200 18165 3205 18195
rect 3235 18165 3240 18195
rect 3200 18035 3240 18165
rect 3200 18005 3205 18035
rect 3235 18005 3240 18035
rect 3200 17875 3240 18005
rect 3200 17845 3205 17875
rect 3235 17845 3240 17875
rect 3200 17715 3240 17845
rect 3200 17685 3205 17715
rect 3235 17685 3240 17715
rect 3200 17555 3240 17685
rect 3200 17525 3205 17555
rect 3235 17525 3240 17555
rect 3200 17395 3240 17525
rect 3200 17365 3205 17395
rect 3235 17365 3240 17395
rect 3200 17235 3240 17365
rect 3200 17205 3205 17235
rect 3235 17205 3240 17235
rect 3200 17200 3240 17205
rect 3280 18195 3320 18200
rect 3280 18165 3285 18195
rect 3315 18165 3320 18195
rect 3280 18035 3320 18165
rect 3280 18005 3285 18035
rect 3315 18005 3320 18035
rect 3280 17875 3320 18005
rect 3280 17845 3285 17875
rect 3315 17845 3320 17875
rect 3280 17715 3320 17845
rect 3280 17685 3285 17715
rect 3315 17685 3320 17715
rect 3280 17555 3320 17685
rect 3280 17525 3285 17555
rect 3315 17525 3320 17555
rect 3280 17395 3320 17525
rect 3280 17365 3285 17395
rect 3315 17365 3320 17395
rect 3280 17235 3320 17365
rect 3280 17205 3285 17235
rect 3315 17205 3320 17235
rect 3280 17200 3320 17205
rect 3360 18195 3400 18200
rect 3360 18165 3365 18195
rect 3395 18165 3400 18195
rect 3360 18035 3400 18165
rect 3360 18005 3365 18035
rect 3395 18005 3400 18035
rect 3360 17875 3400 18005
rect 3360 17845 3365 17875
rect 3395 17845 3400 17875
rect 3360 17715 3400 17845
rect 3360 17685 3365 17715
rect 3395 17685 3400 17715
rect 3360 17555 3400 17685
rect 3360 17525 3365 17555
rect 3395 17525 3400 17555
rect 3360 17395 3400 17525
rect 3360 17365 3365 17395
rect 3395 17365 3400 17395
rect 3360 17235 3400 17365
rect 3360 17205 3365 17235
rect 3395 17205 3400 17235
rect 3360 17200 3400 17205
rect 3440 18195 3480 18200
rect 3440 18165 3445 18195
rect 3475 18165 3480 18195
rect 3440 18035 3480 18165
rect 3440 18005 3445 18035
rect 3475 18005 3480 18035
rect 3440 17875 3480 18005
rect 3440 17845 3445 17875
rect 3475 17845 3480 17875
rect 3440 17715 3480 17845
rect 3440 17685 3445 17715
rect 3475 17685 3480 17715
rect 3440 17555 3480 17685
rect 3440 17525 3445 17555
rect 3475 17525 3480 17555
rect 3440 17395 3480 17525
rect 3440 17365 3445 17395
rect 3475 17365 3480 17395
rect 3440 17235 3480 17365
rect 3440 17205 3445 17235
rect 3475 17205 3480 17235
rect 3440 17200 3480 17205
rect 3520 18195 3560 18200
rect 3520 18165 3525 18195
rect 3555 18165 3560 18195
rect 3520 18035 3560 18165
rect 3520 18005 3525 18035
rect 3555 18005 3560 18035
rect 3520 17875 3560 18005
rect 3520 17845 3525 17875
rect 3555 17845 3560 17875
rect 3520 17715 3560 17845
rect 3520 17685 3525 17715
rect 3555 17685 3560 17715
rect 3520 17555 3560 17685
rect 3520 17525 3525 17555
rect 3555 17525 3560 17555
rect 3520 17395 3560 17525
rect 3520 17365 3525 17395
rect 3555 17365 3560 17395
rect 3520 17235 3560 17365
rect 3520 17205 3525 17235
rect 3555 17205 3560 17235
rect 3520 17200 3560 17205
rect 3600 18195 3640 18200
rect 3600 18165 3605 18195
rect 3635 18165 3640 18195
rect 3600 18035 3640 18165
rect 3600 18005 3605 18035
rect 3635 18005 3640 18035
rect 3600 17875 3640 18005
rect 3600 17845 3605 17875
rect 3635 17845 3640 17875
rect 3600 17715 3640 17845
rect 3600 17685 3605 17715
rect 3635 17685 3640 17715
rect 3600 17555 3640 17685
rect 3600 17525 3605 17555
rect 3635 17525 3640 17555
rect 3600 17395 3640 17525
rect 3600 17365 3605 17395
rect 3635 17365 3640 17395
rect 3600 17235 3640 17365
rect 3600 17205 3605 17235
rect 3635 17205 3640 17235
rect 3600 17200 3640 17205
rect 3680 18195 3720 18200
rect 3680 18165 3685 18195
rect 3715 18165 3720 18195
rect 3680 18035 3720 18165
rect 3680 18005 3685 18035
rect 3715 18005 3720 18035
rect 3680 17875 3720 18005
rect 3680 17845 3685 17875
rect 3715 17845 3720 17875
rect 3680 17715 3720 17845
rect 3680 17685 3685 17715
rect 3715 17685 3720 17715
rect 3680 17555 3720 17685
rect 3680 17525 3685 17555
rect 3715 17525 3720 17555
rect 3680 17395 3720 17525
rect 3680 17365 3685 17395
rect 3715 17365 3720 17395
rect 3680 17235 3720 17365
rect 3680 17205 3685 17235
rect 3715 17205 3720 17235
rect 3680 17200 3720 17205
rect 3760 18195 3800 18200
rect 3760 18165 3765 18195
rect 3795 18165 3800 18195
rect 3760 18035 3800 18165
rect 3760 18005 3765 18035
rect 3795 18005 3800 18035
rect 3760 17875 3800 18005
rect 3760 17845 3765 17875
rect 3795 17845 3800 17875
rect 3760 17715 3800 17845
rect 3760 17685 3765 17715
rect 3795 17685 3800 17715
rect 3760 17555 3800 17685
rect 3760 17525 3765 17555
rect 3795 17525 3800 17555
rect 3760 17395 3800 17525
rect 3760 17365 3765 17395
rect 3795 17365 3800 17395
rect 3760 17235 3800 17365
rect 3760 17205 3765 17235
rect 3795 17205 3800 17235
rect 3760 17200 3800 17205
rect 3840 18195 3880 18200
rect 3840 18165 3845 18195
rect 3875 18165 3880 18195
rect 3840 18035 3880 18165
rect 3840 18005 3845 18035
rect 3875 18005 3880 18035
rect 3840 17875 3880 18005
rect 3840 17845 3845 17875
rect 3875 17845 3880 17875
rect 3840 17715 3880 17845
rect 3840 17685 3845 17715
rect 3875 17685 3880 17715
rect 3840 17555 3880 17685
rect 3840 17525 3845 17555
rect 3875 17525 3880 17555
rect 3840 17395 3880 17525
rect 3840 17365 3845 17395
rect 3875 17365 3880 17395
rect 3840 17235 3880 17365
rect 3840 17205 3845 17235
rect 3875 17205 3880 17235
rect 3840 17200 3880 17205
rect 3920 18195 3960 18200
rect 3920 18165 3925 18195
rect 3955 18165 3960 18195
rect 3920 18035 3960 18165
rect 3920 18005 3925 18035
rect 3955 18005 3960 18035
rect 3920 17875 3960 18005
rect 3920 17845 3925 17875
rect 3955 17845 3960 17875
rect 3920 17715 3960 17845
rect 3920 17685 3925 17715
rect 3955 17685 3960 17715
rect 3920 17555 3960 17685
rect 3920 17525 3925 17555
rect 3955 17525 3960 17555
rect 3920 17395 3960 17525
rect 3920 17365 3925 17395
rect 3955 17365 3960 17395
rect 3920 17235 3960 17365
rect 3920 17205 3925 17235
rect 3955 17205 3960 17235
rect 3920 17200 3960 17205
rect 4000 18195 4040 18200
rect 4000 18165 4005 18195
rect 4035 18165 4040 18195
rect 4000 18035 4040 18165
rect 4000 18005 4005 18035
rect 4035 18005 4040 18035
rect 4000 17875 4040 18005
rect 4000 17845 4005 17875
rect 4035 17845 4040 17875
rect 4000 17715 4040 17845
rect 4000 17685 4005 17715
rect 4035 17685 4040 17715
rect 4000 17555 4040 17685
rect 4000 17525 4005 17555
rect 4035 17525 4040 17555
rect 4000 17395 4040 17525
rect 4000 17365 4005 17395
rect 4035 17365 4040 17395
rect 4000 17235 4040 17365
rect 4000 17205 4005 17235
rect 4035 17205 4040 17235
rect 4000 17200 4040 17205
rect 4080 18195 4120 18200
rect 4080 18165 4085 18195
rect 4115 18165 4120 18195
rect 4080 18035 4120 18165
rect 4080 18005 4085 18035
rect 4115 18005 4120 18035
rect 4080 17875 4120 18005
rect 4080 17845 4085 17875
rect 4115 17845 4120 17875
rect 4080 17715 4120 17845
rect 4080 17685 4085 17715
rect 4115 17685 4120 17715
rect 4080 17555 4120 17685
rect 4080 17525 4085 17555
rect 4115 17525 4120 17555
rect 4080 17395 4120 17525
rect 4080 17365 4085 17395
rect 4115 17365 4120 17395
rect 4080 17235 4120 17365
rect 4080 17205 4085 17235
rect 4115 17205 4120 17235
rect 4080 17200 4120 17205
rect 4160 18195 4200 18200
rect 4160 18165 4165 18195
rect 4195 18165 4200 18195
rect 4160 18035 4200 18165
rect 4160 18005 4165 18035
rect 4195 18005 4200 18035
rect 4160 17875 4200 18005
rect 4160 17845 4165 17875
rect 4195 17845 4200 17875
rect 4160 17715 4200 17845
rect 4160 17685 4165 17715
rect 4195 17685 4200 17715
rect 4160 17555 4200 17685
rect 4160 17525 4165 17555
rect 4195 17525 4200 17555
rect 4160 17395 4200 17525
rect 4160 17365 4165 17395
rect 4195 17365 4200 17395
rect 4160 17235 4200 17365
rect 4160 17205 4165 17235
rect 4195 17205 4200 17235
rect 4160 17200 4200 17205
rect 0 17155 40 17160
rect 0 17125 5 17155
rect 35 17125 40 17155
rect 0 16995 40 17125
rect 0 16965 5 16995
rect 35 16965 40 16995
rect 0 16960 40 16965
rect 80 17155 120 17160
rect 80 17125 85 17155
rect 115 17125 120 17155
rect 80 16995 120 17125
rect 80 16965 85 16995
rect 115 16965 120 16995
rect 80 16960 120 16965
rect 160 17155 200 17160
rect 160 17125 165 17155
rect 195 17125 200 17155
rect 160 16995 200 17125
rect 160 16965 165 16995
rect 195 16965 200 16995
rect 160 16960 200 16965
rect 240 17155 280 17160
rect 240 17125 245 17155
rect 275 17125 280 17155
rect 240 16995 280 17125
rect 240 16965 245 16995
rect 275 16965 280 16995
rect 240 16960 280 16965
rect 320 17155 360 17160
rect 320 17125 325 17155
rect 355 17125 360 17155
rect 320 16995 360 17125
rect 320 16965 325 16995
rect 355 16965 360 16995
rect 320 16960 360 16965
rect 400 17155 440 17160
rect 400 17125 405 17155
rect 435 17125 440 17155
rect 400 16995 440 17125
rect 400 16965 405 16995
rect 435 16965 440 16995
rect 400 16960 440 16965
rect 480 17155 520 17160
rect 480 17125 485 17155
rect 515 17125 520 17155
rect 480 16995 520 17125
rect 480 16965 485 16995
rect 515 16965 520 16995
rect 480 16960 520 16965
rect 560 17155 600 17160
rect 560 17125 565 17155
rect 595 17125 600 17155
rect 560 16995 600 17125
rect 560 16965 565 16995
rect 595 16965 600 16995
rect 560 16960 600 16965
rect 640 17155 680 17160
rect 640 17125 645 17155
rect 675 17125 680 17155
rect 640 16995 680 17125
rect 640 16965 645 16995
rect 675 16965 680 16995
rect 640 16960 680 16965
rect 720 17155 760 17160
rect 720 17125 725 17155
rect 755 17125 760 17155
rect 720 16995 760 17125
rect 720 16965 725 16995
rect 755 16965 760 16995
rect 720 16960 760 16965
rect 800 17155 840 17160
rect 800 17125 805 17155
rect 835 17125 840 17155
rect 800 16995 840 17125
rect 800 16965 805 16995
rect 835 16965 840 16995
rect 800 16960 840 16965
rect 880 17155 920 17160
rect 880 17125 885 17155
rect 915 17125 920 17155
rect 880 16995 920 17125
rect 880 16965 885 16995
rect 915 16965 920 16995
rect 880 16960 920 16965
rect 960 17155 1000 17160
rect 960 17125 965 17155
rect 995 17125 1000 17155
rect 960 16995 1000 17125
rect 960 16965 965 16995
rect 995 16965 1000 16995
rect 960 16960 1000 16965
rect 1040 17155 1080 17160
rect 1040 17125 1045 17155
rect 1075 17125 1080 17155
rect 1040 16995 1080 17125
rect 1040 16965 1045 16995
rect 1075 16965 1080 16995
rect 1040 16960 1080 16965
rect 1120 17155 1160 17160
rect 1120 17125 1125 17155
rect 1155 17125 1160 17155
rect 1120 16995 1160 17125
rect 1120 16965 1125 16995
rect 1155 16965 1160 16995
rect 1120 16960 1160 16965
rect 1200 17155 1240 17160
rect 1200 17125 1205 17155
rect 1235 17125 1240 17155
rect 1200 16995 1240 17125
rect 1200 16965 1205 16995
rect 1235 16965 1240 16995
rect 1200 16960 1240 16965
rect 1280 17155 1320 17160
rect 1280 17125 1285 17155
rect 1315 17125 1320 17155
rect 1280 16995 1320 17125
rect 1280 16965 1285 16995
rect 1315 16965 1320 16995
rect 1280 16960 1320 16965
rect 1360 17155 1400 17160
rect 1360 17125 1365 17155
rect 1395 17125 1400 17155
rect 1360 16995 1400 17125
rect 1360 16965 1365 16995
rect 1395 16965 1400 16995
rect 1360 16960 1400 16965
rect 1440 17155 1480 17160
rect 1440 17125 1445 17155
rect 1475 17125 1480 17155
rect 1440 16995 1480 17125
rect 1440 16965 1445 16995
rect 1475 16965 1480 16995
rect 1440 16960 1480 16965
rect 1520 17155 1560 17160
rect 1520 17125 1525 17155
rect 1555 17125 1560 17155
rect 1520 16995 1560 17125
rect 1520 16965 1525 16995
rect 1555 16965 1560 16995
rect 1520 16960 1560 16965
rect 1600 17155 1640 17160
rect 1600 17125 1605 17155
rect 1635 17125 1640 17155
rect 1600 16995 1640 17125
rect 1600 16965 1605 16995
rect 1635 16965 1640 16995
rect 1600 16960 1640 16965
rect 1680 17155 1720 17160
rect 1680 17125 1685 17155
rect 1715 17125 1720 17155
rect 1680 16995 1720 17125
rect 1680 16965 1685 16995
rect 1715 16965 1720 16995
rect 1680 16960 1720 16965
rect 1760 17155 1800 17160
rect 1760 17125 1765 17155
rect 1795 17125 1800 17155
rect 1760 16995 1800 17125
rect 1760 16965 1765 16995
rect 1795 16965 1800 16995
rect 1760 16960 1800 16965
rect 1840 17155 1880 17160
rect 1840 17125 1845 17155
rect 1875 17125 1880 17155
rect 1840 16995 1880 17125
rect 1840 16965 1845 16995
rect 1875 16965 1880 16995
rect 1840 16960 1880 16965
rect 1920 17155 1960 17160
rect 1920 17125 1925 17155
rect 1955 17125 1960 17155
rect 1920 16995 1960 17125
rect 1920 16965 1925 16995
rect 1955 16965 1960 16995
rect 1920 16960 1960 16965
rect 2000 17155 2040 17160
rect 2000 17125 2005 17155
rect 2035 17125 2040 17155
rect 2000 16995 2040 17125
rect 2000 16965 2005 16995
rect 2035 16965 2040 16995
rect 2000 16960 2040 16965
rect 2080 17155 2120 17160
rect 2080 17125 2085 17155
rect 2115 17125 2120 17155
rect 2080 16995 2120 17125
rect 2080 16965 2085 16995
rect 2115 16965 2120 16995
rect 2080 16960 2120 16965
rect 2160 17155 2200 17160
rect 2160 17125 2165 17155
rect 2195 17125 2200 17155
rect 2160 16995 2200 17125
rect 2160 16965 2165 16995
rect 2195 16965 2200 16995
rect 2160 16960 2200 16965
rect 2240 17155 2280 17160
rect 2240 17125 2245 17155
rect 2275 17125 2280 17155
rect 2240 16995 2280 17125
rect 2240 16965 2245 16995
rect 2275 16965 2280 16995
rect 2240 16960 2280 16965
rect 2320 17155 2360 17160
rect 2320 17125 2325 17155
rect 2355 17125 2360 17155
rect 2320 16995 2360 17125
rect 2320 16965 2325 16995
rect 2355 16965 2360 16995
rect 2320 16960 2360 16965
rect 2400 17155 2440 17160
rect 2400 17125 2405 17155
rect 2435 17125 2440 17155
rect 2400 16995 2440 17125
rect 2400 16965 2405 16995
rect 2435 16965 2440 16995
rect 2400 16960 2440 16965
rect 2480 17155 2520 17160
rect 2480 17125 2485 17155
rect 2515 17125 2520 17155
rect 2480 16995 2520 17125
rect 2480 16965 2485 16995
rect 2515 16965 2520 16995
rect 2480 16960 2520 16965
rect 2560 17155 2600 17160
rect 2560 17125 2565 17155
rect 2595 17125 2600 17155
rect 2560 16995 2600 17125
rect 2560 16965 2565 16995
rect 2595 16965 2600 16995
rect 2560 16960 2600 16965
rect 2640 17155 2680 17160
rect 2640 17125 2645 17155
rect 2675 17125 2680 17155
rect 2640 16995 2680 17125
rect 2640 16965 2645 16995
rect 2675 16965 2680 16995
rect 2640 16960 2680 16965
rect 2720 17155 2760 17160
rect 2720 17125 2725 17155
rect 2755 17125 2760 17155
rect 2720 16995 2760 17125
rect 2720 16965 2725 16995
rect 2755 16965 2760 16995
rect 2720 16960 2760 16965
rect 2800 17155 2840 17160
rect 2800 17125 2805 17155
rect 2835 17125 2840 17155
rect 2800 16995 2840 17125
rect 2800 16965 2805 16995
rect 2835 16965 2840 16995
rect 2800 16960 2840 16965
rect 2880 17155 2920 17160
rect 2880 17125 2885 17155
rect 2915 17125 2920 17155
rect 2880 16995 2920 17125
rect 2880 16965 2885 16995
rect 2915 16965 2920 16995
rect 2880 16960 2920 16965
rect 2960 17155 3000 17160
rect 2960 17125 2965 17155
rect 2995 17125 3000 17155
rect 2960 16995 3000 17125
rect 2960 16965 2965 16995
rect 2995 16965 3000 16995
rect 2960 16960 3000 16965
rect 3040 17155 3080 17160
rect 3040 17125 3045 17155
rect 3075 17125 3080 17155
rect 3040 16995 3080 17125
rect 3040 16965 3045 16995
rect 3075 16965 3080 16995
rect 3040 16960 3080 16965
rect 3120 17155 3160 17160
rect 3120 17125 3125 17155
rect 3155 17125 3160 17155
rect 3120 16995 3160 17125
rect 3120 16965 3125 16995
rect 3155 16965 3160 16995
rect 3120 16960 3160 16965
rect 3200 17155 3240 17160
rect 3200 17125 3205 17155
rect 3235 17125 3240 17155
rect 3200 16995 3240 17125
rect 3200 16965 3205 16995
rect 3235 16965 3240 16995
rect 3200 16960 3240 16965
rect 3280 17155 3320 17160
rect 3280 17125 3285 17155
rect 3315 17125 3320 17155
rect 3280 16995 3320 17125
rect 3280 16965 3285 16995
rect 3315 16965 3320 16995
rect 3280 16960 3320 16965
rect 3360 17155 3400 17160
rect 3360 17125 3365 17155
rect 3395 17125 3400 17155
rect 3360 16995 3400 17125
rect 3360 16965 3365 16995
rect 3395 16965 3400 16995
rect 3360 16960 3400 16965
rect 3440 17155 3480 17160
rect 3440 17125 3445 17155
rect 3475 17125 3480 17155
rect 3440 16995 3480 17125
rect 3440 16965 3445 16995
rect 3475 16965 3480 16995
rect 3440 16960 3480 16965
rect 3520 17155 3560 17160
rect 3520 17125 3525 17155
rect 3555 17125 3560 17155
rect 3520 16995 3560 17125
rect 3520 16965 3525 16995
rect 3555 16965 3560 16995
rect 3520 16960 3560 16965
rect 3600 17155 3640 17160
rect 3600 17125 3605 17155
rect 3635 17125 3640 17155
rect 3600 16995 3640 17125
rect 3600 16965 3605 16995
rect 3635 16965 3640 16995
rect 3600 16960 3640 16965
rect 3680 17155 3720 17160
rect 3680 17125 3685 17155
rect 3715 17125 3720 17155
rect 3680 16995 3720 17125
rect 3680 16965 3685 16995
rect 3715 16965 3720 16995
rect 3680 16960 3720 16965
rect 3760 17155 3800 17160
rect 3760 17125 3765 17155
rect 3795 17125 3800 17155
rect 3760 16995 3800 17125
rect 3760 16965 3765 16995
rect 3795 16965 3800 16995
rect 3760 16960 3800 16965
rect 3840 17155 3880 17160
rect 3840 17125 3845 17155
rect 3875 17125 3880 17155
rect 3840 16995 3880 17125
rect 3840 16965 3845 16995
rect 3875 16965 3880 16995
rect 3840 16960 3880 16965
rect 3920 17155 3960 17160
rect 3920 17125 3925 17155
rect 3955 17125 3960 17155
rect 3920 16995 3960 17125
rect 3920 16965 3925 16995
rect 3955 16965 3960 16995
rect 3920 16960 3960 16965
rect 4000 17155 4040 17160
rect 4000 17125 4005 17155
rect 4035 17125 4040 17155
rect 4000 16995 4040 17125
rect 4000 16965 4005 16995
rect 4035 16965 4040 16995
rect 4000 16960 4040 16965
rect 4080 17155 4120 17160
rect 4080 17125 4085 17155
rect 4115 17125 4120 17155
rect 4080 16995 4120 17125
rect 4080 16965 4085 16995
rect 4115 16965 4120 16995
rect 4080 16960 4120 16965
rect 4160 17155 4200 17160
rect 4160 17125 4165 17155
rect 4195 17125 4200 17155
rect 4160 16995 4200 17125
rect 4160 16965 4165 16995
rect 4195 16965 4200 16995
rect 4160 16960 4200 16965
rect 0 16915 40 16920
rect 0 16885 5 16915
rect 35 16885 40 16915
rect 0 16755 40 16885
rect 0 16725 5 16755
rect 35 16725 40 16755
rect 0 16720 40 16725
rect 80 16915 120 16920
rect 80 16885 85 16915
rect 115 16885 120 16915
rect 80 16755 120 16885
rect 80 16725 85 16755
rect 115 16725 120 16755
rect 80 16720 120 16725
rect 160 16915 200 16920
rect 160 16885 165 16915
rect 195 16885 200 16915
rect 160 16755 200 16885
rect 160 16725 165 16755
rect 195 16725 200 16755
rect 160 16720 200 16725
rect 240 16915 280 16920
rect 240 16885 245 16915
rect 275 16885 280 16915
rect 240 16755 280 16885
rect 240 16725 245 16755
rect 275 16725 280 16755
rect 240 16720 280 16725
rect 320 16915 360 16920
rect 320 16885 325 16915
rect 355 16885 360 16915
rect 320 16755 360 16885
rect 320 16725 325 16755
rect 355 16725 360 16755
rect 320 16720 360 16725
rect 400 16915 440 16920
rect 400 16885 405 16915
rect 435 16885 440 16915
rect 400 16755 440 16885
rect 400 16725 405 16755
rect 435 16725 440 16755
rect 400 16720 440 16725
rect 480 16915 520 16920
rect 480 16885 485 16915
rect 515 16885 520 16915
rect 480 16755 520 16885
rect 480 16725 485 16755
rect 515 16725 520 16755
rect 480 16720 520 16725
rect 560 16915 600 16920
rect 560 16885 565 16915
rect 595 16885 600 16915
rect 560 16755 600 16885
rect 560 16725 565 16755
rect 595 16725 600 16755
rect 560 16720 600 16725
rect 640 16915 680 16920
rect 640 16885 645 16915
rect 675 16885 680 16915
rect 640 16755 680 16885
rect 640 16725 645 16755
rect 675 16725 680 16755
rect 640 16720 680 16725
rect 720 16915 760 16920
rect 720 16885 725 16915
rect 755 16885 760 16915
rect 720 16755 760 16885
rect 720 16725 725 16755
rect 755 16725 760 16755
rect 720 16720 760 16725
rect 800 16915 840 16920
rect 800 16885 805 16915
rect 835 16885 840 16915
rect 800 16755 840 16885
rect 800 16725 805 16755
rect 835 16725 840 16755
rect 800 16720 840 16725
rect 880 16915 920 16920
rect 880 16885 885 16915
rect 915 16885 920 16915
rect 880 16755 920 16885
rect 880 16725 885 16755
rect 915 16725 920 16755
rect 880 16720 920 16725
rect 960 16915 1000 16920
rect 960 16885 965 16915
rect 995 16885 1000 16915
rect 960 16755 1000 16885
rect 960 16725 965 16755
rect 995 16725 1000 16755
rect 960 16720 1000 16725
rect 1040 16915 1080 16920
rect 1040 16885 1045 16915
rect 1075 16885 1080 16915
rect 1040 16755 1080 16885
rect 1040 16725 1045 16755
rect 1075 16725 1080 16755
rect 1040 16720 1080 16725
rect 1120 16915 1160 16920
rect 1120 16885 1125 16915
rect 1155 16885 1160 16915
rect 1120 16755 1160 16885
rect 1120 16725 1125 16755
rect 1155 16725 1160 16755
rect 1120 16720 1160 16725
rect 1200 16915 1240 16920
rect 1200 16885 1205 16915
rect 1235 16885 1240 16915
rect 1200 16755 1240 16885
rect 1200 16725 1205 16755
rect 1235 16725 1240 16755
rect 1200 16720 1240 16725
rect 1280 16915 1320 16920
rect 1280 16885 1285 16915
rect 1315 16885 1320 16915
rect 1280 16755 1320 16885
rect 1280 16725 1285 16755
rect 1315 16725 1320 16755
rect 1280 16720 1320 16725
rect 1360 16915 1400 16920
rect 1360 16885 1365 16915
rect 1395 16885 1400 16915
rect 1360 16755 1400 16885
rect 1360 16725 1365 16755
rect 1395 16725 1400 16755
rect 1360 16720 1400 16725
rect 1440 16915 1480 16920
rect 1440 16885 1445 16915
rect 1475 16885 1480 16915
rect 1440 16755 1480 16885
rect 1440 16725 1445 16755
rect 1475 16725 1480 16755
rect 1440 16720 1480 16725
rect 1520 16915 1560 16920
rect 1520 16885 1525 16915
rect 1555 16885 1560 16915
rect 1520 16755 1560 16885
rect 1520 16725 1525 16755
rect 1555 16725 1560 16755
rect 1520 16720 1560 16725
rect 1600 16915 1640 16920
rect 1600 16885 1605 16915
rect 1635 16885 1640 16915
rect 1600 16755 1640 16885
rect 1600 16725 1605 16755
rect 1635 16725 1640 16755
rect 1600 16720 1640 16725
rect 1680 16915 1720 16920
rect 1680 16885 1685 16915
rect 1715 16885 1720 16915
rect 1680 16755 1720 16885
rect 1680 16725 1685 16755
rect 1715 16725 1720 16755
rect 1680 16720 1720 16725
rect 1760 16915 1800 16920
rect 1760 16885 1765 16915
rect 1795 16885 1800 16915
rect 1760 16755 1800 16885
rect 1760 16725 1765 16755
rect 1795 16725 1800 16755
rect 1760 16720 1800 16725
rect 1840 16915 1880 16920
rect 1840 16885 1845 16915
rect 1875 16885 1880 16915
rect 1840 16755 1880 16885
rect 1840 16725 1845 16755
rect 1875 16725 1880 16755
rect 1840 16720 1880 16725
rect 1920 16915 1960 16920
rect 1920 16885 1925 16915
rect 1955 16885 1960 16915
rect 1920 16755 1960 16885
rect 1920 16725 1925 16755
rect 1955 16725 1960 16755
rect 1920 16720 1960 16725
rect 2000 16915 2040 16920
rect 2000 16885 2005 16915
rect 2035 16885 2040 16915
rect 2000 16755 2040 16885
rect 2000 16725 2005 16755
rect 2035 16725 2040 16755
rect 2000 16720 2040 16725
rect 2080 16915 2120 16920
rect 2080 16885 2085 16915
rect 2115 16885 2120 16915
rect 2080 16755 2120 16885
rect 2080 16725 2085 16755
rect 2115 16725 2120 16755
rect 2080 16720 2120 16725
rect 2160 16915 2200 16920
rect 2160 16885 2165 16915
rect 2195 16885 2200 16915
rect 2160 16755 2200 16885
rect 2160 16725 2165 16755
rect 2195 16725 2200 16755
rect 2160 16720 2200 16725
rect 2240 16915 2280 16920
rect 2240 16885 2245 16915
rect 2275 16885 2280 16915
rect 2240 16755 2280 16885
rect 2240 16725 2245 16755
rect 2275 16725 2280 16755
rect 2240 16720 2280 16725
rect 2320 16915 2360 16920
rect 2320 16885 2325 16915
rect 2355 16885 2360 16915
rect 2320 16755 2360 16885
rect 2320 16725 2325 16755
rect 2355 16725 2360 16755
rect 2320 16720 2360 16725
rect 2400 16915 2440 16920
rect 2400 16885 2405 16915
rect 2435 16885 2440 16915
rect 2400 16755 2440 16885
rect 2400 16725 2405 16755
rect 2435 16725 2440 16755
rect 2400 16720 2440 16725
rect 2480 16915 2520 16920
rect 2480 16885 2485 16915
rect 2515 16885 2520 16915
rect 2480 16755 2520 16885
rect 2480 16725 2485 16755
rect 2515 16725 2520 16755
rect 2480 16720 2520 16725
rect 2560 16915 2600 16920
rect 2560 16885 2565 16915
rect 2595 16885 2600 16915
rect 2560 16755 2600 16885
rect 2560 16725 2565 16755
rect 2595 16725 2600 16755
rect 2560 16720 2600 16725
rect 2640 16915 2680 16920
rect 2640 16885 2645 16915
rect 2675 16885 2680 16915
rect 2640 16755 2680 16885
rect 2640 16725 2645 16755
rect 2675 16725 2680 16755
rect 2640 16720 2680 16725
rect 2720 16915 2760 16920
rect 2720 16885 2725 16915
rect 2755 16885 2760 16915
rect 2720 16755 2760 16885
rect 2720 16725 2725 16755
rect 2755 16725 2760 16755
rect 2720 16720 2760 16725
rect 2800 16915 2840 16920
rect 2800 16885 2805 16915
rect 2835 16885 2840 16915
rect 2800 16755 2840 16885
rect 2800 16725 2805 16755
rect 2835 16725 2840 16755
rect 2800 16720 2840 16725
rect 2880 16915 2920 16920
rect 2880 16885 2885 16915
rect 2915 16885 2920 16915
rect 2880 16755 2920 16885
rect 2880 16725 2885 16755
rect 2915 16725 2920 16755
rect 2880 16720 2920 16725
rect 2960 16915 3000 16920
rect 2960 16885 2965 16915
rect 2995 16885 3000 16915
rect 2960 16755 3000 16885
rect 2960 16725 2965 16755
rect 2995 16725 3000 16755
rect 2960 16720 3000 16725
rect 3040 16915 3080 16920
rect 3040 16885 3045 16915
rect 3075 16885 3080 16915
rect 3040 16755 3080 16885
rect 3040 16725 3045 16755
rect 3075 16725 3080 16755
rect 3040 16720 3080 16725
rect 3120 16915 3160 16920
rect 3120 16885 3125 16915
rect 3155 16885 3160 16915
rect 3120 16755 3160 16885
rect 3120 16725 3125 16755
rect 3155 16725 3160 16755
rect 3120 16720 3160 16725
rect 3200 16915 3240 16920
rect 3200 16885 3205 16915
rect 3235 16885 3240 16915
rect 3200 16755 3240 16885
rect 3200 16725 3205 16755
rect 3235 16725 3240 16755
rect 3200 16720 3240 16725
rect 3280 16915 3320 16920
rect 3280 16885 3285 16915
rect 3315 16885 3320 16915
rect 3280 16755 3320 16885
rect 3280 16725 3285 16755
rect 3315 16725 3320 16755
rect 3280 16720 3320 16725
rect 3360 16915 3400 16920
rect 3360 16885 3365 16915
rect 3395 16885 3400 16915
rect 3360 16755 3400 16885
rect 3360 16725 3365 16755
rect 3395 16725 3400 16755
rect 3360 16720 3400 16725
rect 3440 16915 3480 16920
rect 3440 16885 3445 16915
rect 3475 16885 3480 16915
rect 3440 16755 3480 16885
rect 3440 16725 3445 16755
rect 3475 16725 3480 16755
rect 3440 16720 3480 16725
rect 3520 16915 3560 16920
rect 3520 16885 3525 16915
rect 3555 16885 3560 16915
rect 3520 16755 3560 16885
rect 3520 16725 3525 16755
rect 3555 16725 3560 16755
rect 3520 16720 3560 16725
rect 3600 16915 3640 16920
rect 3600 16885 3605 16915
rect 3635 16885 3640 16915
rect 3600 16755 3640 16885
rect 3600 16725 3605 16755
rect 3635 16725 3640 16755
rect 3600 16720 3640 16725
rect 3680 16915 3720 16920
rect 3680 16885 3685 16915
rect 3715 16885 3720 16915
rect 3680 16755 3720 16885
rect 3680 16725 3685 16755
rect 3715 16725 3720 16755
rect 3680 16720 3720 16725
rect 3760 16915 3800 16920
rect 3760 16885 3765 16915
rect 3795 16885 3800 16915
rect 3760 16755 3800 16885
rect 3760 16725 3765 16755
rect 3795 16725 3800 16755
rect 3760 16720 3800 16725
rect 3840 16915 3880 16920
rect 3840 16885 3845 16915
rect 3875 16885 3880 16915
rect 3840 16755 3880 16885
rect 3840 16725 3845 16755
rect 3875 16725 3880 16755
rect 3840 16720 3880 16725
rect 3920 16915 3960 16920
rect 3920 16885 3925 16915
rect 3955 16885 3960 16915
rect 3920 16755 3960 16885
rect 3920 16725 3925 16755
rect 3955 16725 3960 16755
rect 3920 16720 3960 16725
rect 4000 16915 4040 16920
rect 4000 16885 4005 16915
rect 4035 16885 4040 16915
rect 4000 16755 4040 16885
rect 4000 16725 4005 16755
rect 4035 16725 4040 16755
rect 4000 16720 4040 16725
rect 4080 16915 4120 16920
rect 4080 16885 4085 16915
rect 4115 16885 4120 16915
rect 4080 16755 4120 16885
rect 4080 16725 4085 16755
rect 4115 16725 4120 16755
rect 4080 16720 4120 16725
rect 4160 16915 4200 16920
rect 4160 16885 4165 16915
rect 4195 16885 4200 16915
rect 4160 16755 4200 16885
rect 4160 16725 4165 16755
rect 4195 16725 4200 16755
rect 4160 16720 4200 16725
rect 4240 16720 4280 18485
rect 4320 18595 4360 18720
rect 4320 18565 4325 18595
rect 4355 18565 4360 18595
rect 4320 16720 4360 18565
rect 4400 18675 4440 18720
rect 4400 18645 4405 18675
rect 4435 18645 4440 18675
rect 4400 18515 4440 18645
rect 4400 18485 4405 18515
rect 4435 18485 4440 18515
rect 4400 16720 4440 18485
rect 4480 18435 4520 18720
rect 4480 18405 4485 18435
rect 4515 18405 4520 18435
rect 4480 18275 4520 18405
rect 4480 18245 4485 18275
rect 4515 18245 4520 18275
rect 4480 16720 4520 18245
rect 4560 18355 4600 18720
rect 4560 18325 4565 18355
rect 4595 18325 4600 18355
rect 4560 16720 4600 18325
rect 4640 18435 4680 18720
rect 4640 18405 4645 18435
rect 4675 18405 4680 18435
rect 4640 18275 4680 18405
rect 4640 18245 4645 18275
rect 4675 18245 4680 18275
rect 4640 16720 4680 18245
rect 4720 18195 4760 18720
rect 4720 18165 4725 18195
rect 4755 18165 4760 18195
rect 4720 18035 4760 18165
rect 4720 18005 4725 18035
rect 4755 18005 4760 18035
rect 4720 17875 4760 18005
rect 4720 17845 4725 17875
rect 4755 17845 4760 17875
rect 4720 17715 4760 17845
rect 4720 17685 4725 17715
rect 4755 17685 4760 17715
rect 4720 17555 4760 17685
rect 4720 17525 4725 17555
rect 4755 17525 4760 17555
rect 4720 17395 4760 17525
rect 4720 17365 4725 17395
rect 4755 17365 4760 17395
rect 4720 17235 4760 17365
rect 4720 17205 4725 17235
rect 4755 17205 4760 17235
rect 4720 16720 4760 17205
rect 4800 18115 4840 18720
rect 4800 18085 4805 18115
rect 4835 18085 4840 18115
rect 4800 16720 4840 18085
rect 4880 18195 4920 18720
rect 4880 18165 4885 18195
rect 4915 18165 4920 18195
rect 4880 18035 4920 18165
rect 4880 18005 4885 18035
rect 4915 18005 4920 18035
rect 4880 17875 4920 18005
rect 4880 17845 4885 17875
rect 4915 17845 4920 17875
rect 4880 17715 4920 17845
rect 4880 17685 4885 17715
rect 4915 17685 4920 17715
rect 4880 17555 4920 17685
rect 4880 17525 4885 17555
rect 4915 17525 4920 17555
rect 4880 17395 4920 17525
rect 4880 17365 4885 17395
rect 4915 17365 4920 17395
rect 4880 17235 4920 17365
rect 4880 17205 4885 17235
rect 4915 17205 4920 17235
rect 4880 16720 4920 17205
rect 4960 17955 5000 18720
rect 4960 17925 4965 17955
rect 4995 17925 5000 17955
rect 4960 16720 5000 17925
rect 5040 18195 5080 18720
rect 5040 18165 5045 18195
rect 5075 18165 5080 18195
rect 5040 18035 5080 18165
rect 5040 18005 5045 18035
rect 5075 18005 5080 18035
rect 5040 17875 5080 18005
rect 5040 17845 5045 17875
rect 5075 17845 5080 17875
rect 5040 17715 5080 17845
rect 5040 17685 5045 17715
rect 5075 17685 5080 17715
rect 5040 17555 5080 17685
rect 5040 17525 5045 17555
rect 5075 17525 5080 17555
rect 5040 17395 5080 17525
rect 5040 17365 5045 17395
rect 5075 17365 5080 17395
rect 5040 17235 5080 17365
rect 5040 17205 5045 17235
rect 5075 17205 5080 17235
rect 5040 16720 5080 17205
rect 5120 17795 5160 18720
rect 5120 17765 5125 17795
rect 5155 17765 5160 17795
rect 5120 16720 5160 17765
rect 5200 18195 5240 18720
rect 5200 18165 5205 18195
rect 5235 18165 5240 18195
rect 5200 18035 5240 18165
rect 5200 18005 5205 18035
rect 5235 18005 5240 18035
rect 5200 17875 5240 18005
rect 5200 17845 5205 17875
rect 5235 17845 5240 17875
rect 5200 17715 5240 17845
rect 5200 17685 5205 17715
rect 5235 17685 5240 17715
rect 5200 17555 5240 17685
rect 5200 17525 5205 17555
rect 5235 17525 5240 17555
rect 5200 17395 5240 17525
rect 5200 17365 5205 17395
rect 5235 17365 5240 17395
rect 5200 17235 5240 17365
rect 5200 17205 5205 17235
rect 5235 17205 5240 17235
rect 5200 16720 5240 17205
rect 5280 17635 5320 18720
rect 5280 17605 5285 17635
rect 5315 17605 5320 17635
rect 5280 16720 5320 17605
rect 5360 18195 5400 18720
rect 5360 18165 5365 18195
rect 5395 18165 5400 18195
rect 5360 18035 5400 18165
rect 5360 18005 5365 18035
rect 5395 18005 5400 18035
rect 5360 17875 5400 18005
rect 5360 17845 5365 17875
rect 5395 17845 5400 17875
rect 5360 17715 5400 17845
rect 5360 17685 5365 17715
rect 5395 17685 5400 17715
rect 5360 17555 5400 17685
rect 5360 17525 5365 17555
rect 5395 17525 5400 17555
rect 5360 17395 5400 17525
rect 5360 17365 5365 17395
rect 5395 17365 5400 17395
rect 5360 17235 5400 17365
rect 5360 17205 5365 17235
rect 5395 17205 5400 17235
rect 5360 16720 5400 17205
rect 5440 17475 5480 18720
rect 5440 17445 5445 17475
rect 5475 17445 5480 17475
rect 5440 16720 5480 17445
rect 5520 18195 5560 18720
rect 5520 18165 5525 18195
rect 5555 18165 5560 18195
rect 5520 18035 5560 18165
rect 5520 18005 5525 18035
rect 5555 18005 5560 18035
rect 5520 17875 5560 18005
rect 5520 17845 5525 17875
rect 5555 17845 5560 17875
rect 5520 17715 5560 17845
rect 5520 17685 5525 17715
rect 5555 17685 5560 17715
rect 5520 17555 5560 17685
rect 5520 17525 5525 17555
rect 5555 17525 5560 17555
rect 5520 17395 5560 17525
rect 5520 17365 5525 17395
rect 5555 17365 5560 17395
rect 5520 17235 5560 17365
rect 5520 17205 5525 17235
rect 5555 17205 5560 17235
rect 5520 16720 5560 17205
rect 5600 17315 5640 18720
rect 5600 17285 5605 17315
rect 5635 17285 5640 17315
rect 5600 16720 5640 17285
rect 5680 18195 5720 18720
rect 5680 18165 5685 18195
rect 5715 18165 5720 18195
rect 5680 18035 5720 18165
rect 5680 18005 5685 18035
rect 5715 18005 5720 18035
rect 5680 17875 5720 18005
rect 5680 17845 5685 17875
rect 5715 17845 5720 17875
rect 5680 17715 5720 17845
rect 5680 17685 5685 17715
rect 5715 17685 5720 17715
rect 5680 17555 5720 17685
rect 5680 17525 5685 17555
rect 5715 17525 5720 17555
rect 5680 17395 5720 17525
rect 5680 17365 5685 17395
rect 5715 17365 5720 17395
rect 5680 17235 5720 17365
rect 5680 17205 5685 17235
rect 5715 17205 5720 17235
rect 5680 16720 5720 17205
rect 5760 17155 5800 18720
rect 5760 17125 5765 17155
rect 5795 17125 5800 17155
rect 5760 16995 5800 17125
rect 5760 16965 5765 16995
rect 5795 16965 5800 16995
rect 5760 16720 5800 16965
rect 5840 17075 5880 18720
rect 5840 17045 5845 17075
rect 5875 17045 5880 17075
rect 5840 16720 5880 17045
rect 5920 17155 5960 18720
rect 5920 17125 5925 17155
rect 5955 17125 5960 17155
rect 5920 16995 5960 17125
rect 5920 16965 5925 16995
rect 5955 16965 5960 16995
rect 5920 16720 5960 16965
rect 6000 16915 6040 18720
rect 6000 16885 6005 16915
rect 6035 16885 6040 16915
rect 6000 16755 6040 16885
rect 6000 16725 6005 16755
rect 6035 16725 6040 16755
rect 6000 16720 6040 16725
rect 6080 16835 6120 18720
rect 6080 16805 6085 16835
rect 6115 16805 6120 16835
rect 6080 16720 6120 16805
rect 6160 16915 6200 18720
rect 6240 18675 6280 18680
rect 6240 18645 6245 18675
rect 6275 18645 6280 18675
rect 6240 18515 6280 18645
rect 6240 18485 6245 18515
rect 6275 18485 6280 18515
rect 6240 18480 6280 18485
rect 6320 18675 6360 18680
rect 6320 18645 6325 18675
rect 6355 18645 6360 18675
rect 6320 18515 6360 18645
rect 6320 18485 6325 18515
rect 6355 18485 6360 18515
rect 6320 18480 6360 18485
rect 6400 18675 6440 18680
rect 6400 18645 6405 18675
rect 6435 18645 6440 18675
rect 6400 18515 6440 18645
rect 6400 18485 6405 18515
rect 6435 18485 6440 18515
rect 6400 18480 6440 18485
rect 6480 18675 6520 18680
rect 6480 18645 6485 18675
rect 6515 18645 6520 18675
rect 6480 18515 6520 18645
rect 6480 18485 6485 18515
rect 6515 18485 6520 18515
rect 6480 18480 6520 18485
rect 6560 18675 6600 18680
rect 6560 18645 6565 18675
rect 6595 18645 6600 18675
rect 6560 18515 6600 18645
rect 6560 18485 6565 18515
rect 6595 18485 6600 18515
rect 6560 18480 6600 18485
rect 6640 18675 6680 18680
rect 6640 18645 6645 18675
rect 6675 18645 6680 18675
rect 6640 18515 6680 18645
rect 6640 18485 6645 18515
rect 6675 18485 6680 18515
rect 6640 18480 6680 18485
rect 6720 18675 6760 18680
rect 6720 18645 6725 18675
rect 6755 18645 6760 18675
rect 6720 18515 6760 18645
rect 6720 18485 6725 18515
rect 6755 18485 6760 18515
rect 6720 18480 6760 18485
rect 6800 18675 6840 18680
rect 6800 18645 6805 18675
rect 6835 18645 6840 18675
rect 6800 18515 6840 18645
rect 6800 18485 6805 18515
rect 6835 18485 6840 18515
rect 6800 18480 6840 18485
rect 6880 18675 6920 18680
rect 6880 18645 6885 18675
rect 6915 18645 6920 18675
rect 6880 18515 6920 18645
rect 6880 18485 6885 18515
rect 6915 18485 6920 18515
rect 6880 18480 6920 18485
rect 6960 18675 7000 18680
rect 6960 18645 6965 18675
rect 6995 18645 7000 18675
rect 6960 18515 7000 18645
rect 6960 18485 6965 18515
rect 6995 18485 7000 18515
rect 6960 18480 7000 18485
rect 7040 18675 7080 18680
rect 7040 18645 7045 18675
rect 7075 18645 7080 18675
rect 7040 18515 7080 18645
rect 7040 18485 7045 18515
rect 7075 18485 7080 18515
rect 7040 18480 7080 18485
rect 7120 18675 7160 18680
rect 7120 18645 7125 18675
rect 7155 18645 7160 18675
rect 7120 18515 7160 18645
rect 7120 18485 7125 18515
rect 7155 18485 7160 18515
rect 7120 18480 7160 18485
rect 7200 18675 7240 18680
rect 7200 18645 7205 18675
rect 7235 18645 7240 18675
rect 7200 18515 7240 18645
rect 7200 18485 7205 18515
rect 7235 18485 7240 18515
rect 7200 18480 7240 18485
rect 7280 18675 7320 18680
rect 7280 18645 7285 18675
rect 7315 18645 7320 18675
rect 7280 18515 7320 18645
rect 7280 18485 7285 18515
rect 7315 18485 7320 18515
rect 7280 18480 7320 18485
rect 7360 18675 7400 18680
rect 7360 18645 7365 18675
rect 7395 18645 7400 18675
rect 7360 18515 7400 18645
rect 7360 18485 7365 18515
rect 7395 18485 7400 18515
rect 7360 18480 7400 18485
rect 7440 18675 7480 18680
rect 7440 18645 7445 18675
rect 7475 18645 7480 18675
rect 7440 18515 7480 18645
rect 7440 18485 7445 18515
rect 7475 18485 7480 18515
rect 7440 18480 7480 18485
rect 7520 18675 7560 18680
rect 7520 18645 7525 18675
rect 7555 18645 7560 18675
rect 7520 18515 7560 18645
rect 7520 18485 7525 18515
rect 7555 18485 7560 18515
rect 7520 18480 7560 18485
rect 7600 18675 7640 18680
rect 7600 18645 7605 18675
rect 7635 18645 7640 18675
rect 7600 18515 7640 18645
rect 7600 18485 7605 18515
rect 7635 18485 7640 18515
rect 7600 18480 7640 18485
rect 7680 18675 7720 18680
rect 7680 18645 7685 18675
rect 7715 18645 7720 18675
rect 7680 18515 7720 18645
rect 7680 18485 7685 18515
rect 7715 18485 7720 18515
rect 7680 18480 7720 18485
rect 7760 18675 7800 18680
rect 7760 18645 7765 18675
rect 7795 18645 7800 18675
rect 7760 18515 7800 18645
rect 7760 18485 7765 18515
rect 7795 18485 7800 18515
rect 7760 18480 7800 18485
rect 7840 18675 7880 18680
rect 7840 18645 7845 18675
rect 7875 18645 7880 18675
rect 7840 18515 7880 18645
rect 7840 18485 7845 18515
rect 7875 18485 7880 18515
rect 7840 18480 7880 18485
rect 7920 18675 7960 18680
rect 7920 18645 7925 18675
rect 7955 18645 7960 18675
rect 7920 18515 7960 18645
rect 7920 18485 7925 18515
rect 7955 18485 7960 18515
rect 7920 18480 7960 18485
rect 8000 18675 8040 18680
rect 8000 18645 8005 18675
rect 8035 18645 8040 18675
rect 8000 18515 8040 18645
rect 8000 18485 8005 18515
rect 8035 18485 8040 18515
rect 8000 18480 8040 18485
rect 8080 18675 8120 18680
rect 8080 18645 8085 18675
rect 8115 18645 8120 18675
rect 8080 18515 8120 18645
rect 8080 18485 8085 18515
rect 8115 18485 8120 18515
rect 8080 18480 8120 18485
rect 8160 18675 8200 18680
rect 8160 18645 8165 18675
rect 8195 18645 8200 18675
rect 8160 18515 8200 18645
rect 8160 18485 8165 18515
rect 8195 18485 8200 18515
rect 8160 18480 8200 18485
rect 8240 18675 8280 18680
rect 8240 18645 8245 18675
rect 8275 18645 8280 18675
rect 8240 18515 8280 18645
rect 8240 18485 8245 18515
rect 8275 18485 8280 18515
rect 8240 18480 8280 18485
rect 8320 18675 8360 18680
rect 8320 18645 8325 18675
rect 8355 18645 8360 18675
rect 8320 18515 8360 18645
rect 8320 18485 8325 18515
rect 8355 18485 8360 18515
rect 8320 18480 8360 18485
rect 8400 18675 8440 18680
rect 8400 18645 8405 18675
rect 8435 18645 8440 18675
rect 8400 18515 8440 18645
rect 8400 18485 8405 18515
rect 8435 18485 8440 18515
rect 8400 18480 8440 18485
rect 8480 18675 8520 18680
rect 8480 18645 8485 18675
rect 8515 18645 8520 18675
rect 8480 18515 8520 18645
rect 8480 18485 8485 18515
rect 8515 18485 8520 18515
rect 8480 18480 8520 18485
rect 8560 18675 8600 18680
rect 8560 18645 8565 18675
rect 8595 18645 8600 18675
rect 8560 18515 8600 18645
rect 8560 18485 8565 18515
rect 8595 18485 8600 18515
rect 8560 18480 8600 18485
rect 8640 18675 8680 18680
rect 8640 18645 8645 18675
rect 8675 18645 8680 18675
rect 8640 18515 8680 18645
rect 8640 18485 8645 18515
rect 8675 18485 8680 18515
rect 8640 18480 8680 18485
rect 8720 18675 8760 18680
rect 8720 18645 8725 18675
rect 8755 18645 8760 18675
rect 8720 18515 8760 18645
rect 8720 18485 8725 18515
rect 8755 18485 8760 18515
rect 8720 18480 8760 18485
rect 8800 18675 8840 18680
rect 8800 18645 8805 18675
rect 8835 18645 8840 18675
rect 8800 18515 8840 18645
rect 8800 18485 8805 18515
rect 8835 18485 8840 18515
rect 8800 18480 8840 18485
rect 8880 18675 8920 18680
rect 8880 18645 8885 18675
rect 8915 18645 8920 18675
rect 8880 18515 8920 18645
rect 8880 18485 8885 18515
rect 8915 18485 8920 18515
rect 8880 18480 8920 18485
rect 8960 18675 9000 18680
rect 8960 18645 8965 18675
rect 8995 18645 9000 18675
rect 8960 18515 9000 18645
rect 8960 18485 8965 18515
rect 8995 18485 9000 18515
rect 8960 18480 9000 18485
rect 9040 18675 9080 18680
rect 9040 18645 9045 18675
rect 9075 18645 9080 18675
rect 9040 18515 9080 18645
rect 9040 18485 9045 18515
rect 9075 18485 9080 18515
rect 9040 18480 9080 18485
rect 9120 18675 9160 18680
rect 9120 18645 9125 18675
rect 9155 18645 9160 18675
rect 9120 18515 9160 18645
rect 9120 18485 9125 18515
rect 9155 18485 9160 18515
rect 9120 18480 9160 18485
rect 9200 18675 9240 18680
rect 9200 18645 9205 18675
rect 9235 18645 9240 18675
rect 9200 18515 9240 18645
rect 9200 18485 9205 18515
rect 9235 18485 9240 18515
rect 9200 18480 9240 18485
rect 9280 18675 9320 18680
rect 9280 18645 9285 18675
rect 9315 18645 9320 18675
rect 9280 18515 9320 18645
rect 9280 18485 9285 18515
rect 9315 18485 9320 18515
rect 9280 18480 9320 18485
rect 9360 18675 9400 18680
rect 9360 18645 9365 18675
rect 9395 18645 9400 18675
rect 9360 18515 9400 18645
rect 9360 18485 9365 18515
rect 9395 18485 9400 18515
rect 9360 18480 9400 18485
rect 9440 18675 9480 18680
rect 9440 18645 9445 18675
rect 9475 18645 9480 18675
rect 9440 18515 9480 18645
rect 9440 18485 9445 18515
rect 9475 18485 9480 18515
rect 9440 18480 9480 18485
rect 6240 18435 6280 18440
rect 6240 18405 6245 18435
rect 6275 18405 6280 18435
rect 6240 18275 6280 18405
rect 6240 18245 6245 18275
rect 6275 18245 6280 18275
rect 6240 18240 6280 18245
rect 6320 18435 6360 18440
rect 6320 18405 6325 18435
rect 6355 18405 6360 18435
rect 6320 18275 6360 18405
rect 6320 18245 6325 18275
rect 6355 18245 6360 18275
rect 6320 18240 6360 18245
rect 6400 18435 6440 18440
rect 6400 18405 6405 18435
rect 6435 18405 6440 18435
rect 6400 18275 6440 18405
rect 6400 18245 6405 18275
rect 6435 18245 6440 18275
rect 6400 18240 6440 18245
rect 6480 18435 6520 18440
rect 6480 18405 6485 18435
rect 6515 18405 6520 18435
rect 6480 18275 6520 18405
rect 6480 18245 6485 18275
rect 6515 18245 6520 18275
rect 6480 18240 6520 18245
rect 6560 18435 6600 18440
rect 6560 18405 6565 18435
rect 6595 18405 6600 18435
rect 6560 18275 6600 18405
rect 6560 18245 6565 18275
rect 6595 18245 6600 18275
rect 6560 18240 6600 18245
rect 6640 18435 6680 18440
rect 6640 18405 6645 18435
rect 6675 18405 6680 18435
rect 6640 18275 6680 18405
rect 6640 18245 6645 18275
rect 6675 18245 6680 18275
rect 6640 18240 6680 18245
rect 6720 18435 6760 18440
rect 6720 18405 6725 18435
rect 6755 18405 6760 18435
rect 6720 18275 6760 18405
rect 6720 18245 6725 18275
rect 6755 18245 6760 18275
rect 6720 18240 6760 18245
rect 6800 18435 6840 18440
rect 6800 18405 6805 18435
rect 6835 18405 6840 18435
rect 6800 18275 6840 18405
rect 6800 18245 6805 18275
rect 6835 18245 6840 18275
rect 6800 18240 6840 18245
rect 6880 18435 6920 18440
rect 6880 18405 6885 18435
rect 6915 18405 6920 18435
rect 6880 18275 6920 18405
rect 6880 18245 6885 18275
rect 6915 18245 6920 18275
rect 6880 18240 6920 18245
rect 6960 18435 7000 18440
rect 6960 18405 6965 18435
rect 6995 18405 7000 18435
rect 6960 18275 7000 18405
rect 6960 18245 6965 18275
rect 6995 18245 7000 18275
rect 6960 18240 7000 18245
rect 7040 18435 7080 18440
rect 7040 18405 7045 18435
rect 7075 18405 7080 18435
rect 7040 18275 7080 18405
rect 7040 18245 7045 18275
rect 7075 18245 7080 18275
rect 7040 18240 7080 18245
rect 7120 18435 7160 18440
rect 7120 18405 7125 18435
rect 7155 18405 7160 18435
rect 7120 18275 7160 18405
rect 7120 18245 7125 18275
rect 7155 18245 7160 18275
rect 7120 18240 7160 18245
rect 7200 18435 7240 18440
rect 7200 18405 7205 18435
rect 7235 18405 7240 18435
rect 7200 18275 7240 18405
rect 7200 18245 7205 18275
rect 7235 18245 7240 18275
rect 7200 18240 7240 18245
rect 7280 18435 7320 18440
rect 7280 18405 7285 18435
rect 7315 18405 7320 18435
rect 7280 18275 7320 18405
rect 7280 18245 7285 18275
rect 7315 18245 7320 18275
rect 7280 18240 7320 18245
rect 7360 18435 7400 18440
rect 7360 18405 7365 18435
rect 7395 18405 7400 18435
rect 7360 18275 7400 18405
rect 7360 18245 7365 18275
rect 7395 18245 7400 18275
rect 7360 18240 7400 18245
rect 7440 18435 7480 18440
rect 7440 18405 7445 18435
rect 7475 18405 7480 18435
rect 7440 18275 7480 18405
rect 7440 18245 7445 18275
rect 7475 18245 7480 18275
rect 7440 18240 7480 18245
rect 7520 18435 7560 18440
rect 7520 18405 7525 18435
rect 7555 18405 7560 18435
rect 7520 18275 7560 18405
rect 7520 18245 7525 18275
rect 7555 18245 7560 18275
rect 7520 18240 7560 18245
rect 7600 18435 7640 18440
rect 7600 18405 7605 18435
rect 7635 18405 7640 18435
rect 7600 18275 7640 18405
rect 7600 18245 7605 18275
rect 7635 18245 7640 18275
rect 7600 18240 7640 18245
rect 7680 18435 7720 18440
rect 7680 18405 7685 18435
rect 7715 18405 7720 18435
rect 7680 18275 7720 18405
rect 7680 18245 7685 18275
rect 7715 18245 7720 18275
rect 7680 18240 7720 18245
rect 7760 18435 7800 18440
rect 7760 18405 7765 18435
rect 7795 18405 7800 18435
rect 7760 18275 7800 18405
rect 7760 18245 7765 18275
rect 7795 18245 7800 18275
rect 7760 18240 7800 18245
rect 7840 18435 7880 18440
rect 7840 18405 7845 18435
rect 7875 18405 7880 18435
rect 7840 18275 7880 18405
rect 7840 18245 7845 18275
rect 7875 18245 7880 18275
rect 7840 18240 7880 18245
rect 7920 18435 7960 18440
rect 7920 18405 7925 18435
rect 7955 18405 7960 18435
rect 7920 18275 7960 18405
rect 7920 18245 7925 18275
rect 7955 18245 7960 18275
rect 7920 18240 7960 18245
rect 8000 18435 8040 18440
rect 8000 18405 8005 18435
rect 8035 18405 8040 18435
rect 8000 18275 8040 18405
rect 8000 18245 8005 18275
rect 8035 18245 8040 18275
rect 8000 18240 8040 18245
rect 8080 18435 8120 18440
rect 8080 18405 8085 18435
rect 8115 18405 8120 18435
rect 8080 18275 8120 18405
rect 8080 18245 8085 18275
rect 8115 18245 8120 18275
rect 8080 18240 8120 18245
rect 8160 18435 8200 18440
rect 8160 18405 8165 18435
rect 8195 18405 8200 18435
rect 8160 18275 8200 18405
rect 8160 18245 8165 18275
rect 8195 18245 8200 18275
rect 8160 18240 8200 18245
rect 8240 18435 8280 18440
rect 8240 18405 8245 18435
rect 8275 18405 8280 18435
rect 8240 18275 8280 18405
rect 8240 18245 8245 18275
rect 8275 18245 8280 18275
rect 8240 18240 8280 18245
rect 8320 18435 8360 18440
rect 8320 18405 8325 18435
rect 8355 18405 8360 18435
rect 8320 18275 8360 18405
rect 8320 18245 8325 18275
rect 8355 18245 8360 18275
rect 8320 18240 8360 18245
rect 8400 18435 8440 18440
rect 8400 18405 8405 18435
rect 8435 18405 8440 18435
rect 8400 18275 8440 18405
rect 8400 18245 8405 18275
rect 8435 18245 8440 18275
rect 8400 18240 8440 18245
rect 8480 18435 8520 18440
rect 8480 18405 8485 18435
rect 8515 18405 8520 18435
rect 8480 18275 8520 18405
rect 8480 18245 8485 18275
rect 8515 18245 8520 18275
rect 8480 18240 8520 18245
rect 8560 18435 8600 18440
rect 8560 18405 8565 18435
rect 8595 18405 8600 18435
rect 8560 18275 8600 18405
rect 8560 18245 8565 18275
rect 8595 18245 8600 18275
rect 8560 18240 8600 18245
rect 8640 18435 8680 18440
rect 8640 18405 8645 18435
rect 8675 18405 8680 18435
rect 8640 18275 8680 18405
rect 8640 18245 8645 18275
rect 8675 18245 8680 18275
rect 8640 18240 8680 18245
rect 8720 18435 8760 18440
rect 8720 18405 8725 18435
rect 8755 18405 8760 18435
rect 8720 18275 8760 18405
rect 8720 18245 8725 18275
rect 8755 18245 8760 18275
rect 8720 18240 8760 18245
rect 8800 18435 8840 18440
rect 8800 18405 8805 18435
rect 8835 18405 8840 18435
rect 8800 18275 8840 18405
rect 8800 18245 8805 18275
rect 8835 18245 8840 18275
rect 8800 18240 8840 18245
rect 8880 18435 8920 18440
rect 8880 18405 8885 18435
rect 8915 18405 8920 18435
rect 8880 18275 8920 18405
rect 8880 18245 8885 18275
rect 8915 18245 8920 18275
rect 8880 18240 8920 18245
rect 8960 18435 9000 18440
rect 8960 18405 8965 18435
rect 8995 18405 9000 18435
rect 8960 18275 9000 18405
rect 8960 18245 8965 18275
rect 8995 18245 9000 18275
rect 8960 18240 9000 18245
rect 9040 18435 9080 18440
rect 9040 18405 9045 18435
rect 9075 18405 9080 18435
rect 9040 18275 9080 18405
rect 9040 18245 9045 18275
rect 9075 18245 9080 18275
rect 9040 18240 9080 18245
rect 9120 18435 9160 18440
rect 9120 18405 9125 18435
rect 9155 18405 9160 18435
rect 9120 18275 9160 18405
rect 9120 18245 9125 18275
rect 9155 18245 9160 18275
rect 9120 18240 9160 18245
rect 9200 18435 9240 18440
rect 9200 18405 9205 18435
rect 9235 18405 9240 18435
rect 9200 18275 9240 18405
rect 9200 18245 9205 18275
rect 9235 18245 9240 18275
rect 9200 18240 9240 18245
rect 9280 18435 9320 18440
rect 9280 18405 9285 18435
rect 9315 18405 9320 18435
rect 9280 18275 9320 18405
rect 9280 18245 9285 18275
rect 9315 18245 9320 18275
rect 9280 18240 9320 18245
rect 9360 18435 9400 18440
rect 9360 18405 9365 18435
rect 9395 18405 9400 18435
rect 9360 18275 9400 18405
rect 9360 18245 9365 18275
rect 9395 18245 9400 18275
rect 9360 18240 9400 18245
rect 9440 18435 9480 18440
rect 9440 18405 9445 18435
rect 9475 18405 9480 18435
rect 9440 18275 9480 18405
rect 9440 18245 9445 18275
rect 9475 18245 9480 18275
rect 9440 18240 9480 18245
rect 6240 18195 6280 18200
rect 6240 18165 6245 18195
rect 6275 18165 6280 18195
rect 6240 18035 6280 18165
rect 6240 18005 6245 18035
rect 6275 18005 6280 18035
rect 6240 17875 6280 18005
rect 6240 17845 6245 17875
rect 6275 17845 6280 17875
rect 6240 17715 6280 17845
rect 6240 17685 6245 17715
rect 6275 17685 6280 17715
rect 6240 17555 6280 17685
rect 6240 17525 6245 17555
rect 6275 17525 6280 17555
rect 6240 17395 6280 17525
rect 6240 17365 6245 17395
rect 6275 17365 6280 17395
rect 6240 17235 6280 17365
rect 6240 17205 6245 17235
rect 6275 17205 6280 17235
rect 6240 17200 6280 17205
rect 6320 18195 6360 18200
rect 6320 18165 6325 18195
rect 6355 18165 6360 18195
rect 6320 18035 6360 18165
rect 6320 18005 6325 18035
rect 6355 18005 6360 18035
rect 6320 17875 6360 18005
rect 6320 17845 6325 17875
rect 6355 17845 6360 17875
rect 6320 17715 6360 17845
rect 6320 17685 6325 17715
rect 6355 17685 6360 17715
rect 6320 17555 6360 17685
rect 6320 17525 6325 17555
rect 6355 17525 6360 17555
rect 6320 17395 6360 17525
rect 6320 17365 6325 17395
rect 6355 17365 6360 17395
rect 6320 17235 6360 17365
rect 6320 17205 6325 17235
rect 6355 17205 6360 17235
rect 6320 17200 6360 17205
rect 6400 18195 6440 18200
rect 6400 18165 6405 18195
rect 6435 18165 6440 18195
rect 6400 18035 6440 18165
rect 6400 18005 6405 18035
rect 6435 18005 6440 18035
rect 6400 17875 6440 18005
rect 6400 17845 6405 17875
rect 6435 17845 6440 17875
rect 6400 17715 6440 17845
rect 6400 17685 6405 17715
rect 6435 17685 6440 17715
rect 6400 17555 6440 17685
rect 6400 17525 6405 17555
rect 6435 17525 6440 17555
rect 6400 17395 6440 17525
rect 6400 17365 6405 17395
rect 6435 17365 6440 17395
rect 6400 17235 6440 17365
rect 6400 17205 6405 17235
rect 6435 17205 6440 17235
rect 6400 17200 6440 17205
rect 6480 18195 6520 18200
rect 6480 18165 6485 18195
rect 6515 18165 6520 18195
rect 6480 18035 6520 18165
rect 6480 18005 6485 18035
rect 6515 18005 6520 18035
rect 6480 17875 6520 18005
rect 6480 17845 6485 17875
rect 6515 17845 6520 17875
rect 6480 17715 6520 17845
rect 6480 17685 6485 17715
rect 6515 17685 6520 17715
rect 6480 17555 6520 17685
rect 6480 17525 6485 17555
rect 6515 17525 6520 17555
rect 6480 17395 6520 17525
rect 6480 17365 6485 17395
rect 6515 17365 6520 17395
rect 6480 17235 6520 17365
rect 6480 17205 6485 17235
rect 6515 17205 6520 17235
rect 6480 17200 6520 17205
rect 6560 18195 6600 18200
rect 6560 18165 6565 18195
rect 6595 18165 6600 18195
rect 6560 18035 6600 18165
rect 6560 18005 6565 18035
rect 6595 18005 6600 18035
rect 6560 17875 6600 18005
rect 6560 17845 6565 17875
rect 6595 17845 6600 17875
rect 6560 17715 6600 17845
rect 6560 17685 6565 17715
rect 6595 17685 6600 17715
rect 6560 17555 6600 17685
rect 6560 17525 6565 17555
rect 6595 17525 6600 17555
rect 6560 17395 6600 17525
rect 6560 17365 6565 17395
rect 6595 17365 6600 17395
rect 6560 17235 6600 17365
rect 6560 17205 6565 17235
rect 6595 17205 6600 17235
rect 6560 17200 6600 17205
rect 6640 18195 6680 18200
rect 6640 18165 6645 18195
rect 6675 18165 6680 18195
rect 6640 18035 6680 18165
rect 6640 18005 6645 18035
rect 6675 18005 6680 18035
rect 6640 17875 6680 18005
rect 6640 17845 6645 17875
rect 6675 17845 6680 17875
rect 6640 17715 6680 17845
rect 6640 17685 6645 17715
rect 6675 17685 6680 17715
rect 6640 17555 6680 17685
rect 6640 17525 6645 17555
rect 6675 17525 6680 17555
rect 6640 17395 6680 17525
rect 6640 17365 6645 17395
rect 6675 17365 6680 17395
rect 6640 17235 6680 17365
rect 6640 17205 6645 17235
rect 6675 17205 6680 17235
rect 6640 17200 6680 17205
rect 6720 18195 6760 18200
rect 6720 18165 6725 18195
rect 6755 18165 6760 18195
rect 6720 18035 6760 18165
rect 6720 18005 6725 18035
rect 6755 18005 6760 18035
rect 6720 17875 6760 18005
rect 6720 17845 6725 17875
rect 6755 17845 6760 17875
rect 6720 17715 6760 17845
rect 6720 17685 6725 17715
rect 6755 17685 6760 17715
rect 6720 17555 6760 17685
rect 6720 17525 6725 17555
rect 6755 17525 6760 17555
rect 6720 17395 6760 17525
rect 6720 17365 6725 17395
rect 6755 17365 6760 17395
rect 6720 17235 6760 17365
rect 6720 17205 6725 17235
rect 6755 17205 6760 17235
rect 6720 17200 6760 17205
rect 6800 18195 6840 18200
rect 6800 18165 6805 18195
rect 6835 18165 6840 18195
rect 6800 18035 6840 18165
rect 6800 18005 6805 18035
rect 6835 18005 6840 18035
rect 6800 17875 6840 18005
rect 6800 17845 6805 17875
rect 6835 17845 6840 17875
rect 6800 17715 6840 17845
rect 6800 17685 6805 17715
rect 6835 17685 6840 17715
rect 6800 17555 6840 17685
rect 6800 17525 6805 17555
rect 6835 17525 6840 17555
rect 6800 17395 6840 17525
rect 6800 17365 6805 17395
rect 6835 17365 6840 17395
rect 6800 17235 6840 17365
rect 6800 17205 6805 17235
rect 6835 17205 6840 17235
rect 6800 17200 6840 17205
rect 6880 18195 6920 18200
rect 6880 18165 6885 18195
rect 6915 18165 6920 18195
rect 6880 18035 6920 18165
rect 6880 18005 6885 18035
rect 6915 18005 6920 18035
rect 6880 17875 6920 18005
rect 6880 17845 6885 17875
rect 6915 17845 6920 17875
rect 6880 17715 6920 17845
rect 6880 17685 6885 17715
rect 6915 17685 6920 17715
rect 6880 17555 6920 17685
rect 6880 17525 6885 17555
rect 6915 17525 6920 17555
rect 6880 17395 6920 17525
rect 6880 17365 6885 17395
rect 6915 17365 6920 17395
rect 6880 17235 6920 17365
rect 6880 17205 6885 17235
rect 6915 17205 6920 17235
rect 6880 17200 6920 17205
rect 6960 18195 7000 18200
rect 6960 18165 6965 18195
rect 6995 18165 7000 18195
rect 6960 18035 7000 18165
rect 6960 18005 6965 18035
rect 6995 18005 7000 18035
rect 6960 17875 7000 18005
rect 6960 17845 6965 17875
rect 6995 17845 7000 17875
rect 6960 17715 7000 17845
rect 6960 17685 6965 17715
rect 6995 17685 7000 17715
rect 6960 17555 7000 17685
rect 6960 17525 6965 17555
rect 6995 17525 7000 17555
rect 6960 17395 7000 17525
rect 6960 17365 6965 17395
rect 6995 17365 7000 17395
rect 6960 17235 7000 17365
rect 6960 17205 6965 17235
rect 6995 17205 7000 17235
rect 6960 17200 7000 17205
rect 7040 18195 7080 18200
rect 7040 18165 7045 18195
rect 7075 18165 7080 18195
rect 7040 18035 7080 18165
rect 7040 18005 7045 18035
rect 7075 18005 7080 18035
rect 7040 17875 7080 18005
rect 7040 17845 7045 17875
rect 7075 17845 7080 17875
rect 7040 17715 7080 17845
rect 7040 17685 7045 17715
rect 7075 17685 7080 17715
rect 7040 17555 7080 17685
rect 7040 17525 7045 17555
rect 7075 17525 7080 17555
rect 7040 17395 7080 17525
rect 7040 17365 7045 17395
rect 7075 17365 7080 17395
rect 7040 17235 7080 17365
rect 7040 17205 7045 17235
rect 7075 17205 7080 17235
rect 7040 17200 7080 17205
rect 7120 18195 7160 18200
rect 7120 18165 7125 18195
rect 7155 18165 7160 18195
rect 7120 18035 7160 18165
rect 7120 18005 7125 18035
rect 7155 18005 7160 18035
rect 7120 17875 7160 18005
rect 7120 17845 7125 17875
rect 7155 17845 7160 17875
rect 7120 17715 7160 17845
rect 7120 17685 7125 17715
rect 7155 17685 7160 17715
rect 7120 17555 7160 17685
rect 7120 17525 7125 17555
rect 7155 17525 7160 17555
rect 7120 17395 7160 17525
rect 7120 17365 7125 17395
rect 7155 17365 7160 17395
rect 7120 17235 7160 17365
rect 7120 17205 7125 17235
rect 7155 17205 7160 17235
rect 7120 17200 7160 17205
rect 7200 18195 7240 18200
rect 7200 18165 7205 18195
rect 7235 18165 7240 18195
rect 7200 18035 7240 18165
rect 7200 18005 7205 18035
rect 7235 18005 7240 18035
rect 7200 17875 7240 18005
rect 7200 17845 7205 17875
rect 7235 17845 7240 17875
rect 7200 17715 7240 17845
rect 7200 17685 7205 17715
rect 7235 17685 7240 17715
rect 7200 17555 7240 17685
rect 7200 17525 7205 17555
rect 7235 17525 7240 17555
rect 7200 17395 7240 17525
rect 7200 17365 7205 17395
rect 7235 17365 7240 17395
rect 7200 17235 7240 17365
rect 7200 17205 7205 17235
rect 7235 17205 7240 17235
rect 7200 17200 7240 17205
rect 7280 18195 7320 18200
rect 7280 18165 7285 18195
rect 7315 18165 7320 18195
rect 7280 18035 7320 18165
rect 7280 18005 7285 18035
rect 7315 18005 7320 18035
rect 7280 17875 7320 18005
rect 7280 17845 7285 17875
rect 7315 17845 7320 17875
rect 7280 17715 7320 17845
rect 7280 17685 7285 17715
rect 7315 17685 7320 17715
rect 7280 17555 7320 17685
rect 7280 17525 7285 17555
rect 7315 17525 7320 17555
rect 7280 17395 7320 17525
rect 7280 17365 7285 17395
rect 7315 17365 7320 17395
rect 7280 17235 7320 17365
rect 7280 17205 7285 17235
rect 7315 17205 7320 17235
rect 7280 17200 7320 17205
rect 7360 18195 7400 18200
rect 7360 18165 7365 18195
rect 7395 18165 7400 18195
rect 7360 18035 7400 18165
rect 7360 18005 7365 18035
rect 7395 18005 7400 18035
rect 7360 17875 7400 18005
rect 7360 17845 7365 17875
rect 7395 17845 7400 17875
rect 7360 17715 7400 17845
rect 7360 17685 7365 17715
rect 7395 17685 7400 17715
rect 7360 17555 7400 17685
rect 7360 17525 7365 17555
rect 7395 17525 7400 17555
rect 7360 17395 7400 17525
rect 7360 17365 7365 17395
rect 7395 17365 7400 17395
rect 7360 17235 7400 17365
rect 7360 17205 7365 17235
rect 7395 17205 7400 17235
rect 7360 17200 7400 17205
rect 7440 18195 7480 18200
rect 7440 18165 7445 18195
rect 7475 18165 7480 18195
rect 7440 18035 7480 18165
rect 7440 18005 7445 18035
rect 7475 18005 7480 18035
rect 7440 17875 7480 18005
rect 7440 17845 7445 17875
rect 7475 17845 7480 17875
rect 7440 17715 7480 17845
rect 7440 17685 7445 17715
rect 7475 17685 7480 17715
rect 7440 17555 7480 17685
rect 7440 17525 7445 17555
rect 7475 17525 7480 17555
rect 7440 17395 7480 17525
rect 7440 17365 7445 17395
rect 7475 17365 7480 17395
rect 7440 17235 7480 17365
rect 7440 17205 7445 17235
rect 7475 17205 7480 17235
rect 7440 17200 7480 17205
rect 7520 18195 7560 18200
rect 7520 18165 7525 18195
rect 7555 18165 7560 18195
rect 7520 18035 7560 18165
rect 7520 18005 7525 18035
rect 7555 18005 7560 18035
rect 7520 17875 7560 18005
rect 7520 17845 7525 17875
rect 7555 17845 7560 17875
rect 7520 17715 7560 17845
rect 7520 17685 7525 17715
rect 7555 17685 7560 17715
rect 7520 17555 7560 17685
rect 7520 17525 7525 17555
rect 7555 17525 7560 17555
rect 7520 17395 7560 17525
rect 7520 17365 7525 17395
rect 7555 17365 7560 17395
rect 7520 17235 7560 17365
rect 7520 17205 7525 17235
rect 7555 17205 7560 17235
rect 7520 17200 7560 17205
rect 7600 18195 7640 18200
rect 7600 18165 7605 18195
rect 7635 18165 7640 18195
rect 7600 18035 7640 18165
rect 7600 18005 7605 18035
rect 7635 18005 7640 18035
rect 7600 17875 7640 18005
rect 7600 17845 7605 17875
rect 7635 17845 7640 17875
rect 7600 17715 7640 17845
rect 7600 17685 7605 17715
rect 7635 17685 7640 17715
rect 7600 17555 7640 17685
rect 7600 17525 7605 17555
rect 7635 17525 7640 17555
rect 7600 17395 7640 17525
rect 7600 17365 7605 17395
rect 7635 17365 7640 17395
rect 7600 17235 7640 17365
rect 7600 17205 7605 17235
rect 7635 17205 7640 17235
rect 7600 17200 7640 17205
rect 7680 18195 7720 18200
rect 7680 18165 7685 18195
rect 7715 18165 7720 18195
rect 7680 18035 7720 18165
rect 7680 18005 7685 18035
rect 7715 18005 7720 18035
rect 7680 17875 7720 18005
rect 7680 17845 7685 17875
rect 7715 17845 7720 17875
rect 7680 17715 7720 17845
rect 7680 17685 7685 17715
rect 7715 17685 7720 17715
rect 7680 17555 7720 17685
rect 7680 17525 7685 17555
rect 7715 17525 7720 17555
rect 7680 17395 7720 17525
rect 7680 17365 7685 17395
rect 7715 17365 7720 17395
rect 7680 17235 7720 17365
rect 7680 17205 7685 17235
rect 7715 17205 7720 17235
rect 7680 17200 7720 17205
rect 7760 18195 7800 18200
rect 7760 18165 7765 18195
rect 7795 18165 7800 18195
rect 7760 18035 7800 18165
rect 7760 18005 7765 18035
rect 7795 18005 7800 18035
rect 7760 17875 7800 18005
rect 7760 17845 7765 17875
rect 7795 17845 7800 17875
rect 7760 17715 7800 17845
rect 7760 17685 7765 17715
rect 7795 17685 7800 17715
rect 7760 17555 7800 17685
rect 7760 17525 7765 17555
rect 7795 17525 7800 17555
rect 7760 17395 7800 17525
rect 7760 17365 7765 17395
rect 7795 17365 7800 17395
rect 7760 17235 7800 17365
rect 7760 17205 7765 17235
rect 7795 17205 7800 17235
rect 7760 17200 7800 17205
rect 7840 18195 7880 18200
rect 7840 18165 7845 18195
rect 7875 18165 7880 18195
rect 7840 18035 7880 18165
rect 7840 18005 7845 18035
rect 7875 18005 7880 18035
rect 7840 17875 7880 18005
rect 7840 17845 7845 17875
rect 7875 17845 7880 17875
rect 7840 17715 7880 17845
rect 7840 17685 7845 17715
rect 7875 17685 7880 17715
rect 7840 17555 7880 17685
rect 7840 17525 7845 17555
rect 7875 17525 7880 17555
rect 7840 17395 7880 17525
rect 7840 17365 7845 17395
rect 7875 17365 7880 17395
rect 7840 17235 7880 17365
rect 7840 17205 7845 17235
rect 7875 17205 7880 17235
rect 7840 17200 7880 17205
rect 7920 18195 7960 18200
rect 7920 18165 7925 18195
rect 7955 18165 7960 18195
rect 7920 18035 7960 18165
rect 7920 18005 7925 18035
rect 7955 18005 7960 18035
rect 7920 17875 7960 18005
rect 7920 17845 7925 17875
rect 7955 17845 7960 17875
rect 7920 17715 7960 17845
rect 7920 17685 7925 17715
rect 7955 17685 7960 17715
rect 7920 17555 7960 17685
rect 7920 17525 7925 17555
rect 7955 17525 7960 17555
rect 7920 17395 7960 17525
rect 7920 17365 7925 17395
rect 7955 17365 7960 17395
rect 7920 17235 7960 17365
rect 7920 17205 7925 17235
rect 7955 17205 7960 17235
rect 7920 17200 7960 17205
rect 8000 18195 8040 18200
rect 8000 18165 8005 18195
rect 8035 18165 8040 18195
rect 8000 18035 8040 18165
rect 8000 18005 8005 18035
rect 8035 18005 8040 18035
rect 8000 17875 8040 18005
rect 8000 17845 8005 17875
rect 8035 17845 8040 17875
rect 8000 17715 8040 17845
rect 8000 17685 8005 17715
rect 8035 17685 8040 17715
rect 8000 17555 8040 17685
rect 8000 17525 8005 17555
rect 8035 17525 8040 17555
rect 8000 17395 8040 17525
rect 8000 17365 8005 17395
rect 8035 17365 8040 17395
rect 8000 17235 8040 17365
rect 8000 17205 8005 17235
rect 8035 17205 8040 17235
rect 8000 17200 8040 17205
rect 8080 18195 8120 18200
rect 8080 18165 8085 18195
rect 8115 18165 8120 18195
rect 8080 18035 8120 18165
rect 8080 18005 8085 18035
rect 8115 18005 8120 18035
rect 8080 17875 8120 18005
rect 8080 17845 8085 17875
rect 8115 17845 8120 17875
rect 8080 17715 8120 17845
rect 8080 17685 8085 17715
rect 8115 17685 8120 17715
rect 8080 17555 8120 17685
rect 8080 17525 8085 17555
rect 8115 17525 8120 17555
rect 8080 17395 8120 17525
rect 8080 17365 8085 17395
rect 8115 17365 8120 17395
rect 8080 17235 8120 17365
rect 8080 17205 8085 17235
rect 8115 17205 8120 17235
rect 8080 17200 8120 17205
rect 8160 18195 8200 18200
rect 8160 18165 8165 18195
rect 8195 18165 8200 18195
rect 8160 18035 8200 18165
rect 8160 18005 8165 18035
rect 8195 18005 8200 18035
rect 8160 17875 8200 18005
rect 8160 17845 8165 17875
rect 8195 17845 8200 17875
rect 8160 17715 8200 17845
rect 8160 17685 8165 17715
rect 8195 17685 8200 17715
rect 8160 17555 8200 17685
rect 8160 17525 8165 17555
rect 8195 17525 8200 17555
rect 8160 17395 8200 17525
rect 8160 17365 8165 17395
rect 8195 17365 8200 17395
rect 8160 17235 8200 17365
rect 8160 17205 8165 17235
rect 8195 17205 8200 17235
rect 8160 17200 8200 17205
rect 8240 18195 8280 18200
rect 8240 18165 8245 18195
rect 8275 18165 8280 18195
rect 8240 18035 8280 18165
rect 8240 18005 8245 18035
rect 8275 18005 8280 18035
rect 8240 17875 8280 18005
rect 8240 17845 8245 17875
rect 8275 17845 8280 17875
rect 8240 17715 8280 17845
rect 8240 17685 8245 17715
rect 8275 17685 8280 17715
rect 8240 17555 8280 17685
rect 8240 17525 8245 17555
rect 8275 17525 8280 17555
rect 8240 17395 8280 17525
rect 8240 17365 8245 17395
rect 8275 17365 8280 17395
rect 8240 17235 8280 17365
rect 8240 17205 8245 17235
rect 8275 17205 8280 17235
rect 8240 17200 8280 17205
rect 8320 18195 8360 18200
rect 8320 18165 8325 18195
rect 8355 18165 8360 18195
rect 8320 18035 8360 18165
rect 8320 18005 8325 18035
rect 8355 18005 8360 18035
rect 8320 17875 8360 18005
rect 8320 17845 8325 17875
rect 8355 17845 8360 17875
rect 8320 17715 8360 17845
rect 8320 17685 8325 17715
rect 8355 17685 8360 17715
rect 8320 17555 8360 17685
rect 8320 17525 8325 17555
rect 8355 17525 8360 17555
rect 8320 17395 8360 17525
rect 8320 17365 8325 17395
rect 8355 17365 8360 17395
rect 8320 17235 8360 17365
rect 8320 17205 8325 17235
rect 8355 17205 8360 17235
rect 8320 17200 8360 17205
rect 8400 18195 8440 18200
rect 8400 18165 8405 18195
rect 8435 18165 8440 18195
rect 8400 18035 8440 18165
rect 8400 18005 8405 18035
rect 8435 18005 8440 18035
rect 8400 17875 8440 18005
rect 8400 17845 8405 17875
rect 8435 17845 8440 17875
rect 8400 17715 8440 17845
rect 8400 17685 8405 17715
rect 8435 17685 8440 17715
rect 8400 17555 8440 17685
rect 8400 17525 8405 17555
rect 8435 17525 8440 17555
rect 8400 17395 8440 17525
rect 8400 17365 8405 17395
rect 8435 17365 8440 17395
rect 8400 17235 8440 17365
rect 8400 17205 8405 17235
rect 8435 17205 8440 17235
rect 8400 17200 8440 17205
rect 8480 18195 8520 18200
rect 8480 18165 8485 18195
rect 8515 18165 8520 18195
rect 8480 18035 8520 18165
rect 8480 18005 8485 18035
rect 8515 18005 8520 18035
rect 8480 17875 8520 18005
rect 8480 17845 8485 17875
rect 8515 17845 8520 17875
rect 8480 17715 8520 17845
rect 8480 17685 8485 17715
rect 8515 17685 8520 17715
rect 8480 17555 8520 17685
rect 8480 17525 8485 17555
rect 8515 17525 8520 17555
rect 8480 17395 8520 17525
rect 8480 17365 8485 17395
rect 8515 17365 8520 17395
rect 8480 17235 8520 17365
rect 8480 17205 8485 17235
rect 8515 17205 8520 17235
rect 8480 17200 8520 17205
rect 8560 18195 8600 18200
rect 8560 18165 8565 18195
rect 8595 18165 8600 18195
rect 8560 18035 8600 18165
rect 8560 18005 8565 18035
rect 8595 18005 8600 18035
rect 8560 17875 8600 18005
rect 8560 17845 8565 17875
rect 8595 17845 8600 17875
rect 8560 17715 8600 17845
rect 8560 17685 8565 17715
rect 8595 17685 8600 17715
rect 8560 17555 8600 17685
rect 8560 17525 8565 17555
rect 8595 17525 8600 17555
rect 8560 17395 8600 17525
rect 8560 17365 8565 17395
rect 8595 17365 8600 17395
rect 8560 17235 8600 17365
rect 8560 17205 8565 17235
rect 8595 17205 8600 17235
rect 8560 17200 8600 17205
rect 8640 18195 8680 18200
rect 8640 18165 8645 18195
rect 8675 18165 8680 18195
rect 8640 18035 8680 18165
rect 8640 18005 8645 18035
rect 8675 18005 8680 18035
rect 8640 17875 8680 18005
rect 8640 17845 8645 17875
rect 8675 17845 8680 17875
rect 8640 17715 8680 17845
rect 8640 17685 8645 17715
rect 8675 17685 8680 17715
rect 8640 17555 8680 17685
rect 8640 17525 8645 17555
rect 8675 17525 8680 17555
rect 8640 17395 8680 17525
rect 8640 17365 8645 17395
rect 8675 17365 8680 17395
rect 8640 17235 8680 17365
rect 8640 17205 8645 17235
rect 8675 17205 8680 17235
rect 8640 17200 8680 17205
rect 8720 18195 8760 18200
rect 8720 18165 8725 18195
rect 8755 18165 8760 18195
rect 8720 18035 8760 18165
rect 8720 18005 8725 18035
rect 8755 18005 8760 18035
rect 8720 17875 8760 18005
rect 8720 17845 8725 17875
rect 8755 17845 8760 17875
rect 8720 17715 8760 17845
rect 8720 17685 8725 17715
rect 8755 17685 8760 17715
rect 8720 17555 8760 17685
rect 8720 17525 8725 17555
rect 8755 17525 8760 17555
rect 8720 17395 8760 17525
rect 8720 17365 8725 17395
rect 8755 17365 8760 17395
rect 8720 17235 8760 17365
rect 8720 17205 8725 17235
rect 8755 17205 8760 17235
rect 8720 17200 8760 17205
rect 8800 18195 8840 18200
rect 8800 18165 8805 18195
rect 8835 18165 8840 18195
rect 8800 18035 8840 18165
rect 8800 18005 8805 18035
rect 8835 18005 8840 18035
rect 8800 17875 8840 18005
rect 8800 17845 8805 17875
rect 8835 17845 8840 17875
rect 8800 17715 8840 17845
rect 8800 17685 8805 17715
rect 8835 17685 8840 17715
rect 8800 17555 8840 17685
rect 8800 17525 8805 17555
rect 8835 17525 8840 17555
rect 8800 17395 8840 17525
rect 8800 17365 8805 17395
rect 8835 17365 8840 17395
rect 8800 17235 8840 17365
rect 8800 17205 8805 17235
rect 8835 17205 8840 17235
rect 8800 17200 8840 17205
rect 8880 18195 8920 18200
rect 8880 18165 8885 18195
rect 8915 18165 8920 18195
rect 8880 18035 8920 18165
rect 8880 18005 8885 18035
rect 8915 18005 8920 18035
rect 8880 17875 8920 18005
rect 8880 17845 8885 17875
rect 8915 17845 8920 17875
rect 8880 17715 8920 17845
rect 8880 17685 8885 17715
rect 8915 17685 8920 17715
rect 8880 17555 8920 17685
rect 8880 17525 8885 17555
rect 8915 17525 8920 17555
rect 8880 17395 8920 17525
rect 8880 17365 8885 17395
rect 8915 17365 8920 17395
rect 8880 17235 8920 17365
rect 8880 17205 8885 17235
rect 8915 17205 8920 17235
rect 8880 17200 8920 17205
rect 8960 18195 9000 18200
rect 8960 18165 8965 18195
rect 8995 18165 9000 18195
rect 8960 18035 9000 18165
rect 8960 18005 8965 18035
rect 8995 18005 9000 18035
rect 8960 17875 9000 18005
rect 8960 17845 8965 17875
rect 8995 17845 9000 17875
rect 8960 17715 9000 17845
rect 8960 17685 8965 17715
rect 8995 17685 9000 17715
rect 8960 17555 9000 17685
rect 8960 17525 8965 17555
rect 8995 17525 9000 17555
rect 8960 17395 9000 17525
rect 8960 17365 8965 17395
rect 8995 17365 9000 17395
rect 8960 17235 9000 17365
rect 8960 17205 8965 17235
rect 8995 17205 9000 17235
rect 8960 17200 9000 17205
rect 9040 18195 9080 18200
rect 9040 18165 9045 18195
rect 9075 18165 9080 18195
rect 9040 18035 9080 18165
rect 9040 18005 9045 18035
rect 9075 18005 9080 18035
rect 9040 17875 9080 18005
rect 9040 17845 9045 17875
rect 9075 17845 9080 17875
rect 9040 17715 9080 17845
rect 9040 17685 9045 17715
rect 9075 17685 9080 17715
rect 9040 17555 9080 17685
rect 9040 17525 9045 17555
rect 9075 17525 9080 17555
rect 9040 17395 9080 17525
rect 9040 17365 9045 17395
rect 9075 17365 9080 17395
rect 9040 17235 9080 17365
rect 9040 17205 9045 17235
rect 9075 17205 9080 17235
rect 9040 17200 9080 17205
rect 9120 18195 9160 18200
rect 9120 18165 9125 18195
rect 9155 18165 9160 18195
rect 9120 18035 9160 18165
rect 9120 18005 9125 18035
rect 9155 18005 9160 18035
rect 9120 17875 9160 18005
rect 9120 17845 9125 17875
rect 9155 17845 9160 17875
rect 9120 17715 9160 17845
rect 9120 17685 9125 17715
rect 9155 17685 9160 17715
rect 9120 17555 9160 17685
rect 9120 17525 9125 17555
rect 9155 17525 9160 17555
rect 9120 17395 9160 17525
rect 9120 17365 9125 17395
rect 9155 17365 9160 17395
rect 9120 17235 9160 17365
rect 9120 17205 9125 17235
rect 9155 17205 9160 17235
rect 9120 17200 9160 17205
rect 9200 18195 9240 18200
rect 9200 18165 9205 18195
rect 9235 18165 9240 18195
rect 9200 18035 9240 18165
rect 9200 18005 9205 18035
rect 9235 18005 9240 18035
rect 9200 17875 9240 18005
rect 9200 17845 9205 17875
rect 9235 17845 9240 17875
rect 9200 17715 9240 17845
rect 9200 17685 9205 17715
rect 9235 17685 9240 17715
rect 9200 17555 9240 17685
rect 9200 17525 9205 17555
rect 9235 17525 9240 17555
rect 9200 17395 9240 17525
rect 9200 17365 9205 17395
rect 9235 17365 9240 17395
rect 9200 17235 9240 17365
rect 9200 17205 9205 17235
rect 9235 17205 9240 17235
rect 9200 17200 9240 17205
rect 9280 18195 9320 18200
rect 9280 18165 9285 18195
rect 9315 18165 9320 18195
rect 9280 18035 9320 18165
rect 9280 18005 9285 18035
rect 9315 18005 9320 18035
rect 9280 17875 9320 18005
rect 9280 17845 9285 17875
rect 9315 17845 9320 17875
rect 9280 17715 9320 17845
rect 9280 17685 9285 17715
rect 9315 17685 9320 17715
rect 9280 17555 9320 17685
rect 9280 17525 9285 17555
rect 9315 17525 9320 17555
rect 9280 17395 9320 17525
rect 9280 17365 9285 17395
rect 9315 17365 9320 17395
rect 9280 17235 9320 17365
rect 9280 17205 9285 17235
rect 9315 17205 9320 17235
rect 9280 17200 9320 17205
rect 9360 18195 9400 18200
rect 9360 18165 9365 18195
rect 9395 18165 9400 18195
rect 9360 18035 9400 18165
rect 9360 18005 9365 18035
rect 9395 18005 9400 18035
rect 9360 17875 9400 18005
rect 9360 17845 9365 17875
rect 9395 17845 9400 17875
rect 9360 17715 9400 17845
rect 9360 17685 9365 17715
rect 9395 17685 9400 17715
rect 9360 17555 9400 17685
rect 9360 17525 9365 17555
rect 9395 17525 9400 17555
rect 9360 17395 9400 17525
rect 9360 17365 9365 17395
rect 9395 17365 9400 17395
rect 9360 17235 9400 17365
rect 9360 17205 9365 17235
rect 9395 17205 9400 17235
rect 9360 17200 9400 17205
rect 9440 18195 9480 18200
rect 9440 18165 9445 18195
rect 9475 18165 9480 18195
rect 9440 18035 9480 18165
rect 9440 18005 9445 18035
rect 9475 18005 9480 18035
rect 9440 17875 9480 18005
rect 9440 17845 9445 17875
rect 9475 17845 9480 17875
rect 9440 17715 9480 17845
rect 9440 17685 9445 17715
rect 9475 17685 9480 17715
rect 9440 17555 9480 17685
rect 9440 17525 9445 17555
rect 9475 17525 9480 17555
rect 9440 17395 9480 17525
rect 9440 17365 9445 17395
rect 9475 17365 9480 17395
rect 9440 17235 9480 17365
rect 9440 17205 9445 17235
rect 9475 17205 9480 17235
rect 9440 17200 9480 17205
rect 6240 17155 6280 17160
rect 6240 17125 6245 17155
rect 6275 17125 6280 17155
rect 6240 16995 6280 17125
rect 6240 16965 6245 16995
rect 6275 16965 6280 16995
rect 6240 16960 6280 16965
rect 6320 17155 6360 17160
rect 6320 17125 6325 17155
rect 6355 17125 6360 17155
rect 6320 16995 6360 17125
rect 6320 16965 6325 16995
rect 6355 16965 6360 16995
rect 6320 16960 6360 16965
rect 6400 17155 6440 17160
rect 6400 17125 6405 17155
rect 6435 17125 6440 17155
rect 6400 16995 6440 17125
rect 6400 16965 6405 16995
rect 6435 16965 6440 16995
rect 6400 16960 6440 16965
rect 6480 17155 6520 17160
rect 6480 17125 6485 17155
rect 6515 17125 6520 17155
rect 6480 16995 6520 17125
rect 6480 16965 6485 16995
rect 6515 16965 6520 16995
rect 6480 16960 6520 16965
rect 6560 17155 6600 17160
rect 6560 17125 6565 17155
rect 6595 17125 6600 17155
rect 6560 16995 6600 17125
rect 6560 16965 6565 16995
rect 6595 16965 6600 16995
rect 6560 16960 6600 16965
rect 6640 17155 6680 17160
rect 6640 17125 6645 17155
rect 6675 17125 6680 17155
rect 6640 16995 6680 17125
rect 6640 16965 6645 16995
rect 6675 16965 6680 16995
rect 6640 16960 6680 16965
rect 6720 17155 6760 17160
rect 6720 17125 6725 17155
rect 6755 17125 6760 17155
rect 6720 16995 6760 17125
rect 6720 16965 6725 16995
rect 6755 16965 6760 16995
rect 6720 16960 6760 16965
rect 6800 17155 6840 17160
rect 6800 17125 6805 17155
rect 6835 17125 6840 17155
rect 6800 16995 6840 17125
rect 6800 16965 6805 16995
rect 6835 16965 6840 16995
rect 6800 16960 6840 16965
rect 6880 17155 6920 17160
rect 6880 17125 6885 17155
rect 6915 17125 6920 17155
rect 6880 16995 6920 17125
rect 6880 16965 6885 16995
rect 6915 16965 6920 16995
rect 6880 16960 6920 16965
rect 6960 17155 7000 17160
rect 6960 17125 6965 17155
rect 6995 17125 7000 17155
rect 6960 16995 7000 17125
rect 6960 16965 6965 16995
rect 6995 16965 7000 16995
rect 6960 16960 7000 16965
rect 7040 17155 7080 17160
rect 7040 17125 7045 17155
rect 7075 17125 7080 17155
rect 7040 16995 7080 17125
rect 7040 16965 7045 16995
rect 7075 16965 7080 16995
rect 7040 16960 7080 16965
rect 7120 17155 7160 17160
rect 7120 17125 7125 17155
rect 7155 17125 7160 17155
rect 7120 16995 7160 17125
rect 7120 16965 7125 16995
rect 7155 16965 7160 16995
rect 7120 16960 7160 16965
rect 7200 17155 7240 17160
rect 7200 17125 7205 17155
rect 7235 17125 7240 17155
rect 7200 16995 7240 17125
rect 7200 16965 7205 16995
rect 7235 16965 7240 16995
rect 7200 16960 7240 16965
rect 7280 17155 7320 17160
rect 7280 17125 7285 17155
rect 7315 17125 7320 17155
rect 7280 16995 7320 17125
rect 7280 16965 7285 16995
rect 7315 16965 7320 16995
rect 7280 16960 7320 16965
rect 7360 17155 7400 17160
rect 7360 17125 7365 17155
rect 7395 17125 7400 17155
rect 7360 16995 7400 17125
rect 7360 16965 7365 16995
rect 7395 16965 7400 16995
rect 7360 16960 7400 16965
rect 7440 17155 7480 17160
rect 7440 17125 7445 17155
rect 7475 17125 7480 17155
rect 7440 16995 7480 17125
rect 7440 16965 7445 16995
rect 7475 16965 7480 16995
rect 7440 16960 7480 16965
rect 7520 17155 7560 17160
rect 7520 17125 7525 17155
rect 7555 17125 7560 17155
rect 7520 16995 7560 17125
rect 7520 16965 7525 16995
rect 7555 16965 7560 16995
rect 7520 16960 7560 16965
rect 7600 17155 7640 17160
rect 7600 17125 7605 17155
rect 7635 17125 7640 17155
rect 7600 16995 7640 17125
rect 7600 16965 7605 16995
rect 7635 16965 7640 16995
rect 7600 16960 7640 16965
rect 7680 17155 7720 17160
rect 7680 17125 7685 17155
rect 7715 17125 7720 17155
rect 7680 16995 7720 17125
rect 7680 16965 7685 16995
rect 7715 16965 7720 16995
rect 7680 16960 7720 16965
rect 7760 17155 7800 17160
rect 7760 17125 7765 17155
rect 7795 17125 7800 17155
rect 7760 16995 7800 17125
rect 7760 16965 7765 16995
rect 7795 16965 7800 16995
rect 7760 16960 7800 16965
rect 7840 17155 7880 17160
rect 7840 17125 7845 17155
rect 7875 17125 7880 17155
rect 7840 16995 7880 17125
rect 7840 16965 7845 16995
rect 7875 16965 7880 16995
rect 7840 16960 7880 16965
rect 7920 17155 7960 17160
rect 7920 17125 7925 17155
rect 7955 17125 7960 17155
rect 7920 16995 7960 17125
rect 7920 16965 7925 16995
rect 7955 16965 7960 16995
rect 7920 16960 7960 16965
rect 8000 17155 8040 17160
rect 8000 17125 8005 17155
rect 8035 17125 8040 17155
rect 8000 16995 8040 17125
rect 8000 16965 8005 16995
rect 8035 16965 8040 16995
rect 8000 16960 8040 16965
rect 8080 17155 8120 17160
rect 8080 17125 8085 17155
rect 8115 17125 8120 17155
rect 8080 16995 8120 17125
rect 8080 16965 8085 16995
rect 8115 16965 8120 16995
rect 8080 16960 8120 16965
rect 8160 17155 8200 17160
rect 8160 17125 8165 17155
rect 8195 17125 8200 17155
rect 8160 16995 8200 17125
rect 8160 16965 8165 16995
rect 8195 16965 8200 16995
rect 8160 16960 8200 16965
rect 8240 17155 8280 17160
rect 8240 17125 8245 17155
rect 8275 17125 8280 17155
rect 8240 16995 8280 17125
rect 8240 16965 8245 16995
rect 8275 16965 8280 16995
rect 8240 16960 8280 16965
rect 8320 17155 8360 17160
rect 8320 17125 8325 17155
rect 8355 17125 8360 17155
rect 8320 16995 8360 17125
rect 8320 16965 8325 16995
rect 8355 16965 8360 16995
rect 8320 16960 8360 16965
rect 8400 17155 8440 17160
rect 8400 17125 8405 17155
rect 8435 17125 8440 17155
rect 8400 16995 8440 17125
rect 8400 16965 8405 16995
rect 8435 16965 8440 16995
rect 8400 16960 8440 16965
rect 8480 17155 8520 17160
rect 8480 17125 8485 17155
rect 8515 17125 8520 17155
rect 8480 16995 8520 17125
rect 8480 16965 8485 16995
rect 8515 16965 8520 16995
rect 8480 16960 8520 16965
rect 8560 17155 8600 17160
rect 8560 17125 8565 17155
rect 8595 17125 8600 17155
rect 8560 16995 8600 17125
rect 8560 16965 8565 16995
rect 8595 16965 8600 16995
rect 8560 16960 8600 16965
rect 8640 17155 8680 17160
rect 8640 17125 8645 17155
rect 8675 17125 8680 17155
rect 8640 16995 8680 17125
rect 8640 16965 8645 16995
rect 8675 16965 8680 16995
rect 8640 16960 8680 16965
rect 8720 17155 8760 17160
rect 8720 17125 8725 17155
rect 8755 17125 8760 17155
rect 8720 16995 8760 17125
rect 8720 16965 8725 16995
rect 8755 16965 8760 16995
rect 8720 16960 8760 16965
rect 8800 17155 8840 17160
rect 8800 17125 8805 17155
rect 8835 17125 8840 17155
rect 8800 16995 8840 17125
rect 8800 16965 8805 16995
rect 8835 16965 8840 16995
rect 8800 16960 8840 16965
rect 8880 17155 8920 17160
rect 8880 17125 8885 17155
rect 8915 17125 8920 17155
rect 8880 16995 8920 17125
rect 8880 16965 8885 16995
rect 8915 16965 8920 16995
rect 8880 16960 8920 16965
rect 8960 17155 9000 17160
rect 8960 17125 8965 17155
rect 8995 17125 9000 17155
rect 8960 16995 9000 17125
rect 8960 16965 8965 16995
rect 8995 16965 9000 16995
rect 8960 16960 9000 16965
rect 9040 17155 9080 17160
rect 9040 17125 9045 17155
rect 9075 17125 9080 17155
rect 9040 16995 9080 17125
rect 9040 16965 9045 16995
rect 9075 16965 9080 16995
rect 9040 16960 9080 16965
rect 9120 17155 9160 17160
rect 9120 17125 9125 17155
rect 9155 17125 9160 17155
rect 9120 16995 9160 17125
rect 9120 16965 9125 16995
rect 9155 16965 9160 16995
rect 9120 16960 9160 16965
rect 9200 17155 9240 17160
rect 9200 17125 9205 17155
rect 9235 17125 9240 17155
rect 9200 16995 9240 17125
rect 9200 16965 9205 16995
rect 9235 16965 9240 16995
rect 9200 16960 9240 16965
rect 9280 17155 9320 17160
rect 9280 17125 9285 17155
rect 9315 17125 9320 17155
rect 9280 16995 9320 17125
rect 9280 16965 9285 16995
rect 9315 16965 9320 16995
rect 9280 16960 9320 16965
rect 9360 17155 9400 17160
rect 9360 17125 9365 17155
rect 9395 17125 9400 17155
rect 9360 16995 9400 17125
rect 9360 16965 9365 16995
rect 9395 16965 9400 16995
rect 9360 16960 9400 16965
rect 9440 17155 9480 17160
rect 9440 17125 9445 17155
rect 9475 17125 9480 17155
rect 9440 16995 9480 17125
rect 9440 16965 9445 16995
rect 9475 16965 9480 16995
rect 9440 16960 9480 16965
rect 6160 16885 6165 16915
rect 6195 16885 6200 16915
rect 6160 16755 6200 16885
rect 6160 16725 6165 16755
rect 6195 16725 6200 16755
rect 6160 16720 6200 16725
rect 6240 16915 6280 16920
rect 6240 16885 6245 16915
rect 6275 16885 6280 16915
rect 6240 16755 6280 16885
rect 6240 16725 6245 16755
rect 6275 16725 6280 16755
rect 6240 16720 6280 16725
rect 6320 16915 6360 16920
rect 6320 16885 6325 16915
rect 6355 16885 6360 16915
rect 6320 16755 6360 16885
rect 6320 16725 6325 16755
rect 6355 16725 6360 16755
rect 6320 16720 6360 16725
rect 6400 16915 6440 16920
rect 6400 16885 6405 16915
rect 6435 16885 6440 16915
rect 6400 16755 6440 16885
rect 6400 16725 6405 16755
rect 6435 16725 6440 16755
rect 6400 16720 6440 16725
rect 6480 16915 6520 16920
rect 6480 16885 6485 16915
rect 6515 16885 6520 16915
rect 6480 16755 6520 16885
rect 6480 16725 6485 16755
rect 6515 16725 6520 16755
rect 6480 16720 6520 16725
rect 6560 16915 6600 16920
rect 6560 16885 6565 16915
rect 6595 16885 6600 16915
rect 6560 16755 6600 16885
rect 6560 16725 6565 16755
rect 6595 16725 6600 16755
rect 6560 16720 6600 16725
rect 6640 16915 6680 16920
rect 6640 16885 6645 16915
rect 6675 16885 6680 16915
rect 6640 16755 6680 16885
rect 6640 16725 6645 16755
rect 6675 16725 6680 16755
rect 6640 16720 6680 16725
rect 6720 16915 6760 16920
rect 6720 16885 6725 16915
rect 6755 16885 6760 16915
rect 6720 16755 6760 16885
rect 6720 16725 6725 16755
rect 6755 16725 6760 16755
rect 6720 16720 6760 16725
rect 6800 16915 6840 16920
rect 6800 16885 6805 16915
rect 6835 16885 6840 16915
rect 6800 16755 6840 16885
rect 6800 16725 6805 16755
rect 6835 16725 6840 16755
rect 6800 16720 6840 16725
rect 6880 16915 6920 16920
rect 6880 16885 6885 16915
rect 6915 16885 6920 16915
rect 6880 16755 6920 16885
rect 6880 16725 6885 16755
rect 6915 16725 6920 16755
rect 6880 16720 6920 16725
rect 6960 16915 7000 16920
rect 6960 16885 6965 16915
rect 6995 16885 7000 16915
rect 6960 16755 7000 16885
rect 6960 16725 6965 16755
rect 6995 16725 7000 16755
rect 6960 16720 7000 16725
rect 7040 16915 7080 16920
rect 7040 16885 7045 16915
rect 7075 16885 7080 16915
rect 7040 16755 7080 16885
rect 7040 16725 7045 16755
rect 7075 16725 7080 16755
rect 7040 16720 7080 16725
rect 7120 16915 7160 16920
rect 7120 16885 7125 16915
rect 7155 16885 7160 16915
rect 7120 16755 7160 16885
rect 7120 16725 7125 16755
rect 7155 16725 7160 16755
rect 7120 16720 7160 16725
rect 7200 16915 7240 16920
rect 7200 16885 7205 16915
rect 7235 16885 7240 16915
rect 7200 16755 7240 16885
rect 7200 16725 7205 16755
rect 7235 16725 7240 16755
rect 7200 16720 7240 16725
rect 7280 16915 7320 16920
rect 7280 16885 7285 16915
rect 7315 16885 7320 16915
rect 7280 16755 7320 16885
rect 7280 16725 7285 16755
rect 7315 16725 7320 16755
rect 7280 16720 7320 16725
rect 7360 16915 7400 16920
rect 7360 16885 7365 16915
rect 7395 16885 7400 16915
rect 7360 16755 7400 16885
rect 7360 16725 7365 16755
rect 7395 16725 7400 16755
rect 7360 16720 7400 16725
rect 7440 16915 7480 16920
rect 7440 16885 7445 16915
rect 7475 16885 7480 16915
rect 7440 16755 7480 16885
rect 7440 16725 7445 16755
rect 7475 16725 7480 16755
rect 7440 16720 7480 16725
rect 7520 16915 7560 16920
rect 7520 16885 7525 16915
rect 7555 16885 7560 16915
rect 7520 16755 7560 16885
rect 7520 16725 7525 16755
rect 7555 16725 7560 16755
rect 7520 16720 7560 16725
rect 7600 16915 7640 16920
rect 7600 16885 7605 16915
rect 7635 16885 7640 16915
rect 7600 16755 7640 16885
rect 7600 16725 7605 16755
rect 7635 16725 7640 16755
rect 7600 16720 7640 16725
rect 7680 16915 7720 16920
rect 7680 16885 7685 16915
rect 7715 16885 7720 16915
rect 7680 16755 7720 16885
rect 7680 16725 7685 16755
rect 7715 16725 7720 16755
rect 7680 16720 7720 16725
rect 7760 16915 7800 16920
rect 7760 16885 7765 16915
rect 7795 16885 7800 16915
rect 7760 16755 7800 16885
rect 7760 16725 7765 16755
rect 7795 16725 7800 16755
rect 7760 16720 7800 16725
rect 7840 16915 7880 16920
rect 7840 16885 7845 16915
rect 7875 16885 7880 16915
rect 7840 16755 7880 16885
rect 7840 16725 7845 16755
rect 7875 16725 7880 16755
rect 7840 16720 7880 16725
rect 7920 16915 7960 16920
rect 7920 16885 7925 16915
rect 7955 16885 7960 16915
rect 7920 16755 7960 16885
rect 7920 16725 7925 16755
rect 7955 16725 7960 16755
rect 7920 16720 7960 16725
rect 8000 16915 8040 16920
rect 8000 16885 8005 16915
rect 8035 16885 8040 16915
rect 8000 16755 8040 16885
rect 8000 16725 8005 16755
rect 8035 16725 8040 16755
rect 8000 16720 8040 16725
rect 8080 16915 8120 16920
rect 8080 16885 8085 16915
rect 8115 16885 8120 16915
rect 8080 16755 8120 16885
rect 8080 16725 8085 16755
rect 8115 16725 8120 16755
rect 8080 16720 8120 16725
rect 8160 16915 8200 16920
rect 8160 16885 8165 16915
rect 8195 16885 8200 16915
rect 8160 16755 8200 16885
rect 8160 16725 8165 16755
rect 8195 16725 8200 16755
rect 8160 16720 8200 16725
rect 8240 16915 8280 16920
rect 8240 16885 8245 16915
rect 8275 16885 8280 16915
rect 8240 16755 8280 16885
rect 8240 16725 8245 16755
rect 8275 16725 8280 16755
rect 8240 16720 8280 16725
rect 8320 16915 8360 16920
rect 8320 16885 8325 16915
rect 8355 16885 8360 16915
rect 8320 16755 8360 16885
rect 8320 16725 8325 16755
rect 8355 16725 8360 16755
rect 8320 16720 8360 16725
rect 8400 16915 8440 16920
rect 8400 16885 8405 16915
rect 8435 16885 8440 16915
rect 8400 16755 8440 16885
rect 8400 16725 8405 16755
rect 8435 16725 8440 16755
rect 8400 16720 8440 16725
rect 8480 16915 8520 16920
rect 8480 16885 8485 16915
rect 8515 16885 8520 16915
rect 8480 16755 8520 16885
rect 8480 16725 8485 16755
rect 8515 16725 8520 16755
rect 8480 16720 8520 16725
rect 8560 16915 8600 16920
rect 8560 16885 8565 16915
rect 8595 16885 8600 16915
rect 8560 16755 8600 16885
rect 8560 16725 8565 16755
rect 8595 16725 8600 16755
rect 8560 16720 8600 16725
rect 8640 16915 8680 16920
rect 8640 16885 8645 16915
rect 8675 16885 8680 16915
rect 8640 16755 8680 16885
rect 8640 16725 8645 16755
rect 8675 16725 8680 16755
rect 8640 16720 8680 16725
rect 8720 16915 8760 16920
rect 8720 16885 8725 16915
rect 8755 16885 8760 16915
rect 8720 16755 8760 16885
rect 8720 16725 8725 16755
rect 8755 16725 8760 16755
rect 8720 16720 8760 16725
rect 8800 16915 8840 16920
rect 8800 16885 8805 16915
rect 8835 16885 8840 16915
rect 8800 16755 8840 16885
rect 8800 16725 8805 16755
rect 8835 16725 8840 16755
rect 8800 16720 8840 16725
rect 8880 16915 8920 16920
rect 8880 16885 8885 16915
rect 8915 16885 8920 16915
rect 8880 16755 8920 16885
rect 8880 16725 8885 16755
rect 8915 16725 8920 16755
rect 8880 16720 8920 16725
rect 8960 16915 9000 16920
rect 8960 16885 8965 16915
rect 8995 16885 9000 16915
rect 8960 16755 9000 16885
rect 8960 16725 8965 16755
rect 8995 16725 9000 16755
rect 8960 16720 9000 16725
rect 9040 16915 9080 16920
rect 9040 16885 9045 16915
rect 9075 16885 9080 16915
rect 9040 16755 9080 16885
rect 9040 16725 9045 16755
rect 9075 16725 9080 16755
rect 9040 16720 9080 16725
rect 9120 16915 9160 16920
rect 9120 16885 9125 16915
rect 9155 16885 9160 16915
rect 9120 16755 9160 16885
rect 9120 16725 9125 16755
rect 9155 16725 9160 16755
rect 9120 16720 9160 16725
rect 9200 16915 9240 16920
rect 9200 16885 9205 16915
rect 9235 16885 9240 16915
rect 9200 16755 9240 16885
rect 9200 16725 9205 16755
rect 9235 16725 9240 16755
rect 9200 16720 9240 16725
rect 9280 16915 9320 16920
rect 9280 16885 9285 16915
rect 9315 16885 9320 16915
rect 9280 16755 9320 16885
rect 9280 16725 9285 16755
rect 9315 16725 9320 16755
rect 9280 16720 9320 16725
rect 9360 16915 9400 16920
rect 9360 16885 9365 16915
rect 9395 16885 9400 16915
rect 9360 16755 9400 16885
rect 9360 16725 9365 16755
rect 9395 16725 9400 16755
rect 9360 16720 9400 16725
rect 9440 16915 9480 16920
rect 9440 16885 9445 16915
rect 9475 16885 9480 16915
rect 9440 16755 9480 16885
rect 9440 16725 9445 16755
rect 9475 16725 9480 16755
rect 9440 16720 9480 16725
rect 9520 16915 9560 18680
rect 9520 16885 9525 16915
rect 9555 16885 9560 16915
rect 9520 16755 9560 16885
rect 9520 16725 9525 16755
rect 9555 16725 9560 16755
rect 0 16675 40 16680
rect 0 16645 5 16675
rect 35 16645 40 16675
rect 0 16515 40 16645
rect 0 16485 5 16515
rect 35 16485 40 16515
rect 0 16480 40 16485
rect 80 16675 120 16680
rect 80 16645 85 16675
rect 115 16645 120 16675
rect 80 16515 120 16645
rect 80 16485 85 16515
rect 115 16485 120 16515
rect 80 16480 120 16485
rect 160 16675 200 16680
rect 160 16645 165 16675
rect 195 16645 200 16675
rect 160 16515 200 16645
rect 160 16485 165 16515
rect 195 16485 200 16515
rect 160 16480 200 16485
rect 240 16675 280 16680
rect 240 16645 245 16675
rect 275 16645 280 16675
rect 240 16515 280 16645
rect 240 16485 245 16515
rect 275 16485 280 16515
rect 240 16480 280 16485
rect 320 16675 360 16680
rect 320 16645 325 16675
rect 355 16645 360 16675
rect 320 16515 360 16645
rect 320 16485 325 16515
rect 355 16485 360 16515
rect 320 16480 360 16485
rect 400 16675 440 16680
rect 400 16645 405 16675
rect 435 16645 440 16675
rect 400 16515 440 16645
rect 400 16485 405 16515
rect 435 16485 440 16515
rect 400 16480 440 16485
rect 480 16675 520 16680
rect 480 16645 485 16675
rect 515 16645 520 16675
rect 480 16515 520 16645
rect 480 16485 485 16515
rect 515 16485 520 16515
rect 480 16480 520 16485
rect 560 16675 600 16680
rect 560 16645 565 16675
rect 595 16645 600 16675
rect 560 16515 600 16645
rect 560 16485 565 16515
rect 595 16485 600 16515
rect 560 16480 600 16485
rect 640 16675 680 16680
rect 640 16645 645 16675
rect 675 16645 680 16675
rect 640 16515 680 16645
rect 640 16485 645 16515
rect 675 16485 680 16515
rect 640 16480 680 16485
rect 720 16675 760 16680
rect 720 16645 725 16675
rect 755 16645 760 16675
rect 720 16515 760 16645
rect 720 16485 725 16515
rect 755 16485 760 16515
rect 720 16480 760 16485
rect 800 16675 840 16680
rect 800 16645 805 16675
rect 835 16645 840 16675
rect 800 16515 840 16645
rect 800 16485 805 16515
rect 835 16485 840 16515
rect 800 16480 840 16485
rect 880 16675 920 16680
rect 880 16645 885 16675
rect 915 16645 920 16675
rect 880 16515 920 16645
rect 880 16485 885 16515
rect 915 16485 920 16515
rect 880 16480 920 16485
rect 960 16675 1000 16680
rect 960 16645 965 16675
rect 995 16645 1000 16675
rect 960 16515 1000 16645
rect 960 16485 965 16515
rect 995 16485 1000 16515
rect 960 16480 1000 16485
rect 1040 16675 1080 16680
rect 1040 16645 1045 16675
rect 1075 16645 1080 16675
rect 1040 16515 1080 16645
rect 1040 16485 1045 16515
rect 1075 16485 1080 16515
rect 1040 16480 1080 16485
rect 1120 16675 1160 16680
rect 1120 16645 1125 16675
rect 1155 16645 1160 16675
rect 1120 16515 1160 16645
rect 1120 16485 1125 16515
rect 1155 16485 1160 16515
rect 1120 16480 1160 16485
rect 1200 16675 1240 16680
rect 1200 16645 1205 16675
rect 1235 16645 1240 16675
rect 1200 16515 1240 16645
rect 1200 16485 1205 16515
rect 1235 16485 1240 16515
rect 1200 16480 1240 16485
rect 1280 16675 1320 16680
rect 1280 16645 1285 16675
rect 1315 16645 1320 16675
rect 1280 16515 1320 16645
rect 1280 16485 1285 16515
rect 1315 16485 1320 16515
rect 1280 16480 1320 16485
rect 1360 16675 1400 16680
rect 1360 16645 1365 16675
rect 1395 16645 1400 16675
rect 1360 16515 1400 16645
rect 1360 16485 1365 16515
rect 1395 16485 1400 16515
rect 1360 16480 1400 16485
rect 1440 16675 1480 16680
rect 1440 16645 1445 16675
rect 1475 16645 1480 16675
rect 1440 16515 1480 16645
rect 1440 16485 1445 16515
rect 1475 16485 1480 16515
rect 1440 16480 1480 16485
rect 1520 16675 1560 16680
rect 1520 16645 1525 16675
rect 1555 16645 1560 16675
rect 1520 16515 1560 16645
rect 1520 16485 1525 16515
rect 1555 16485 1560 16515
rect 1520 16480 1560 16485
rect 1600 16675 1640 16680
rect 1600 16645 1605 16675
rect 1635 16645 1640 16675
rect 1600 16515 1640 16645
rect 1600 16485 1605 16515
rect 1635 16485 1640 16515
rect 1600 16480 1640 16485
rect 1680 16675 1720 16680
rect 1680 16645 1685 16675
rect 1715 16645 1720 16675
rect 1680 16515 1720 16645
rect 1680 16485 1685 16515
rect 1715 16485 1720 16515
rect 1680 16480 1720 16485
rect 1760 16675 1800 16680
rect 1760 16645 1765 16675
rect 1795 16645 1800 16675
rect 1760 16515 1800 16645
rect 1760 16485 1765 16515
rect 1795 16485 1800 16515
rect 1760 16480 1800 16485
rect 1840 16675 1880 16680
rect 1840 16645 1845 16675
rect 1875 16645 1880 16675
rect 1840 16515 1880 16645
rect 1840 16485 1845 16515
rect 1875 16485 1880 16515
rect 1840 16480 1880 16485
rect 1920 16675 1960 16680
rect 1920 16645 1925 16675
rect 1955 16645 1960 16675
rect 1920 16515 1960 16645
rect 1920 16485 1925 16515
rect 1955 16485 1960 16515
rect 1920 16480 1960 16485
rect 2000 16675 2040 16680
rect 2000 16645 2005 16675
rect 2035 16645 2040 16675
rect 2000 16515 2040 16645
rect 2000 16485 2005 16515
rect 2035 16485 2040 16515
rect 2000 16480 2040 16485
rect 2080 16675 2120 16680
rect 2080 16645 2085 16675
rect 2115 16645 2120 16675
rect 2080 16515 2120 16645
rect 2080 16485 2085 16515
rect 2115 16485 2120 16515
rect 2080 16480 2120 16485
rect 2160 16675 2200 16680
rect 2160 16645 2165 16675
rect 2195 16645 2200 16675
rect 2160 16515 2200 16645
rect 2160 16485 2165 16515
rect 2195 16485 2200 16515
rect 2160 16480 2200 16485
rect 2240 16675 2280 16680
rect 2240 16645 2245 16675
rect 2275 16645 2280 16675
rect 2240 16515 2280 16645
rect 2240 16485 2245 16515
rect 2275 16485 2280 16515
rect 2240 16480 2280 16485
rect 2320 16675 2360 16680
rect 2320 16645 2325 16675
rect 2355 16645 2360 16675
rect 2320 16515 2360 16645
rect 2320 16485 2325 16515
rect 2355 16485 2360 16515
rect 2320 16480 2360 16485
rect 2400 16675 2440 16680
rect 2400 16645 2405 16675
rect 2435 16645 2440 16675
rect 2400 16515 2440 16645
rect 2400 16485 2405 16515
rect 2435 16485 2440 16515
rect 2400 16480 2440 16485
rect 2480 16675 2520 16680
rect 2480 16645 2485 16675
rect 2515 16645 2520 16675
rect 2480 16515 2520 16645
rect 2480 16485 2485 16515
rect 2515 16485 2520 16515
rect 2480 16480 2520 16485
rect 2560 16675 2600 16680
rect 2560 16645 2565 16675
rect 2595 16645 2600 16675
rect 2560 16515 2600 16645
rect 2560 16485 2565 16515
rect 2595 16485 2600 16515
rect 2560 16480 2600 16485
rect 2640 16675 2680 16680
rect 2640 16645 2645 16675
rect 2675 16645 2680 16675
rect 2640 16515 2680 16645
rect 2640 16485 2645 16515
rect 2675 16485 2680 16515
rect 2640 16480 2680 16485
rect 2720 16675 2760 16680
rect 2720 16645 2725 16675
rect 2755 16645 2760 16675
rect 2720 16515 2760 16645
rect 2720 16485 2725 16515
rect 2755 16485 2760 16515
rect 2720 16480 2760 16485
rect 2800 16675 2840 16680
rect 2800 16645 2805 16675
rect 2835 16645 2840 16675
rect 2800 16515 2840 16645
rect 2800 16485 2805 16515
rect 2835 16485 2840 16515
rect 2800 16480 2840 16485
rect 2880 16675 2920 16680
rect 2880 16645 2885 16675
rect 2915 16645 2920 16675
rect 2880 16515 2920 16645
rect 2880 16485 2885 16515
rect 2915 16485 2920 16515
rect 2880 16480 2920 16485
rect 2960 16675 3000 16680
rect 2960 16645 2965 16675
rect 2995 16645 3000 16675
rect 2960 16515 3000 16645
rect 2960 16485 2965 16515
rect 2995 16485 3000 16515
rect 2960 16480 3000 16485
rect 3040 16675 3080 16680
rect 3040 16645 3045 16675
rect 3075 16645 3080 16675
rect 3040 16515 3080 16645
rect 3040 16485 3045 16515
rect 3075 16485 3080 16515
rect 3040 16480 3080 16485
rect 3120 16675 3160 16680
rect 3120 16645 3125 16675
rect 3155 16645 3160 16675
rect 3120 16515 3160 16645
rect 3120 16485 3125 16515
rect 3155 16485 3160 16515
rect 3120 16480 3160 16485
rect 3200 16675 3240 16680
rect 3200 16645 3205 16675
rect 3235 16645 3240 16675
rect 3200 16515 3240 16645
rect 3200 16485 3205 16515
rect 3235 16485 3240 16515
rect 3200 16480 3240 16485
rect 3280 16675 3320 16680
rect 3280 16645 3285 16675
rect 3315 16645 3320 16675
rect 3280 16515 3320 16645
rect 3280 16485 3285 16515
rect 3315 16485 3320 16515
rect 3280 16480 3320 16485
rect 3360 16675 3400 16680
rect 3360 16645 3365 16675
rect 3395 16645 3400 16675
rect 3360 16515 3400 16645
rect 3360 16485 3365 16515
rect 3395 16485 3400 16515
rect 3360 16480 3400 16485
rect 3440 16675 3480 16680
rect 3440 16645 3445 16675
rect 3475 16645 3480 16675
rect 3440 16515 3480 16645
rect 3440 16485 3445 16515
rect 3475 16485 3480 16515
rect 3440 16480 3480 16485
rect 3520 16675 3560 16680
rect 3520 16645 3525 16675
rect 3555 16645 3560 16675
rect 3520 16515 3560 16645
rect 3520 16485 3525 16515
rect 3555 16485 3560 16515
rect 3520 16480 3560 16485
rect 3600 16675 3640 16680
rect 3600 16645 3605 16675
rect 3635 16645 3640 16675
rect 3600 16515 3640 16645
rect 3600 16485 3605 16515
rect 3635 16485 3640 16515
rect 3600 16480 3640 16485
rect 3680 16675 3720 16680
rect 3680 16645 3685 16675
rect 3715 16645 3720 16675
rect 3680 16515 3720 16645
rect 3680 16485 3685 16515
rect 3715 16485 3720 16515
rect 3680 16480 3720 16485
rect 3760 16675 3800 16680
rect 3760 16645 3765 16675
rect 3795 16645 3800 16675
rect 3760 16515 3800 16645
rect 3760 16485 3765 16515
rect 3795 16485 3800 16515
rect 3760 16480 3800 16485
rect 3840 16675 3880 16680
rect 3840 16645 3845 16675
rect 3875 16645 3880 16675
rect 3840 16515 3880 16645
rect 3840 16485 3845 16515
rect 3875 16485 3880 16515
rect 3840 16480 3880 16485
rect 3920 16675 3960 16680
rect 3920 16645 3925 16675
rect 3955 16645 3960 16675
rect 3920 16515 3960 16645
rect 3920 16485 3925 16515
rect 3955 16485 3960 16515
rect 3920 16480 3960 16485
rect 4000 16675 4040 16680
rect 4000 16645 4005 16675
rect 4035 16645 4040 16675
rect 4000 16515 4040 16645
rect 4000 16485 4005 16515
rect 4035 16485 4040 16515
rect 4000 16480 4040 16485
rect 4080 16675 4120 16680
rect 4080 16645 4085 16675
rect 4115 16645 4120 16675
rect 4080 16515 4120 16645
rect 4080 16485 4085 16515
rect 4115 16485 4120 16515
rect 4080 16480 4120 16485
rect 4160 16675 4200 16680
rect 4160 16645 4165 16675
rect 4195 16645 4200 16675
rect 4160 16515 4200 16645
rect 4160 16485 4165 16515
rect 4195 16485 4200 16515
rect 4160 16480 4200 16485
rect 4240 16675 4280 16680
rect 4240 16645 4245 16675
rect 4275 16645 4280 16675
rect 4240 16515 4280 16645
rect 4240 16485 4245 16515
rect 4275 16485 4280 16515
rect 0 16435 40 16440
rect 0 16405 5 16435
rect 35 16405 40 16435
rect 0 16275 40 16405
rect 0 16245 5 16275
rect 35 16245 40 16275
rect 0 16240 40 16245
rect 80 16435 120 16440
rect 80 16405 85 16435
rect 115 16405 120 16435
rect 80 16275 120 16405
rect 80 16245 85 16275
rect 115 16245 120 16275
rect 80 16240 120 16245
rect 160 16435 200 16440
rect 160 16405 165 16435
rect 195 16405 200 16435
rect 160 16275 200 16405
rect 160 16245 165 16275
rect 195 16245 200 16275
rect 160 16240 200 16245
rect 240 16435 280 16440
rect 240 16405 245 16435
rect 275 16405 280 16435
rect 240 16275 280 16405
rect 240 16245 245 16275
rect 275 16245 280 16275
rect 240 16240 280 16245
rect 320 16435 360 16440
rect 320 16405 325 16435
rect 355 16405 360 16435
rect 320 16275 360 16405
rect 320 16245 325 16275
rect 355 16245 360 16275
rect 320 16240 360 16245
rect 400 16435 440 16440
rect 400 16405 405 16435
rect 435 16405 440 16435
rect 400 16275 440 16405
rect 400 16245 405 16275
rect 435 16245 440 16275
rect 400 16240 440 16245
rect 480 16435 520 16440
rect 480 16405 485 16435
rect 515 16405 520 16435
rect 480 16275 520 16405
rect 480 16245 485 16275
rect 515 16245 520 16275
rect 480 16240 520 16245
rect 560 16435 600 16440
rect 560 16405 565 16435
rect 595 16405 600 16435
rect 560 16275 600 16405
rect 560 16245 565 16275
rect 595 16245 600 16275
rect 560 16240 600 16245
rect 640 16435 680 16440
rect 640 16405 645 16435
rect 675 16405 680 16435
rect 640 16275 680 16405
rect 640 16245 645 16275
rect 675 16245 680 16275
rect 640 16240 680 16245
rect 720 16435 760 16440
rect 720 16405 725 16435
rect 755 16405 760 16435
rect 720 16275 760 16405
rect 720 16245 725 16275
rect 755 16245 760 16275
rect 720 16240 760 16245
rect 800 16435 840 16440
rect 800 16405 805 16435
rect 835 16405 840 16435
rect 800 16275 840 16405
rect 800 16245 805 16275
rect 835 16245 840 16275
rect 800 16240 840 16245
rect 880 16435 920 16440
rect 880 16405 885 16435
rect 915 16405 920 16435
rect 880 16275 920 16405
rect 880 16245 885 16275
rect 915 16245 920 16275
rect 880 16240 920 16245
rect 960 16435 1000 16440
rect 960 16405 965 16435
rect 995 16405 1000 16435
rect 960 16275 1000 16405
rect 960 16245 965 16275
rect 995 16245 1000 16275
rect 960 16240 1000 16245
rect 1040 16435 1080 16440
rect 1040 16405 1045 16435
rect 1075 16405 1080 16435
rect 1040 16275 1080 16405
rect 1040 16245 1045 16275
rect 1075 16245 1080 16275
rect 1040 16240 1080 16245
rect 1120 16435 1160 16440
rect 1120 16405 1125 16435
rect 1155 16405 1160 16435
rect 1120 16275 1160 16405
rect 1120 16245 1125 16275
rect 1155 16245 1160 16275
rect 1120 16240 1160 16245
rect 1200 16435 1240 16440
rect 1200 16405 1205 16435
rect 1235 16405 1240 16435
rect 1200 16275 1240 16405
rect 1200 16245 1205 16275
rect 1235 16245 1240 16275
rect 1200 16240 1240 16245
rect 1280 16435 1320 16440
rect 1280 16405 1285 16435
rect 1315 16405 1320 16435
rect 1280 16275 1320 16405
rect 1280 16245 1285 16275
rect 1315 16245 1320 16275
rect 1280 16240 1320 16245
rect 1360 16435 1400 16440
rect 1360 16405 1365 16435
rect 1395 16405 1400 16435
rect 1360 16275 1400 16405
rect 1360 16245 1365 16275
rect 1395 16245 1400 16275
rect 1360 16240 1400 16245
rect 1440 16435 1480 16440
rect 1440 16405 1445 16435
rect 1475 16405 1480 16435
rect 1440 16275 1480 16405
rect 1440 16245 1445 16275
rect 1475 16245 1480 16275
rect 1440 16240 1480 16245
rect 1520 16435 1560 16440
rect 1520 16405 1525 16435
rect 1555 16405 1560 16435
rect 1520 16275 1560 16405
rect 1520 16245 1525 16275
rect 1555 16245 1560 16275
rect 1520 16240 1560 16245
rect 1600 16435 1640 16440
rect 1600 16405 1605 16435
rect 1635 16405 1640 16435
rect 1600 16275 1640 16405
rect 1600 16245 1605 16275
rect 1635 16245 1640 16275
rect 1600 16240 1640 16245
rect 1680 16435 1720 16440
rect 1680 16405 1685 16435
rect 1715 16405 1720 16435
rect 1680 16275 1720 16405
rect 1680 16245 1685 16275
rect 1715 16245 1720 16275
rect 1680 16240 1720 16245
rect 1760 16435 1800 16440
rect 1760 16405 1765 16435
rect 1795 16405 1800 16435
rect 1760 16275 1800 16405
rect 1760 16245 1765 16275
rect 1795 16245 1800 16275
rect 1760 16240 1800 16245
rect 1840 16435 1880 16440
rect 1840 16405 1845 16435
rect 1875 16405 1880 16435
rect 1840 16275 1880 16405
rect 1840 16245 1845 16275
rect 1875 16245 1880 16275
rect 1840 16240 1880 16245
rect 1920 16435 1960 16440
rect 1920 16405 1925 16435
rect 1955 16405 1960 16435
rect 1920 16275 1960 16405
rect 1920 16245 1925 16275
rect 1955 16245 1960 16275
rect 1920 16240 1960 16245
rect 2000 16435 2040 16440
rect 2000 16405 2005 16435
rect 2035 16405 2040 16435
rect 2000 16275 2040 16405
rect 2000 16245 2005 16275
rect 2035 16245 2040 16275
rect 2000 16240 2040 16245
rect 2080 16435 2120 16440
rect 2080 16405 2085 16435
rect 2115 16405 2120 16435
rect 2080 16275 2120 16405
rect 2080 16245 2085 16275
rect 2115 16245 2120 16275
rect 2080 16240 2120 16245
rect 2160 16435 2200 16440
rect 2160 16405 2165 16435
rect 2195 16405 2200 16435
rect 2160 16275 2200 16405
rect 2160 16245 2165 16275
rect 2195 16245 2200 16275
rect 2160 16240 2200 16245
rect 2240 16435 2280 16440
rect 2240 16405 2245 16435
rect 2275 16405 2280 16435
rect 2240 16275 2280 16405
rect 2240 16245 2245 16275
rect 2275 16245 2280 16275
rect 2240 16240 2280 16245
rect 2320 16435 2360 16440
rect 2320 16405 2325 16435
rect 2355 16405 2360 16435
rect 2320 16275 2360 16405
rect 2320 16245 2325 16275
rect 2355 16245 2360 16275
rect 2320 16240 2360 16245
rect 2400 16435 2440 16440
rect 2400 16405 2405 16435
rect 2435 16405 2440 16435
rect 2400 16275 2440 16405
rect 2400 16245 2405 16275
rect 2435 16245 2440 16275
rect 2400 16240 2440 16245
rect 2480 16435 2520 16440
rect 2480 16405 2485 16435
rect 2515 16405 2520 16435
rect 2480 16275 2520 16405
rect 2480 16245 2485 16275
rect 2515 16245 2520 16275
rect 2480 16240 2520 16245
rect 2560 16435 2600 16440
rect 2560 16405 2565 16435
rect 2595 16405 2600 16435
rect 2560 16275 2600 16405
rect 2560 16245 2565 16275
rect 2595 16245 2600 16275
rect 2560 16240 2600 16245
rect 2640 16435 2680 16440
rect 2640 16405 2645 16435
rect 2675 16405 2680 16435
rect 2640 16275 2680 16405
rect 2640 16245 2645 16275
rect 2675 16245 2680 16275
rect 2640 16240 2680 16245
rect 2720 16435 2760 16440
rect 2720 16405 2725 16435
rect 2755 16405 2760 16435
rect 2720 16275 2760 16405
rect 2720 16245 2725 16275
rect 2755 16245 2760 16275
rect 2720 16240 2760 16245
rect 2800 16435 2840 16440
rect 2800 16405 2805 16435
rect 2835 16405 2840 16435
rect 2800 16275 2840 16405
rect 2800 16245 2805 16275
rect 2835 16245 2840 16275
rect 2800 16240 2840 16245
rect 2880 16435 2920 16440
rect 2880 16405 2885 16435
rect 2915 16405 2920 16435
rect 2880 16275 2920 16405
rect 2880 16245 2885 16275
rect 2915 16245 2920 16275
rect 2880 16240 2920 16245
rect 2960 16435 3000 16440
rect 2960 16405 2965 16435
rect 2995 16405 3000 16435
rect 2960 16275 3000 16405
rect 2960 16245 2965 16275
rect 2995 16245 3000 16275
rect 2960 16240 3000 16245
rect 3040 16435 3080 16440
rect 3040 16405 3045 16435
rect 3075 16405 3080 16435
rect 3040 16275 3080 16405
rect 3040 16245 3045 16275
rect 3075 16245 3080 16275
rect 3040 16240 3080 16245
rect 3120 16435 3160 16440
rect 3120 16405 3125 16435
rect 3155 16405 3160 16435
rect 3120 16275 3160 16405
rect 3120 16245 3125 16275
rect 3155 16245 3160 16275
rect 3120 16240 3160 16245
rect 3200 16435 3240 16440
rect 3200 16405 3205 16435
rect 3235 16405 3240 16435
rect 3200 16275 3240 16405
rect 3200 16245 3205 16275
rect 3235 16245 3240 16275
rect 3200 16240 3240 16245
rect 3280 16435 3320 16440
rect 3280 16405 3285 16435
rect 3315 16405 3320 16435
rect 3280 16275 3320 16405
rect 3280 16245 3285 16275
rect 3315 16245 3320 16275
rect 3280 16240 3320 16245
rect 3360 16435 3400 16440
rect 3360 16405 3365 16435
rect 3395 16405 3400 16435
rect 3360 16275 3400 16405
rect 3360 16245 3365 16275
rect 3395 16245 3400 16275
rect 3360 16240 3400 16245
rect 3440 16435 3480 16440
rect 3440 16405 3445 16435
rect 3475 16405 3480 16435
rect 3440 16275 3480 16405
rect 3440 16245 3445 16275
rect 3475 16245 3480 16275
rect 3440 16240 3480 16245
rect 3520 16435 3560 16440
rect 3520 16405 3525 16435
rect 3555 16405 3560 16435
rect 3520 16275 3560 16405
rect 3520 16245 3525 16275
rect 3555 16245 3560 16275
rect 3520 16240 3560 16245
rect 3600 16435 3640 16440
rect 3600 16405 3605 16435
rect 3635 16405 3640 16435
rect 3600 16275 3640 16405
rect 3600 16245 3605 16275
rect 3635 16245 3640 16275
rect 3600 16240 3640 16245
rect 3680 16435 3720 16440
rect 3680 16405 3685 16435
rect 3715 16405 3720 16435
rect 3680 16275 3720 16405
rect 3680 16245 3685 16275
rect 3715 16245 3720 16275
rect 3680 16240 3720 16245
rect 3760 16435 3800 16440
rect 3760 16405 3765 16435
rect 3795 16405 3800 16435
rect 3760 16275 3800 16405
rect 3760 16245 3765 16275
rect 3795 16245 3800 16275
rect 3760 16240 3800 16245
rect 3840 16435 3880 16440
rect 3840 16405 3845 16435
rect 3875 16405 3880 16435
rect 3840 16275 3880 16405
rect 3840 16245 3845 16275
rect 3875 16245 3880 16275
rect 3840 16240 3880 16245
rect 3920 16435 3960 16440
rect 3920 16405 3925 16435
rect 3955 16405 3960 16435
rect 3920 16275 3960 16405
rect 3920 16245 3925 16275
rect 3955 16245 3960 16275
rect 3920 16240 3960 16245
rect 4000 16435 4040 16440
rect 4000 16405 4005 16435
rect 4035 16405 4040 16435
rect 4000 16275 4040 16405
rect 4000 16245 4005 16275
rect 4035 16245 4040 16275
rect 4000 16240 4040 16245
rect 4080 16435 4120 16440
rect 4080 16405 4085 16435
rect 4115 16405 4120 16435
rect 4080 16275 4120 16405
rect 4080 16245 4085 16275
rect 4115 16245 4120 16275
rect 4080 16240 4120 16245
rect 4160 16435 4200 16440
rect 4160 16405 4165 16435
rect 4195 16405 4200 16435
rect 4160 16275 4200 16405
rect 4160 16245 4165 16275
rect 4195 16245 4200 16275
rect 4160 16240 4200 16245
rect 0 16195 40 16200
rect 0 16165 5 16195
rect 35 16165 40 16195
rect 0 16035 40 16165
rect 0 16005 5 16035
rect 35 16005 40 16035
rect 0 15875 40 16005
rect 0 15845 5 15875
rect 35 15845 40 15875
rect 0 15715 40 15845
rect 0 15685 5 15715
rect 35 15685 40 15715
rect 0 15555 40 15685
rect 0 15525 5 15555
rect 35 15525 40 15555
rect 0 15395 40 15525
rect 0 15365 5 15395
rect 35 15365 40 15395
rect 0 15235 40 15365
rect 0 15205 5 15235
rect 35 15205 40 15235
rect 0 15200 40 15205
rect 80 16195 120 16200
rect 80 16165 85 16195
rect 115 16165 120 16195
rect 80 16035 120 16165
rect 80 16005 85 16035
rect 115 16005 120 16035
rect 80 15875 120 16005
rect 80 15845 85 15875
rect 115 15845 120 15875
rect 80 15715 120 15845
rect 80 15685 85 15715
rect 115 15685 120 15715
rect 80 15555 120 15685
rect 80 15525 85 15555
rect 115 15525 120 15555
rect 80 15395 120 15525
rect 80 15365 85 15395
rect 115 15365 120 15395
rect 80 15235 120 15365
rect 80 15205 85 15235
rect 115 15205 120 15235
rect 80 15200 120 15205
rect 160 16195 200 16200
rect 160 16165 165 16195
rect 195 16165 200 16195
rect 160 16035 200 16165
rect 160 16005 165 16035
rect 195 16005 200 16035
rect 160 15875 200 16005
rect 160 15845 165 15875
rect 195 15845 200 15875
rect 160 15715 200 15845
rect 160 15685 165 15715
rect 195 15685 200 15715
rect 160 15555 200 15685
rect 160 15525 165 15555
rect 195 15525 200 15555
rect 160 15395 200 15525
rect 160 15365 165 15395
rect 195 15365 200 15395
rect 160 15235 200 15365
rect 160 15205 165 15235
rect 195 15205 200 15235
rect 160 15200 200 15205
rect 240 16195 280 16200
rect 240 16165 245 16195
rect 275 16165 280 16195
rect 240 16035 280 16165
rect 240 16005 245 16035
rect 275 16005 280 16035
rect 240 15875 280 16005
rect 240 15845 245 15875
rect 275 15845 280 15875
rect 240 15715 280 15845
rect 240 15685 245 15715
rect 275 15685 280 15715
rect 240 15555 280 15685
rect 240 15525 245 15555
rect 275 15525 280 15555
rect 240 15395 280 15525
rect 240 15365 245 15395
rect 275 15365 280 15395
rect 240 15235 280 15365
rect 240 15205 245 15235
rect 275 15205 280 15235
rect 240 15200 280 15205
rect 320 16195 360 16200
rect 320 16165 325 16195
rect 355 16165 360 16195
rect 320 16035 360 16165
rect 320 16005 325 16035
rect 355 16005 360 16035
rect 320 15875 360 16005
rect 320 15845 325 15875
rect 355 15845 360 15875
rect 320 15715 360 15845
rect 320 15685 325 15715
rect 355 15685 360 15715
rect 320 15555 360 15685
rect 320 15525 325 15555
rect 355 15525 360 15555
rect 320 15395 360 15525
rect 320 15365 325 15395
rect 355 15365 360 15395
rect 320 15235 360 15365
rect 320 15205 325 15235
rect 355 15205 360 15235
rect 320 15200 360 15205
rect 400 16195 440 16200
rect 400 16165 405 16195
rect 435 16165 440 16195
rect 400 16035 440 16165
rect 400 16005 405 16035
rect 435 16005 440 16035
rect 400 15875 440 16005
rect 400 15845 405 15875
rect 435 15845 440 15875
rect 400 15715 440 15845
rect 400 15685 405 15715
rect 435 15685 440 15715
rect 400 15555 440 15685
rect 400 15525 405 15555
rect 435 15525 440 15555
rect 400 15395 440 15525
rect 400 15365 405 15395
rect 435 15365 440 15395
rect 400 15235 440 15365
rect 400 15205 405 15235
rect 435 15205 440 15235
rect 400 15200 440 15205
rect 480 16195 520 16200
rect 480 16165 485 16195
rect 515 16165 520 16195
rect 480 16035 520 16165
rect 480 16005 485 16035
rect 515 16005 520 16035
rect 480 15875 520 16005
rect 480 15845 485 15875
rect 515 15845 520 15875
rect 480 15715 520 15845
rect 480 15685 485 15715
rect 515 15685 520 15715
rect 480 15555 520 15685
rect 480 15525 485 15555
rect 515 15525 520 15555
rect 480 15395 520 15525
rect 480 15365 485 15395
rect 515 15365 520 15395
rect 480 15235 520 15365
rect 480 15205 485 15235
rect 515 15205 520 15235
rect 480 15200 520 15205
rect 560 16195 600 16200
rect 560 16165 565 16195
rect 595 16165 600 16195
rect 560 16035 600 16165
rect 560 16005 565 16035
rect 595 16005 600 16035
rect 560 15875 600 16005
rect 560 15845 565 15875
rect 595 15845 600 15875
rect 560 15715 600 15845
rect 560 15685 565 15715
rect 595 15685 600 15715
rect 560 15555 600 15685
rect 560 15525 565 15555
rect 595 15525 600 15555
rect 560 15395 600 15525
rect 560 15365 565 15395
rect 595 15365 600 15395
rect 560 15235 600 15365
rect 560 15205 565 15235
rect 595 15205 600 15235
rect 560 15200 600 15205
rect 640 16195 680 16200
rect 640 16165 645 16195
rect 675 16165 680 16195
rect 640 16035 680 16165
rect 640 16005 645 16035
rect 675 16005 680 16035
rect 640 15875 680 16005
rect 640 15845 645 15875
rect 675 15845 680 15875
rect 640 15715 680 15845
rect 640 15685 645 15715
rect 675 15685 680 15715
rect 640 15555 680 15685
rect 640 15525 645 15555
rect 675 15525 680 15555
rect 640 15395 680 15525
rect 640 15365 645 15395
rect 675 15365 680 15395
rect 640 15235 680 15365
rect 640 15205 645 15235
rect 675 15205 680 15235
rect 640 15200 680 15205
rect 720 16195 760 16200
rect 720 16165 725 16195
rect 755 16165 760 16195
rect 720 16035 760 16165
rect 720 16005 725 16035
rect 755 16005 760 16035
rect 720 15875 760 16005
rect 720 15845 725 15875
rect 755 15845 760 15875
rect 720 15715 760 15845
rect 720 15685 725 15715
rect 755 15685 760 15715
rect 720 15555 760 15685
rect 720 15525 725 15555
rect 755 15525 760 15555
rect 720 15395 760 15525
rect 720 15365 725 15395
rect 755 15365 760 15395
rect 720 15235 760 15365
rect 720 15205 725 15235
rect 755 15205 760 15235
rect 720 15200 760 15205
rect 800 16195 840 16200
rect 800 16165 805 16195
rect 835 16165 840 16195
rect 800 16035 840 16165
rect 800 16005 805 16035
rect 835 16005 840 16035
rect 800 15875 840 16005
rect 800 15845 805 15875
rect 835 15845 840 15875
rect 800 15715 840 15845
rect 800 15685 805 15715
rect 835 15685 840 15715
rect 800 15555 840 15685
rect 800 15525 805 15555
rect 835 15525 840 15555
rect 800 15395 840 15525
rect 800 15365 805 15395
rect 835 15365 840 15395
rect 800 15235 840 15365
rect 800 15205 805 15235
rect 835 15205 840 15235
rect 800 15200 840 15205
rect 880 16195 920 16200
rect 880 16165 885 16195
rect 915 16165 920 16195
rect 880 16035 920 16165
rect 880 16005 885 16035
rect 915 16005 920 16035
rect 880 15875 920 16005
rect 880 15845 885 15875
rect 915 15845 920 15875
rect 880 15715 920 15845
rect 880 15685 885 15715
rect 915 15685 920 15715
rect 880 15555 920 15685
rect 880 15525 885 15555
rect 915 15525 920 15555
rect 880 15395 920 15525
rect 880 15365 885 15395
rect 915 15365 920 15395
rect 880 15235 920 15365
rect 880 15205 885 15235
rect 915 15205 920 15235
rect 880 15200 920 15205
rect 960 16195 1000 16200
rect 960 16165 965 16195
rect 995 16165 1000 16195
rect 960 16035 1000 16165
rect 960 16005 965 16035
rect 995 16005 1000 16035
rect 960 15875 1000 16005
rect 960 15845 965 15875
rect 995 15845 1000 15875
rect 960 15715 1000 15845
rect 960 15685 965 15715
rect 995 15685 1000 15715
rect 960 15555 1000 15685
rect 960 15525 965 15555
rect 995 15525 1000 15555
rect 960 15395 1000 15525
rect 960 15365 965 15395
rect 995 15365 1000 15395
rect 960 15235 1000 15365
rect 960 15205 965 15235
rect 995 15205 1000 15235
rect 960 15200 1000 15205
rect 1040 16195 1080 16200
rect 1040 16165 1045 16195
rect 1075 16165 1080 16195
rect 1040 16035 1080 16165
rect 1040 16005 1045 16035
rect 1075 16005 1080 16035
rect 1040 15875 1080 16005
rect 1040 15845 1045 15875
rect 1075 15845 1080 15875
rect 1040 15715 1080 15845
rect 1040 15685 1045 15715
rect 1075 15685 1080 15715
rect 1040 15555 1080 15685
rect 1040 15525 1045 15555
rect 1075 15525 1080 15555
rect 1040 15395 1080 15525
rect 1040 15365 1045 15395
rect 1075 15365 1080 15395
rect 1040 15235 1080 15365
rect 1040 15205 1045 15235
rect 1075 15205 1080 15235
rect 1040 15200 1080 15205
rect 1120 16195 1160 16200
rect 1120 16165 1125 16195
rect 1155 16165 1160 16195
rect 1120 16035 1160 16165
rect 1120 16005 1125 16035
rect 1155 16005 1160 16035
rect 1120 15875 1160 16005
rect 1120 15845 1125 15875
rect 1155 15845 1160 15875
rect 1120 15715 1160 15845
rect 1120 15685 1125 15715
rect 1155 15685 1160 15715
rect 1120 15555 1160 15685
rect 1120 15525 1125 15555
rect 1155 15525 1160 15555
rect 1120 15395 1160 15525
rect 1120 15365 1125 15395
rect 1155 15365 1160 15395
rect 1120 15235 1160 15365
rect 1120 15205 1125 15235
rect 1155 15205 1160 15235
rect 1120 15200 1160 15205
rect 1200 16195 1240 16200
rect 1200 16165 1205 16195
rect 1235 16165 1240 16195
rect 1200 16035 1240 16165
rect 1200 16005 1205 16035
rect 1235 16005 1240 16035
rect 1200 15875 1240 16005
rect 1200 15845 1205 15875
rect 1235 15845 1240 15875
rect 1200 15715 1240 15845
rect 1200 15685 1205 15715
rect 1235 15685 1240 15715
rect 1200 15555 1240 15685
rect 1200 15525 1205 15555
rect 1235 15525 1240 15555
rect 1200 15395 1240 15525
rect 1200 15365 1205 15395
rect 1235 15365 1240 15395
rect 1200 15235 1240 15365
rect 1200 15205 1205 15235
rect 1235 15205 1240 15235
rect 1200 15200 1240 15205
rect 1280 16195 1320 16200
rect 1280 16165 1285 16195
rect 1315 16165 1320 16195
rect 1280 16035 1320 16165
rect 1280 16005 1285 16035
rect 1315 16005 1320 16035
rect 1280 15875 1320 16005
rect 1280 15845 1285 15875
rect 1315 15845 1320 15875
rect 1280 15715 1320 15845
rect 1280 15685 1285 15715
rect 1315 15685 1320 15715
rect 1280 15555 1320 15685
rect 1280 15525 1285 15555
rect 1315 15525 1320 15555
rect 1280 15395 1320 15525
rect 1280 15365 1285 15395
rect 1315 15365 1320 15395
rect 1280 15235 1320 15365
rect 1280 15205 1285 15235
rect 1315 15205 1320 15235
rect 1280 15200 1320 15205
rect 1360 16195 1400 16200
rect 1360 16165 1365 16195
rect 1395 16165 1400 16195
rect 1360 16035 1400 16165
rect 1360 16005 1365 16035
rect 1395 16005 1400 16035
rect 1360 15875 1400 16005
rect 1360 15845 1365 15875
rect 1395 15845 1400 15875
rect 1360 15715 1400 15845
rect 1360 15685 1365 15715
rect 1395 15685 1400 15715
rect 1360 15555 1400 15685
rect 1360 15525 1365 15555
rect 1395 15525 1400 15555
rect 1360 15395 1400 15525
rect 1360 15365 1365 15395
rect 1395 15365 1400 15395
rect 1360 15235 1400 15365
rect 1360 15205 1365 15235
rect 1395 15205 1400 15235
rect 1360 15200 1400 15205
rect 1440 16195 1480 16200
rect 1440 16165 1445 16195
rect 1475 16165 1480 16195
rect 1440 16035 1480 16165
rect 1440 16005 1445 16035
rect 1475 16005 1480 16035
rect 1440 15875 1480 16005
rect 1440 15845 1445 15875
rect 1475 15845 1480 15875
rect 1440 15715 1480 15845
rect 1440 15685 1445 15715
rect 1475 15685 1480 15715
rect 1440 15555 1480 15685
rect 1440 15525 1445 15555
rect 1475 15525 1480 15555
rect 1440 15395 1480 15525
rect 1440 15365 1445 15395
rect 1475 15365 1480 15395
rect 1440 15235 1480 15365
rect 1440 15205 1445 15235
rect 1475 15205 1480 15235
rect 1440 15200 1480 15205
rect 1520 16195 1560 16200
rect 1520 16165 1525 16195
rect 1555 16165 1560 16195
rect 1520 16035 1560 16165
rect 1520 16005 1525 16035
rect 1555 16005 1560 16035
rect 1520 15875 1560 16005
rect 1520 15845 1525 15875
rect 1555 15845 1560 15875
rect 1520 15715 1560 15845
rect 1520 15685 1525 15715
rect 1555 15685 1560 15715
rect 1520 15555 1560 15685
rect 1520 15525 1525 15555
rect 1555 15525 1560 15555
rect 1520 15395 1560 15525
rect 1520 15365 1525 15395
rect 1555 15365 1560 15395
rect 1520 15235 1560 15365
rect 1520 15205 1525 15235
rect 1555 15205 1560 15235
rect 1520 15200 1560 15205
rect 1600 16195 1640 16200
rect 1600 16165 1605 16195
rect 1635 16165 1640 16195
rect 1600 16035 1640 16165
rect 1600 16005 1605 16035
rect 1635 16005 1640 16035
rect 1600 15875 1640 16005
rect 1600 15845 1605 15875
rect 1635 15845 1640 15875
rect 1600 15715 1640 15845
rect 1600 15685 1605 15715
rect 1635 15685 1640 15715
rect 1600 15555 1640 15685
rect 1600 15525 1605 15555
rect 1635 15525 1640 15555
rect 1600 15395 1640 15525
rect 1600 15365 1605 15395
rect 1635 15365 1640 15395
rect 1600 15235 1640 15365
rect 1600 15205 1605 15235
rect 1635 15205 1640 15235
rect 1600 15200 1640 15205
rect 1680 16195 1720 16200
rect 1680 16165 1685 16195
rect 1715 16165 1720 16195
rect 1680 16035 1720 16165
rect 1680 16005 1685 16035
rect 1715 16005 1720 16035
rect 1680 15875 1720 16005
rect 1680 15845 1685 15875
rect 1715 15845 1720 15875
rect 1680 15715 1720 15845
rect 1680 15685 1685 15715
rect 1715 15685 1720 15715
rect 1680 15555 1720 15685
rect 1680 15525 1685 15555
rect 1715 15525 1720 15555
rect 1680 15395 1720 15525
rect 1680 15365 1685 15395
rect 1715 15365 1720 15395
rect 1680 15235 1720 15365
rect 1680 15205 1685 15235
rect 1715 15205 1720 15235
rect 1680 15200 1720 15205
rect 1760 16195 1800 16200
rect 1760 16165 1765 16195
rect 1795 16165 1800 16195
rect 1760 16035 1800 16165
rect 1760 16005 1765 16035
rect 1795 16005 1800 16035
rect 1760 15875 1800 16005
rect 1760 15845 1765 15875
rect 1795 15845 1800 15875
rect 1760 15715 1800 15845
rect 1760 15685 1765 15715
rect 1795 15685 1800 15715
rect 1760 15555 1800 15685
rect 1760 15525 1765 15555
rect 1795 15525 1800 15555
rect 1760 15395 1800 15525
rect 1760 15365 1765 15395
rect 1795 15365 1800 15395
rect 1760 15235 1800 15365
rect 1760 15205 1765 15235
rect 1795 15205 1800 15235
rect 1760 15200 1800 15205
rect 1840 16195 1880 16200
rect 1840 16165 1845 16195
rect 1875 16165 1880 16195
rect 1840 16035 1880 16165
rect 1840 16005 1845 16035
rect 1875 16005 1880 16035
rect 1840 15875 1880 16005
rect 1840 15845 1845 15875
rect 1875 15845 1880 15875
rect 1840 15715 1880 15845
rect 1840 15685 1845 15715
rect 1875 15685 1880 15715
rect 1840 15555 1880 15685
rect 1840 15525 1845 15555
rect 1875 15525 1880 15555
rect 1840 15395 1880 15525
rect 1840 15365 1845 15395
rect 1875 15365 1880 15395
rect 1840 15235 1880 15365
rect 1840 15205 1845 15235
rect 1875 15205 1880 15235
rect 1840 15200 1880 15205
rect 1920 16195 1960 16200
rect 1920 16165 1925 16195
rect 1955 16165 1960 16195
rect 1920 16035 1960 16165
rect 1920 16005 1925 16035
rect 1955 16005 1960 16035
rect 1920 15875 1960 16005
rect 1920 15845 1925 15875
rect 1955 15845 1960 15875
rect 1920 15715 1960 15845
rect 1920 15685 1925 15715
rect 1955 15685 1960 15715
rect 1920 15555 1960 15685
rect 1920 15525 1925 15555
rect 1955 15525 1960 15555
rect 1920 15395 1960 15525
rect 1920 15365 1925 15395
rect 1955 15365 1960 15395
rect 1920 15235 1960 15365
rect 1920 15205 1925 15235
rect 1955 15205 1960 15235
rect 1920 15200 1960 15205
rect 2000 16195 2040 16200
rect 2000 16165 2005 16195
rect 2035 16165 2040 16195
rect 2000 16035 2040 16165
rect 2000 16005 2005 16035
rect 2035 16005 2040 16035
rect 2000 15875 2040 16005
rect 2000 15845 2005 15875
rect 2035 15845 2040 15875
rect 2000 15715 2040 15845
rect 2000 15685 2005 15715
rect 2035 15685 2040 15715
rect 2000 15555 2040 15685
rect 2000 15525 2005 15555
rect 2035 15525 2040 15555
rect 2000 15395 2040 15525
rect 2000 15365 2005 15395
rect 2035 15365 2040 15395
rect 2000 15235 2040 15365
rect 2000 15205 2005 15235
rect 2035 15205 2040 15235
rect 2000 15200 2040 15205
rect 2080 16195 2120 16200
rect 2080 16165 2085 16195
rect 2115 16165 2120 16195
rect 2080 16035 2120 16165
rect 2080 16005 2085 16035
rect 2115 16005 2120 16035
rect 2080 15875 2120 16005
rect 2080 15845 2085 15875
rect 2115 15845 2120 15875
rect 2080 15715 2120 15845
rect 2080 15685 2085 15715
rect 2115 15685 2120 15715
rect 2080 15555 2120 15685
rect 2080 15525 2085 15555
rect 2115 15525 2120 15555
rect 2080 15395 2120 15525
rect 2080 15365 2085 15395
rect 2115 15365 2120 15395
rect 2080 15235 2120 15365
rect 2080 15205 2085 15235
rect 2115 15205 2120 15235
rect 2080 15200 2120 15205
rect 2160 16195 2200 16200
rect 2160 16165 2165 16195
rect 2195 16165 2200 16195
rect 2160 16035 2200 16165
rect 2160 16005 2165 16035
rect 2195 16005 2200 16035
rect 2160 15875 2200 16005
rect 2160 15845 2165 15875
rect 2195 15845 2200 15875
rect 2160 15715 2200 15845
rect 2160 15685 2165 15715
rect 2195 15685 2200 15715
rect 2160 15555 2200 15685
rect 2160 15525 2165 15555
rect 2195 15525 2200 15555
rect 2160 15395 2200 15525
rect 2160 15365 2165 15395
rect 2195 15365 2200 15395
rect 2160 15235 2200 15365
rect 2160 15205 2165 15235
rect 2195 15205 2200 15235
rect 2160 15200 2200 15205
rect 2240 16195 2280 16200
rect 2240 16165 2245 16195
rect 2275 16165 2280 16195
rect 2240 16035 2280 16165
rect 2240 16005 2245 16035
rect 2275 16005 2280 16035
rect 2240 15875 2280 16005
rect 2240 15845 2245 15875
rect 2275 15845 2280 15875
rect 2240 15715 2280 15845
rect 2240 15685 2245 15715
rect 2275 15685 2280 15715
rect 2240 15555 2280 15685
rect 2240 15525 2245 15555
rect 2275 15525 2280 15555
rect 2240 15395 2280 15525
rect 2240 15365 2245 15395
rect 2275 15365 2280 15395
rect 2240 15235 2280 15365
rect 2240 15205 2245 15235
rect 2275 15205 2280 15235
rect 2240 15200 2280 15205
rect 2320 16195 2360 16200
rect 2320 16165 2325 16195
rect 2355 16165 2360 16195
rect 2320 16035 2360 16165
rect 2320 16005 2325 16035
rect 2355 16005 2360 16035
rect 2320 15875 2360 16005
rect 2320 15845 2325 15875
rect 2355 15845 2360 15875
rect 2320 15715 2360 15845
rect 2320 15685 2325 15715
rect 2355 15685 2360 15715
rect 2320 15555 2360 15685
rect 2320 15525 2325 15555
rect 2355 15525 2360 15555
rect 2320 15395 2360 15525
rect 2320 15365 2325 15395
rect 2355 15365 2360 15395
rect 2320 15235 2360 15365
rect 2320 15205 2325 15235
rect 2355 15205 2360 15235
rect 2320 15200 2360 15205
rect 2400 16195 2440 16200
rect 2400 16165 2405 16195
rect 2435 16165 2440 16195
rect 2400 16035 2440 16165
rect 2400 16005 2405 16035
rect 2435 16005 2440 16035
rect 2400 15875 2440 16005
rect 2400 15845 2405 15875
rect 2435 15845 2440 15875
rect 2400 15715 2440 15845
rect 2400 15685 2405 15715
rect 2435 15685 2440 15715
rect 2400 15555 2440 15685
rect 2400 15525 2405 15555
rect 2435 15525 2440 15555
rect 2400 15395 2440 15525
rect 2400 15365 2405 15395
rect 2435 15365 2440 15395
rect 2400 15235 2440 15365
rect 2400 15205 2405 15235
rect 2435 15205 2440 15235
rect 2400 15200 2440 15205
rect 2480 16195 2520 16200
rect 2480 16165 2485 16195
rect 2515 16165 2520 16195
rect 2480 16035 2520 16165
rect 2480 16005 2485 16035
rect 2515 16005 2520 16035
rect 2480 15875 2520 16005
rect 2480 15845 2485 15875
rect 2515 15845 2520 15875
rect 2480 15715 2520 15845
rect 2480 15685 2485 15715
rect 2515 15685 2520 15715
rect 2480 15555 2520 15685
rect 2480 15525 2485 15555
rect 2515 15525 2520 15555
rect 2480 15395 2520 15525
rect 2480 15365 2485 15395
rect 2515 15365 2520 15395
rect 2480 15235 2520 15365
rect 2480 15205 2485 15235
rect 2515 15205 2520 15235
rect 2480 15200 2520 15205
rect 2560 16195 2600 16200
rect 2560 16165 2565 16195
rect 2595 16165 2600 16195
rect 2560 16035 2600 16165
rect 2560 16005 2565 16035
rect 2595 16005 2600 16035
rect 2560 15875 2600 16005
rect 2560 15845 2565 15875
rect 2595 15845 2600 15875
rect 2560 15715 2600 15845
rect 2560 15685 2565 15715
rect 2595 15685 2600 15715
rect 2560 15555 2600 15685
rect 2560 15525 2565 15555
rect 2595 15525 2600 15555
rect 2560 15395 2600 15525
rect 2560 15365 2565 15395
rect 2595 15365 2600 15395
rect 2560 15235 2600 15365
rect 2560 15205 2565 15235
rect 2595 15205 2600 15235
rect 2560 15200 2600 15205
rect 2640 16195 2680 16200
rect 2640 16165 2645 16195
rect 2675 16165 2680 16195
rect 2640 16035 2680 16165
rect 2640 16005 2645 16035
rect 2675 16005 2680 16035
rect 2640 15875 2680 16005
rect 2640 15845 2645 15875
rect 2675 15845 2680 15875
rect 2640 15715 2680 15845
rect 2640 15685 2645 15715
rect 2675 15685 2680 15715
rect 2640 15555 2680 15685
rect 2640 15525 2645 15555
rect 2675 15525 2680 15555
rect 2640 15395 2680 15525
rect 2640 15365 2645 15395
rect 2675 15365 2680 15395
rect 2640 15235 2680 15365
rect 2640 15205 2645 15235
rect 2675 15205 2680 15235
rect 2640 15200 2680 15205
rect 2720 16195 2760 16200
rect 2720 16165 2725 16195
rect 2755 16165 2760 16195
rect 2720 16035 2760 16165
rect 2720 16005 2725 16035
rect 2755 16005 2760 16035
rect 2720 15875 2760 16005
rect 2720 15845 2725 15875
rect 2755 15845 2760 15875
rect 2720 15715 2760 15845
rect 2720 15685 2725 15715
rect 2755 15685 2760 15715
rect 2720 15555 2760 15685
rect 2720 15525 2725 15555
rect 2755 15525 2760 15555
rect 2720 15395 2760 15525
rect 2720 15365 2725 15395
rect 2755 15365 2760 15395
rect 2720 15235 2760 15365
rect 2720 15205 2725 15235
rect 2755 15205 2760 15235
rect 2720 15200 2760 15205
rect 2800 16195 2840 16200
rect 2800 16165 2805 16195
rect 2835 16165 2840 16195
rect 2800 16035 2840 16165
rect 2800 16005 2805 16035
rect 2835 16005 2840 16035
rect 2800 15875 2840 16005
rect 2800 15845 2805 15875
rect 2835 15845 2840 15875
rect 2800 15715 2840 15845
rect 2800 15685 2805 15715
rect 2835 15685 2840 15715
rect 2800 15555 2840 15685
rect 2800 15525 2805 15555
rect 2835 15525 2840 15555
rect 2800 15395 2840 15525
rect 2800 15365 2805 15395
rect 2835 15365 2840 15395
rect 2800 15235 2840 15365
rect 2800 15205 2805 15235
rect 2835 15205 2840 15235
rect 2800 15200 2840 15205
rect 2880 16195 2920 16200
rect 2880 16165 2885 16195
rect 2915 16165 2920 16195
rect 2880 16035 2920 16165
rect 2880 16005 2885 16035
rect 2915 16005 2920 16035
rect 2880 15875 2920 16005
rect 2880 15845 2885 15875
rect 2915 15845 2920 15875
rect 2880 15715 2920 15845
rect 2880 15685 2885 15715
rect 2915 15685 2920 15715
rect 2880 15555 2920 15685
rect 2880 15525 2885 15555
rect 2915 15525 2920 15555
rect 2880 15395 2920 15525
rect 2880 15365 2885 15395
rect 2915 15365 2920 15395
rect 2880 15235 2920 15365
rect 2880 15205 2885 15235
rect 2915 15205 2920 15235
rect 2880 15200 2920 15205
rect 2960 16195 3000 16200
rect 2960 16165 2965 16195
rect 2995 16165 3000 16195
rect 2960 16035 3000 16165
rect 2960 16005 2965 16035
rect 2995 16005 3000 16035
rect 2960 15875 3000 16005
rect 2960 15845 2965 15875
rect 2995 15845 3000 15875
rect 2960 15715 3000 15845
rect 2960 15685 2965 15715
rect 2995 15685 3000 15715
rect 2960 15555 3000 15685
rect 2960 15525 2965 15555
rect 2995 15525 3000 15555
rect 2960 15395 3000 15525
rect 2960 15365 2965 15395
rect 2995 15365 3000 15395
rect 2960 15235 3000 15365
rect 2960 15205 2965 15235
rect 2995 15205 3000 15235
rect 2960 15200 3000 15205
rect 3040 16195 3080 16200
rect 3040 16165 3045 16195
rect 3075 16165 3080 16195
rect 3040 16035 3080 16165
rect 3040 16005 3045 16035
rect 3075 16005 3080 16035
rect 3040 15875 3080 16005
rect 3040 15845 3045 15875
rect 3075 15845 3080 15875
rect 3040 15715 3080 15845
rect 3040 15685 3045 15715
rect 3075 15685 3080 15715
rect 3040 15555 3080 15685
rect 3040 15525 3045 15555
rect 3075 15525 3080 15555
rect 3040 15395 3080 15525
rect 3040 15365 3045 15395
rect 3075 15365 3080 15395
rect 3040 15235 3080 15365
rect 3040 15205 3045 15235
rect 3075 15205 3080 15235
rect 3040 15200 3080 15205
rect 3120 16195 3160 16200
rect 3120 16165 3125 16195
rect 3155 16165 3160 16195
rect 3120 16035 3160 16165
rect 3120 16005 3125 16035
rect 3155 16005 3160 16035
rect 3120 15875 3160 16005
rect 3120 15845 3125 15875
rect 3155 15845 3160 15875
rect 3120 15715 3160 15845
rect 3120 15685 3125 15715
rect 3155 15685 3160 15715
rect 3120 15555 3160 15685
rect 3120 15525 3125 15555
rect 3155 15525 3160 15555
rect 3120 15395 3160 15525
rect 3120 15365 3125 15395
rect 3155 15365 3160 15395
rect 3120 15235 3160 15365
rect 3120 15205 3125 15235
rect 3155 15205 3160 15235
rect 3120 15200 3160 15205
rect 3200 16195 3240 16200
rect 3200 16165 3205 16195
rect 3235 16165 3240 16195
rect 3200 16035 3240 16165
rect 3200 16005 3205 16035
rect 3235 16005 3240 16035
rect 3200 15875 3240 16005
rect 3200 15845 3205 15875
rect 3235 15845 3240 15875
rect 3200 15715 3240 15845
rect 3200 15685 3205 15715
rect 3235 15685 3240 15715
rect 3200 15555 3240 15685
rect 3200 15525 3205 15555
rect 3235 15525 3240 15555
rect 3200 15395 3240 15525
rect 3200 15365 3205 15395
rect 3235 15365 3240 15395
rect 3200 15235 3240 15365
rect 3200 15205 3205 15235
rect 3235 15205 3240 15235
rect 3200 15200 3240 15205
rect 3280 16195 3320 16200
rect 3280 16165 3285 16195
rect 3315 16165 3320 16195
rect 3280 16035 3320 16165
rect 3280 16005 3285 16035
rect 3315 16005 3320 16035
rect 3280 15875 3320 16005
rect 3280 15845 3285 15875
rect 3315 15845 3320 15875
rect 3280 15715 3320 15845
rect 3280 15685 3285 15715
rect 3315 15685 3320 15715
rect 3280 15555 3320 15685
rect 3280 15525 3285 15555
rect 3315 15525 3320 15555
rect 3280 15395 3320 15525
rect 3280 15365 3285 15395
rect 3315 15365 3320 15395
rect 3280 15235 3320 15365
rect 3280 15205 3285 15235
rect 3315 15205 3320 15235
rect 3280 15200 3320 15205
rect 3360 16195 3400 16200
rect 3360 16165 3365 16195
rect 3395 16165 3400 16195
rect 3360 16035 3400 16165
rect 3360 16005 3365 16035
rect 3395 16005 3400 16035
rect 3360 15875 3400 16005
rect 3360 15845 3365 15875
rect 3395 15845 3400 15875
rect 3360 15715 3400 15845
rect 3360 15685 3365 15715
rect 3395 15685 3400 15715
rect 3360 15555 3400 15685
rect 3360 15525 3365 15555
rect 3395 15525 3400 15555
rect 3360 15395 3400 15525
rect 3360 15365 3365 15395
rect 3395 15365 3400 15395
rect 3360 15235 3400 15365
rect 3360 15205 3365 15235
rect 3395 15205 3400 15235
rect 3360 15200 3400 15205
rect 3440 16195 3480 16200
rect 3440 16165 3445 16195
rect 3475 16165 3480 16195
rect 3440 16035 3480 16165
rect 3440 16005 3445 16035
rect 3475 16005 3480 16035
rect 3440 15875 3480 16005
rect 3440 15845 3445 15875
rect 3475 15845 3480 15875
rect 3440 15715 3480 15845
rect 3440 15685 3445 15715
rect 3475 15685 3480 15715
rect 3440 15555 3480 15685
rect 3440 15525 3445 15555
rect 3475 15525 3480 15555
rect 3440 15395 3480 15525
rect 3440 15365 3445 15395
rect 3475 15365 3480 15395
rect 3440 15235 3480 15365
rect 3440 15205 3445 15235
rect 3475 15205 3480 15235
rect 3440 15200 3480 15205
rect 3520 16195 3560 16200
rect 3520 16165 3525 16195
rect 3555 16165 3560 16195
rect 3520 16035 3560 16165
rect 3520 16005 3525 16035
rect 3555 16005 3560 16035
rect 3520 15875 3560 16005
rect 3520 15845 3525 15875
rect 3555 15845 3560 15875
rect 3520 15715 3560 15845
rect 3520 15685 3525 15715
rect 3555 15685 3560 15715
rect 3520 15555 3560 15685
rect 3520 15525 3525 15555
rect 3555 15525 3560 15555
rect 3520 15395 3560 15525
rect 3520 15365 3525 15395
rect 3555 15365 3560 15395
rect 3520 15235 3560 15365
rect 3520 15205 3525 15235
rect 3555 15205 3560 15235
rect 3520 15200 3560 15205
rect 3600 16195 3640 16200
rect 3600 16165 3605 16195
rect 3635 16165 3640 16195
rect 3600 16035 3640 16165
rect 3600 16005 3605 16035
rect 3635 16005 3640 16035
rect 3600 15875 3640 16005
rect 3600 15845 3605 15875
rect 3635 15845 3640 15875
rect 3600 15715 3640 15845
rect 3600 15685 3605 15715
rect 3635 15685 3640 15715
rect 3600 15555 3640 15685
rect 3600 15525 3605 15555
rect 3635 15525 3640 15555
rect 3600 15395 3640 15525
rect 3600 15365 3605 15395
rect 3635 15365 3640 15395
rect 3600 15235 3640 15365
rect 3600 15205 3605 15235
rect 3635 15205 3640 15235
rect 3600 15200 3640 15205
rect 3680 16195 3720 16200
rect 3680 16165 3685 16195
rect 3715 16165 3720 16195
rect 3680 16035 3720 16165
rect 3680 16005 3685 16035
rect 3715 16005 3720 16035
rect 3680 15875 3720 16005
rect 3680 15845 3685 15875
rect 3715 15845 3720 15875
rect 3680 15715 3720 15845
rect 3680 15685 3685 15715
rect 3715 15685 3720 15715
rect 3680 15555 3720 15685
rect 3680 15525 3685 15555
rect 3715 15525 3720 15555
rect 3680 15395 3720 15525
rect 3680 15365 3685 15395
rect 3715 15365 3720 15395
rect 3680 15235 3720 15365
rect 3680 15205 3685 15235
rect 3715 15205 3720 15235
rect 3680 15200 3720 15205
rect 3760 16195 3800 16200
rect 3760 16165 3765 16195
rect 3795 16165 3800 16195
rect 3760 16035 3800 16165
rect 3760 16005 3765 16035
rect 3795 16005 3800 16035
rect 3760 15875 3800 16005
rect 3760 15845 3765 15875
rect 3795 15845 3800 15875
rect 3760 15715 3800 15845
rect 3760 15685 3765 15715
rect 3795 15685 3800 15715
rect 3760 15555 3800 15685
rect 3760 15525 3765 15555
rect 3795 15525 3800 15555
rect 3760 15395 3800 15525
rect 3760 15365 3765 15395
rect 3795 15365 3800 15395
rect 3760 15235 3800 15365
rect 3760 15205 3765 15235
rect 3795 15205 3800 15235
rect 3760 15200 3800 15205
rect 3840 16195 3880 16200
rect 3840 16165 3845 16195
rect 3875 16165 3880 16195
rect 3840 16035 3880 16165
rect 3840 16005 3845 16035
rect 3875 16005 3880 16035
rect 3840 15875 3880 16005
rect 3840 15845 3845 15875
rect 3875 15845 3880 15875
rect 3840 15715 3880 15845
rect 3840 15685 3845 15715
rect 3875 15685 3880 15715
rect 3840 15555 3880 15685
rect 3840 15525 3845 15555
rect 3875 15525 3880 15555
rect 3840 15395 3880 15525
rect 3840 15365 3845 15395
rect 3875 15365 3880 15395
rect 3840 15235 3880 15365
rect 3840 15205 3845 15235
rect 3875 15205 3880 15235
rect 3840 15200 3880 15205
rect 3920 16195 3960 16200
rect 3920 16165 3925 16195
rect 3955 16165 3960 16195
rect 3920 16035 3960 16165
rect 3920 16005 3925 16035
rect 3955 16005 3960 16035
rect 3920 15875 3960 16005
rect 3920 15845 3925 15875
rect 3955 15845 3960 15875
rect 3920 15715 3960 15845
rect 3920 15685 3925 15715
rect 3955 15685 3960 15715
rect 3920 15555 3960 15685
rect 3920 15525 3925 15555
rect 3955 15525 3960 15555
rect 3920 15395 3960 15525
rect 3920 15365 3925 15395
rect 3955 15365 3960 15395
rect 3920 15235 3960 15365
rect 3920 15205 3925 15235
rect 3955 15205 3960 15235
rect 3920 15200 3960 15205
rect 4000 16195 4040 16200
rect 4000 16165 4005 16195
rect 4035 16165 4040 16195
rect 4000 16035 4040 16165
rect 4000 16005 4005 16035
rect 4035 16005 4040 16035
rect 4000 15875 4040 16005
rect 4000 15845 4005 15875
rect 4035 15845 4040 15875
rect 4000 15715 4040 15845
rect 4000 15685 4005 15715
rect 4035 15685 4040 15715
rect 4000 15555 4040 15685
rect 4000 15525 4005 15555
rect 4035 15525 4040 15555
rect 4000 15395 4040 15525
rect 4000 15365 4005 15395
rect 4035 15365 4040 15395
rect 4000 15235 4040 15365
rect 4000 15205 4005 15235
rect 4035 15205 4040 15235
rect 4000 15200 4040 15205
rect 4080 16195 4120 16200
rect 4080 16165 4085 16195
rect 4115 16165 4120 16195
rect 4080 16035 4120 16165
rect 4080 16005 4085 16035
rect 4115 16005 4120 16035
rect 4080 15875 4120 16005
rect 4080 15845 4085 15875
rect 4115 15845 4120 15875
rect 4080 15715 4120 15845
rect 4080 15685 4085 15715
rect 4115 15685 4120 15715
rect 4080 15555 4120 15685
rect 4080 15525 4085 15555
rect 4115 15525 4120 15555
rect 4080 15395 4120 15525
rect 4080 15365 4085 15395
rect 4115 15365 4120 15395
rect 4080 15235 4120 15365
rect 4080 15205 4085 15235
rect 4115 15205 4120 15235
rect 4080 15200 4120 15205
rect 4160 16195 4200 16200
rect 4160 16165 4165 16195
rect 4195 16165 4200 16195
rect 4160 16035 4200 16165
rect 4160 16005 4165 16035
rect 4195 16005 4200 16035
rect 4160 15875 4200 16005
rect 4160 15845 4165 15875
rect 4195 15845 4200 15875
rect 4160 15715 4200 15845
rect 4160 15685 4165 15715
rect 4195 15685 4200 15715
rect 4160 15555 4200 15685
rect 4160 15525 4165 15555
rect 4195 15525 4200 15555
rect 4160 15395 4200 15525
rect 4160 15365 4165 15395
rect 4195 15365 4200 15395
rect 4160 15235 4200 15365
rect 4160 15205 4165 15235
rect 4195 15205 4200 15235
rect 4160 15200 4200 15205
rect 0 15155 40 15160
rect 0 15125 5 15155
rect 35 15125 40 15155
rect 0 14995 40 15125
rect 0 14965 5 14995
rect 35 14965 40 14995
rect 0 14960 40 14965
rect 80 15155 120 15160
rect 80 15125 85 15155
rect 115 15125 120 15155
rect 80 14995 120 15125
rect 80 14965 85 14995
rect 115 14965 120 14995
rect 80 14960 120 14965
rect 160 15155 200 15160
rect 160 15125 165 15155
rect 195 15125 200 15155
rect 160 14995 200 15125
rect 160 14965 165 14995
rect 195 14965 200 14995
rect 160 14960 200 14965
rect 240 15155 280 15160
rect 240 15125 245 15155
rect 275 15125 280 15155
rect 240 14995 280 15125
rect 240 14965 245 14995
rect 275 14965 280 14995
rect 240 14960 280 14965
rect 320 15155 360 15160
rect 320 15125 325 15155
rect 355 15125 360 15155
rect 320 14995 360 15125
rect 320 14965 325 14995
rect 355 14965 360 14995
rect 320 14960 360 14965
rect 400 15155 440 15160
rect 400 15125 405 15155
rect 435 15125 440 15155
rect 400 14995 440 15125
rect 400 14965 405 14995
rect 435 14965 440 14995
rect 400 14960 440 14965
rect 480 15155 520 15160
rect 480 15125 485 15155
rect 515 15125 520 15155
rect 480 14995 520 15125
rect 480 14965 485 14995
rect 515 14965 520 14995
rect 480 14960 520 14965
rect 560 15155 600 15160
rect 560 15125 565 15155
rect 595 15125 600 15155
rect 560 14995 600 15125
rect 560 14965 565 14995
rect 595 14965 600 14995
rect 560 14960 600 14965
rect 640 15155 680 15160
rect 640 15125 645 15155
rect 675 15125 680 15155
rect 640 14995 680 15125
rect 640 14965 645 14995
rect 675 14965 680 14995
rect 640 14960 680 14965
rect 720 15155 760 15160
rect 720 15125 725 15155
rect 755 15125 760 15155
rect 720 14995 760 15125
rect 720 14965 725 14995
rect 755 14965 760 14995
rect 720 14960 760 14965
rect 800 15155 840 15160
rect 800 15125 805 15155
rect 835 15125 840 15155
rect 800 14995 840 15125
rect 800 14965 805 14995
rect 835 14965 840 14995
rect 800 14960 840 14965
rect 880 15155 920 15160
rect 880 15125 885 15155
rect 915 15125 920 15155
rect 880 14995 920 15125
rect 880 14965 885 14995
rect 915 14965 920 14995
rect 880 14960 920 14965
rect 960 15155 1000 15160
rect 960 15125 965 15155
rect 995 15125 1000 15155
rect 960 14995 1000 15125
rect 960 14965 965 14995
rect 995 14965 1000 14995
rect 960 14960 1000 14965
rect 1040 15155 1080 15160
rect 1040 15125 1045 15155
rect 1075 15125 1080 15155
rect 1040 14995 1080 15125
rect 1040 14965 1045 14995
rect 1075 14965 1080 14995
rect 1040 14960 1080 14965
rect 1120 15155 1160 15160
rect 1120 15125 1125 15155
rect 1155 15125 1160 15155
rect 1120 14995 1160 15125
rect 1120 14965 1125 14995
rect 1155 14965 1160 14995
rect 1120 14960 1160 14965
rect 1200 15155 1240 15160
rect 1200 15125 1205 15155
rect 1235 15125 1240 15155
rect 1200 14995 1240 15125
rect 1200 14965 1205 14995
rect 1235 14965 1240 14995
rect 1200 14960 1240 14965
rect 1280 15155 1320 15160
rect 1280 15125 1285 15155
rect 1315 15125 1320 15155
rect 1280 14995 1320 15125
rect 1280 14965 1285 14995
rect 1315 14965 1320 14995
rect 1280 14960 1320 14965
rect 1360 15155 1400 15160
rect 1360 15125 1365 15155
rect 1395 15125 1400 15155
rect 1360 14995 1400 15125
rect 1360 14965 1365 14995
rect 1395 14965 1400 14995
rect 1360 14960 1400 14965
rect 1440 15155 1480 15160
rect 1440 15125 1445 15155
rect 1475 15125 1480 15155
rect 1440 14995 1480 15125
rect 1440 14965 1445 14995
rect 1475 14965 1480 14995
rect 1440 14960 1480 14965
rect 1520 15155 1560 15160
rect 1520 15125 1525 15155
rect 1555 15125 1560 15155
rect 1520 14995 1560 15125
rect 1520 14965 1525 14995
rect 1555 14965 1560 14995
rect 1520 14960 1560 14965
rect 1600 15155 1640 15160
rect 1600 15125 1605 15155
rect 1635 15125 1640 15155
rect 1600 14995 1640 15125
rect 1600 14965 1605 14995
rect 1635 14965 1640 14995
rect 1600 14960 1640 14965
rect 1680 15155 1720 15160
rect 1680 15125 1685 15155
rect 1715 15125 1720 15155
rect 1680 14995 1720 15125
rect 1680 14965 1685 14995
rect 1715 14965 1720 14995
rect 1680 14960 1720 14965
rect 1760 15155 1800 15160
rect 1760 15125 1765 15155
rect 1795 15125 1800 15155
rect 1760 14995 1800 15125
rect 1760 14965 1765 14995
rect 1795 14965 1800 14995
rect 1760 14960 1800 14965
rect 1840 15155 1880 15160
rect 1840 15125 1845 15155
rect 1875 15125 1880 15155
rect 1840 14995 1880 15125
rect 1840 14965 1845 14995
rect 1875 14965 1880 14995
rect 1840 14960 1880 14965
rect 1920 15155 1960 15160
rect 1920 15125 1925 15155
rect 1955 15125 1960 15155
rect 1920 14995 1960 15125
rect 1920 14965 1925 14995
rect 1955 14965 1960 14995
rect 1920 14960 1960 14965
rect 2000 15155 2040 15160
rect 2000 15125 2005 15155
rect 2035 15125 2040 15155
rect 2000 14995 2040 15125
rect 2000 14965 2005 14995
rect 2035 14965 2040 14995
rect 2000 14960 2040 14965
rect 2080 15155 2120 15160
rect 2080 15125 2085 15155
rect 2115 15125 2120 15155
rect 2080 14995 2120 15125
rect 2080 14965 2085 14995
rect 2115 14965 2120 14995
rect 2080 14960 2120 14965
rect 2160 15155 2200 15160
rect 2160 15125 2165 15155
rect 2195 15125 2200 15155
rect 2160 14995 2200 15125
rect 2160 14965 2165 14995
rect 2195 14965 2200 14995
rect 2160 14960 2200 14965
rect 2240 15155 2280 15160
rect 2240 15125 2245 15155
rect 2275 15125 2280 15155
rect 2240 14995 2280 15125
rect 2240 14965 2245 14995
rect 2275 14965 2280 14995
rect 2240 14960 2280 14965
rect 2320 15155 2360 15160
rect 2320 15125 2325 15155
rect 2355 15125 2360 15155
rect 2320 14995 2360 15125
rect 2320 14965 2325 14995
rect 2355 14965 2360 14995
rect 2320 14960 2360 14965
rect 2400 15155 2440 15160
rect 2400 15125 2405 15155
rect 2435 15125 2440 15155
rect 2400 14995 2440 15125
rect 2400 14965 2405 14995
rect 2435 14965 2440 14995
rect 2400 14960 2440 14965
rect 2480 15155 2520 15160
rect 2480 15125 2485 15155
rect 2515 15125 2520 15155
rect 2480 14995 2520 15125
rect 2480 14965 2485 14995
rect 2515 14965 2520 14995
rect 2480 14960 2520 14965
rect 2560 15155 2600 15160
rect 2560 15125 2565 15155
rect 2595 15125 2600 15155
rect 2560 14995 2600 15125
rect 2560 14965 2565 14995
rect 2595 14965 2600 14995
rect 2560 14960 2600 14965
rect 2640 15155 2680 15160
rect 2640 15125 2645 15155
rect 2675 15125 2680 15155
rect 2640 14995 2680 15125
rect 2640 14965 2645 14995
rect 2675 14965 2680 14995
rect 2640 14960 2680 14965
rect 2720 15155 2760 15160
rect 2720 15125 2725 15155
rect 2755 15125 2760 15155
rect 2720 14995 2760 15125
rect 2720 14965 2725 14995
rect 2755 14965 2760 14995
rect 2720 14960 2760 14965
rect 2800 15155 2840 15160
rect 2800 15125 2805 15155
rect 2835 15125 2840 15155
rect 2800 14995 2840 15125
rect 2800 14965 2805 14995
rect 2835 14965 2840 14995
rect 2800 14960 2840 14965
rect 2880 15155 2920 15160
rect 2880 15125 2885 15155
rect 2915 15125 2920 15155
rect 2880 14995 2920 15125
rect 2880 14965 2885 14995
rect 2915 14965 2920 14995
rect 2880 14960 2920 14965
rect 2960 15155 3000 15160
rect 2960 15125 2965 15155
rect 2995 15125 3000 15155
rect 2960 14995 3000 15125
rect 2960 14965 2965 14995
rect 2995 14965 3000 14995
rect 2960 14960 3000 14965
rect 3040 15155 3080 15160
rect 3040 15125 3045 15155
rect 3075 15125 3080 15155
rect 3040 14995 3080 15125
rect 3040 14965 3045 14995
rect 3075 14965 3080 14995
rect 3040 14960 3080 14965
rect 3120 15155 3160 15160
rect 3120 15125 3125 15155
rect 3155 15125 3160 15155
rect 3120 14995 3160 15125
rect 3120 14965 3125 14995
rect 3155 14965 3160 14995
rect 3120 14960 3160 14965
rect 3200 15155 3240 15160
rect 3200 15125 3205 15155
rect 3235 15125 3240 15155
rect 3200 14995 3240 15125
rect 3200 14965 3205 14995
rect 3235 14965 3240 14995
rect 3200 14960 3240 14965
rect 3280 15155 3320 15160
rect 3280 15125 3285 15155
rect 3315 15125 3320 15155
rect 3280 14995 3320 15125
rect 3280 14965 3285 14995
rect 3315 14965 3320 14995
rect 3280 14960 3320 14965
rect 3360 15155 3400 15160
rect 3360 15125 3365 15155
rect 3395 15125 3400 15155
rect 3360 14995 3400 15125
rect 3360 14965 3365 14995
rect 3395 14965 3400 14995
rect 3360 14960 3400 14965
rect 3440 15155 3480 15160
rect 3440 15125 3445 15155
rect 3475 15125 3480 15155
rect 3440 14995 3480 15125
rect 3440 14965 3445 14995
rect 3475 14965 3480 14995
rect 3440 14960 3480 14965
rect 3520 15155 3560 15160
rect 3520 15125 3525 15155
rect 3555 15125 3560 15155
rect 3520 14995 3560 15125
rect 3520 14965 3525 14995
rect 3555 14965 3560 14995
rect 3520 14960 3560 14965
rect 3600 15155 3640 15160
rect 3600 15125 3605 15155
rect 3635 15125 3640 15155
rect 3600 14995 3640 15125
rect 3600 14965 3605 14995
rect 3635 14965 3640 14995
rect 3600 14960 3640 14965
rect 3680 15155 3720 15160
rect 3680 15125 3685 15155
rect 3715 15125 3720 15155
rect 3680 14995 3720 15125
rect 3680 14965 3685 14995
rect 3715 14965 3720 14995
rect 3680 14960 3720 14965
rect 3760 15155 3800 15160
rect 3760 15125 3765 15155
rect 3795 15125 3800 15155
rect 3760 14995 3800 15125
rect 3760 14965 3765 14995
rect 3795 14965 3800 14995
rect 3760 14960 3800 14965
rect 3840 15155 3880 15160
rect 3840 15125 3845 15155
rect 3875 15125 3880 15155
rect 3840 14995 3880 15125
rect 3840 14965 3845 14995
rect 3875 14965 3880 14995
rect 3840 14960 3880 14965
rect 3920 15155 3960 15160
rect 3920 15125 3925 15155
rect 3955 15125 3960 15155
rect 3920 14995 3960 15125
rect 3920 14965 3925 14995
rect 3955 14965 3960 14995
rect 3920 14960 3960 14965
rect 4000 15155 4040 15160
rect 4000 15125 4005 15155
rect 4035 15125 4040 15155
rect 4000 14995 4040 15125
rect 4000 14965 4005 14995
rect 4035 14965 4040 14995
rect 4000 14960 4040 14965
rect 4080 15155 4120 15160
rect 4080 15125 4085 15155
rect 4115 15125 4120 15155
rect 4080 14995 4120 15125
rect 4080 14965 4085 14995
rect 4115 14965 4120 14995
rect 4080 14960 4120 14965
rect 4160 15155 4200 15160
rect 4160 15125 4165 15155
rect 4195 15125 4200 15155
rect 4160 14995 4200 15125
rect 4160 14965 4165 14995
rect 4195 14965 4200 14995
rect 4160 14960 4200 14965
rect 0 14915 40 14920
rect 0 14885 5 14915
rect 35 14885 40 14915
rect 0 14755 40 14885
rect 0 14725 5 14755
rect 35 14725 40 14755
rect 0 14720 40 14725
rect 80 14915 120 14920
rect 80 14885 85 14915
rect 115 14885 120 14915
rect 80 14755 120 14885
rect 80 14725 85 14755
rect 115 14725 120 14755
rect 80 14720 120 14725
rect 160 14915 200 14920
rect 160 14885 165 14915
rect 195 14885 200 14915
rect 160 14755 200 14885
rect 160 14725 165 14755
rect 195 14725 200 14755
rect 160 14720 200 14725
rect 240 14915 280 14920
rect 240 14885 245 14915
rect 275 14885 280 14915
rect 240 14755 280 14885
rect 240 14725 245 14755
rect 275 14725 280 14755
rect 240 14720 280 14725
rect 320 14915 360 14920
rect 320 14885 325 14915
rect 355 14885 360 14915
rect 320 14755 360 14885
rect 320 14725 325 14755
rect 355 14725 360 14755
rect 320 14720 360 14725
rect 400 14915 440 14920
rect 400 14885 405 14915
rect 435 14885 440 14915
rect 400 14755 440 14885
rect 400 14725 405 14755
rect 435 14725 440 14755
rect 400 14720 440 14725
rect 480 14915 520 14920
rect 480 14885 485 14915
rect 515 14885 520 14915
rect 480 14755 520 14885
rect 480 14725 485 14755
rect 515 14725 520 14755
rect 480 14720 520 14725
rect 560 14915 600 14920
rect 560 14885 565 14915
rect 595 14885 600 14915
rect 560 14755 600 14885
rect 560 14725 565 14755
rect 595 14725 600 14755
rect 560 14720 600 14725
rect 640 14915 680 14920
rect 640 14885 645 14915
rect 675 14885 680 14915
rect 640 14755 680 14885
rect 640 14725 645 14755
rect 675 14725 680 14755
rect 640 14720 680 14725
rect 720 14915 760 14920
rect 720 14885 725 14915
rect 755 14885 760 14915
rect 720 14755 760 14885
rect 720 14725 725 14755
rect 755 14725 760 14755
rect 720 14720 760 14725
rect 800 14915 840 14920
rect 800 14885 805 14915
rect 835 14885 840 14915
rect 800 14755 840 14885
rect 800 14725 805 14755
rect 835 14725 840 14755
rect 800 14720 840 14725
rect 880 14915 920 14920
rect 880 14885 885 14915
rect 915 14885 920 14915
rect 880 14755 920 14885
rect 880 14725 885 14755
rect 915 14725 920 14755
rect 880 14720 920 14725
rect 960 14915 1000 14920
rect 960 14885 965 14915
rect 995 14885 1000 14915
rect 960 14755 1000 14885
rect 960 14725 965 14755
rect 995 14725 1000 14755
rect 960 14720 1000 14725
rect 1040 14915 1080 14920
rect 1040 14885 1045 14915
rect 1075 14885 1080 14915
rect 1040 14755 1080 14885
rect 1040 14725 1045 14755
rect 1075 14725 1080 14755
rect 1040 14720 1080 14725
rect 1120 14915 1160 14920
rect 1120 14885 1125 14915
rect 1155 14885 1160 14915
rect 1120 14755 1160 14885
rect 1120 14725 1125 14755
rect 1155 14725 1160 14755
rect 1120 14720 1160 14725
rect 1200 14915 1240 14920
rect 1200 14885 1205 14915
rect 1235 14885 1240 14915
rect 1200 14755 1240 14885
rect 1200 14725 1205 14755
rect 1235 14725 1240 14755
rect 1200 14720 1240 14725
rect 1280 14915 1320 14920
rect 1280 14885 1285 14915
rect 1315 14885 1320 14915
rect 1280 14755 1320 14885
rect 1280 14725 1285 14755
rect 1315 14725 1320 14755
rect 1280 14720 1320 14725
rect 1360 14915 1400 14920
rect 1360 14885 1365 14915
rect 1395 14885 1400 14915
rect 1360 14755 1400 14885
rect 1360 14725 1365 14755
rect 1395 14725 1400 14755
rect 1360 14720 1400 14725
rect 1440 14915 1480 14920
rect 1440 14885 1445 14915
rect 1475 14885 1480 14915
rect 1440 14755 1480 14885
rect 1440 14725 1445 14755
rect 1475 14725 1480 14755
rect 1440 14720 1480 14725
rect 1520 14915 1560 14920
rect 1520 14885 1525 14915
rect 1555 14885 1560 14915
rect 1520 14755 1560 14885
rect 1520 14725 1525 14755
rect 1555 14725 1560 14755
rect 1520 14720 1560 14725
rect 1600 14915 1640 14920
rect 1600 14885 1605 14915
rect 1635 14885 1640 14915
rect 1600 14755 1640 14885
rect 1600 14725 1605 14755
rect 1635 14725 1640 14755
rect 1600 14720 1640 14725
rect 1680 14915 1720 14920
rect 1680 14885 1685 14915
rect 1715 14885 1720 14915
rect 1680 14755 1720 14885
rect 1680 14725 1685 14755
rect 1715 14725 1720 14755
rect 1680 14720 1720 14725
rect 1760 14915 1800 14920
rect 1760 14885 1765 14915
rect 1795 14885 1800 14915
rect 1760 14755 1800 14885
rect 1760 14725 1765 14755
rect 1795 14725 1800 14755
rect 1760 14720 1800 14725
rect 1840 14915 1880 14920
rect 1840 14885 1845 14915
rect 1875 14885 1880 14915
rect 1840 14755 1880 14885
rect 1840 14725 1845 14755
rect 1875 14725 1880 14755
rect 1840 14720 1880 14725
rect 1920 14915 1960 14920
rect 1920 14885 1925 14915
rect 1955 14885 1960 14915
rect 1920 14755 1960 14885
rect 1920 14725 1925 14755
rect 1955 14725 1960 14755
rect 1920 14720 1960 14725
rect 2000 14915 2040 14920
rect 2000 14885 2005 14915
rect 2035 14885 2040 14915
rect 2000 14755 2040 14885
rect 2000 14725 2005 14755
rect 2035 14725 2040 14755
rect 2000 14720 2040 14725
rect 2080 14915 2120 14920
rect 2080 14885 2085 14915
rect 2115 14885 2120 14915
rect 2080 14755 2120 14885
rect 2080 14725 2085 14755
rect 2115 14725 2120 14755
rect 2080 14720 2120 14725
rect 2160 14915 2200 14920
rect 2160 14885 2165 14915
rect 2195 14885 2200 14915
rect 2160 14755 2200 14885
rect 2160 14725 2165 14755
rect 2195 14725 2200 14755
rect 2160 14720 2200 14725
rect 2240 14915 2280 14920
rect 2240 14885 2245 14915
rect 2275 14885 2280 14915
rect 2240 14755 2280 14885
rect 2240 14725 2245 14755
rect 2275 14725 2280 14755
rect 2240 14720 2280 14725
rect 2320 14915 2360 14920
rect 2320 14885 2325 14915
rect 2355 14885 2360 14915
rect 2320 14755 2360 14885
rect 2320 14725 2325 14755
rect 2355 14725 2360 14755
rect 2320 14720 2360 14725
rect 2400 14915 2440 14920
rect 2400 14885 2405 14915
rect 2435 14885 2440 14915
rect 2400 14755 2440 14885
rect 2400 14725 2405 14755
rect 2435 14725 2440 14755
rect 2400 14720 2440 14725
rect 2480 14915 2520 14920
rect 2480 14885 2485 14915
rect 2515 14885 2520 14915
rect 2480 14755 2520 14885
rect 2480 14725 2485 14755
rect 2515 14725 2520 14755
rect 2480 14720 2520 14725
rect 2560 14915 2600 14920
rect 2560 14885 2565 14915
rect 2595 14885 2600 14915
rect 2560 14755 2600 14885
rect 2560 14725 2565 14755
rect 2595 14725 2600 14755
rect 2560 14720 2600 14725
rect 2640 14915 2680 14920
rect 2640 14885 2645 14915
rect 2675 14885 2680 14915
rect 2640 14755 2680 14885
rect 2640 14725 2645 14755
rect 2675 14725 2680 14755
rect 2640 14720 2680 14725
rect 2720 14915 2760 14920
rect 2720 14885 2725 14915
rect 2755 14885 2760 14915
rect 2720 14755 2760 14885
rect 2720 14725 2725 14755
rect 2755 14725 2760 14755
rect 2720 14720 2760 14725
rect 2800 14915 2840 14920
rect 2800 14885 2805 14915
rect 2835 14885 2840 14915
rect 2800 14755 2840 14885
rect 2800 14725 2805 14755
rect 2835 14725 2840 14755
rect 2800 14720 2840 14725
rect 2880 14915 2920 14920
rect 2880 14885 2885 14915
rect 2915 14885 2920 14915
rect 2880 14755 2920 14885
rect 2880 14725 2885 14755
rect 2915 14725 2920 14755
rect 2880 14720 2920 14725
rect 2960 14915 3000 14920
rect 2960 14885 2965 14915
rect 2995 14885 3000 14915
rect 2960 14755 3000 14885
rect 2960 14725 2965 14755
rect 2995 14725 3000 14755
rect 2960 14720 3000 14725
rect 3040 14915 3080 14920
rect 3040 14885 3045 14915
rect 3075 14885 3080 14915
rect 3040 14755 3080 14885
rect 3040 14725 3045 14755
rect 3075 14725 3080 14755
rect 3040 14720 3080 14725
rect 3120 14915 3160 14920
rect 3120 14885 3125 14915
rect 3155 14885 3160 14915
rect 3120 14755 3160 14885
rect 3120 14725 3125 14755
rect 3155 14725 3160 14755
rect 3120 14720 3160 14725
rect 3200 14915 3240 14920
rect 3200 14885 3205 14915
rect 3235 14885 3240 14915
rect 3200 14755 3240 14885
rect 3200 14725 3205 14755
rect 3235 14725 3240 14755
rect 3200 14720 3240 14725
rect 3280 14915 3320 14920
rect 3280 14885 3285 14915
rect 3315 14885 3320 14915
rect 3280 14755 3320 14885
rect 3280 14725 3285 14755
rect 3315 14725 3320 14755
rect 3280 14720 3320 14725
rect 3360 14915 3400 14920
rect 3360 14885 3365 14915
rect 3395 14885 3400 14915
rect 3360 14755 3400 14885
rect 3360 14725 3365 14755
rect 3395 14725 3400 14755
rect 3360 14720 3400 14725
rect 3440 14915 3480 14920
rect 3440 14885 3445 14915
rect 3475 14885 3480 14915
rect 3440 14755 3480 14885
rect 3440 14725 3445 14755
rect 3475 14725 3480 14755
rect 3440 14720 3480 14725
rect 3520 14915 3560 14920
rect 3520 14885 3525 14915
rect 3555 14885 3560 14915
rect 3520 14755 3560 14885
rect 3520 14725 3525 14755
rect 3555 14725 3560 14755
rect 3520 14720 3560 14725
rect 3600 14915 3640 14920
rect 3600 14885 3605 14915
rect 3635 14885 3640 14915
rect 3600 14755 3640 14885
rect 3600 14725 3605 14755
rect 3635 14725 3640 14755
rect 3600 14720 3640 14725
rect 3680 14915 3720 14920
rect 3680 14885 3685 14915
rect 3715 14885 3720 14915
rect 3680 14755 3720 14885
rect 3680 14725 3685 14755
rect 3715 14725 3720 14755
rect 3680 14720 3720 14725
rect 3760 14915 3800 14920
rect 3760 14885 3765 14915
rect 3795 14885 3800 14915
rect 3760 14755 3800 14885
rect 3760 14725 3765 14755
rect 3795 14725 3800 14755
rect 3760 14720 3800 14725
rect 3840 14915 3880 14920
rect 3840 14885 3845 14915
rect 3875 14885 3880 14915
rect 3840 14755 3880 14885
rect 3840 14725 3845 14755
rect 3875 14725 3880 14755
rect 3840 14720 3880 14725
rect 3920 14915 3960 14920
rect 3920 14885 3925 14915
rect 3955 14885 3960 14915
rect 3920 14755 3960 14885
rect 3920 14725 3925 14755
rect 3955 14725 3960 14755
rect 3920 14720 3960 14725
rect 4000 14915 4040 14920
rect 4000 14885 4005 14915
rect 4035 14885 4040 14915
rect 4000 14755 4040 14885
rect 4000 14725 4005 14755
rect 4035 14725 4040 14755
rect 4000 14720 4040 14725
rect 4080 14915 4120 14920
rect 4080 14885 4085 14915
rect 4115 14885 4120 14915
rect 4080 14755 4120 14885
rect 4080 14725 4085 14755
rect 4115 14725 4120 14755
rect 4080 14720 4120 14725
rect 4160 14915 4200 14920
rect 4160 14885 4165 14915
rect 4195 14885 4200 14915
rect 4160 14755 4200 14885
rect 4160 14725 4165 14755
rect 4195 14725 4200 14755
rect 4160 14720 4200 14725
rect 4240 14680 4280 16485
rect 4320 16595 4360 16680
rect 4320 16565 4325 16595
rect 4355 16565 4360 16595
rect 4320 14680 4360 16565
rect 4400 16675 4440 16680
rect 4400 16645 4405 16675
rect 4435 16645 4440 16675
rect 4400 16515 4440 16645
rect 4400 16485 4405 16515
rect 4435 16485 4440 16515
rect 4400 14680 4440 16485
rect 4480 16435 4520 16680
rect 4480 16405 4485 16435
rect 4515 16405 4520 16435
rect 4480 16275 4520 16405
rect 4480 16245 4485 16275
rect 4515 16245 4520 16275
rect 4480 14680 4520 16245
rect 4560 16355 4600 16680
rect 4560 16325 4565 16355
rect 4595 16325 4600 16355
rect 4560 14680 4600 16325
rect 4640 16435 4680 16680
rect 4640 16405 4645 16435
rect 4675 16405 4680 16435
rect 4640 16275 4680 16405
rect 4640 16245 4645 16275
rect 4675 16245 4680 16275
rect 4640 14680 4680 16245
rect 4720 16195 4760 16680
rect 4720 16165 4725 16195
rect 4755 16165 4760 16195
rect 4720 16035 4760 16165
rect 4720 16005 4725 16035
rect 4755 16005 4760 16035
rect 4720 15875 4760 16005
rect 4720 15845 4725 15875
rect 4755 15845 4760 15875
rect 4720 15715 4760 15845
rect 4720 15685 4725 15715
rect 4755 15685 4760 15715
rect 4720 15555 4760 15685
rect 4720 15525 4725 15555
rect 4755 15525 4760 15555
rect 4720 15395 4760 15525
rect 4720 15365 4725 15395
rect 4755 15365 4760 15395
rect 4720 15235 4760 15365
rect 4720 15205 4725 15235
rect 4755 15205 4760 15235
rect 4720 14680 4760 15205
rect 4800 16115 4840 16680
rect 4800 16085 4805 16115
rect 4835 16085 4840 16115
rect 4800 14680 4840 16085
rect 4880 16195 4920 16680
rect 4880 16165 4885 16195
rect 4915 16165 4920 16195
rect 4880 16035 4920 16165
rect 4880 16005 4885 16035
rect 4915 16005 4920 16035
rect 4880 15875 4920 16005
rect 4880 15845 4885 15875
rect 4915 15845 4920 15875
rect 4880 15715 4920 15845
rect 4880 15685 4885 15715
rect 4915 15685 4920 15715
rect 4880 15555 4920 15685
rect 4880 15525 4885 15555
rect 4915 15525 4920 15555
rect 4880 15395 4920 15525
rect 4880 15365 4885 15395
rect 4915 15365 4920 15395
rect 4880 15235 4920 15365
rect 4880 15205 4885 15235
rect 4915 15205 4920 15235
rect 4880 14680 4920 15205
rect 4960 15955 5000 16680
rect 4960 15925 4965 15955
rect 4995 15925 5000 15955
rect 4960 14680 5000 15925
rect 5040 16195 5080 16680
rect 5040 16165 5045 16195
rect 5075 16165 5080 16195
rect 5040 16035 5080 16165
rect 5040 16005 5045 16035
rect 5075 16005 5080 16035
rect 5040 15875 5080 16005
rect 5040 15845 5045 15875
rect 5075 15845 5080 15875
rect 5040 15715 5080 15845
rect 5040 15685 5045 15715
rect 5075 15685 5080 15715
rect 5040 15555 5080 15685
rect 5040 15525 5045 15555
rect 5075 15525 5080 15555
rect 5040 15395 5080 15525
rect 5040 15365 5045 15395
rect 5075 15365 5080 15395
rect 5040 15235 5080 15365
rect 5040 15205 5045 15235
rect 5075 15205 5080 15235
rect 5040 14680 5080 15205
rect 5120 15795 5160 16680
rect 5120 15765 5125 15795
rect 5155 15765 5160 15795
rect 5120 14680 5160 15765
rect 5200 16195 5240 16680
rect 5200 16165 5205 16195
rect 5235 16165 5240 16195
rect 5200 16035 5240 16165
rect 5200 16005 5205 16035
rect 5235 16005 5240 16035
rect 5200 15875 5240 16005
rect 5200 15845 5205 15875
rect 5235 15845 5240 15875
rect 5200 15715 5240 15845
rect 5200 15685 5205 15715
rect 5235 15685 5240 15715
rect 5200 15555 5240 15685
rect 5200 15525 5205 15555
rect 5235 15525 5240 15555
rect 5200 15395 5240 15525
rect 5200 15365 5205 15395
rect 5235 15365 5240 15395
rect 5200 15235 5240 15365
rect 5200 15205 5205 15235
rect 5235 15205 5240 15235
rect 5200 14680 5240 15205
rect 5280 15635 5320 16680
rect 5280 15605 5285 15635
rect 5315 15605 5320 15635
rect 5280 14680 5320 15605
rect 5360 16195 5400 16680
rect 5360 16165 5365 16195
rect 5395 16165 5400 16195
rect 5360 16035 5400 16165
rect 5360 16005 5365 16035
rect 5395 16005 5400 16035
rect 5360 15875 5400 16005
rect 5360 15845 5365 15875
rect 5395 15845 5400 15875
rect 5360 15715 5400 15845
rect 5360 15685 5365 15715
rect 5395 15685 5400 15715
rect 5360 15555 5400 15685
rect 5360 15525 5365 15555
rect 5395 15525 5400 15555
rect 5360 15395 5400 15525
rect 5360 15365 5365 15395
rect 5395 15365 5400 15395
rect 5360 15235 5400 15365
rect 5360 15205 5365 15235
rect 5395 15205 5400 15235
rect 5360 14680 5400 15205
rect 5440 15475 5480 16680
rect 5440 15445 5445 15475
rect 5475 15445 5480 15475
rect 5440 14680 5480 15445
rect 5520 16195 5560 16680
rect 5520 16165 5525 16195
rect 5555 16165 5560 16195
rect 5520 16035 5560 16165
rect 5520 16005 5525 16035
rect 5555 16005 5560 16035
rect 5520 15875 5560 16005
rect 5520 15845 5525 15875
rect 5555 15845 5560 15875
rect 5520 15715 5560 15845
rect 5520 15685 5525 15715
rect 5555 15685 5560 15715
rect 5520 15555 5560 15685
rect 5520 15525 5525 15555
rect 5555 15525 5560 15555
rect 5520 15395 5560 15525
rect 5520 15365 5525 15395
rect 5555 15365 5560 15395
rect 5520 15235 5560 15365
rect 5520 15205 5525 15235
rect 5555 15205 5560 15235
rect 5520 14680 5560 15205
rect 5600 15315 5640 16680
rect 5600 15285 5605 15315
rect 5635 15285 5640 15315
rect 5600 14680 5640 15285
rect 5680 16195 5720 16680
rect 5680 16165 5685 16195
rect 5715 16165 5720 16195
rect 5680 16035 5720 16165
rect 5680 16005 5685 16035
rect 5715 16005 5720 16035
rect 5680 15875 5720 16005
rect 5680 15845 5685 15875
rect 5715 15845 5720 15875
rect 5680 15715 5720 15845
rect 5680 15685 5685 15715
rect 5715 15685 5720 15715
rect 5680 15555 5720 15685
rect 5680 15525 5685 15555
rect 5715 15525 5720 15555
rect 5680 15395 5720 15525
rect 5680 15365 5685 15395
rect 5715 15365 5720 15395
rect 5680 15235 5720 15365
rect 5680 15205 5685 15235
rect 5715 15205 5720 15235
rect 5680 14680 5720 15205
rect 5760 15155 5800 16680
rect 5760 15125 5765 15155
rect 5795 15125 5800 15155
rect 5760 14995 5800 15125
rect 5760 14965 5765 14995
rect 5795 14965 5800 14995
rect 5760 14680 5800 14965
rect 5840 15075 5880 16680
rect 5840 15045 5845 15075
rect 5875 15045 5880 15075
rect 5840 14680 5880 15045
rect 5920 15155 5960 16680
rect 5920 15125 5925 15155
rect 5955 15125 5960 15155
rect 5920 14995 5960 15125
rect 5920 14965 5925 14995
rect 5955 14965 5960 14995
rect 5920 14680 5960 14965
rect 6000 14915 6040 16680
rect 6000 14885 6005 14915
rect 6035 14885 6040 14915
rect 6000 14755 6040 14885
rect 6000 14725 6005 14755
rect 6035 14725 6040 14755
rect 6000 14680 6040 14725
rect 6080 14835 6120 16680
rect 6080 14805 6085 14835
rect 6115 14805 6120 14835
rect 6080 14680 6120 14805
rect 6160 14915 6200 16680
rect 6240 16675 6280 16680
rect 6240 16645 6245 16675
rect 6275 16645 6280 16675
rect 6240 16515 6280 16645
rect 6240 16485 6245 16515
rect 6275 16485 6280 16515
rect 6240 16480 6280 16485
rect 6320 16675 6360 16680
rect 6320 16645 6325 16675
rect 6355 16645 6360 16675
rect 6320 16515 6360 16645
rect 6320 16485 6325 16515
rect 6355 16485 6360 16515
rect 6320 16480 6360 16485
rect 6400 16675 6440 16680
rect 6400 16645 6405 16675
rect 6435 16645 6440 16675
rect 6400 16515 6440 16645
rect 6400 16485 6405 16515
rect 6435 16485 6440 16515
rect 6400 16480 6440 16485
rect 6480 16675 6520 16680
rect 6480 16645 6485 16675
rect 6515 16645 6520 16675
rect 6480 16515 6520 16645
rect 6480 16485 6485 16515
rect 6515 16485 6520 16515
rect 6480 16480 6520 16485
rect 6560 16675 6600 16680
rect 6560 16645 6565 16675
rect 6595 16645 6600 16675
rect 6560 16515 6600 16645
rect 6560 16485 6565 16515
rect 6595 16485 6600 16515
rect 6560 16480 6600 16485
rect 6640 16675 6680 16680
rect 6640 16645 6645 16675
rect 6675 16645 6680 16675
rect 6640 16515 6680 16645
rect 6640 16485 6645 16515
rect 6675 16485 6680 16515
rect 6640 16480 6680 16485
rect 6720 16675 6760 16680
rect 6720 16645 6725 16675
rect 6755 16645 6760 16675
rect 6720 16515 6760 16645
rect 6720 16485 6725 16515
rect 6755 16485 6760 16515
rect 6720 16480 6760 16485
rect 6800 16675 6840 16680
rect 6800 16645 6805 16675
rect 6835 16645 6840 16675
rect 6800 16515 6840 16645
rect 6800 16485 6805 16515
rect 6835 16485 6840 16515
rect 6800 16480 6840 16485
rect 6880 16675 6920 16680
rect 6880 16645 6885 16675
rect 6915 16645 6920 16675
rect 6880 16515 6920 16645
rect 6880 16485 6885 16515
rect 6915 16485 6920 16515
rect 6880 16480 6920 16485
rect 6960 16675 7000 16680
rect 6960 16645 6965 16675
rect 6995 16645 7000 16675
rect 6960 16515 7000 16645
rect 6960 16485 6965 16515
rect 6995 16485 7000 16515
rect 6960 16480 7000 16485
rect 7040 16675 7080 16680
rect 7040 16645 7045 16675
rect 7075 16645 7080 16675
rect 7040 16515 7080 16645
rect 7040 16485 7045 16515
rect 7075 16485 7080 16515
rect 7040 16480 7080 16485
rect 7120 16675 7160 16680
rect 7120 16645 7125 16675
rect 7155 16645 7160 16675
rect 7120 16515 7160 16645
rect 7120 16485 7125 16515
rect 7155 16485 7160 16515
rect 7120 16480 7160 16485
rect 7200 16675 7240 16680
rect 7200 16645 7205 16675
rect 7235 16645 7240 16675
rect 7200 16515 7240 16645
rect 7200 16485 7205 16515
rect 7235 16485 7240 16515
rect 7200 16480 7240 16485
rect 7280 16675 7320 16680
rect 7280 16645 7285 16675
rect 7315 16645 7320 16675
rect 7280 16515 7320 16645
rect 7280 16485 7285 16515
rect 7315 16485 7320 16515
rect 7280 16480 7320 16485
rect 7360 16675 7400 16680
rect 7360 16645 7365 16675
rect 7395 16645 7400 16675
rect 7360 16515 7400 16645
rect 7360 16485 7365 16515
rect 7395 16485 7400 16515
rect 7360 16480 7400 16485
rect 7440 16675 7480 16680
rect 7440 16645 7445 16675
rect 7475 16645 7480 16675
rect 7440 16515 7480 16645
rect 7440 16485 7445 16515
rect 7475 16485 7480 16515
rect 7440 16480 7480 16485
rect 7520 16675 7560 16680
rect 7520 16645 7525 16675
rect 7555 16645 7560 16675
rect 7520 16515 7560 16645
rect 7520 16485 7525 16515
rect 7555 16485 7560 16515
rect 7520 16480 7560 16485
rect 7600 16675 7640 16680
rect 7600 16645 7605 16675
rect 7635 16645 7640 16675
rect 7600 16515 7640 16645
rect 7600 16485 7605 16515
rect 7635 16485 7640 16515
rect 7600 16480 7640 16485
rect 7680 16675 7720 16680
rect 7680 16645 7685 16675
rect 7715 16645 7720 16675
rect 7680 16515 7720 16645
rect 7680 16485 7685 16515
rect 7715 16485 7720 16515
rect 7680 16480 7720 16485
rect 7760 16675 7800 16680
rect 7760 16645 7765 16675
rect 7795 16645 7800 16675
rect 7760 16515 7800 16645
rect 7760 16485 7765 16515
rect 7795 16485 7800 16515
rect 7760 16480 7800 16485
rect 7840 16675 7880 16680
rect 7840 16645 7845 16675
rect 7875 16645 7880 16675
rect 7840 16515 7880 16645
rect 7840 16485 7845 16515
rect 7875 16485 7880 16515
rect 7840 16480 7880 16485
rect 7920 16675 7960 16680
rect 7920 16645 7925 16675
rect 7955 16645 7960 16675
rect 7920 16515 7960 16645
rect 7920 16485 7925 16515
rect 7955 16485 7960 16515
rect 7920 16480 7960 16485
rect 8000 16675 8040 16680
rect 8000 16645 8005 16675
rect 8035 16645 8040 16675
rect 8000 16515 8040 16645
rect 8000 16485 8005 16515
rect 8035 16485 8040 16515
rect 8000 16480 8040 16485
rect 8080 16675 8120 16680
rect 8080 16645 8085 16675
rect 8115 16645 8120 16675
rect 8080 16515 8120 16645
rect 8080 16485 8085 16515
rect 8115 16485 8120 16515
rect 8080 16480 8120 16485
rect 8160 16675 8200 16680
rect 8160 16645 8165 16675
rect 8195 16645 8200 16675
rect 8160 16515 8200 16645
rect 8160 16485 8165 16515
rect 8195 16485 8200 16515
rect 8160 16480 8200 16485
rect 8240 16675 8280 16680
rect 8240 16645 8245 16675
rect 8275 16645 8280 16675
rect 8240 16515 8280 16645
rect 8240 16485 8245 16515
rect 8275 16485 8280 16515
rect 8240 16480 8280 16485
rect 8320 16675 8360 16680
rect 8320 16645 8325 16675
rect 8355 16645 8360 16675
rect 8320 16515 8360 16645
rect 8320 16485 8325 16515
rect 8355 16485 8360 16515
rect 8320 16480 8360 16485
rect 8400 16675 8440 16680
rect 8400 16645 8405 16675
rect 8435 16645 8440 16675
rect 8400 16515 8440 16645
rect 8400 16485 8405 16515
rect 8435 16485 8440 16515
rect 8400 16480 8440 16485
rect 8480 16675 8520 16680
rect 8480 16645 8485 16675
rect 8515 16645 8520 16675
rect 8480 16515 8520 16645
rect 8480 16485 8485 16515
rect 8515 16485 8520 16515
rect 8480 16480 8520 16485
rect 8560 16675 8600 16680
rect 8560 16645 8565 16675
rect 8595 16645 8600 16675
rect 8560 16515 8600 16645
rect 8560 16485 8565 16515
rect 8595 16485 8600 16515
rect 8560 16480 8600 16485
rect 8640 16675 8680 16680
rect 8640 16645 8645 16675
rect 8675 16645 8680 16675
rect 8640 16515 8680 16645
rect 8640 16485 8645 16515
rect 8675 16485 8680 16515
rect 8640 16480 8680 16485
rect 8720 16675 8760 16680
rect 8720 16645 8725 16675
rect 8755 16645 8760 16675
rect 8720 16515 8760 16645
rect 8720 16485 8725 16515
rect 8755 16485 8760 16515
rect 8720 16480 8760 16485
rect 8800 16675 8840 16680
rect 8800 16645 8805 16675
rect 8835 16645 8840 16675
rect 8800 16515 8840 16645
rect 8800 16485 8805 16515
rect 8835 16485 8840 16515
rect 8800 16480 8840 16485
rect 8880 16675 8920 16680
rect 8880 16645 8885 16675
rect 8915 16645 8920 16675
rect 8880 16515 8920 16645
rect 8880 16485 8885 16515
rect 8915 16485 8920 16515
rect 8880 16480 8920 16485
rect 8960 16675 9000 16680
rect 8960 16645 8965 16675
rect 8995 16645 9000 16675
rect 8960 16515 9000 16645
rect 8960 16485 8965 16515
rect 8995 16485 9000 16515
rect 8960 16480 9000 16485
rect 9040 16675 9080 16680
rect 9040 16645 9045 16675
rect 9075 16645 9080 16675
rect 9040 16515 9080 16645
rect 9040 16485 9045 16515
rect 9075 16485 9080 16515
rect 9040 16480 9080 16485
rect 9120 16675 9160 16680
rect 9120 16645 9125 16675
rect 9155 16645 9160 16675
rect 9120 16515 9160 16645
rect 9120 16485 9125 16515
rect 9155 16485 9160 16515
rect 9120 16480 9160 16485
rect 9200 16675 9240 16680
rect 9200 16645 9205 16675
rect 9235 16645 9240 16675
rect 9200 16515 9240 16645
rect 9200 16485 9205 16515
rect 9235 16485 9240 16515
rect 9200 16480 9240 16485
rect 9280 16675 9320 16680
rect 9280 16645 9285 16675
rect 9315 16645 9320 16675
rect 9280 16515 9320 16645
rect 9280 16485 9285 16515
rect 9315 16485 9320 16515
rect 9280 16480 9320 16485
rect 9360 16675 9400 16680
rect 9360 16645 9365 16675
rect 9395 16645 9400 16675
rect 9360 16515 9400 16645
rect 9360 16485 9365 16515
rect 9395 16485 9400 16515
rect 9360 16480 9400 16485
rect 9440 16675 9480 16680
rect 9440 16645 9445 16675
rect 9475 16645 9480 16675
rect 9440 16515 9480 16645
rect 9440 16485 9445 16515
rect 9475 16485 9480 16515
rect 9440 16480 9480 16485
rect 9520 16675 9560 16725
rect 9520 16645 9525 16675
rect 9555 16645 9560 16675
rect 9520 16515 9560 16645
rect 9520 16485 9525 16515
rect 9555 16485 9560 16515
rect 6240 16435 6280 16440
rect 6240 16405 6245 16435
rect 6275 16405 6280 16435
rect 6240 16275 6280 16405
rect 6240 16245 6245 16275
rect 6275 16245 6280 16275
rect 6240 16240 6280 16245
rect 6320 16435 6360 16440
rect 6320 16405 6325 16435
rect 6355 16405 6360 16435
rect 6320 16275 6360 16405
rect 6320 16245 6325 16275
rect 6355 16245 6360 16275
rect 6320 16240 6360 16245
rect 6400 16435 6440 16440
rect 6400 16405 6405 16435
rect 6435 16405 6440 16435
rect 6400 16275 6440 16405
rect 6400 16245 6405 16275
rect 6435 16245 6440 16275
rect 6400 16240 6440 16245
rect 6480 16435 6520 16440
rect 6480 16405 6485 16435
rect 6515 16405 6520 16435
rect 6480 16275 6520 16405
rect 6480 16245 6485 16275
rect 6515 16245 6520 16275
rect 6480 16240 6520 16245
rect 6560 16435 6600 16440
rect 6560 16405 6565 16435
rect 6595 16405 6600 16435
rect 6560 16275 6600 16405
rect 6560 16245 6565 16275
rect 6595 16245 6600 16275
rect 6560 16240 6600 16245
rect 6640 16435 6680 16440
rect 6640 16405 6645 16435
rect 6675 16405 6680 16435
rect 6640 16275 6680 16405
rect 6640 16245 6645 16275
rect 6675 16245 6680 16275
rect 6640 16240 6680 16245
rect 6720 16435 6760 16440
rect 6720 16405 6725 16435
rect 6755 16405 6760 16435
rect 6720 16275 6760 16405
rect 6720 16245 6725 16275
rect 6755 16245 6760 16275
rect 6720 16240 6760 16245
rect 6800 16435 6840 16440
rect 6800 16405 6805 16435
rect 6835 16405 6840 16435
rect 6800 16275 6840 16405
rect 6800 16245 6805 16275
rect 6835 16245 6840 16275
rect 6800 16240 6840 16245
rect 6880 16435 6920 16440
rect 6880 16405 6885 16435
rect 6915 16405 6920 16435
rect 6880 16275 6920 16405
rect 6880 16245 6885 16275
rect 6915 16245 6920 16275
rect 6880 16240 6920 16245
rect 6960 16435 7000 16440
rect 6960 16405 6965 16435
rect 6995 16405 7000 16435
rect 6960 16275 7000 16405
rect 6960 16245 6965 16275
rect 6995 16245 7000 16275
rect 6960 16240 7000 16245
rect 7040 16435 7080 16440
rect 7040 16405 7045 16435
rect 7075 16405 7080 16435
rect 7040 16275 7080 16405
rect 7040 16245 7045 16275
rect 7075 16245 7080 16275
rect 7040 16240 7080 16245
rect 7120 16435 7160 16440
rect 7120 16405 7125 16435
rect 7155 16405 7160 16435
rect 7120 16275 7160 16405
rect 7120 16245 7125 16275
rect 7155 16245 7160 16275
rect 7120 16240 7160 16245
rect 7200 16435 7240 16440
rect 7200 16405 7205 16435
rect 7235 16405 7240 16435
rect 7200 16275 7240 16405
rect 7200 16245 7205 16275
rect 7235 16245 7240 16275
rect 7200 16240 7240 16245
rect 7280 16435 7320 16440
rect 7280 16405 7285 16435
rect 7315 16405 7320 16435
rect 7280 16275 7320 16405
rect 7280 16245 7285 16275
rect 7315 16245 7320 16275
rect 7280 16240 7320 16245
rect 7360 16435 7400 16440
rect 7360 16405 7365 16435
rect 7395 16405 7400 16435
rect 7360 16275 7400 16405
rect 7360 16245 7365 16275
rect 7395 16245 7400 16275
rect 7360 16240 7400 16245
rect 7440 16435 7480 16440
rect 7440 16405 7445 16435
rect 7475 16405 7480 16435
rect 7440 16275 7480 16405
rect 7440 16245 7445 16275
rect 7475 16245 7480 16275
rect 7440 16240 7480 16245
rect 7520 16435 7560 16440
rect 7520 16405 7525 16435
rect 7555 16405 7560 16435
rect 7520 16275 7560 16405
rect 7520 16245 7525 16275
rect 7555 16245 7560 16275
rect 7520 16240 7560 16245
rect 7600 16435 7640 16440
rect 7600 16405 7605 16435
rect 7635 16405 7640 16435
rect 7600 16275 7640 16405
rect 7600 16245 7605 16275
rect 7635 16245 7640 16275
rect 7600 16240 7640 16245
rect 7680 16435 7720 16440
rect 7680 16405 7685 16435
rect 7715 16405 7720 16435
rect 7680 16275 7720 16405
rect 7680 16245 7685 16275
rect 7715 16245 7720 16275
rect 7680 16240 7720 16245
rect 7760 16435 7800 16440
rect 7760 16405 7765 16435
rect 7795 16405 7800 16435
rect 7760 16275 7800 16405
rect 7760 16245 7765 16275
rect 7795 16245 7800 16275
rect 7760 16240 7800 16245
rect 7840 16435 7880 16440
rect 7840 16405 7845 16435
rect 7875 16405 7880 16435
rect 7840 16275 7880 16405
rect 7840 16245 7845 16275
rect 7875 16245 7880 16275
rect 7840 16240 7880 16245
rect 7920 16435 7960 16440
rect 7920 16405 7925 16435
rect 7955 16405 7960 16435
rect 7920 16275 7960 16405
rect 7920 16245 7925 16275
rect 7955 16245 7960 16275
rect 7920 16240 7960 16245
rect 8000 16435 8040 16440
rect 8000 16405 8005 16435
rect 8035 16405 8040 16435
rect 8000 16275 8040 16405
rect 8000 16245 8005 16275
rect 8035 16245 8040 16275
rect 8000 16240 8040 16245
rect 8080 16435 8120 16440
rect 8080 16405 8085 16435
rect 8115 16405 8120 16435
rect 8080 16275 8120 16405
rect 8080 16245 8085 16275
rect 8115 16245 8120 16275
rect 8080 16240 8120 16245
rect 8160 16435 8200 16440
rect 8160 16405 8165 16435
rect 8195 16405 8200 16435
rect 8160 16275 8200 16405
rect 8160 16245 8165 16275
rect 8195 16245 8200 16275
rect 8160 16240 8200 16245
rect 8240 16435 8280 16440
rect 8240 16405 8245 16435
rect 8275 16405 8280 16435
rect 8240 16275 8280 16405
rect 8240 16245 8245 16275
rect 8275 16245 8280 16275
rect 8240 16240 8280 16245
rect 8320 16435 8360 16440
rect 8320 16405 8325 16435
rect 8355 16405 8360 16435
rect 8320 16275 8360 16405
rect 8320 16245 8325 16275
rect 8355 16245 8360 16275
rect 8320 16240 8360 16245
rect 8400 16435 8440 16440
rect 8400 16405 8405 16435
rect 8435 16405 8440 16435
rect 8400 16275 8440 16405
rect 8400 16245 8405 16275
rect 8435 16245 8440 16275
rect 8400 16240 8440 16245
rect 8480 16435 8520 16440
rect 8480 16405 8485 16435
rect 8515 16405 8520 16435
rect 8480 16275 8520 16405
rect 8480 16245 8485 16275
rect 8515 16245 8520 16275
rect 8480 16240 8520 16245
rect 8560 16435 8600 16440
rect 8560 16405 8565 16435
rect 8595 16405 8600 16435
rect 8560 16275 8600 16405
rect 8560 16245 8565 16275
rect 8595 16245 8600 16275
rect 8560 16240 8600 16245
rect 8640 16435 8680 16440
rect 8640 16405 8645 16435
rect 8675 16405 8680 16435
rect 8640 16275 8680 16405
rect 8640 16245 8645 16275
rect 8675 16245 8680 16275
rect 8640 16240 8680 16245
rect 8720 16435 8760 16440
rect 8720 16405 8725 16435
rect 8755 16405 8760 16435
rect 8720 16275 8760 16405
rect 8720 16245 8725 16275
rect 8755 16245 8760 16275
rect 8720 16240 8760 16245
rect 8800 16435 8840 16440
rect 8800 16405 8805 16435
rect 8835 16405 8840 16435
rect 8800 16275 8840 16405
rect 8800 16245 8805 16275
rect 8835 16245 8840 16275
rect 8800 16240 8840 16245
rect 8880 16435 8920 16440
rect 8880 16405 8885 16435
rect 8915 16405 8920 16435
rect 8880 16275 8920 16405
rect 8880 16245 8885 16275
rect 8915 16245 8920 16275
rect 8880 16240 8920 16245
rect 8960 16435 9000 16440
rect 8960 16405 8965 16435
rect 8995 16405 9000 16435
rect 8960 16275 9000 16405
rect 8960 16245 8965 16275
rect 8995 16245 9000 16275
rect 8960 16240 9000 16245
rect 9040 16435 9080 16440
rect 9040 16405 9045 16435
rect 9075 16405 9080 16435
rect 9040 16275 9080 16405
rect 9040 16245 9045 16275
rect 9075 16245 9080 16275
rect 9040 16240 9080 16245
rect 9120 16435 9160 16440
rect 9120 16405 9125 16435
rect 9155 16405 9160 16435
rect 9120 16275 9160 16405
rect 9120 16245 9125 16275
rect 9155 16245 9160 16275
rect 9120 16240 9160 16245
rect 9200 16435 9240 16440
rect 9200 16405 9205 16435
rect 9235 16405 9240 16435
rect 9200 16275 9240 16405
rect 9200 16245 9205 16275
rect 9235 16245 9240 16275
rect 9200 16240 9240 16245
rect 9280 16435 9320 16440
rect 9280 16405 9285 16435
rect 9315 16405 9320 16435
rect 9280 16275 9320 16405
rect 9280 16245 9285 16275
rect 9315 16245 9320 16275
rect 9280 16240 9320 16245
rect 9360 16435 9400 16440
rect 9360 16405 9365 16435
rect 9395 16405 9400 16435
rect 9360 16275 9400 16405
rect 9360 16245 9365 16275
rect 9395 16245 9400 16275
rect 9360 16240 9400 16245
rect 9440 16435 9480 16440
rect 9440 16405 9445 16435
rect 9475 16405 9480 16435
rect 9440 16275 9480 16405
rect 9440 16245 9445 16275
rect 9475 16245 9480 16275
rect 9440 16240 9480 16245
rect 6240 16195 6280 16200
rect 6240 16165 6245 16195
rect 6275 16165 6280 16195
rect 6240 16035 6280 16165
rect 6240 16005 6245 16035
rect 6275 16005 6280 16035
rect 6240 15875 6280 16005
rect 6240 15845 6245 15875
rect 6275 15845 6280 15875
rect 6240 15715 6280 15845
rect 6240 15685 6245 15715
rect 6275 15685 6280 15715
rect 6240 15555 6280 15685
rect 6240 15525 6245 15555
rect 6275 15525 6280 15555
rect 6240 15395 6280 15525
rect 6240 15365 6245 15395
rect 6275 15365 6280 15395
rect 6240 15235 6280 15365
rect 6240 15205 6245 15235
rect 6275 15205 6280 15235
rect 6240 15200 6280 15205
rect 6320 16195 6360 16200
rect 6320 16165 6325 16195
rect 6355 16165 6360 16195
rect 6320 16035 6360 16165
rect 6320 16005 6325 16035
rect 6355 16005 6360 16035
rect 6320 15875 6360 16005
rect 6320 15845 6325 15875
rect 6355 15845 6360 15875
rect 6320 15715 6360 15845
rect 6320 15685 6325 15715
rect 6355 15685 6360 15715
rect 6320 15555 6360 15685
rect 6320 15525 6325 15555
rect 6355 15525 6360 15555
rect 6320 15395 6360 15525
rect 6320 15365 6325 15395
rect 6355 15365 6360 15395
rect 6320 15235 6360 15365
rect 6320 15205 6325 15235
rect 6355 15205 6360 15235
rect 6320 15200 6360 15205
rect 6400 16195 6440 16200
rect 6400 16165 6405 16195
rect 6435 16165 6440 16195
rect 6400 16035 6440 16165
rect 6400 16005 6405 16035
rect 6435 16005 6440 16035
rect 6400 15875 6440 16005
rect 6400 15845 6405 15875
rect 6435 15845 6440 15875
rect 6400 15715 6440 15845
rect 6400 15685 6405 15715
rect 6435 15685 6440 15715
rect 6400 15555 6440 15685
rect 6400 15525 6405 15555
rect 6435 15525 6440 15555
rect 6400 15395 6440 15525
rect 6400 15365 6405 15395
rect 6435 15365 6440 15395
rect 6400 15235 6440 15365
rect 6400 15205 6405 15235
rect 6435 15205 6440 15235
rect 6400 15200 6440 15205
rect 6480 16195 6520 16200
rect 6480 16165 6485 16195
rect 6515 16165 6520 16195
rect 6480 16035 6520 16165
rect 6480 16005 6485 16035
rect 6515 16005 6520 16035
rect 6480 15875 6520 16005
rect 6480 15845 6485 15875
rect 6515 15845 6520 15875
rect 6480 15715 6520 15845
rect 6480 15685 6485 15715
rect 6515 15685 6520 15715
rect 6480 15555 6520 15685
rect 6480 15525 6485 15555
rect 6515 15525 6520 15555
rect 6480 15395 6520 15525
rect 6480 15365 6485 15395
rect 6515 15365 6520 15395
rect 6480 15235 6520 15365
rect 6480 15205 6485 15235
rect 6515 15205 6520 15235
rect 6480 15200 6520 15205
rect 6560 16195 6600 16200
rect 6560 16165 6565 16195
rect 6595 16165 6600 16195
rect 6560 16035 6600 16165
rect 6560 16005 6565 16035
rect 6595 16005 6600 16035
rect 6560 15875 6600 16005
rect 6560 15845 6565 15875
rect 6595 15845 6600 15875
rect 6560 15715 6600 15845
rect 6560 15685 6565 15715
rect 6595 15685 6600 15715
rect 6560 15555 6600 15685
rect 6560 15525 6565 15555
rect 6595 15525 6600 15555
rect 6560 15395 6600 15525
rect 6560 15365 6565 15395
rect 6595 15365 6600 15395
rect 6560 15235 6600 15365
rect 6560 15205 6565 15235
rect 6595 15205 6600 15235
rect 6560 15200 6600 15205
rect 6640 16195 6680 16200
rect 6640 16165 6645 16195
rect 6675 16165 6680 16195
rect 6640 16035 6680 16165
rect 6640 16005 6645 16035
rect 6675 16005 6680 16035
rect 6640 15875 6680 16005
rect 6640 15845 6645 15875
rect 6675 15845 6680 15875
rect 6640 15715 6680 15845
rect 6640 15685 6645 15715
rect 6675 15685 6680 15715
rect 6640 15555 6680 15685
rect 6640 15525 6645 15555
rect 6675 15525 6680 15555
rect 6640 15395 6680 15525
rect 6640 15365 6645 15395
rect 6675 15365 6680 15395
rect 6640 15235 6680 15365
rect 6640 15205 6645 15235
rect 6675 15205 6680 15235
rect 6640 15200 6680 15205
rect 6720 16195 6760 16200
rect 6720 16165 6725 16195
rect 6755 16165 6760 16195
rect 6720 16035 6760 16165
rect 6720 16005 6725 16035
rect 6755 16005 6760 16035
rect 6720 15875 6760 16005
rect 6720 15845 6725 15875
rect 6755 15845 6760 15875
rect 6720 15715 6760 15845
rect 6720 15685 6725 15715
rect 6755 15685 6760 15715
rect 6720 15555 6760 15685
rect 6720 15525 6725 15555
rect 6755 15525 6760 15555
rect 6720 15395 6760 15525
rect 6720 15365 6725 15395
rect 6755 15365 6760 15395
rect 6720 15235 6760 15365
rect 6720 15205 6725 15235
rect 6755 15205 6760 15235
rect 6720 15200 6760 15205
rect 6800 16195 6840 16200
rect 6800 16165 6805 16195
rect 6835 16165 6840 16195
rect 6800 16035 6840 16165
rect 6800 16005 6805 16035
rect 6835 16005 6840 16035
rect 6800 15875 6840 16005
rect 6800 15845 6805 15875
rect 6835 15845 6840 15875
rect 6800 15715 6840 15845
rect 6800 15685 6805 15715
rect 6835 15685 6840 15715
rect 6800 15555 6840 15685
rect 6800 15525 6805 15555
rect 6835 15525 6840 15555
rect 6800 15395 6840 15525
rect 6800 15365 6805 15395
rect 6835 15365 6840 15395
rect 6800 15235 6840 15365
rect 6800 15205 6805 15235
rect 6835 15205 6840 15235
rect 6800 15200 6840 15205
rect 6880 16195 6920 16200
rect 6880 16165 6885 16195
rect 6915 16165 6920 16195
rect 6880 16035 6920 16165
rect 6880 16005 6885 16035
rect 6915 16005 6920 16035
rect 6880 15875 6920 16005
rect 6880 15845 6885 15875
rect 6915 15845 6920 15875
rect 6880 15715 6920 15845
rect 6880 15685 6885 15715
rect 6915 15685 6920 15715
rect 6880 15555 6920 15685
rect 6880 15525 6885 15555
rect 6915 15525 6920 15555
rect 6880 15395 6920 15525
rect 6880 15365 6885 15395
rect 6915 15365 6920 15395
rect 6880 15235 6920 15365
rect 6880 15205 6885 15235
rect 6915 15205 6920 15235
rect 6880 15200 6920 15205
rect 6960 16195 7000 16200
rect 6960 16165 6965 16195
rect 6995 16165 7000 16195
rect 6960 16035 7000 16165
rect 6960 16005 6965 16035
rect 6995 16005 7000 16035
rect 6960 15875 7000 16005
rect 6960 15845 6965 15875
rect 6995 15845 7000 15875
rect 6960 15715 7000 15845
rect 6960 15685 6965 15715
rect 6995 15685 7000 15715
rect 6960 15555 7000 15685
rect 6960 15525 6965 15555
rect 6995 15525 7000 15555
rect 6960 15395 7000 15525
rect 6960 15365 6965 15395
rect 6995 15365 7000 15395
rect 6960 15235 7000 15365
rect 6960 15205 6965 15235
rect 6995 15205 7000 15235
rect 6960 15200 7000 15205
rect 7040 16195 7080 16200
rect 7040 16165 7045 16195
rect 7075 16165 7080 16195
rect 7040 16035 7080 16165
rect 7040 16005 7045 16035
rect 7075 16005 7080 16035
rect 7040 15875 7080 16005
rect 7040 15845 7045 15875
rect 7075 15845 7080 15875
rect 7040 15715 7080 15845
rect 7040 15685 7045 15715
rect 7075 15685 7080 15715
rect 7040 15555 7080 15685
rect 7040 15525 7045 15555
rect 7075 15525 7080 15555
rect 7040 15395 7080 15525
rect 7040 15365 7045 15395
rect 7075 15365 7080 15395
rect 7040 15235 7080 15365
rect 7040 15205 7045 15235
rect 7075 15205 7080 15235
rect 7040 15200 7080 15205
rect 7120 16195 7160 16200
rect 7120 16165 7125 16195
rect 7155 16165 7160 16195
rect 7120 16035 7160 16165
rect 7120 16005 7125 16035
rect 7155 16005 7160 16035
rect 7120 15875 7160 16005
rect 7120 15845 7125 15875
rect 7155 15845 7160 15875
rect 7120 15715 7160 15845
rect 7120 15685 7125 15715
rect 7155 15685 7160 15715
rect 7120 15555 7160 15685
rect 7120 15525 7125 15555
rect 7155 15525 7160 15555
rect 7120 15395 7160 15525
rect 7120 15365 7125 15395
rect 7155 15365 7160 15395
rect 7120 15235 7160 15365
rect 7120 15205 7125 15235
rect 7155 15205 7160 15235
rect 7120 15200 7160 15205
rect 7200 16195 7240 16200
rect 7200 16165 7205 16195
rect 7235 16165 7240 16195
rect 7200 16035 7240 16165
rect 7200 16005 7205 16035
rect 7235 16005 7240 16035
rect 7200 15875 7240 16005
rect 7200 15845 7205 15875
rect 7235 15845 7240 15875
rect 7200 15715 7240 15845
rect 7200 15685 7205 15715
rect 7235 15685 7240 15715
rect 7200 15555 7240 15685
rect 7200 15525 7205 15555
rect 7235 15525 7240 15555
rect 7200 15395 7240 15525
rect 7200 15365 7205 15395
rect 7235 15365 7240 15395
rect 7200 15235 7240 15365
rect 7200 15205 7205 15235
rect 7235 15205 7240 15235
rect 7200 15200 7240 15205
rect 7280 16195 7320 16200
rect 7280 16165 7285 16195
rect 7315 16165 7320 16195
rect 7280 16035 7320 16165
rect 7280 16005 7285 16035
rect 7315 16005 7320 16035
rect 7280 15875 7320 16005
rect 7280 15845 7285 15875
rect 7315 15845 7320 15875
rect 7280 15715 7320 15845
rect 7280 15685 7285 15715
rect 7315 15685 7320 15715
rect 7280 15555 7320 15685
rect 7280 15525 7285 15555
rect 7315 15525 7320 15555
rect 7280 15395 7320 15525
rect 7280 15365 7285 15395
rect 7315 15365 7320 15395
rect 7280 15235 7320 15365
rect 7280 15205 7285 15235
rect 7315 15205 7320 15235
rect 7280 15200 7320 15205
rect 7360 16195 7400 16200
rect 7360 16165 7365 16195
rect 7395 16165 7400 16195
rect 7360 16035 7400 16165
rect 7360 16005 7365 16035
rect 7395 16005 7400 16035
rect 7360 15875 7400 16005
rect 7360 15845 7365 15875
rect 7395 15845 7400 15875
rect 7360 15715 7400 15845
rect 7360 15685 7365 15715
rect 7395 15685 7400 15715
rect 7360 15555 7400 15685
rect 7360 15525 7365 15555
rect 7395 15525 7400 15555
rect 7360 15395 7400 15525
rect 7360 15365 7365 15395
rect 7395 15365 7400 15395
rect 7360 15235 7400 15365
rect 7360 15205 7365 15235
rect 7395 15205 7400 15235
rect 7360 15200 7400 15205
rect 7440 16195 7480 16200
rect 7440 16165 7445 16195
rect 7475 16165 7480 16195
rect 7440 16035 7480 16165
rect 7440 16005 7445 16035
rect 7475 16005 7480 16035
rect 7440 15875 7480 16005
rect 7440 15845 7445 15875
rect 7475 15845 7480 15875
rect 7440 15715 7480 15845
rect 7440 15685 7445 15715
rect 7475 15685 7480 15715
rect 7440 15555 7480 15685
rect 7440 15525 7445 15555
rect 7475 15525 7480 15555
rect 7440 15395 7480 15525
rect 7440 15365 7445 15395
rect 7475 15365 7480 15395
rect 7440 15235 7480 15365
rect 7440 15205 7445 15235
rect 7475 15205 7480 15235
rect 7440 15200 7480 15205
rect 7520 16195 7560 16200
rect 7520 16165 7525 16195
rect 7555 16165 7560 16195
rect 7520 16035 7560 16165
rect 7520 16005 7525 16035
rect 7555 16005 7560 16035
rect 7520 15875 7560 16005
rect 7520 15845 7525 15875
rect 7555 15845 7560 15875
rect 7520 15715 7560 15845
rect 7520 15685 7525 15715
rect 7555 15685 7560 15715
rect 7520 15555 7560 15685
rect 7520 15525 7525 15555
rect 7555 15525 7560 15555
rect 7520 15395 7560 15525
rect 7520 15365 7525 15395
rect 7555 15365 7560 15395
rect 7520 15235 7560 15365
rect 7520 15205 7525 15235
rect 7555 15205 7560 15235
rect 7520 15200 7560 15205
rect 7600 16195 7640 16200
rect 7600 16165 7605 16195
rect 7635 16165 7640 16195
rect 7600 16035 7640 16165
rect 7600 16005 7605 16035
rect 7635 16005 7640 16035
rect 7600 15875 7640 16005
rect 7600 15845 7605 15875
rect 7635 15845 7640 15875
rect 7600 15715 7640 15845
rect 7600 15685 7605 15715
rect 7635 15685 7640 15715
rect 7600 15555 7640 15685
rect 7600 15525 7605 15555
rect 7635 15525 7640 15555
rect 7600 15395 7640 15525
rect 7600 15365 7605 15395
rect 7635 15365 7640 15395
rect 7600 15235 7640 15365
rect 7600 15205 7605 15235
rect 7635 15205 7640 15235
rect 7600 15200 7640 15205
rect 7680 16195 7720 16200
rect 7680 16165 7685 16195
rect 7715 16165 7720 16195
rect 7680 16035 7720 16165
rect 7680 16005 7685 16035
rect 7715 16005 7720 16035
rect 7680 15875 7720 16005
rect 7680 15845 7685 15875
rect 7715 15845 7720 15875
rect 7680 15715 7720 15845
rect 7680 15685 7685 15715
rect 7715 15685 7720 15715
rect 7680 15555 7720 15685
rect 7680 15525 7685 15555
rect 7715 15525 7720 15555
rect 7680 15395 7720 15525
rect 7680 15365 7685 15395
rect 7715 15365 7720 15395
rect 7680 15235 7720 15365
rect 7680 15205 7685 15235
rect 7715 15205 7720 15235
rect 7680 15200 7720 15205
rect 7760 16195 7800 16200
rect 7760 16165 7765 16195
rect 7795 16165 7800 16195
rect 7760 16035 7800 16165
rect 7760 16005 7765 16035
rect 7795 16005 7800 16035
rect 7760 15875 7800 16005
rect 7760 15845 7765 15875
rect 7795 15845 7800 15875
rect 7760 15715 7800 15845
rect 7760 15685 7765 15715
rect 7795 15685 7800 15715
rect 7760 15555 7800 15685
rect 7760 15525 7765 15555
rect 7795 15525 7800 15555
rect 7760 15395 7800 15525
rect 7760 15365 7765 15395
rect 7795 15365 7800 15395
rect 7760 15235 7800 15365
rect 7760 15205 7765 15235
rect 7795 15205 7800 15235
rect 7760 15200 7800 15205
rect 7840 16195 7880 16200
rect 7840 16165 7845 16195
rect 7875 16165 7880 16195
rect 7840 16035 7880 16165
rect 7840 16005 7845 16035
rect 7875 16005 7880 16035
rect 7840 15875 7880 16005
rect 7840 15845 7845 15875
rect 7875 15845 7880 15875
rect 7840 15715 7880 15845
rect 7840 15685 7845 15715
rect 7875 15685 7880 15715
rect 7840 15555 7880 15685
rect 7840 15525 7845 15555
rect 7875 15525 7880 15555
rect 7840 15395 7880 15525
rect 7840 15365 7845 15395
rect 7875 15365 7880 15395
rect 7840 15235 7880 15365
rect 7840 15205 7845 15235
rect 7875 15205 7880 15235
rect 7840 15200 7880 15205
rect 7920 16195 7960 16200
rect 7920 16165 7925 16195
rect 7955 16165 7960 16195
rect 7920 16035 7960 16165
rect 7920 16005 7925 16035
rect 7955 16005 7960 16035
rect 7920 15875 7960 16005
rect 7920 15845 7925 15875
rect 7955 15845 7960 15875
rect 7920 15715 7960 15845
rect 7920 15685 7925 15715
rect 7955 15685 7960 15715
rect 7920 15555 7960 15685
rect 7920 15525 7925 15555
rect 7955 15525 7960 15555
rect 7920 15395 7960 15525
rect 7920 15365 7925 15395
rect 7955 15365 7960 15395
rect 7920 15235 7960 15365
rect 7920 15205 7925 15235
rect 7955 15205 7960 15235
rect 7920 15200 7960 15205
rect 8000 16195 8040 16200
rect 8000 16165 8005 16195
rect 8035 16165 8040 16195
rect 8000 16035 8040 16165
rect 8000 16005 8005 16035
rect 8035 16005 8040 16035
rect 8000 15875 8040 16005
rect 8000 15845 8005 15875
rect 8035 15845 8040 15875
rect 8000 15715 8040 15845
rect 8000 15685 8005 15715
rect 8035 15685 8040 15715
rect 8000 15555 8040 15685
rect 8000 15525 8005 15555
rect 8035 15525 8040 15555
rect 8000 15395 8040 15525
rect 8000 15365 8005 15395
rect 8035 15365 8040 15395
rect 8000 15235 8040 15365
rect 8000 15205 8005 15235
rect 8035 15205 8040 15235
rect 8000 15200 8040 15205
rect 8080 16195 8120 16200
rect 8080 16165 8085 16195
rect 8115 16165 8120 16195
rect 8080 16035 8120 16165
rect 8080 16005 8085 16035
rect 8115 16005 8120 16035
rect 8080 15875 8120 16005
rect 8080 15845 8085 15875
rect 8115 15845 8120 15875
rect 8080 15715 8120 15845
rect 8080 15685 8085 15715
rect 8115 15685 8120 15715
rect 8080 15555 8120 15685
rect 8080 15525 8085 15555
rect 8115 15525 8120 15555
rect 8080 15395 8120 15525
rect 8080 15365 8085 15395
rect 8115 15365 8120 15395
rect 8080 15235 8120 15365
rect 8080 15205 8085 15235
rect 8115 15205 8120 15235
rect 8080 15200 8120 15205
rect 8160 16195 8200 16200
rect 8160 16165 8165 16195
rect 8195 16165 8200 16195
rect 8160 16035 8200 16165
rect 8160 16005 8165 16035
rect 8195 16005 8200 16035
rect 8160 15875 8200 16005
rect 8160 15845 8165 15875
rect 8195 15845 8200 15875
rect 8160 15715 8200 15845
rect 8160 15685 8165 15715
rect 8195 15685 8200 15715
rect 8160 15555 8200 15685
rect 8160 15525 8165 15555
rect 8195 15525 8200 15555
rect 8160 15395 8200 15525
rect 8160 15365 8165 15395
rect 8195 15365 8200 15395
rect 8160 15235 8200 15365
rect 8160 15205 8165 15235
rect 8195 15205 8200 15235
rect 8160 15200 8200 15205
rect 8240 16195 8280 16200
rect 8240 16165 8245 16195
rect 8275 16165 8280 16195
rect 8240 16035 8280 16165
rect 8240 16005 8245 16035
rect 8275 16005 8280 16035
rect 8240 15875 8280 16005
rect 8240 15845 8245 15875
rect 8275 15845 8280 15875
rect 8240 15715 8280 15845
rect 8240 15685 8245 15715
rect 8275 15685 8280 15715
rect 8240 15555 8280 15685
rect 8240 15525 8245 15555
rect 8275 15525 8280 15555
rect 8240 15395 8280 15525
rect 8240 15365 8245 15395
rect 8275 15365 8280 15395
rect 8240 15235 8280 15365
rect 8240 15205 8245 15235
rect 8275 15205 8280 15235
rect 8240 15200 8280 15205
rect 8320 16195 8360 16200
rect 8320 16165 8325 16195
rect 8355 16165 8360 16195
rect 8320 16035 8360 16165
rect 8320 16005 8325 16035
rect 8355 16005 8360 16035
rect 8320 15875 8360 16005
rect 8320 15845 8325 15875
rect 8355 15845 8360 15875
rect 8320 15715 8360 15845
rect 8320 15685 8325 15715
rect 8355 15685 8360 15715
rect 8320 15555 8360 15685
rect 8320 15525 8325 15555
rect 8355 15525 8360 15555
rect 8320 15395 8360 15525
rect 8320 15365 8325 15395
rect 8355 15365 8360 15395
rect 8320 15235 8360 15365
rect 8320 15205 8325 15235
rect 8355 15205 8360 15235
rect 8320 15200 8360 15205
rect 8400 16195 8440 16200
rect 8400 16165 8405 16195
rect 8435 16165 8440 16195
rect 8400 16035 8440 16165
rect 8400 16005 8405 16035
rect 8435 16005 8440 16035
rect 8400 15875 8440 16005
rect 8400 15845 8405 15875
rect 8435 15845 8440 15875
rect 8400 15715 8440 15845
rect 8400 15685 8405 15715
rect 8435 15685 8440 15715
rect 8400 15555 8440 15685
rect 8400 15525 8405 15555
rect 8435 15525 8440 15555
rect 8400 15395 8440 15525
rect 8400 15365 8405 15395
rect 8435 15365 8440 15395
rect 8400 15235 8440 15365
rect 8400 15205 8405 15235
rect 8435 15205 8440 15235
rect 8400 15200 8440 15205
rect 8480 16195 8520 16200
rect 8480 16165 8485 16195
rect 8515 16165 8520 16195
rect 8480 16035 8520 16165
rect 8480 16005 8485 16035
rect 8515 16005 8520 16035
rect 8480 15875 8520 16005
rect 8480 15845 8485 15875
rect 8515 15845 8520 15875
rect 8480 15715 8520 15845
rect 8480 15685 8485 15715
rect 8515 15685 8520 15715
rect 8480 15555 8520 15685
rect 8480 15525 8485 15555
rect 8515 15525 8520 15555
rect 8480 15395 8520 15525
rect 8480 15365 8485 15395
rect 8515 15365 8520 15395
rect 8480 15235 8520 15365
rect 8480 15205 8485 15235
rect 8515 15205 8520 15235
rect 8480 15200 8520 15205
rect 8560 16195 8600 16200
rect 8560 16165 8565 16195
rect 8595 16165 8600 16195
rect 8560 16035 8600 16165
rect 8560 16005 8565 16035
rect 8595 16005 8600 16035
rect 8560 15875 8600 16005
rect 8560 15845 8565 15875
rect 8595 15845 8600 15875
rect 8560 15715 8600 15845
rect 8560 15685 8565 15715
rect 8595 15685 8600 15715
rect 8560 15555 8600 15685
rect 8560 15525 8565 15555
rect 8595 15525 8600 15555
rect 8560 15395 8600 15525
rect 8560 15365 8565 15395
rect 8595 15365 8600 15395
rect 8560 15235 8600 15365
rect 8560 15205 8565 15235
rect 8595 15205 8600 15235
rect 8560 15200 8600 15205
rect 8640 16195 8680 16200
rect 8640 16165 8645 16195
rect 8675 16165 8680 16195
rect 8640 16035 8680 16165
rect 8640 16005 8645 16035
rect 8675 16005 8680 16035
rect 8640 15875 8680 16005
rect 8640 15845 8645 15875
rect 8675 15845 8680 15875
rect 8640 15715 8680 15845
rect 8640 15685 8645 15715
rect 8675 15685 8680 15715
rect 8640 15555 8680 15685
rect 8640 15525 8645 15555
rect 8675 15525 8680 15555
rect 8640 15395 8680 15525
rect 8640 15365 8645 15395
rect 8675 15365 8680 15395
rect 8640 15235 8680 15365
rect 8640 15205 8645 15235
rect 8675 15205 8680 15235
rect 8640 15200 8680 15205
rect 8720 16195 8760 16200
rect 8720 16165 8725 16195
rect 8755 16165 8760 16195
rect 8720 16035 8760 16165
rect 8720 16005 8725 16035
rect 8755 16005 8760 16035
rect 8720 15875 8760 16005
rect 8720 15845 8725 15875
rect 8755 15845 8760 15875
rect 8720 15715 8760 15845
rect 8720 15685 8725 15715
rect 8755 15685 8760 15715
rect 8720 15555 8760 15685
rect 8720 15525 8725 15555
rect 8755 15525 8760 15555
rect 8720 15395 8760 15525
rect 8720 15365 8725 15395
rect 8755 15365 8760 15395
rect 8720 15235 8760 15365
rect 8720 15205 8725 15235
rect 8755 15205 8760 15235
rect 8720 15200 8760 15205
rect 8800 16195 8840 16200
rect 8800 16165 8805 16195
rect 8835 16165 8840 16195
rect 8800 16035 8840 16165
rect 8800 16005 8805 16035
rect 8835 16005 8840 16035
rect 8800 15875 8840 16005
rect 8800 15845 8805 15875
rect 8835 15845 8840 15875
rect 8800 15715 8840 15845
rect 8800 15685 8805 15715
rect 8835 15685 8840 15715
rect 8800 15555 8840 15685
rect 8800 15525 8805 15555
rect 8835 15525 8840 15555
rect 8800 15395 8840 15525
rect 8800 15365 8805 15395
rect 8835 15365 8840 15395
rect 8800 15235 8840 15365
rect 8800 15205 8805 15235
rect 8835 15205 8840 15235
rect 8800 15200 8840 15205
rect 8880 16195 8920 16200
rect 8880 16165 8885 16195
rect 8915 16165 8920 16195
rect 8880 16035 8920 16165
rect 8880 16005 8885 16035
rect 8915 16005 8920 16035
rect 8880 15875 8920 16005
rect 8880 15845 8885 15875
rect 8915 15845 8920 15875
rect 8880 15715 8920 15845
rect 8880 15685 8885 15715
rect 8915 15685 8920 15715
rect 8880 15555 8920 15685
rect 8880 15525 8885 15555
rect 8915 15525 8920 15555
rect 8880 15395 8920 15525
rect 8880 15365 8885 15395
rect 8915 15365 8920 15395
rect 8880 15235 8920 15365
rect 8880 15205 8885 15235
rect 8915 15205 8920 15235
rect 8880 15200 8920 15205
rect 8960 16195 9000 16200
rect 8960 16165 8965 16195
rect 8995 16165 9000 16195
rect 8960 16035 9000 16165
rect 8960 16005 8965 16035
rect 8995 16005 9000 16035
rect 8960 15875 9000 16005
rect 8960 15845 8965 15875
rect 8995 15845 9000 15875
rect 8960 15715 9000 15845
rect 8960 15685 8965 15715
rect 8995 15685 9000 15715
rect 8960 15555 9000 15685
rect 8960 15525 8965 15555
rect 8995 15525 9000 15555
rect 8960 15395 9000 15525
rect 8960 15365 8965 15395
rect 8995 15365 9000 15395
rect 8960 15235 9000 15365
rect 8960 15205 8965 15235
rect 8995 15205 9000 15235
rect 8960 15200 9000 15205
rect 9040 16195 9080 16200
rect 9040 16165 9045 16195
rect 9075 16165 9080 16195
rect 9040 16035 9080 16165
rect 9040 16005 9045 16035
rect 9075 16005 9080 16035
rect 9040 15875 9080 16005
rect 9040 15845 9045 15875
rect 9075 15845 9080 15875
rect 9040 15715 9080 15845
rect 9040 15685 9045 15715
rect 9075 15685 9080 15715
rect 9040 15555 9080 15685
rect 9040 15525 9045 15555
rect 9075 15525 9080 15555
rect 9040 15395 9080 15525
rect 9040 15365 9045 15395
rect 9075 15365 9080 15395
rect 9040 15235 9080 15365
rect 9040 15205 9045 15235
rect 9075 15205 9080 15235
rect 9040 15200 9080 15205
rect 9120 16195 9160 16200
rect 9120 16165 9125 16195
rect 9155 16165 9160 16195
rect 9120 16035 9160 16165
rect 9120 16005 9125 16035
rect 9155 16005 9160 16035
rect 9120 15875 9160 16005
rect 9120 15845 9125 15875
rect 9155 15845 9160 15875
rect 9120 15715 9160 15845
rect 9120 15685 9125 15715
rect 9155 15685 9160 15715
rect 9120 15555 9160 15685
rect 9120 15525 9125 15555
rect 9155 15525 9160 15555
rect 9120 15395 9160 15525
rect 9120 15365 9125 15395
rect 9155 15365 9160 15395
rect 9120 15235 9160 15365
rect 9120 15205 9125 15235
rect 9155 15205 9160 15235
rect 9120 15200 9160 15205
rect 9200 16195 9240 16200
rect 9200 16165 9205 16195
rect 9235 16165 9240 16195
rect 9200 16035 9240 16165
rect 9200 16005 9205 16035
rect 9235 16005 9240 16035
rect 9200 15875 9240 16005
rect 9200 15845 9205 15875
rect 9235 15845 9240 15875
rect 9200 15715 9240 15845
rect 9200 15685 9205 15715
rect 9235 15685 9240 15715
rect 9200 15555 9240 15685
rect 9200 15525 9205 15555
rect 9235 15525 9240 15555
rect 9200 15395 9240 15525
rect 9200 15365 9205 15395
rect 9235 15365 9240 15395
rect 9200 15235 9240 15365
rect 9200 15205 9205 15235
rect 9235 15205 9240 15235
rect 9200 15200 9240 15205
rect 9280 16195 9320 16200
rect 9280 16165 9285 16195
rect 9315 16165 9320 16195
rect 9280 16035 9320 16165
rect 9280 16005 9285 16035
rect 9315 16005 9320 16035
rect 9280 15875 9320 16005
rect 9280 15845 9285 15875
rect 9315 15845 9320 15875
rect 9280 15715 9320 15845
rect 9280 15685 9285 15715
rect 9315 15685 9320 15715
rect 9280 15555 9320 15685
rect 9280 15525 9285 15555
rect 9315 15525 9320 15555
rect 9280 15395 9320 15525
rect 9280 15365 9285 15395
rect 9315 15365 9320 15395
rect 9280 15235 9320 15365
rect 9280 15205 9285 15235
rect 9315 15205 9320 15235
rect 9280 15200 9320 15205
rect 9360 16195 9400 16200
rect 9360 16165 9365 16195
rect 9395 16165 9400 16195
rect 9360 16035 9400 16165
rect 9360 16005 9365 16035
rect 9395 16005 9400 16035
rect 9360 15875 9400 16005
rect 9360 15845 9365 15875
rect 9395 15845 9400 15875
rect 9360 15715 9400 15845
rect 9360 15685 9365 15715
rect 9395 15685 9400 15715
rect 9360 15555 9400 15685
rect 9360 15525 9365 15555
rect 9395 15525 9400 15555
rect 9360 15395 9400 15525
rect 9360 15365 9365 15395
rect 9395 15365 9400 15395
rect 9360 15235 9400 15365
rect 9360 15205 9365 15235
rect 9395 15205 9400 15235
rect 9360 15200 9400 15205
rect 9440 16195 9480 16200
rect 9440 16165 9445 16195
rect 9475 16165 9480 16195
rect 9440 16035 9480 16165
rect 9440 16005 9445 16035
rect 9475 16005 9480 16035
rect 9440 15875 9480 16005
rect 9440 15845 9445 15875
rect 9475 15845 9480 15875
rect 9440 15715 9480 15845
rect 9440 15685 9445 15715
rect 9475 15685 9480 15715
rect 9440 15555 9480 15685
rect 9440 15525 9445 15555
rect 9475 15525 9480 15555
rect 9440 15395 9480 15525
rect 9440 15365 9445 15395
rect 9475 15365 9480 15395
rect 9440 15235 9480 15365
rect 9440 15205 9445 15235
rect 9475 15205 9480 15235
rect 9440 15200 9480 15205
rect 6240 15155 6280 15160
rect 6240 15125 6245 15155
rect 6275 15125 6280 15155
rect 6240 14995 6280 15125
rect 6240 14965 6245 14995
rect 6275 14965 6280 14995
rect 6240 14960 6280 14965
rect 6320 15155 6360 15160
rect 6320 15125 6325 15155
rect 6355 15125 6360 15155
rect 6320 14995 6360 15125
rect 6320 14965 6325 14995
rect 6355 14965 6360 14995
rect 6320 14960 6360 14965
rect 6400 15155 6440 15160
rect 6400 15125 6405 15155
rect 6435 15125 6440 15155
rect 6400 14995 6440 15125
rect 6400 14965 6405 14995
rect 6435 14965 6440 14995
rect 6400 14960 6440 14965
rect 6480 15155 6520 15160
rect 6480 15125 6485 15155
rect 6515 15125 6520 15155
rect 6480 14995 6520 15125
rect 6480 14965 6485 14995
rect 6515 14965 6520 14995
rect 6480 14960 6520 14965
rect 6560 15155 6600 15160
rect 6560 15125 6565 15155
rect 6595 15125 6600 15155
rect 6560 14995 6600 15125
rect 6560 14965 6565 14995
rect 6595 14965 6600 14995
rect 6560 14960 6600 14965
rect 6640 15155 6680 15160
rect 6640 15125 6645 15155
rect 6675 15125 6680 15155
rect 6640 14995 6680 15125
rect 6640 14965 6645 14995
rect 6675 14965 6680 14995
rect 6640 14960 6680 14965
rect 6720 15155 6760 15160
rect 6720 15125 6725 15155
rect 6755 15125 6760 15155
rect 6720 14995 6760 15125
rect 6720 14965 6725 14995
rect 6755 14965 6760 14995
rect 6720 14960 6760 14965
rect 6800 15155 6840 15160
rect 6800 15125 6805 15155
rect 6835 15125 6840 15155
rect 6800 14995 6840 15125
rect 6800 14965 6805 14995
rect 6835 14965 6840 14995
rect 6800 14960 6840 14965
rect 6880 15155 6920 15160
rect 6880 15125 6885 15155
rect 6915 15125 6920 15155
rect 6880 14995 6920 15125
rect 6880 14965 6885 14995
rect 6915 14965 6920 14995
rect 6880 14960 6920 14965
rect 6960 15155 7000 15160
rect 6960 15125 6965 15155
rect 6995 15125 7000 15155
rect 6960 14995 7000 15125
rect 6960 14965 6965 14995
rect 6995 14965 7000 14995
rect 6960 14960 7000 14965
rect 7040 15155 7080 15160
rect 7040 15125 7045 15155
rect 7075 15125 7080 15155
rect 7040 14995 7080 15125
rect 7040 14965 7045 14995
rect 7075 14965 7080 14995
rect 7040 14960 7080 14965
rect 7120 15155 7160 15160
rect 7120 15125 7125 15155
rect 7155 15125 7160 15155
rect 7120 14995 7160 15125
rect 7120 14965 7125 14995
rect 7155 14965 7160 14995
rect 7120 14960 7160 14965
rect 7200 15155 7240 15160
rect 7200 15125 7205 15155
rect 7235 15125 7240 15155
rect 7200 14995 7240 15125
rect 7200 14965 7205 14995
rect 7235 14965 7240 14995
rect 7200 14960 7240 14965
rect 7280 15155 7320 15160
rect 7280 15125 7285 15155
rect 7315 15125 7320 15155
rect 7280 14995 7320 15125
rect 7280 14965 7285 14995
rect 7315 14965 7320 14995
rect 7280 14960 7320 14965
rect 7360 15155 7400 15160
rect 7360 15125 7365 15155
rect 7395 15125 7400 15155
rect 7360 14995 7400 15125
rect 7360 14965 7365 14995
rect 7395 14965 7400 14995
rect 7360 14960 7400 14965
rect 7440 15155 7480 15160
rect 7440 15125 7445 15155
rect 7475 15125 7480 15155
rect 7440 14995 7480 15125
rect 7440 14965 7445 14995
rect 7475 14965 7480 14995
rect 7440 14960 7480 14965
rect 7520 15155 7560 15160
rect 7520 15125 7525 15155
rect 7555 15125 7560 15155
rect 7520 14995 7560 15125
rect 7520 14965 7525 14995
rect 7555 14965 7560 14995
rect 7520 14960 7560 14965
rect 7600 15155 7640 15160
rect 7600 15125 7605 15155
rect 7635 15125 7640 15155
rect 7600 14995 7640 15125
rect 7600 14965 7605 14995
rect 7635 14965 7640 14995
rect 7600 14960 7640 14965
rect 7680 15155 7720 15160
rect 7680 15125 7685 15155
rect 7715 15125 7720 15155
rect 7680 14995 7720 15125
rect 7680 14965 7685 14995
rect 7715 14965 7720 14995
rect 7680 14960 7720 14965
rect 7760 15155 7800 15160
rect 7760 15125 7765 15155
rect 7795 15125 7800 15155
rect 7760 14995 7800 15125
rect 7760 14965 7765 14995
rect 7795 14965 7800 14995
rect 7760 14960 7800 14965
rect 7840 15155 7880 15160
rect 7840 15125 7845 15155
rect 7875 15125 7880 15155
rect 7840 14995 7880 15125
rect 7840 14965 7845 14995
rect 7875 14965 7880 14995
rect 7840 14960 7880 14965
rect 7920 15155 7960 15160
rect 7920 15125 7925 15155
rect 7955 15125 7960 15155
rect 7920 14995 7960 15125
rect 7920 14965 7925 14995
rect 7955 14965 7960 14995
rect 7920 14960 7960 14965
rect 8000 15155 8040 15160
rect 8000 15125 8005 15155
rect 8035 15125 8040 15155
rect 8000 14995 8040 15125
rect 8000 14965 8005 14995
rect 8035 14965 8040 14995
rect 8000 14960 8040 14965
rect 8080 15155 8120 15160
rect 8080 15125 8085 15155
rect 8115 15125 8120 15155
rect 8080 14995 8120 15125
rect 8080 14965 8085 14995
rect 8115 14965 8120 14995
rect 8080 14960 8120 14965
rect 8160 15155 8200 15160
rect 8160 15125 8165 15155
rect 8195 15125 8200 15155
rect 8160 14995 8200 15125
rect 8160 14965 8165 14995
rect 8195 14965 8200 14995
rect 8160 14960 8200 14965
rect 8240 15155 8280 15160
rect 8240 15125 8245 15155
rect 8275 15125 8280 15155
rect 8240 14995 8280 15125
rect 8240 14965 8245 14995
rect 8275 14965 8280 14995
rect 8240 14960 8280 14965
rect 8320 15155 8360 15160
rect 8320 15125 8325 15155
rect 8355 15125 8360 15155
rect 8320 14995 8360 15125
rect 8320 14965 8325 14995
rect 8355 14965 8360 14995
rect 8320 14960 8360 14965
rect 8400 15155 8440 15160
rect 8400 15125 8405 15155
rect 8435 15125 8440 15155
rect 8400 14995 8440 15125
rect 8400 14965 8405 14995
rect 8435 14965 8440 14995
rect 8400 14960 8440 14965
rect 8480 15155 8520 15160
rect 8480 15125 8485 15155
rect 8515 15125 8520 15155
rect 8480 14995 8520 15125
rect 8480 14965 8485 14995
rect 8515 14965 8520 14995
rect 8480 14960 8520 14965
rect 8560 15155 8600 15160
rect 8560 15125 8565 15155
rect 8595 15125 8600 15155
rect 8560 14995 8600 15125
rect 8560 14965 8565 14995
rect 8595 14965 8600 14995
rect 8560 14960 8600 14965
rect 8640 15155 8680 15160
rect 8640 15125 8645 15155
rect 8675 15125 8680 15155
rect 8640 14995 8680 15125
rect 8640 14965 8645 14995
rect 8675 14965 8680 14995
rect 8640 14960 8680 14965
rect 8720 15155 8760 15160
rect 8720 15125 8725 15155
rect 8755 15125 8760 15155
rect 8720 14995 8760 15125
rect 8720 14965 8725 14995
rect 8755 14965 8760 14995
rect 8720 14960 8760 14965
rect 8800 15155 8840 15160
rect 8800 15125 8805 15155
rect 8835 15125 8840 15155
rect 8800 14995 8840 15125
rect 8800 14965 8805 14995
rect 8835 14965 8840 14995
rect 8800 14960 8840 14965
rect 8880 15155 8920 15160
rect 8880 15125 8885 15155
rect 8915 15125 8920 15155
rect 8880 14995 8920 15125
rect 8880 14965 8885 14995
rect 8915 14965 8920 14995
rect 8880 14960 8920 14965
rect 8960 15155 9000 15160
rect 8960 15125 8965 15155
rect 8995 15125 9000 15155
rect 8960 14995 9000 15125
rect 8960 14965 8965 14995
rect 8995 14965 9000 14995
rect 8960 14960 9000 14965
rect 9040 15155 9080 15160
rect 9040 15125 9045 15155
rect 9075 15125 9080 15155
rect 9040 14995 9080 15125
rect 9040 14965 9045 14995
rect 9075 14965 9080 14995
rect 9040 14960 9080 14965
rect 9120 15155 9160 15160
rect 9120 15125 9125 15155
rect 9155 15125 9160 15155
rect 9120 14995 9160 15125
rect 9120 14965 9125 14995
rect 9155 14965 9160 14995
rect 9120 14960 9160 14965
rect 9200 15155 9240 15160
rect 9200 15125 9205 15155
rect 9235 15125 9240 15155
rect 9200 14995 9240 15125
rect 9200 14965 9205 14995
rect 9235 14965 9240 14995
rect 9200 14960 9240 14965
rect 9280 15155 9320 15160
rect 9280 15125 9285 15155
rect 9315 15125 9320 15155
rect 9280 14995 9320 15125
rect 9280 14965 9285 14995
rect 9315 14965 9320 14995
rect 9280 14960 9320 14965
rect 9360 15155 9400 15160
rect 9360 15125 9365 15155
rect 9395 15125 9400 15155
rect 9360 14995 9400 15125
rect 9360 14965 9365 14995
rect 9395 14965 9400 14995
rect 9360 14960 9400 14965
rect 9440 15155 9480 15160
rect 9440 15125 9445 15155
rect 9475 15125 9480 15155
rect 9440 14995 9480 15125
rect 9440 14965 9445 14995
rect 9475 14965 9480 14995
rect 9440 14960 9480 14965
rect 6160 14885 6165 14915
rect 6195 14885 6200 14915
rect 6160 14755 6200 14885
rect 6160 14725 6165 14755
rect 6195 14725 6200 14755
rect 6160 14680 6200 14725
rect 6240 14915 6280 14920
rect 6240 14885 6245 14915
rect 6275 14885 6280 14915
rect 6240 14755 6280 14885
rect 6240 14725 6245 14755
rect 6275 14725 6280 14755
rect 6240 14720 6280 14725
rect 6320 14915 6360 14920
rect 6320 14885 6325 14915
rect 6355 14885 6360 14915
rect 6320 14755 6360 14885
rect 6320 14725 6325 14755
rect 6355 14725 6360 14755
rect 6320 14720 6360 14725
rect 6400 14915 6440 14920
rect 6400 14885 6405 14915
rect 6435 14885 6440 14915
rect 6400 14755 6440 14885
rect 6400 14725 6405 14755
rect 6435 14725 6440 14755
rect 6400 14720 6440 14725
rect 6480 14915 6520 14920
rect 6480 14885 6485 14915
rect 6515 14885 6520 14915
rect 6480 14755 6520 14885
rect 6480 14725 6485 14755
rect 6515 14725 6520 14755
rect 6480 14720 6520 14725
rect 6560 14915 6600 14920
rect 6560 14885 6565 14915
rect 6595 14885 6600 14915
rect 6560 14755 6600 14885
rect 6560 14725 6565 14755
rect 6595 14725 6600 14755
rect 6560 14720 6600 14725
rect 6640 14915 6680 14920
rect 6640 14885 6645 14915
rect 6675 14885 6680 14915
rect 6640 14755 6680 14885
rect 6640 14725 6645 14755
rect 6675 14725 6680 14755
rect 6640 14720 6680 14725
rect 6720 14915 6760 14920
rect 6720 14885 6725 14915
rect 6755 14885 6760 14915
rect 6720 14755 6760 14885
rect 6720 14725 6725 14755
rect 6755 14725 6760 14755
rect 6720 14720 6760 14725
rect 6800 14915 6840 14920
rect 6800 14885 6805 14915
rect 6835 14885 6840 14915
rect 6800 14755 6840 14885
rect 6800 14725 6805 14755
rect 6835 14725 6840 14755
rect 6800 14720 6840 14725
rect 6880 14915 6920 14920
rect 6880 14885 6885 14915
rect 6915 14885 6920 14915
rect 6880 14755 6920 14885
rect 6880 14725 6885 14755
rect 6915 14725 6920 14755
rect 6880 14720 6920 14725
rect 6960 14915 7000 14920
rect 6960 14885 6965 14915
rect 6995 14885 7000 14915
rect 6960 14755 7000 14885
rect 6960 14725 6965 14755
rect 6995 14725 7000 14755
rect 6960 14720 7000 14725
rect 7040 14915 7080 14920
rect 7040 14885 7045 14915
rect 7075 14885 7080 14915
rect 7040 14755 7080 14885
rect 7040 14725 7045 14755
rect 7075 14725 7080 14755
rect 7040 14720 7080 14725
rect 7120 14915 7160 14920
rect 7120 14885 7125 14915
rect 7155 14885 7160 14915
rect 7120 14755 7160 14885
rect 7120 14725 7125 14755
rect 7155 14725 7160 14755
rect 7120 14720 7160 14725
rect 7200 14915 7240 14920
rect 7200 14885 7205 14915
rect 7235 14885 7240 14915
rect 7200 14755 7240 14885
rect 7200 14725 7205 14755
rect 7235 14725 7240 14755
rect 7200 14720 7240 14725
rect 7280 14915 7320 14920
rect 7280 14885 7285 14915
rect 7315 14885 7320 14915
rect 7280 14755 7320 14885
rect 7280 14725 7285 14755
rect 7315 14725 7320 14755
rect 7280 14720 7320 14725
rect 7360 14915 7400 14920
rect 7360 14885 7365 14915
rect 7395 14885 7400 14915
rect 7360 14755 7400 14885
rect 7360 14725 7365 14755
rect 7395 14725 7400 14755
rect 7360 14720 7400 14725
rect 7440 14915 7480 14920
rect 7440 14885 7445 14915
rect 7475 14885 7480 14915
rect 7440 14755 7480 14885
rect 7440 14725 7445 14755
rect 7475 14725 7480 14755
rect 7440 14720 7480 14725
rect 7520 14915 7560 14920
rect 7520 14885 7525 14915
rect 7555 14885 7560 14915
rect 7520 14755 7560 14885
rect 7520 14725 7525 14755
rect 7555 14725 7560 14755
rect 7520 14720 7560 14725
rect 7600 14915 7640 14920
rect 7600 14885 7605 14915
rect 7635 14885 7640 14915
rect 7600 14755 7640 14885
rect 7600 14725 7605 14755
rect 7635 14725 7640 14755
rect 7600 14720 7640 14725
rect 7680 14915 7720 14920
rect 7680 14885 7685 14915
rect 7715 14885 7720 14915
rect 7680 14755 7720 14885
rect 7680 14725 7685 14755
rect 7715 14725 7720 14755
rect 7680 14720 7720 14725
rect 7760 14915 7800 14920
rect 7760 14885 7765 14915
rect 7795 14885 7800 14915
rect 7760 14755 7800 14885
rect 7760 14725 7765 14755
rect 7795 14725 7800 14755
rect 7760 14720 7800 14725
rect 7840 14915 7880 14920
rect 7840 14885 7845 14915
rect 7875 14885 7880 14915
rect 7840 14755 7880 14885
rect 7840 14725 7845 14755
rect 7875 14725 7880 14755
rect 7840 14720 7880 14725
rect 7920 14915 7960 14920
rect 7920 14885 7925 14915
rect 7955 14885 7960 14915
rect 7920 14755 7960 14885
rect 7920 14725 7925 14755
rect 7955 14725 7960 14755
rect 7920 14720 7960 14725
rect 8000 14915 8040 14920
rect 8000 14885 8005 14915
rect 8035 14885 8040 14915
rect 8000 14755 8040 14885
rect 8000 14725 8005 14755
rect 8035 14725 8040 14755
rect 8000 14720 8040 14725
rect 8080 14915 8120 14920
rect 8080 14885 8085 14915
rect 8115 14885 8120 14915
rect 8080 14755 8120 14885
rect 8080 14725 8085 14755
rect 8115 14725 8120 14755
rect 8080 14720 8120 14725
rect 8160 14915 8200 14920
rect 8160 14885 8165 14915
rect 8195 14885 8200 14915
rect 8160 14755 8200 14885
rect 8160 14725 8165 14755
rect 8195 14725 8200 14755
rect 8160 14720 8200 14725
rect 8240 14915 8280 14920
rect 8240 14885 8245 14915
rect 8275 14885 8280 14915
rect 8240 14755 8280 14885
rect 8240 14725 8245 14755
rect 8275 14725 8280 14755
rect 8240 14720 8280 14725
rect 8320 14915 8360 14920
rect 8320 14885 8325 14915
rect 8355 14885 8360 14915
rect 8320 14755 8360 14885
rect 8320 14725 8325 14755
rect 8355 14725 8360 14755
rect 8320 14720 8360 14725
rect 8400 14915 8440 14920
rect 8400 14885 8405 14915
rect 8435 14885 8440 14915
rect 8400 14755 8440 14885
rect 8400 14725 8405 14755
rect 8435 14725 8440 14755
rect 8400 14720 8440 14725
rect 8480 14915 8520 14920
rect 8480 14885 8485 14915
rect 8515 14885 8520 14915
rect 8480 14755 8520 14885
rect 8480 14725 8485 14755
rect 8515 14725 8520 14755
rect 8480 14720 8520 14725
rect 8560 14915 8600 14920
rect 8560 14885 8565 14915
rect 8595 14885 8600 14915
rect 8560 14755 8600 14885
rect 8560 14725 8565 14755
rect 8595 14725 8600 14755
rect 8560 14720 8600 14725
rect 8640 14915 8680 14920
rect 8640 14885 8645 14915
rect 8675 14885 8680 14915
rect 8640 14755 8680 14885
rect 8640 14725 8645 14755
rect 8675 14725 8680 14755
rect 8640 14720 8680 14725
rect 8720 14915 8760 14920
rect 8720 14885 8725 14915
rect 8755 14885 8760 14915
rect 8720 14755 8760 14885
rect 8720 14725 8725 14755
rect 8755 14725 8760 14755
rect 8720 14720 8760 14725
rect 8800 14915 8840 14920
rect 8800 14885 8805 14915
rect 8835 14885 8840 14915
rect 8800 14755 8840 14885
rect 8800 14725 8805 14755
rect 8835 14725 8840 14755
rect 8800 14720 8840 14725
rect 8880 14915 8920 14920
rect 8880 14885 8885 14915
rect 8915 14885 8920 14915
rect 8880 14755 8920 14885
rect 8880 14725 8885 14755
rect 8915 14725 8920 14755
rect 8880 14720 8920 14725
rect 8960 14915 9000 14920
rect 8960 14885 8965 14915
rect 8995 14885 9000 14915
rect 8960 14755 9000 14885
rect 8960 14725 8965 14755
rect 8995 14725 9000 14755
rect 8960 14720 9000 14725
rect 9040 14915 9080 14920
rect 9040 14885 9045 14915
rect 9075 14885 9080 14915
rect 9040 14755 9080 14885
rect 9040 14725 9045 14755
rect 9075 14725 9080 14755
rect 9040 14720 9080 14725
rect 9120 14915 9160 14920
rect 9120 14885 9125 14915
rect 9155 14885 9160 14915
rect 9120 14755 9160 14885
rect 9120 14725 9125 14755
rect 9155 14725 9160 14755
rect 9120 14720 9160 14725
rect 9200 14915 9240 14920
rect 9200 14885 9205 14915
rect 9235 14885 9240 14915
rect 9200 14755 9240 14885
rect 9200 14725 9205 14755
rect 9235 14725 9240 14755
rect 9200 14720 9240 14725
rect 9280 14915 9320 14920
rect 9280 14885 9285 14915
rect 9315 14885 9320 14915
rect 9280 14755 9320 14885
rect 9280 14725 9285 14755
rect 9315 14725 9320 14755
rect 9280 14720 9320 14725
rect 9360 14915 9400 14920
rect 9360 14885 9365 14915
rect 9395 14885 9400 14915
rect 9360 14755 9400 14885
rect 9360 14725 9365 14755
rect 9395 14725 9400 14755
rect 9360 14720 9400 14725
rect 9440 14915 9480 14920
rect 9440 14885 9445 14915
rect 9475 14885 9480 14915
rect 9440 14755 9480 14885
rect 9440 14725 9445 14755
rect 9475 14725 9480 14755
rect 9440 14720 9480 14725
rect 9520 14720 9560 16485
rect 9600 16835 9640 18680
rect 9600 16805 9605 16835
rect 9635 16805 9640 16835
rect 9600 16595 9640 16805
rect 9600 16565 9605 16595
rect 9635 16565 9640 16595
rect 9600 14720 9640 16565
rect 9680 16915 9720 18680
rect 9680 16885 9685 16915
rect 9715 16885 9720 16915
rect 9680 16755 9720 16885
rect 9680 16725 9685 16755
rect 9715 16725 9720 16755
rect 9680 16675 9720 16725
rect 9680 16645 9685 16675
rect 9715 16645 9720 16675
rect 9680 16515 9720 16645
rect 9680 16485 9685 16515
rect 9715 16485 9720 16515
rect 9680 14720 9720 16485
rect 9760 17155 9800 18680
rect 9760 17125 9765 17155
rect 9795 17125 9800 17155
rect 9760 16995 9800 17125
rect 9760 16965 9765 16995
rect 9795 16965 9800 16995
rect 9760 16435 9800 16965
rect 9760 16405 9765 16435
rect 9795 16405 9800 16435
rect 9760 16275 9800 16405
rect 9760 16245 9765 16275
rect 9795 16245 9800 16275
rect 9760 14720 9800 16245
rect 9840 17075 9880 18680
rect 9840 17045 9845 17075
rect 9875 17045 9880 17075
rect 9840 16355 9880 17045
rect 9840 16325 9845 16355
rect 9875 16325 9880 16355
rect 9840 14720 9880 16325
rect 9920 17155 9960 18680
rect 9920 17125 9925 17155
rect 9955 17125 9960 17155
rect 9920 16995 9960 17125
rect 9920 16965 9925 16995
rect 9955 16965 9960 16995
rect 9920 16435 9960 16965
rect 9920 16405 9925 16435
rect 9955 16405 9960 16435
rect 9920 16275 9960 16405
rect 9920 16245 9925 16275
rect 9955 16245 9960 16275
rect 9920 14720 9960 16245
rect 10000 18195 10040 18680
rect 10000 18165 10005 18195
rect 10035 18165 10040 18195
rect 10000 18035 10040 18165
rect 10000 18005 10005 18035
rect 10035 18005 10040 18035
rect 10000 17875 10040 18005
rect 10000 17845 10005 17875
rect 10035 17845 10040 17875
rect 10000 17715 10040 17845
rect 10000 17685 10005 17715
rect 10035 17685 10040 17715
rect 10000 17555 10040 17685
rect 10000 17525 10005 17555
rect 10035 17525 10040 17555
rect 10000 17395 10040 17525
rect 10000 17365 10005 17395
rect 10035 17365 10040 17395
rect 10000 17235 10040 17365
rect 10000 17205 10005 17235
rect 10035 17205 10040 17235
rect 10000 16195 10040 17205
rect 10000 16165 10005 16195
rect 10035 16165 10040 16195
rect 10000 16035 10040 16165
rect 10000 16005 10005 16035
rect 10035 16005 10040 16035
rect 10000 15875 10040 16005
rect 10000 15845 10005 15875
rect 10035 15845 10040 15875
rect 10000 15715 10040 15845
rect 10000 15685 10005 15715
rect 10035 15685 10040 15715
rect 10000 15555 10040 15685
rect 10000 15525 10005 15555
rect 10035 15525 10040 15555
rect 10000 15395 10040 15525
rect 10000 15365 10005 15395
rect 10035 15365 10040 15395
rect 10000 15235 10040 15365
rect 10000 15205 10005 15235
rect 10035 15205 10040 15235
rect 10000 14720 10040 15205
rect 10080 17315 10120 18680
rect 10080 17285 10085 17315
rect 10115 17285 10120 17315
rect 10080 16115 10120 17285
rect 10080 16085 10085 16115
rect 10115 16085 10120 16115
rect 10080 14720 10120 16085
rect 10160 18195 10200 18680
rect 10160 18165 10165 18195
rect 10195 18165 10200 18195
rect 10160 18035 10200 18165
rect 10160 18005 10165 18035
rect 10195 18005 10200 18035
rect 10160 17875 10200 18005
rect 10160 17845 10165 17875
rect 10195 17845 10200 17875
rect 10160 17715 10200 17845
rect 10160 17685 10165 17715
rect 10195 17685 10200 17715
rect 10160 17555 10200 17685
rect 10160 17525 10165 17555
rect 10195 17525 10200 17555
rect 10160 17395 10200 17525
rect 10160 17365 10165 17395
rect 10195 17365 10200 17395
rect 10160 17235 10200 17365
rect 10160 17205 10165 17235
rect 10195 17205 10200 17235
rect 10160 16195 10200 17205
rect 10160 16165 10165 16195
rect 10195 16165 10200 16195
rect 10160 16035 10200 16165
rect 10160 16005 10165 16035
rect 10195 16005 10200 16035
rect 10160 15875 10200 16005
rect 10160 15845 10165 15875
rect 10195 15845 10200 15875
rect 10160 15715 10200 15845
rect 10160 15685 10165 15715
rect 10195 15685 10200 15715
rect 10160 15555 10200 15685
rect 10160 15525 10165 15555
rect 10195 15525 10200 15555
rect 10160 15395 10200 15525
rect 10160 15365 10165 15395
rect 10195 15365 10200 15395
rect 10160 15235 10200 15365
rect 10160 15205 10165 15235
rect 10195 15205 10200 15235
rect 10160 14720 10200 15205
rect 10240 17475 10280 18680
rect 10240 17445 10245 17475
rect 10275 17445 10280 17475
rect 10240 15955 10280 17445
rect 10240 15925 10245 15955
rect 10275 15925 10280 15955
rect 10240 14720 10280 15925
rect 10320 18195 10360 18680
rect 10320 18165 10325 18195
rect 10355 18165 10360 18195
rect 10320 18035 10360 18165
rect 10320 18005 10325 18035
rect 10355 18005 10360 18035
rect 10320 17875 10360 18005
rect 10320 17845 10325 17875
rect 10355 17845 10360 17875
rect 10320 17715 10360 17845
rect 10320 17685 10325 17715
rect 10355 17685 10360 17715
rect 10320 17555 10360 17685
rect 10320 17525 10325 17555
rect 10355 17525 10360 17555
rect 10320 17395 10360 17525
rect 10320 17365 10325 17395
rect 10355 17365 10360 17395
rect 10320 17235 10360 17365
rect 10320 17205 10325 17235
rect 10355 17205 10360 17235
rect 10320 16195 10360 17205
rect 10320 16165 10325 16195
rect 10355 16165 10360 16195
rect 10320 16035 10360 16165
rect 10320 16005 10325 16035
rect 10355 16005 10360 16035
rect 10320 15875 10360 16005
rect 10320 15845 10325 15875
rect 10355 15845 10360 15875
rect 10320 15715 10360 15845
rect 10320 15685 10325 15715
rect 10355 15685 10360 15715
rect 10320 15555 10360 15685
rect 10320 15525 10325 15555
rect 10355 15525 10360 15555
rect 10320 15395 10360 15525
rect 10320 15365 10325 15395
rect 10355 15365 10360 15395
rect 10320 15235 10360 15365
rect 10320 15205 10325 15235
rect 10355 15205 10360 15235
rect 10320 14720 10360 15205
rect 10400 17635 10440 18680
rect 10400 17605 10405 17635
rect 10435 17605 10440 17635
rect 10400 15795 10440 17605
rect 10400 15765 10405 15795
rect 10435 15765 10440 15795
rect 10400 14720 10440 15765
rect 10480 18195 10520 18680
rect 10480 18165 10485 18195
rect 10515 18165 10520 18195
rect 10480 18035 10520 18165
rect 10480 18005 10485 18035
rect 10515 18005 10520 18035
rect 10480 17875 10520 18005
rect 10480 17845 10485 17875
rect 10515 17845 10520 17875
rect 10480 17715 10520 17845
rect 10480 17685 10485 17715
rect 10515 17685 10520 17715
rect 10480 17555 10520 17685
rect 10480 17525 10485 17555
rect 10515 17525 10520 17555
rect 10480 17395 10520 17525
rect 10480 17365 10485 17395
rect 10515 17365 10520 17395
rect 10480 17235 10520 17365
rect 10480 17205 10485 17235
rect 10515 17205 10520 17235
rect 10480 16195 10520 17205
rect 10480 16165 10485 16195
rect 10515 16165 10520 16195
rect 10480 16035 10520 16165
rect 10480 16005 10485 16035
rect 10515 16005 10520 16035
rect 10480 15875 10520 16005
rect 10480 15845 10485 15875
rect 10515 15845 10520 15875
rect 10480 15715 10520 15845
rect 10480 15685 10485 15715
rect 10515 15685 10520 15715
rect 10480 15555 10520 15685
rect 10480 15525 10485 15555
rect 10515 15525 10520 15555
rect 10480 15395 10520 15525
rect 10480 15365 10485 15395
rect 10515 15365 10520 15395
rect 10480 15235 10520 15365
rect 10480 15205 10485 15235
rect 10515 15205 10520 15235
rect 10480 14720 10520 15205
rect 10560 17795 10600 18680
rect 10560 17765 10565 17795
rect 10595 17765 10600 17795
rect 10560 15635 10600 17765
rect 10560 15605 10565 15635
rect 10595 15605 10600 15635
rect 10560 14720 10600 15605
rect 10640 18195 10680 18680
rect 10640 18165 10645 18195
rect 10675 18165 10680 18195
rect 10640 18035 10680 18165
rect 10640 18005 10645 18035
rect 10675 18005 10680 18035
rect 10640 17875 10680 18005
rect 10640 17845 10645 17875
rect 10675 17845 10680 17875
rect 10640 17715 10680 17845
rect 10640 17685 10645 17715
rect 10675 17685 10680 17715
rect 10640 17555 10680 17685
rect 10640 17525 10645 17555
rect 10675 17525 10680 17555
rect 10640 17395 10680 17525
rect 10640 17365 10645 17395
rect 10675 17365 10680 17395
rect 10640 17235 10680 17365
rect 10640 17205 10645 17235
rect 10675 17205 10680 17235
rect 10640 16195 10680 17205
rect 10640 16165 10645 16195
rect 10675 16165 10680 16195
rect 10640 16035 10680 16165
rect 10640 16005 10645 16035
rect 10675 16005 10680 16035
rect 10640 15875 10680 16005
rect 10640 15845 10645 15875
rect 10675 15845 10680 15875
rect 10640 15715 10680 15845
rect 10640 15685 10645 15715
rect 10675 15685 10680 15715
rect 10640 15555 10680 15685
rect 10640 15525 10645 15555
rect 10675 15525 10680 15555
rect 10640 15395 10680 15525
rect 10640 15365 10645 15395
rect 10675 15365 10680 15395
rect 10640 15235 10680 15365
rect 10640 15205 10645 15235
rect 10675 15205 10680 15235
rect 10640 14720 10680 15205
rect 10720 17955 10760 18680
rect 10720 17925 10725 17955
rect 10755 17925 10760 17955
rect 10720 15475 10760 17925
rect 10720 15445 10725 15475
rect 10755 15445 10760 15475
rect 10720 14720 10760 15445
rect 10800 18195 10840 18680
rect 10800 18165 10805 18195
rect 10835 18165 10840 18195
rect 10800 18035 10840 18165
rect 10800 18005 10805 18035
rect 10835 18005 10840 18035
rect 10800 17875 10840 18005
rect 10800 17845 10805 17875
rect 10835 17845 10840 17875
rect 10800 17715 10840 17845
rect 10800 17685 10805 17715
rect 10835 17685 10840 17715
rect 10800 17555 10840 17685
rect 10800 17525 10805 17555
rect 10835 17525 10840 17555
rect 10800 17395 10840 17525
rect 10800 17365 10805 17395
rect 10835 17365 10840 17395
rect 10800 17235 10840 17365
rect 10800 17205 10805 17235
rect 10835 17205 10840 17235
rect 10800 16195 10840 17205
rect 10800 16165 10805 16195
rect 10835 16165 10840 16195
rect 10800 16035 10840 16165
rect 10800 16005 10805 16035
rect 10835 16005 10840 16035
rect 10800 15875 10840 16005
rect 10800 15845 10805 15875
rect 10835 15845 10840 15875
rect 10800 15715 10840 15845
rect 10800 15685 10805 15715
rect 10835 15685 10840 15715
rect 10800 15555 10840 15685
rect 10800 15525 10805 15555
rect 10835 15525 10840 15555
rect 10800 15395 10840 15525
rect 10800 15365 10805 15395
rect 10835 15365 10840 15395
rect 10800 15235 10840 15365
rect 10800 15205 10805 15235
rect 10835 15205 10840 15235
rect 10800 14720 10840 15205
rect 10880 18115 10920 18680
rect 10880 18085 10885 18115
rect 10915 18085 10920 18115
rect 10880 15315 10920 18085
rect 10880 15285 10885 15315
rect 10915 15285 10920 15315
rect 10880 14720 10920 15285
rect 10960 18195 11000 18680
rect 10960 18165 10965 18195
rect 10995 18165 11000 18195
rect 10960 18035 11000 18165
rect 10960 18005 10965 18035
rect 10995 18005 11000 18035
rect 10960 17875 11000 18005
rect 10960 17845 10965 17875
rect 10995 17845 11000 17875
rect 10960 17715 11000 17845
rect 10960 17685 10965 17715
rect 10995 17685 11000 17715
rect 10960 17555 11000 17685
rect 10960 17525 10965 17555
rect 10995 17525 11000 17555
rect 10960 17395 11000 17525
rect 10960 17365 10965 17395
rect 10995 17365 11000 17395
rect 10960 17235 11000 17365
rect 10960 17205 10965 17235
rect 10995 17205 11000 17235
rect 10960 16195 11000 17205
rect 10960 16165 10965 16195
rect 10995 16165 11000 16195
rect 10960 16035 11000 16165
rect 10960 16005 10965 16035
rect 10995 16005 11000 16035
rect 10960 15875 11000 16005
rect 10960 15845 10965 15875
rect 10995 15845 11000 15875
rect 10960 15715 11000 15845
rect 10960 15685 10965 15715
rect 10995 15685 11000 15715
rect 10960 15555 11000 15685
rect 10960 15525 10965 15555
rect 10995 15525 11000 15555
rect 10960 15395 11000 15525
rect 10960 15365 10965 15395
rect 10995 15365 11000 15395
rect 10960 15235 11000 15365
rect 10960 15205 10965 15235
rect 10995 15205 11000 15235
rect 10960 14720 11000 15205
rect 11040 18435 11080 18680
rect 11040 18405 11045 18435
rect 11075 18405 11080 18435
rect 11040 18275 11080 18405
rect 11040 18245 11045 18275
rect 11075 18245 11080 18275
rect 11040 15155 11080 18245
rect 11040 15125 11045 15155
rect 11075 15125 11080 15155
rect 11040 14995 11080 15125
rect 11040 14965 11045 14995
rect 11075 14965 11080 14995
rect 11040 14720 11080 14965
rect 11120 18355 11160 18680
rect 11120 18325 11125 18355
rect 11155 18325 11160 18355
rect 11120 15075 11160 18325
rect 11120 15045 11125 15075
rect 11155 15045 11160 15075
rect 11120 14720 11160 15045
rect 11200 18435 11240 18680
rect 11200 18405 11205 18435
rect 11235 18405 11240 18435
rect 11200 18275 11240 18405
rect 11200 18245 11205 18275
rect 11235 18245 11240 18275
rect 11200 15155 11240 18245
rect 11200 15125 11205 15155
rect 11235 15125 11240 15155
rect 11200 14995 11240 15125
rect 11200 14965 11205 14995
rect 11235 14965 11240 14995
rect 11200 14720 11240 14965
rect 11280 18675 11320 18680
rect 11280 18645 11285 18675
rect 11315 18645 11320 18675
rect 11280 18515 11320 18645
rect 11280 18485 11285 18515
rect 11315 18485 11320 18515
rect 11280 14915 11320 18485
rect 11280 14885 11285 14915
rect 11315 14885 11320 14915
rect 11280 14755 11320 14885
rect 11280 14725 11285 14755
rect 11315 14725 11320 14755
rect 11280 14720 11320 14725
rect 11360 18595 11400 18680
rect 11360 18565 11365 18595
rect 11395 18565 11400 18595
rect 11360 14835 11400 18565
rect 11360 14805 11365 14835
rect 11395 14805 11400 14835
rect 11360 14720 11400 14805
rect 11440 18675 11480 18680
rect 11440 18645 11445 18675
rect 11475 18645 11480 18675
rect 11440 18515 11480 18645
rect 11440 18485 11445 18515
rect 11475 18485 11480 18515
rect 11440 14915 11480 18485
rect 11560 18675 11600 18680
rect 11560 18645 11565 18675
rect 11595 18645 11600 18675
rect 11560 18515 11600 18645
rect 11560 18485 11565 18515
rect 11595 18485 11600 18515
rect 11560 18480 11600 18485
rect 11640 18675 11680 18680
rect 11640 18645 11645 18675
rect 11675 18645 11680 18675
rect 11640 18515 11680 18645
rect 11640 18485 11645 18515
rect 11675 18485 11680 18515
rect 11640 18480 11680 18485
rect 11720 18675 11760 18680
rect 11720 18645 11725 18675
rect 11755 18645 11760 18675
rect 11720 18515 11760 18645
rect 11720 18485 11725 18515
rect 11755 18485 11760 18515
rect 11720 18480 11760 18485
rect 11800 18675 11840 18680
rect 11800 18645 11805 18675
rect 11835 18645 11840 18675
rect 11800 18515 11840 18645
rect 11800 18485 11805 18515
rect 11835 18485 11840 18515
rect 11800 18480 11840 18485
rect 11880 18675 11920 18680
rect 11880 18645 11885 18675
rect 11915 18645 11920 18675
rect 11880 18515 11920 18645
rect 11880 18485 11885 18515
rect 11915 18485 11920 18515
rect 11880 18480 11920 18485
rect 11960 18675 12000 18680
rect 11960 18645 11965 18675
rect 11995 18645 12000 18675
rect 11960 18515 12000 18645
rect 11960 18485 11965 18515
rect 11995 18485 12000 18515
rect 11960 18480 12000 18485
rect 12040 18675 12080 18680
rect 12040 18645 12045 18675
rect 12075 18645 12080 18675
rect 12040 18515 12080 18645
rect 12040 18485 12045 18515
rect 12075 18485 12080 18515
rect 12040 18480 12080 18485
rect 12120 18675 12160 18680
rect 12120 18645 12125 18675
rect 12155 18645 12160 18675
rect 12120 18515 12160 18645
rect 12120 18485 12125 18515
rect 12155 18485 12160 18515
rect 12120 18480 12160 18485
rect 12200 18675 12240 18680
rect 12200 18645 12205 18675
rect 12235 18645 12240 18675
rect 12200 18515 12240 18645
rect 12200 18485 12205 18515
rect 12235 18485 12240 18515
rect 12200 18480 12240 18485
rect 12280 18675 12320 18680
rect 12280 18645 12285 18675
rect 12315 18645 12320 18675
rect 12280 18515 12320 18645
rect 12280 18485 12285 18515
rect 12315 18485 12320 18515
rect 12280 18480 12320 18485
rect 12360 18675 12400 18680
rect 12360 18645 12365 18675
rect 12395 18645 12400 18675
rect 12360 18515 12400 18645
rect 12360 18485 12365 18515
rect 12395 18485 12400 18515
rect 12360 18480 12400 18485
rect 12440 18675 12480 18680
rect 12440 18645 12445 18675
rect 12475 18645 12480 18675
rect 12440 18515 12480 18645
rect 12440 18485 12445 18515
rect 12475 18485 12480 18515
rect 12440 18480 12480 18485
rect 12520 18675 12560 18680
rect 12520 18645 12525 18675
rect 12555 18645 12560 18675
rect 12520 18515 12560 18645
rect 12520 18485 12525 18515
rect 12555 18485 12560 18515
rect 12520 18480 12560 18485
rect 12600 18675 12640 18680
rect 12600 18645 12605 18675
rect 12635 18645 12640 18675
rect 12600 18515 12640 18645
rect 12600 18485 12605 18515
rect 12635 18485 12640 18515
rect 12600 18480 12640 18485
rect 12680 18675 12720 18680
rect 12680 18645 12685 18675
rect 12715 18645 12720 18675
rect 12680 18515 12720 18645
rect 12680 18485 12685 18515
rect 12715 18485 12720 18515
rect 12680 18480 12720 18485
rect 12760 18675 12800 18680
rect 12760 18645 12765 18675
rect 12795 18645 12800 18675
rect 12760 18515 12800 18645
rect 12760 18485 12765 18515
rect 12795 18485 12800 18515
rect 12760 18480 12800 18485
rect 12840 18675 12880 18680
rect 12840 18645 12845 18675
rect 12875 18645 12880 18675
rect 12840 18515 12880 18645
rect 12840 18485 12845 18515
rect 12875 18485 12880 18515
rect 12840 18480 12880 18485
rect 12920 18675 12960 18680
rect 12920 18645 12925 18675
rect 12955 18645 12960 18675
rect 12920 18515 12960 18645
rect 12920 18485 12925 18515
rect 12955 18485 12960 18515
rect 12920 18480 12960 18485
rect 13000 18675 13040 18680
rect 13000 18645 13005 18675
rect 13035 18645 13040 18675
rect 13000 18515 13040 18645
rect 13000 18485 13005 18515
rect 13035 18485 13040 18515
rect 13000 18480 13040 18485
rect 13080 18675 13120 18680
rect 13080 18645 13085 18675
rect 13115 18645 13120 18675
rect 13080 18515 13120 18645
rect 13080 18485 13085 18515
rect 13115 18485 13120 18515
rect 13080 18480 13120 18485
rect 13160 18675 13200 18680
rect 13160 18645 13165 18675
rect 13195 18645 13200 18675
rect 13160 18515 13200 18645
rect 13160 18485 13165 18515
rect 13195 18485 13200 18515
rect 13160 18480 13200 18485
rect 13240 18675 13280 18680
rect 13240 18645 13245 18675
rect 13275 18645 13280 18675
rect 13240 18515 13280 18645
rect 13240 18485 13245 18515
rect 13275 18485 13280 18515
rect 13240 18480 13280 18485
rect 13320 18675 13360 18680
rect 13320 18645 13325 18675
rect 13355 18645 13360 18675
rect 13320 18515 13360 18645
rect 13320 18485 13325 18515
rect 13355 18485 13360 18515
rect 13320 18480 13360 18485
rect 13400 18675 13440 18680
rect 13400 18645 13405 18675
rect 13435 18645 13440 18675
rect 13400 18515 13440 18645
rect 13400 18485 13405 18515
rect 13435 18485 13440 18515
rect 13400 18480 13440 18485
rect 13480 18675 13520 18680
rect 13480 18645 13485 18675
rect 13515 18645 13520 18675
rect 13480 18515 13520 18645
rect 13480 18485 13485 18515
rect 13515 18485 13520 18515
rect 13480 18480 13520 18485
rect 13560 18675 13600 18680
rect 13560 18645 13565 18675
rect 13595 18645 13600 18675
rect 13560 18515 13600 18645
rect 13560 18485 13565 18515
rect 13595 18485 13600 18515
rect 13560 18480 13600 18485
rect 13640 18675 13680 18680
rect 13640 18645 13645 18675
rect 13675 18645 13680 18675
rect 13640 18515 13680 18645
rect 13640 18485 13645 18515
rect 13675 18485 13680 18515
rect 13640 18480 13680 18485
rect 13720 18675 13760 18680
rect 13720 18645 13725 18675
rect 13755 18645 13760 18675
rect 13720 18515 13760 18645
rect 13720 18485 13725 18515
rect 13755 18485 13760 18515
rect 13720 18480 13760 18485
rect 13800 18675 13840 18680
rect 13800 18645 13805 18675
rect 13835 18645 13840 18675
rect 13800 18515 13840 18645
rect 13800 18485 13805 18515
rect 13835 18485 13840 18515
rect 13800 18480 13840 18485
rect 13880 18675 13920 18680
rect 13880 18645 13885 18675
rect 13915 18645 13920 18675
rect 13880 18515 13920 18645
rect 13880 18485 13885 18515
rect 13915 18485 13920 18515
rect 13880 18480 13920 18485
rect 13960 18675 14000 18680
rect 13960 18645 13965 18675
rect 13995 18645 14000 18675
rect 13960 18515 14000 18645
rect 13960 18485 13965 18515
rect 13995 18485 14000 18515
rect 13960 18480 14000 18485
rect 14040 18675 14080 18680
rect 14040 18645 14045 18675
rect 14075 18645 14080 18675
rect 14040 18515 14080 18645
rect 14040 18485 14045 18515
rect 14075 18485 14080 18515
rect 14040 18480 14080 18485
rect 14120 18675 14160 18680
rect 14120 18645 14125 18675
rect 14155 18645 14160 18675
rect 14120 18515 14160 18645
rect 14120 18485 14125 18515
rect 14155 18485 14160 18515
rect 14120 18480 14160 18485
rect 14200 18675 14240 18680
rect 14200 18645 14205 18675
rect 14235 18645 14240 18675
rect 14200 18515 14240 18645
rect 14200 18485 14205 18515
rect 14235 18485 14240 18515
rect 14200 18480 14240 18485
rect 14280 18675 14320 18680
rect 14280 18645 14285 18675
rect 14315 18645 14320 18675
rect 14280 18515 14320 18645
rect 14280 18485 14285 18515
rect 14315 18485 14320 18515
rect 14280 18480 14320 18485
rect 14360 18675 14400 18680
rect 14360 18645 14365 18675
rect 14395 18645 14400 18675
rect 14360 18515 14400 18645
rect 14360 18485 14365 18515
rect 14395 18485 14400 18515
rect 14360 18480 14400 18485
rect 14440 18675 14480 18680
rect 14440 18645 14445 18675
rect 14475 18645 14480 18675
rect 14440 18515 14480 18645
rect 14440 18485 14445 18515
rect 14475 18485 14480 18515
rect 14440 18480 14480 18485
rect 14520 18675 14560 18680
rect 14520 18645 14525 18675
rect 14555 18645 14560 18675
rect 14520 18515 14560 18645
rect 14520 18485 14525 18515
rect 14555 18485 14560 18515
rect 14520 18480 14560 18485
rect 14600 18675 14640 18680
rect 14600 18645 14605 18675
rect 14635 18645 14640 18675
rect 14600 18515 14640 18645
rect 14600 18485 14605 18515
rect 14635 18485 14640 18515
rect 14600 18480 14640 18485
rect 14680 18675 14720 18680
rect 14680 18645 14685 18675
rect 14715 18645 14720 18675
rect 14680 18515 14720 18645
rect 14680 18485 14685 18515
rect 14715 18485 14720 18515
rect 14680 18480 14720 18485
rect 11560 18435 11600 18440
rect 11560 18405 11565 18435
rect 11595 18405 11600 18435
rect 11560 18275 11600 18405
rect 11560 18245 11565 18275
rect 11595 18245 11600 18275
rect 11560 18240 11600 18245
rect 11640 18435 11680 18440
rect 11640 18405 11645 18435
rect 11675 18405 11680 18435
rect 11640 18275 11680 18405
rect 11640 18245 11645 18275
rect 11675 18245 11680 18275
rect 11640 18240 11680 18245
rect 11720 18435 11760 18440
rect 11720 18405 11725 18435
rect 11755 18405 11760 18435
rect 11720 18275 11760 18405
rect 11720 18245 11725 18275
rect 11755 18245 11760 18275
rect 11720 18240 11760 18245
rect 11800 18435 11840 18440
rect 11800 18405 11805 18435
rect 11835 18405 11840 18435
rect 11800 18275 11840 18405
rect 11800 18245 11805 18275
rect 11835 18245 11840 18275
rect 11800 18240 11840 18245
rect 11880 18435 11920 18440
rect 11880 18405 11885 18435
rect 11915 18405 11920 18435
rect 11880 18275 11920 18405
rect 11880 18245 11885 18275
rect 11915 18245 11920 18275
rect 11880 18240 11920 18245
rect 11960 18435 12000 18440
rect 11960 18405 11965 18435
rect 11995 18405 12000 18435
rect 11960 18275 12000 18405
rect 11960 18245 11965 18275
rect 11995 18245 12000 18275
rect 11960 18240 12000 18245
rect 12040 18435 12080 18440
rect 12040 18405 12045 18435
rect 12075 18405 12080 18435
rect 12040 18275 12080 18405
rect 12040 18245 12045 18275
rect 12075 18245 12080 18275
rect 12040 18240 12080 18245
rect 12120 18435 12160 18440
rect 12120 18405 12125 18435
rect 12155 18405 12160 18435
rect 12120 18275 12160 18405
rect 12120 18245 12125 18275
rect 12155 18245 12160 18275
rect 12120 18240 12160 18245
rect 12200 18435 12240 18440
rect 12200 18405 12205 18435
rect 12235 18405 12240 18435
rect 12200 18275 12240 18405
rect 12200 18245 12205 18275
rect 12235 18245 12240 18275
rect 12200 18240 12240 18245
rect 12280 18435 12320 18440
rect 12280 18405 12285 18435
rect 12315 18405 12320 18435
rect 12280 18275 12320 18405
rect 12280 18245 12285 18275
rect 12315 18245 12320 18275
rect 12280 18240 12320 18245
rect 12360 18435 12400 18440
rect 12360 18405 12365 18435
rect 12395 18405 12400 18435
rect 12360 18275 12400 18405
rect 12360 18245 12365 18275
rect 12395 18245 12400 18275
rect 12360 18240 12400 18245
rect 12440 18435 12480 18440
rect 12440 18405 12445 18435
rect 12475 18405 12480 18435
rect 12440 18275 12480 18405
rect 12440 18245 12445 18275
rect 12475 18245 12480 18275
rect 12440 18240 12480 18245
rect 12520 18435 12560 18440
rect 12520 18405 12525 18435
rect 12555 18405 12560 18435
rect 12520 18275 12560 18405
rect 12520 18245 12525 18275
rect 12555 18245 12560 18275
rect 12520 18240 12560 18245
rect 12600 18435 12640 18440
rect 12600 18405 12605 18435
rect 12635 18405 12640 18435
rect 12600 18275 12640 18405
rect 12600 18245 12605 18275
rect 12635 18245 12640 18275
rect 12600 18240 12640 18245
rect 12680 18435 12720 18440
rect 12680 18405 12685 18435
rect 12715 18405 12720 18435
rect 12680 18275 12720 18405
rect 12680 18245 12685 18275
rect 12715 18245 12720 18275
rect 12680 18240 12720 18245
rect 12760 18435 12800 18440
rect 12760 18405 12765 18435
rect 12795 18405 12800 18435
rect 12760 18275 12800 18405
rect 12760 18245 12765 18275
rect 12795 18245 12800 18275
rect 12760 18240 12800 18245
rect 12840 18435 12880 18440
rect 12840 18405 12845 18435
rect 12875 18405 12880 18435
rect 12840 18275 12880 18405
rect 12840 18245 12845 18275
rect 12875 18245 12880 18275
rect 12840 18240 12880 18245
rect 12920 18435 12960 18440
rect 12920 18405 12925 18435
rect 12955 18405 12960 18435
rect 12920 18275 12960 18405
rect 12920 18245 12925 18275
rect 12955 18245 12960 18275
rect 12920 18240 12960 18245
rect 13000 18435 13040 18440
rect 13000 18405 13005 18435
rect 13035 18405 13040 18435
rect 13000 18275 13040 18405
rect 13000 18245 13005 18275
rect 13035 18245 13040 18275
rect 13000 18240 13040 18245
rect 13080 18435 13120 18440
rect 13080 18405 13085 18435
rect 13115 18405 13120 18435
rect 13080 18275 13120 18405
rect 13080 18245 13085 18275
rect 13115 18245 13120 18275
rect 13080 18240 13120 18245
rect 13160 18435 13200 18440
rect 13160 18405 13165 18435
rect 13195 18405 13200 18435
rect 13160 18275 13200 18405
rect 13160 18245 13165 18275
rect 13195 18245 13200 18275
rect 13160 18240 13200 18245
rect 13240 18435 13280 18440
rect 13240 18405 13245 18435
rect 13275 18405 13280 18435
rect 13240 18275 13280 18405
rect 13240 18245 13245 18275
rect 13275 18245 13280 18275
rect 13240 18240 13280 18245
rect 13320 18435 13360 18440
rect 13320 18405 13325 18435
rect 13355 18405 13360 18435
rect 13320 18275 13360 18405
rect 13320 18245 13325 18275
rect 13355 18245 13360 18275
rect 13320 18240 13360 18245
rect 13400 18435 13440 18440
rect 13400 18405 13405 18435
rect 13435 18405 13440 18435
rect 13400 18275 13440 18405
rect 13400 18245 13405 18275
rect 13435 18245 13440 18275
rect 13400 18240 13440 18245
rect 13480 18435 13520 18440
rect 13480 18405 13485 18435
rect 13515 18405 13520 18435
rect 13480 18275 13520 18405
rect 13480 18245 13485 18275
rect 13515 18245 13520 18275
rect 13480 18240 13520 18245
rect 13560 18435 13600 18440
rect 13560 18405 13565 18435
rect 13595 18405 13600 18435
rect 13560 18275 13600 18405
rect 13560 18245 13565 18275
rect 13595 18245 13600 18275
rect 13560 18240 13600 18245
rect 13640 18435 13680 18440
rect 13640 18405 13645 18435
rect 13675 18405 13680 18435
rect 13640 18275 13680 18405
rect 13640 18245 13645 18275
rect 13675 18245 13680 18275
rect 13640 18240 13680 18245
rect 13720 18435 13760 18440
rect 13720 18405 13725 18435
rect 13755 18405 13760 18435
rect 13720 18275 13760 18405
rect 13720 18245 13725 18275
rect 13755 18245 13760 18275
rect 13720 18240 13760 18245
rect 13800 18435 13840 18440
rect 13800 18405 13805 18435
rect 13835 18405 13840 18435
rect 13800 18275 13840 18405
rect 13800 18245 13805 18275
rect 13835 18245 13840 18275
rect 13800 18240 13840 18245
rect 13880 18435 13920 18440
rect 13880 18405 13885 18435
rect 13915 18405 13920 18435
rect 13880 18275 13920 18405
rect 13880 18245 13885 18275
rect 13915 18245 13920 18275
rect 13880 18240 13920 18245
rect 13960 18435 14000 18440
rect 13960 18405 13965 18435
rect 13995 18405 14000 18435
rect 13960 18275 14000 18405
rect 13960 18245 13965 18275
rect 13995 18245 14000 18275
rect 13960 18240 14000 18245
rect 14040 18435 14080 18440
rect 14040 18405 14045 18435
rect 14075 18405 14080 18435
rect 14040 18275 14080 18405
rect 14040 18245 14045 18275
rect 14075 18245 14080 18275
rect 14040 18240 14080 18245
rect 14120 18435 14160 18440
rect 14120 18405 14125 18435
rect 14155 18405 14160 18435
rect 14120 18275 14160 18405
rect 14120 18245 14125 18275
rect 14155 18245 14160 18275
rect 14120 18240 14160 18245
rect 14200 18435 14240 18440
rect 14200 18405 14205 18435
rect 14235 18405 14240 18435
rect 14200 18275 14240 18405
rect 14200 18245 14205 18275
rect 14235 18245 14240 18275
rect 14200 18240 14240 18245
rect 14280 18435 14320 18440
rect 14280 18405 14285 18435
rect 14315 18405 14320 18435
rect 14280 18275 14320 18405
rect 14280 18245 14285 18275
rect 14315 18245 14320 18275
rect 14280 18240 14320 18245
rect 14360 18435 14400 18440
rect 14360 18405 14365 18435
rect 14395 18405 14400 18435
rect 14360 18275 14400 18405
rect 14360 18245 14365 18275
rect 14395 18245 14400 18275
rect 14360 18240 14400 18245
rect 14440 18435 14480 18440
rect 14440 18405 14445 18435
rect 14475 18405 14480 18435
rect 14440 18275 14480 18405
rect 14440 18245 14445 18275
rect 14475 18245 14480 18275
rect 14440 18240 14480 18245
rect 14520 18435 14560 18440
rect 14520 18405 14525 18435
rect 14555 18405 14560 18435
rect 14520 18275 14560 18405
rect 14520 18245 14525 18275
rect 14555 18245 14560 18275
rect 14520 18240 14560 18245
rect 14600 18435 14640 18440
rect 14600 18405 14605 18435
rect 14635 18405 14640 18435
rect 14600 18275 14640 18405
rect 14600 18245 14605 18275
rect 14635 18245 14640 18275
rect 14600 18240 14640 18245
rect 14680 18435 14720 18440
rect 14680 18405 14685 18435
rect 14715 18405 14720 18435
rect 14680 18275 14720 18405
rect 14680 18245 14685 18275
rect 14715 18245 14720 18275
rect 14680 18240 14720 18245
rect 11560 18195 11600 18200
rect 11560 18165 11565 18195
rect 11595 18165 11600 18195
rect 11560 18035 11600 18165
rect 11560 18005 11565 18035
rect 11595 18005 11600 18035
rect 11560 17875 11600 18005
rect 11560 17845 11565 17875
rect 11595 17845 11600 17875
rect 11560 17715 11600 17845
rect 11560 17685 11565 17715
rect 11595 17685 11600 17715
rect 11560 17555 11600 17685
rect 11560 17525 11565 17555
rect 11595 17525 11600 17555
rect 11560 17395 11600 17525
rect 11560 17365 11565 17395
rect 11595 17365 11600 17395
rect 11560 17235 11600 17365
rect 11560 17205 11565 17235
rect 11595 17205 11600 17235
rect 11560 17200 11600 17205
rect 11640 18195 11680 18200
rect 11640 18165 11645 18195
rect 11675 18165 11680 18195
rect 11640 18035 11680 18165
rect 11640 18005 11645 18035
rect 11675 18005 11680 18035
rect 11640 17875 11680 18005
rect 11640 17845 11645 17875
rect 11675 17845 11680 17875
rect 11640 17715 11680 17845
rect 11640 17685 11645 17715
rect 11675 17685 11680 17715
rect 11640 17555 11680 17685
rect 11640 17525 11645 17555
rect 11675 17525 11680 17555
rect 11640 17395 11680 17525
rect 11640 17365 11645 17395
rect 11675 17365 11680 17395
rect 11640 17235 11680 17365
rect 11640 17205 11645 17235
rect 11675 17205 11680 17235
rect 11640 17200 11680 17205
rect 11720 18195 11760 18200
rect 11720 18165 11725 18195
rect 11755 18165 11760 18195
rect 11720 18035 11760 18165
rect 11720 18005 11725 18035
rect 11755 18005 11760 18035
rect 11720 17875 11760 18005
rect 11720 17845 11725 17875
rect 11755 17845 11760 17875
rect 11720 17715 11760 17845
rect 11720 17685 11725 17715
rect 11755 17685 11760 17715
rect 11720 17555 11760 17685
rect 11720 17525 11725 17555
rect 11755 17525 11760 17555
rect 11720 17395 11760 17525
rect 11720 17365 11725 17395
rect 11755 17365 11760 17395
rect 11720 17235 11760 17365
rect 11720 17205 11725 17235
rect 11755 17205 11760 17235
rect 11720 17200 11760 17205
rect 11800 18195 11840 18200
rect 11800 18165 11805 18195
rect 11835 18165 11840 18195
rect 11800 18035 11840 18165
rect 11800 18005 11805 18035
rect 11835 18005 11840 18035
rect 11800 17875 11840 18005
rect 11800 17845 11805 17875
rect 11835 17845 11840 17875
rect 11800 17715 11840 17845
rect 11800 17685 11805 17715
rect 11835 17685 11840 17715
rect 11800 17555 11840 17685
rect 11800 17525 11805 17555
rect 11835 17525 11840 17555
rect 11800 17395 11840 17525
rect 11800 17365 11805 17395
rect 11835 17365 11840 17395
rect 11800 17235 11840 17365
rect 11800 17205 11805 17235
rect 11835 17205 11840 17235
rect 11800 17200 11840 17205
rect 11880 18195 11920 18200
rect 11880 18165 11885 18195
rect 11915 18165 11920 18195
rect 11880 18035 11920 18165
rect 11880 18005 11885 18035
rect 11915 18005 11920 18035
rect 11880 17875 11920 18005
rect 11880 17845 11885 17875
rect 11915 17845 11920 17875
rect 11880 17715 11920 17845
rect 11880 17685 11885 17715
rect 11915 17685 11920 17715
rect 11880 17555 11920 17685
rect 11880 17525 11885 17555
rect 11915 17525 11920 17555
rect 11880 17395 11920 17525
rect 11880 17365 11885 17395
rect 11915 17365 11920 17395
rect 11880 17235 11920 17365
rect 11880 17205 11885 17235
rect 11915 17205 11920 17235
rect 11880 17200 11920 17205
rect 11960 18195 12000 18200
rect 11960 18165 11965 18195
rect 11995 18165 12000 18195
rect 11960 18035 12000 18165
rect 11960 18005 11965 18035
rect 11995 18005 12000 18035
rect 11960 17875 12000 18005
rect 11960 17845 11965 17875
rect 11995 17845 12000 17875
rect 11960 17715 12000 17845
rect 11960 17685 11965 17715
rect 11995 17685 12000 17715
rect 11960 17555 12000 17685
rect 11960 17525 11965 17555
rect 11995 17525 12000 17555
rect 11960 17395 12000 17525
rect 11960 17365 11965 17395
rect 11995 17365 12000 17395
rect 11960 17235 12000 17365
rect 11960 17205 11965 17235
rect 11995 17205 12000 17235
rect 11960 17200 12000 17205
rect 12040 18195 12080 18200
rect 12040 18165 12045 18195
rect 12075 18165 12080 18195
rect 12040 18035 12080 18165
rect 12040 18005 12045 18035
rect 12075 18005 12080 18035
rect 12040 17875 12080 18005
rect 12040 17845 12045 17875
rect 12075 17845 12080 17875
rect 12040 17715 12080 17845
rect 12040 17685 12045 17715
rect 12075 17685 12080 17715
rect 12040 17555 12080 17685
rect 12040 17525 12045 17555
rect 12075 17525 12080 17555
rect 12040 17395 12080 17525
rect 12040 17365 12045 17395
rect 12075 17365 12080 17395
rect 12040 17235 12080 17365
rect 12040 17205 12045 17235
rect 12075 17205 12080 17235
rect 12040 17200 12080 17205
rect 12120 18195 12160 18200
rect 12120 18165 12125 18195
rect 12155 18165 12160 18195
rect 12120 18035 12160 18165
rect 12120 18005 12125 18035
rect 12155 18005 12160 18035
rect 12120 17875 12160 18005
rect 12120 17845 12125 17875
rect 12155 17845 12160 17875
rect 12120 17715 12160 17845
rect 12120 17685 12125 17715
rect 12155 17685 12160 17715
rect 12120 17555 12160 17685
rect 12120 17525 12125 17555
rect 12155 17525 12160 17555
rect 12120 17395 12160 17525
rect 12120 17365 12125 17395
rect 12155 17365 12160 17395
rect 12120 17235 12160 17365
rect 12120 17205 12125 17235
rect 12155 17205 12160 17235
rect 12120 17200 12160 17205
rect 12200 18195 12240 18200
rect 12200 18165 12205 18195
rect 12235 18165 12240 18195
rect 12200 18035 12240 18165
rect 12200 18005 12205 18035
rect 12235 18005 12240 18035
rect 12200 17875 12240 18005
rect 12200 17845 12205 17875
rect 12235 17845 12240 17875
rect 12200 17715 12240 17845
rect 12200 17685 12205 17715
rect 12235 17685 12240 17715
rect 12200 17555 12240 17685
rect 12200 17525 12205 17555
rect 12235 17525 12240 17555
rect 12200 17395 12240 17525
rect 12200 17365 12205 17395
rect 12235 17365 12240 17395
rect 12200 17235 12240 17365
rect 12200 17205 12205 17235
rect 12235 17205 12240 17235
rect 12200 17200 12240 17205
rect 12280 18195 12320 18200
rect 12280 18165 12285 18195
rect 12315 18165 12320 18195
rect 12280 18035 12320 18165
rect 12280 18005 12285 18035
rect 12315 18005 12320 18035
rect 12280 17875 12320 18005
rect 12280 17845 12285 17875
rect 12315 17845 12320 17875
rect 12280 17715 12320 17845
rect 12280 17685 12285 17715
rect 12315 17685 12320 17715
rect 12280 17555 12320 17685
rect 12280 17525 12285 17555
rect 12315 17525 12320 17555
rect 12280 17395 12320 17525
rect 12280 17365 12285 17395
rect 12315 17365 12320 17395
rect 12280 17235 12320 17365
rect 12280 17205 12285 17235
rect 12315 17205 12320 17235
rect 12280 17200 12320 17205
rect 12360 18195 12400 18200
rect 12360 18165 12365 18195
rect 12395 18165 12400 18195
rect 12360 18035 12400 18165
rect 12360 18005 12365 18035
rect 12395 18005 12400 18035
rect 12360 17875 12400 18005
rect 12360 17845 12365 17875
rect 12395 17845 12400 17875
rect 12360 17715 12400 17845
rect 12360 17685 12365 17715
rect 12395 17685 12400 17715
rect 12360 17555 12400 17685
rect 12360 17525 12365 17555
rect 12395 17525 12400 17555
rect 12360 17395 12400 17525
rect 12360 17365 12365 17395
rect 12395 17365 12400 17395
rect 12360 17235 12400 17365
rect 12360 17205 12365 17235
rect 12395 17205 12400 17235
rect 12360 17200 12400 17205
rect 12440 18195 12480 18200
rect 12440 18165 12445 18195
rect 12475 18165 12480 18195
rect 12440 18035 12480 18165
rect 12440 18005 12445 18035
rect 12475 18005 12480 18035
rect 12440 17875 12480 18005
rect 12440 17845 12445 17875
rect 12475 17845 12480 17875
rect 12440 17715 12480 17845
rect 12440 17685 12445 17715
rect 12475 17685 12480 17715
rect 12440 17555 12480 17685
rect 12440 17525 12445 17555
rect 12475 17525 12480 17555
rect 12440 17395 12480 17525
rect 12440 17365 12445 17395
rect 12475 17365 12480 17395
rect 12440 17235 12480 17365
rect 12440 17205 12445 17235
rect 12475 17205 12480 17235
rect 12440 17200 12480 17205
rect 12520 18195 12560 18200
rect 12520 18165 12525 18195
rect 12555 18165 12560 18195
rect 12520 18035 12560 18165
rect 12520 18005 12525 18035
rect 12555 18005 12560 18035
rect 12520 17875 12560 18005
rect 12520 17845 12525 17875
rect 12555 17845 12560 17875
rect 12520 17715 12560 17845
rect 12520 17685 12525 17715
rect 12555 17685 12560 17715
rect 12520 17555 12560 17685
rect 12520 17525 12525 17555
rect 12555 17525 12560 17555
rect 12520 17395 12560 17525
rect 12520 17365 12525 17395
rect 12555 17365 12560 17395
rect 12520 17235 12560 17365
rect 12520 17205 12525 17235
rect 12555 17205 12560 17235
rect 12520 17200 12560 17205
rect 12600 18195 12640 18200
rect 12600 18165 12605 18195
rect 12635 18165 12640 18195
rect 12600 18035 12640 18165
rect 12600 18005 12605 18035
rect 12635 18005 12640 18035
rect 12600 17875 12640 18005
rect 12600 17845 12605 17875
rect 12635 17845 12640 17875
rect 12600 17715 12640 17845
rect 12600 17685 12605 17715
rect 12635 17685 12640 17715
rect 12600 17555 12640 17685
rect 12600 17525 12605 17555
rect 12635 17525 12640 17555
rect 12600 17395 12640 17525
rect 12600 17365 12605 17395
rect 12635 17365 12640 17395
rect 12600 17235 12640 17365
rect 12600 17205 12605 17235
rect 12635 17205 12640 17235
rect 12600 17200 12640 17205
rect 12680 18195 12720 18200
rect 12680 18165 12685 18195
rect 12715 18165 12720 18195
rect 12680 18035 12720 18165
rect 12680 18005 12685 18035
rect 12715 18005 12720 18035
rect 12680 17875 12720 18005
rect 12680 17845 12685 17875
rect 12715 17845 12720 17875
rect 12680 17715 12720 17845
rect 12680 17685 12685 17715
rect 12715 17685 12720 17715
rect 12680 17555 12720 17685
rect 12680 17525 12685 17555
rect 12715 17525 12720 17555
rect 12680 17395 12720 17525
rect 12680 17365 12685 17395
rect 12715 17365 12720 17395
rect 12680 17235 12720 17365
rect 12680 17205 12685 17235
rect 12715 17205 12720 17235
rect 12680 17200 12720 17205
rect 12760 18195 12800 18200
rect 12760 18165 12765 18195
rect 12795 18165 12800 18195
rect 12760 18035 12800 18165
rect 12760 18005 12765 18035
rect 12795 18005 12800 18035
rect 12760 17875 12800 18005
rect 12760 17845 12765 17875
rect 12795 17845 12800 17875
rect 12760 17715 12800 17845
rect 12760 17685 12765 17715
rect 12795 17685 12800 17715
rect 12760 17555 12800 17685
rect 12760 17525 12765 17555
rect 12795 17525 12800 17555
rect 12760 17395 12800 17525
rect 12760 17365 12765 17395
rect 12795 17365 12800 17395
rect 12760 17235 12800 17365
rect 12760 17205 12765 17235
rect 12795 17205 12800 17235
rect 12760 17200 12800 17205
rect 12840 18195 12880 18200
rect 12840 18165 12845 18195
rect 12875 18165 12880 18195
rect 12840 18035 12880 18165
rect 12840 18005 12845 18035
rect 12875 18005 12880 18035
rect 12840 17875 12880 18005
rect 12840 17845 12845 17875
rect 12875 17845 12880 17875
rect 12840 17715 12880 17845
rect 12840 17685 12845 17715
rect 12875 17685 12880 17715
rect 12840 17555 12880 17685
rect 12840 17525 12845 17555
rect 12875 17525 12880 17555
rect 12840 17395 12880 17525
rect 12840 17365 12845 17395
rect 12875 17365 12880 17395
rect 12840 17235 12880 17365
rect 12840 17205 12845 17235
rect 12875 17205 12880 17235
rect 12840 17200 12880 17205
rect 12920 18195 12960 18200
rect 12920 18165 12925 18195
rect 12955 18165 12960 18195
rect 12920 18035 12960 18165
rect 12920 18005 12925 18035
rect 12955 18005 12960 18035
rect 12920 17875 12960 18005
rect 12920 17845 12925 17875
rect 12955 17845 12960 17875
rect 12920 17715 12960 17845
rect 12920 17685 12925 17715
rect 12955 17685 12960 17715
rect 12920 17555 12960 17685
rect 12920 17525 12925 17555
rect 12955 17525 12960 17555
rect 12920 17395 12960 17525
rect 12920 17365 12925 17395
rect 12955 17365 12960 17395
rect 12920 17235 12960 17365
rect 12920 17205 12925 17235
rect 12955 17205 12960 17235
rect 12920 17200 12960 17205
rect 13000 18195 13040 18200
rect 13000 18165 13005 18195
rect 13035 18165 13040 18195
rect 13000 18035 13040 18165
rect 13000 18005 13005 18035
rect 13035 18005 13040 18035
rect 13000 17875 13040 18005
rect 13000 17845 13005 17875
rect 13035 17845 13040 17875
rect 13000 17715 13040 17845
rect 13000 17685 13005 17715
rect 13035 17685 13040 17715
rect 13000 17555 13040 17685
rect 13000 17525 13005 17555
rect 13035 17525 13040 17555
rect 13000 17395 13040 17525
rect 13000 17365 13005 17395
rect 13035 17365 13040 17395
rect 13000 17235 13040 17365
rect 13000 17205 13005 17235
rect 13035 17205 13040 17235
rect 13000 17200 13040 17205
rect 13080 18195 13120 18200
rect 13080 18165 13085 18195
rect 13115 18165 13120 18195
rect 13080 18035 13120 18165
rect 13080 18005 13085 18035
rect 13115 18005 13120 18035
rect 13080 17875 13120 18005
rect 13080 17845 13085 17875
rect 13115 17845 13120 17875
rect 13080 17715 13120 17845
rect 13080 17685 13085 17715
rect 13115 17685 13120 17715
rect 13080 17555 13120 17685
rect 13080 17525 13085 17555
rect 13115 17525 13120 17555
rect 13080 17395 13120 17525
rect 13080 17365 13085 17395
rect 13115 17365 13120 17395
rect 13080 17235 13120 17365
rect 13080 17205 13085 17235
rect 13115 17205 13120 17235
rect 13080 17200 13120 17205
rect 13160 18195 13200 18200
rect 13160 18165 13165 18195
rect 13195 18165 13200 18195
rect 13160 18035 13200 18165
rect 13160 18005 13165 18035
rect 13195 18005 13200 18035
rect 13160 17875 13200 18005
rect 13160 17845 13165 17875
rect 13195 17845 13200 17875
rect 13160 17715 13200 17845
rect 13160 17685 13165 17715
rect 13195 17685 13200 17715
rect 13160 17555 13200 17685
rect 13160 17525 13165 17555
rect 13195 17525 13200 17555
rect 13160 17395 13200 17525
rect 13160 17365 13165 17395
rect 13195 17365 13200 17395
rect 13160 17235 13200 17365
rect 13160 17205 13165 17235
rect 13195 17205 13200 17235
rect 13160 17200 13200 17205
rect 13240 18195 13280 18200
rect 13240 18165 13245 18195
rect 13275 18165 13280 18195
rect 13240 18035 13280 18165
rect 13240 18005 13245 18035
rect 13275 18005 13280 18035
rect 13240 17875 13280 18005
rect 13240 17845 13245 17875
rect 13275 17845 13280 17875
rect 13240 17715 13280 17845
rect 13240 17685 13245 17715
rect 13275 17685 13280 17715
rect 13240 17555 13280 17685
rect 13240 17525 13245 17555
rect 13275 17525 13280 17555
rect 13240 17395 13280 17525
rect 13240 17365 13245 17395
rect 13275 17365 13280 17395
rect 13240 17235 13280 17365
rect 13240 17205 13245 17235
rect 13275 17205 13280 17235
rect 13240 17200 13280 17205
rect 13320 18195 13360 18200
rect 13320 18165 13325 18195
rect 13355 18165 13360 18195
rect 13320 18035 13360 18165
rect 13320 18005 13325 18035
rect 13355 18005 13360 18035
rect 13320 17875 13360 18005
rect 13320 17845 13325 17875
rect 13355 17845 13360 17875
rect 13320 17715 13360 17845
rect 13320 17685 13325 17715
rect 13355 17685 13360 17715
rect 13320 17555 13360 17685
rect 13320 17525 13325 17555
rect 13355 17525 13360 17555
rect 13320 17395 13360 17525
rect 13320 17365 13325 17395
rect 13355 17365 13360 17395
rect 13320 17235 13360 17365
rect 13320 17205 13325 17235
rect 13355 17205 13360 17235
rect 13320 17200 13360 17205
rect 13400 18195 13440 18200
rect 13400 18165 13405 18195
rect 13435 18165 13440 18195
rect 13400 18035 13440 18165
rect 13400 18005 13405 18035
rect 13435 18005 13440 18035
rect 13400 17875 13440 18005
rect 13400 17845 13405 17875
rect 13435 17845 13440 17875
rect 13400 17715 13440 17845
rect 13400 17685 13405 17715
rect 13435 17685 13440 17715
rect 13400 17555 13440 17685
rect 13400 17525 13405 17555
rect 13435 17525 13440 17555
rect 13400 17395 13440 17525
rect 13400 17365 13405 17395
rect 13435 17365 13440 17395
rect 13400 17235 13440 17365
rect 13400 17205 13405 17235
rect 13435 17205 13440 17235
rect 13400 17200 13440 17205
rect 13480 18195 13520 18200
rect 13480 18165 13485 18195
rect 13515 18165 13520 18195
rect 13480 18035 13520 18165
rect 13480 18005 13485 18035
rect 13515 18005 13520 18035
rect 13480 17875 13520 18005
rect 13480 17845 13485 17875
rect 13515 17845 13520 17875
rect 13480 17715 13520 17845
rect 13480 17685 13485 17715
rect 13515 17685 13520 17715
rect 13480 17555 13520 17685
rect 13480 17525 13485 17555
rect 13515 17525 13520 17555
rect 13480 17395 13520 17525
rect 13480 17365 13485 17395
rect 13515 17365 13520 17395
rect 13480 17235 13520 17365
rect 13480 17205 13485 17235
rect 13515 17205 13520 17235
rect 13480 17200 13520 17205
rect 13560 18195 13600 18200
rect 13560 18165 13565 18195
rect 13595 18165 13600 18195
rect 13560 18035 13600 18165
rect 13560 18005 13565 18035
rect 13595 18005 13600 18035
rect 13560 17875 13600 18005
rect 13560 17845 13565 17875
rect 13595 17845 13600 17875
rect 13560 17715 13600 17845
rect 13560 17685 13565 17715
rect 13595 17685 13600 17715
rect 13560 17555 13600 17685
rect 13560 17525 13565 17555
rect 13595 17525 13600 17555
rect 13560 17395 13600 17525
rect 13560 17365 13565 17395
rect 13595 17365 13600 17395
rect 13560 17235 13600 17365
rect 13560 17205 13565 17235
rect 13595 17205 13600 17235
rect 13560 17200 13600 17205
rect 13640 18195 13680 18200
rect 13640 18165 13645 18195
rect 13675 18165 13680 18195
rect 13640 18035 13680 18165
rect 13640 18005 13645 18035
rect 13675 18005 13680 18035
rect 13640 17875 13680 18005
rect 13640 17845 13645 17875
rect 13675 17845 13680 17875
rect 13640 17715 13680 17845
rect 13640 17685 13645 17715
rect 13675 17685 13680 17715
rect 13640 17555 13680 17685
rect 13640 17525 13645 17555
rect 13675 17525 13680 17555
rect 13640 17395 13680 17525
rect 13640 17365 13645 17395
rect 13675 17365 13680 17395
rect 13640 17235 13680 17365
rect 13640 17205 13645 17235
rect 13675 17205 13680 17235
rect 13640 17200 13680 17205
rect 13720 18195 13760 18200
rect 13720 18165 13725 18195
rect 13755 18165 13760 18195
rect 13720 18035 13760 18165
rect 13720 18005 13725 18035
rect 13755 18005 13760 18035
rect 13720 17875 13760 18005
rect 13720 17845 13725 17875
rect 13755 17845 13760 17875
rect 13720 17715 13760 17845
rect 13720 17685 13725 17715
rect 13755 17685 13760 17715
rect 13720 17555 13760 17685
rect 13720 17525 13725 17555
rect 13755 17525 13760 17555
rect 13720 17395 13760 17525
rect 13720 17365 13725 17395
rect 13755 17365 13760 17395
rect 13720 17235 13760 17365
rect 13720 17205 13725 17235
rect 13755 17205 13760 17235
rect 13720 17200 13760 17205
rect 13800 18195 13840 18200
rect 13800 18165 13805 18195
rect 13835 18165 13840 18195
rect 13800 18035 13840 18165
rect 13800 18005 13805 18035
rect 13835 18005 13840 18035
rect 13800 17875 13840 18005
rect 13800 17845 13805 17875
rect 13835 17845 13840 17875
rect 13800 17715 13840 17845
rect 13800 17685 13805 17715
rect 13835 17685 13840 17715
rect 13800 17555 13840 17685
rect 13800 17525 13805 17555
rect 13835 17525 13840 17555
rect 13800 17395 13840 17525
rect 13800 17365 13805 17395
rect 13835 17365 13840 17395
rect 13800 17235 13840 17365
rect 13800 17205 13805 17235
rect 13835 17205 13840 17235
rect 13800 17200 13840 17205
rect 13880 18195 13920 18200
rect 13880 18165 13885 18195
rect 13915 18165 13920 18195
rect 13880 18035 13920 18165
rect 13880 18005 13885 18035
rect 13915 18005 13920 18035
rect 13880 17875 13920 18005
rect 13880 17845 13885 17875
rect 13915 17845 13920 17875
rect 13880 17715 13920 17845
rect 13880 17685 13885 17715
rect 13915 17685 13920 17715
rect 13880 17555 13920 17685
rect 13880 17525 13885 17555
rect 13915 17525 13920 17555
rect 13880 17395 13920 17525
rect 13880 17365 13885 17395
rect 13915 17365 13920 17395
rect 13880 17235 13920 17365
rect 13880 17205 13885 17235
rect 13915 17205 13920 17235
rect 13880 17200 13920 17205
rect 13960 18195 14000 18200
rect 13960 18165 13965 18195
rect 13995 18165 14000 18195
rect 13960 18035 14000 18165
rect 13960 18005 13965 18035
rect 13995 18005 14000 18035
rect 13960 17875 14000 18005
rect 13960 17845 13965 17875
rect 13995 17845 14000 17875
rect 13960 17715 14000 17845
rect 13960 17685 13965 17715
rect 13995 17685 14000 17715
rect 13960 17555 14000 17685
rect 13960 17525 13965 17555
rect 13995 17525 14000 17555
rect 13960 17395 14000 17525
rect 13960 17365 13965 17395
rect 13995 17365 14000 17395
rect 13960 17235 14000 17365
rect 13960 17205 13965 17235
rect 13995 17205 14000 17235
rect 13960 17200 14000 17205
rect 14040 18195 14080 18200
rect 14040 18165 14045 18195
rect 14075 18165 14080 18195
rect 14040 18035 14080 18165
rect 14040 18005 14045 18035
rect 14075 18005 14080 18035
rect 14040 17875 14080 18005
rect 14040 17845 14045 17875
rect 14075 17845 14080 17875
rect 14040 17715 14080 17845
rect 14040 17685 14045 17715
rect 14075 17685 14080 17715
rect 14040 17555 14080 17685
rect 14040 17525 14045 17555
rect 14075 17525 14080 17555
rect 14040 17395 14080 17525
rect 14040 17365 14045 17395
rect 14075 17365 14080 17395
rect 14040 17235 14080 17365
rect 14040 17205 14045 17235
rect 14075 17205 14080 17235
rect 14040 17200 14080 17205
rect 14120 18195 14160 18200
rect 14120 18165 14125 18195
rect 14155 18165 14160 18195
rect 14120 18035 14160 18165
rect 14120 18005 14125 18035
rect 14155 18005 14160 18035
rect 14120 17875 14160 18005
rect 14120 17845 14125 17875
rect 14155 17845 14160 17875
rect 14120 17715 14160 17845
rect 14120 17685 14125 17715
rect 14155 17685 14160 17715
rect 14120 17555 14160 17685
rect 14120 17525 14125 17555
rect 14155 17525 14160 17555
rect 14120 17395 14160 17525
rect 14120 17365 14125 17395
rect 14155 17365 14160 17395
rect 14120 17235 14160 17365
rect 14120 17205 14125 17235
rect 14155 17205 14160 17235
rect 14120 17200 14160 17205
rect 14200 18195 14240 18200
rect 14200 18165 14205 18195
rect 14235 18165 14240 18195
rect 14200 18035 14240 18165
rect 14200 18005 14205 18035
rect 14235 18005 14240 18035
rect 14200 17875 14240 18005
rect 14200 17845 14205 17875
rect 14235 17845 14240 17875
rect 14200 17715 14240 17845
rect 14200 17685 14205 17715
rect 14235 17685 14240 17715
rect 14200 17555 14240 17685
rect 14200 17525 14205 17555
rect 14235 17525 14240 17555
rect 14200 17395 14240 17525
rect 14200 17365 14205 17395
rect 14235 17365 14240 17395
rect 14200 17235 14240 17365
rect 14200 17205 14205 17235
rect 14235 17205 14240 17235
rect 14200 17200 14240 17205
rect 14280 18195 14320 18200
rect 14280 18165 14285 18195
rect 14315 18165 14320 18195
rect 14280 18035 14320 18165
rect 14280 18005 14285 18035
rect 14315 18005 14320 18035
rect 14280 17875 14320 18005
rect 14280 17845 14285 17875
rect 14315 17845 14320 17875
rect 14280 17715 14320 17845
rect 14280 17685 14285 17715
rect 14315 17685 14320 17715
rect 14280 17555 14320 17685
rect 14280 17525 14285 17555
rect 14315 17525 14320 17555
rect 14280 17395 14320 17525
rect 14280 17365 14285 17395
rect 14315 17365 14320 17395
rect 14280 17235 14320 17365
rect 14280 17205 14285 17235
rect 14315 17205 14320 17235
rect 14280 17200 14320 17205
rect 14360 18195 14400 18200
rect 14360 18165 14365 18195
rect 14395 18165 14400 18195
rect 14360 18035 14400 18165
rect 14360 18005 14365 18035
rect 14395 18005 14400 18035
rect 14360 17875 14400 18005
rect 14360 17845 14365 17875
rect 14395 17845 14400 17875
rect 14360 17715 14400 17845
rect 14360 17685 14365 17715
rect 14395 17685 14400 17715
rect 14360 17555 14400 17685
rect 14360 17525 14365 17555
rect 14395 17525 14400 17555
rect 14360 17395 14400 17525
rect 14360 17365 14365 17395
rect 14395 17365 14400 17395
rect 14360 17235 14400 17365
rect 14360 17205 14365 17235
rect 14395 17205 14400 17235
rect 14360 17200 14400 17205
rect 14440 18195 14480 18200
rect 14440 18165 14445 18195
rect 14475 18165 14480 18195
rect 14440 18035 14480 18165
rect 14440 18005 14445 18035
rect 14475 18005 14480 18035
rect 14440 17875 14480 18005
rect 14440 17845 14445 17875
rect 14475 17845 14480 17875
rect 14440 17715 14480 17845
rect 14440 17685 14445 17715
rect 14475 17685 14480 17715
rect 14440 17555 14480 17685
rect 14440 17525 14445 17555
rect 14475 17525 14480 17555
rect 14440 17395 14480 17525
rect 14440 17365 14445 17395
rect 14475 17365 14480 17395
rect 14440 17235 14480 17365
rect 14440 17205 14445 17235
rect 14475 17205 14480 17235
rect 14440 17200 14480 17205
rect 14520 18195 14560 18200
rect 14520 18165 14525 18195
rect 14555 18165 14560 18195
rect 14520 18035 14560 18165
rect 14520 18005 14525 18035
rect 14555 18005 14560 18035
rect 14520 17875 14560 18005
rect 14520 17845 14525 17875
rect 14555 17845 14560 17875
rect 14520 17715 14560 17845
rect 14520 17685 14525 17715
rect 14555 17685 14560 17715
rect 14520 17555 14560 17685
rect 14520 17525 14525 17555
rect 14555 17525 14560 17555
rect 14520 17395 14560 17525
rect 14520 17365 14525 17395
rect 14555 17365 14560 17395
rect 14520 17235 14560 17365
rect 14520 17205 14525 17235
rect 14555 17205 14560 17235
rect 14520 17200 14560 17205
rect 14600 18195 14640 18200
rect 14600 18165 14605 18195
rect 14635 18165 14640 18195
rect 14600 18035 14640 18165
rect 14600 18005 14605 18035
rect 14635 18005 14640 18035
rect 14600 17875 14640 18005
rect 14600 17845 14605 17875
rect 14635 17845 14640 17875
rect 14600 17715 14640 17845
rect 14600 17685 14605 17715
rect 14635 17685 14640 17715
rect 14600 17555 14640 17685
rect 14600 17525 14605 17555
rect 14635 17525 14640 17555
rect 14600 17395 14640 17525
rect 14600 17365 14605 17395
rect 14635 17365 14640 17395
rect 14600 17235 14640 17365
rect 14600 17205 14605 17235
rect 14635 17205 14640 17235
rect 14600 17200 14640 17205
rect 14680 18195 14720 18200
rect 14680 18165 14685 18195
rect 14715 18165 14720 18195
rect 14680 18035 14720 18165
rect 14680 18005 14685 18035
rect 14715 18005 14720 18035
rect 14680 17875 14720 18005
rect 14680 17845 14685 17875
rect 14715 17845 14720 17875
rect 14680 17715 14720 17845
rect 14680 17685 14685 17715
rect 14715 17685 14720 17715
rect 14680 17555 14720 17685
rect 14680 17525 14685 17555
rect 14715 17525 14720 17555
rect 14680 17395 14720 17525
rect 14680 17365 14685 17395
rect 14715 17365 14720 17395
rect 14680 17235 14720 17365
rect 14680 17205 14685 17235
rect 14715 17205 14720 17235
rect 14680 17200 14720 17205
rect 11560 17155 11600 17160
rect 11560 17125 11565 17155
rect 11595 17125 11600 17155
rect 11560 16995 11600 17125
rect 11560 16965 11565 16995
rect 11595 16965 11600 16995
rect 11560 16960 11600 16965
rect 11640 17155 11680 17160
rect 11640 17125 11645 17155
rect 11675 17125 11680 17155
rect 11640 16995 11680 17125
rect 11640 16965 11645 16995
rect 11675 16965 11680 16995
rect 11640 16960 11680 16965
rect 11720 17155 11760 17160
rect 11720 17125 11725 17155
rect 11755 17125 11760 17155
rect 11720 16995 11760 17125
rect 11720 16965 11725 16995
rect 11755 16965 11760 16995
rect 11720 16960 11760 16965
rect 11800 17155 11840 17160
rect 11800 17125 11805 17155
rect 11835 17125 11840 17155
rect 11800 16995 11840 17125
rect 11800 16965 11805 16995
rect 11835 16965 11840 16995
rect 11800 16960 11840 16965
rect 11880 17155 11920 17160
rect 11880 17125 11885 17155
rect 11915 17125 11920 17155
rect 11880 16995 11920 17125
rect 11880 16965 11885 16995
rect 11915 16965 11920 16995
rect 11880 16960 11920 16965
rect 11960 17155 12000 17160
rect 11960 17125 11965 17155
rect 11995 17125 12000 17155
rect 11960 16995 12000 17125
rect 11960 16965 11965 16995
rect 11995 16965 12000 16995
rect 11960 16960 12000 16965
rect 12040 17155 12080 17160
rect 12040 17125 12045 17155
rect 12075 17125 12080 17155
rect 12040 16995 12080 17125
rect 12040 16965 12045 16995
rect 12075 16965 12080 16995
rect 12040 16960 12080 16965
rect 12120 17155 12160 17160
rect 12120 17125 12125 17155
rect 12155 17125 12160 17155
rect 12120 16995 12160 17125
rect 12120 16965 12125 16995
rect 12155 16965 12160 16995
rect 12120 16960 12160 16965
rect 12200 17155 12240 17160
rect 12200 17125 12205 17155
rect 12235 17125 12240 17155
rect 12200 16995 12240 17125
rect 12200 16965 12205 16995
rect 12235 16965 12240 16995
rect 12200 16960 12240 16965
rect 12280 17155 12320 17160
rect 12280 17125 12285 17155
rect 12315 17125 12320 17155
rect 12280 16995 12320 17125
rect 12280 16965 12285 16995
rect 12315 16965 12320 16995
rect 12280 16960 12320 16965
rect 12360 17155 12400 17160
rect 12360 17125 12365 17155
rect 12395 17125 12400 17155
rect 12360 16995 12400 17125
rect 12360 16965 12365 16995
rect 12395 16965 12400 16995
rect 12360 16960 12400 16965
rect 12440 17155 12480 17160
rect 12440 17125 12445 17155
rect 12475 17125 12480 17155
rect 12440 16995 12480 17125
rect 12440 16965 12445 16995
rect 12475 16965 12480 16995
rect 12440 16960 12480 16965
rect 12520 17155 12560 17160
rect 12520 17125 12525 17155
rect 12555 17125 12560 17155
rect 12520 16995 12560 17125
rect 12520 16965 12525 16995
rect 12555 16965 12560 16995
rect 12520 16960 12560 16965
rect 12600 17155 12640 17160
rect 12600 17125 12605 17155
rect 12635 17125 12640 17155
rect 12600 16995 12640 17125
rect 12600 16965 12605 16995
rect 12635 16965 12640 16995
rect 12600 16960 12640 16965
rect 12680 17155 12720 17160
rect 12680 17125 12685 17155
rect 12715 17125 12720 17155
rect 12680 16995 12720 17125
rect 12680 16965 12685 16995
rect 12715 16965 12720 16995
rect 12680 16960 12720 16965
rect 12760 17155 12800 17160
rect 12760 17125 12765 17155
rect 12795 17125 12800 17155
rect 12760 16995 12800 17125
rect 12760 16965 12765 16995
rect 12795 16965 12800 16995
rect 12760 16960 12800 16965
rect 12840 17155 12880 17160
rect 12840 17125 12845 17155
rect 12875 17125 12880 17155
rect 12840 16995 12880 17125
rect 12840 16965 12845 16995
rect 12875 16965 12880 16995
rect 12840 16960 12880 16965
rect 12920 17155 12960 17160
rect 12920 17125 12925 17155
rect 12955 17125 12960 17155
rect 12920 16995 12960 17125
rect 12920 16965 12925 16995
rect 12955 16965 12960 16995
rect 12920 16960 12960 16965
rect 13000 17155 13040 17160
rect 13000 17125 13005 17155
rect 13035 17125 13040 17155
rect 13000 16995 13040 17125
rect 13000 16965 13005 16995
rect 13035 16965 13040 16995
rect 13000 16960 13040 16965
rect 13080 17155 13120 17160
rect 13080 17125 13085 17155
rect 13115 17125 13120 17155
rect 13080 16995 13120 17125
rect 13080 16965 13085 16995
rect 13115 16965 13120 16995
rect 13080 16960 13120 16965
rect 13160 17155 13200 17160
rect 13160 17125 13165 17155
rect 13195 17125 13200 17155
rect 13160 16995 13200 17125
rect 13160 16965 13165 16995
rect 13195 16965 13200 16995
rect 13160 16960 13200 16965
rect 13240 17155 13280 17160
rect 13240 17125 13245 17155
rect 13275 17125 13280 17155
rect 13240 16995 13280 17125
rect 13240 16965 13245 16995
rect 13275 16965 13280 16995
rect 13240 16960 13280 16965
rect 13320 17155 13360 17160
rect 13320 17125 13325 17155
rect 13355 17125 13360 17155
rect 13320 16995 13360 17125
rect 13320 16965 13325 16995
rect 13355 16965 13360 16995
rect 13320 16960 13360 16965
rect 13400 17155 13440 17160
rect 13400 17125 13405 17155
rect 13435 17125 13440 17155
rect 13400 16995 13440 17125
rect 13400 16965 13405 16995
rect 13435 16965 13440 16995
rect 13400 16960 13440 16965
rect 13480 17155 13520 17160
rect 13480 17125 13485 17155
rect 13515 17125 13520 17155
rect 13480 16995 13520 17125
rect 13480 16965 13485 16995
rect 13515 16965 13520 16995
rect 13480 16960 13520 16965
rect 13560 17155 13600 17160
rect 13560 17125 13565 17155
rect 13595 17125 13600 17155
rect 13560 16995 13600 17125
rect 13560 16965 13565 16995
rect 13595 16965 13600 16995
rect 13560 16960 13600 16965
rect 13640 17155 13680 17160
rect 13640 17125 13645 17155
rect 13675 17125 13680 17155
rect 13640 16995 13680 17125
rect 13640 16965 13645 16995
rect 13675 16965 13680 16995
rect 13640 16960 13680 16965
rect 13720 17155 13760 17160
rect 13720 17125 13725 17155
rect 13755 17125 13760 17155
rect 13720 16995 13760 17125
rect 13720 16965 13725 16995
rect 13755 16965 13760 16995
rect 13720 16960 13760 16965
rect 13800 17155 13840 17160
rect 13800 17125 13805 17155
rect 13835 17125 13840 17155
rect 13800 16995 13840 17125
rect 13800 16965 13805 16995
rect 13835 16965 13840 16995
rect 13800 16960 13840 16965
rect 13880 17155 13920 17160
rect 13880 17125 13885 17155
rect 13915 17125 13920 17155
rect 13880 16995 13920 17125
rect 13880 16965 13885 16995
rect 13915 16965 13920 16995
rect 13880 16960 13920 16965
rect 13960 17155 14000 17160
rect 13960 17125 13965 17155
rect 13995 17125 14000 17155
rect 13960 16995 14000 17125
rect 13960 16965 13965 16995
rect 13995 16965 14000 16995
rect 13960 16960 14000 16965
rect 14040 17155 14080 17160
rect 14040 17125 14045 17155
rect 14075 17125 14080 17155
rect 14040 16995 14080 17125
rect 14040 16965 14045 16995
rect 14075 16965 14080 16995
rect 14040 16960 14080 16965
rect 14120 17155 14160 17160
rect 14120 17125 14125 17155
rect 14155 17125 14160 17155
rect 14120 16995 14160 17125
rect 14120 16965 14125 16995
rect 14155 16965 14160 16995
rect 14120 16960 14160 16965
rect 14200 17155 14240 17160
rect 14200 17125 14205 17155
rect 14235 17125 14240 17155
rect 14200 16995 14240 17125
rect 14200 16965 14205 16995
rect 14235 16965 14240 16995
rect 14200 16960 14240 16965
rect 14280 17155 14320 17160
rect 14280 17125 14285 17155
rect 14315 17125 14320 17155
rect 14280 16995 14320 17125
rect 14280 16965 14285 16995
rect 14315 16965 14320 16995
rect 14280 16960 14320 16965
rect 14360 17155 14400 17160
rect 14360 17125 14365 17155
rect 14395 17125 14400 17155
rect 14360 16995 14400 17125
rect 14360 16965 14365 16995
rect 14395 16965 14400 16995
rect 14360 16960 14400 16965
rect 14440 17155 14480 17160
rect 14440 17125 14445 17155
rect 14475 17125 14480 17155
rect 14440 16995 14480 17125
rect 14440 16965 14445 16995
rect 14475 16965 14480 16995
rect 14440 16960 14480 16965
rect 14520 17155 14560 17160
rect 14520 17125 14525 17155
rect 14555 17125 14560 17155
rect 14520 16995 14560 17125
rect 14520 16965 14525 16995
rect 14555 16965 14560 16995
rect 14520 16960 14560 16965
rect 14600 17155 14640 17160
rect 14600 17125 14605 17155
rect 14635 17125 14640 17155
rect 14600 16995 14640 17125
rect 14600 16965 14605 16995
rect 14635 16965 14640 16995
rect 14600 16960 14640 16965
rect 14680 17155 14720 17160
rect 14680 17125 14685 17155
rect 14715 17125 14720 17155
rect 14680 16995 14720 17125
rect 14680 16965 14685 16995
rect 14715 16965 14720 16995
rect 14680 16960 14720 16965
rect 11560 16915 11600 16920
rect 11560 16885 11565 16915
rect 11595 16885 11600 16915
rect 11560 16755 11600 16885
rect 11560 16725 11565 16755
rect 11595 16725 11600 16755
rect 11560 16720 11600 16725
rect 11640 16915 11680 16920
rect 11640 16885 11645 16915
rect 11675 16885 11680 16915
rect 11640 16755 11680 16885
rect 11640 16725 11645 16755
rect 11675 16725 11680 16755
rect 11640 16720 11680 16725
rect 11720 16915 11760 16920
rect 11720 16885 11725 16915
rect 11755 16885 11760 16915
rect 11720 16755 11760 16885
rect 11720 16725 11725 16755
rect 11755 16725 11760 16755
rect 11720 16720 11760 16725
rect 11800 16915 11840 16920
rect 11800 16885 11805 16915
rect 11835 16885 11840 16915
rect 11800 16755 11840 16885
rect 11800 16725 11805 16755
rect 11835 16725 11840 16755
rect 11800 16720 11840 16725
rect 11880 16915 11920 16920
rect 11880 16885 11885 16915
rect 11915 16885 11920 16915
rect 11880 16755 11920 16885
rect 11880 16725 11885 16755
rect 11915 16725 11920 16755
rect 11880 16720 11920 16725
rect 11960 16915 12000 16920
rect 11960 16885 11965 16915
rect 11995 16885 12000 16915
rect 11960 16755 12000 16885
rect 11960 16725 11965 16755
rect 11995 16725 12000 16755
rect 11960 16720 12000 16725
rect 12040 16915 12080 16920
rect 12040 16885 12045 16915
rect 12075 16885 12080 16915
rect 12040 16755 12080 16885
rect 12040 16725 12045 16755
rect 12075 16725 12080 16755
rect 12040 16720 12080 16725
rect 12120 16915 12160 16920
rect 12120 16885 12125 16915
rect 12155 16885 12160 16915
rect 12120 16755 12160 16885
rect 12120 16725 12125 16755
rect 12155 16725 12160 16755
rect 12120 16720 12160 16725
rect 12200 16915 12240 16920
rect 12200 16885 12205 16915
rect 12235 16885 12240 16915
rect 12200 16755 12240 16885
rect 12200 16725 12205 16755
rect 12235 16725 12240 16755
rect 12200 16720 12240 16725
rect 12280 16915 12320 16920
rect 12280 16885 12285 16915
rect 12315 16885 12320 16915
rect 12280 16755 12320 16885
rect 12280 16725 12285 16755
rect 12315 16725 12320 16755
rect 12280 16720 12320 16725
rect 12360 16915 12400 16920
rect 12360 16885 12365 16915
rect 12395 16885 12400 16915
rect 12360 16755 12400 16885
rect 12360 16725 12365 16755
rect 12395 16725 12400 16755
rect 12360 16720 12400 16725
rect 12440 16915 12480 16920
rect 12440 16885 12445 16915
rect 12475 16885 12480 16915
rect 12440 16755 12480 16885
rect 12440 16725 12445 16755
rect 12475 16725 12480 16755
rect 12440 16720 12480 16725
rect 12520 16915 12560 16920
rect 12520 16885 12525 16915
rect 12555 16885 12560 16915
rect 12520 16755 12560 16885
rect 12520 16725 12525 16755
rect 12555 16725 12560 16755
rect 12520 16720 12560 16725
rect 12600 16915 12640 16920
rect 12600 16885 12605 16915
rect 12635 16885 12640 16915
rect 12600 16755 12640 16885
rect 12600 16725 12605 16755
rect 12635 16725 12640 16755
rect 12600 16720 12640 16725
rect 12680 16915 12720 16920
rect 12680 16885 12685 16915
rect 12715 16885 12720 16915
rect 12680 16755 12720 16885
rect 12680 16725 12685 16755
rect 12715 16725 12720 16755
rect 12680 16720 12720 16725
rect 12760 16915 12800 16920
rect 12760 16885 12765 16915
rect 12795 16885 12800 16915
rect 12760 16755 12800 16885
rect 12760 16725 12765 16755
rect 12795 16725 12800 16755
rect 12760 16720 12800 16725
rect 12840 16915 12880 16920
rect 12840 16885 12845 16915
rect 12875 16885 12880 16915
rect 12840 16755 12880 16885
rect 12840 16725 12845 16755
rect 12875 16725 12880 16755
rect 12840 16720 12880 16725
rect 12920 16915 12960 16920
rect 12920 16885 12925 16915
rect 12955 16885 12960 16915
rect 12920 16755 12960 16885
rect 12920 16725 12925 16755
rect 12955 16725 12960 16755
rect 12920 16720 12960 16725
rect 13000 16915 13040 16920
rect 13000 16885 13005 16915
rect 13035 16885 13040 16915
rect 13000 16755 13040 16885
rect 13000 16725 13005 16755
rect 13035 16725 13040 16755
rect 13000 16720 13040 16725
rect 13080 16915 13120 16920
rect 13080 16885 13085 16915
rect 13115 16885 13120 16915
rect 13080 16755 13120 16885
rect 13080 16725 13085 16755
rect 13115 16725 13120 16755
rect 13080 16720 13120 16725
rect 13160 16915 13200 16920
rect 13160 16885 13165 16915
rect 13195 16885 13200 16915
rect 13160 16755 13200 16885
rect 13160 16725 13165 16755
rect 13195 16725 13200 16755
rect 13160 16720 13200 16725
rect 13240 16915 13280 16920
rect 13240 16885 13245 16915
rect 13275 16885 13280 16915
rect 13240 16755 13280 16885
rect 13240 16725 13245 16755
rect 13275 16725 13280 16755
rect 13240 16720 13280 16725
rect 13320 16915 13360 16920
rect 13320 16885 13325 16915
rect 13355 16885 13360 16915
rect 13320 16755 13360 16885
rect 13320 16725 13325 16755
rect 13355 16725 13360 16755
rect 13320 16720 13360 16725
rect 13400 16915 13440 16920
rect 13400 16885 13405 16915
rect 13435 16885 13440 16915
rect 13400 16755 13440 16885
rect 13400 16725 13405 16755
rect 13435 16725 13440 16755
rect 13400 16720 13440 16725
rect 13480 16915 13520 16920
rect 13480 16885 13485 16915
rect 13515 16885 13520 16915
rect 13480 16755 13520 16885
rect 13480 16725 13485 16755
rect 13515 16725 13520 16755
rect 13480 16720 13520 16725
rect 13560 16915 13600 16920
rect 13560 16885 13565 16915
rect 13595 16885 13600 16915
rect 13560 16755 13600 16885
rect 13560 16725 13565 16755
rect 13595 16725 13600 16755
rect 13560 16720 13600 16725
rect 13640 16915 13680 16920
rect 13640 16885 13645 16915
rect 13675 16885 13680 16915
rect 13640 16755 13680 16885
rect 13640 16725 13645 16755
rect 13675 16725 13680 16755
rect 13640 16720 13680 16725
rect 13720 16915 13760 16920
rect 13720 16885 13725 16915
rect 13755 16885 13760 16915
rect 13720 16755 13760 16885
rect 13720 16725 13725 16755
rect 13755 16725 13760 16755
rect 13720 16720 13760 16725
rect 13800 16915 13840 16920
rect 13800 16885 13805 16915
rect 13835 16885 13840 16915
rect 13800 16755 13840 16885
rect 13800 16725 13805 16755
rect 13835 16725 13840 16755
rect 13800 16720 13840 16725
rect 13880 16915 13920 16920
rect 13880 16885 13885 16915
rect 13915 16885 13920 16915
rect 13880 16755 13920 16885
rect 13880 16725 13885 16755
rect 13915 16725 13920 16755
rect 13880 16720 13920 16725
rect 13960 16915 14000 16920
rect 13960 16885 13965 16915
rect 13995 16885 14000 16915
rect 13960 16755 14000 16885
rect 13960 16725 13965 16755
rect 13995 16725 14000 16755
rect 13960 16720 14000 16725
rect 14040 16915 14080 16920
rect 14040 16885 14045 16915
rect 14075 16885 14080 16915
rect 14040 16755 14080 16885
rect 14040 16725 14045 16755
rect 14075 16725 14080 16755
rect 14040 16720 14080 16725
rect 14120 16915 14160 16920
rect 14120 16885 14125 16915
rect 14155 16885 14160 16915
rect 14120 16755 14160 16885
rect 14120 16725 14125 16755
rect 14155 16725 14160 16755
rect 14120 16720 14160 16725
rect 14200 16915 14240 16920
rect 14200 16885 14205 16915
rect 14235 16885 14240 16915
rect 14200 16755 14240 16885
rect 14200 16725 14205 16755
rect 14235 16725 14240 16755
rect 14200 16720 14240 16725
rect 14280 16915 14320 16920
rect 14280 16885 14285 16915
rect 14315 16885 14320 16915
rect 14280 16755 14320 16885
rect 14280 16725 14285 16755
rect 14315 16725 14320 16755
rect 14280 16720 14320 16725
rect 14360 16915 14400 16920
rect 14360 16885 14365 16915
rect 14395 16885 14400 16915
rect 14360 16755 14400 16885
rect 14360 16725 14365 16755
rect 14395 16725 14400 16755
rect 14360 16720 14400 16725
rect 14440 16915 14480 16920
rect 14440 16885 14445 16915
rect 14475 16885 14480 16915
rect 14440 16755 14480 16885
rect 14440 16725 14445 16755
rect 14475 16725 14480 16755
rect 14440 16720 14480 16725
rect 14520 16915 14560 16920
rect 14520 16885 14525 16915
rect 14555 16885 14560 16915
rect 14520 16755 14560 16885
rect 14520 16725 14525 16755
rect 14555 16725 14560 16755
rect 14520 16720 14560 16725
rect 14600 16915 14640 16920
rect 14600 16885 14605 16915
rect 14635 16885 14640 16915
rect 14600 16755 14640 16885
rect 14600 16725 14605 16755
rect 14635 16725 14640 16755
rect 14600 16720 14640 16725
rect 14680 16915 14720 16920
rect 14680 16885 14685 16915
rect 14715 16885 14720 16915
rect 14680 16755 14720 16885
rect 14680 16725 14685 16755
rect 14715 16725 14720 16755
rect 14680 16720 14720 16725
rect 14760 16915 14800 18720
rect 14760 16885 14765 16915
rect 14795 16885 14800 16915
rect 14760 16755 14800 16885
rect 14760 16725 14765 16755
rect 14795 16725 14800 16755
rect 14760 16720 14800 16725
rect 14840 16835 14880 18720
rect 14840 16805 14845 16835
rect 14875 16805 14880 16835
rect 14840 16720 14880 16805
rect 14920 16915 14960 18720
rect 14920 16885 14925 16915
rect 14955 16885 14960 16915
rect 14920 16755 14960 16885
rect 14920 16725 14925 16755
rect 14955 16725 14960 16755
rect 14920 16720 14960 16725
rect 15000 17155 15040 18720
rect 15000 17125 15005 17155
rect 15035 17125 15040 17155
rect 15000 16995 15040 17125
rect 15000 16965 15005 16995
rect 15035 16965 15040 16995
rect 15000 16720 15040 16965
rect 15080 17075 15120 18720
rect 15080 17045 15085 17075
rect 15115 17045 15120 17075
rect 15080 16720 15120 17045
rect 15160 17155 15200 18720
rect 15160 17125 15165 17155
rect 15195 17125 15200 17155
rect 15160 16995 15200 17125
rect 15160 16965 15165 16995
rect 15195 16965 15200 16995
rect 15160 16720 15200 16965
rect 15240 18195 15280 18720
rect 15240 18165 15245 18195
rect 15275 18165 15280 18195
rect 15240 18035 15280 18165
rect 15240 18005 15245 18035
rect 15275 18005 15280 18035
rect 15240 17875 15280 18005
rect 15240 17845 15245 17875
rect 15275 17845 15280 17875
rect 15240 17715 15280 17845
rect 15240 17685 15245 17715
rect 15275 17685 15280 17715
rect 15240 17555 15280 17685
rect 15240 17525 15245 17555
rect 15275 17525 15280 17555
rect 15240 17395 15280 17525
rect 15240 17365 15245 17395
rect 15275 17365 15280 17395
rect 15240 17235 15280 17365
rect 15240 17205 15245 17235
rect 15275 17205 15280 17235
rect 15240 16720 15280 17205
rect 15320 17315 15360 18720
rect 15320 17285 15325 17315
rect 15355 17285 15360 17315
rect 15320 16720 15360 17285
rect 15400 18195 15440 18720
rect 15400 18165 15405 18195
rect 15435 18165 15440 18195
rect 15400 18035 15440 18165
rect 15400 18005 15405 18035
rect 15435 18005 15440 18035
rect 15400 17875 15440 18005
rect 15400 17845 15405 17875
rect 15435 17845 15440 17875
rect 15400 17715 15440 17845
rect 15400 17685 15405 17715
rect 15435 17685 15440 17715
rect 15400 17555 15440 17685
rect 15400 17525 15405 17555
rect 15435 17525 15440 17555
rect 15400 17395 15440 17525
rect 15400 17365 15405 17395
rect 15435 17365 15440 17395
rect 15400 17235 15440 17365
rect 15400 17205 15405 17235
rect 15435 17205 15440 17235
rect 15400 16720 15440 17205
rect 15480 17475 15520 18720
rect 15480 17445 15485 17475
rect 15515 17445 15520 17475
rect 15480 16720 15520 17445
rect 15560 18195 15600 18720
rect 15560 18165 15565 18195
rect 15595 18165 15600 18195
rect 15560 18035 15600 18165
rect 15560 18005 15565 18035
rect 15595 18005 15600 18035
rect 15560 17875 15600 18005
rect 15560 17845 15565 17875
rect 15595 17845 15600 17875
rect 15560 17715 15600 17845
rect 15560 17685 15565 17715
rect 15595 17685 15600 17715
rect 15560 17555 15600 17685
rect 15560 17525 15565 17555
rect 15595 17525 15600 17555
rect 15560 17395 15600 17525
rect 15560 17365 15565 17395
rect 15595 17365 15600 17395
rect 15560 17235 15600 17365
rect 15560 17205 15565 17235
rect 15595 17205 15600 17235
rect 15560 16720 15600 17205
rect 15640 17635 15680 18720
rect 15640 17605 15645 17635
rect 15675 17605 15680 17635
rect 15640 16720 15680 17605
rect 15720 18195 15760 18720
rect 15720 18165 15725 18195
rect 15755 18165 15760 18195
rect 15720 18035 15760 18165
rect 15720 18005 15725 18035
rect 15755 18005 15760 18035
rect 15720 17875 15760 18005
rect 15720 17845 15725 17875
rect 15755 17845 15760 17875
rect 15720 17715 15760 17845
rect 15720 17685 15725 17715
rect 15755 17685 15760 17715
rect 15720 17555 15760 17685
rect 15720 17525 15725 17555
rect 15755 17525 15760 17555
rect 15720 17395 15760 17525
rect 15720 17365 15725 17395
rect 15755 17365 15760 17395
rect 15720 17235 15760 17365
rect 15720 17205 15725 17235
rect 15755 17205 15760 17235
rect 15720 16720 15760 17205
rect 15800 17795 15840 18720
rect 15800 17765 15805 17795
rect 15835 17765 15840 17795
rect 15800 16720 15840 17765
rect 15880 18195 15920 18720
rect 15880 18165 15885 18195
rect 15915 18165 15920 18195
rect 15880 18035 15920 18165
rect 15880 18005 15885 18035
rect 15915 18005 15920 18035
rect 15880 17875 15920 18005
rect 15880 17845 15885 17875
rect 15915 17845 15920 17875
rect 15880 17715 15920 17845
rect 15880 17685 15885 17715
rect 15915 17685 15920 17715
rect 15880 17555 15920 17685
rect 15880 17525 15885 17555
rect 15915 17525 15920 17555
rect 15880 17395 15920 17525
rect 15880 17365 15885 17395
rect 15915 17365 15920 17395
rect 15880 17235 15920 17365
rect 15880 17205 15885 17235
rect 15915 17205 15920 17235
rect 15880 16720 15920 17205
rect 15960 17955 16000 18720
rect 15960 17925 15965 17955
rect 15995 17925 16000 17955
rect 15960 16720 16000 17925
rect 16040 18195 16080 18720
rect 16040 18165 16045 18195
rect 16075 18165 16080 18195
rect 16040 18035 16080 18165
rect 16040 18005 16045 18035
rect 16075 18005 16080 18035
rect 16040 17875 16080 18005
rect 16040 17845 16045 17875
rect 16075 17845 16080 17875
rect 16040 17715 16080 17845
rect 16040 17685 16045 17715
rect 16075 17685 16080 17715
rect 16040 17555 16080 17685
rect 16040 17525 16045 17555
rect 16075 17525 16080 17555
rect 16040 17395 16080 17525
rect 16040 17365 16045 17395
rect 16075 17365 16080 17395
rect 16040 17235 16080 17365
rect 16040 17205 16045 17235
rect 16075 17205 16080 17235
rect 16040 16720 16080 17205
rect 16120 18115 16160 18720
rect 16120 18085 16125 18115
rect 16155 18085 16160 18115
rect 16120 16720 16160 18085
rect 16200 18195 16240 18720
rect 16200 18165 16205 18195
rect 16235 18165 16240 18195
rect 16200 18035 16240 18165
rect 16200 18005 16205 18035
rect 16235 18005 16240 18035
rect 16200 17875 16240 18005
rect 16200 17845 16205 17875
rect 16235 17845 16240 17875
rect 16200 17715 16240 17845
rect 16200 17685 16205 17715
rect 16235 17685 16240 17715
rect 16200 17555 16240 17685
rect 16200 17525 16205 17555
rect 16235 17525 16240 17555
rect 16200 17395 16240 17525
rect 16200 17365 16205 17395
rect 16235 17365 16240 17395
rect 16200 17235 16240 17365
rect 16200 17205 16205 17235
rect 16235 17205 16240 17235
rect 16200 16720 16240 17205
rect 16280 18435 16320 18720
rect 16280 18405 16285 18435
rect 16315 18405 16320 18435
rect 16280 18275 16320 18405
rect 16280 18245 16285 18275
rect 16315 18245 16320 18275
rect 16280 16720 16320 18245
rect 16360 18355 16400 18720
rect 16360 18325 16365 18355
rect 16395 18325 16400 18355
rect 16360 16720 16400 18325
rect 16440 18435 16480 18720
rect 16440 18405 16445 18435
rect 16475 18405 16480 18435
rect 16440 18275 16480 18405
rect 16440 18245 16445 18275
rect 16475 18245 16480 18275
rect 16440 16720 16480 18245
rect 16520 18675 16560 18720
rect 16520 18645 16525 18675
rect 16555 18645 16560 18675
rect 16520 18515 16560 18645
rect 16520 18485 16525 18515
rect 16555 18485 16560 18515
rect 16520 16720 16560 18485
rect 16600 18595 16640 18720
rect 16600 18565 16605 18595
rect 16635 18565 16640 18595
rect 16600 16720 16640 18565
rect 16680 18675 16720 18720
rect 16680 18645 16685 18675
rect 16715 18645 16720 18675
rect 16680 18515 16720 18645
rect 16680 18485 16685 18515
rect 16715 18485 16720 18515
rect 16680 16720 16720 18485
rect 16760 18675 16800 18680
rect 16760 18645 16765 18675
rect 16795 18645 16800 18675
rect 16760 18515 16800 18645
rect 16760 18485 16765 18515
rect 16795 18485 16800 18515
rect 16760 18480 16800 18485
rect 16840 18675 16880 18680
rect 16840 18645 16845 18675
rect 16875 18645 16880 18675
rect 16840 18515 16880 18645
rect 16840 18485 16845 18515
rect 16875 18485 16880 18515
rect 16840 18480 16880 18485
rect 16920 18675 16960 18680
rect 16920 18645 16925 18675
rect 16955 18645 16960 18675
rect 16920 18515 16960 18645
rect 16920 18485 16925 18515
rect 16955 18485 16960 18515
rect 16920 18480 16960 18485
rect 17000 18675 17040 18680
rect 17000 18645 17005 18675
rect 17035 18645 17040 18675
rect 17000 18515 17040 18645
rect 17000 18485 17005 18515
rect 17035 18485 17040 18515
rect 17000 18480 17040 18485
rect 17080 18675 17120 18680
rect 17080 18645 17085 18675
rect 17115 18645 17120 18675
rect 17080 18515 17120 18645
rect 17080 18485 17085 18515
rect 17115 18485 17120 18515
rect 17080 18480 17120 18485
rect 17160 18675 17200 18680
rect 17160 18645 17165 18675
rect 17195 18645 17200 18675
rect 17160 18515 17200 18645
rect 17160 18485 17165 18515
rect 17195 18485 17200 18515
rect 17160 18480 17200 18485
rect 17240 18675 17280 18680
rect 17240 18645 17245 18675
rect 17275 18645 17280 18675
rect 17240 18515 17280 18645
rect 17240 18485 17245 18515
rect 17275 18485 17280 18515
rect 17240 18480 17280 18485
rect 17320 18675 17360 18680
rect 17320 18645 17325 18675
rect 17355 18645 17360 18675
rect 17320 18515 17360 18645
rect 17320 18485 17325 18515
rect 17355 18485 17360 18515
rect 17320 18480 17360 18485
rect 17400 18675 17440 18680
rect 17400 18645 17405 18675
rect 17435 18645 17440 18675
rect 17400 18515 17440 18645
rect 17400 18485 17405 18515
rect 17435 18485 17440 18515
rect 17400 18480 17440 18485
rect 17480 18675 17520 18680
rect 17480 18645 17485 18675
rect 17515 18645 17520 18675
rect 17480 18515 17520 18645
rect 17480 18485 17485 18515
rect 17515 18485 17520 18515
rect 17480 18480 17520 18485
rect 17560 18675 17600 18680
rect 17560 18645 17565 18675
rect 17595 18645 17600 18675
rect 17560 18515 17600 18645
rect 17560 18485 17565 18515
rect 17595 18485 17600 18515
rect 17560 18480 17600 18485
rect 17640 18675 17680 18680
rect 17640 18645 17645 18675
rect 17675 18645 17680 18675
rect 17640 18515 17680 18645
rect 17640 18485 17645 18515
rect 17675 18485 17680 18515
rect 17640 18480 17680 18485
rect 17720 18675 17760 18680
rect 17720 18645 17725 18675
rect 17755 18645 17760 18675
rect 17720 18515 17760 18645
rect 17720 18485 17725 18515
rect 17755 18485 17760 18515
rect 17720 18480 17760 18485
rect 17800 18675 17840 18680
rect 17800 18645 17805 18675
rect 17835 18645 17840 18675
rect 17800 18515 17840 18645
rect 17800 18485 17805 18515
rect 17835 18485 17840 18515
rect 17800 18480 17840 18485
rect 17880 18675 17920 18680
rect 17880 18645 17885 18675
rect 17915 18645 17920 18675
rect 17880 18515 17920 18645
rect 17880 18485 17885 18515
rect 17915 18485 17920 18515
rect 17880 18480 17920 18485
rect 17960 18675 18000 18680
rect 17960 18645 17965 18675
rect 17995 18645 18000 18675
rect 17960 18515 18000 18645
rect 17960 18485 17965 18515
rect 17995 18485 18000 18515
rect 17960 18480 18000 18485
rect 18040 18675 18080 18680
rect 18040 18645 18045 18675
rect 18075 18645 18080 18675
rect 18040 18515 18080 18645
rect 18040 18485 18045 18515
rect 18075 18485 18080 18515
rect 18040 18480 18080 18485
rect 18120 18675 18160 18680
rect 18120 18645 18125 18675
rect 18155 18645 18160 18675
rect 18120 18515 18160 18645
rect 18120 18485 18125 18515
rect 18155 18485 18160 18515
rect 18120 18480 18160 18485
rect 18200 18675 18240 18680
rect 18200 18645 18205 18675
rect 18235 18645 18240 18675
rect 18200 18515 18240 18645
rect 18200 18485 18205 18515
rect 18235 18485 18240 18515
rect 18200 18480 18240 18485
rect 18280 18675 18320 18680
rect 18280 18645 18285 18675
rect 18315 18645 18320 18675
rect 18280 18515 18320 18645
rect 18280 18485 18285 18515
rect 18315 18485 18320 18515
rect 18280 18480 18320 18485
rect 18360 18675 18400 18680
rect 18360 18645 18365 18675
rect 18395 18645 18400 18675
rect 18360 18515 18400 18645
rect 18360 18485 18365 18515
rect 18395 18485 18400 18515
rect 18360 18480 18400 18485
rect 18440 18675 18480 18680
rect 18440 18645 18445 18675
rect 18475 18645 18480 18675
rect 18440 18515 18480 18645
rect 18440 18485 18445 18515
rect 18475 18485 18480 18515
rect 18440 18480 18480 18485
rect 18520 18675 18560 18680
rect 18520 18645 18525 18675
rect 18555 18645 18560 18675
rect 18520 18515 18560 18645
rect 18520 18485 18525 18515
rect 18555 18485 18560 18515
rect 18520 18480 18560 18485
rect 18600 18675 18640 18680
rect 18600 18645 18605 18675
rect 18635 18645 18640 18675
rect 18600 18515 18640 18645
rect 18600 18485 18605 18515
rect 18635 18485 18640 18515
rect 18600 18480 18640 18485
rect 18680 18675 18720 18680
rect 18680 18645 18685 18675
rect 18715 18645 18720 18675
rect 18680 18515 18720 18645
rect 18680 18485 18685 18515
rect 18715 18485 18720 18515
rect 18680 18480 18720 18485
rect 18760 18675 18800 18680
rect 18760 18645 18765 18675
rect 18795 18645 18800 18675
rect 18760 18515 18800 18645
rect 18760 18485 18765 18515
rect 18795 18485 18800 18515
rect 18760 18480 18800 18485
rect 18840 18675 18880 18680
rect 18840 18645 18845 18675
rect 18875 18645 18880 18675
rect 18840 18515 18880 18645
rect 18840 18485 18845 18515
rect 18875 18485 18880 18515
rect 18840 18480 18880 18485
rect 18920 18675 18960 18680
rect 18920 18645 18925 18675
rect 18955 18645 18960 18675
rect 18920 18515 18960 18645
rect 18920 18485 18925 18515
rect 18955 18485 18960 18515
rect 18920 18480 18960 18485
rect 19000 18675 19040 18680
rect 19000 18645 19005 18675
rect 19035 18645 19040 18675
rect 19000 18515 19040 18645
rect 19000 18485 19005 18515
rect 19035 18485 19040 18515
rect 19000 18480 19040 18485
rect 19080 18675 19120 18680
rect 19080 18645 19085 18675
rect 19115 18645 19120 18675
rect 19080 18515 19120 18645
rect 19080 18485 19085 18515
rect 19115 18485 19120 18515
rect 19080 18480 19120 18485
rect 19160 18675 19200 18680
rect 19160 18645 19165 18675
rect 19195 18645 19200 18675
rect 19160 18515 19200 18645
rect 19160 18485 19165 18515
rect 19195 18485 19200 18515
rect 19160 18480 19200 18485
rect 19240 18675 19280 18680
rect 19240 18645 19245 18675
rect 19275 18645 19280 18675
rect 19240 18515 19280 18645
rect 19240 18485 19245 18515
rect 19275 18485 19280 18515
rect 19240 18480 19280 18485
rect 19320 18675 19360 18680
rect 19320 18645 19325 18675
rect 19355 18645 19360 18675
rect 19320 18515 19360 18645
rect 19320 18485 19325 18515
rect 19355 18485 19360 18515
rect 19320 18480 19360 18485
rect 19400 18675 19440 18680
rect 19400 18645 19405 18675
rect 19435 18645 19440 18675
rect 19400 18515 19440 18645
rect 19400 18485 19405 18515
rect 19435 18485 19440 18515
rect 19400 18480 19440 18485
rect 19480 18675 19520 18680
rect 19480 18645 19485 18675
rect 19515 18645 19520 18675
rect 19480 18515 19520 18645
rect 19480 18485 19485 18515
rect 19515 18485 19520 18515
rect 19480 18480 19520 18485
rect 19560 18675 19600 18680
rect 19560 18645 19565 18675
rect 19595 18645 19600 18675
rect 19560 18515 19600 18645
rect 19560 18485 19565 18515
rect 19595 18485 19600 18515
rect 19560 18480 19600 18485
rect 19640 18675 19680 18680
rect 19640 18645 19645 18675
rect 19675 18645 19680 18675
rect 19640 18515 19680 18645
rect 19640 18485 19645 18515
rect 19675 18485 19680 18515
rect 19640 18480 19680 18485
rect 19720 18675 19760 18680
rect 19720 18645 19725 18675
rect 19755 18645 19760 18675
rect 19720 18515 19760 18645
rect 19720 18485 19725 18515
rect 19755 18485 19760 18515
rect 19720 18480 19760 18485
rect 19800 18675 19840 18680
rect 19800 18645 19805 18675
rect 19835 18645 19840 18675
rect 19800 18515 19840 18645
rect 19800 18485 19805 18515
rect 19835 18485 19840 18515
rect 19800 18480 19840 18485
rect 19880 18675 19920 18680
rect 19880 18645 19885 18675
rect 19915 18645 19920 18675
rect 19880 18515 19920 18645
rect 19880 18485 19885 18515
rect 19915 18485 19920 18515
rect 19880 18480 19920 18485
rect 19960 18675 20000 18680
rect 19960 18645 19965 18675
rect 19995 18645 20000 18675
rect 19960 18515 20000 18645
rect 19960 18485 19965 18515
rect 19995 18485 20000 18515
rect 19960 18480 20000 18485
rect 20040 18675 20080 18680
rect 20040 18645 20045 18675
rect 20075 18645 20080 18675
rect 20040 18515 20080 18645
rect 20040 18485 20045 18515
rect 20075 18485 20080 18515
rect 20040 18480 20080 18485
rect 20120 18675 20160 18680
rect 20120 18645 20125 18675
rect 20155 18645 20160 18675
rect 20120 18515 20160 18645
rect 20120 18485 20125 18515
rect 20155 18485 20160 18515
rect 20120 18480 20160 18485
rect 20200 18675 20240 18680
rect 20200 18645 20205 18675
rect 20235 18645 20240 18675
rect 20200 18515 20240 18645
rect 20200 18485 20205 18515
rect 20235 18485 20240 18515
rect 20200 18480 20240 18485
rect 20280 18675 20320 18680
rect 20280 18645 20285 18675
rect 20315 18645 20320 18675
rect 20280 18515 20320 18645
rect 20280 18485 20285 18515
rect 20315 18485 20320 18515
rect 20280 18480 20320 18485
rect 20360 18675 20400 18680
rect 20360 18645 20365 18675
rect 20395 18645 20400 18675
rect 20360 18515 20400 18645
rect 20360 18485 20365 18515
rect 20395 18485 20400 18515
rect 20360 18480 20400 18485
rect 20440 18675 20480 18680
rect 20440 18645 20445 18675
rect 20475 18645 20480 18675
rect 20440 18515 20480 18645
rect 20440 18485 20445 18515
rect 20475 18485 20480 18515
rect 20440 18480 20480 18485
rect 20520 18675 20560 18680
rect 20520 18645 20525 18675
rect 20555 18645 20560 18675
rect 20520 18515 20560 18645
rect 20520 18485 20525 18515
rect 20555 18485 20560 18515
rect 20520 18480 20560 18485
rect 20600 18675 20640 18680
rect 20600 18645 20605 18675
rect 20635 18645 20640 18675
rect 20600 18515 20640 18645
rect 20600 18485 20605 18515
rect 20635 18485 20640 18515
rect 20600 18480 20640 18485
rect 20680 18675 20720 18680
rect 20680 18645 20685 18675
rect 20715 18645 20720 18675
rect 20680 18515 20720 18645
rect 20680 18485 20685 18515
rect 20715 18485 20720 18515
rect 20680 18480 20720 18485
rect 20760 18675 20800 18680
rect 20760 18645 20765 18675
rect 20795 18645 20800 18675
rect 20760 18515 20800 18645
rect 20760 18485 20765 18515
rect 20795 18485 20800 18515
rect 20760 18480 20800 18485
rect 20840 18675 20880 18680
rect 20840 18645 20845 18675
rect 20875 18645 20880 18675
rect 20840 18515 20880 18645
rect 20840 18485 20845 18515
rect 20875 18485 20880 18515
rect 20840 18480 20880 18485
rect 20920 18675 20960 18680
rect 20920 18645 20925 18675
rect 20955 18645 20960 18675
rect 20920 18515 20960 18645
rect 20920 18485 20925 18515
rect 20955 18485 20960 18515
rect 20920 18480 20960 18485
rect 16760 18435 16800 18440
rect 16760 18405 16765 18435
rect 16795 18405 16800 18435
rect 16760 18275 16800 18405
rect 16760 18245 16765 18275
rect 16795 18245 16800 18275
rect 16760 18240 16800 18245
rect 16840 18435 16880 18440
rect 16840 18405 16845 18435
rect 16875 18405 16880 18435
rect 16840 18275 16880 18405
rect 16840 18245 16845 18275
rect 16875 18245 16880 18275
rect 16840 18240 16880 18245
rect 16920 18435 16960 18440
rect 16920 18405 16925 18435
rect 16955 18405 16960 18435
rect 16920 18275 16960 18405
rect 16920 18245 16925 18275
rect 16955 18245 16960 18275
rect 16920 18240 16960 18245
rect 17000 18435 17040 18440
rect 17000 18405 17005 18435
rect 17035 18405 17040 18435
rect 17000 18275 17040 18405
rect 17000 18245 17005 18275
rect 17035 18245 17040 18275
rect 17000 18240 17040 18245
rect 17080 18435 17120 18440
rect 17080 18405 17085 18435
rect 17115 18405 17120 18435
rect 17080 18275 17120 18405
rect 17080 18245 17085 18275
rect 17115 18245 17120 18275
rect 17080 18240 17120 18245
rect 17160 18435 17200 18440
rect 17160 18405 17165 18435
rect 17195 18405 17200 18435
rect 17160 18275 17200 18405
rect 17160 18245 17165 18275
rect 17195 18245 17200 18275
rect 17160 18240 17200 18245
rect 17240 18435 17280 18440
rect 17240 18405 17245 18435
rect 17275 18405 17280 18435
rect 17240 18275 17280 18405
rect 17240 18245 17245 18275
rect 17275 18245 17280 18275
rect 17240 18240 17280 18245
rect 17320 18435 17360 18440
rect 17320 18405 17325 18435
rect 17355 18405 17360 18435
rect 17320 18275 17360 18405
rect 17320 18245 17325 18275
rect 17355 18245 17360 18275
rect 17320 18240 17360 18245
rect 17400 18435 17440 18440
rect 17400 18405 17405 18435
rect 17435 18405 17440 18435
rect 17400 18275 17440 18405
rect 17400 18245 17405 18275
rect 17435 18245 17440 18275
rect 17400 18240 17440 18245
rect 17480 18435 17520 18440
rect 17480 18405 17485 18435
rect 17515 18405 17520 18435
rect 17480 18275 17520 18405
rect 17480 18245 17485 18275
rect 17515 18245 17520 18275
rect 17480 18240 17520 18245
rect 17560 18435 17600 18440
rect 17560 18405 17565 18435
rect 17595 18405 17600 18435
rect 17560 18275 17600 18405
rect 17560 18245 17565 18275
rect 17595 18245 17600 18275
rect 17560 18240 17600 18245
rect 17640 18435 17680 18440
rect 17640 18405 17645 18435
rect 17675 18405 17680 18435
rect 17640 18275 17680 18405
rect 17640 18245 17645 18275
rect 17675 18245 17680 18275
rect 17640 18240 17680 18245
rect 17720 18435 17760 18440
rect 17720 18405 17725 18435
rect 17755 18405 17760 18435
rect 17720 18275 17760 18405
rect 17720 18245 17725 18275
rect 17755 18245 17760 18275
rect 17720 18240 17760 18245
rect 17800 18435 17840 18440
rect 17800 18405 17805 18435
rect 17835 18405 17840 18435
rect 17800 18275 17840 18405
rect 17800 18245 17805 18275
rect 17835 18245 17840 18275
rect 17800 18240 17840 18245
rect 17880 18435 17920 18440
rect 17880 18405 17885 18435
rect 17915 18405 17920 18435
rect 17880 18275 17920 18405
rect 17880 18245 17885 18275
rect 17915 18245 17920 18275
rect 17880 18240 17920 18245
rect 17960 18435 18000 18440
rect 17960 18405 17965 18435
rect 17995 18405 18000 18435
rect 17960 18275 18000 18405
rect 17960 18245 17965 18275
rect 17995 18245 18000 18275
rect 17960 18240 18000 18245
rect 18040 18435 18080 18440
rect 18040 18405 18045 18435
rect 18075 18405 18080 18435
rect 18040 18275 18080 18405
rect 18040 18245 18045 18275
rect 18075 18245 18080 18275
rect 18040 18240 18080 18245
rect 18120 18435 18160 18440
rect 18120 18405 18125 18435
rect 18155 18405 18160 18435
rect 18120 18275 18160 18405
rect 18120 18245 18125 18275
rect 18155 18245 18160 18275
rect 18120 18240 18160 18245
rect 18200 18435 18240 18440
rect 18200 18405 18205 18435
rect 18235 18405 18240 18435
rect 18200 18275 18240 18405
rect 18200 18245 18205 18275
rect 18235 18245 18240 18275
rect 18200 18240 18240 18245
rect 18280 18435 18320 18440
rect 18280 18405 18285 18435
rect 18315 18405 18320 18435
rect 18280 18275 18320 18405
rect 18280 18245 18285 18275
rect 18315 18245 18320 18275
rect 18280 18240 18320 18245
rect 18360 18435 18400 18440
rect 18360 18405 18365 18435
rect 18395 18405 18400 18435
rect 18360 18275 18400 18405
rect 18360 18245 18365 18275
rect 18395 18245 18400 18275
rect 18360 18240 18400 18245
rect 18440 18435 18480 18440
rect 18440 18405 18445 18435
rect 18475 18405 18480 18435
rect 18440 18275 18480 18405
rect 18440 18245 18445 18275
rect 18475 18245 18480 18275
rect 18440 18240 18480 18245
rect 18520 18435 18560 18440
rect 18520 18405 18525 18435
rect 18555 18405 18560 18435
rect 18520 18275 18560 18405
rect 18520 18245 18525 18275
rect 18555 18245 18560 18275
rect 18520 18240 18560 18245
rect 18600 18435 18640 18440
rect 18600 18405 18605 18435
rect 18635 18405 18640 18435
rect 18600 18275 18640 18405
rect 18600 18245 18605 18275
rect 18635 18245 18640 18275
rect 18600 18240 18640 18245
rect 18680 18435 18720 18440
rect 18680 18405 18685 18435
rect 18715 18405 18720 18435
rect 18680 18275 18720 18405
rect 18680 18245 18685 18275
rect 18715 18245 18720 18275
rect 18680 18240 18720 18245
rect 18760 18435 18800 18440
rect 18760 18405 18765 18435
rect 18795 18405 18800 18435
rect 18760 18275 18800 18405
rect 18760 18245 18765 18275
rect 18795 18245 18800 18275
rect 18760 18240 18800 18245
rect 18840 18435 18880 18440
rect 18840 18405 18845 18435
rect 18875 18405 18880 18435
rect 18840 18275 18880 18405
rect 18840 18245 18845 18275
rect 18875 18245 18880 18275
rect 18840 18240 18880 18245
rect 18920 18435 18960 18440
rect 18920 18405 18925 18435
rect 18955 18405 18960 18435
rect 18920 18275 18960 18405
rect 18920 18245 18925 18275
rect 18955 18245 18960 18275
rect 18920 18240 18960 18245
rect 19000 18435 19040 18440
rect 19000 18405 19005 18435
rect 19035 18405 19040 18435
rect 19000 18275 19040 18405
rect 19000 18245 19005 18275
rect 19035 18245 19040 18275
rect 19000 18240 19040 18245
rect 19080 18435 19120 18440
rect 19080 18405 19085 18435
rect 19115 18405 19120 18435
rect 19080 18275 19120 18405
rect 19080 18245 19085 18275
rect 19115 18245 19120 18275
rect 19080 18240 19120 18245
rect 19160 18435 19200 18440
rect 19160 18405 19165 18435
rect 19195 18405 19200 18435
rect 19160 18275 19200 18405
rect 19160 18245 19165 18275
rect 19195 18245 19200 18275
rect 19160 18240 19200 18245
rect 19240 18435 19280 18440
rect 19240 18405 19245 18435
rect 19275 18405 19280 18435
rect 19240 18275 19280 18405
rect 19240 18245 19245 18275
rect 19275 18245 19280 18275
rect 19240 18240 19280 18245
rect 19320 18435 19360 18440
rect 19320 18405 19325 18435
rect 19355 18405 19360 18435
rect 19320 18275 19360 18405
rect 19320 18245 19325 18275
rect 19355 18245 19360 18275
rect 19320 18240 19360 18245
rect 19400 18435 19440 18440
rect 19400 18405 19405 18435
rect 19435 18405 19440 18435
rect 19400 18275 19440 18405
rect 19400 18245 19405 18275
rect 19435 18245 19440 18275
rect 19400 18240 19440 18245
rect 19480 18435 19520 18440
rect 19480 18405 19485 18435
rect 19515 18405 19520 18435
rect 19480 18275 19520 18405
rect 19480 18245 19485 18275
rect 19515 18245 19520 18275
rect 19480 18240 19520 18245
rect 19560 18435 19600 18440
rect 19560 18405 19565 18435
rect 19595 18405 19600 18435
rect 19560 18275 19600 18405
rect 19560 18245 19565 18275
rect 19595 18245 19600 18275
rect 19560 18240 19600 18245
rect 19640 18435 19680 18440
rect 19640 18405 19645 18435
rect 19675 18405 19680 18435
rect 19640 18275 19680 18405
rect 19640 18245 19645 18275
rect 19675 18245 19680 18275
rect 19640 18240 19680 18245
rect 19720 18435 19760 18440
rect 19720 18405 19725 18435
rect 19755 18405 19760 18435
rect 19720 18275 19760 18405
rect 19720 18245 19725 18275
rect 19755 18245 19760 18275
rect 19720 18240 19760 18245
rect 19800 18435 19840 18440
rect 19800 18405 19805 18435
rect 19835 18405 19840 18435
rect 19800 18275 19840 18405
rect 19800 18245 19805 18275
rect 19835 18245 19840 18275
rect 19800 18240 19840 18245
rect 19880 18435 19920 18440
rect 19880 18405 19885 18435
rect 19915 18405 19920 18435
rect 19880 18275 19920 18405
rect 19880 18245 19885 18275
rect 19915 18245 19920 18275
rect 19880 18240 19920 18245
rect 19960 18435 20000 18440
rect 19960 18405 19965 18435
rect 19995 18405 20000 18435
rect 19960 18275 20000 18405
rect 19960 18245 19965 18275
rect 19995 18245 20000 18275
rect 19960 18240 20000 18245
rect 20040 18435 20080 18440
rect 20040 18405 20045 18435
rect 20075 18405 20080 18435
rect 20040 18275 20080 18405
rect 20040 18245 20045 18275
rect 20075 18245 20080 18275
rect 20040 18240 20080 18245
rect 20120 18435 20160 18440
rect 20120 18405 20125 18435
rect 20155 18405 20160 18435
rect 20120 18275 20160 18405
rect 20120 18245 20125 18275
rect 20155 18245 20160 18275
rect 20120 18240 20160 18245
rect 20200 18435 20240 18440
rect 20200 18405 20205 18435
rect 20235 18405 20240 18435
rect 20200 18275 20240 18405
rect 20200 18245 20205 18275
rect 20235 18245 20240 18275
rect 20200 18240 20240 18245
rect 20280 18435 20320 18440
rect 20280 18405 20285 18435
rect 20315 18405 20320 18435
rect 20280 18275 20320 18405
rect 20280 18245 20285 18275
rect 20315 18245 20320 18275
rect 20280 18240 20320 18245
rect 20360 18435 20400 18440
rect 20360 18405 20365 18435
rect 20395 18405 20400 18435
rect 20360 18275 20400 18405
rect 20360 18245 20365 18275
rect 20395 18245 20400 18275
rect 20360 18240 20400 18245
rect 20440 18435 20480 18440
rect 20440 18405 20445 18435
rect 20475 18405 20480 18435
rect 20440 18275 20480 18405
rect 20440 18245 20445 18275
rect 20475 18245 20480 18275
rect 20440 18240 20480 18245
rect 20520 18435 20560 18440
rect 20520 18405 20525 18435
rect 20555 18405 20560 18435
rect 20520 18275 20560 18405
rect 20520 18245 20525 18275
rect 20555 18245 20560 18275
rect 20520 18240 20560 18245
rect 20600 18435 20640 18440
rect 20600 18405 20605 18435
rect 20635 18405 20640 18435
rect 20600 18275 20640 18405
rect 20600 18245 20605 18275
rect 20635 18245 20640 18275
rect 20600 18240 20640 18245
rect 20680 18435 20720 18440
rect 20680 18405 20685 18435
rect 20715 18405 20720 18435
rect 20680 18275 20720 18405
rect 20680 18245 20685 18275
rect 20715 18245 20720 18275
rect 20680 18240 20720 18245
rect 20760 18435 20800 18440
rect 20760 18405 20765 18435
rect 20795 18405 20800 18435
rect 20760 18275 20800 18405
rect 20760 18245 20765 18275
rect 20795 18245 20800 18275
rect 20760 18240 20800 18245
rect 20840 18435 20880 18440
rect 20840 18405 20845 18435
rect 20875 18405 20880 18435
rect 20840 18275 20880 18405
rect 20840 18245 20845 18275
rect 20875 18245 20880 18275
rect 20840 18240 20880 18245
rect 20920 18435 20960 18440
rect 20920 18405 20925 18435
rect 20955 18405 20960 18435
rect 20920 18275 20960 18405
rect 20920 18245 20925 18275
rect 20955 18245 20960 18275
rect 20920 18240 20960 18245
rect 16760 18195 16800 18200
rect 16760 18165 16765 18195
rect 16795 18165 16800 18195
rect 16760 18035 16800 18165
rect 16760 18005 16765 18035
rect 16795 18005 16800 18035
rect 16760 17875 16800 18005
rect 16760 17845 16765 17875
rect 16795 17845 16800 17875
rect 16760 17715 16800 17845
rect 16760 17685 16765 17715
rect 16795 17685 16800 17715
rect 16760 17555 16800 17685
rect 16760 17525 16765 17555
rect 16795 17525 16800 17555
rect 16760 17395 16800 17525
rect 16760 17365 16765 17395
rect 16795 17365 16800 17395
rect 16760 17235 16800 17365
rect 16760 17205 16765 17235
rect 16795 17205 16800 17235
rect 16760 17200 16800 17205
rect 16840 18195 16880 18200
rect 16840 18165 16845 18195
rect 16875 18165 16880 18195
rect 16840 18035 16880 18165
rect 16840 18005 16845 18035
rect 16875 18005 16880 18035
rect 16840 17875 16880 18005
rect 16840 17845 16845 17875
rect 16875 17845 16880 17875
rect 16840 17715 16880 17845
rect 16840 17685 16845 17715
rect 16875 17685 16880 17715
rect 16840 17555 16880 17685
rect 16840 17525 16845 17555
rect 16875 17525 16880 17555
rect 16840 17395 16880 17525
rect 16840 17365 16845 17395
rect 16875 17365 16880 17395
rect 16840 17235 16880 17365
rect 16840 17205 16845 17235
rect 16875 17205 16880 17235
rect 16840 17200 16880 17205
rect 16920 18195 16960 18200
rect 16920 18165 16925 18195
rect 16955 18165 16960 18195
rect 16920 18035 16960 18165
rect 16920 18005 16925 18035
rect 16955 18005 16960 18035
rect 16920 17875 16960 18005
rect 16920 17845 16925 17875
rect 16955 17845 16960 17875
rect 16920 17715 16960 17845
rect 16920 17685 16925 17715
rect 16955 17685 16960 17715
rect 16920 17555 16960 17685
rect 16920 17525 16925 17555
rect 16955 17525 16960 17555
rect 16920 17395 16960 17525
rect 16920 17365 16925 17395
rect 16955 17365 16960 17395
rect 16920 17235 16960 17365
rect 16920 17205 16925 17235
rect 16955 17205 16960 17235
rect 16920 17200 16960 17205
rect 17000 18195 17040 18200
rect 17000 18165 17005 18195
rect 17035 18165 17040 18195
rect 17000 18035 17040 18165
rect 17000 18005 17005 18035
rect 17035 18005 17040 18035
rect 17000 17875 17040 18005
rect 17000 17845 17005 17875
rect 17035 17845 17040 17875
rect 17000 17715 17040 17845
rect 17000 17685 17005 17715
rect 17035 17685 17040 17715
rect 17000 17555 17040 17685
rect 17000 17525 17005 17555
rect 17035 17525 17040 17555
rect 17000 17395 17040 17525
rect 17000 17365 17005 17395
rect 17035 17365 17040 17395
rect 17000 17235 17040 17365
rect 17000 17205 17005 17235
rect 17035 17205 17040 17235
rect 17000 17200 17040 17205
rect 17080 18195 17120 18200
rect 17080 18165 17085 18195
rect 17115 18165 17120 18195
rect 17080 18035 17120 18165
rect 17080 18005 17085 18035
rect 17115 18005 17120 18035
rect 17080 17875 17120 18005
rect 17080 17845 17085 17875
rect 17115 17845 17120 17875
rect 17080 17715 17120 17845
rect 17080 17685 17085 17715
rect 17115 17685 17120 17715
rect 17080 17555 17120 17685
rect 17080 17525 17085 17555
rect 17115 17525 17120 17555
rect 17080 17395 17120 17525
rect 17080 17365 17085 17395
rect 17115 17365 17120 17395
rect 17080 17235 17120 17365
rect 17080 17205 17085 17235
rect 17115 17205 17120 17235
rect 17080 17200 17120 17205
rect 17160 18195 17200 18200
rect 17160 18165 17165 18195
rect 17195 18165 17200 18195
rect 17160 18035 17200 18165
rect 17160 18005 17165 18035
rect 17195 18005 17200 18035
rect 17160 17875 17200 18005
rect 17160 17845 17165 17875
rect 17195 17845 17200 17875
rect 17160 17715 17200 17845
rect 17160 17685 17165 17715
rect 17195 17685 17200 17715
rect 17160 17555 17200 17685
rect 17160 17525 17165 17555
rect 17195 17525 17200 17555
rect 17160 17395 17200 17525
rect 17160 17365 17165 17395
rect 17195 17365 17200 17395
rect 17160 17235 17200 17365
rect 17160 17205 17165 17235
rect 17195 17205 17200 17235
rect 17160 17200 17200 17205
rect 17240 18195 17280 18200
rect 17240 18165 17245 18195
rect 17275 18165 17280 18195
rect 17240 18035 17280 18165
rect 17240 18005 17245 18035
rect 17275 18005 17280 18035
rect 17240 17875 17280 18005
rect 17240 17845 17245 17875
rect 17275 17845 17280 17875
rect 17240 17715 17280 17845
rect 17240 17685 17245 17715
rect 17275 17685 17280 17715
rect 17240 17555 17280 17685
rect 17240 17525 17245 17555
rect 17275 17525 17280 17555
rect 17240 17395 17280 17525
rect 17240 17365 17245 17395
rect 17275 17365 17280 17395
rect 17240 17235 17280 17365
rect 17240 17205 17245 17235
rect 17275 17205 17280 17235
rect 17240 17200 17280 17205
rect 17320 18195 17360 18200
rect 17320 18165 17325 18195
rect 17355 18165 17360 18195
rect 17320 18035 17360 18165
rect 17320 18005 17325 18035
rect 17355 18005 17360 18035
rect 17320 17875 17360 18005
rect 17320 17845 17325 17875
rect 17355 17845 17360 17875
rect 17320 17715 17360 17845
rect 17320 17685 17325 17715
rect 17355 17685 17360 17715
rect 17320 17555 17360 17685
rect 17320 17525 17325 17555
rect 17355 17525 17360 17555
rect 17320 17395 17360 17525
rect 17320 17365 17325 17395
rect 17355 17365 17360 17395
rect 17320 17235 17360 17365
rect 17320 17205 17325 17235
rect 17355 17205 17360 17235
rect 17320 17200 17360 17205
rect 17400 18195 17440 18200
rect 17400 18165 17405 18195
rect 17435 18165 17440 18195
rect 17400 18035 17440 18165
rect 17400 18005 17405 18035
rect 17435 18005 17440 18035
rect 17400 17875 17440 18005
rect 17400 17845 17405 17875
rect 17435 17845 17440 17875
rect 17400 17715 17440 17845
rect 17400 17685 17405 17715
rect 17435 17685 17440 17715
rect 17400 17555 17440 17685
rect 17400 17525 17405 17555
rect 17435 17525 17440 17555
rect 17400 17395 17440 17525
rect 17400 17365 17405 17395
rect 17435 17365 17440 17395
rect 17400 17235 17440 17365
rect 17400 17205 17405 17235
rect 17435 17205 17440 17235
rect 17400 17200 17440 17205
rect 17480 18195 17520 18200
rect 17480 18165 17485 18195
rect 17515 18165 17520 18195
rect 17480 18035 17520 18165
rect 17480 18005 17485 18035
rect 17515 18005 17520 18035
rect 17480 17875 17520 18005
rect 17480 17845 17485 17875
rect 17515 17845 17520 17875
rect 17480 17715 17520 17845
rect 17480 17685 17485 17715
rect 17515 17685 17520 17715
rect 17480 17555 17520 17685
rect 17480 17525 17485 17555
rect 17515 17525 17520 17555
rect 17480 17395 17520 17525
rect 17480 17365 17485 17395
rect 17515 17365 17520 17395
rect 17480 17235 17520 17365
rect 17480 17205 17485 17235
rect 17515 17205 17520 17235
rect 17480 17200 17520 17205
rect 17560 18195 17600 18200
rect 17560 18165 17565 18195
rect 17595 18165 17600 18195
rect 17560 18035 17600 18165
rect 17560 18005 17565 18035
rect 17595 18005 17600 18035
rect 17560 17875 17600 18005
rect 17560 17845 17565 17875
rect 17595 17845 17600 17875
rect 17560 17715 17600 17845
rect 17560 17685 17565 17715
rect 17595 17685 17600 17715
rect 17560 17555 17600 17685
rect 17560 17525 17565 17555
rect 17595 17525 17600 17555
rect 17560 17395 17600 17525
rect 17560 17365 17565 17395
rect 17595 17365 17600 17395
rect 17560 17235 17600 17365
rect 17560 17205 17565 17235
rect 17595 17205 17600 17235
rect 17560 17200 17600 17205
rect 17640 18195 17680 18200
rect 17640 18165 17645 18195
rect 17675 18165 17680 18195
rect 17640 18035 17680 18165
rect 17640 18005 17645 18035
rect 17675 18005 17680 18035
rect 17640 17875 17680 18005
rect 17640 17845 17645 17875
rect 17675 17845 17680 17875
rect 17640 17715 17680 17845
rect 17640 17685 17645 17715
rect 17675 17685 17680 17715
rect 17640 17555 17680 17685
rect 17640 17525 17645 17555
rect 17675 17525 17680 17555
rect 17640 17395 17680 17525
rect 17640 17365 17645 17395
rect 17675 17365 17680 17395
rect 17640 17235 17680 17365
rect 17640 17205 17645 17235
rect 17675 17205 17680 17235
rect 17640 17200 17680 17205
rect 17720 18195 17760 18200
rect 17720 18165 17725 18195
rect 17755 18165 17760 18195
rect 17720 18035 17760 18165
rect 17720 18005 17725 18035
rect 17755 18005 17760 18035
rect 17720 17875 17760 18005
rect 17720 17845 17725 17875
rect 17755 17845 17760 17875
rect 17720 17715 17760 17845
rect 17720 17685 17725 17715
rect 17755 17685 17760 17715
rect 17720 17555 17760 17685
rect 17720 17525 17725 17555
rect 17755 17525 17760 17555
rect 17720 17395 17760 17525
rect 17720 17365 17725 17395
rect 17755 17365 17760 17395
rect 17720 17235 17760 17365
rect 17720 17205 17725 17235
rect 17755 17205 17760 17235
rect 17720 17200 17760 17205
rect 17800 18195 17840 18200
rect 17800 18165 17805 18195
rect 17835 18165 17840 18195
rect 17800 18035 17840 18165
rect 17800 18005 17805 18035
rect 17835 18005 17840 18035
rect 17800 17875 17840 18005
rect 17800 17845 17805 17875
rect 17835 17845 17840 17875
rect 17800 17715 17840 17845
rect 17800 17685 17805 17715
rect 17835 17685 17840 17715
rect 17800 17555 17840 17685
rect 17800 17525 17805 17555
rect 17835 17525 17840 17555
rect 17800 17395 17840 17525
rect 17800 17365 17805 17395
rect 17835 17365 17840 17395
rect 17800 17235 17840 17365
rect 17800 17205 17805 17235
rect 17835 17205 17840 17235
rect 17800 17200 17840 17205
rect 17880 18195 17920 18200
rect 17880 18165 17885 18195
rect 17915 18165 17920 18195
rect 17880 18035 17920 18165
rect 17880 18005 17885 18035
rect 17915 18005 17920 18035
rect 17880 17875 17920 18005
rect 17880 17845 17885 17875
rect 17915 17845 17920 17875
rect 17880 17715 17920 17845
rect 17880 17685 17885 17715
rect 17915 17685 17920 17715
rect 17880 17555 17920 17685
rect 17880 17525 17885 17555
rect 17915 17525 17920 17555
rect 17880 17395 17920 17525
rect 17880 17365 17885 17395
rect 17915 17365 17920 17395
rect 17880 17235 17920 17365
rect 17880 17205 17885 17235
rect 17915 17205 17920 17235
rect 17880 17200 17920 17205
rect 17960 18195 18000 18200
rect 17960 18165 17965 18195
rect 17995 18165 18000 18195
rect 17960 18035 18000 18165
rect 17960 18005 17965 18035
rect 17995 18005 18000 18035
rect 17960 17875 18000 18005
rect 17960 17845 17965 17875
rect 17995 17845 18000 17875
rect 17960 17715 18000 17845
rect 17960 17685 17965 17715
rect 17995 17685 18000 17715
rect 17960 17555 18000 17685
rect 17960 17525 17965 17555
rect 17995 17525 18000 17555
rect 17960 17395 18000 17525
rect 17960 17365 17965 17395
rect 17995 17365 18000 17395
rect 17960 17235 18000 17365
rect 17960 17205 17965 17235
rect 17995 17205 18000 17235
rect 17960 17200 18000 17205
rect 18040 18195 18080 18200
rect 18040 18165 18045 18195
rect 18075 18165 18080 18195
rect 18040 18035 18080 18165
rect 18040 18005 18045 18035
rect 18075 18005 18080 18035
rect 18040 17875 18080 18005
rect 18040 17845 18045 17875
rect 18075 17845 18080 17875
rect 18040 17715 18080 17845
rect 18040 17685 18045 17715
rect 18075 17685 18080 17715
rect 18040 17555 18080 17685
rect 18040 17525 18045 17555
rect 18075 17525 18080 17555
rect 18040 17395 18080 17525
rect 18040 17365 18045 17395
rect 18075 17365 18080 17395
rect 18040 17235 18080 17365
rect 18040 17205 18045 17235
rect 18075 17205 18080 17235
rect 18040 17200 18080 17205
rect 18120 18195 18160 18200
rect 18120 18165 18125 18195
rect 18155 18165 18160 18195
rect 18120 18035 18160 18165
rect 18120 18005 18125 18035
rect 18155 18005 18160 18035
rect 18120 17875 18160 18005
rect 18120 17845 18125 17875
rect 18155 17845 18160 17875
rect 18120 17715 18160 17845
rect 18120 17685 18125 17715
rect 18155 17685 18160 17715
rect 18120 17555 18160 17685
rect 18120 17525 18125 17555
rect 18155 17525 18160 17555
rect 18120 17395 18160 17525
rect 18120 17365 18125 17395
rect 18155 17365 18160 17395
rect 18120 17235 18160 17365
rect 18120 17205 18125 17235
rect 18155 17205 18160 17235
rect 18120 17200 18160 17205
rect 18200 18195 18240 18200
rect 18200 18165 18205 18195
rect 18235 18165 18240 18195
rect 18200 18035 18240 18165
rect 18200 18005 18205 18035
rect 18235 18005 18240 18035
rect 18200 17875 18240 18005
rect 18200 17845 18205 17875
rect 18235 17845 18240 17875
rect 18200 17715 18240 17845
rect 18200 17685 18205 17715
rect 18235 17685 18240 17715
rect 18200 17555 18240 17685
rect 18200 17525 18205 17555
rect 18235 17525 18240 17555
rect 18200 17395 18240 17525
rect 18200 17365 18205 17395
rect 18235 17365 18240 17395
rect 18200 17235 18240 17365
rect 18200 17205 18205 17235
rect 18235 17205 18240 17235
rect 18200 17200 18240 17205
rect 18280 18195 18320 18200
rect 18280 18165 18285 18195
rect 18315 18165 18320 18195
rect 18280 18035 18320 18165
rect 18280 18005 18285 18035
rect 18315 18005 18320 18035
rect 18280 17875 18320 18005
rect 18280 17845 18285 17875
rect 18315 17845 18320 17875
rect 18280 17715 18320 17845
rect 18280 17685 18285 17715
rect 18315 17685 18320 17715
rect 18280 17555 18320 17685
rect 18280 17525 18285 17555
rect 18315 17525 18320 17555
rect 18280 17395 18320 17525
rect 18280 17365 18285 17395
rect 18315 17365 18320 17395
rect 18280 17235 18320 17365
rect 18280 17205 18285 17235
rect 18315 17205 18320 17235
rect 18280 17200 18320 17205
rect 18360 18195 18400 18200
rect 18360 18165 18365 18195
rect 18395 18165 18400 18195
rect 18360 18035 18400 18165
rect 18360 18005 18365 18035
rect 18395 18005 18400 18035
rect 18360 17875 18400 18005
rect 18360 17845 18365 17875
rect 18395 17845 18400 17875
rect 18360 17715 18400 17845
rect 18360 17685 18365 17715
rect 18395 17685 18400 17715
rect 18360 17555 18400 17685
rect 18360 17525 18365 17555
rect 18395 17525 18400 17555
rect 18360 17395 18400 17525
rect 18360 17365 18365 17395
rect 18395 17365 18400 17395
rect 18360 17235 18400 17365
rect 18360 17205 18365 17235
rect 18395 17205 18400 17235
rect 18360 17200 18400 17205
rect 18440 18195 18480 18200
rect 18440 18165 18445 18195
rect 18475 18165 18480 18195
rect 18440 18035 18480 18165
rect 18440 18005 18445 18035
rect 18475 18005 18480 18035
rect 18440 17875 18480 18005
rect 18440 17845 18445 17875
rect 18475 17845 18480 17875
rect 18440 17715 18480 17845
rect 18440 17685 18445 17715
rect 18475 17685 18480 17715
rect 18440 17555 18480 17685
rect 18440 17525 18445 17555
rect 18475 17525 18480 17555
rect 18440 17395 18480 17525
rect 18440 17365 18445 17395
rect 18475 17365 18480 17395
rect 18440 17235 18480 17365
rect 18440 17205 18445 17235
rect 18475 17205 18480 17235
rect 18440 17200 18480 17205
rect 18520 18195 18560 18200
rect 18520 18165 18525 18195
rect 18555 18165 18560 18195
rect 18520 18035 18560 18165
rect 18520 18005 18525 18035
rect 18555 18005 18560 18035
rect 18520 17875 18560 18005
rect 18520 17845 18525 17875
rect 18555 17845 18560 17875
rect 18520 17715 18560 17845
rect 18520 17685 18525 17715
rect 18555 17685 18560 17715
rect 18520 17555 18560 17685
rect 18520 17525 18525 17555
rect 18555 17525 18560 17555
rect 18520 17395 18560 17525
rect 18520 17365 18525 17395
rect 18555 17365 18560 17395
rect 18520 17235 18560 17365
rect 18520 17205 18525 17235
rect 18555 17205 18560 17235
rect 18520 17200 18560 17205
rect 18600 18195 18640 18200
rect 18600 18165 18605 18195
rect 18635 18165 18640 18195
rect 18600 18035 18640 18165
rect 18600 18005 18605 18035
rect 18635 18005 18640 18035
rect 18600 17875 18640 18005
rect 18600 17845 18605 17875
rect 18635 17845 18640 17875
rect 18600 17715 18640 17845
rect 18600 17685 18605 17715
rect 18635 17685 18640 17715
rect 18600 17555 18640 17685
rect 18600 17525 18605 17555
rect 18635 17525 18640 17555
rect 18600 17395 18640 17525
rect 18600 17365 18605 17395
rect 18635 17365 18640 17395
rect 18600 17235 18640 17365
rect 18600 17205 18605 17235
rect 18635 17205 18640 17235
rect 18600 17200 18640 17205
rect 18680 18195 18720 18200
rect 18680 18165 18685 18195
rect 18715 18165 18720 18195
rect 18680 18035 18720 18165
rect 18680 18005 18685 18035
rect 18715 18005 18720 18035
rect 18680 17875 18720 18005
rect 18680 17845 18685 17875
rect 18715 17845 18720 17875
rect 18680 17715 18720 17845
rect 18680 17685 18685 17715
rect 18715 17685 18720 17715
rect 18680 17555 18720 17685
rect 18680 17525 18685 17555
rect 18715 17525 18720 17555
rect 18680 17395 18720 17525
rect 18680 17365 18685 17395
rect 18715 17365 18720 17395
rect 18680 17235 18720 17365
rect 18680 17205 18685 17235
rect 18715 17205 18720 17235
rect 18680 17200 18720 17205
rect 18760 18195 18800 18200
rect 18760 18165 18765 18195
rect 18795 18165 18800 18195
rect 18760 18035 18800 18165
rect 18760 18005 18765 18035
rect 18795 18005 18800 18035
rect 18760 17875 18800 18005
rect 18760 17845 18765 17875
rect 18795 17845 18800 17875
rect 18760 17715 18800 17845
rect 18760 17685 18765 17715
rect 18795 17685 18800 17715
rect 18760 17555 18800 17685
rect 18760 17525 18765 17555
rect 18795 17525 18800 17555
rect 18760 17395 18800 17525
rect 18760 17365 18765 17395
rect 18795 17365 18800 17395
rect 18760 17235 18800 17365
rect 18760 17205 18765 17235
rect 18795 17205 18800 17235
rect 18760 17200 18800 17205
rect 18840 18195 18880 18200
rect 18840 18165 18845 18195
rect 18875 18165 18880 18195
rect 18840 18035 18880 18165
rect 18840 18005 18845 18035
rect 18875 18005 18880 18035
rect 18840 17875 18880 18005
rect 18840 17845 18845 17875
rect 18875 17845 18880 17875
rect 18840 17715 18880 17845
rect 18840 17685 18845 17715
rect 18875 17685 18880 17715
rect 18840 17555 18880 17685
rect 18840 17525 18845 17555
rect 18875 17525 18880 17555
rect 18840 17395 18880 17525
rect 18840 17365 18845 17395
rect 18875 17365 18880 17395
rect 18840 17235 18880 17365
rect 18840 17205 18845 17235
rect 18875 17205 18880 17235
rect 18840 17200 18880 17205
rect 18920 18195 18960 18200
rect 18920 18165 18925 18195
rect 18955 18165 18960 18195
rect 18920 18035 18960 18165
rect 18920 18005 18925 18035
rect 18955 18005 18960 18035
rect 18920 17875 18960 18005
rect 18920 17845 18925 17875
rect 18955 17845 18960 17875
rect 18920 17715 18960 17845
rect 18920 17685 18925 17715
rect 18955 17685 18960 17715
rect 18920 17555 18960 17685
rect 18920 17525 18925 17555
rect 18955 17525 18960 17555
rect 18920 17395 18960 17525
rect 18920 17365 18925 17395
rect 18955 17365 18960 17395
rect 18920 17235 18960 17365
rect 18920 17205 18925 17235
rect 18955 17205 18960 17235
rect 18920 17200 18960 17205
rect 19000 18195 19040 18200
rect 19000 18165 19005 18195
rect 19035 18165 19040 18195
rect 19000 18035 19040 18165
rect 19000 18005 19005 18035
rect 19035 18005 19040 18035
rect 19000 17875 19040 18005
rect 19000 17845 19005 17875
rect 19035 17845 19040 17875
rect 19000 17715 19040 17845
rect 19000 17685 19005 17715
rect 19035 17685 19040 17715
rect 19000 17555 19040 17685
rect 19000 17525 19005 17555
rect 19035 17525 19040 17555
rect 19000 17395 19040 17525
rect 19000 17365 19005 17395
rect 19035 17365 19040 17395
rect 19000 17235 19040 17365
rect 19000 17205 19005 17235
rect 19035 17205 19040 17235
rect 19000 17200 19040 17205
rect 19080 18195 19120 18200
rect 19080 18165 19085 18195
rect 19115 18165 19120 18195
rect 19080 18035 19120 18165
rect 19080 18005 19085 18035
rect 19115 18005 19120 18035
rect 19080 17875 19120 18005
rect 19080 17845 19085 17875
rect 19115 17845 19120 17875
rect 19080 17715 19120 17845
rect 19080 17685 19085 17715
rect 19115 17685 19120 17715
rect 19080 17555 19120 17685
rect 19080 17525 19085 17555
rect 19115 17525 19120 17555
rect 19080 17395 19120 17525
rect 19080 17365 19085 17395
rect 19115 17365 19120 17395
rect 19080 17235 19120 17365
rect 19080 17205 19085 17235
rect 19115 17205 19120 17235
rect 19080 17200 19120 17205
rect 19160 18195 19200 18200
rect 19160 18165 19165 18195
rect 19195 18165 19200 18195
rect 19160 18035 19200 18165
rect 19160 18005 19165 18035
rect 19195 18005 19200 18035
rect 19160 17875 19200 18005
rect 19160 17845 19165 17875
rect 19195 17845 19200 17875
rect 19160 17715 19200 17845
rect 19160 17685 19165 17715
rect 19195 17685 19200 17715
rect 19160 17555 19200 17685
rect 19160 17525 19165 17555
rect 19195 17525 19200 17555
rect 19160 17395 19200 17525
rect 19160 17365 19165 17395
rect 19195 17365 19200 17395
rect 19160 17235 19200 17365
rect 19160 17205 19165 17235
rect 19195 17205 19200 17235
rect 19160 17200 19200 17205
rect 19240 18195 19280 18200
rect 19240 18165 19245 18195
rect 19275 18165 19280 18195
rect 19240 18035 19280 18165
rect 19240 18005 19245 18035
rect 19275 18005 19280 18035
rect 19240 17875 19280 18005
rect 19240 17845 19245 17875
rect 19275 17845 19280 17875
rect 19240 17715 19280 17845
rect 19240 17685 19245 17715
rect 19275 17685 19280 17715
rect 19240 17555 19280 17685
rect 19240 17525 19245 17555
rect 19275 17525 19280 17555
rect 19240 17395 19280 17525
rect 19240 17365 19245 17395
rect 19275 17365 19280 17395
rect 19240 17235 19280 17365
rect 19240 17205 19245 17235
rect 19275 17205 19280 17235
rect 19240 17200 19280 17205
rect 19320 18195 19360 18200
rect 19320 18165 19325 18195
rect 19355 18165 19360 18195
rect 19320 18035 19360 18165
rect 19320 18005 19325 18035
rect 19355 18005 19360 18035
rect 19320 17875 19360 18005
rect 19320 17845 19325 17875
rect 19355 17845 19360 17875
rect 19320 17715 19360 17845
rect 19320 17685 19325 17715
rect 19355 17685 19360 17715
rect 19320 17555 19360 17685
rect 19320 17525 19325 17555
rect 19355 17525 19360 17555
rect 19320 17395 19360 17525
rect 19320 17365 19325 17395
rect 19355 17365 19360 17395
rect 19320 17235 19360 17365
rect 19320 17205 19325 17235
rect 19355 17205 19360 17235
rect 19320 17200 19360 17205
rect 19400 18195 19440 18200
rect 19400 18165 19405 18195
rect 19435 18165 19440 18195
rect 19400 18035 19440 18165
rect 19400 18005 19405 18035
rect 19435 18005 19440 18035
rect 19400 17875 19440 18005
rect 19400 17845 19405 17875
rect 19435 17845 19440 17875
rect 19400 17715 19440 17845
rect 19400 17685 19405 17715
rect 19435 17685 19440 17715
rect 19400 17555 19440 17685
rect 19400 17525 19405 17555
rect 19435 17525 19440 17555
rect 19400 17395 19440 17525
rect 19400 17365 19405 17395
rect 19435 17365 19440 17395
rect 19400 17235 19440 17365
rect 19400 17205 19405 17235
rect 19435 17205 19440 17235
rect 19400 17200 19440 17205
rect 19480 18195 19520 18200
rect 19480 18165 19485 18195
rect 19515 18165 19520 18195
rect 19480 18035 19520 18165
rect 19480 18005 19485 18035
rect 19515 18005 19520 18035
rect 19480 17875 19520 18005
rect 19480 17845 19485 17875
rect 19515 17845 19520 17875
rect 19480 17715 19520 17845
rect 19480 17685 19485 17715
rect 19515 17685 19520 17715
rect 19480 17555 19520 17685
rect 19480 17525 19485 17555
rect 19515 17525 19520 17555
rect 19480 17395 19520 17525
rect 19480 17365 19485 17395
rect 19515 17365 19520 17395
rect 19480 17235 19520 17365
rect 19480 17205 19485 17235
rect 19515 17205 19520 17235
rect 19480 17200 19520 17205
rect 19560 18195 19600 18200
rect 19560 18165 19565 18195
rect 19595 18165 19600 18195
rect 19560 18035 19600 18165
rect 19560 18005 19565 18035
rect 19595 18005 19600 18035
rect 19560 17875 19600 18005
rect 19560 17845 19565 17875
rect 19595 17845 19600 17875
rect 19560 17715 19600 17845
rect 19560 17685 19565 17715
rect 19595 17685 19600 17715
rect 19560 17555 19600 17685
rect 19560 17525 19565 17555
rect 19595 17525 19600 17555
rect 19560 17395 19600 17525
rect 19560 17365 19565 17395
rect 19595 17365 19600 17395
rect 19560 17235 19600 17365
rect 19560 17205 19565 17235
rect 19595 17205 19600 17235
rect 19560 17200 19600 17205
rect 19640 18195 19680 18200
rect 19640 18165 19645 18195
rect 19675 18165 19680 18195
rect 19640 18035 19680 18165
rect 19640 18005 19645 18035
rect 19675 18005 19680 18035
rect 19640 17875 19680 18005
rect 19640 17845 19645 17875
rect 19675 17845 19680 17875
rect 19640 17715 19680 17845
rect 19640 17685 19645 17715
rect 19675 17685 19680 17715
rect 19640 17555 19680 17685
rect 19640 17525 19645 17555
rect 19675 17525 19680 17555
rect 19640 17395 19680 17525
rect 19640 17365 19645 17395
rect 19675 17365 19680 17395
rect 19640 17235 19680 17365
rect 19640 17205 19645 17235
rect 19675 17205 19680 17235
rect 19640 17200 19680 17205
rect 19720 18195 19760 18200
rect 19720 18165 19725 18195
rect 19755 18165 19760 18195
rect 19720 18035 19760 18165
rect 19720 18005 19725 18035
rect 19755 18005 19760 18035
rect 19720 17875 19760 18005
rect 19720 17845 19725 17875
rect 19755 17845 19760 17875
rect 19720 17715 19760 17845
rect 19720 17685 19725 17715
rect 19755 17685 19760 17715
rect 19720 17555 19760 17685
rect 19720 17525 19725 17555
rect 19755 17525 19760 17555
rect 19720 17395 19760 17525
rect 19720 17365 19725 17395
rect 19755 17365 19760 17395
rect 19720 17235 19760 17365
rect 19720 17205 19725 17235
rect 19755 17205 19760 17235
rect 19720 17200 19760 17205
rect 19800 18195 19840 18200
rect 19800 18165 19805 18195
rect 19835 18165 19840 18195
rect 19800 18035 19840 18165
rect 19800 18005 19805 18035
rect 19835 18005 19840 18035
rect 19800 17875 19840 18005
rect 19800 17845 19805 17875
rect 19835 17845 19840 17875
rect 19800 17715 19840 17845
rect 19800 17685 19805 17715
rect 19835 17685 19840 17715
rect 19800 17555 19840 17685
rect 19800 17525 19805 17555
rect 19835 17525 19840 17555
rect 19800 17395 19840 17525
rect 19800 17365 19805 17395
rect 19835 17365 19840 17395
rect 19800 17235 19840 17365
rect 19800 17205 19805 17235
rect 19835 17205 19840 17235
rect 19800 17200 19840 17205
rect 19880 18195 19920 18200
rect 19880 18165 19885 18195
rect 19915 18165 19920 18195
rect 19880 18035 19920 18165
rect 19880 18005 19885 18035
rect 19915 18005 19920 18035
rect 19880 17875 19920 18005
rect 19880 17845 19885 17875
rect 19915 17845 19920 17875
rect 19880 17715 19920 17845
rect 19880 17685 19885 17715
rect 19915 17685 19920 17715
rect 19880 17555 19920 17685
rect 19880 17525 19885 17555
rect 19915 17525 19920 17555
rect 19880 17395 19920 17525
rect 19880 17365 19885 17395
rect 19915 17365 19920 17395
rect 19880 17235 19920 17365
rect 19880 17205 19885 17235
rect 19915 17205 19920 17235
rect 19880 17200 19920 17205
rect 19960 18195 20000 18200
rect 19960 18165 19965 18195
rect 19995 18165 20000 18195
rect 19960 18035 20000 18165
rect 19960 18005 19965 18035
rect 19995 18005 20000 18035
rect 19960 17875 20000 18005
rect 19960 17845 19965 17875
rect 19995 17845 20000 17875
rect 19960 17715 20000 17845
rect 19960 17685 19965 17715
rect 19995 17685 20000 17715
rect 19960 17555 20000 17685
rect 19960 17525 19965 17555
rect 19995 17525 20000 17555
rect 19960 17395 20000 17525
rect 19960 17365 19965 17395
rect 19995 17365 20000 17395
rect 19960 17235 20000 17365
rect 19960 17205 19965 17235
rect 19995 17205 20000 17235
rect 19960 17200 20000 17205
rect 20040 18195 20080 18200
rect 20040 18165 20045 18195
rect 20075 18165 20080 18195
rect 20040 18035 20080 18165
rect 20040 18005 20045 18035
rect 20075 18005 20080 18035
rect 20040 17875 20080 18005
rect 20040 17845 20045 17875
rect 20075 17845 20080 17875
rect 20040 17715 20080 17845
rect 20040 17685 20045 17715
rect 20075 17685 20080 17715
rect 20040 17555 20080 17685
rect 20040 17525 20045 17555
rect 20075 17525 20080 17555
rect 20040 17395 20080 17525
rect 20040 17365 20045 17395
rect 20075 17365 20080 17395
rect 20040 17235 20080 17365
rect 20040 17205 20045 17235
rect 20075 17205 20080 17235
rect 20040 17200 20080 17205
rect 20120 18195 20160 18200
rect 20120 18165 20125 18195
rect 20155 18165 20160 18195
rect 20120 18035 20160 18165
rect 20120 18005 20125 18035
rect 20155 18005 20160 18035
rect 20120 17875 20160 18005
rect 20120 17845 20125 17875
rect 20155 17845 20160 17875
rect 20120 17715 20160 17845
rect 20120 17685 20125 17715
rect 20155 17685 20160 17715
rect 20120 17555 20160 17685
rect 20120 17525 20125 17555
rect 20155 17525 20160 17555
rect 20120 17395 20160 17525
rect 20120 17365 20125 17395
rect 20155 17365 20160 17395
rect 20120 17235 20160 17365
rect 20120 17205 20125 17235
rect 20155 17205 20160 17235
rect 20120 17200 20160 17205
rect 20200 18195 20240 18200
rect 20200 18165 20205 18195
rect 20235 18165 20240 18195
rect 20200 18035 20240 18165
rect 20200 18005 20205 18035
rect 20235 18005 20240 18035
rect 20200 17875 20240 18005
rect 20200 17845 20205 17875
rect 20235 17845 20240 17875
rect 20200 17715 20240 17845
rect 20200 17685 20205 17715
rect 20235 17685 20240 17715
rect 20200 17555 20240 17685
rect 20200 17525 20205 17555
rect 20235 17525 20240 17555
rect 20200 17395 20240 17525
rect 20200 17365 20205 17395
rect 20235 17365 20240 17395
rect 20200 17235 20240 17365
rect 20200 17205 20205 17235
rect 20235 17205 20240 17235
rect 20200 17200 20240 17205
rect 20280 18195 20320 18200
rect 20280 18165 20285 18195
rect 20315 18165 20320 18195
rect 20280 18035 20320 18165
rect 20280 18005 20285 18035
rect 20315 18005 20320 18035
rect 20280 17875 20320 18005
rect 20280 17845 20285 17875
rect 20315 17845 20320 17875
rect 20280 17715 20320 17845
rect 20280 17685 20285 17715
rect 20315 17685 20320 17715
rect 20280 17555 20320 17685
rect 20280 17525 20285 17555
rect 20315 17525 20320 17555
rect 20280 17395 20320 17525
rect 20280 17365 20285 17395
rect 20315 17365 20320 17395
rect 20280 17235 20320 17365
rect 20280 17205 20285 17235
rect 20315 17205 20320 17235
rect 20280 17200 20320 17205
rect 20360 18195 20400 18200
rect 20360 18165 20365 18195
rect 20395 18165 20400 18195
rect 20360 18035 20400 18165
rect 20360 18005 20365 18035
rect 20395 18005 20400 18035
rect 20360 17875 20400 18005
rect 20360 17845 20365 17875
rect 20395 17845 20400 17875
rect 20360 17715 20400 17845
rect 20360 17685 20365 17715
rect 20395 17685 20400 17715
rect 20360 17555 20400 17685
rect 20360 17525 20365 17555
rect 20395 17525 20400 17555
rect 20360 17395 20400 17525
rect 20360 17365 20365 17395
rect 20395 17365 20400 17395
rect 20360 17235 20400 17365
rect 20360 17205 20365 17235
rect 20395 17205 20400 17235
rect 20360 17200 20400 17205
rect 20440 18195 20480 18200
rect 20440 18165 20445 18195
rect 20475 18165 20480 18195
rect 20440 18035 20480 18165
rect 20440 18005 20445 18035
rect 20475 18005 20480 18035
rect 20440 17875 20480 18005
rect 20440 17845 20445 17875
rect 20475 17845 20480 17875
rect 20440 17715 20480 17845
rect 20440 17685 20445 17715
rect 20475 17685 20480 17715
rect 20440 17555 20480 17685
rect 20440 17525 20445 17555
rect 20475 17525 20480 17555
rect 20440 17395 20480 17525
rect 20440 17365 20445 17395
rect 20475 17365 20480 17395
rect 20440 17235 20480 17365
rect 20440 17205 20445 17235
rect 20475 17205 20480 17235
rect 20440 17200 20480 17205
rect 20520 18195 20560 18200
rect 20520 18165 20525 18195
rect 20555 18165 20560 18195
rect 20520 18035 20560 18165
rect 20520 18005 20525 18035
rect 20555 18005 20560 18035
rect 20520 17875 20560 18005
rect 20520 17845 20525 17875
rect 20555 17845 20560 17875
rect 20520 17715 20560 17845
rect 20520 17685 20525 17715
rect 20555 17685 20560 17715
rect 20520 17555 20560 17685
rect 20520 17525 20525 17555
rect 20555 17525 20560 17555
rect 20520 17395 20560 17525
rect 20520 17365 20525 17395
rect 20555 17365 20560 17395
rect 20520 17235 20560 17365
rect 20520 17205 20525 17235
rect 20555 17205 20560 17235
rect 20520 17200 20560 17205
rect 20600 18195 20640 18200
rect 20600 18165 20605 18195
rect 20635 18165 20640 18195
rect 20600 18035 20640 18165
rect 20600 18005 20605 18035
rect 20635 18005 20640 18035
rect 20600 17875 20640 18005
rect 20600 17845 20605 17875
rect 20635 17845 20640 17875
rect 20600 17715 20640 17845
rect 20600 17685 20605 17715
rect 20635 17685 20640 17715
rect 20600 17555 20640 17685
rect 20600 17525 20605 17555
rect 20635 17525 20640 17555
rect 20600 17395 20640 17525
rect 20600 17365 20605 17395
rect 20635 17365 20640 17395
rect 20600 17235 20640 17365
rect 20600 17205 20605 17235
rect 20635 17205 20640 17235
rect 20600 17200 20640 17205
rect 20680 18195 20720 18200
rect 20680 18165 20685 18195
rect 20715 18165 20720 18195
rect 20680 18035 20720 18165
rect 20680 18005 20685 18035
rect 20715 18005 20720 18035
rect 20680 17875 20720 18005
rect 20680 17845 20685 17875
rect 20715 17845 20720 17875
rect 20680 17715 20720 17845
rect 20680 17685 20685 17715
rect 20715 17685 20720 17715
rect 20680 17555 20720 17685
rect 20680 17525 20685 17555
rect 20715 17525 20720 17555
rect 20680 17395 20720 17525
rect 20680 17365 20685 17395
rect 20715 17365 20720 17395
rect 20680 17235 20720 17365
rect 20680 17205 20685 17235
rect 20715 17205 20720 17235
rect 20680 17200 20720 17205
rect 20760 18195 20800 18200
rect 20760 18165 20765 18195
rect 20795 18165 20800 18195
rect 20760 18035 20800 18165
rect 20760 18005 20765 18035
rect 20795 18005 20800 18035
rect 20760 17875 20800 18005
rect 20760 17845 20765 17875
rect 20795 17845 20800 17875
rect 20760 17715 20800 17845
rect 20760 17685 20765 17715
rect 20795 17685 20800 17715
rect 20760 17555 20800 17685
rect 20760 17525 20765 17555
rect 20795 17525 20800 17555
rect 20760 17395 20800 17525
rect 20760 17365 20765 17395
rect 20795 17365 20800 17395
rect 20760 17235 20800 17365
rect 20760 17205 20765 17235
rect 20795 17205 20800 17235
rect 20760 17200 20800 17205
rect 20840 18195 20880 18200
rect 20840 18165 20845 18195
rect 20875 18165 20880 18195
rect 20840 18035 20880 18165
rect 20840 18005 20845 18035
rect 20875 18005 20880 18035
rect 20840 17875 20880 18005
rect 20840 17845 20845 17875
rect 20875 17845 20880 17875
rect 20840 17715 20880 17845
rect 20840 17685 20845 17715
rect 20875 17685 20880 17715
rect 20840 17555 20880 17685
rect 20840 17525 20845 17555
rect 20875 17525 20880 17555
rect 20840 17395 20880 17525
rect 20840 17365 20845 17395
rect 20875 17365 20880 17395
rect 20840 17235 20880 17365
rect 20840 17205 20845 17235
rect 20875 17205 20880 17235
rect 20840 17200 20880 17205
rect 20920 18195 20960 18200
rect 20920 18165 20925 18195
rect 20955 18165 20960 18195
rect 20920 18035 20960 18165
rect 20920 18005 20925 18035
rect 20955 18005 20960 18035
rect 20920 17875 20960 18005
rect 20920 17845 20925 17875
rect 20955 17845 20960 17875
rect 20920 17715 20960 17845
rect 20920 17685 20925 17715
rect 20955 17685 20960 17715
rect 20920 17555 20960 17685
rect 20920 17525 20925 17555
rect 20955 17525 20960 17555
rect 20920 17395 20960 17525
rect 20920 17365 20925 17395
rect 20955 17365 20960 17395
rect 20920 17235 20960 17365
rect 20920 17205 20925 17235
rect 20955 17205 20960 17235
rect 20920 17200 20960 17205
rect 16760 17155 16800 17160
rect 16760 17125 16765 17155
rect 16795 17125 16800 17155
rect 16760 16995 16800 17125
rect 16760 16965 16765 16995
rect 16795 16965 16800 16995
rect 16760 16960 16800 16965
rect 16840 17155 16880 17160
rect 16840 17125 16845 17155
rect 16875 17125 16880 17155
rect 16840 16995 16880 17125
rect 16840 16965 16845 16995
rect 16875 16965 16880 16995
rect 16840 16960 16880 16965
rect 16920 17155 16960 17160
rect 16920 17125 16925 17155
rect 16955 17125 16960 17155
rect 16920 16995 16960 17125
rect 16920 16965 16925 16995
rect 16955 16965 16960 16995
rect 16920 16960 16960 16965
rect 17000 17155 17040 17160
rect 17000 17125 17005 17155
rect 17035 17125 17040 17155
rect 17000 16995 17040 17125
rect 17000 16965 17005 16995
rect 17035 16965 17040 16995
rect 17000 16960 17040 16965
rect 17080 17155 17120 17160
rect 17080 17125 17085 17155
rect 17115 17125 17120 17155
rect 17080 16995 17120 17125
rect 17080 16965 17085 16995
rect 17115 16965 17120 16995
rect 17080 16960 17120 16965
rect 17160 17155 17200 17160
rect 17160 17125 17165 17155
rect 17195 17125 17200 17155
rect 17160 16995 17200 17125
rect 17160 16965 17165 16995
rect 17195 16965 17200 16995
rect 17160 16960 17200 16965
rect 17240 17155 17280 17160
rect 17240 17125 17245 17155
rect 17275 17125 17280 17155
rect 17240 16995 17280 17125
rect 17240 16965 17245 16995
rect 17275 16965 17280 16995
rect 17240 16960 17280 16965
rect 17320 17155 17360 17160
rect 17320 17125 17325 17155
rect 17355 17125 17360 17155
rect 17320 16995 17360 17125
rect 17320 16965 17325 16995
rect 17355 16965 17360 16995
rect 17320 16960 17360 16965
rect 17400 17155 17440 17160
rect 17400 17125 17405 17155
rect 17435 17125 17440 17155
rect 17400 16995 17440 17125
rect 17400 16965 17405 16995
rect 17435 16965 17440 16995
rect 17400 16960 17440 16965
rect 17480 17155 17520 17160
rect 17480 17125 17485 17155
rect 17515 17125 17520 17155
rect 17480 16995 17520 17125
rect 17480 16965 17485 16995
rect 17515 16965 17520 16995
rect 17480 16960 17520 16965
rect 17560 17155 17600 17160
rect 17560 17125 17565 17155
rect 17595 17125 17600 17155
rect 17560 16995 17600 17125
rect 17560 16965 17565 16995
rect 17595 16965 17600 16995
rect 17560 16960 17600 16965
rect 17640 17155 17680 17160
rect 17640 17125 17645 17155
rect 17675 17125 17680 17155
rect 17640 16995 17680 17125
rect 17640 16965 17645 16995
rect 17675 16965 17680 16995
rect 17640 16960 17680 16965
rect 17720 17155 17760 17160
rect 17720 17125 17725 17155
rect 17755 17125 17760 17155
rect 17720 16995 17760 17125
rect 17720 16965 17725 16995
rect 17755 16965 17760 16995
rect 17720 16960 17760 16965
rect 17800 17155 17840 17160
rect 17800 17125 17805 17155
rect 17835 17125 17840 17155
rect 17800 16995 17840 17125
rect 17800 16965 17805 16995
rect 17835 16965 17840 16995
rect 17800 16960 17840 16965
rect 17880 17155 17920 17160
rect 17880 17125 17885 17155
rect 17915 17125 17920 17155
rect 17880 16995 17920 17125
rect 17880 16965 17885 16995
rect 17915 16965 17920 16995
rect 17880 16960 17920 16965
rect 17960 17155 18000 17160
rect 17960 17125 17965 17155
rect 17995 17125 18000 17155
rect 17960 16995 18000 17125
rect 17960 16965 17965 16995
rect 17995 16965 18000 16995
rect 17960 16960 18000 16965
rect 18040 17155 18080 17160
rect 18040 17125 18045 17155
rect 18075 17125 18080 17155
rect 18040 16995 18080 17125
rect 18040 16965 18045 16995
rect 18075 16965 18080 16995
rect 18040 16960 18080 16965
rect 18120 17155 18160 17160
rect 18120 17125 18125 17155
rect 18155 17125 18160 17155
rect 18120 16995 18160 17125
rect 18120 16965 18125 16995
rect 18155 16965 18160 16995
rect 18120 16960 18160 16965
rect 18200 17155 18240 17160
rect 18200 17125 18205 17155
rect 18235 17125 18240 17155
rect 18200 16995 18240 17125
rect 18200 16965 18205 16995
rect 18235 16965 18240 16995
rect 18200 16960 18240 16965
rect 18280 17155 18320 17160
rect 18280 17125 18285 17155
rect 18315 17125 18320 17155
rect 18280 16995 18320 17125
rect 18280 16965 18285 16995
rect 18315 16965 18320 16995
rect 18280 16960 18320 16965
rect 18360 17155 18400 17160
rect 18360 17125 18365 17155
rect 18395 17125 18400 17155
rect 18360 16995 18400 17125
rect 18360 16965 18365 16995
rect 18395 16965 18400 16995
rect 18360 16960 18400 16965
rect 18440 17155 18480 17160
rect 18440 17125 18445 17155
rect 18475 17125 18480 17155
rect 18440 16995 18480 17125
rect 18440 16965 18445 16995
rect 18475 16965 18480 16995
rect 18440 16960 18480 16965
rect 18520 17155 18560 17160
rect 18520 17125 18525 17155
rect 18555 17125 18560 17155
rect 18520 16995 18560 17125
rect 18520 16965 18525 16995
rect 18555 16965 18560 16995
rect 18520 16960 18560 16965
rect 18600 17155 18640 17160
rect 18600 17125 18605 17155
rect 18635 17125 18640 17155
rect 18600 16995 18640 17125
rect 18600 16965 18605 16995
rect 18635 16965 18640 16995
rect 18600 16960 18640 16965
rect 18680 17155 18720 17160
rect 18680 17125 18685 17155
rect 18715 17125 18720 17155
rect 18680 16995 18720 17125
rect 18680 16965 18685 16995
rect 18715 16965 18720 16995
rect 18680 16960 18720 16965
rect 18760 17155 18800 17160
rect 18760 17125 18765 17155
rect 18795 17125 18800 17155
rect 18760 16995 18800 17125
rect 18760 16965 18765 16995
rect 18795 16965 18800 16995
rect 18760 16960 18800 16965
rect 18840 17155 18880 17160
rect 18840 17125 18845 17155
rect 18875 17125 18880 17155
rect 18840 16995 18880 17125
rect 18840 16965 18845 16995
rect 18875 16965 18880 16995
rect 18840 16960 18880 16965
rect 18920 17155 18960 17160
rect 18920 17125 18925 17155
rect 18955 17125 18960 17155
rect 18920 16995 18960 17125
rect 18920 16965 18925 16995
rect 18955 16965 18960 16995
rect 18920 16960 18960 16965
rect 19000 17155 19040 17160
rect 19000 17125 19005 17155
rect 19035 17125 19040 17155
rect 19000 16995 19040 17125
rect 19000 16965 19005 16995
rect 19035 16965 19040 16995
rect 19000 16960 19040 16965
rect 19080 17155 19120 17160
rect 19080 17125 19085 17155
rect 19115 17125 19120 17155
rect 19080 16995 19120 17125
rect 19080 16965 19085 16995
rect 19115 16965 19120 16995
rect 19080 16960 19120 16965
rect 19160 17155 19200 17160
rect 19160 17125 19165 17155
rect 19195 17125 19200 17155
rect 19160 16995 19200 17125
rect 19160 16965 19165 16995
rect 19195 16965 19200 16995
rect 19160 16960 19200 16965
rect 19240 17155 19280 17160
rect 19240 17125 19245 17155
rect 19275 17125 19280 17155
rect 19240 16995 19280 17125
rect 19240 16965 19245 16995
rect 19275 16965 19280 16995
rect 19240 16960 19280 16965
rect 19320 17155 19360 17160
rect 19320 17125 19325 17155
rect 19355 17125 19360 17155
rect 19320 16995 19360 17125
rect 19320 16965 19325 16995
rect 19355 16965 19360 16995
rect 19320 16960 19360 16965
rect 19400 17155 19440 17160
rect 19400 17125 19405 17155
rect 19435 17125 19440 17155
rect 19400 16995 19440 17125
rect 19400 16965 19405 16995
rect 19435 16965 19440 16995
rect 19400 16960 19440 16965
rect 19480 17155 19520 17160
rect 19480 17125 19485 17155
rect 19515 17125 19520 17155
rect 19480 16995 19520 17125
rect 19480 16965 19485 16995
rect 19515 16965 19520 16995
rect 19480 16960 19520 16965
rect 19560 17155 19600 17160
rect 19560 17125 19565 17155
rect 19595 17125 19600 17155
rect 19560 16995 19600 17125
rect 19560 16965 19565 16995
rect 19595 16965 19600 16995
rect 19560 16960 19600 16965
rect 19640 17155 19680 17160
rect 19640 17125 19645 17155
rect 19675 17125 19680 17155
rect 19640 16995 19680 17125
rect 19640 16965 19645 16995
rect 19675 16965 19680 16995
rect 19640 16960 19680 16965
rect 19720 17155 19760 17160
rect 19720 17125 19725 17155
rect 19755 17125 19760 17155
rect 19720 16995 19760 17125
rect 19720 16965 19725 16995
rect 19755 16965 19760 16995
rect 19720 16960 19760 16965
rect 19800 17155 19840 17160
rect 19800 17125 19805 17155
rect 19835 17125 19840 17155
rect 19800 16995 19840 17125
rect 19800 16965 19805 16995
rect 19835 16965 19840 16995
rect 19800 16960 19840 16965
rect 19880 17155 19920 17160
rect 19880 17125 19885 17155
rect 19915 17125 19920 17155
rect 19880 16995 19920 17125
rect 19880 16965 19885 16995
rect 19915 16965 19920 16995
rect 19880 16960 19920 16965
rect 19960 17155 20000 17160
rect 19960 17125 19965 17155
rect 19995 17125 20000 17155
rect 19960 16995 20000 17125
rect 19960 16965 19965 16995
rect 19995 16965 20000 16995
rect 19960 16960 20000 16965
rect 20040 17155 20080 17160
rect 20040 17125 20045 17155
rect 20075 17125 20080 17155
rect 20040 16995 20080 17125
rect 20040 16965 20045 16995
rect 20075 16965 20080 16995
rect 20040 16960 20080 16965
rect 20120 17155 20160 17160
rect 20120 17125 20125 17155
rect 20155 17125 20160 17155
rect 20120 16995 20160 17125
rect 20120 16965 20125 16995
rect 20155 16965 20160 16995
rect 20120 16960 20160 16965
rect 20200 17155 20240 17160
rect 20200 17125 20205 17155
rect 20235 17125 20240 17155
rect 20200 16995 20240 17125
rect 20200 16965 20205 16995
rect 20235 16965 20240 16995
rect 20200 16960 20240 16965
rect 20280 17155 20320 17160
rect 20280 17125 20285 17155
rect 20315 17125 20320 17155
rect 20280 16995 20320 17125
rect 20280 16965 20285 16995
rect 20315 16965 20320 16995
rect 20280 16960 20320 16965
rect 20360 17155 20400 17160
rect 20360 17125 20365 17155
rect 20395 17125 20400 17155
rect 20360 16995 20400 17125
rect 20360 16965 20365 16995
rect 20395 16965 20400 16995
rect 20360 16960 20400 16965
rect 20440 17155 20480 17160
rect 20440 17125 20445 17155
rect 20475 17125 20480 17155
rect 20440 16995 20480 17125
rect 20440 16965 20445 16995
rect 20475 16965 20480 16995
rect 20440 16960 20480 16965
rect 20520 17155 20560 17160
rect 20520 17125 20525 17155
rect 20555 17125 20560 17155
rect 20520 16995 20560 17125
rect 20520 16965 20525 16995
rect 20555 16965 20560 16995
rect 20520 16960 20560 16965
rect 20600 17155 20640 17160
rect 20600 17125 20605 17155
rect 20635 17125 20640 17155
rect 20600 16995 20640 17125
rect 20600 16965 20605 16995
rect 20635 16965 20640 16995
rect 20600 16960 20640 16965
rect 20680 17155 20720 17160
rect 20680 17125 20685 17155
rect 20715 17125 20720 17155
rect 20680 16995 20720 17125
rect 20680 16965 20685 16995
rect 20715 16965 20720 16995
rect 20680 16960 20720 16965
rect 20760 17155 20800 17160
rect 20760 17125 20765 17155
rect 20795 17125 20800 17155
rect 20760 16995 20800 17125
rect 20760 16965 20765 16995
rect 20795 16965 20800 16995
rect 20760 16960 20800 16965
rect 20840 17155 20880 17160
rect 20840 17125 20845 17155
rect 20875 17125 20880 17155
rect 20840 16995 20880 17125
rect 20840 16965 20845 16995
rect 20875 16965 20880 16995
rect 20840 16960 20880 16965
rect 20920 17155 20960 17160
rect 20920 17125 20925 17155
rect 20955 17125 20960 17155
rect 20920 16995 20960 17125
rect 20920 16965 20925 16995
rect 20955 16965 20960 16995
rect 20920 16960 20960 16965
rect 16760 16915 16800 16920
rect 16760 16885 16765 16915
rect 16795 16885 16800 16915
rect 16760 16755 16800 16885
rect 16760 16725 16765 16755
rect 16795 16725 16800 16755
rect 16760 16720 16800 16725
rect 16840 16915 16880 16920
rect 16840 16885 16845 16915
rect 16875 16885 16880 16915
rect 16840 16755 16880 16885
rect 16840 16725 16845 16755
rect 16875 16725 16880 16755
rect 16840 16720 16880 16725
rect 16920 16915 16960 16920
rect 16920 16885 16925 16915
rect 16955 16885 16960 16915
rect 16920 16755 16960 16885
rect 16920 16725 16925 16755
rect 16955 16725 16960 16755
rect 16920 16720 16960 16725
rect 17000 16915 17040 16920
rect 17000 16885 17005 16915
rect 17035 16885 17040 16915
rect 17000 16755 17040 16885
rect 17000 16725 17005 16755
rect 17035 16725 17040 16755
rect 17000 16720 17040 16725
rect 17080 16915 17120 16920
rect 17080 16885 17085 16915
rect 17115 16885 17120 16915
rect 17080 16755 17120 16885
rect 17080 16725 17085 16755
rect 17115 16725 17120 16755
rect 17080 16720 17120 16725
rect 17160 16915 17200 16920
rect 17160 16885 17165 16915
rect 17195 16885 17200 16915
rect 17160 16755 17200 16885
rect 17160 16725 17165 16755
rect 17195 16725 17200 16755
rect 17160 16720 17200 16725
rect 17240 16915 17280 16920
rect 17240 16885 17245 16915
rect 17275 16885 17280 16915
rect 17240 16755 17280 16885
rect 17240 16725 17245 16755
rect 17275 16725 17280 16755
rect 17240 16720 17280 16725
rect 17320 16915 17360 16920
rect 17320 16885 17325 16915
rect 17355 16885 17360 16915
rect 17320 16755 17360 16885
rect 17320 16725 17325 16755
rect 17355 16725 17360 16755
rect 17320 16720 17360 16725
rect 17400 16915 17440 16920
rect 17400 16885 17405 16915
rect 17435 16885 17440 16915
rect 17400 16755 17440 16885
rect 17400 16725 17405 16755
rect 17435 16725 17440 16755
rect 17400 16720 17440 16725
rect 17480 16915 17520 16920
rect 17480 16885 17485 16915
rect 17515 16885 17520 16915
rect 17480 16755 17520 16885
rect 17480 16725 17485 16755
rect 17515 16725 17520 16755
rect 17480 16720 17520 16725
rect 17560 16915 17600 16920
rect 17560 16885 17565 16915
rect 17595 16885 17600 16915
rect 17560 16755 17600 16885
rect 17560 16725 17565 16755
rect 17595 16725 17600 16755
rect 17560 16720 17600 16725
rect 17640 16915 17680 16920
rect 17640 16885 17645 16915
rect 17675 16885 17680 16915
rect 17640 16755 17680 16885
rect 17640 16725 17645 16755
rect 17675 16725 17680 16755
rect 17640 16720 17680 16725
rect 17720 16915 17760 16920
rect 17720 16885 17725 16915
rect 17755 16885 17760 16915
rect 17720 16755 17760 16885
rect 17720 16725 17725 16755
rect 17755 16725 17760 16755
rect 17720 16720 17760 16725
rect 17800 16915 17840 16920
rect 17800 16885 17805 16915
rect 17835 16885 17840 16915
rect 17800 16755 17840 16885
rect 17800 16725 17805 16755
rect 17835 16725 17840 16755
rect 17800 16720 17840 16725
rect 17880 16915 17920 16920
rect 17880 16885 17885 16915
rect 17915 16885 17920 16915
rect 17880 16755 17920 16885
rect 17880 16725 17885 16755
rect 17915 16725 17920 16755
rect 17880 16720 17920 16725
rect 17960 16915 18000 16920
rect 17960 16885 17965 16915
rect 17995 16885 18000 16915
rect 17960 16755 18000 16885
rect 17960 16725 17965 16755
rect 17995 16725 18000 16755
rect 17960 16720 18000 16725
rect 18040 16915 18080 16920
rect 18040 16885 18045 16915
rect 18075 16885 18080 16915
rect 18040 16755 18080 16885
rect 18040 16725 18045 16755
rect 18075 16725 18080 16755
rect 18040 16720 18080 16725
rect 18120 16915 18160 16920
rect 18120 16885 18125 16915
rect 18155 16885 18160 16915
rect 18120 16755 18160 16885
rect 18120 16725 18125 16755
rect 18155 16725 18160 16755
rect 18120 16720 18160 16725
rect 18200 16915 18240 16920
rect 18200 16885 18205 16915
rect 18235 16885 18240 16915
rect 18200 16755 18240 16885
rect 18200 16725 18205 16755
rect 18235 16725 18240 16755
rect 18200 16720 18240 16725
rect 18280 16915 18320 16920
rect 18280 16885 18285 16915
rect 18315 16885 18320 16915
rect 18280 16755 18320 16885
rect 18280 16725 18285 16755
rect 18315 16725 18320 16755
rect 18280 16720 18320 16725
rect 18360 16915 18400 16920
rect 18360 16885 18365 16915
rect 18395 16885 18400 16915
rect 18360 16755 18400 16885
rect 18360 16725 18365 16755
rect 18395 16725 18400 16755
rect 18360 16720 18400 16725
rect 18440 16915 18480 16920
rect 18440 16885 18445 16915
rect 18475 16885 18480 16915
rect 18440 16755 18480 16885
rect 18440 16725 18445 16755
rect 18475 16725 18480 16755
rect 18440 16720 18480 16725
rect 18520 16915 18560 16920
rect 18520 16885 18525 16915
rect 18555 16885 18560 16915
rect 18520 16755 18560 16885
rect 18520 16725 18525 16755
rect 18555 16725 18560 16755
rect 18520 16720 18560 16725
rect 18600 16915 18640 16920
rect 18600 16885 18605 16915
rect 18635 16885 18640 16915
rect 18600 16755 18640 16885
rect 18600 16725 18605 16755
rect 18635 16725 18640 16755
rect 18600 16720 18640 16725
rect 18680 16915 18720 16920
rect 18680 16885 18685 16915
rect 18715 16885 18720 16915
rect 18680 16755 18720 16885
rect 18680 16725 18685 16755
rect 18715 16725 18720 16755
rect 18680 16720 18720 16725
rect 18760 16915 18800 16920
rect 18760 16885 18765 16915
rect 18795 16885 18800 16915
rect 18760 16755 18800 16885
rect 18760 16725 18765 16755
rect 18795 16725 18800 16755
rect 18760 16720 18800 16725
rect 18840 16915 18880 16920
rect 18840 16885 18845 16915
rect 18875 16885 18880 16915
rect 18840 16755 18880 16885
rect 18840 16725 18845 16755
rect 18875 16725 18880 16755
rect 18840 16720 18880 16725
rect 18920 16915 18960 16920
rect 18920 16885 18925 16915
rect 18955 16885 18960 16915
rect 18920 16755 18960 16885
rect 18920 16725 18925 16755
rect 18955 16725 18960 16755
rect 18920 16720 18960 16725
rect 19000 16915 19040 16920
rect 19000 16885 19005 16915
rect 19035 16885 19040 16915
rect 19000 16755 19040 16885
rect 19000 16725 19005 16755
rect 19035 16725 19040 16755
rect 19000 16720 19040 16725
rect 19080 16915 19120 16920
rect 19080 16885 19085 16915
rect 19115 16885 19120 16915
rect 19080 16755 19120 16885
rect 19080 16725 19085 16755
rect 19115 16725 19120 16755
rect 19080 16720 19120 16725
rect 19160 16915 19200 16920
rect 19160 16885 19165 16915
rect 19195 16885 19200 16915
rect 19160 16755 19200 16885
rect 19160 16725 19165 16755
rect 19195 16725 19200 16755
rect 19160 16720 19200 16725
rect 19240 16915 19280 16920
rect 19240 16885 19245 16915
rect 19275 16885 19280 16915
rect 19240 16755 19280 16885
rect 19240 16725 19245 16755
rect 19275 16725 19280 16755
rect 19240 16720 19280 16725
rect 19320 16915 19360 16920
rect 19320 16885 19325 16915
rect 19355 16885 19360 16915
rect 19320 16755 19360 16885
rect 19320 16725 19325 16755
rect 19355 16725 19360 16755
rect 19320 16720 19360 16725
rect 19400 16915 19440 16920
rect 19400 16885 19405 16915
rect 19435 16885 19440 16915
rect 19400 16755 19440 16885
rect 19400 16725 19405 16755
rect 19435 16725 19440 16755
rect 19400 16720 19440 16725
rect 19480 16915 19520 16920
rect 19480 16885 19485 16915
rect 19515 16885 19520 16915
rect 19480 16755 19520 16885
rect 19480 16725 19485 16755
rect 19515 16725 19520 16755
rect 19480 16720 19520 16725
rect 19560 16915 19600 16920
rect 19560 16885 19565 16915
rect 19595 16885 19600 16915
rect 19560 16755 19600 16885
rect 19560 16725 19565 16755
rect 19595 16725 19600 16755
rect 19560 16720 19600 16725
rect 19640 16915 19680 16920
rect 19640 16885 19645 16915
rect 19675 16885 19680 16915
rect 19640 16755 19680 16885
rect 19640 16725 19645 16755
rect 19675 16725 19680 16755
rect 19640 16720 19680 16725
rect 19720 16915 19760 16920
rect 19720 16885 19725 16915
rect 19755 16885 19760 16915
rect 19720 16755 19760 16885
rect 19720 16725 19725 16755
rect 19755 16725 19760 16755
rect 19720 16720 19760 16725
rect 19800 16915 19840 16920
rect 19800 16885 19805 16915
rect 19835 16885 19840 16915
rect 19800 16755 19840 16885
rect 19800 16725 19805 16755
rect 19835 16725 19840 16755
rect 19800 16720 19840 16725
rect 19880 16915 19920 16920
rect 19880 16885 19885 16915
rect 19915 16885 19920 16915
rect 19880 16755 19920 16885
rect 19880 16725 19885 16755
rect 19915 16725 19920 16755
rect 19880 16720 19920 16725
rect 19960 16915 20000 16920
rect 19960 16885 19965 16915
rect 19995 16885 20000 16915
rect 19960 16755 20000 16885
rect 19960 16725 19965 16755
rect 19995 16725 20000 16755
rect 19960 16720 20000 16725
rect 20040 16915 20080 16920
rect 20040 16885 20045 16915
rect 20075 16885 20080 16915
rect 20040 16755 20080 16885
rect 20040 16725 20045 16755
rect 20075 16725 20080 16755
rect 20040 16720 20080 16725
rect 20120 16915 20160 16920
rect 20120 16885 20125 16915
rect 20155 16885 20160 16915
rect 20120 16755 20160 16885
rect 20120 16725 20125 16755
rect 20155 16725 20160 16755
rect 20120 16720 20160 16725
rect 20200 16915 20240 16920
rect 20200 16885 20205 16915
rect 20235 16885 20240 16915
rect 20200 16755 20240 16885
rect 20200 16725 20205 16755
rect 20235 16725 20240 16755
rect 20200 16720 20240 16725
rect 20280 16915 20320 16920
rect 20280 16885 20285 16915
rect 20315 16885 20320 16915
rect 20280 16755 20320 16885
rect 20280 16725 20285 16755
rect 20315 16725 20320 16755
rect 20280 16720 20320 16725
rect 20360 16915 20400 16920
rect 20360 16885 20365 16915
rect 20395 16885 20400 16915
rect 20360 16755 20400 16885
rect 20360 16725 20365 16755
rect 20395 16725 20400 16755
rect 20360 16720 20400 16725
rect 20440 16915 20480 16920
rect 20440 16885 20445 16915
rect 20475 16885 20480 16915
rect 20440 16755 20480 16885
rect 20440 16725 20445 16755
rect 20475 16725 20480 16755
rect 20440 16720 20480 16725
rect 20520 16915 20560 16920
rect 20520 16885 20525 16915
rect 20555 16885 20560 16915
rect 20520 16755 20560 16885
rect 20520 16725 20525 16755
rect 20555 16725 20560 16755
rect 20520 16720 20560 16725
rect 20600 16915 20640 16920
rect 20600 16885 20605 16915
rect 20635 16885 20640 16915
rect 20600 16755 20640 16885
rect 20600 16725 20605 16755
rect 20635 16725 20640 16755
rect 20600 16720 20640 16725
rect 20680 16915 20720 16920
rect 20680 16885 20685 16915
rect 20715 16885 20720 16915
rect 20680 16755 20720 16885
rect 20680 16725 20685 16755
rect 20715 16725 20720 16755
rect 20680 16720 20720 16725
rect 20760 16915 20800 16920
rect 20760 16885 20765 16915
rect 20795 16885 20800 16915
rect 20760 16755 20800 16885
rect 20760 16725 20765 16755
rect 20795 16725 20800 16755
rect 20760 16720 20800 16725
rect 20840 16915 20880 16920
rect 20840 16885 20845 16915
rect 20875 16885 20880 16915
rect 20840 16755 20880 16885
rect 20840 16725 20845 16755
rect 20875 16725 20880 16755
rect 20840 16720 20880 16725
rect 20920 16915 20960 16920
rect 20920 16885 20925 16915
rect 20955 16885 20960 16915
rect 20920 16755 20960 16885
rect 20920 16725 20925 16755
rect 20955 16725 20960 16755
rect 20920 16720 20960 16725
rect 11560 16675 11600 16680
rect 11560 16645 11565 16675
rect 11595 16645 11600 16675
rect 11560 16515 11600 16645
rect 11560 16485 11565 16515
rect 11595 16485 11600 16515
rect 11560 16480 11600 16485
rect 11640 16675 11680 16680
rect 11640 16645 11645 16675
rect 11675 16645 11680 16675
rect 11640 16515 11680 16645
rect 11640 16485 11645 16515
rect 11675 16485 11680 16515
rect 11640 16480 11680 16485
rect 11720 16675 11760 16680
rect 11720 16645 11725 16675
rect 11755 16645 11760 16675
rect 11720 16515 11760 16645
rect 11720 16485 11725 16515
rect 11755 16485 11760 16515
rect 11720 16480 11760 16485
rect 11800 16675 11840 16680
rect 11800 16645 11805 16675
rect 11835 16645 11840 16675
rect 11800 16515 11840 16645
rect 11800 16485 11805 16515
rect 11835 16485 11840 16515
rect 11800 16480 11840 16485
rect 11880 16675 11920 16680
rect 11880 16645 11885 16675
rect 11915 16645 11920 16675
rect 11880 16515 11920 16645
rect 11880 16485 11885 16515
rect 11915 16485 11920 16515
rect 11880 16480 11920 16485
rect 11960 16675 12000 16680
rect 11960 16645 11965 16675
rect 11995 16645 12000 16675
rect 11960 16515 12000 16645
rect 11960 16485 11965 16515
rect 11995 16485 12000 16515
rect 11960 16480 12000 16485
rect 12040 16675 12080 16680
rect 12040 16645 12045 16675
rect 12075 16645 12080 16675
rect 12040 16515 12080 16645
rect 12040 16485 12045 16515
rect 12075 16485 12080 16515
rect 12040 16480 12080 16485
rect 12120 16675 12160 16680
rect 12120 16645 12125 16675
rect 12155 16645 12160 16675
rect 12120 16515 12160 16645
rect 12120 16485 12125 16515
rect 12155 16485 12160 16515
rect 12120 16480 12160 16485
rect 12200 16675 12240 16680
rect 12200 16645 12205 16675
rect 12235 16645 12240 16675
rect 12200 16515 12240 16645
rect 12200 16485 12205 16515
rect 12235 16485 12240 16515
rect 12200 16480 12240 16485
rect 12280 16675 12320 16680
rect 12280 16645 12285 16675
rect 12315 16645 12320 16675
rect 12280 16515 12320 16645
rect 12280 16485 12285 16515
rect 12315 16485 12320 16515
rect 12280 16480 12320 16485
rect 12360 16675 12400 16680
rect 12360 16645 12365 16675
rect 12395 16645 12400 16675
rect 12360 16515 12400 16645
rect 12360 16485 12365 16515
rect 12395 16485 12400 16515
rect 12360 16480 12400 16485
rect 12440 16675 12480 16680
rect 12440 16645 12445 16675
rect 12475 16645 12480 16675
rect 12440 16515 12480 16645
rect 12440 16485 12445 16515
rect 12475 16485 12480 16515
rect 12440 16480 12480 16485
rect 12520 16675 12560 16680
rect 12520 16645 12525 16675
rect 12555 16645 12560 16675
rect 12520 16515 12560 16645
rect 12520 16485 12525 16515
rect 12555 16485 12560 16515
rect 12520 16480 12560 16485
rect 12600 16675 12640 16680
rect 12600 16645 12605 16675
rect 12635 16645 12640 16675
rect 12600 16515 12640 16645
rect 12600 16485 12605 16515
rect 12635 16485 12640 16515
rect 12600 16480 12640 16485
rect 12680 16675 12720 16680
rect 12680 16645 12685 16675
rect 12715 16645 12720 16675
rect 12680 16515 12720 16645
rect 12680 16485 12685 16515
rect 12715 16485 12720 16515
rect 12680 16480 12720 16485
rect 12760 16675 12800 16680
rect 12760 16645 12765 16675
rect 12795 16645 12800 16675
rect 12760 16515 12800 16645
rect 12760 16485 12765 16515
rect 12795 16485 12800 16515
rect 12760 16480 12800 16485
rect 12840 16675 12880 16680
rect 12840 16645 12845 16675
rect 12875 16645 12880 16675
rect 12840 16515 12880 16645
rect 12840 16485 12845 16515
rect 12875 16485 12880 16515
rect 12840 16480 12880 16485
rect 12920 16675 12960 16680
rect 12920 16645 12925 16675
rect 12955 16645 12960 16675
rect 12920 16515 12960 16645
rect 12920 16485 12925 16515
rect 12955 16485 12960 16515
rect 12920 16480 12960 16485
rect 13000 16675 13040 16680
rect 13000 16645 13005 16675
rect 13035 16645 13040 16675
rect 13000 16515 13040 16645
rect 13000 16485 13005 16515
rect 13035 16485 13040 16515
rect 13000 16480 13040 16485
rect 13080 16675 13120 16680
rect 13080 16645 13085 16675
rect 13115 16645 13120 16675
rect 13080 16515 13120 16645
rect 13080 16485 13085 16515
rect 13115 16485 13120 16515
rect 13080 16480 13120 16485
rect 13160 16675 13200 16680
rect 13160 16645 13165 16675
rect 13195 16645 13200 16675
rect 13160 16515 13200 16645
rect 13160 16485 13165 16515
rect 13195 16485 13200 16515
rect 13160 16480 13200 16485
rect 13240 16675 13280 16680
rect 13240 16645 13245 16675
rect 13275 16645 13280 16675
rect 13240 16515 13280 16645
rect 13240 16485 13245 16515
rect 13275 16485 13280 16515
rect 13240 16480 13280 16485
rect 13320 16675 13360 16680
rect 13320 16645 13325 16675
rect 13355 16645 13360 16675
rect 13320 16515 13360 16645
rect 13320 16485 13325 16515
rect 13355 16485 13360 16515
rect 13320 16480 13360 16485
rect 13400 16675 13440 16680
rect 13400 16645 13405 16675
rect 13435 16645 13440 16675
rect 13400 16515 13440 16645
rect 13400 16485 13405 16515
rect 13435 16485 13440 16515
rect 13400 16480 13440 16485
rect 13480 16675 13520 16680
rect 13480 16645 13485 16675
rect 13515 16645 13520 16675
rect 13480 16515 13520 16645
rect 13480 16485 13485 16515
rect 13515 16485 13520 16515
rect 13480 16480 13520 16485
rect 13560 16675 13600 16680
rect 13560 16645 13565 16675
rect 13595 16645 13600 16675
rect 13560 16515 13600 16645
rect 13560 16485 13565 16515
rect 13595 16485 13600 16515
rect 13560 16480 13600 16485
rect 13640 16675 13680 16680
rect 13640 16645 13645 16675
rect 13675 16645 13680 16675
rect 13640 16515 13680 16645
rect 13640 16485 13645 16515
rect 13675 16485 13680 16515
rect 13640 16480 13680 16485
rect 13720 16675 13760 16680
rect 13720 16645 13725 16675
rect 13755 16645 13760 16675
rect 13720 16515 13760 16645
rect 13720 16485 13725 16515
rect 13755 16485 13760 16515
rect 13720 16480 13760 16485
rect 13800 16675 13840 16680
rect 13800 16645 13805 16675
rect 13835 16645 13840 16675
rect 13800 16515 13840 16645
rect 13800 16485 13805 16515
rect 13835 16485 13840 16515
rect 13800 16480 13840 16485
rect 13880 16675 13920 16680
rect 13880 16645 13885 16675
rect 13915 16645 13920 16675
rect 13880 16515 13920 16645
rect 13880 16485 13885 16515
rect 13915 16485 13920 16515
rect 13880 16480 13920 16485
rect 13960 16675 14000 16680
rect 13960 16645 13965 16675
rect 13995 16645 14000 16675
rect 13960 16515 14000 16645
rect 13960 16485 13965 16515
rect 13995 16485 14000 16515
rect 13960 16480 14000 16485
rect 14040 16675 14080 16680
rect 14040 16645 14045 16675
rect 14075 16645 14080 16675
rect 14040 16515 14080 16645
rect 14040 16485 14045 16515
rect 14075 16485 14080 16515
rect 14040 16480 14080 16485
rect 14120 16675 14160 16680
rect 14120 16645 14125 16675
rect 14155 16645 14160 16675
rect 14120 16515 14160 16645
rect 14120 16485 14125 16515
rect 14155 16485 14160 16515
rect 14120 16480 14160 16485
rect 14200 16675 14240 16680
rect 14200 16645 14205 16675
rect 14235 16645 14240 16675
rect 14200 16515 14240 16645
rect 14200 16485 14205 16515
rect 14235 16485 14240 16515
rect 14200 16480 14240 16485
rect 14280 16675 14320 16680
rect 14280 16645 14285 16675
rect 14315 16645 14320 16675
rect 14280 16515 14320 16645
rect 14280 16485 14285 16515
rect 14315 16485 14320 16515
rect 14280 16480 14320 16485
rect 14360 16675 14400 16680
rect 14360 16645 14365 16675
rect 14395 16645 14400 16675
rect 14360 16515 14400 16645
rect 14360 16485 14365 16515
rect 14395 16485 14400 16515
rect 14360 16480 14400 16485
rect 14440 16675 14480 16680
rect 14440 16645 14445 16675
rect 14475 16645 14480 16675
rect 14440 16515 14480 16645
rect 14440 16485 14445 16515
rect 14475 16485 14480 16515
rect 14440 16480 14480 16485
rect 14520 16675 14560 16680
rect 14520 16645 14525 16675
rect 14555 16645 14560 16675
rect 14520 16515 14560 16645
rect 14520 16485 14525 16515
rect 14555 16485 14560 16515
rect 14520 16480 14560 16485
rect 14600 16675 14640 16680
rect 14600 16645 14605 16675
rect 14635 16645 14640 16675
rect 14600 16515 14640 16645
rect 14600 16485 14605 16515
rect 14635 16485 14640 16515
rect 14600 16480 14640 16485
rect 14680 16675 14720 16680
rect 14680 16645 14685 16675
rect 14715 16645 14720 16675
rect 14680 16515 14720 16645
rect 14680 16485 14685 16515
rect 14715 16485 14720 16515
rect 14680 16480 14720 16485
rect 11560 16435 11600 16440
rect 11560 16405 11565 16435
rect 11595 16405 11600 16435
rect 11560 16275 11600 16405
rect 11560 16245 11565 16275
rect 11595 16245 11600 16275
rect 11560 16240 11600 16245
rect 11640 16435 11680 16440
rect 11640 16405 11645 16435
rect 11675 16405 11680 16435
rect 11640 16275 11680 16405
rect 11640 16245 11645 16275
rect 11675 16245 11680 16275
rect 11640 16240 11680 16245
rect 11720 16435 11760 16440
rect 11720 16405 11725 16435
rect 11755 16405 11760 16435
rect 11720 16275 11760 16405
rect 11720 16245 11725 16275
rect 11755 16245 11760 16275
rect 11720 16240 11760 16245
rect 11800 16435 11840 16440
rect 11800 16405 11805 16435
rect 11835 16405 11840 16435
rect 11800 16275 11840 16405
rect 11800 16245 11805 16275
rect 11835 16245 11840 16275
rect 11800 16240 11840 16245
rect 11880 16435 11920 16440
rect 11880 16405 11885 16435
rect 11915 16405 11920 16435
rect 11880 16275 11920 16405
rect 11880 16245 11885 16275
rect 11915 16245 11920 16275
rect 11880 16240 11920 16245
rect 11960 16435 12000 16440
rect 11960 16405 11965 16435
rect 11995 16405 12000 16435
rect 11960 16275 12000 16405
rect 11960 16245 11965 16275
rect 11995 16245 12000 16275
rect 11960 16240 12000 16245
rect 12040 16435 12080 16440
rect 12040 16405 12045 16435
rect 12075 16405 12080 16435
rect 12040 16275 12080 16405
rect 12040 16245 12045 16275
rect 12075 16245 12080 16275
rect 12040 16240 12080 16245
rect 12120 16435 12160 16440
rect 12120 16405 12125 16435
rect 12155 16405 12160 16435
rect 12120 16275 12160 16405
rect 12120 16245 12125 16275
rect 12155 16245 12160 16275
rect 12120 16240 12160 16245
rect 12200 16435 12240 16440
rect 12200 16405 12205 16435
rect 12235 16405 12240 16435
rect 12200 16275 12240 16405
rect 12200 16245 12205 16275
rect 12235 16245 12240 16275
rect 12200 16240 12240 16245
rect 12280 16435 12320 16440
rect 12280 16405 12285 16435
rect 12315 16405 12320 16435
rect 12280 16275 12320 16405
rect 12280 16245 12285 16275
rect 12315 16245 12320 16275
rect 12280 16240 12320 16245
rect 12360 16435 12400 16440
rect 12360 16405 12365 16435
rect 12395 16405 12400 16435
rect 12360 16275 12400 16405
rect 12360 16245 12365 16275
rect 12395 16245 12400 16275
rect 12360 16240 12400 16245
rect 12440 16435 12480 16440
rect 12440 16405 12445 16435
rect 12475 16405 12480 16435
rect 12440 16275 12480 16405
rect 12440 16245 12445 16275
rect 12475 16245 12480 16275
rect 12440 16240 12480 16245
rect 12520 16435 12560 16440
rect 12520 16405 12525 16435
rect 12555 16405 12560 16435
rect 12520 16275 12560 16405
rect 12520 16245 12525 16275
rect 12555 16245 12560 16275
rect 12520 16240 12560 16245
rect 12600 16435 12640 16440
rect 12600 16405 12605 16435
rect 12635 16405 12640 16435
rect 12600 16275 12640 16405
rect 12600 16245 12605 16275
rect 12635 16245 12640 16275
rect 12600 16240 12640 16245
rect 12680 16435 12720 16440
rect 12680 16405 12685 16435
rect 12715 16405 12720 16435
rect 12680 16275 12720 16405
rect 12680 16245 12685 16275
rect 12715 16245 12720 16275
rect 12680 16240 12720 16245
rect 12760 16435 12800 16440
rect 12760 16405 12765 16435
rect 12795 16405 12800 16435
rect 12760 16275 12800 16405
rect 12760 16245 12765 16275
rect 12795 16245 12800 16275
rect 12760 16240 12800 16245
rect 12840 16435 12880 16440
rect 12840 16405 12845 16435
rect 12875 16405 12880 16435
rect 12840 16275 12880 16405
rect 12840 16245 12845 16275
rect 12875 16245 12880 16275
rect 12840 16240 12880 16245
rect 12920 16435 12960 16440
rect 12920 16405 12925 16435
rect 12955 16405 12960 16435
rect 12920 16275 12960 16405
rect 12920 16245 12925 16275
rect 12955 16245 12960 16275
rect 12920 16240 12960 16245
rect 13000 16435 13040 16440
rect 13000 16405 13005 16435
rect 13035 16405 13040 16435
rect 13000 16275 13040 16405
rect 13000 16245 13005 16275
rect 13035 16245 13040 16275
rect 13000 16240 13040 16245
rect 13080 16435 13120 16440
rect 13080 16405 13085 16435
rect 13115 16405 13120 16435
rect 13080 16275 13120 16405
rect 13080 16245 13085 16275
rect 13115 16245 13120 16275
rect 13080 16240 13120 16245
rect 13160 16435 13200 16440
rect 13160 16405 13165 16435
rect 13195 16405 13200 16435
rect 13160 16275 13200 16405
rect 13160 16245 13165 16275
rect 13195 16245 13200 16275
rect 13160 16240 13200 16245
rect 13240 16435 13280 16440
rect 13240 16405 13245 16435
rect 13275 16405 13280 16435
rect 13240 16275 13280 16405
rect 13240 16245 13245 16275
rect 13275 16245 13280 16275
rect 13240 16240 13280 16245
rect 13320 16435 13360 16440
rect 13320 16405 13325 16435
rect 13355 16405 13360 16435
rect 13320 16275 13360 16405
rect 13320 16245 13325 16275
rect 13355 16245 13360 16275
rect 13320 16240 13360 16245
rect 13400 16435 13440 16440
rect 13400 16405 13405 16435
rect 13435 16405 13440 16435
rect 13400 16275 13440 16405
rect 13400 16245 13405 16275
rect 13435 16245 13440 16275
rect 13400 16240 13440 16245
rect 13480 16435 13520 16440
rect 13480 16405 13485 16435
rect 13515 16405 13520 16435
rect 13480 16275 13520 16405
rect 13480 16245 13485 16275
rect 13515 16245 13520 16275
rect 13480 16240 13520 16245
rect 13560 16435 13600 16440
rect 13560 16405 13565 16435
rect 13595 16405 13600 16435
rect 13560 16275 13600 16405
rect 13560 16245 13565 16275
rect 13595 16245 13600 16275
rect 13560 16240 13600 16245
rect 13640 16435 13680 16440
rect 13640 16405 13645 16435
rect 13675 16405 13680 16435
rect 13640 16275 13680 16405
rect 13640 16245 13645 16275
rect 13675 16245 13680 16275
rect 13640 16240 13680 16245
rect 13720 16435 13760 16440
rect 13720 16405 13725 16435
rect 13755 16405 13760 16435
rect 13720 16275 13760 16405
rect 13720 16245 13725 16275
rect 13755 16245 13760 16275
rect 13720 16240 13760 16245
rect 13800 16435 13840 16440
rect 13800 16405 13805 16435
rect 13835 16405 13840 16435
rect 13800 16275 13840 16405
rect 13800 16245 13805 16275
rect 13835 16245 13840 16275
rect 13800 16240 13840 16245
rect 13880 16435 13920 16440
rect 13880 16405 13885 16435
rect 13915 16405 13920 16435
rect 13880 16275 13920 16405
rect 13880 16245 13885 16275
rect 13915 16245 13920 16275
rect 13880 16240 13920 16245
rect 13960 16435 14000 16440
rect 13960 16405 13965 16435
rect 13995 16405 14000 16435
rect 13960 16275 14000 16405
rect 13960 16245 13965 16275
rect 13995 16245 14000 16275
rect 13960 16240 14000 16245
rect 14040 16435 14080 16440
rect 14040 16405 14045 16435
rect 14075 16405 14080 16435
rect 14040 16275 14080 16405
rect 14040 16245 14045 16275
rect 14075 16245 14080 16275
rect 14040 16240 14080 16245
rect 14120 16435 14160 16440
rect 14120 16405 14125 16435
rect 14155 16405 14160 16435
rect 14120 16275 14160 16405
rect 14120 16245 14125 16275
rect 14155 16245 14160 16275
rect 14120 16240 14160 16245
rect 14200 16435 14240 16440
rect 14200 16405 14205 16435
rect 14235 16405 14240 16435
rect 14200 16275 14240 16405
rect 14200 16245 14205 16275
rect 14235 16245 14240 16275
rect 14200 16240 14240 16245
rect 14280 16435 14320 16440
rect 14280 16405 14285 16435
rect 14315 16405 14320 16435
rect 14280 16275 14320 16405
rect 14280 16245 14285 16275
rect 14315 16245 14320 16275
rect 14280 16240 14320 16245
rect 14360 16435 14400 16440
rect 14360 16405 14365 16435
rect 14395 16405 14400 16435
rect 14360 16275 14400 16405
rect 14360 16245 14365 16275
rect 14395 16245 14400 16275
rect 14360 16240 14400 16245
rect 14440 16435 14480 16440
rect 14440 16405 14445 16435
rect 14475 16405 14480 16435
rect 14440 16275 14480 16405
rect 14440 16245 14445 16275
rect 14475 16245 14480 16275
rect 14440 16240 14480 16245
rect 14520 16435 14560 16440
rect 14520 16405 14525 16435
rect 14555 16405 14560 16435
rect 14520 16275 14560 16405
rect 14520 16245 14525 16275
rect 14555 16245 14560 16275
rect 14520 16240 14560 16245
rect 14600 16435 14640 16440
rect 14600 16405 14605 16435
rect 14635 16405 14640 16435
rect 14600 16275 14640 16405
rect 14600 16245 14605 16275
rect 14635 16245 14640 16275
rect 14600 16240 14640 16245
rect 14680 16435 14720 16440
rect 14680 16405 14685 16435
rect 14715 16405 14720 16435
rect 14680 16275 14720 16405
rect 14680 16245 14685 16275
rect 14715 16245 14720 16275
rect 14680 16240 14720 16245
rect 11560 16195 11600 16200
rect 11560 16165 11565 16195
rect 11595 16165 11600 16195
rect 11560 16035 11600 16165
rect 11560 16005 11565 16035
rect 11595 16005 11600 16035
rect 11560 15875 11600 16005
rect 11560 15845 11565 15875
rect 11595 15845 11600 15875
rect 11560 15715 11600 15845
rect 11560 15685 11565 15715
rect 11595 15685 11600 15715
rect 11560 15555 11600 15685
rect 11560 15525 11565 15555
rect 11595 15525 11600 15555
rect 11560 15395 11600 15525
rect 11560 15365 11565 15395
rect 11595 15365 11600 15395
rect 11560 15235 11600 15365
rect 11560 15205 11565 15235
rect 11595 15205 11600 15235
rect 11560 15200 11600 15205
rect 11640 16195 11680 16200
rect 11640 16165 11645 16195
rect 11675 16165 11680 16195
rect 11640 16035 11680 16165
rect 11640 16005 11645 16035
rect 11675 16005 11680 16035
rect 11640 15875 11680 16005
rect 11640 15845 11645 15875
rect 11675 15845 11680 15875
rect 11640 15715 11680 15845
rect 11640 15685 11645 15715
rect 11675 15685 11680 15715
rect 11640 15555 11680 15685
rect 11640 15525 11645 15555
rect 11675 15525 11680 15555
rect 11640 15395 11680 15525
rect 11640 15365 11645 15395
rect 11675 15365 11680 15395
rect 11640 15235 11680 15365
rect 11640 15205 11645 15235
rect 11675 15205 11680 15235
rect 11640 15200 11680 15205
rect 11720 16195 11760 16200
rect 11720 16165 11725 16195
rect 11755 16165 11760 16195
rect 11720 16035 11760 16165
rect 11720 16005 11725 16035
rect 11755 16005 11760 16035
rect 11720 15875 11760 16005
rect 11720 15845 11725 15875
rect 11755 15845 11760 15875
rect 11720 15715 11760 15845
rect 11720 15685 11725 15715
rect 11755 15685 11760 15715
rect 11720 15555 11760 15685
rect 11720 15525 11725 15555
rect 11755 15525 11760 15555
rect 11720 15395 11760 15525
rect 11720 15365 11725 15395
rect 11755 15365 11760 15395
rect 11720 15235 11760 15365
rect 11720 15205 11725 15235
rect 11755 15205 11760 15235
rect 11720 15200 11760 15205
rect 11800 16195 11840 16200
rect 11800 16165 11805 16195
rect 11835 16165 11840 16195
rect 11800 16035 11840 16165
rect 11800 16005 11805 16035
rect 11835 16005 11840 16035
rect 11800 15875 11840 16005
rect 11800 15845 11805 15875
rect 11835 15845 11840 15875
rect 11800 15715 11840 15845
rect 11800 15685 11805 15715
rect 11835 15685 11840 15715
rect 11800 15555 11840 15685
rect 11800 15525 11805 15555
rect 11835 15525 11840 15555
rect 11800 15395 11840 15525
rect 11800 15365 11805 15395
rect 11835 15365 11840 15395
rect 11800 15235 11840 15365
rect 11800 15205 11805 15235
rect 11835 15205 11840 15235
rect 11800 15200 11840 15205
rect 11880 16195 11920 16200
rect 11880 16165 11885 16195
rect 11915 16165 11920 16195
rect 11880 16035 11920 16165
rect 11880 16005 11885 16035
rect 11915 16005 11920 16035
rect 11880 15875 11920 16005
rect 11880 15845 11885 15875
rect 11915 15845 11920 15875
rect 11880 15715 11920 15845
rect 11880 15685 11885 15715
rect 11915 15685 11920 15715
rect 11880 15555 11920 15685
rect 11880 15525 11885 15555
rect 11915 15525 11920 15555
rect 11880 15395 11920 15525
rect 11880 15365 11885 15395
rect 11915 15365 11920 15395
rect 11880 15235 11920 15365
rect 11880 15205 11885 15235
rect 11915 15205 11920 15235
rect 11880 15200 11920 15205
rect 11960 16195 12000 16200
rect 11960 16165 11965 16195
rect 11995 16165 12000 16195
rect 11960 16035 12000 16165
rect 11960 16005 11965 16035
rect 11995 16005 12000 16035
rect 11960 15875 12000 16005
rect 11960 15845 11965 15875
rect 11995 15845 12000 15875
rect 11960 15715 12000 15845
rect 11960 15685 11965 15715
rect 11995 15685 12000 15715
rect 11960 15555 12000 15685
rect 11960 15525 11965 15555
rect 11995 15525 12000 15555
rect 11960 15395 12000 15525
rect 11960 15365 11965 15395
rect 11995 15365 12000 15395
rect 11960 15235 12000 15365
rect 11960 15205 11965 15235
rect 11995 15205 12000 15235
rect 11960 15200 12000 15205
rect 12040 16195 12080 16200
rect 12040 16165 12045 16195
rect 12075 16165 12080 16195
rect 12040 16035 12080 16165
rect 12040 16005 12045 16035
rect 12075 16005 12080 16035
rect 12040 15875 12080 16005
rect 12040 15845 12045 15875
rect 12075 15845 12080 15875
rect 12040 15715 12080 15845
rect 12040 15685 12045 15715
rect 12075 15685 12080 15715
rect 12040 15555 12080 15685
rect 12040 15525 12045 15555
rect 12075 15525 12080 15555
rect 12040 15395 12080 15525
rect 12040 15365 12045 15395
rect 12075 15365 12080 15395
rect 12040 15235 12080 15365
rect 12040 15205 12045 15235
rect 12075 15205 12080 15235
rect 12040 15200 12080 15205
rect 12120 16195 12160 16200
rect 12120 16165 12125 16195
rect 12155 16165 12160 16195
rect 12120 16035 12160 16165
rect 12120 16005 12125 16035
rect 12155 16005 12160 16035
rect 12120 15875 12160 16005
rect 12120 15845 12125 15875
rect 12155 15845 12160 15875
rect 12120 15715 12160 15845
rect 12120 15685 12125 15715
rect 12155 15685 12160 15715
rect 12120 15555 12160 15685
rect 12120 15525 12125 15555
rect 12155 15525 12160 15555
rect 12120 15395 12160 15525
rect 12120 15365 12125 15395
rect 12155 15365 12160 15395
rect 12120 15235 12160 15365
rect 12120 15205 12125 15235
rect 12155 15205 12160 15235
rect 12120 15200 12160 15205
rect 12200 16195 12240 16200
rect 12200 16165 12205 16195
rect 12235 16165 12240 16195
rect 12200 16035 12240 16165
rect 12200 16005 12205 16035
rect 12235 16005 12240 16035
rect 12200 15875 12240 16005
rect 12200 15845 12205 15875
rect 12235 15845 12240 15875
rect 12200 15715 12240 15845
rect 12200 15685 12205 15715
rect 12235 15685 12240 15715
rect 12200 15555 12240 15685
rect 12200 15525 12205 15555
rect 12235 15525 12240 15555
rect 12200 15395 12240 15525
rect 12200 15365 12205 15395
rect 12235 15365 12240 15395
rect 12200 15235 12240 15365
rect 12200 15205 12205 15235
rect 12235 15205 12240 15235
rect 12200 15200 12240 15205
rect 12280 16195 12320 16200
rect 12280 16165 12285 16195
rect 12315 16165 12320 16195
rect 12280 16035 12320 16165
rect 12280 16005 12285 16035
rect 12315 16005 12320 16035
rect 12280 15875 12320 16005
rect 12280 15845 12285 15875
rect 12315 15845 12320 15875
rect 12280 15715 12320 15845
rect 12280 15685 12285 15715
rect 12315 15685 12320 15715
rect 12280 15555 12320 15685
rect 12280 15525 12285 15555
rect 12315 15525 12320 15555
rect 12280 15395 12320 15525
rect 12280 15365 12285 15395
rect 12315 15365 12320 15395
rect 12280 15235 12320 15365
rect 12280 15205 12285 15235
rect 12315 15205 12320 15235
rect 12280 15200 12320 15205
rect 12360 16195 12400 16200
rect 12360 16165 12365 16195
rect 12395 16165 12400 16195
rect 12360 16035 12400 16165
rect 12360 16005 12365 16035
rect 12395 16005 12400 16035
rect 12360 15875 12400 16005
rect 12360 15845 12365 15875
rect 12395 15845 12400 15875
rect 12360 15715 12400 15845
rect 12360 15685 12365 15715
rect 12395 15685 12400 15715
rect 12360 15555 12400 15685
rect 12360 15525 12365 15555
rect 12395 15525 12400 15555
rect 12360 15395 12400 15525
rect 12360 15365 12365 15395
rect 12395 15365 12400 15395
rect 12360 15235 12400 15365
rect 12360 15205 12365 15235
rect 12395 15205 12400 15235
rect 12360 15200 12400 15205
rect 12440 16195 12480 16200
rect 12440 16165 12445 16195
rect 12475 16165 12480 16195
rect 12440 16035 12480 16165
rect 12440 16005 12445 16035
rect 12475 16005 12480 16035
rect 12440 15875 12480 16005
rect 12440 15845 12445 15875
rect 12475 15845 12480 15875
rect 12440 15715 12480 15845
rect 12440 15685 12445 15715
rect 12475 15685 12480 15715
rect 12440 15555 12480 15685
rect 12440 15525 12445 15555
rect 12475 15525 12480 15555
rect 12440 15395 12480 15525
rect 12440 15365 12445 15395
rect 12475 15365 12480 15395
rect 12440 15235 12480 15365
rect 12440 15205 12445 15235
rect 12475 15205 12480 15235
rect 12440 15200 12480 15205
rect 12520 16195 12560 16200
rect 12520 16165 12525 16195
rect 12555 16165 12560 16195
rect 12520 16035 12560 16165
rect 12520 16005 12525 16035
rect 12555 16005 12560 16035
rect 12520 15875 12560 16005
rect 12520 15845 12525 15875
rect 12555 15845 12560 15875
rect 12520 15715 12560 15845
rect 12520 15685 12525 15715
rect 12555 15685 12560 15715
rect 12520 15555 12560 15685
rect 12520 15525 12525 15555
rect 12555 15525 12560 15555
rect 12520 15395 12560 15525
rect 12520 15365 12525 15395
rect 12555 15365 12560 15395
rect 12520 15235 12560 15365
rect 12520 15205 12525 15235
rect 12555 15205 12560 15235
rect 12520 15200 12560 15205
rect 12600 16195 12640 16200
rect 12600 16165 12605 16195
rect 12635 16165 12640 16195
rect 12600 16035 12640 16165
rect 12600 16005 12605 16035
rect 12635 16005 12640 16035
rect 12600 15875 12640 16005
rect 12600 15845 12605 15875
rect 12635 15845 12640 15875
rect 12600 15715 12640 15845
rect 12600 15685 12605 15715
rect 12635 15685 12640 15715
rect 12600 15555 12640 15685
rect 12600 15525 12605 15555
rect 12635 15525 12640 15555
rect 12600 15395 12640 15525
rect 12600 15365 12605 15395
rect 12635 15365 12640 15395
rect 12600 15235 12640 15365
rect 12600 15205 12605 15235
rect 12635 15205 12640 15235
rect 12600 15200 12640 15205
rect 12680 16195 12720 16200
rect 12680 16165 12685 16195
rect 12715 16165 12720 16195
rect 12680 16035 12720 16165
rect 12680 16005 12685 16035
rect 12715 16005 12720 16035
rect 12680 15875 12720 16005
rect 12680 15845 12685 15875
rect 12715 15845 12720 15875
rect 12680 15715 12720 15845
rect 12680 15685 12685 15715
rect 12715 15685 12720 15715
rect 12680 15555 12720 15685
rect 12680 15525 12685 15555
rect 12715 15525 12720 15555
rect 12680 15395 12720 15525
rect 12680 15365 12685 15395
rect 12715 15365 12720 15395
rect 12680 15235 12720 15365
rect 12680 15205 12685 15235
rect 12715 15205 12720 15235
rect 12680 15200 12720 15205
rect 12760 16195 12800 16200
rect 12760 16165 12765 16195
rect 12795 16165 12800 16195
rect 12760 16035 12800 16165
rect 12760 16005 12765 16035
rect 12795 16005 12800 16035
rect 12760 15875 12800 16005
rect 12760 15845 12765 15875
rect 12795 15845 12800 15875
rect 12760 15715 12800 15845
rect 12760 15685 12765 15715
rect 12795 15685 12800 15715
rect 12760 15555 12800 15685
rect 12760 15525 12765 15555
rect 12795 15525 12800 15555
rect 12760 15395 12800 15525
rect 12760 15365 12765 15395
rect 12795 15365 12800 15395
rect 12760 15235 12800 15365
rect 12760 15205 12765 15235
rect 12795 15205 12800 15235
rect 12760 15200 12800 15205
rect 12840 16195 12880 16200
rect 12840 16165 12845 16195
rect 12875 16165 12880 16195
rect 12840 16035 12880 16165
rect 12840 16005 12845 16035
rect 12875 16005 12880 16035
rect 12840 15875 12880 16005
rect 12840 15845 12845 15875
rect 12875 15845 12880 15875
rect 12840 15715 12880 15845
rect 12840 15685 12845 15715
rect 12875 15685 12880 15715
rect 12840 15555 12880 15685
rect 12840 15525 12845 15555
rect 12875 15525 12880 15555
rect 12840 15395 12880 15525
rect 12840 15365 12845 15395
rect 12875 15365 12880 15395
rect 12840 15235 12880 15365
rect 12840 15205 12845 15235
rect 12875 15205 12880 15235
rect 12840 15200 12880 15205
rect 12920 16195 12960 16200
rect 12920 16165 12925 16195
rect 12955 16165 12960 16195
rect 12920 16035 12960 16165
rect 12920 16005 12925 16035
rect 12955 16005 12960 16035
rect 12920 15875 12960 16005
rect 12920 15845 12925 15875
rect 12955 15845 12960 15875
rect 12920 15715 12960 15845
rect 12920 15685 12925 15715
rect 12955 15685 12960 15715
rect 12920 15555 12960 15685
rect 12920 15525 12925 15555
rect 12955 15525 12960 15555
rect 12920 15395 12960 15525
rect 12920 15365 12925 15395
rect 12955 15365 12960 15395
rect 12920 15235 12960 15365
rect 12920 15205 12925 15235
rect 12955 15205 12960 15235
rect 12920 15200 12960 15205
rect 13000 16195 13040 16200
rect 13000 16165 13005 16195
rect 13035 16165 13040 16195
rect 13000 16035 13040 16165
rect 13000 16005 13005 16035
rect 13035 16005 13040 16035
rect 13000 15875 13040 16005
rect 13000 15845 13005 15875
rect 13035 15845 13040 15875
rect 13000 15715 13040 15845
rect 13000 15685 13005 15715
rect 13035 15685 13040 15715
rect 13000 15555 13040 15685
rect 13000 15525 13005 15555
rect 13035 15525 13040 15555
rect 13000 15395 13040 15525
rect 13000 15365 13005 15395
rect 13035 15365 13040 15395
rect 13000 15235 13040 15365
rect 13000 15205 13005 15235
rect 13035 15205 13040 15235
rect 13000 15200 13040 15205
rect 13080 16195 13120 16200
rect 13080 16165 13085 16195
rect 13115 16165 13120 16195
rect 13080 16035 13120 16165
rect 13080 16005 13085 16035
rect 13115 16005 13120 16035
rect 13080 15875 13120 16005
rect 13080 15845 13085 15875
rect 13115 15845 13120 15875
rect 13080 15715 13120 15845
rect 13080 15685 13085 15715
rect 13115 15685 13120 15715
rect 13080 15555 13120 15685
rect 13080 15525 13085 15555
rect 13115 15525 13120 15555
rect 13080 15395 13120 15525
rect 13080 15365 13085 15395
rect 13115 15365 13120 15395
rect 13080 15235 13120 15365
rect 13080 15205 13085 15235
rect 13115 15205 13120 15235
rect 13080 15200 13120 15205
rect 13160 16195 13200 16200
rect 13160 16165 13165 16195
rect 13195 16165 13200 16195
rect 13160 16035 13200 16165
rect 13160 16005 13165 16035
rect 13195 16005 13200 16035
rect 13160 15875 13200 16005
rect 13160 15845 13165 15875
rect 13195 15845 13200 15875
rect 13160 15715 13200 15845
rect 13160 15685 13165 15715
rect 13195 15685 13200 15715
rect 13160 15555 13200 15685
rect 13160 15525 13165 15555
rect 13195 15525 13200 15555
rect 13160 15395 13200 15525
rect 13160 15365 13165 15395
rect 13195 15365 13200 15395
rect 13160 15235 13200 15365
rect 13160 15205 13165 15235
rect 13195 15205 13200 15235
rect 13160 15200 13200 15205
rect 13240 16195 13280 16200
rect 13240 16165 13245 16195
rect 13275 16165 13280 16195
rect 13240 16035 13280 16165
rect 13240 16005 13245 16035
rect 13275 16005 13280 16035
rect 13240 15875 13280 16005
rect 13240 15845 13245 15875
rect 13275 15845 13280 15875
rect 13240 15715 13280 15845
rect 13240 15685 13245 15715
rect 13275 15685 13280 15715
rect 13240 15555 13280 15685
rect 13240 15525 13245 15555
rect 13275 15525 13280 15555
rect 13240 15395 13280 15525
rect 13240 15365 13245 15395
rect 13275 15365 13280 15395
rect 13240 15235 13280 15365
rect 13240 15205 13245 15235
rect 13275 15205 13280 15235
rect 13240 15200 13280 15205
rect 13320 16195 13360 16200
rect 13320 16165 13325 16195
rect 13355 16165 13360 16195
rect 13320 16035 13360 16165
rect 13320 16005 13325 16035
rect 13355 16005 13360 16035
rect 13320 15875 13360 16005
rect 13320 15845 13325 15875
rect 13355 15845 13360 15875
rect 13320 15715 13360 15845
rect 13320 15685 13325 15715
rect 13355 15685 13360 15715
rect 13320 15555 13360 15685
rect 13320 15525 13325 15555
rect 13355 15525 13360 15555
rect 13320 15395 13360 15525
rect 13320 15365 13325 15395
rect 13355 15365 13360 15395
rect 13320 15235 13360 15365
rect 13320 15205 13325 15235
rect 13355 15205 13360 15235
rect 13320 15200 13360 15205
rect 13400 16195 13440 16200
rect 13400 16165 13405 16195
rect 13435 16165 13440 16195
rect 13400 16035 13440 16165
rect 13400 16005 13405 16035
rect 13435 16005 13440 16035
rect 13400 15875 13440 16005
rect 13400 15845 13405 15875
rect 13435 15845 13440 15875
rect 13400 15715 13440 15845
rect 13400 15685 13405 15715
rect 13435 15685 13440 15715
rect 13400 15555 13440 15685
rect 13400 15525 13405 15555
rect 13435 15525 13440 15555
rect 13400 15395 13440 15525
rect 13400 15365 13405 15395
rect 13435 15365 13440 15395
rect 13400 15235 13440 15365
rect 13400 15205 13405 15235
rect 13435 15205 13440 15235
rect 13400 15200 13440 15205
rect 13480 16195 13520 16200
rect 13480 16165 13485 16195
rect 13515 16165 13520 16195
rect 13480 16035 13520 16165
rect 13480 16005 13485 16035
rect 13515 16005 13520 16035
rect 13480 15875 13520 16005
rect 13480 15845 13485 15875
rect 13515 15845 13520 15875
rect 13480 15715 13520 15845
rect 13480 15685 13485 15715
rect 13515 15685 13520 15715
rect 13480 15555 13520 15685
rect 13480 15525 13485 15555
rect 13515 15525 13520 15555
rect 13480 15395 13520 15525
rect 13480 15365 13485 15395
rect 13515 15365 13520 15395
rect 13480 15235 13520 15365
rect 13480 15205 13485 15235
rect 13515 15205 13520 15235
rect 13480 15200 13520 15205
rect 13560 16195 13600 16200
rect 13560 16165 13565 16195
rect 13595 16165 13600 16195
rect 13560 16035 13600 16165
rect 13560 16005 13565 16035
rect 13595 16005 13600 16035
rect 13560 15875 13600 16005
rect 13560 15845 13565 15875
rect 13595 15845 13600 15875
rect 13560 15715 13600 15845
rect 13560 15685 13565 15715
rect 13595 15685 13600 15715
rect 13560 15555 13600 15685
rect 13560 15525 13565 15555
rect 13595 15525 13600 15555
rect 13560 15395 13600 15525
rect 13560 15365 13565 15395
rect 13595 15365 13600 15395
rect 13560 15235 13600 15365
rect 13560 15205 13565 15235
rect 13595 15205 13600 15235
rect 13560 15200 13600 15205
rect 13640 16195 13680 16200
rect 13640 16165 13645 16195
rect 13675 16165 13680 16195
rect 13640 16035 13680 16165
rect 13640 16005 13645 16035
rect 13675 16005 13680 16035
rect 13640 15875 13680 16005
rect 13640 15845 13645 15875
rect 13675 15845 13680 15875
rect 13640 15715 13680 15845
rect 13640 15685 13645 15715
rect 13675 15685 13680 15715
rect 13640 15555 13680 15685
rect 13640 15525 13645 15555
rect 13675 15525 13680 15555
rect 13640 15395 13680 15525
rect 13640 15365 13645 15395
rect 13675 15365 13680 15395
rect 13640 15235 13680 15365
rect 13640 15205 13645 15235
rect 13675 15205 13680 15235
rect 13640 15200 13680 15205
rect 13720 16195 13760 16200
rect 13720 16165 13725 16195
rect 13755 16165 13760 16195
rect 13720 16035 13760 16165
rect 13720 16005 13725 16035
rect 13755 16005 13760 16035
rect 13720 15875 13760 16005
rect 13720 15845 13725 15875
rect 13755 15845 13760 15875
rect 13720 15715 13760 15845
rect 13720 15685 13725 15715
rect 13755 15685 13760 15715
rect 13720 15555 13760 15685
rect 13720 15525 13725 15555
rect 13755 15525 13760 15555
rect 13720 15395 13760 15525
rect 13720 15365 13725 15395
rect 13755 15365 13760 15395
rect 13720 15235 13760 15365
rect 13720 15205 13725 15235
rect 13755 15205 13760 15235
rect 13720 15200 13760 15205
rect 13800 16195 13840 16200
rect 13800 16165 13805 16195
rect 13835 16165 13840 16195
rect 13800 16035 13840 16165
rect 13800 16005 13805 16035
rect 13835 16005 13840 16035
rect 13800 15875 13840 16005
rect 13800 15845 13805 15875
rect 13835 15845 13840 15875
rect 13800 15715 13840 15845
rect 13800 15685 13805 15715
rect 13835 15685 13840 15715
rect 13800 15555 13840 15685
rect 13800 15525 13805 15555
rect 13835 15525 13840 15555
rect 13800 15395 13840 15525
rect 13800 15365 13805 15395
rect 13835 15365 13840 15395
rect 13800 15235 13840 15365
rect 13800 15205 13805 15235
rect 13835 15205 13840 15235
rect 13800 15200 13840 15205
rect 13880 16195 13920 16200
rect 13880 16165 13885 16195
rect 13915 16165 13920 16195
rect 13880 16035 13920 16165
rect 13880 16005 13885 16035
rect 13915 16005 13920 16035
rect 13880 15875 13920 16005
rect 13880 15845 13885 15875
rect 13915 15845 13920 15875
rect 13880 15715 13920 15845
rect 13880 15685 13885 15715
rect 13915 15685 13920 15715
rect 13880 15555 13920 15685
rect 13880 15525 13885 15555
rect 13915 15525 13920 15555
rect 13880 15395 13920 15525
rect 13880 15365 13885 15395
rect 13915 15365 13920 15395
rect 13880 15235 13920 15365
rect 13880 15205 13885 15235
rect 13915 15205 13920 15235
rect 13880 15200 13920 15205
rect 13960 16195 14000 16200
rect 13960 16165 13965 16195
rect 13995 16165 14000 16195
rect 13960 16035 14000 16165
rect 13960 16005 13965 16035
rect 13995 16005 14000 16035
rect 13960 15875 14000 16005
rect 13960 15845 13965 15875
rect 13995 15845 14000 15875
rect 13960 15715 14000 15845
rect 13960 15685 13965 15715
rect 13995 15685 14000 15715
rect 13960 15555 14000 15685
rect 13960 15525 13965 15555
rect 13995 15525 14000 15555
rect 13960 15395 14000 15525
rect 13960 15365 13965 15395
rect 13995 15365 14000 15395
rect 13960 15235 14000 15365
rect 13960 15205 13965 15235
rect 13995 15205 14000 15235
rect 13960 15200 14000 15205
rect 14040 16195 14080 16200
rect 14040 16165 14045 16195
rect 14075 16165 14080 16195
rect 14040 16035 14080 16165
rect 14040 16005 14045 16035
rect 14075 16005 14080 16035
rect 14040 15875 14080 16005
rect 14040 15845 14045 15875
rect 14075 15845 14080 15875
rect 14040 15715 14080 15845
rect 14040 15685 14045 15715
rect 14075 15685 14080 15715
rect 14040 15555 14080 15685
rect 14040 15525 14045 15555
rect 14075 15525 14080 15555
rect 14040 15395 14080 15525
rect 14040 15365 14045 15395
rect 14075 15365 14080 15395
rect 14040 15235 14080 15365
rect 14040 15205 14045 15235
rect 14075 15205 14080 15235
rect 14040 15200 14080 15205
rect 14120 16195 14160 16200
rect 14120 16165 14125 16195
rect 14155 16165 14160 16195
rect 14120 16035 14160 16165
rect 14120 16005 14125 16035
rect 14155 16005 14160 16035
rect 14120 15875 14160 16005
rect 14120 15845 14125 15875
rect 14155 15845 14160 15875
rect 14120 15715 14160 15845
rect 14120 15685 14125 15715
rect 14155 15685 14160 15715
rect 14120 15555 14160 15685
rect 14120 15525 14125 15555
rect 14155 15525 14160 15555
rect 14120 15395 14160 15525
rect 14120 15365 14125 15395
rect 14155 15365 14160 15395
rect 14120 15235 14160 15365
rect 14120 15205 14125 15235
rect 14155 15205 14160 15235
rect 14120 15200 14160 15205
rect 14200 16195 14240 16200
rect 14200 16165 14205 16195
rect 14235 16165 14240 16195
rect 14200 16035 14240 16165
rect 14200 16005 14205 16035
rect 14235 16005 14240 16035
rect 14200 15875 14240 16005
rect 14200 15845 14205 15875
rect 14235 15845 14240 15875
rect 14200 15715 14240 15845
rect 14200 15685 14205 15715
rect 14235 15685 14240 15715
rect 14200 15555 14240 15685
rect 14200 15525 14205 15555
rect 14235 15525 14240 15555
rect 14200 15395 14240 15525
rect 14200 15365 14205 15395
rect 14235 15365 14240 15395
rect 14200 15235 14240 15365
rect 14200 15205 14205 15235
rect 14235 15205 14240 15235
rect 14200 15200 14240 15205
rect 14280 16195 14320 16200
rect 14280 16165 14285 16195
rect 14315 16165 14320 16195
rect 14280 16035 14320 16165
rect 14280 16005 14285 16035
rect 14315 16005 14320 16035
rect 14280 15875 14320 16005
rect 14280 15845 14285 15875
rect 14315 15845 14320 15875
rect 14280 15715 14320 15845
rect 14280 15685 14285 15715
rect 14315 15685 14320 15715
rect 14280 15555 14320 15685
rect 14280 15525 14285 15555
rect 14315 15525 14320 15555
rect 14280 15395 14320 15525
rect 14280 15365 14285 15395
rect 14315 15365 14320 15395
rect 14280 15235 14320 15365
rect 14280 15205 14285 15235
rect 14315 15205 14320 15235
rect 14280 15200 14320 15205
rect 14360 16195 14400 16200
rect 14360 16165 14365 16195
rect 14395 16165 14400 16195
rect 14360 16035 14400 16165
rect 14360 16005 14365 16035
rect 14395 16005 14400 16035
rect 14360 15875 14400 16005
rect 14360 15845 14365 15875
rect 14395 15845 14400 15875
rect 14360 15715 14400 15845
rect 14360 15685 14365 15715
rect 14395 15685 14400 15715
rect 14360 15555 14400 15685
rect 14360 15525 14365 15555
rect 14395 15525 14400 15555
rect 14360 15395 14400 15525
rect 14360 15365 14365 15395
rect 14395 15365 14400 15395
rect 14360 15235 14400 15365
rect 14360 15205 14365 15235
rect 14395 15205 14400 15235
rect 14360 15200 14400 15205
rect 14440 16195 14480 16200
rect 14440 16165 14445 16195
rect 14475 16165 14480 16195
rect 14440 16035 14480 16165
rect 14440 16005 14445 16035
rect 14475 16005 14480 16035
rect 14440 15875 14480 16005
rect 14440 15845 14445 15875
rect 14475 15845 14480 15875
rect 14440 15715 14480 15845
rect 14440 15685 14445 15715
rect 14475 15685 14480 15715
rect 14440 15555 14480 15685
rect 14440 15525 14445 15555
rect 14475 15525 14480 15555
rect 14440 15395 14480 15525
rect 14440 15365 14445 15395
rect 14475 15365 14480 15395
rect 14440 15235 14480 15365
rect 14440 15205 14445 15235
rect 14475 15205 14480 15235
rect 14440 15200 14480 15205
rect 14520 16195 14560 16200
rect 14520 16165 14525 16195
rect 14555 16165 14560 16195
rect 14520 16035 14560 16165
rect 14520 16005 14525 16035
rect 14555 16005 14560 16035
rect 14520 15875 14560 16005
rect 14520 15845 14525 15875
rect 14555 15845 14560 15875
rect 14520 15715 14560 15845
rect 14520 15685 14525 15715
rect 14555 15685 14560 15715
rect 14520 15555 14560 15685
rect 14520 15525 14525 15555
rect 14555 15525 14560 15555
rect 14520 15395 14560 15525
rect 14520 15365 14525 15395
rect 14555 15365 14560 15395
rect 14520 15235 14560 15365
rect 14520 15205 14525 15235
rect 14555 15205 14560 15235
rect 14520 15200 14560 15205
rect 14600 16195 14640 16200
rect 14600 16165 14605 16195
rect 14635 16165 14640 16195
rect 14600 16035 14640 16165
rect 14600 16005 14605 16035
rect 14635 16005 14640 16035
rect 14600 15875 14640 16005
rect 14600 15845 14605 15875
rect 14635 15845 14640 15875
rect 14600 15715 14640 15845
rect 14600 15685 14605 15715
rect 14635 15685 14640 15715
rect 14600 15555 14640 15685
rect 14600 15525 14605 15555
rect 14635 15525 14640 15555
rect 14600 15395 14640 15525
rect 14600 15365 14605 15395
rect 14635 15365 14640 15395
rect 14600 15235 14640 15365
rect 14600 15205 14605 15235
rect 14635 15205 14640 15235
rect 14600 15200 14640 15205
rect 14680 16195 14720 16200
rect 14680 16165 14685 16195
rect 14715 16165 14720 16195
rect 14680 16035 14720 16165
rect 14680 16005 14685 16035
rect 14715 16005 14720 16035
rect 14680 15875 14720 16005
rect 14680 15845 14685 15875
rect 14715 15845 14720 15875
rect 14680 15715 14720 15845
rect 14680 15685 14685 15715
rect 14715 15685 14720 15715
rect 14680 15555 14720 15685
rect 14680 15525 14685 15555
rect 14715 15525 14720 15555
rect 14680 15395 14720 15525
rect 14680 15365 14685 15395
rect 14715 15365 14720 15395
rect 14680 15235 14720 15365
rect 14680 15205 14685 15235
rect 14715 15205 14720 15235
rect 14680 15200 14720 15205
rect 11560 15155 11600 15160
rect 11560 15125 11565 15155
rect 11595 15125 11600 15155
rect 11560 14995 11600 15125
rect 11560 14965 11565 14995
rect 11595 14965 11600 14995
rect 11560 14960 11600 14965
rect 11640 15155 11680 15160
rect 11640 15125 11645 15155
rect 11675 15125 11680 15155
rect 11640 14995 11680 15125
rect 11640 14965 11645 14995
rect 11675 14965 11680 14995
rect 11640 14960 11680 14965
rect 11720 15155 11760 15160
rect 11720 15125 11725 15155
rect 11755 15125 11760 15155
rect 11720 14995 11760 15125
rect 11720 14965 11725 14995
rect 11755 14965 11760 14995
rect 11720 14960 11760 14965
rect 11800 15155 11840 15160
rect 11800 15125 11805 15155
rect 11835 15125 11840 15155
rect 11800 14995 11840 15125
rect 11800 14965 11805 14995
rect 11835 14965 11840 14995
rect 11800 14960 11840 14965
rect 11880 15155 11920 15160
rect 11880 15125 11885 15155
rect 11915 15125 11920 15155
rect 11880 14995 11920 15125
rect 11880 14965 11885 14995
rect 11915 14965 11920 14995
rect 11880 14960 11920 14965
rect 11960 15155 12000 15160
rect 11960 15125 11965 15155
rect 11995 15125 12000 15155
rect 11960 14995 12000 15125
rect 11960 14965 11965 14995
rect 11995 14965 12000 14995
rect 11960 14960 12000 14965
rect 12040 15155 12080 15160
rect 12040 15125 12045 15155
rect 12075 15125 12080 15155
rect 12040 14995 12080 15125
rect 12040 14965 12045 14995
rect 12075 14965 12080 14995
rect 12040 14960 12080 14965
rect 12120 15155 12160 15160
rect 12120 15125 12125 15155
rect 12155 15125 12160 15155
rect 12120 14995 12160 15125
rect 12120 14965 12125 14995
rect 12155 14965 12160 14995
rect 12120 14960 12160 14965
rect 12200 15155 12240 15160
rect 12200 15125 12205 15155
rect 12235 15125 12240 15155
rect 12200 14995 12240 15125
rect 12200 14965 12205 14995
rect 12235 14965 12240 14995
rect 12200 14960 12240 14965
rect 12280 15155 12320 15160
rect 12280 15125 12285 15155
rect 12315 15125 12320 15155
rect 12280 14995 12320 15125
rect 12280 14965 12285 14995
rect 12315 14965 12320 14995
rect 12280 14960 12320 14965
rect 12360 15155 12400 15160
rect 12360 15125 12365 15155
rect 12395 15125 12400 15155
rect 12360 14995 12400 15125
rect 12360 14965 12365 14995
rect 12395 14965 12400 14995
rect 12360 14960 12400 14965
rect 12440 15155 12480 15160
rect 12440 15125 12445 15155
rect 12475 15125 12480 15155
rect 12440 14995 12480 15125
rect 12440 14965 12445 14995
rect 12475 14965 12480 14995
rect 12440 14960 12480 14965
rect 12520 15155 12560 15160
rect 12520 15125 12525 15155
rect 12555 15125 12560 15155
rect 12520 14995 12560 15125
rect 12520 14965 12525 14995
rect 12555 14965 12560 14995
rect 12520 14960 12560 14965
rect 12600 15155 12640 15160
rect 12600 15125 12605 15155
rect 12635 15125 12640 15155
rect 12600 14995 12640 15125
rect 12600 14965 12605 14995
rect 12635 14965 12640 14995
rect 12600 14960 12640 14965
rect 12680 15155 12720 15160
rect 12680 15125 12685 15155
rect 12715 15125 12720 15155
rect 12680 14995 12720 15125
rect 12680 14965 12685 14995
rect 12715 14965 12720 14995
rect 12680 14960 12720 14965
rect 12760 15155 12800 15160
rect 12760 15125 12765 15155
rect 12795 15125 12800 15155
rect 12760 14995 12800 15125
rect 12760 14965 12765 14995
rect 12795 14965 12800 14995
rect 12760 14960 12800 14965
rect 12840 15155 12880 15160
rect 12840 15125 12845 15155
rect 12875 15125 12880 15155
rect 12840 14995 12880 15125
rect 12840 14965 12845 14995
rect 12875 14965 12880 14995
rect 12840 14960 12880 14965
rect 12920 15155 12960 15160
rect 12920 15125 12925 15155
rect 12955 15125 12960 15155
rect 12920 14995 12960 15125
rect 12920 14965 12925 14995
rect 12955 14965 12960 14995
rect 12920 14960 12960 14965
rect 13000 15155 13040 15160
rect 13000 15125 13005 15155
rect 13035 15125 13040 15155
rect 13000 14995 13040 15125
rect 13000 14965 13005 14995
rect 13035 14965 13040 14995
rect 13000 14960 13040 14965
rect 13080 15155 13120 15160
rect 13080 15125 13085 15155
rect 13115 15125 13120 15155
rect 13080 14995 13120 15125
rect 13080 14965 13085 14995
rect 13115 14965 13120 14995
rect 13080 14960 13120 14965
rect 13160 15155 13200 15160
rect 13160 15125 13165 15155
rect 13195 15125 13200 15155
rect 13160 14995 13200 15125
rect 13160 14965 13165 14995
rect 13195 14965 13200 14995
rect 13160 14960 13200 14965
rect 13240 15155 13280 15160
rect 13240 15125 13245 15155
rect 13275 15125 13280 15155
rect 13240 14995 13280 15125
rect 13240 14965 13245 14995
rect 13275 14965 13280 14995
rect 13240 14960 13280 14965
rect 13320 15155 13360 15160
rect 13320 15125 13325 15155
rect 13355 15125 13360 15155
rect 13320 14995 13360 15125
rect 13320 14965 13325 14995
rect 13355 14965 13360 14995
rect 13320 14960 13360 14965
rect 13400 15155 13440 15160
rect 13400 15125 13405 15155
rect 13435 15125 13440 15155
rect 13400 14995 13440 15125
rect 13400 14965 13405 14995
rect 13435 14965 13440 14995
rect 13400 14960 13440 14965
rect 13480 15155 13520 15160
rect 13480 15125 13485 15155
rect 13515 15125 13520 15155
rect 13480 14995 13520 15125
rect 13480 14965 13485 14995
rect 13515 14965 13520 14995
rect 13480 14960 13520 14965
rect 13560 15155 13600 15160
rect 13560 15125 13565 15155
rect 13595 15125 13600 15155
rect 13560 14995 13600 15125
rect 13560 14965 13565 14995
rect 13595 14965 13600 14995
rect 13560 14960 13600 14965
rect 13640 15155 13680 15160
rect 13640 15125 13645 15155
rect 13675 15125 13680 15155
rect 13640 14995 13680 15125
rect 13640 14965 13645 14995
rect 13675 14965 13680 14995
rect 13640 14960 13680 14965
rect 13720 15155 13760 15160
rect 13720 15125 13725 15155
rect 13755 15125 13760 15155
rect 13720 14995 13760 15125
rect 13720 14965 13725 14995
rect 13755 14965 13760 14995
rect 13720 14960 13760 14965
rect 13800 15155 13840 15160
rect 13800 15125 13805 15155
rect 13835 15125 13840 15155
rect 13800 14995 13840 15125
rect 13800 14965 13805 14995
rect 13835 14965 13840 14995
rect 13800 14960 13840 14965
rect 13880 15155 13920 15160
rect 13880 15125 13885 15155
rect 13915 15125 13920 15155
rect 13880 14995 13920 15125
rect 13880 14965 13885 14995
rect 13915 14965 13920 14995
rect 13880 14960 13920 14965
rect 13960 15155 14000 15160
rect 13960 15125 13965 15155
rect 13995 15125 14000 15155
rect 13960 14995 14000 15125
rect 13960 14965 13965 14995
rect 13995 14965 14000 14995
rect 13960 14960 14000 14965
rect 14040 15155 14080 15160
rect 14040 15125 14045 15155
rect 14075 15125 14080 15155
rect 14040 14995 14080 15125
rect 14040 14965 14045 14995
rect 14075 14965 14080 14995
rect 14040 14960 14080 14965
rect 14120 15155 14160 15160
rect 14120 15125 14125 15155
rect 14155 15125 14160 15155
rect 14120 14995 14160 15125
rect 14120 14965 14125 14995
rect 14155 14965 14160 14995
rect 14120 14960 14160 14965
rect 14200 15155 14240 15160
rect 14200 15125 14205 15155
rect 14235 15125 14240 15155
rect 14200 14995 14240 15125
rect 14200 14965 14205 14995
rect 14235 14965 14240 14995
rect 14200 14960 14240 14965
rect 14280 15155 14320 15160
rect 14280 15125 14285 15155
rect 14315 15125 14320 15155
rect 14280 14995 14320 15125
rect 14280 14965 14285 14995
rect 14315 14965 14320 14995
rect 14280 14960 14320 14965
rect 14360 15155 14400 15160
rect 14360 15125 14365 15155
rect 14395 15125 14400 15155
rect 14360 14995 14400 15125
rect 14360 14965 14365 14995
rect 14395 14965 14400 14995
rect 14360 14960 14400 14965
rect 14440 15155 14480 15160
rect 14440 15125 14445 15155
rect 14475 15125 14480 15155
rect 14440 14995 14480 15125
rect 14440 14965 14445 14995
rect 14475 14965 14480 14995
rect 14440 14960 14480 14965
rect 14520 15155 14560 15160
rect 14520 15125 14525 15155
rect 14555 15125 14560 15155
rect 14520 14995 14560 15125
rect 14520 14965 14525 14995
rect 14555 14965 14560 14995
rect 14520 14960 14560 14965
rect 14600 15155 14640 15160
rect 14600 15125 14605 15155
rect 14635 15125 14640 15155
rect 14600 14995 14640 15125
rect 14600 14965 14605 14995
rect 14635 14965 14640 14995
rect 14600 14960 14640 14965
rect 14680 15155 14720 15160
rect 14680 15125 14685 15155
rect 14715 15125 14720 15155
rect 14680 14995 14720 15125
rect 14680 14965 14685 14995
rect 14715 14965 14720 14995
rect 14680 14960 14720 14965
rect 11440 14885 11445 14915
rect 11475 14885 11480 14915
rect 11440 14755 11480 14885
rect 11440 14725 11445 14755
rect 11475 14725 11480 14755
rect 11440 14720 11480 14725
rect 11560 14915 11600 14920
rect 11560 14885 11565 14915
rect 11595 14885 11600 14915
rect 11560 14755 11600 14885
rect 11560 14725 11565 14755
rect 11595 14725 11600 14755
rect 11560 14720 11600 14725
rect 11640 14915 11680 14920
rect 11640 14885 11645 14915
rect 11675 14885 11680 14915
rect 11640 14755 11680 14885
rect 11640 14725 11645 14755
rect 11675 14725 11680 14755
rect 11640 14720 11680 14725
rect 11720 14915 11760 14920
rect 11720 14885 11725 14915
rect 11755 14885 11760 14915
rect 11720 14755 11760 14885
rect 11720 14725 11725 14755
rect 11755 14725 11760 14755
rect 11720 14720 11760 14725
rect 11800 14915 11840 14920
rect 11800 14885 11805 14915
rect 11835 14885 11840 14915
rect 11800 14755 11840 14885
rect 11800 14725 11805 14755
rect 11835 14725 11840 14755
rect 11800 14720 11840 14725
rect 11880 14915 11920 14920
rect 11880 14885 11885 14915
rect 11915 14885 11920 14915
rect 11880 14755 11920 14885
rect 11880 14725 11885 14755
rect 11915 14725 11920 14755
rect 11880 14720 11920 14725
rect 11960 14915 12000 14920
rect 11960 14885 11965 14915
rect 11995 14885 12000 14915
rect 11960 14755 12000 14885
rect 11960 14725 11965 14755
rect 11995 14725 12000 14755
rect 11960 14720 12000 14725
rect 12040 14915 12080 14920
rect 12040 14885 12045 14915
rect 12075 14885 12080 14915
rect 12040 14755 12080 14885
rect 12040 14725 12045 14755
rect 12075 14725 12080 14755
rect 12040 14720 12080 14725
rect 12120 14915 12160 14920
rect 12120 14885 12125 14915
rect 12155 14885 12160 14915
rect 12120 14755 12160 14885
rect 12120 14725 12125 14755
rect 12155 14725 12160 14755
rect 12120 14720 12160 14725
rect 12200 14915 12240 14920
rect 12200 14885 12205 14915
rect 12235 14885 12240 14915
rect 12200 14755 12240 14885
rect 12200 14725 12205 14755
rect 12235 14725 12240 14755
rect 12200 14720 12240 14725
rect 12280 14915 12320 14920
rect 12280 14885 12285 14915
rect 12315 14885 12320 14915
rect 12280 14755 12320 14885
rect 12280 14725 12285 14755
rect 12315 14725 12320 14755
rect 12280 14720 12320 14725
rect 12360 14915 12400 14920
rect 12360 14885 12365 14915
rect 12395 14885 12400 14915
rect 12360 14755 12400 14885
rect 12360 14725 12365 14755
rect 12395 14725 12400 14755
rect 12360 14720 12400 14725
rect 12440 14915 12480 14920
rect 12440 14885 12445 14915
rect 12475 14885 12480 14915
rect 12440 14755 12480 14885
rect 12440 14725 12445 14755
rect 12475 14725 12480 14755
rect 12440 14720 12480 14725
rect 12520 14915 12560 14920
rect 12520 14885 12525 14915
rect 12555 14885 12560 14915
rect 12520 14755 12560 14885
rect 12520 14725 12525 14755
rect 12555 14725 12560 14755
rect 12520 14720 12560 14725
rect 12600 14915 12640 14920
rect 12600 14885 12605 14915
rect 12635 14885 12640 14915
rect 12600 14755 12640 14885
rect 12600 14725 12605 14755
rect 12635 14725 12640 14755
rect 12600 14720 12640 14725
rect 12680 14915 12720 14920
rect 12680 14885 12685 14915
rect 12715 14885 12720 14915
rect 12680 14755 12720 14885
rect 12680 14725 12685 14755
rect 12715 14725 12720 14755
rect 12680 14720 12720 14725
rect 12760 14915 12800 14920
rect 12760 14885 12765 14915
rect 12795 14885 12800 14915
rect 12760 14755 12800 14885
rect 12760 14725 12765 14755
rect 12795 14725 12800 14755
rect 12760 14720 12800 14725
rect 12840 14915 12880 14920
rect 12840 14885 12845 14915
rect 12875 14885 12880 14915
rect 12840 14755 12880 14885
rect 12840 14725 12845 14755
rect 12875 14725 12880 14755
rect 12840 14720 12880 14725
rect 12920 14915 12960 14920
rect 12920 14885 12925 14915
rect 12955 14885 12960 14915
rect 12920 14755 12960 14885
rect 12920 14725 12925 14755
rect 12955 14725 12960 14755
rect 12920 14720 12960 14725
rect 13000 14915 13040 14920
rect 13000 14885 13005 14915
rect 13035 14885 13040 14915
rect 13000 14755 13040 14885
rect 13000 14725 13005 14755
rect 13035 14725 13040 14755
rect 13000 14720 13040 14725
rect 13080 14915 13120 14920
rect 13080 14885 13085 14915
rect 13115 14885 13120 14915
rect 13080 14755 13120 14885
rect 13080 14725 13085 14755
rect 13115 14725 13120 14755
rect 13080 14720 13120 14725
rect 13160 14915 13200 14920
rect 13160 14885 13165 14915
rect 13195 14885 13200 14915
rect 13160 14755 13200 14885
rect 13160 14725 13165 14755
rect 13195 14725 13200 14755
rect 13160 14720 13200 14725
rect 13240 14915 13280 14920
rect 13240 14885 13245 14915
rect 13275 14885 13280 14915
rect 13240 14755 13280 14885
rect 13240 14725 13245 14755
rect 13275 14725 13280 14755
rect 13240 14720 13280 14725
rect 13320 14915 13360 14920
rect 13320 14885 13325 14915
rect 13355 14885 13360 14915
rect 13320 14755 13360 14885
rect 13320 14725 13325 14755
rect 13355 14725 13360 14755
rect 13320 14720 13360 14725
rect 13400 14915 13440 14920
rect 13400 14885 13405 14915
rect 13435 14885 13440 14915
rect 13400 14755 13440 14885
rect 13400 14725 13405 14755
rect 13435 14725 13440 14755
rect 13400 14720 13440 14725
rect 13480 14915 13520 14920
rect 13480 14885 13485 14915
rect 13515 14885 13520 14915
rect 13480 14755 13520 14885
rect 13480 14725 13485 14755
rect 13515 14725 13520 14755
rect 13480 14720 13520 14725
rect 13560 14915 13600 14920
rect 13560 14885 13565 14915
rect 13595 14885 13600 14915
rect 13560 14755 13600 14885
rect 13560 14725 13565 14755
rect 13595 14725 13600 14755
rect 13560 14720 13600 14725
rect 13640 14915 13680 14920
rect 13640 14885 13645 14915
rect 13675 14885 13680 14915
rect 13640 14755 13680 14885
rect 13640 14725 13645 14755
rect 13675 14725 13680 14755
rect 13640 14720 13680 14725
rect 13720 14915 13760 14920
rect 13720 14885 13725 14915
rect 13755 14885 13760 14915
rect 13720 14755 13760 14885
rect 13720 14725 13725 14755
rect 13755 14725 13760 14755
rect 13720 14720 13760 14725
rect 13800 14915 13840 14920
rect 13800 14885 13805 14915
rect 13835 14885 13840 14915
rect 13800 14755 13840 14885
rect 13800 14725 13805 14755
rect 13835 14725 13840 14755
rect 13800 14720 13840 14725
rect 13880 14915 13920 14920
rect 13880 14885 13885 14915
rect 13915 14885 13920 14915
rect 13880 14755 13920 14885
rect 13880 14725 13885 14755
rect 13915 14725 13920 14755
rect 13880 14720 13920 14725
rect 13960 14915 14000 14920
rect 13960 14885 13965 14915
rect 13995 14885 14000 14915
rect 13960 14755 14000 14885
rect 13960 14725 13965 14755
rect 13995 14725 14000 14755
rect 13960 14720 14000 14725
rect 14040 14915 14080 14920
rect 14040 14885 14045 14915
rect 14075 14885 14080 14915
rect 14040 14755 14080 14885
rect 14040 14725 14045 14755
rect 14075 14725 14080 14755
rect 14040 14720 14080 14725
rect 14120 14915 14160 14920
rect 14120 14885 14125 14915
rect 14155 14885 14160 14915
rect 14120 14755 14160 14885
rect 14120 14725 14125 14755
rect 14155 14725 14160 14755
rect 14120 14720 14160 14725
rect 14200 14915 14240 14920
rect 14200 14885 14205 14915
rect 14235 14885 14240 14915
rect 14200 14755 14240 14885
rect 14200 14725 14205 14755
rect 14235 14725 14240 14755
rect 14200 14720 14240 14725
rect 14280 14915 14320 14920
rect 14280 14885 14285 14915
rect 14315 14885 14320 14915
rect 14280 14755 14320 14885
rect 14280 14725 14285 14755
rect 14315 14725 14320 14755
rect 14280 14720 14320 14725
rect 14360 14915 14400 14920
rect 14360 14885 14365 14915
rect 14395 14885 14400 14915
rect 14360 14755 14400 14885
rect 14360 14725 14365 14755
rect 14395 14725 14400 14755
rect 14360 14720 14400 14725
rect 14440 14915 14480 14920
rect 14440 14885 14445 14915
rect 14475 14885 14480 14915
rect 14440 14755 14480 14885
rect 14440 14725 14445 14755
rect 14475 14725 14480 14755
rect 14440 14720 14480 14725
rect 14520 14915 14560 14920
rect 14520 14885 14525 14915
rect 14555 14885 14560 14915
rect 14520 14755 14560 14885
rect 14520 14725 14525 14755
rect 14555 14725 14560 14755
rect 14520 14720 14560 14725
rect 14600 14915 14640 14920
rect 14600 14885 14605 14915
rect 14635 14885 14640 14915
rect 14600 14755 14640 14885
rect 14600 14725 14605 14755
rect 14635 14725 14640 14755
rect 14600 14720 14640 14725
rect 14680 14915 14720 14920
rect 14680 14885 14685 14915
rect 14715 14885 14720 14915
rect 14680 14755 14720 14885
rect 14680 14725 14685 14755
rect 14715 14725 14720 14755
rect 14680 14720 14720 14725
rect 14760 14915 14800 16680
rect 14760 14885 14765 14915
rect 14795 14885 14800 14915
rect 14760 14755 14800 14885
rect 14760 14725 14765 14755
rect 14795 14725 14800 14755
rect 14760 14680 14800 14725
rect 14840 14835 14880 16680
rect 14840 14805 14845 14835
rect 14875 14805 14880 14835
rect 14840 14680 14880 14805
rect 14920 14915 14960 16680
rect 14920 14885 14925 14915
rect 14955 14885 14960 14915
rect 14920 14755 14960 14885
rect 14920 14725 14925 14755
rect 14955 14725 14960 14755
rect 14920 14680 14960 14725
rect 15000 15155 15040 16680
rect 15000 15125 15005 15155
rect 15035 15125 15040 15155
rect 15000 14995 15040 15125
rect 15000 14965 15005 14995
rect 15035 14965 15040 14995
rect 15000 14680 15040 14965
rect 15080 15075 15120 16680
rect 15080 15045 15085 15075
rect 15115 15045 15120 15075
rect 15080 14680 15120 15045
rect 15160 15155 15200 16680
rect 15160 15125 15165 15155
rect 15195 15125 15200 15155
rect 15160 14995 15200 15125
rect 15160 14965 15165 14995
rect 15195 14965 15200 14995
rect 15160 14680 15200 14965
rect 15240 16195 15280 16680
rect 15240 16165 15245 16195
rect 15275 16165 15280 16195
rect 15240 16035 15280 16165
rect 15240 16005 15245 16035
rect 15275 16005 15280 16035
rect 15240 15875 15280 16005
rect 15240 15845 15245 15875
rect 15275 15845 15280 15875
rect 15240 15715 15280 15845
rect 15240 15685 15245 15715
rect 15275 15685 15280 15715
rect 15240 15555 15280 15685
rect 15240 15525 15245 15555
rect 15275 15525 15280 15555
rect 15240 15395 15280 15525
rect 15240 15365 15245 15395
rect 15275 15365 15280 15395
rect 15240 15235 15280 15365
rect 15240 15205 15245 15235
rect 15275 15205 15280 15235
rect 15240 14680 15280 15205
rect 15320 15315 15360 16680
rect 15320 15285 15325 15315
rect 15355 15285 15360 15315
rect 15320 14680 15360 15285
rect 15400 16195 15440 16680
rect 15400 16165 15405 16195
rect 15435 16165 15440 16195
rect 15400 16035 15440 16165
rect 15400 16005 15405 16035
rect 15435 16005 15440 16035
rect 15400 15875 15440 16005
rect 15400 15845 15405 15875
rect 15435 15845 15440 15875
rect 15400 15715 15440 15845
rect 15400 15685 15405 15715
rect 15435 15685 15440 15715
rect 15400 15555 15440 15685
rect 15400 15525 15405 15555
rect 15435 15525 15440 15555
rect 15400 15395 15440 15525
rect 15400 15365 15405 15395
rect 15435 15365 15440 15395
rect 15400 15235 15440 15365
rect 15400 15205 15405 15235
rect 15435 15205 15440 15235
rect 15400 14680 15440 15205
rect 15480 15475 15520 16680
rect 15480 15445 15485 15475
rect 15515 15445 15520 15475
rect 15480 14680 15520 15445
rect 15560 16195 15600 16680
rect 15560 16165 15565 16195
rect 15595 16165 15600 16195
rect 15560 16035 15600 16165
rect 15560 16005 15565 16035
rect 15595 16005 15600 16035
rect 15560 15875 15600 16005
rect 15560 15845 15565 15875
rect 15595 15845 15600 15875
rect 15560 15715 15600 15845
rect 15560 15685 15565 15715
rect 15595 15685 15600 15715
rect 15560 15555 15600 15685
rect 15560 15525 15565 15555
rect 15595 15525 15600 15555
rect 15560 15395 15600 15525
rect 15560 15365 15565 15395
rect 15595 15365 15600 15395
rect 15560 15235 15600 15365
rect 15560 15205 15565 15235
rect 15595 15205 15600 15235
rect 15560 14680 15600 15205
rect 15640 15635 15680 16680
rect 15640 15605 15645 15635
rect 15675 15605 15680 15635
rect 15640 14680 15680 15605
rect 15720 16195 15760 16680
rect 15720 16165 15725 16195
rect 15755 16165 15760 16195
rect 15720 16035 15760 16165
rect 15720 16005 15725 16035
rect 15755 16005 15760 16035
rect 15720 15875 15760 16005
rect 15720 15845 15725 15875
rect 15755 15845 15760 15875
rect 15720 15715 15760 15845
rect 15720 15685 15725 15715
rect 15755 15685 15760 15715
rect 15720 15555 15760 15685
rect 15720 15525 15725 15555
rect 15755 15525 15760 15555
rect 15720 15395 15760 15525
rect 15720 15365 15725 15395
rect 15755 15365 15760 15395
rect 15720 15235 15760 15365
rect 15720 15205 15725 15235
rect 15755 15205 15760 15235
rect 15720 14680 15760 15205
rect 15800 15795 15840 16680
rect 15800 15765 15805 15795
rect 15835 15765 15840 15795
rect 15800 14680 15840 15765
rect 15880 16195 15920 16680
rect 15880 16165 15885 16195
rect 15915 16165 15920 16195
rect 15880 16035 15920 16165
rect 15880 16005 15885 16035
rect 15915 16005 15920 16035
rect 15880 15875 15920 16005
rect 15880 15845 15885 15875
rect 15915 15845 15920 15875
rect 15880 15715 15920 15845
rect 15880 15685 15885 15715
rect 15915 15685 15920 15715
rect 15880 15555 15920 15685
rect 15880 15525 15885 15555
rect 15915 15525 15920 15555
rect 15880 15395 15920 15525
rect 15880 15365 15885 15395
rect 15915 15365 15920 15395
rect 15880 15235 15920 15365
rect 15880 15205 15885 15235
rect 15915 15205 15920 15235
rect 15880 14680 15920 15205
rect 15960 15955 16000 16680
rect 15960 15925 15965 15955
rect 15995 15925 16000 15955
rect 15960 14680 16000 15925
rect 16040 16195 16080 16680
rect 16040 16165 16045 16195
rect 16075 16165 16080 16195
rect 16040 16035 16080 16165
rect 16040 16005 16045 16035
rect 16075 16005 16080 16035
rect 16040 15875 16080 16005
rect 16040 15845 16045 15875
rect 16075 15845 16080 15875
rect 16040 15715 16080 15845
rect 16040 15685 16045 15715
rect 16075 15685 16080 15715
rect 16040 15555 16080 15685
rect 16040 15525 16045 15555
rect 16075 15525 16080 15555
rect 16040 15395 16080 15525
rect 16040 15365 16045 15395
rect 16075 15365 16080 15395
rect 16040 15235 16080 15365
rect 16040 15205 16045 15235
rect 16075 15205 16080 15235
rect 16040 14680 16080 15205
rect 16120 16115 16160 16680
rect 16120 16085 16125 16115
rect 16155 16085 16160 16115
rect 16120 14680 16160 16085
rect 16200 16195 16240 16680
rect 16200 16165 16205 16195
rect 16235 16165 16240 16195
rect 16200 16035 16240 16165
rect 16200 16005 16205 16035
rect 16235 16005 16240 16035
rect 16200 15875 16240 16005
rect 16200 15845 16205 15875
rect 16235 15845 16240 15875
rect 16200 15715 16240 15845
rect 16200 15685 16205 15715
rect 16235 15685 16240 15715
rect 16200 15555 16240 15685
rect 16200 15525 16205 15555
rect 16235 15525 16240 15555
rect 16200 15395 16240 15525
rect 16200 15365 16205 15395
rect 16235 15365 16240 15395
rect 16200 15235 16240 15365
rect 16200 15205 16205 15235
rect 16235 15205 16240 15235
rect 16200 14680 16240 15205
rect 16280 16435 16320 16680
rect 16280 16405 16285 16435
rect 16315 16405 16320 16435
rect 16280 16275 16320 16405
rect 16280 16245 16285 16275
rect 16315 16245 16320 16275
rect 16280 14680 16320 16245
rect 16360 16355 16400 16680
rect 16360 16325 16365 16355
rect 16395 16325 16400 16355
rect 16360 14680 16400 16325
rect 16440 16435 16480 16680
rect 16440 16405 16445 16435
rect 16475 16405 16480 16435
rect 16440 16275 16480 16405
rect 16440 16245 16445 16275
rect 16475 16245 16480 16275
rect 16440 14680 16480 16245
rect 16520 16675 16560 16680
rect 16520 16645 16525 16675
rect 16555 16645 16560 16675
rect 16520 16515 16560 16645
rect 16520 16485 16525 16515
rect 16555 16485 16560 16515
rect 16520 14680 16560 16485
rect 16600 16595 16640 16680
rect 16600 16565 16605 16595
rect 16635 16565 16640 16595
rect 16600 14680 16640 16565
rect 16680 16675 16720 16680
rect 16680 16645 16685 16675
rect 16715 16645 16720 16675
rect 16680 16515 16720 16645
rect 16680 16485 16685 16515
rect 16715 16485 16720 16515
rect 16680 14680 16720 16485
rect 16760 16675 16800 16680
rect 16760 16645 16765 16675
rect 16795 16645 16800 16675
rect 16760 16515 16800 16645
rect 16760 16485 16765 16515
rect 16795 16485 16800 16515
rect 16760 16480 16800 16485
rect 16840 16675 16880 16680
rect 16840 16645 16845 16675
rect 16875 16645 16880 16675
rect 16840 16515 16880 16645
rect 16840 16485 16845 16515
rect 16875 16485 16880 16515
rect 16840 16480 16880 16485
rect 16920 16675 16960 16680
rect 16920 16645 16925 16675
rect 16955 16645 16960 16675
rect 16920 16515 16960 16645
rect 16920 16485 16925 16515
rect 16955 16485 16960 16515
rect 16920 16480 16960 16485
rect 17000 16675 17040 16680
rect 17000 16645 17005 16675
rect 17035 16645 17040 16675
rect 17000 16515 17040 16645
rect 17000 16485 17005 16515
rect 17035 16485 17040 16515
rect 17000 16480 17040 16485
rect 17080 16675 17120 16680
rect 17080 16645 17085 16675
rect 17115 16645 17120 16675
rect 17080 16515 17120 16645
rect 17080 16485 17085 16515
rect 17115 16485 17120 16515
rect 17080 16480 17120 16485
rect 17160 16675 17200 16680
rect 17160 16645 17165 16675
rect 17195 16645 17200 16675
rect 17160 16515 17200 16645
rect 17160 16485 17165 16515
rect 17195 16485 17200 16515
rect 17160 16480 17200 16485
rect 17240 16675 17280 16680
rect 17240 16645 17245 16675
rect 17275 16645 17280 16675
rect 17240 16515 17280 16645
rect 17240 16485 17245 16515
rect 17275 16485 17280 16515
rect 17240 16480 17280 16485
rect 17320 16675 17360 16680
rect 17320 16645 17325 16675
rect 17355 16645 17360 16675
rect 17320 16515 17360 16645
rect 17320 16485 17325 16515
rect 17355 16485 17360 16515
rect 17320 16480 17360 16485
rect 17400 16675 17440 16680
rect 17400 16645 17405 16675
rect 17435 16645 17440 16675
rect 17400 16515 17440 16645
rect 17400 16485 17405 16515
rect 17435 16485 17440 16515
rect 17400 16480 17440 16485
rect 17480 16675 17520 16680
rect 17480 16645 17485 16675
rect 17515 16645 17520 16675
rect 17480 16515 17520 16645
rect 17480 16485 17485 16515
rect 17515 16485 17520 16515
rect 17480 16480 17520 16485
rect 17560 16675 17600 16680
rect 17560 16645 17565 16675
rect 17595 16645 17600 16675
rect 17560 16515 17600 16645
rect 17560 16485 17565 16515
rect 17595 16485 17600 16515
rect 17560 16480 17600 16485
rect 17640 16675 17680 16680
rect 17640 16645 17645 16675
rect 17675 16645 17680 16675
rect 17640 16515 17680 16645
rect 17640 16485 17645 16515
rect 17675 16485 17680 16515
rect 17640 16480 17680 16485
rect 17720 16675 17760 16680
rect 17720 16645 17725 16675
rect 17755 16645 17760 16675
rect 17720 16515 17760 16645
rect 17720 16485 17725 16515
rect 17755 16485 17760 16515
rect 17720 16480 17760 16485
rect 17800 16675 17840 16680
rect 17800 16645 17805 16675
rect 17835 16645 17840 16675
rect 17800 16515 17840 16645
rect 17800 16485 17805 16515
rect 17835 16485 17840 16515
rect 17800 16480 17840 16485
rect 17880 16675 17920 16680
rect 17880 16645 17885 16675
rect 17915 16645 17920 16675
rect 17880 16515 17920 16645
rect 17880 16485 17885 16515
rect 17915 16485 17920 16515
rect 17880 16480 17920 16485
rect 17960 16675 18000 16680
rect 17960 16645 17965 16675
rect 17995 16645 18000 16675
rect 17960 16515 18000 16645
rect 17960 16485 17965 16515
rect 17995 16485 18000 16515
rect 17960 16480 18000 16485
rect 18040 16675 18080 16680
rect 18040 16645 18045 16675
rect 18075 16645 18080 16675
rect 18040 16515 18080 16645
rect 18040 16485 18045 16515
rect 18075 16485 18080 16515
rect 18040 16480 18080 16485
rect 18120 16675 18160 16680
rect 18120 16645 18125 16675
rect 18155 16645 18160 16675
rect 18120 16515 18160 16645
rect 18120 16485 18125 16515
rect 18155 16485 18160 16515
rect 18120 16480 18160 16485
rect 18200 16675 18240 16680
rect 18200 16645 18205 16675
rect 18235 16645 18240 16675
rect 18200 16515 18240 16645
rect 18200 16485 18205 16515
rect 18235 16485 18240 16515
rect 18200 16480 18240 16485
rect 18280 16675 18320 16680
rect 18280 16645 18285 16675
rect 18315 16645 18320 16675
rect 18280 16515 18320 16645
rect 18280 16485 18285 16515
rect 18315 16485 18320 16515
rect 18280 16480 18320 16485
rect 18360 16675 18400 16680
rect 18360 16645 18365 16675
rect 18395 16645 18400 16675
rect 18360 16515 18400 16645
rect 18360 16485 18365 16515
rect 18395 16485 18400 16515
rect 18360 16480 18400 16485
rect 18440 16675 18480 16680
rect 18440 16645 18445 16675
rect 18475 16645 18480 16675
rect 18440 16515 18480 16645
rect 18440 16485 18445 16515
rect 18475 16485 18480 16515
rect 18440 16480 18480 16485
rect 18520 16675 18560 16680
rect 18520 16645 18525 16675
rect 18555 16645 18560 16675
rect 18520 16515 18560 16645
rect 18520 16485 18525 16515
rect 18555 16485 18560 16515
rect 18520 16480 18560 16485
rect 18600 16675 18640 16680
rect 18600 16645 18605 16675
rect 18635 16645 18640 16675
rect 18600 16515 18640 16645
rect 18600 16485 18605 16515
rect 18635 16485 18640 16515
rect 18600 16480 18640 16485
rect 18680 16675 18720 16680
rect 18680 16645 18685 16675
rect 18715 16645 18720 16675
rect 18680 16515 18720 16645
rect 18680 16485 18685 16515
rect 18715 16485 18720 16515
rect 18680 16480 18720 16485
rect 18760 16675 18800 16680
rect 18760 16645 18765 16675
rect 18795 16645 18800 16675
rect 18760 16515 18800 16645
rect 18760 16485 18765 16515
rect 18795 16485 18800 16515
rect 18760 16480 18800 16485
rect 18840 16675 18880 16680
rect 18840 16645 18845 16675
rect 18875 16645 18880 16675
rect 18840 16515 18880 16645
rect 18840 16485 18845 16515
rect 18875 16485 18880 16515
rect 18840 16480 18880 16485
rect 18920 16675 18960 16680
rect 18920 16645 18925 16675
rect 18955 16645 18960 16675
rect 18920 16515 18960 16645
rect 18920 16485 18925 16515
rect 18955 16485 18960 16515
rect 18920 16480 18960 16485
rect 19000 16675 19040 16680
rect 19000 16645 19005 16675
rect 19035 16645 19040 16675
rect 19000 16515 19040 16645
rect 19000 16485 19005 16515
rect 19035 16485 19040 16515
rect 19000 16480 19040 16485
rect 19080 16675 19120 16680
rect 19080 16645 19085 16675
rect 19115 16645 19120 16675
rect 19080 16515 19120 16645
rect 19080 16485 19085 16515
rect 19115 16485 19120 16515
rect 19080 16480 19120 16485
rect 19160 16675 19200 16680
rect 19160 16645 19165 16675
rect 19195 16645 19200 16675
rect 19160 16515 19200 16645
rect 19160 16485 19165 16515
rect 19195 16485 19200 16515
rect 19160 16480 19200 16485
rect 19240 16675 19280 16680
rect 19240 16645 19245 16675
rect 19275 16645 19280 16675
rect 19240 16515 19280 16645
rect 19240 16485 19245 16515
rect 19275 16485 19280 16515
rect 19240 16480 19280 16485
rect 19320 16675 19360 16680
rect 19320 16645 19325 16675
rect 19355 16645 19360 16675
rect 19320 16515 19360 16645
rect 19320 16485 19325 16515
rect 19355 16485 19360 16515
rect 19320 16480 19360 16485
rect 19400 16675 19440 16680
rect 19400 16645 19405 16675
rect 19435 16645 19440 16675
rect 19400 16515 19440 16645
rect 19400 16485 19405 16515
rect 19435 16485 19440 16515
rect 19400 16480 19440 16485
rect 19480 16675 19520 16680
rect 19480 16645 19485 16675
rect 19515 16645 19520 16675
rect 19480 16515 19520 16645
rect 19480 16485 19485 16515
rect 19515 16485 19520 16515
rect 19480 16480 19520 16485
rect 19560 16675 19600 16680
rect 19560 16645 19565 16675
rect 19595 16645 19600 16675
rect 19560 16515 19600 16645
rect 19560 16485 19565 16515
rect 19595 16485 19600 16515
rect 19560 16480 19600 16485
rect 19640 16675 19680 16680
rect 19640 16645 19645 16675
rect 19675 16645 19680 16675
rect 19640 16515 19680 16645
rect 19640 16485 19645 16515
rect 19675 16485 19680 16515
rect 19640 16480 19680 16485
rect 19720 16675 19760 16680
rect 19720 16645 19725 16675
rect 19755 16645 19760 16675
rect 19720 16515 19760 16645
rect 19720 16485 19725 16515
rect 19755 16485 19760 16515
rect 19720 16480 19760 16485
rect 19800 16675 19840 16680
rect 19800 16645 19805 16675
rect 19835 16645 19840 16675
rect 19800 16515 19840 16645
rect 19800 16485 19805 16515
rect 19835 16485 19840 16515
rect 19800 16480 19840 16485
rect 19880 16675 19920 16680
rect 19880 16645 19885 16675
rect 19915 16645 19920 16675
rect 19880 16515 19920 16645
rect 19880 16485 19885 16515
rect 19915 16485 19920 16515
rect 19880 16480 19920 16485
rect 19960 16675 20000 16680
rect 19960 16645 19965 16675
rect 19995 16645 20000 16675
rect 19960 16515 20000 16645
rect 19960 16485 19965 16515
rect 19995 16485 20000 16515
rect 19960 16480 20000 16485
rect 20040 16675 20080 16680
rect 20040 16645 20045 16675
rect 20075 16645 20080 16675
rect 20040 16515 20080 16645
rect 20040 16485 20045 16515
rect 20075 16485 20080 16515
rect 20040 16480 20080 16485
rect 20120 16675 20160 16680
rect 20120 16645 20125 16675
rect 20155 16645 20160 16675
rect 20120 16515 20160 16645
rect 20120 16485 20125 16515
rect 20155 16485 20160 16515
rect 20120 16480 20160 16485
rect 20200 16675 20240 16680
rect 20200 16645 20205 16675
rect 20235 16645 20240 16675
rect 20200 16515 20240 16645
rect 20200 16485 20205 16515
rect 20235 16485 20240 16515
rect 20200 16480 20240 16485
rect 20280 16675 20320 16680
rect 20280 16645 20285 16675
rect 20315 16645 20320 16675
rect 20280 16515 20320 16645
rect 20280 16485 20285 16515
rect 20315 16485 20320 16515
rect 20280 16480 20320 16485
rect 20360 16675 20400 16680
rect 20360 16645 20365 16675
rect 20395 16645 20400 16675
rect 20360 16515 20400 16645
rect 20360 16485 20365 16515
rect 20395 16485 20400 16515
rect 20360 16480 20400 16485
rect 20440 16675 20480 16680
rect 20440 16645 20445 16675
rect 20475 16645 20480 16675
rect 20440 16515 20480 16645
rect 20440 16485 20445 16515
rect 20475 16485 20480 16515
rect 20440 16480 20480 16485
rect 20520 16675 20560 16680
rect 20520 16645 20525 16675
rect 20555 16645 20560 16675
rect 20520 16515 20560 16645
rect 20520 16485 20525 16515
rect 20555 16485 20560 16515
rect 20520 16480 20560 16485
rect 20600 16675 20640 16680
rect 20600 16645 20605 16675
rect 20635 16645 20640 16675
rect 20600 16515 20640 16645
rect 20600 16485 20605 16515
rect 20635 16485 20640 16515
rect 20600 16480 20640 16485
rect 20680 16675 20720 16680
rect 20680 16645 20685 16675
rect 20715 16645 20720 16675
rect 20680 16515 20720 16645
rect 20680 16485 20685 16515
rect 20715 16485 20720 16515
rect 20680 16480 20720 16485
rect 20760 16675 20800 16680
rect 20760 16645 20765 16675
rect 20795 16645 20800 16675
rect 20760 16515 20800 16645
rect 20760 16485 20765 16515
rect 20795 16485 20800 16515
rect 20760 16480 20800 16485
rect 20840 16675 20880 16680
rect 20840 16645 20845 16675
rect 20875 16645 20880 16675
rect 20840 16515 20880 16645
rect 20840 16485 20845 16515
rect 20875 16485 20880 16515
rect 20840 16480 20880 16485
rect 20920 16675 20960 16680
rect 20920 16645 20925 16675
rect 20955 16645 20960 16675
rect 20920 16515 20960 16645
rect 20920 16485 20925 16515
rect 20955 16485 20960 16515
rect 20920 16480 20960 16485
rect 16760 16435 16800 16440
rect 16760 16405 16765 16435
rect 16795 16405 16800 16435
rect 16760 16275 16800 16405
rect 16760 16245 16765 16275
rect 16795 16245 16800 16275
rect 16760 16240 16800 16245
rect 16840 16435 16880 16440
rect 16840 16405 16845 16435
rect 16875 16405 16880 16435
rect 16840 16275 16880 16405
rect 16840 16245 16845 16275
rect 16875 16245 16880 16275
rect 16840 16240 16880 16245
rect 16920 16435 16960 16440
rect 16920 16405 16925 16435
rect 16955 16405 16960 16435
rect 16920 16275 16960 16405
rect 16920 16245 16925 16275
rect 16955 16245 16960 16275
rect 16920 16240 16960 16245
rect 17000 16435 17040 16440
rect 17000 16405 17005 16435
rect 17035 16405 17040 16435
rect 17000 16275 17040 16405
rect 17000 16245 17005 16275
rect 17035 16245 17040 16275
rect 17000 16240 17040 16245
rect 17080 16435 17120 16440
rect 17080 16405 17085 16435
rect 17115 16405 17120 16435
rect 17080 16275 17120 16405
rect 17080 16245 17085 16275
rect 17115 16245 17120 16275
rect 17080 16240 17120 16245
rect 17160 16435 17200 16440
rect 17160 16405 17165 16435
rect 17195 16405 17200 16435
rect 17160 16275 17200 16405
rect 17160 16245 17165 16275
rect 17195 16245 17200 16275
rect 17160 16240 17200 16245
rect 17240 16435 17280 16440
rect 17240 16405 17245 16435
rect 17275 16405 17280 16435
rect 17240 16275 17280 16405
rect 17240 16245 17245 16275
rect 17275 16245 17280 16275
rect 17240 16240 17280 16245
rect 17320 16435 17360 16440
rect 17320 16405 17325 16435
rect 17355 16405 17360 16435
rect 17320 16275 17360 16405
rect 17320 16245 17325 16275
rect 17355 16245 17360 16275
rect 17320 16240 17360 16245
rect 17400 16435 17440 16440
rect 17400 16405 17405 16435
rect 17435 16405 17440 16435
rect 17400 16275 17440 16405
rect 17400 16245 17405 16275
rect 17435 16245 17440 16275
rect 17400 16240 17440 16245
rect 17480 16435 17520 16440
rect 17480 16405 17485 16435
rect 17515 16405 17520 16435
rect 17480 16275 17520 16405
rect 17480 16245 17485 16275
rect 17515 16245 17520 16275
rect 17480 16240 17520 16245
rect 17560 16435 17600 16440
rect 17560 16405 17565 16435
rect 17595 16405 17600 16435
rect 17560 16275 17600 16405
rect 17560 16245 17565 16275
rect 17595 16245 17600 16275
rect 17560 16240 17600 16245
rect 17640 16435 17680 16440
rect 17640 16405 17645 16435
rect 17675 16405 17680 16435
rect 17640 16275 17680 16405
rect 17640 16245 17645 16275
rect 17675 16245 17680 16275
rect 17640 16240 17680 16245
rect 17720 16435 17760 16440
rect 17720 16405 17725 16435
rect 17755 16405 17760 16435
rect 17720 16275 17760 16405
rect 17720 16245 17725 16275
rect 17755 16245 17760 16275
rect 17720 16240 17760 16245
rect 17800 16435 17840 16440
rect 17800 16405 17805 16435
rect 17835 16405 17840 16435
rect 17800 16275 17840 16405
rect 17800 16245 17805 16275
rect 17835 16245 17840 16275
rect 17800 16240 17840 16245
rect 17880 16435 17920 16440
rect 17880 16405 17885 16435
rect 17915 16405 17920 16435
rect 17880 16275 17920 16405
rect 17880 16245 17885 16275
rect 17915 16245 17920 16275
rect 17880 16240 17920 16245
rect 17960 16435 18000 16440
rect 17960 16405 17965 16435
rect 17995 16405 18000 16435
rect 17960 16275 18000 16405
rect 17960 16245 17965 16275
rect 17995 16245 18000 16275
rect 17960 16240 18000 16245
rect 18040 16435 18080 16440
rect 18040 16405 18045 16435
rect 18075 16405 18080 16435
rect 18040 16275 18080 16405
rect 18040 16245 18045 16275
rect 18075 16245 18080 16275
rect 18040 16240 18080 16245
rect 18120 16435 18160 16440
rect 18120 16405 18125 16435
rect 18155 16405 18160 16435
rect 18120 16275 18160 16405
rect 18120 16245 18125 16275
rect 18155 16245 18160 16275
rect 18120 16240 18160 16245
rect 18200 16435 18240 16440
rect 18200 16405 18205 16435
rect 18235 16405 18240 16435
rect 18200 16275 18240 16405
rect 18200 16245 18205 16275
rect 18235 16245 18240 16275
rect 18200 16240 18240 16245
rect 18280 16435 18320 16440
rect 18280 16405 18285 16435
rect 18315 16405 18320 16435
rect 18280 16275 18320 16405
rect 18280 16245 18285 16275
rect 18315 16245 18320 16275
rect 18280 16240 18320 16245
rect 18360 16435 18400 16440
rect 18360 16405 18365 16435
rect 18395 16405 18400 16435
rect 18360 16275 18400 16405
rect 18360 16245 18365 16275
rect 18395 16245 18400 16275
rect 18360 16240 18400 16245
rect 18440 16435 18480 16440
rect 18440 16405 18445 16435
rect 18475 16405 18480 16435
rect 18440 16275 18480 16405
rect 18440 16245 18445 16275
rect 18475 16245 18480 16275
rect 18440 16240 18480 16245
rect 18520 16435 18560 16440
rect 18520 16405 18525 16435
rect 18555 16405 18560 16435
rect 18520 16275 18560 16405
rect 18520 16245 18525 16275
rect 18555 16245 18560 16275
rect 18520 16240 18560 16245
rect 18600 16435 18640 16440
rect 18600 16405 18605 16435
rect 18635 16405 18640 16435
rect 18600 16275 18640 16405
rect 18600 16245 18605 16275
rect 18635 16245 18640 16275
rect 18600 16240 18640 16245
rect 18680 16435 18720 16440
rect 18680 16405 18685 16435
rect 18715 16405 18720 16435
rect 18680 16275 18720 16405
rect 18680 16245 18685 16275
rect 18715 16245 18720 16275
rect 18680 16240 18720 16245
rect 18760 16435 18800 16440
rect 18760 16405 18765 16435
rect 18795 16405 18800 16435
rect 18760 16275 18800 16405
rect 18760 16245 18765 16275
rect 18795 16245 18800 16275
rect 18760 16240 18800 16245
rect 18840 16435 18880 16440
rect 18840 16405 18845 16435
rect 18875 16405 18880 16435
rect 18840 16275 18880 16405
rect 18840 16245 18845 16275
rect 18875 16245 18880 16275
rect 18840 16240 18880 16245
rect 18920 16435 18960 16440
rect 18920 16405 18925 16435
rect 18955 16405 18960 16435
rect 18920 16275 18960 16405
rect 18920 16245 18925 16275
rect 18955 16245 18960 16275
rect 18920 16240 18960 16245
rect 19000 16435 19040 16440
rect 19000 16405 19005 16435
rect 19035 16405 19040 16435
rect 19000 16275 19040 16405
rect 19000 16245 19005 16275
rect 19035 16245 19040 16275
rect 19000 16240 19040 16245
rect 19080 16435 19120 16440
rect 19080 16405 19085 16435
rect 19115 16405 19120 16435
rect 19080 16275 19120 16405
rect 19080 16245 19085 16275
rect 19115 16245 19120 16275
rect 19080 16240 19120 16245
rect 19160 16435 19200 16440
rect 19160 16405 19165 16435
rect 19195 16405 19200 16435
rect 19160 16275 19200 16405
rect 19160 16245 19165 16275
rect 19195 16245 19200 16275
rect 19160 16240 19200 16245
rect 19240 16435 19280 16440
rect 19240 16405 19245 16435
rect 19275 16405 19280 16435
rect 19240 16275 19280 16405
rect 19240 16245 19245 16275
rect 19275 16245 19280 16275
rect 19240 16240 19280 16245
rect 19320 16435 19360 16440
rect 19320 16405 19325 16435
rect 19355 16405 19360 16435
rect 19320 16275 19360 16405
rect 19320 16245 19325 16275
rect 19355 16245 19360 16275
rect 19320 16240 19360 16245
rect 19400 16435 19440 16440
rect 19400 16405 19405 16435
rect 19435 16405 19440 16435
rect 19400 16275 19440 16405
rect 19400 16245 19405 16275
rect 19435 16245 19440 16275
rect 19400 16240 19440 16245
rect 19480 16435 19520 16440
rect 19480 16405 19485 16435
rect 19515 16405 19520 16435
rect 19480 16275 19520 16405
rect 19480 16245 19485 16275
rect 19515 16245 19520 16275
rect 19480 16240 19520 16245
rect 19560 16435 19600 16440
rect 19560 16405 19565 16435
rect 19595 16405 19600 16435
rect 19560 16275 19600 16405
rect 19560 16245 19565 16275
rect 19595 16245 19600 16275
rect 19560 16240 19600 16245
rect 19640 16435 19680 16440
rect 19640 16405 19645 16435
rect 19675 16405 19680 16435
rect 19640 16275 19680 16405
rect 19640 16245 19645 16275
rect 19675 16245 19680 16275
rect 19640 16240 19680 16245
rect 19720 16435 19760 16440
rect 19720 16405 19725 16435
rect 19755 16405 19760 16435
rect 19720 16275 19760 16405
rect 19720 16245 19725 16275
rect 19755 16245 19760 16275
rect 19720 16240 19760 16245
rect 19800 16435 19840 16440
rect 19800 16405 19805 16435
rect 19835 16405 19840 16435
rect 19800 16275 19840 16405
rect 19800 16245 19805 16275
rect 19835 16245 19840 16275
rect 19800 16240 19840 16245
rect 19880 16435 19920 16440
rect 19880 16405 19885 16435
rect 19915 16405 19920 16435
rect 19880 16275 19920 16405
rect 19880 16245 19885 16275
rect 19915 16245 19920 16275
rect 19880 16240 19920 16245
rect 19960 16435 20000 16440
rect 19960 16405 19965 16435
rect 19995 16405 20000 16435
rect 19960 16275 20000 16405
rect 19960 16245 19965 16275
rect 19995 16245 20000 16275
rect 19960 16240 20000 16245
rect 20040 16435 20080 16440
rect 20040 16405 20045 16435
rect 20075 16405 20080 16435
rect 20040 16275 20080 16405
rect 20040 16245 20045 16275
rect 20075 16245 20080 16275
rect 20040 16240 20080 16245
rect 20120 16435 20160 16440
rect 20120 16405 20125 16435
rect 20155 16405 20160 16435
rect 20120 16275 20160 16405
rect 20120 16245 20125 16275
rect 20155 16245 20160 16275
rect 20120 16240 20160 16245
rect 20200 16435 20240 16440
rect 20200 16405 20205 16435
rect 20235 16405 20240 16435
rect 20200 16275 20240 16405
rect 20200 16245 20205 16275
rect 20235 16245 20240 16275
rect 20200 16240 20240 16245
rect 20280 16435 20320 16440
rect 20280 16405 20285 16435
rect 20315 16405 20320 16435
rect 20280 16275 20320 16405
rect 20280 16245 20285 16275
rect 20315 16245 20320 16275
rect 20280 16240 20320 16245
rect 20360 16435 20400 16440
rect 20360 16405 20365 16435
rect 20395 16405 20400 16435
rect 20360 16275 20400 16405
rect 20360 16245 20365 16275
rect 20395 16245 20400 16275
rect 20360 16240 20400 16245
rect 20440 16435 20480 16440
rect 20440 16405 20445 16435
rect 20475 16405 20480 16435
rect 20440 16275 20480 16405
rect 20440 16245 20445 16275
rect 20475 16245 20480 16275
rect 20440 16240 20480 16245
rect 20520 16435 20560 16440
rect 20520 16405 20525 16435
rect 20555 16405 20560 16435
rect 20520 16275 20560 16405
rect 20520 16245 20525 16275
rect 20555 16245 20560 16275
rect 20520 16240 20560 16245
rect 20600 16435 20640 16440
rect 20600 16405 20605 16435
rect 20635 16405 20640 16435
rect 20600 16275 20640 16405
rect 20600 16245 20605 16275
rect 20635 16245 20640 16275
rect 20600 16240 20640 16245
rect 20680 16435 20720 16440
rect 20680 16405 20685 16435
rect 20715 16405 20720 16435
rect 20680 16275 20720 16405
rect 20680 16245 20685 16275
rect 20715 16245 20720 16275
rect 20680 16240 20720 16245
rect 20760 16435 20800 16440
rect 20760 16405 20765 16435
rect 20795 16405 20800 16435
rect 20760 16275 20800 16405
rect 20760 16245 20765 16275
rect 20795 16245 20800 16275
rect 20760 16240 20800 16245
rect 20840 16435 20880 16440
rect 20840 16405 20845 16435
rect 20875 16405 20880 16435
rect 20840 16275 20880 16405
rect 20840 16245 20845 16275
rect 20875 16245 20880 16275
rect 20840 16240 20880 16245
rect 20920 16435 20960 16440
rect 20920 16405 20925 16435
rect 20955 16405 20960 16435
rect 20920 16275 20960 16405
rect 20920 16245 20925 16275
rect 20955 16245 20960 16275
rect 20920 16240 20960 16245
rect 16760 16195 16800 16200
rect 16760 16165 16765 16195
rect 16795 16165 16800 16195
rect 16760 16035 16800 16165
rect 16760 16005 16765 16035
rect 16795 16005 16800 16035
rect 16760 15875 16800 16005
rect 16760 15845 16765 15875
rect 16795 15845 16800 15875
rect 16760 15715 16800 15845
rect 16760 15685 16765 15715
rect 16795 15685 16800 15715
rect 16760 15555 16800 15685
rect 16760 15525 16765 15555
rect 16795 15525 16800 15555
rect 16760 15395 16800 15525
rect 16760 15365 16765 15395
rect 16795 15365 16800 15395
rect 16760 15235 16800 15365
rect 16760 15205 16765 15235
rect 16795 15205 16800 15235
rect 16760 15200 16800 15205
rect 16840 16195 16880 16200
rect 16840 16165 16845 16195
rect 16875 16165 16880 16195
rect 16840 16035 16880 16165
rect 16840 16005 16845 16035
rect 16875 16005 16880 16035
rect 16840 15875 16880 16005
rect 16840 15845 16845 15875
rect 16875 15845 16880 15875
rect 16840 15715 16880 15845
rect 16840 15685 16845 15715
rect 16875 15685 16880 15715
rect 16840 15555 16880 15685
rect 16840 15525 16845 15555
rect 16875 15525 16880 15555
rect 16840 15395 16880 15525
rect 16840 15365 16845 15395
rect 16875 15365 16880 15395
rect 16840 15235 16880 15365
rect 16840 15205 16845 15235
rect 16875 15205 16880 15235
rect 16840 15200 16880 15205
rect 16920 16195 16960 16200
rect 16920 16165 16925 16195
rect 16955 16165 16960 16195
rect 16920 16035 16960 16165
rect 16920 16005 16925 16035
rect 16955 16005 16960 16035
rect 16920 15875 16960 16005
rect 16920 15845 16925 15875
rect 16955 15845 16960 15875
rect 16920 15715 16960 15845
rect 16920 15685 16925 15715
rect 16955 15685 16960 15715
rect 16920 15555 16960 15685
rect 16920 15525 16925 15555
rect 16955 15525 16960 15555
rect 16920 15395 16960 15525
rect 16920 15365 16925 15395
rect 16955 15365 16960 15395
rect 16920 15235 16960 15365
rect 16920 15205 16925 15235
rect 16955 15205 16960 15235
rect 16920 15200 16960 15205
rect 17000 16195 17040 16200
rect 17000 16165 17005 16195
rect 17035 16165 17040 16195
rect 17000 16035 17040 16165
rect 17000 16005 17005 16035
rect 17035 16005 17040 16035
rect 17000 15875 17040 16005
rect 17000 15845 17005 15875
rect 17035 15845 17040 15875
rect 17000 15715 17040 15845
rect 17000 15685 17005 15715
rect 17035 15685 17040 15715
rect 17000 15555 17040 15685
rect 17000 15525 17005 15555
rect 17035 15525 17040 15555
rect 17000 15395 17040 15525
rect 17000 15365 17005 15395
rect 17035 15365 17040 15395
rect 17000 15235 17040 15365
rect 17000 15205 17005 15235
rect 17035 15205 17040 15235
rect 17000 15200 17040 15205
rect 17080 16195 17120 16200
rect 17080 16165 17085 16195
rect 17115 16165 17120 16195
rect 17080 16035 17120 16165
rect 17080 16005 17085 16035
rect 17115 16005 17120 16035
rect 17080 15875 17120 16005
rect 17080 15845 17085 15875
rect 17115 15845 17120 15875
rect 17080 15715 17120 15845
rect 17080 15685 17085 15715
rect 17115 15685 17120 15715
rect 17080 15555 17120 15685
rect 17080 15525 17085 15555
rect 17115 15525 17120 15555
rect 17080 15395 17120 15525
rect 17080 15365 17085 15395
rect 17115 15365 17120 15395
rect 17080 15235 17120 15365
rect 17080 15205 17085 15235
rect 17115 15205 17120 15235
rect 17080 15200 17120 15205
rect 17160 16195 17200 16200
rect 17160 16165 17165 16195
rect 17195 16165 17200 16195
rect 17160 16035 17200 16165
rect 17160 16005 17165 16035
rect 17195 16005 17200 16035
rect 17160 15875 17200 16005
rect 17160 15845 17165 15875
rect 17195 15845 17200 15875
rect 17160 15715 17200 15845
rect 17160 15685 17165 15715
rect 17195 15685 17200 15715
rect 17160 15555 17200 15685
rect 17160 15525 17165 15555
rect 17195 15525 17200 15555
rect 17160 15395 17200 15525
rect 17160 15365 17165 15395
rect 17195 15365 17200 15395
rect 17160 15235 17200 15365
rect 17160 15205 17165 15235
rect 17195 15205 17200 15235
rect 17160 15200 17200 15205
rect 17240 16195 17280 16200
rect 17240 16165 17245 16195
rect 17275 16165 17280 16195
rect 17240 16035 17280 16165
rect 17240 16005 17245 16035
rect 17275 16005 17280 16035
rect 17240 15875 17280 16005
rect 17240 15845 17245 15875
rect 17275 15845 17280 15875
rect 17240 15715 17280 15845
rect 17240 15685 17245 15715
rect 17275 15685 17280 15715
rect 17240 15555 17280 15685
rect 17240 15525 17245 15555
rect 17275 15525 17280 15555
rect 17240 15395 17280 15525
rect 17240 15365 17245 15395
rect 17275 15365 17280 15395
rect 17240 15235 17280 15365
rect 17240 15205 17245 15235
rect 17275 15205 17280 15235
rect 17240 15200 17280 15205
rect 17320 16195 17360 16200
rect 17320 16165 17325 16195
rect 17355 16165 17360 16195
rect 17320 16035 17360 16165
rect 17320 16005 17325 16035
rect 17355 16005 17360 16035
rect 17320 15875 17360 16005
rect 17320 15845 17325 15875
rect 17355 15845 17360 15875
rect 17320 15715 17360 15845
rect 17320 15685 17325 15715
rect 17355 15685 17360 15715
rect 17320 15555 17360 15685
rect 17320 15525 17325 15555
rect 17355 15525 17360 15555
rect 17320 15395 17360 15525
rect 17320 15365 17325 15395
rect 17355 15365 17360 15395
rect 17320 15235 17360 15365
rect 17320 15205 17325 15235
rect 17355 15205 17360 15235
rect 17320 15200 17360 15205
rect 17400 16195 17440 16200
rect 17400 16165 17405 16195
rect 17435 16165 17440 16195
rect 17400 16035 17440 16165
rect 17400 16005 17405 16035
rect 17435 16005 17440 16035
rect 17400 15875 17440 16005
rect 17400 15845 17405 15875
rect 17435 15845 17440 15875
rect 17400 15715 17440 15845
rect 17400 15685 17405 15715
rect 17435 15685 17440 15715
rect 17400 15555 17440 15685
rect 17400 15525 17405 15555
rect 17435 15525 17440 15555
rect 17400 15395 17440 15525
rect 17400 15365 17405 15395
rect 17435 15365 17440 15395
rect 17400 15235 17440 15365
rect 17400 15205 17405 15235
rect 17435 15205 17440 15235
rect 17400 15200 17440 15205
rect 17480 16195 17520 16200
rect 17480 16165 17485 16195
rect 17515 16165 17520 16195
rect 17480 16035 17520 16165
rect 17480 16005 17485 16035
rect 17515 16005 17520 16035
rect 17480 15875 17520 16005
rect 17480 15845 17485 15875
rect 17515 15845 17520 15875
rect 17480 15715 17520 15845
rect 17480 15685 17485 15715
rect 17515 15685 17520 15715
rect 17480 15555 17520 15685
rect 17480 15525 17485 15555
rect 17515 15525 17520 15555
rect 17480 15395 17520 15525
rect 17480 15365 17485 15395
rect 17515 15365 17520 15395
rect 17480 15235 17520 15365
rect 17480 15205 17485 15235
rect 17515 15205 17520 15235
rect 17480 15200 17520 15205
rect 17560 16195 17600 16200
rect 17560 16165 17565 16195
rect 17595 16165 17600 16195
rect 17560 16035 17600 16165
rect 17560 16005 17565 16035
rect 17595 16005 17600 16035
rect 17560 15875 17600 16005
rect 17560 15845 17565 15875
rect 17595 15845 17600 15875
rect 17560 15715 17600 15845
rect 17560 15685 17565 15715
rect 17595 15685 17600 15715
rect 17560 15555 17600 15685
rect 17560 15525 17565 15555
rect 17595 15525 17600 15555
rect 17560 15395 17600 15525
rect 17560 15365 17565 15395
rect 17595 15365 17600 15395
rect 17560 15235 17600 15365
rect 17560 15205 17565 15235
rect 17595 15205 17600 15235
rect 17560 15200 17600 15205
rect 17640 16195 17680 16200
rect 17640 16165 17645 16195
rect 17675 16165 17680 16195
rect 17640 16035 17680 16165
rect 17640 16005 17645 16035
rect 17675 16005 17680 16035
rect 17640 15875 17680 16005
rect 17640 15845 17645 15875
rect 17675 15845 17680 15875
rect 17640 15715 17680 15845
rect 17640 15685 17645 15715
rect 17675 15685 17680 15715
rect 17640 15555 17680 15685
rect 17640 15525 17645 15555
rect 17675 15525 17680 15555
rect 17640 15395 17680 15525
rect 17640 15365 17645 15395
rect 17675 15365 17680 15395
rect 17640 15235 17680 15365
rect 17640 15205 17645 15235
rect 17675 15205 17680 15235
rect 17640 15200 17680 15205
rect 17720 16195 17760 16200
rect 17720 16165 17725 16195
rect 17755 16165 17760 16195
rect 17720 16035 17760 16165
rect 17720 16005 17725 16035
rect 17755 16005 17760 16035
rect 17720 15875 17760 16005
rect 17720 15845 17725 15875
rect 17755 15845 17760 15875
rect 17720 15715 17760 15845
rect 17720 15685 17725 15715
rect 17755 15685 17760 15715
rect 17720 15555 17760 15685
rect 17720 15525 17725 15555
rect 17755 15525 17760 15555
rect 17720 15395 17760 15525
rect 17720 15365 17725 15395
rect 17755 15365 17760 15395
rect 17720 15235 17760 15365
rect 17720 15205 17725 15235
rect 17755 15205 17760 15235
rect 17720 15200 17760 15205
rect 17800 16195 17840 16200
rect 17800 16165 17805 16195
rect 17835 16165 17840 16195
rect 17800 16035 17840 16165
rect 17800 16005 17805 16035
rect 17835 16005 17840 16035
rect 17800 15875 17840 16005
rect 17800 15845 17805 15875
rect 17835 15845 17840 15875
rect 17800 15715 17840 15845
rect 17800 15685 17805 15715
rect 17835 15685 17840 15715
rect 17800 15555 17840 15685
rect 17800 15525 17805 15555
rect 17835 15525 17840 15555
rect 17800 15395 17840 15525
rect 17800 15365 17805 15395
rect 17835 15365 17840 15395
rect 17800 15235 17840 15365
rect 17800 15205 17805 15235
rect 17835 15205 17840 15235
rect 17800 15200 17840 15205
rect 17880 16195 17920 16200
rect 17880 16165 17885 16195
rect 17915 16165 17920 16195
rect 17880 16035 17920 16165
rect 17880 16005 17885 16035
rect 17915 16005 17920 16035
rect 17880 15875 17920 16005
rect 17880 15845 17885 15875
rect 17915 15845 17920 15875
rect 17880 15715 17920 15845
rect 17880 15685 17885 15715
rect 17915 15685 17920 15715
rect 17880 15555 17920 15685
rect 17880 15525 17885 15555
rect 17915 15525 17920 15555
rect 17880 15395 17920 15525
rect 17880 15365 17885 15395
rect 17915 15365 17920 15395
rect 17880 15235 17920 15365
rect 17880 15205 17885 15235
rect 17915 15205 17920 15235
rect 17880 15200 17920 15205
rect 17960 16195 18000 16200
rect 17960 16165 17965 16195
rect 17995 16165 18000 16195
rect 17960 16035 18000 16165
rect 17960 16005 17965 16035
rect 17995 16005 18000 16035
rect 17960 15875 18000 16005
rect 17960 15845 17965 15875
rect 17995 15845 18000 15875
rect 17960 15715 18000 15845
rect 17960 15685 17965 15715
rect 17995 15685 18000 15715
rect 17960 15555 18000 15685
rect 17960 15525 17965 15555
rect 17995 15525 18000 15555
rect 17960 15395 18000 15525
rect 17960 15365 17965 15395
rect 17995 15365 18000 15395
rect 17960 15235 18000 15365
rect 17960 15205 17965 15235
rect 17995 15205 18000 15235
rect 17960 15200 18000 15205
rect 18040 16195 18080 16200
rect 18040 16165 18045 16195
rect 18075 16165 18080 16195
rect 18040 16035 18080 16165
rect 18040 16005 18045 16035
rect 18075 16005 18080 16035
rect 18040 15875 18080 16005
rect 18040 15845 18045 15875
rect 18075 15845 18080 15875
rect 18040 15715 18080 15845
rect 18040 15685 18045 15715
rect 18075 15685 18080 15715
rect 18040 15555 18080 15685
rect 18040 15525 18045 15555
rect 18075 15525 18080 15555
rect 18040 15395 18080 15525
rect 18040 15365 18045 15395
rect 18075 15365 18080 15395
rect 18040 15235 18080 15365
rect 18040 15205 18045 15235
rect 18075 15205 18080 15235
rect 18040 15200 18080 15205
rect 18120 16195 18160 16200
rect 18120 16165 18125 16195
rect 18155 16165 18160 16195
rect 18120 16035 18160 16165
rect 18120 16005 18125 16035
rect 18155 16005 18160 16035
rect 18120 15875 18160 16005
rect 18120 15845 18125 15875
rect 18155 15845 18160 15875
rect 18120 15715 18160 15845
rect 18120 15685 18125 15715
rect 18155 15685 18160 15715
rect 18120 15555 18160 15685
rect 18120 15525 18125 15555
rect 18155 15525 18160 15555
rect 18120 15395 18160 15525
rect 18120 15365 18125 15395
rect 18155 15365 18160 15395
rect 18120 15235 18160 15365
rect 18120 15205 18125 15235
rect 18155 15205 18160 15235
rect 18120 15200 18160 15205
rect 18200 16195 18240 16200
rect 18200 16165 18205 16195
rect 18235 16165 18240 16195
rect 18200 16035 18240 16165
rect 18200 16005 18205 16035
rect 18235 16005 18240 16035
rect 18200 15875 18240 16005
rect 18200 15845 18205 15875
rect 18235 15845 18240 15875
rect 18200 15715 18240 15845
rect 18200 15685 18205 15715
rect 18235 15685 18240 15715
rect 18200 15555 18240 15685
rect 18200 15525 18205 15555
rect 18235 15525 18240 15555
rect 18200 15395 18240 15525
rect 18200 15365 18205 15395
rect 18235 15365 18240 15395
rect 18200 15235 18240 15365
rect 18200 15205 18205 15235
rect 18235 15205 18240 15235
rect 18200 15200 18240 15205
rect 18280 16195 18320 16200
rect 18280 16165 18285 16195
rect 18315 16165 18320 16195
rect 18280 16035 18320 16165
rect 18280 16005 18285 16035
rect 18315 16005 18320 16035
rect 18280 15875 18320 16005
rect 18280 15845 18285 15875
rect 18315 15845 18320 15875
rect 18280 15715 18320 15845
rect 18280 15685 18285 15715
rect 18315 15685 18320 15715
rect 18280 15555 18320 15685
rect 18280 15525 18285 15555
rect 18315 15525 18320 15555
rect 18280 15395 18320 15525
rect 18280 15365 18285 15395
rect 18315 15365 18320 15395
rect 18280 15235 18320 15365
rect 18280 15205 18285 15235
rect 18315 15205 18320 15235
rect 18280 15200 18320 15205
rect 18360 16195 18400 16200
rect 18360 16165 18365 16195
rect 18395 16165 18400 16195
rect 18360 16035 18400 16165
rect 18360 16005 18365 16035
rect 18395 16005 18400 16035
rect 18360 15875 18400 16005
rect 18360 15845 18365 15875
rect 18395 15845 18400 15875
rect 18360 15715 18400 15845
rect 18360 15685 18365 15715
rect 18395 15685 18400 15715
rect 18360 15555 18400 15685
rect 18360 15525 18365 15555
rect 18395 15525 18400 15555
rect 18360 15395 18400 15525
rect 18360 15365 18365 15395
rect 18395 15365 18400 15395
rect 18360 15235 18400 15365
rect 18360 15205 18365 15235
rect 18395 15205 18400 15235
rect 18360 15200 18400 15205
rect 18440 16195 18480 16200
rect 18440 16165 18445 16195
rect 18475 16165 18480 16195
rect 18440 16035 18480 16165
rect 18440 16005 18445 16035
rect 18475 16005 18480 16035
rect 18440 15875 18480 16005
rect 18440 15845 18445 15875
rect 18475 15845 18480 15875
rect 18440 15715 18480 15845
rect 18440 15685 18445 15715
rect 18475 15685 18480 15715
rect 18440 15555 18480 15685
rect 18440 15525 18445 15555
rect 18475 15525 18480 15555
rect 18440 15395 18480 15525
rect 18440 15365 18445 15395
rect 18475 15365 18480 15395
rect 18440 15235 18480 15365
rect 18440 15205 18445 15235
rect 18475 15205 18480 15235
rect 18440 15200 18480 15205
rect 18520 16195 18560 16200
rect 18520 16165 18525 16195
rect 18555 16165 18560 16195
rect 18520 16035 18560 16165
rect 18520 16005 18525 16035
rect 18555 16005 18560 16035
rect 18520 15875 18560 16005
rect 18520 15845 18525 15875
rect 18555 15845 18560 15875
rect 18520 15715 18560 15845
rect 18520 15685 18525 15715
rect 18555 15685 18560 15715
rect 18520 15555 18560 15685
rect 18520 15525 18525 15555
rect 18555 15525 18560 15555
rect 18520 15395 18560 15525
rect 18520 15365 18525 15395
rect 18555 15365 18560 15395
rect 18520 15235 18560 15365
rect 18520 15205 18525 15235
rect 18555 15205 18560 15235
rect 18520 15200 18560 15205
rect 18600 16195 18640 16200
rect 18600 16165 18605 16195
rect 18635 16165 18640 16195
rect 18600 16035 18640 16165
rect 18600 16005 18605 16035
rect 18635 16005 18640 16035
rect 18600 15875 18640 16005
rect 18600 15845 18605 15875
rect 18635 15845 18640 15875
rect 18600 15715 18640 15845
rect 18600 15685 18605 15715
rect 18635 15685 18640 15715
rect 18600 15555 18640 15685
rect 18600 15525 18605 15555
rect 18635 15525 18640 15555
rect 18600 15395 18640 15525
rect 18600 15365 18605 15395
rect 18635 15365 18640 15395
rect 18600 15235 18640 15365
rect 18600 15205 18605 15235
rect 18635 15205 18640 15235
rect 18600 15200 18640 15205
rect 18680 16195 18720 16200
rect 18680 16165 18685 16195
rect 18715 16165 18720 16195
rect 18680 16035 18720 16165
rect 18680 16005 18685 16035
rect 18715 16005 18720 16035
rect 18680 15875 18720 16005
rect 18680 15845 18685 15875
rect 18715 15845 18720 15875
rect 18680 15715 18720 15845
rect 18680 15685 18685 15715
rect 18715 15685 18720 15715
rect 18680 15555 18720 15685
rect 18680 15525 18685 15555
rect 18715 15525 18720 15555
rect 18680 15395 18720 15525
rect 18680 15365 18685 15395
rect 18715 15365 18720 15395
rect 18680 15235 18720 15365
rect 18680 15205 18685 15235
rect 18715 15205 18720 15235
rect 18680 15200 18720 15205
rect 18760 16195 18800 16200
rect 18760 16165 18765 16195
rect 18795 16165 18800 16195
rect 18760 16035 18800 16165
rect 18760 16005 18765 16035
rect 18795 16005 18800 16035
rect 18760 15875 18800 16005
rect 18760 15845 18765 15875
rect 18795 15845 18800 15875
rect 18760 15715 18800 15845
rect 18760 15685 18765 15715
rect 18795 15685 18800 15715
rect 18760 15555 18800 15685
rect 18760 15525 18765 15555
rect 18795 15525 18800 15555
rect 18760 15395 18800 15525
rect 18760 15365 18765 15395
rect 18795 15365 18800 15395
rect 18760 15235 18800 15365
rect 18760 15205 18765 15235
rect 18795 15205 18800 15235
rect 18760 15200 18800 15205
rect 18840 16195 18880 16200
rect 18840 16165 18845 16195
rect 18875 16165 18880 16195
rect 18840 16035 18880 16165
rect 18840 16005 18845 16035
rect 18875 16005 18880 16035
rect 18840 15875 18880 16005
rect 18840 15845 18845 15875
rect 18875 15845 18880 15875
rect 18840 15715 18880 15845
rect 18840 15685 18845 15715
rect 18875 15685 18880 15715
rect 18840 15555 18880 15685
rect 18840 15525 18845 15555
rect 18875 15525 18880 15555
rect 18840 15395 18880 15525
rect 18840 15365 18845 15395
rect 18875 15365 18880 15395
rect 18840 15235 18880 15365
rect 18840 15205 18845 15235
rect 18875 15205 18880 15235
rect 18840 15200 18880 15205
rect 18920 16195 18960 16200
rect 18920 16165 18925 16195
rect 18955 16165 18960 16195
rect 18920 16035 18960 16165
rect 18920 16005 18925 16035
rect 18955 16005 18960 16035
rect 18920 15875 18960 16005
rect 18920 15845 18925 15875
rect 18955 15845 18960 15875
rect 18920 15715 18960 15845
rect 18920 15685 18925 15715
rect 18955 15685 18960 15715
rect 18920 15555 18960 15685
rect 18920 15525 18925 15555
rect 18955 15525 18960 15555
rect 18920 15395 18960 15525
rect 18920 15365 18925 15395
rect 18955 15365 18960 15395
rect 18920 15235 18960 15365
rect 18920 15205 18925 15235
rect 18955 15205 18960 15235
rect 18920 15200 18960 15205
rect 19000 16195 19040 16200
rect 19000 16165 19005 16195
rect 19035 16165 19040 16195
rect 19000 16035 19040 16165
rect 19000 16005 19005 16035
rect 19035 16005 19040 16035
rect 19000 15875 19040 16005
rect 19000 15845 19005 15875
rect 19035 15845 19040 15875
rect 19000 15715 19040 15845
rect 19000 15685 19005 15715
rect 19035 15685 19040 15715
rect 19000 15555 19040 15685
rect 19000 15525 19005 15555
rect 19035 15525 19040 15555
rect 19000 15395 19040 15525
rect 19000 15365 19005 15395
rect 19035 15365 19040 15395
rect 19000 15235 19040 15365
rect 19000 15205 19005 15235
rect 19035 15205 19040 15235
rect 19000 15200 19040 15205
rect 19080 16195 19120 16200
rect 19080 16165 19085 16195
rect 19115 16165 19120 16195
rect 19080 16035 19120 16165
rect 19080 16005 19085 16035
rect 19115 16005 19120 16035
rect 19080 15875 19120 16005
rect 19080 15845 19085 15875
rect 19115 15845 19120 15875
rect 19080 15715 19120 15845
rect 19080 15685 19085 15715
rect 19115 15685 19120 15715
rect 19080 15555 19120 15685
rect 19080 15525 19085 15555
rect 19115 15525 19120 15555
rect 19080 15395 19120 15525
rect 19080 15365 19085 15395
rect 19115 15365 19120 15395
rect 19080 15235 19120 15365
rect 19080 15205 19085 15235
rect 19115 15205 19120 15235
rect 19080 15200 19120 15205
rect 19160 16195 19200 16200
rect 19160 16165 19165 16195
rect 19195 16165 19200 16195
rect 19160 16035 19200 16165
rect 19160 16005 19165 16035
rect 19195 16005 19200 16035
rect 19160 15875 19200 16005
rect 19160 15845 19165 15875
rect 19195 15845 19200 15875
rect 19160 15715 19200 15845
rect 19160 15685 19165 15715
rect 19195 15685 19200 15715
rect 19160 15555 19200 15685
rect 19160 15525 19165 15555
rect 19195 15525 19200 15555
rect 19160 15395 19200 15525
rect 19160 15365 19165 15395
rect 19195 15365 19200 15395
rect 19160 15235 19200 15365
rect 19160 15205 19165 15235
rect 19195 15205 19200 15235
rect 19160 15200 19200 15205
rect 19240 16195 19280 16200
rect 19240 16165 19245 16195
rect 19275 16165 19280 16195
rect 19240 16035 19280 16165
rect 19240 16005 19245 16035
rect 19275 16005 19280 16035
rect 19240 15875 19280 16005
rect 19240 15845 19245 15875
rect 19275 15845 19280 15875
rect 19240 15715 19280 15845
rect 19240 15685 19245 15715
rect 19275 15685 19280 15715
rect 19240 15555 19280 15685
rect 19240 15525 19245 15555
rect 19275 15525 19280 15555
rect 19240 15395 19280 15525
rect 19240 15365 19245 15395
rect 19275 15365 19280 15395
rect 19240 15235 19280 15365
rect 19240 15205 19245 15235
rect 19275 15205 19280 15235
rect 19240 15200 19280 15205
rect 19320 16195 19360 16200
rect 19320 16165 19325 16195
rect 19355 16165 19360 16195
rect 19320 16035 19360 16165
rect 19320 16005 19325 16035
rect 19355 16005 19360 16035
rect 19320 15875 19360 16005
rect 19320 15845 19325 15875
rect 19355 15845 19360 15875
rect 19320 15715 19360 15845
rect 19320 15685 19325 15715
rect 19355 15685 19360 15715
rect 19320 15555 19360 15685
rect 19320 15525 19325 15555
rect 19355 15525 19360 15555
rect 19320 15395 19360 15525
rect 19320 15365 19325 15395
rect 19355 15365 19360 15395
rect 19320 15235 19360 15365
rect 19320 15205 19325 15235
rect 19355 15205 19360 15235
rect 19320 15200 19360 15205
rect 19400 16195 19440 16200
rect 19400 16165 19405 16195
rect 19435 16165 19440 16195
rect 19400 16035 19440 16165
rect 19400 16005 19405 16035
rect 19435 16005 19440 16035
rect 19400 15875 19440 16005
rect 19400 15845 19405 15875
rect 19435 15845 19440 15875
rect 19400 15715 19440 15845
rect 19400 15685 19405 15715
rect 19435 15685 19440 15715
rect 19400 15555 19440 15685
rect 19400 15525 19405 15555
rect 19435 15525 19440 15555
rect 19400 15395 19440 15525
rect 19400 15365 19405 15395
rect 19435 15365 19440 15395
rect 19400 15235 19440 15365
rect 19400 15205 19405 15235
rect 19435 15205 19440 15235
rect 19400 15200 19440 15205
rect 19480 16195 19520 16200
rect 19480 16165 19485 16195
rect 19515 16165 19520 16195
rect 19480 16035 19520 16165
rect 19480 16005 19485 16035
rect 19515 16005 19520 16035
rect 19480 15875 19520 16005
rect 19480 15845 19485 15875
rect 19515 15845 19520 15875
rect 19480 15715 19520 15845
rect 19480 15685 19485 15715
rect 19515 15685 19520 15715
rect 19480 15555 19520 15685
rect 19480 15525 19485 15555
rect 19515 15525 19520 15555
rect 19480 15395 19520 15525
rect 19480 15365 19485 15395
rect 19515 15365 19520 15395
rect 19480 15235 19520 15365
rect 19480 15205 19485 15235
rect 19515 15205 19520 15235
rect 19480 15200 19520 15205
rect 19560 16195 19600 16200
rect 19560 16165 19565 16195
rect 19595 16165 19600 16195
rect 19560 16035 19600 16165
rect 19560 16005 19565 16035
rect 19595 16005 19600 16035
rect 19560 15875 19600 16005
rect 19560 15845 19565 15875
rect 19595 15845 19600 15875
rect 19560 15715 19600 15845
rect 19560 15685 19565 15715
rect 19595 15685 19600 15715
rect 19560 15555 19600 15685
rect 19560 15525 19565 15555
rect 19595 15525 19600 15555
rect 19560 15395 19600 15525
rect 19560 15365 19565 15395
rect 19595 15365 19600 15395
rect 19560 15235 19600 15365
rect 19560 15205 19565 15235
rect 19595 15205 19600 15235
rect 19560 15200 19600 15205
rect 19640 16195 19680 16200
rect 19640 16165 19645 16195
rect 19675 16165 19680 16195
rect 19640 16035 19680 16165
rect 19640 16005 19645 16035
rect 19675 16005 19680 16035
rect 19640 15875 19680 16005
rect 19640 15845 19645 15875
rect 19675 15845 19680 15875
rect 19640 15715 19680 15845
rect 19640 15685 19645 15715
rect 19675 15685 19680 15715
rect 19640 15555 19680 15685
rect 19640 15525 19645 15555
rect 19675 15525 19680 15555
rect 19640 15395 19680 15525
rect 19640 15365 19645 15395
rect 19675 15365 19680 15395
rect 19640 15235 19680 15365
rect 19640 15205 19645 15235
rect 19675 15205 19680 15235
rect 19640 15200 19680 15205
rect 19720 16195 19760 16200
rect 19720 16165 19725 16195
rect 19755 16165 19760 16195
rect 19720 16035 19760 16165
rect 19720 16005 19725 16035
rect 19755 16005 19760 16035
rect 19720 15875 19760 16005
rect 19720 15845 19725 15875
rect 19755 15845 19760 15875
rect 19720 15715 19760 15845
rect 19720 15685 19725 15715
rect 19755 15685 19760 15715
rect 19720 15555 19760 15685
rect 19720 15525 19725 15555
rect 19755 15525 19760 15555
rect 19720 15395 19760 15525
rect 19720 15365 19725 15395
rect 19755 15365 19760 15395
rect 19720 15235 19760 15365
rect 19720 15205 19725 15235
rect 19755 15205 19760 15235
rect 19720 15200 19760 15205
rect 19800 16195 19840 16200
rect 19800 16165 19805 16195
rect 19835 16165 19840 16195
rect 19800 16035 19840 16165
rect 19800 16005 19805 16035
rect 19835 16005 19840 16035
rect 19800 15875 19840 16005
rect 19800 15845 19805 15875
rect 19835 15845 19840 15875
rect 19800 15715 19840 15845
rect 19800 15685 19805 15715
rect 19835 15685 19840 15715
rect 19800 15555 19840 15685
rect 19800 15525 19805 15555
rect 19835 15525 19840 15555
rect 19800 15395 19840 15525
rect 19800 15365 19805 15395
rect 19835 15365 19840 15395
rect 19800 15235 19840 15365
rect 19800 15205 19805 15235
rect 19835 15205 19840 15235
rect 19800 15200 19840 15205
rect 19880 16195 19920 16200
rect 19880 16165 19885 16195
rect 19915 16165 19920 16195
rect 19880 16035 19920 16165
rect 19880 16005 19885 16035
rect 19915 16005 19920 16035
rect 19880 15875 19920 16005
rect 19880 15845 19885 15875
rect 19915 15845 19920 15875
rect 19880 15715 19920 15845
rect 19880 15685 19885 15715
rect 19915 15685 19920 15715
rect 19880 15555 19920 15685
rect 19880 15525 19885 15555
rect 19915 15525 19920 15555
rect 19880 15395 19920 15525
rect 19880 15365 19885 15395
rect 19915 15365 19920 15395
rect 19880 15235 19920 15365
rect 19880 15205 19885 15235
rect 19915 15205 19920 15235
rect 19880 15200 19920 15205
rect 19960 16195 20000 16200
rect 19960 16165 19965 16195
rect 19995 16165 20000 16195
rect 19960 16035 20000 16165
rect 19960 16005 19965 16035
rect 19995 16005 20000 16035
rect 19960 15875 20000 16005
rect 19960 15845 19965 15875
rect 19995 15845 20000 15875
rect 19960 15715 20000 15845
rect 19960 15685 19965 15715
rect 19995 15685 20000 15715
rect 19960 15555 20000 15685
rect 19960 15525 19965 15555
rect 19995 15525 20000 15555
rect 19960 15395 20000 15525
rect 19960 15365 19965 15395
rect 19995 15365 20000 15395
rect 19960 15235 20000 15365
rect 19960 15205 19965 15235
rect 19995 15205 20000 15235
rect 19960 15200 20000 15205
rect 20040 16195 20080 16200
rect 20040 16165 20045 16195
rect 20075 16165 20080 16195
rect 20040 16035 20080 16165
rect 20040 16005 20045 16035
rect 20075 16005 20080 16035
rect 20040 15875 20080 16005
rect 20040 15845 20045 15875
rect 20075 15845 20080 15875
rect 20040 15715 20080 15845
rect 20040 15685 20045 15715
rect 20075 15685 20080 15715
rect 20040 15555 20080 15685
rect 20040 15525 20045 15555
rect 20075 15525 20080 15555
rect 20040 15395 20080 15525
rect 20040 15365 20045 15395
rect 20075 15365 20080 15395
rect 20040 15235 20080 15365
rect 20040 15205 20045 15235
rect 20075 15205 20080 15235
rect 20040 15200 20080 15205
rect 20120 16195 20160 16200
rect 20120 16165 20125 16195
rect 20155 16165 20160 16195
rect 20120 16035 20160 16165
rect 20120 16005 20125 16035
rect 20155 16005 20160 16035
rect 20120 15875 20160 16005
rect 20120 15845 20125 15875
rect 20155 15845 20160 15875
rect 20120 15715 20160 15845
rect 20120 15685 20125 15715
rect 20155 15685 20160 15715
rect 20120 15555 20160 15685
rect 20120 15525 20125 15555
rect 20155 15525 20160 15555
rect 20120 15395 20160 15525
rect 20120 15365 20125 15395
rect 20155 15365 20160 15395
rect 20120 15235 20160 15365
rect 20120 15205 20125 15235
rect 20155 15205 20160 15235
rect 20120 15200 20160 15205
rect 20200 16195 20240 16200
rect 20200 16165 20205 16195
rect 20235 16165 20240 16195
rect 20200 16035 20240 16165
rect 20200 16005 20205 16035
rect 20235 16005 20240 16035
rect 20200 15875 20240 16005
rect 20200 15845 20205 15875
rect 20235 15845 20240 15875
rect 20200 15715 20240 15845
rect 20200 15685 20205 15715
rect 20235 15685 20240 15715
rect 20200 15555 20240 15685
rect 20200 15525 20205 15555
rect 20235 15525 20240 15555
rect 20200 15395 20240 15525
rect 20200 15365 20205 15395
rect 20235 15365 20240 15395
rect 20200 15235 20240 15365
rect 20200 15205 20205 15235
rect 20235 15205 20240 15235
rect 20200 15200 20240 15205
rect 20280 16195 20320 16200
rect 20280 16165 20285 16195
rect 20315 16165 20320 16195
rect 20280 16035 20320 16165
rect 20280 16005 20285 16035
rect 20315 16005 20320 16035
rect 20280 15875 20320 16005
rect 20280 15845 20285 15875
rect 20315 15845 20320 15875
rect 20280 15715 20320 15845
rect 20280 15685 20285 15715
rect 20315 15685 20320 15715
rect 20280 15555 20320 15685
rect 20280 15525 20285 15555
rect 20315 15525 20320 15555
rect 20280 15395 20320 15525
rect 20280 15365 20285 15395
rect 20315 15365 20320 15395
rect 20280 15235 20320 15365
rect 20280 15205 20285 15235
rect 20315 15205 20320 15235
rect 20280 15200 20320 15205
rect 20360 16195 20400 16200
rect 20360 16165 20365 16195
rect 20395 16165 20400 16195
rect 20360 16035 20400 16165
rect 20360 16005 20365 16035
rect 20395 16005 20400 16035
rect 20360 15875 20400 16005
rect 20360 15845 20365 15875
rect 20395 15845 20400 15875
rect 20360 15715 20400 15845
rect 20360 15685 20365 15715
rect 20395 15685 20400 15715
rect 20360 15555 20400 15685
rect 20360 15525 20365 15555
rect 20395 15525 20400 15555
rect 20360 15395 20400 15525
rect 20360 15365 20365 15395
rect 20395 15365 20400 15395
rect 20360 15235 20400 15365
rect 20360 15205 20365 15235
rect 20395 15205 20400 15235
rect 20360 15200 20400 15205
rect 20440 16195 20480 16200
rect 20440 16165 20445 16195
rect 20475 16165 20480 16195
rect 20440 16035 20480 16165
rect 20440 16005 20445 16035
rect 20475 16005 20480 16035
rect 20440 15875 20480 16005
rect 20440 15845 20445 15875
rect 20475 15845 20480 15875
rect 20440 15715 20480 15845
rect 20440 15685 20445 15715
rect 20475 15685 20480 15715
rect 20440 15555 20480 15685
rect 20440 15525 20445 15555
rect 20475 15525 20480 15555
rect 20440 15395 20480 15525
rect 20440 15365 20445 15395
rect 20475 15365 20480 15395
rect 20440 15235 20480 15365
rect 20440 15205 20445 15235
rect 20475 15205 20480 15235
rect 20440 15200 20480 15205
rect 20520 16195 20560 16200
rect 20520 16165 20525 16195
rect 20555 16165 20560 16195
rect 20520 16035 20560 16165
rect 20520 16005 20525 16035
rect 20555 16005 20560 16035
rect 20520 15875 20560 16005
rect 20520 15845 20525 15875
rect 20555 15845 20560 15875
rect 20520 15715 20560 15845
rect 20520 15685 20525 15715
rect 20555 15685 20560 15715
rect 20520 15555 20560 15685
rect 20520 15525 20525 15555
rect 20555 15525 20560 15555
rect 20520 15395 20560 15525
rect 20520 15365 20525 15395
rect 20555 15365 20560 15395
rect 20520 15235 20560 15365
rect 20520 15205 20525 15235
rect 20555 15205 20560 15235
rect 20520 15200 20560 15205
rect 20600 16195 20640 16200
rect 20600 16165 20605 16195
rect 20635 16165 20640 16195
rect 20600 16035 20640 16165
rect 20600 16005 20605 16035
rect 20635 16005 20640 16035
rect 20600 15875 20640 16005
rect 20600 15845 20605 15875
rect 20635 15845 20640 15875
rect 20600 15715 20640 15845
rect 20600 15685 20605 15715
rect 20635 15685 20640 15715
rect 20600 15555 20640 15685
rect 20600 15525 20605 15555
rect 20635 15525 20640 15555
rect 20600 15395 20640 15525
rect 20600 15365 20605 15395
rect 20635 15365 20640 15395
rect 20600 15235 20640 15365
rect 20600 15205 20605 15235
rect 20635 15205 20640 15235
rect 20600 15200 20640 15205
rect 20680 16195 20720 16200
rect 20680 16165 20685 16195
rect 20715 16165 20720 16195
rect 20680 16035 20720 16165
rect 20680 16005 20685 16035
rect 20715 16005 20720 16035
rect 20680 15875 20720 16005
rect 20680 15845 20685 15875
rect 20715 15845 20720 15875
rect 20680 15715 20720 15845
rect 20680 15685 20685 15715
rect 20715 15685 20720 15715
rect 20680 15555 20720 15685
rect 20680 15525 20685 15555
rect 20715 15525 20720 15555
rect 20680 15395 20720 15525
rect 20680 15365 20685 15395
rect 20715 15365 20720 15395
rect 20680 15235 20720 15365
rect 20680 15205 20685 15235
rect 20715 15205 20720 15235
rect 20680 15200 20720 15205
rect 20760 16195 20800 16200
rect 20760 16165 20765 16195
rect 20795 16165 20800 16195
rect 20760 16035 20800 16165
rect 20760 16005 20765 16035
rect 20795 16005 20800 16035
rect 20760 15875 20800 16005
rect 20760 15845 20765 15875
rect 20795 15845 20800 15875
rect 20760 15715 20800 15845
rect 20760 15685 20765 15715
rect 20795 15685 20800 15715
rect 20760 15555 20800 15685
rect 20760 15525 20765 15555
rect 20795 15525 20800 15555
rect 20760 15395 20800 15525
rect 20760 15365 20765 15395
rect 20795 15365 20800 15395
rect 20760 15235 20800 15365
rect 20760 15205 20765 15235
rect 20795 15205 20800 15235
rect 20760 15200 20800 15205
rect 20840 16195 20880 16200
rect 20840 16165 20845 16195
rect 20875 16165 20880 16195
rect 20840 16035 20880 16165
rect 20840 16005 20845 16035
rect 20875 16005 20880 16035
rect 20840 15875 20880 16005
rect 20840 15845 20845 15875
rect 20875 15845 20880 15875
rect 20840 15715 20880 15845
rect 20840 15685 20845 15715
rect 20875 15685 20880 15715
rect 20840 15555 20880 15685
rect 20840 15525 20845 15555
rect 20875 15525 20880 15555
rect 20840 15395 20880 15525
rect 20840 15365 20845 15395
rect 20875 15365 20880 15395
rect 20840 15235 20880 15365
rect 20840 15205 20845 15235
rect 20875 15205 20880 15235
rect 20840 15200 20880 15205
rect 20920 16195 20960 16200
rect 20920 16165 20925 16195
rect 20955 16165 20960 16195
rect 20920 16035 20960 16165
rect 20920 16005 20925 16035
rect 20955 16005 20960 16035
rect 20920 15875 20960 16005
rect 20920 15845 20925 15875
rect 20955 15845 20960 15875
rect 20920 15715 20960 15845
rect 20920 15685 20925 15715
rect 20955 15685 20960 15715
rect 20920 15555 20960 15685
rect 20920 15525 20925 15555
rect 20955 15525 20960 15555
rect 20920 15395 20960 15525
rect 20920 15365 20925 15395
rect 20955 15365 20960 15395
rect 20920 15235 20960 15365
rect 20920 15205 20925 15235
rect 20955 15205 20960 15235
rect 20920 15200 20960 15205
rect 16760 15155 16800 15160
rect 16760 15125 16765 15155
rect 16795 15125 16800 15155
rect 16760 14995 16800 15125
rect 16760 14965 16765 14995
rect 16795 14965 16800 14995
rect 16760 14960 16800 14965
rect 16840 15155 16880 15160
rect 16840 15125 16845 15155
rect 16875 15125 16880 15155
rect 16840 14995 16880 15125
rect 16840 14965 16845 14995
rect 16875 14965 16880 14995
rect 16840 14960 16880 14965
rect 16920 15155 16960 15160
rect 16920 15125 16925 15155
rect 16955 15125 16960 15155
rect 16920 14995 16960 15125
rect 16920 14965 16925 14995
rect 16955 14965 16960 14995
rect 16920 14960 16960 14965
rect 17000 15155 17040 15160
rect 17000 15125 17005 15155
rect 17035 15125 17040 15155
rect 17000 14995 17040 15125
rect 17000 14965 17005 14995
rect 17035 14965 17040 14995
rect 17000 14960 17040 14965
rect 17080 15155 17120 15160
rect 17080 15125 17085 15155
rect 17115 15125 17120 15155
rect 17080 14995 17120 15125
rect 17080 14965 17085 14995
rect 17115 14965 17120 14995
rect 17080 14960 17120 14965
rect 17160 15155 17200 15160
rect 17160 15125 17165 15155
rect 17195 15125 17200 15155
rect 17160 14995 17200 15125
rect 17160 14965 17165 14995
rect 17195 14965 17200 14995
rect 17160 14960 17200 14965
rect 17240 15155 17280 15160
rect 17240 15125 17245 15155
rect 17275 15125 17280 15155
rect 17240 14995 17280 15125
rect 17240 14965 17245 14995
rect 17275 14965 17280 14995
rect 17240 14960 17280 14965
rect 17320 15155 17360 15160
rect 17320 15125 17325 15155
rect 17355 15125 17360 15155
rect 17320 14995 17360 15125
rect 17320 14965 17325 14995
rect 17355 14965 17360 14995
rect 17320 14960 17360 14965
rect 17400 15155 17440 15160
rect 17400 15125 17405 15155
rect 17435 15125 17440 15155
rect 17400 14995 17440 15125
rect 17400 14965 17405 14995
rect 17435 14965 17440 14995
rect 17400 14960 17440 14965
rect 17480 15155 17520 15160
rect 17480 15125 17485 15155
rect 17515 15125 17520 15155
rect 17480 14995 17520 15125
rect 17480 14965 17485 14995
rect 17515 14965 17520 14995
rect 17480 14960 17520 14965
rect 17560 15155 17600 15160
rect 17560 15125 17565 15155
rect 17595 15125 17600 15155
rect 17560 14995 17600 15125
rect 17560 14965 17565 14995
rect 17595 14965 17600 14995
rect 17560 14960 17600 14965
rect 17640 15155 17680 15160
rect 17640 15125 17645 15155
rect 17675 15125 17680 15155
rect 17640 14995 17680 15125
rect 17640 14965 17645 14995
rect 17675 14965 17680 14995
rect 17640 14960 17680 14965
rect 17720 15155 17760 15160
rect 17720 15125 17725 15155
rect 17755 15125 17760 15155
rect 17720 14995 17760 15125
rect 17720 14965 17725 14995
rect 17755 14965 17760 14995
rect 17720 14960 17760 14965
rect 17800 15155 17840 15160
rect 17800 15125 17805 15155
rect 17835 15125 17840 15155
rect 17800 14995 17840 15125
rect 17800 14965 17805 14995
rect 17835 14965 17840 14995
rect 17800 14960 17840 14965
rect 17880 15155 17920 15160
rect 17880 15125 17885 15155
rect 17915 15125 17920 15155
rect 17880 14995 17920 15125
rect 17880 14965 17885 14995
rect 17915 14965 17920 14995
rect 17880 14960 17920 14965
rect 17960 15155 18000 15160
rect 17960 15125 17965 15155
rect 17995 15125 18000 15155
rect 17960 14995 18000 15125
rect 17960 14965 17965 14995
rect 17995 14965 18000 14995
rect 17960 14960 18000 14965
rect 18040 15155 18080 15160
rect 18040 15125 18045 15155
rect 18075 15125 18080 15155
rect 18040 14995 18080 15125
rect 18040 14965 18045 14995
rect 18075 14965 18080 14995
rect 18040 14960 18080 14965
rect 18120 15155 18160 15160
rect 18120 15125 18125 15155
rect 18155 15125 18160 15155
rect 18120 14995 18160 15125
rect 18120 14965 18125 14995
rect 18155 14965 18160 14995
rect 18120 14960 18160 14965
rect 18200 15155 18240 15160
rect 18200 15125 18205 15155
rect 18235 15125 18240 15155
rect 18200 14995 18240 15125
rect 18200 14965 18205 14995
rect 18235 14965 18240 14995
rect 18200 14960 18240 14965
rect 18280 15155 18320 15160
rect 18280 15125 18285 15155
rect 18315 15125 18320 15155
rect 18280 14995 18320 15125
rect 18280 14965 18285 14995
rect 18315 14965 18320 14995
rect 18280 14960 18320 14965
rect 18360 15155 18400 15160
rect 18360 15125 18365 15155
rect 18395 15125 18400 15155
rect 18360 14995 18400 15125
rect 18360 14965 18365 14995
rect 18395 14965 18400 14995
rect 18360 14960 18400 14965
rect 18440 15155 18480 15160
rect 18440 15125 18445 15155
rect 18475 15125 18480 15155
rect 18440 14995 18480 15125
rect 18440 14965 18445 14995
rect 18475 14965 18480 14995
rect 18440 14960 18480 14965
rect 18520 15155 18560 15160
rect 18520 15125 18525 15155
rect 18555 15125 18560 15155
rect 18520 14995 18560 15125
rect 18520 14965 18525 14995
rect 18555 14965 18560 14995
rect 18520 14960 18560 14965
rect 18600 15155 18640 15160
rect 18600 15125 18605 15155
rect 18635 15125 18640 15155
rect 18600 14995 18640 15125
rect 18600 14965 18605 14995
rect 18635 14965 18640 14995
rect 18600 14960 18640 14965
rect 18680 15155 18720 15160
rect 18680 15125 18685 15155
rect 18715 15125 18720 15155
rect 18680 14995 18720 15125
rect 18680 14965 18685 14995
rect 18715 14965 18720 14995
rect 18680 14960 18720 14965
rect 18760 15155 18800 15160
rect 18760 15125 18765 15155
rect 18795 15125 18800 15155
rect 18760 14995 18800 15125
rect 18760 14965 18765 14995
rect 18795 14965 18800 14995
rect 18760 14960 18800 14965
rect 18840 15155 18880 15160
rect 18840 15125 18845 15155
rect 18875 15125 18880 15155
rect 18840 14995 18880 15125
rect 18840 14965 18845 14995
rect 18875 14965 18880 14995
rect 18840 14960 18880 14965
rect 18920 15155 18960 15160
rect 18920 15125 18925 15155
rect 18955 15125 18960 15155
rect 18920 14995 18960 15125
rect 18920 14965 18925 14995
rect 18955 14965 18960 14995
rect 18920 14960 18960 14965
rect 19000 15155 19040 15160
rect 19000 15125 19005 15155
rect 19035 15125 19040 15155
rect 19000 14995 19040 15125
rect 19000 14965 19005 14995
rect 19035 14965 19040 14995
rect 19000 14960 19040 14965
rect 19080 15155 19120 15160
rect 19080 15125 19085 15155
rect 19115 15125 19120 15155
rect 19080 14995 19120 15125
rect 19080 14965 19085 14995
rect 19115 14965 19120 14995
rect 19080 14960 19120 14965
rect 19160 15155 19200 15160
rect 19160 15125 19165 15155
rect 19195 15125 19200 15155
rect 19160 14995 19200 15125
rect 19160 14965 19165 14995
rect 19195 14965 19200 14995
rect 19160 14960 19200 14965
rect 19240 15155 19280 15160
rect 19240 15125 19245 15155
rect 19275 15125 19280 15155
rect 19240 14995 19280 15125
rect 19240 14965 19245 14995
rect 19275 14965 19280 14995
rect 19240 14960 19280 14965
rect 19320 15155 19360 15160
rect 19320 15125 19325 15155
rect 19355 15125 19360 15155
rect 19320 14995 19360 15125
rect 19320 14965 19325 14995
rect 19355 14965 19360 14995
rect 19320 14960 19360 14965
rect 19400 15155 19440 15160
rect 19400 15125 19405 15155
rect 19435 15125 19440 15155
rect 19400 14995 19440 15125
rect 19400 14965 19405 14995
rect 19435 14965 19440 14995
rect 19400 14960 19440 14965
rect 19480 15155 19520 15160
rect 19480 15125 19485 15155
rect 19515 15125 19520 15155
rect 19480 14995 19520 15125
rect 19480 14965 19485 14995
rect 19515 14965 19520 14995
rect 19480 14960 19520 14965
rect 19560 15155 19600 15160
rect 19560 15125 19565 15155
rect 19595 15125 19600 15155
rect 19560 14995 19600 15125
rect 19560 14965 19565 14995
rect 19595 14965 19600 14995
rect 19560 14960 19600 14965
rect 19640 15155 19680 15160
rect 19640 15125 19645 15155
rect 19675 15125 19680 15155
rect 19640 14995 19680 15125
rect 19640 14965 19645 14995
rect 19675 14965 19680 14995
rect 19640 14960 19680 14965
rect 19720 15155 19760 15160
rect 19720 15125 19725 15155
rect 19755 15125 19760 15155
rect 19720 14995 19760 15125
rect 19720 14965 19725 14995
rect 19755 14965 19760 14995
rect 19720 14960 19760 14965
rect 19800 15155 19840 15160
rect 19800 15125 19805 15155
rect 19835 15125 19840 15155
rect 19800 14995 19840 15125
rect 19800 14965 19805 14995
rect 19835 14965 19840 14995
rect 19800 14960 19840 14965
rect 19880 15155 19920 15160
rect 19880 15125 19885 15155
rect 19915 15125 19920 15155
rect 19880 14995 19920 15125
rect 19880 14965 19885 14995
rect 19915 14965 19920 14995
rect 19880 14960 19920 14965
rect 19960 15155 20000 15160
rect 19960 15125 19965 15155
rect 19995 15125 20000 15155
rect 19960 14995 20000 15125
rect 19960 14965 19965 14995
rect 19995 14965 20000 14995
rect 19960 14960 20000 14965
rect 20040 15155 20080 15160
rect 20040 15125 20045 15155
rect 20075 15125 20080 15155
rect 20040 14995 20080 15125
rect 20040 14965 20045 14995
rect 20075 14965 20080 14995
rect 20040 14960 20080 14965
rect 20120 15155 20160 15160
rect 20120 15125 20125 15155
rect 20155 15125 20160 15155
rect 20120 14995 20160 15125
rect 20120 14965 20125 14995
rect 20155 14965 20160 14995
rect 20120 14960 20160 14965
rect 20200 15155 20240 15160
rect 20200 15125 20205 15155
rect 20235 15125 20240 15155
rect 20200 14995 20240 15125
rect 20200 14965 20205 14995
rect 20235 14965 20240 14995
rect 20200 14960 20240 14965
rect 20280 15155 20320 15160
rect 20280 15125 20285 15155
rect 20315 15125 20320 15155
rect 20280 14995 20320 15125
rect 20280 14965 20285 14995
rect 20315 14965 20320 14995
rect 20280 14960 20320 14965
rect 20360 15155 20400 15160
rect 20360 15125 20365 15155
rect 20395 15125 20400 15155
rect 20360 14995 20400 15125
rect 20360 14965 20365 14995
rect 20395 14965 20400 14995
rect 20360 14960 20400 14965
rect 20440 15155 20480 15160
rect 20440 15125 20445 15155
rect 20475 15125 20480 15155
rect 20440 14995 20480 15125
rect 20440 14965 20445 14995
rect 20475 14965 20480 14995
rect 20440 14960 20480 14965
rect 20520 15155 20560 15160
rect 20520 15125 20525 15155
rect 20555 15125 20560 15155
rect 20520 14995 20560 15125
rect 20520 14965 20525 14995
rect 20555 14965 20560 14995
rect 20520 14960 20560 14965
rect 20600 15155 20640 15160
rect 20600 15125 20605 15155
rect 20635 15125 20640 15155
rect 20600 14995 20640 15125
rect 20600 14965 20605 14995
rect 20635 14965 20640 14995
rect 20600 14960 20640 14965
rect 20680 15155 20720 15160
rect 20680 15125 20685 15155
rect 20715 15125 20720 15155
rect 20680 14995 20720 15125
rect 20680 14965 20685 14995
rect 20715 14965 20720 14995
rect 20680 14960 20720 14965
rect 20760 15155 20800 15160
rect 20760 15125 20765 15155
rect 20795 15125 20800 15155
rect 20760 14995 20800 15125
rect 20760 14965 20765 14995
rect 20795 14965 20800 14995
rect 20760 14960 20800 14965
rect 20840 15155 20880 15160
rect 20840 15125 20845 15155
rect 20875 15125 20880 15155
rect 20840 14995 20880 15125
rect 20840 14965 20845 14995
rect 20875 14965 20880 14995
rect 20840 14960 20880 14965
rect 20920 15155 20960 15160
rect 20920 15125 20925 15155
rect 20955 15125 20960 15155
rect 20920 14995 20960 15125
rect 20920 14965 20925 14995
rect 20955 14965 20960 14995
rect 20920 14960 20960 14965
rect 16760 14915 16800 14920
rect 16760 14885 16765 14915
rect 16795 14885 16800 14915
rect 16760 14755 16800 14885
rect 16760 14725 16765 14755
rect 16795 14725 16800 14755
rect 16760 14720 16800 14725
rect 16840 14915 16880 14920
rect 16840 14885 16845 14915
rect 16875 14885 16880 14915
rect 16840 14755 16880 14885
rect 16840 14725 16845 14755
rect 16875 14725 16880 14755
rect 16840 14720 16880 14725
rect 16920 14915 16960 14920
rect 16920 14885 16925 14915
rect 16955 14885 16960 14915
rect 16920 14755 16960 14885
rect 16920 14725 16925 14755
rect 16955 14725 16960 14755
rect 16920 14720 16960 14725
rect 17000 14915 17040 14920
rect 17000 14885 17005 14915
rect 17035 14885 17040 14915
rect 17000 14755 17040 14885
rect 17000 14725 17005 14755
rect 17035 14725 17040 14755
rect 17000 14720 17040 14725
rect 17080 14915 17120 14920
rect 17080 14885 17085 14915
rect 17115 14885 17120 14915
rect 17080 14755 17120 14885
rect 17080 14725 17085 14755
rect 17115 14725 17120 14755
rect 17080 14720 17120 14725
rect 17160 14915 17200 14920
rect 17160 14885 17165 14915
rect 17195 14885 17200 14915
rect 17160 14755 17200 14885
rect 17160 14725 17165 14755
rect 17195 14725 17200 14755
rect 17160 14720 17200 14725
rect 17240 14915 17280 14920
rect 17240 14885 17245 14915
rect 17275 14885 17280 14915
rect 17240 14755 17280 14885
rect 17240 14725 17245 14755
rect 17275 14725 17280 14755
rect 17240 14720 17280 14725
rect 17320 14915 17360 14920
rect 17320 14885 17325 14915
rect 17355 14885 17360 14915
rect 17320 14755 17360 14885
rect 17320 14725 17325 14755
rect 17355 14725 17360 14755
rect 17320 14720 17360 14725
rect 17400 14915 17440 14920
rect 17400 14885 17405 14915
rect 17435 14885 17440 14915
rect 17400 14755 17440 14885
rect 17400 14725 17405 14755
rect 17435 14725 17440 14755
rect 17400 14720 17440 14725
rect 17480 14915 17520 14920
rect 17480 14885 17485 14915
rect 17515 14885 17520 14915
rect 17480 14755 17520 14885
rect 17480 14725 17485 14755
rect 17515 14725 17520 14755
rect 17480 14720 17520 14725
rect 17560 14915 17600 14920
rect 17560 14885 17565 14915
rect 17595 14885 17600 14915
rect 17560 14755 17600 14885
rect 17560 14725 17565 14755
rect 17595 14725 17600 14755
rect 17560 14720 17600 14725
rect 17640 14915 17680 14920
rect 17640 14885 17645 14915
rect 17675 14885 17680 14915
rect 17640 14755 17680 14885
rect 17640 14725 17645 14755
rect 17675 14725 17680 14755
rect 17640 14720 17680 14725
rect 17720 14915 17760 14920
rect 17720 14885 17725 14915
rect 17755 14885 17760 14915
rect 17720 14755 17760 14885
rect 17720 14725 17725 14755
rect 17755 14725 17760 14755
rect 17720 14720 17760 14725
rect 17800 14915 17840 14920
rect 17800 14885 17805 14915
rect 17835 14885 17840 14915
rect 17800 14755 17840 14885
rect 17800 14725 17805 14755
rect 17835 14725 17840 14755
rect 17800 14720 17840 14725
rect 17880 14915 17920 14920
rect 17880 14885 17885 14915
rect 17915 14885 17920 14915
rect 17880 14755 17920 14885
rect 17880 14725 17885 14755
rect 17915 14725 17920 14755
rect 17880 14720 17920 14725
rect 17960 14915 18000 14920
rect 17960 14885 17965 14915
rect 17995 14885 18000 14915
rect 17960 14755 18000 14885
rect 17960 14725 17965 14755
rect 17995 14725 18000 14755
rect 17960 14720 18000 14725
rect 18040 14915 18080 14920
rect 18040 14885 18045 14915
rect 18075 14885 18080 14915
rect 18040 14755 18080 14885
rect 18040 14725 18045 14755
rect 18075 14725 18080 14755
rect 18040 14720 18080 14725
rect 18120 14915 18160 14920
rect 18120 14885 18125 14915
rect 18155 14885 18160 14915
rect 18120 14755 18160 14885
rect 18120 14725 18125 14755
rect 18155 14725 18160 14755
rect 18120 14720 18160 14725
rect 18200 14915 18240 14920
rect 18200 14885 18205 14915
rect 18235 14885 18240 14915
rect 18200 14755 18240 14885
rect 18200 14725 18205 14755
rect 18235 14725 18240 14755
rect 18200 14720 18240 14725
rect 18280 14915 18320 14920
rect 18280 14885 18285 14915
rect 18315 14885 18320 14915
rect 18280 14755 18320 14885
rect 18280 14725 18285 14755
rect 18315 14725 18320 14755
rect 18280 14720 18320 14725
rect 18360 14915 18400 14920
rect 18360 14885 18365 14915
rect 18395 14885 18400 14915
rect 18360 14755 18400 14885
rect 18360 14725 18365 14755
rect 18395 14725 18400 14755
rect 18360 14720 18400 14725
rect 18440 14915 18480 14920
rect 18440 14885 18445 14915
rect 18475 14885 18480 14915
rect 18440 14755 18480 14885
rect 18440 14725 18445 14755
rect 18475 14725 18480 14755
rect 18440 14720 18480 14725
rect 18520 14915 18560 14920
rect 18520 14885 18525 14915
rect 18555 14885 18560 14915
rect 18520 14755 18560 14885
rect 18520 14725 18525 14755
rect 18555 14725 18560 14755
rect 18520 14720 18560 14725
rect 18600 14915 18640 14920
rect 18600 14885 18605 14915
rect 18635 14885 18640 14915
rect 18600 14755 18640 14885
rect 18600 14725 18605 14755
rect 18635 14725 18640 14755
rect 18600 14720 18640 14725
rect 18680 14915 18720 14920
rect 18680 14885 18685 14915
rect 18715 14885 18720 14915
rect 18680 14755 18720 14885
rect 18680 14725 18685 14755
rect 18715 14725 18720 14755
rect 18680 14720 18720 14725
rect 18760 14915 18800 14920
rect 18760 14885 18765 14915
rect 18795 14885 18800 14915
rect 18760 14755 18800 14885
rect 18760 14725 18765 14755
rect 18795 14725 18800 14755
rect 18760 14720 18800 14725
rect 18840 14915 18880 14920
rect 18840 14885 18845 14915
rect 18875 14885 18880 14915
rect 18840 14755 18880 14885
rect 18840 14725 18845 14755
rect 18875 14725 18880 14755
rect 18840 14720 18880 14725
rect 18920 14915 18960 14920
rect 18920 14885 18925 14915
rect 18955 14885 18960 14915
rect 18920 14755 18960 14885
rect 18920 14725 18925 14755
rect 18955 14725 18960 14755
rect 18920 14720 18960 14725
rect 19000 14915 19040 14920
rect 19000 14885 19005 14915
rect 19035 14885 19040 14915
rect 19000 14755 19040 14885
rect 19000 14725 19005 14755
rect 19035 14725 19040 14755
rect 19000 14720 19040 14725
rect 19080 14915 19120 14920
rect 19080 14885 19085 14915
rect 19115 14885 19120 14915
rect 19080 14755 19120 14885
rect 19080 14725 19085 14755
rect 19115 14725 19120 14755
rect 19080 14720 19120 14725
rect 19160 14915 19200 14920
rect 19160 14885 19165 14915
rect 19195 14885 19200 14915
rect 19160 14755 19200 14885
rect 19160 14725 19165 14755
rect 19195 14725 19200 14755
rect 19160 14720 19200 14725
rect 19240 14915 19280 14920
rect 19240 14885 19245 14915
rect 19275 14885 19280 14915
rect 19240 14755 19280 14885
rect 19240 14725 19245 14755
rect 19275 14725 19280 14755
rect 19240 14720 19280 14725
rect 19320 14915 19360 14920
rect 19320 14885 19325 14915
rect 19355 14885 19360 14915
rect 19320 14755 19360 14885
rect 19320 14725 19325 14755
rect 19355 14725 19360 14755
rect 19320 14720 19360 14725
rect 19400 14915 19440 14920
rect 19400 14885 19405 14915
rect 19435 14885 19440 14915
rect 19400 14755 19440 14885
rect 19400 14725 19405 14755
rect 19435 14725 19440 14755
rect 19400 14720 19440 14725
rect 19480 14915 19520 14920
rect 19480 14885 19485 14915
rect 19515 14885 19520 14915
rect 19480 14755 19520 14885
rect 19480 14725 19485 14755
rect 19515 14725 19520 14755
rect 19480 14720 19520 14725
rect 19560 14915 19600 14920
rect 19560 14885 19565 14915
rect 19595 14885 19600 14915
rect 19560 14755 19600 14885
rect 19560 14725 19565 14755
rect 19595 14725 19600 14755
rect 19560 14720 19600 14725
rect 19640 14915 19680 14920
rect 19640 14885 19645 14915
rect 19675 14885 19680 14915
rect 19640 14755 19680 14885
rect 19640 14725 19645 14755
rect 19675 14725 19680 14755
rect 19640 14720 19680 14725
rect 19720 14915 19760 14920
rect 19720 14885 19725 14915
rect 19755 14885 19760 14915
rect 19720 14755 19760 14885
rect 19720 14725 19725 14755
rect 19755 14725 19760 14755
rect 19720 14720 19760 14725
rect 19800 14915 19840 14920
rect 19800 14885 19805 14915
rect 19835 14885 19840 14915
rect 19800 14755 19840 14885
rect 19800 14725 19805 14755
rect 19835 14725 19840 14755
rect 19800 14720 19840 14725
rect 19880 14915 19920 14920
rect 19880 14885 19885 14915
rect 19915 14885 19920 14915
rect 19880 14755 19920 14885
rect 19880 14725 19885 14755
rect 19915 14725 19920 14755
rect 19880 14720 19920 14725
rect 19960 14915 20000 14920
rect 19960 14885 19965 14915
rect 19995 14885 20000 14915
rect 19960 14755 20000 14885
rect 19960 14725 19965 14755
rect 19995 14725 20000 14755
rect 19960 14720 20000 14725
rect 20040 14915 20080 14920
rect 20040 14885 20045 14915
rect 20075 14885 20080 14915
rect 20040 14755 20080 14885
rect 20040 14725 20045 14755
rect 20075 14725 20080 14755
rect 20040 14720 20080 14725
rect 20120 14915 20160 14920
rect 20120 14885 20125 14915
rect 20155 14885 20160 14915
rect 20120 14755 20160 14885
rect 20120 14725 20125 14755
rect 20155 14725 20160 14755
rect 20120 14720 20160 14725
rect 20200 14915 20240 14920
rect 20200 14885 20205 14915
rect 20235 14885 20240 14915
rect 20200 14755 20240 14885
rect 20200 14725 20205 14755
rect 20235 14725 20240 14755
rect 20200 14720 20240 14725
rect 20280 14915 20320 14920
rect 20280 14885 20285 14915
rect 20315 14885 20320 14915
rect 20280 14755 20320 14885
rect 20280 14725 20285 14755
rect 20315 14725 20320 14755
rect 20280 14720 20320 14725
rect 20360 14915 20400 14920
rect 20360 14885 20365 14915
rect 20395 14885 20400 14915
rect 20360 14755 20400 14885
rect 20360 14725 20365 14755
rect 20395 14725 20400 14755
rect 20360 14720 20400 14725
rect 20440 14915 20480 14920
rect 20440 14885 20445 14915
rect 20475 14885 20480 14915
rect 20440 14755 20480 14885
rect 20440 14725 20445 14755
rect 20475 14725 20480 14755
rect 20440 14720 20480 14725
rect 20520 14915 20560 14920
rect 20520 14885 20525 14915
rect 20555 14885 20560 14915
rect 20520 14755 20560 14885
rect 20520 14725 20525 14755
rect 20555 14725 20560 14755
rect 20520 14720 20560 14725
rect 20600 14915 20640 14920
rect 20600 14885 20605 14915
rect 20635 14885 20640 14915
rect 20600 14755 20640 14885
rect 20600 14725 20605 14755
rect 20635 14725 20640 14755
rect 20600 14720 20640 14725
rect 20680 14915 20720 14920
rect 20680 14885 20685 14915
rect 20715 14885 20720 14915
rect 20680 14755 20720 14885
rect 20680 14725 20685 14755
rect 20715 14725 20720 14755
rect 20680 14720 20720 14725
rect 20760 14915 20800 14920
rect 20760 14885 20765 14915
rect 20795 14885 20800 14915
rect 20760 14755 20800 14885
rect 20760 14725 20765 14755
rect 20795 14725 20800 14755
rect 20760 14720 20800 14725
rect 20840 14915 20880 14920
rect 20840 14885 20845 14915
rect 20875 14885 20880 14915
rect 20840 14755 20880 14885
rect 20840 14725 20845 14755
rect 20875 14725 20880 14755
rect 20840 14720 20880 14725
rect 20920 14915 20960 14920
rect 20920 14885 20925 14915
rect 20955 14885 20960 14915
rect 20920 14755 20960 14885
rect 20920 14725 20925 14755
rect 20955 14725 20960 14755
rect 20920 14720 20960 14725
<< metal4 >>
rect 0 35240 40 35440
rect 10440 35240 10520 35440
rect 0 35000 40 35200
rect 10440 35000 10520 35200
rect 0 34760 40 34960
rect 10440 34760 10520 34960
rect 0 34520 40 34720
rect 10440 34520 10520 34720
rect 10440 -1320 10520 -1120
rect 10440 -1560 10520 -1360
rect 10440 -1800 10520 -1600
rect 10440 -2040 10520 -1840
<< metal5 >>
rect 80 14720 280 18680
rect 560 14720 760 18680
rect 1040 14720 1240 18680
rect 1520 14720 1720 18680
rect 2000 14720 2200 18680
rect 2480 14720 2680 18680
rect 2960 14720 3160 18680
rect 3440 14720 3640 18680
rect 3920 14720 4120 18680
rect 6320 14720 6520 18680
rect 6800 14720 7000 18680
rect 7280 14720 7480 18680
rect 7760 14720 7960 18680
rect 8240 14720 8440 18680
rect 8720 14720 8920 18680
rect 9200 14720 9400 18680
rect 9680 14720 9880 18680
rect 10160 14720 10360 18680
rect 10600 14720 10800 18680
rect 11080 14720 11280 18680
rect 11560 14720 11760 18680
rect 12040 14720 12240 18680
rect 12520 14720 12720 18680
rect 13000 14720 13200 18680
rect 13480 14720 13680 18680
rect 13960 14720 14160 18680
rect 14440 14720 14640 18680
rect 16840 14720 17040 18680
rect 17320 14720 17520 18680
rect 17800 14720 18000 18680
rect 18280 14720 18480 18680
rect 18760 14720 18960 18680
rect 19240 14720 19440 18680
rect 19720 14720 19920 18680
rect 20200 14720 20400 18680
rect 20680 14720 20880 18680
use ota_core  4
timestamp 1638019703
transform 1 0 10520 0 1 -1080
box 0 -2320 10440 15800
use ota_core  3
timestamp 1638019703
transform -1 0 10440 0 1 -1080
box 0 -2320 10440 15800
use ota_core  2
timestamp 1638019703
transform -1 0 20960 0 -1 34480
box 0 -2320 10440 15800
use ota_core  1
timestamp 1638019703
transform 1 0 0 0 -1 34480
box 0 -2320 10440 15800
<< labels >>
rlabel metal2 0 16080 40 16120 0 im
port 0 nsew
rlabel metal2 0 18080 40 18120 0 ip
port 1 nsew
rlabel metal2 0 15920 40 15960 0 op
port 2 nsew
rlabel metal2 0 17920 40 17960 0 om
port 3 nsew
rlabel metal2 0 18560 40 18600 0 ib
port 4 nsew
rlabel metal2 0 16800 40 16840 0 q
port 5 nsew
rlabel metal2 0 18320 40 18360 0 bp
rlabel metal2 0 17760 40 17800 0 x
rlabel metal2 0 17600 40 17640 0 y
rlabel metal4 0 34520 40 34720 0 vdda
port 6 nsew
rlabel metal4 0 35000 40 35200 0 gnda
port 7 nsew
rlabel metal4 0 35240 40 35440 0 vssa
port 8 nsew
rlabel metal4 0 34760 40 34960 0 vddx
rlabel metal3 5840 18680 5880 18720 0 z
<< end >>
