* iref testbench

* Include SkyWater sky130 device models
.lib "/usr/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.param mc_mm_switch=0
.include "iref.spice"


.param pVDD = 1.8

VDD vdd 0 dc {pVDD} pulse(10m {pVDD} 1m 1m 10u 1 1)
VSS vss 0 0

* DUT
X0 vdd vss dp iref
VDP dp vss 0

.save I(VDP) I(VDD)
.save VDD X0.X X0.Y X0.Z X0.N X0.P0 X0.P1 X0.P2 X0.HI

.option gmin=1e-12
.option scale=1e-6
.control

	op
	print X0.X X0.Y X0.Z X0.N
	print i(vdp) i(vdd)

    dc VDD 0.3 1.8 10m
    let vdd_io = i(vdp)
    let vdd_idd = i(vdd)
    wrdata iref_vdd_io.txt vdd_io
    let vdd_psrr = 20*log10(abs(deriv(I(VDP))/I(VDP)))
    wrdata iref_psrr.txt
    plot vdd_io
    plot vdd_idd
    plot vdd_psrr

	dc temp -55 125 1
	let temp_io = i(vdp)
	wrdata iref_temp_io.txt temp_io
    
	tran 10u 10m
	let tran_io  = i(vdp)
	let tran_vdd = vdd
	wrdata iref_tran_io.txt tran_io 
	wrdata iref_tran_vdd.txt tran_vdd
	plot tran_io
    
.endc

.end
