* NGSPICE file created from iref.ext - technology: sky130A

.subckt iref VDDA VSSA DP
X0 P1 LO N VSSA sky130_fd_pr__nfet_01v8 ad=1.6e+12p pd=1.12e+07u as=1.6e+12p ps=1.12e+07u w=1e+06u l=500000u
X1 a_11370_3380# Y a_11190_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X2 VSSA N a_15320_100# VSSA sky130_fd_pr__nfet_01v8 ad=1.05e+13p pd=7.3e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X3 a_16770_100# N a_16590_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X4 a_17130_1980# P2 a_16950_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X5 a_3980_1980# P2 a_3800_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X6 a_14960_100# N a_14780_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X7 a_4520_3380# N a_4340_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X8 a_2360_3380# Z a_2180_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X9 VDDA P0 a_15320_1500# VDDA sky130_fd_pr__pfet_01v8 ad=9.7e+12p pd=6.74e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X10 a_18930_1980# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=1.6e+12p ps=1.12e+07u w=1e+06u l=500000u
X11 VSSA a_n620_3280# a_200_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X12 a_20370_1980# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X13 a_12800_100# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X14 a_13340_1500# P0 a_13160_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X15 a_200_1500# a_n620_1400# a_20_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X16 a_16770_1980# P2 Y VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X17 P0 P2 a_11000_1500# VDDA sky130_fd_pr__pfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X18 Z Y a_17130_3380# VSSA sky130_fd_pr__nfet_01v8 ad=3.2e+12p pd=2.24e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X19 VSSA N a_14970_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X20 Z X a_4160_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X21 a_20_100# a_n620_70# a_n620_70# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X22 a_12980_1500# P0 a_12800_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X23 a_1820_1500# P2 a_1640_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X24 a_16950_3380# Y a_16770_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X25 a_20550_3380# X a_20370_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X26 a_14790_3380# N a_14610_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X27 VSSA N a_5960_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X28 a_1640_100# X Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X29 a_7230_1980# P2 a_7050_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X30 a_18390_1980# P1 a_18210_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X31 a_19650_100# Z a_19470_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X32 P0 Y a_11000_100# VSSA sky130_fd_pr__nfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X33 a_20550_100# Z a_20370_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X34 a_5780_3380# N a_5600_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X35 a_n520_100# a_n620_70# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X36 a_5600_1500# P2 a_5420_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X37 VDDA P0 a_8850_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X38 a_20_1500# a_n620_1400# a_n620_1400# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X39 a_6870_1980# P0 a_6690_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X40 a_3440_1500# P1 a_3260_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X41 a_1280_1500# P2 a_1100_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X42 VSSA N a_9200_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X43 a_16950_100# N a_16770_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X44 a_7410_3380# N a_7230_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X45 a_18570_3380# X a_18390_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X46 a_22170_3380# a_21350_3280# a_21990_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X47 a_11010_1980# P2 a_10830_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X48 a_16230_1500# P2 a_16050_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X49 a_7220_100# N a_7040_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X50 a_3080_1500# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X51 a_7050_3380# N a_6870_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X52 a_6680_100# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X53 a_21630_1500# a_21350_1400# a_21450_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X54 a_18030_1500# P2 a_17850_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X55 a_2000_1980# P2 DP VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X56 a_15870_1500# P2 a_15690_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X57 a_7220_1500# P1 a_7040_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X58 a_8490_1980# P0 a_8310_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X59 a_4520_100# Y Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X60 a_3980_100# X a_3800_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X61 a_12630_1980# P1 a_12450_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X62 a_9020_1500# P2 a_8840_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X63 a_6860_1500# P1 a_6680_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X64 P0 P2 a_10290_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X65 a_1820_100# X a_1640_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X66 a_11000_1500# P2 a_10820_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X67 a_8670_3380# N a_8490_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X68 a_19650_1500# P2 a_19470_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X69 a_3620_1980# P2 a_3440_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X70 VSSA Z a_19650_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X71 a_11360_100# Y P0 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X72 a_20730_100# Z a_20550_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X73 a_17490_1500# P2 a_17310_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X74 a_1460_1980# P2 a_1280_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X75 a_12810_3380# N a_12630_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X76 a_10650_3380# Y P0 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X77 a_16410_1980# P2 a_16230_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X78 a_14250_1980# P2 a_14070_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X79 a_9560_100# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X80 a_8480_1500# P2 N VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=1.6e+12p ps=1.12e+07u w=1e+06u l=500000u
X81 a_3800_3380# N a_3620_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X82 a_1640_3380# Z a_1460_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X83 a_21350_1950# a_21350_1950# a_21630_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X84 a_7400_100# N a_7220_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X85 VDDA P0 a_12440_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X86 a_16050_1980# P2 a_15870_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X87 a_10460_1500# P0 a_10280_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X88 a_13890_1980# P2 N VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X89 a_5240_1980# P2 a_5060_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X90 a_6860_100# N a_6680_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X91 a_14430_3380# N a_14250_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X92 VSSA N a_12090_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X93 a_n620_1400# a_n620_1400# a_n340_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X94 a_4700_100# Y a_4520_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X95 a_4880_1980# P2 P2 VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X96 a_14070_3380# N a_13890_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X97 P2 N a_5240_3380# VSSA sky130_fd_pr__nfet_01v8 ad=1.6e+12p pd=1.12e+07u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X98 a_14240_100# N P1 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X99 VSSA Z a_3080_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X100 a_19830_1980# P1 a_19650_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X101 VDDA LO a_21090_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X102 a_6510_1980# P0 a_6330_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X103 a_2000_100# X a_1820_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X104 a_14240_1500# P2 P1 VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=8e+11p ps=5.6e+06u w=1e+06u l=500000u
X105 a_17670_1980# P1 a_17490_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X106 a_18210_3380# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X107 a_5060_3380# N a_4880_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X108 a_20010_100# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X109 a_11540_100# Y a_11360_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X110 a_20910_100# Z a_20730_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X111 a_13880_1500# P2 a_13700_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X112 a_2720_1500# P2 a_2540_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X113 VDDA LO a_560_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X114 a_20010_3380# X a_19830_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X115 a_17850_3380# X a_17670_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X116 a_21450_3380# a_21350_3280# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X117 a_15690_3380# X a_15510_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X118 VSSA N a_9560_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X119 a_8130_1980# P2 a_7950_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X120 a_19290_1980# P1 a_19110_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X121 LO N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=8e+11p pd=5.6e+06u as=0p ps=0u w=1e+06u l=500000u
X122 a_20910_1500# P1 a_20730_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X123 a_n340_1980# a_n620_1950# a_n520_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X124 a_7040_100# N a_6860_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X125 VDDA P1 a_6320_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X126 a_10110_1980# P2 a_9930_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X127 a_9930_1980# P2 a_9750_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X128 VSSA N a_18210_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X129 a_4340_1500# P1 a_4160_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X130 a_7770_1980# P2 P1 VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X131 VDDA P1 a_2000_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X132 a_8310_3380# N a_8130_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X133 X X a_19290_3380# VSSA sky130_fd_pr__nfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X134 VDDA P0 a_11730_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X135 P2 N a_16050_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X136 a_17130_1500# P2 P2 VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X137 a_1100_1980# P1 a_920_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X138 a_n520_3380# a_n620_3280# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X139 a_3980_1500# P1 a_3800_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X140 a_14420_100# N a_14240_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X141 a_15690_100# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X142 a_7950_3380# N a_7770_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X143 a_13880_100# N a_13700_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X144 a_18930_1500# P1 a_18750_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X145 a_2900_1980# P1 a_2720_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X146 a_920_1980# P1 a_740_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X147 a_20370_1500# P2 a_20190_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X148 a_16770_1500# P2 a_16590_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X149 a_8120_1500# N N VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X150 a_9390_1980# P0 a_9210_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X151 a_11720_100# Y a_11540_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X152 a_10100_1500# P0 a_9920_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X153 a_13530_1980# N N VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X154 a_9920_1500# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X155 a_3260_100# X a_3080_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X156 a_7760_1500# P2 a_7580_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X157 a_11370_1980# P0 a_11190_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X158 a_9920_100# Y VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X159 a_1100_100# X a_920_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X160 a_11900_1500# P2 a_11720_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X161 a_9570_3380# Y a_9390_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X162 a_22170_100# a_21350_70# a_21990_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X163 a_4520_1980# P2 a_4340_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X164 VDDA P2 a_18210_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X165 a_2360_1980# P2 a_2180_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X166 a_19110_100# Z a_18930_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X167 VDDA a_n620_1950# a_200_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X168 N LO P1 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X169 a_11550_3380# Y a_11370_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X170 a_18570_100# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X171 a_17310_1980# P2 a_17130_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X172 VDDA P1 a_14970_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X173 a_9380_1500# P1 a_9200_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X174 a_4700_3380# N a_4520_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X175 a_16410_100# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X176 a_2540_3380# Z a_2360_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X177 a_560_3380# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X178 a_14600_100# N a_14420_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X179 a_13520_1500# P2 a_13340_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X180 a_20550_1980# P2 a_20370_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X181 a_16950_1980# P2 a_16770_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X182 a_15870_100# N a_15690_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X183 a_11360_1500# P2 P0 VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X184 a_14790_1980# P1 a_14610_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X185 VDDA P2 a_5960_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X186 P1 N a_13880_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X187 a_15330_3380# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X188 a_6140_100# X a_5960_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X189 a_13170_3380# N a_12990_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X190 a_2000_1500# P1 a_1820_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X191 a_11900_100# Y a_11720_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X192 a_5780_1980# P2 a_5600_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X193 a_20730_3380# X a_20550_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X194 a_14970_3380# N a_14790_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X195 a_3440_100# X a_3260_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X196 a_4160_3380# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X197 a_22170_1980# a_21350_1950# a_21990_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X198 a_7410_1980# P2 a_7230_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X199 a_15140_1500# P0 a_14960_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X200 a_18570_1980# P2 a_18390_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X201 VSSA a_21350_70# a_22170_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X202 a_19110_3380# X a_18930_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X203 a_5960_3380# N a_5780_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X204 a_14780_1500# P2 a_14600_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X205 VDDA P1 a_3440_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X206 a_7050_1980# P2 a_6870_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X207 X P2 a_1280_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X208 Z X a_18570_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X209 VSSA a_21350_3280# a_22170_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X210 a_18750_100# Z a_18570_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X211 a_10280_100# Y a_10100_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X212 Y Y a_16410_3380# VSSA sky130_fd_pr__nfet_01v8 ad=8e+11p pd=5.6e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X213 Z X a_20010_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X214 a_16410_1500# P2 a_16230_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X215 a_21990_3380# a_21350_3280# a_21350_3280# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X216 a_8480_100# N N VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X217 a_16050_100# N a_15870_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X218 a_21350_1400# a_21350_1400# a_21630_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X219 a_16050_1500# P2 a_15870_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X220 a_7400_1500# P2 a_7220_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X221 a_6320_100# X a_6140_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X222 a_5240_1500# P2 Y VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X223 a_8670_1980# P0 a_8490_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X224 a_9210_3380# Y VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X225 Z Y a_5600_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X226 a_12810_1980# P2 a_12630_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X227 a_7040_1500# P1 a_6860_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X228 a_10650_1980# P2 P0 VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X229 a_4880_1500# P2 a_4700_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X230 VSSA X a_3440_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X231 a_8850_3380# N a_8670_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X232 a_3800_1980# P2 a_3620_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X233 a_6690_3380# N a_6510_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X234 a_3080_100# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X235 VSSA a_n620_70# a_200_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X236 DP P2 a_19650_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X237 VDDA P1 a_21090_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X238 a_17670_1500# P2 a_17490_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X239 a_1640_1980# P2 a_1460_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X240 a_13160_100# N a_12980_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X241 a_10830_3380# Y a_10650_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X242 a_200_3380# a_n620_3280# a_20_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X243 a_21990_100# a_21350_70# a_21350_70# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X244 a_14430_1980# P2 a_14250_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X245 a_18930_100# Z a_18750_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X246 a_8660_1500# P2 a_8480_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X247 a_12270_1980# P1 a_12090_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X248 a_10460_100# Y a_10280_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X249 VSSA Z a_1640_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X250 a_9200_100# N a_9020_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X251 a_12800_1500# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X252 a_10640_1500# P2 a_10460_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X253 a_14070_1980# P2 a_13890_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X254 a_5420_1980# P2 a_5240_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X255 a_8660_100# N a_8480_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X256 a_19290_1500# P2 a_19110_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X257 VDDA P1 a_3080_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X258 a_14610_3380# N a_14430_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X259 a_12450_3380# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X260 a_n340_1500# a_n620_1400# a_n520_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X261 a_10290_3380# Y a_10110_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X262 VSSA X a_6320_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X263 a_18210_1980# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X264 a_5060_1980# P2 a_4880_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X265 a_5960_100# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X266 a_5600_3380# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X267 a_20_3380# a_n620_3280# a_n620_3280# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X268 a_12090_3380# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X269 a_20010_1980# P2 a_19830_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X270 a_3440_3380# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X271 a_1280_3380# Z a_1100_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X272 a_14420_1500# P2 a_14240_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X273 a_21450_1980# a_21350_1950# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X274 a_17850_1980# P1 a_17670_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X275 a_3800_100# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X276 a_1100_1500# P1 a_920_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X277 a_12260_1500# P0 a_12080_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X278 a_15690_1980# P1 a_15510_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X279 LO N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X280 a_16230_3380# Y a_16050_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X281 a_3080_3380# Z a_2900_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X282 a_13340_100# N a_13160_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X283 P1 P2 a_13880_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X284 X P2 a_2720_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X285 a_21090_1980# LO VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X286 a_920_1500# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X287 VSSA X a_17850_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X288 a_21630_3380# a_21350_3280# a_21450_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X289 Z X a_15690_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X290 a_10640_100# Y a_10460_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X291 a_8310_1980# P2 a_8130_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X292 VDDA P1 a_19290_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X293 X X a_2000_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X294 a_n520_1980# a_n620_1950# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X295 a_8840_100# N a_8660_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X296 a_4520_1500# P2 a_4340_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X297 a_7950_1980# P2 a_7770_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X298 a_2360_1500# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X299 VDDA a_n620_1400# a_200_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X300 a_19650_3380# X X VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X301 a_6330_3380# N VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X302 a_17490_3380# X Z VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X303 a_17310_1500# P2 a_17130_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X304 a_17490_100# N a_17310_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X305 a_20550_1500# P2 a_20370_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X306 P2 P2 a_16770_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X307 N N a_8120_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X308 VSSA N LO VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X309 a_6140_1500# P1 a_5960_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X310 a_9570_1980# P0 a_9390_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X311 a_13520_100# N a_13340_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X312 N N a_13530_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X313 a_12980_100# N a_12800_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X314 N P2 a_7760_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X315 a_11550_1980# P0 a_11370_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X316 a_5780_1500# P2 a_5600_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X317 a_n620_3280# a_n620_3280# a_n340_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X318 a_10820_100# Y a_10640_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X319 a_9750_3380# Y a_9570_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X320 P1 N a_7410_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X321 P2 P2 a_4520_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X322 a_22170_1500# a_21350_1400# a_21990_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X323 a_18570_1500# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X324 a_2540_1980# P2 a_2360_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X325 a_2360_100# X X VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X326 a_560_1980# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X327 a_9020_100# N a_8840_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X328 a_11730_3380# Y a_11550_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X329 VSSA Z a_21090_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X330 a_15330_1980# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X331 a_9560_1500# P1 a_9380_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X332 a_13170_1980# P2 a_12990_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X333 a_18210_100# N a_18030_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X334 a_740_3380# Z a_560_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X335 a_2720_3380# Z a_2540_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X336 a_13700_1500# P2 a_13520_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X337 a_20730_1980# P1 a_20550_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X338 P2 N a_17490_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X339 a_11540_1500# P2 a_11360_1500# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X340 a_14970_1980# P1 a_14790_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X341 a_4160_1980# P2 a_3980_1980# VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X342 a_15510_3380# X a_15330_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X343 N N a_13170_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X344 a_920_100# X VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X345 a_11190_3380# Y a_11010_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X346 a_13700_100# N a_13520_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X347 a_19110_1980# P2 a_18930_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X348 a_5960_1980# P2 a_5780_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X349 VSSA X a_20730_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X350 a_12990_3380# N a_12810_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X351 a_5240_100# Y Y VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X352 a_4340_3380# N a_4160_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X353 a_2180_3380# Z a_2000_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X354 a_15320_1500# P0 a_15140_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X355 VDDA a_21350_1950# a_22170_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X356 X P2 a_18570_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X357 a_11000_100# Y a_10820_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X358 X P2 a_20010_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X359 a_13160_1500# P0 a_12980_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X360 Y P2 a_16410_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X361 a_17130_3380# Y a_16950_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X362 P2 N a_3800_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X363 a_2540_100# X a_2360_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X364 a_14960_1500# P0 a_14780_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X365 a_3800_1500# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X366 a_21990_1980# a_21350_1950# a_21350_1950# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X367 a_1640_1500# P2 X VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X368 a_18930_3380# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X369 a_21450_100# a_21350_70# VSSA VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X370 a_16770_3380# Y Y VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X371 a_20370_3380# X Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X372 a_9210_1980# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X373 a_17850_100# N P2 VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X374 P1 LO N VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X375 a_5420_1500# P2 a_5240_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X376 a_8850_1980# P0 a_8670_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X377 a_3260_1500# P2 a_3080_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X378 a_6690_1980# P0 a_6510_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X379 a_7230_3380# N a_7050_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X380 a_7580_100# N a_7400_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X381 a_18390_3380# X a_18210_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X382 a_10830_1980# P2 a_10650_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X383 a_18210_1500# P2 a_18030_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X384 Y P2 a_4880_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X385 a_200_1980# a_n620_1950# a_20_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X386 a_5420_100# Y a_5240_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X387 VSSA N a_8850_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X388 a_6870_3380# N a_6690_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X389 a_4880_100# Y a_4700_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X390 a_20010_1500# P2 DP VDDA sky130_fd_pr__pfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X391 a_21450_1500# a_21350_1400# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X392 a_17850_1500# P2 a_17670_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X393 DP P2 a_1640_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X394 a_9200_1500# P1 a_9020_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X395 a_15690_1500# P2 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X396 a_11010_3380# Y a_10830_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X397 a_2720_100# X a_2540_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X398 a_14610_1980# P1 a_14430_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X399 a_21090_1500# P1 a_20910_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X400 a_8840_1500# P2 a_8660_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X401 a_12450_1980# P1 a_12270_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X402 a_12260_100# Y a_12080_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X403 a_21630_100# a_21350_70# a_21450_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X404 a_6680_1500# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X405 a_10290_1980# P2 a_10110_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X406 a_2000_3380# Z VSSA VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X407 a_10100_100# Y a_9920_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X408 a_21090_100# Z a_20910_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X409 a_10820_1500# P2 a_10640_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X410 a_8490_3380# N a_8310_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X411 a_12090_1980# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X412 a_5600_1980# P2 a_5420_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X413 a_20_1980# a_n620_1950# a_n620_1950# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X414 a_19470_1500# P2 a_19290_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X415 a_3440_1980# P2 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X416 a_18030_100# N a_17850_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X417 a_1280_1980# P2 a_1100_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X418 a_12630_3380# N a_12450_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X419 a_n520_1500# a_n620_1400# VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X420 P0 Y a_10290_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X421 N LO P1 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X422 a_16230_1980# P2 a_16050_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X423 a_3080_1980# P1 a_2900_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X424 a_7760_100# N a_7580_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X425 a_3620_3380# N a_3440_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X426 a_1460_3380# Z a_1280_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X427 a_14600_1500# P2 a_14420_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X428 a_21630_1980# a_21350_1950# a_21450_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X429 VDDA P1 a_17850_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X430 a_5600_100# Y a_5420_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X431 a_12440_1500# P0 a_12260_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X432 a_15870_1980# P1 a_15690_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X433 a_10280_1500# P0 a_10100_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X434 Y Y a_4880_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X435 a_16410_3380# Y a_16230_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X436 a_15140_100# N a_14960_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X437 a_14250_3380# N a_14070_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X438 Z X a_2720_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X439 a_200_100# a_n620_70# a_20_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X440 a_12080_1500# P0 a_11900_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X441 a_21350_3280# a_21350_3280# a_21630_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X442 a_16050_3380# Y Z VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X443 a_13890_3380# N N VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X444 a_21350_70# a_21350_70# a_21630_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X445 a_5240_3380# N a_5060_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X446 a_12440_100# Y a_12260_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X447 a_19650_1980# P1 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X448 a_6330_1980# P0 VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X449 a_17490_1980# P1 a_17310_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X450 a_4880_3380# N a_4700_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X451 a_4700_1500# P2 a_4520_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X452 a_2540_1500# P1 a_2360_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X453 a_560_1500# LO VDDA VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X454 a_19830_3380# X a_19650_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X455 a_6510_3380# N a_6330_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X456 a_17670_3380# X a_17490_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X457 VSSA N LO VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X458 a_1280_100# X a_1100_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X459 N N a_7760_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X460 a_19290_100# Z a_19110_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X461 a_20190_100# Z a_20010_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X462 a_n620_70# a_n620_70# a_n340_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X463 a_20730_1500# P1 a_20550_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X464 a_n620_1950# a_n620_1950# a_n340_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X465 a_17130_100# N a_16950_100# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X466 a_6320_1500# P1 a_6140_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X467 a_9750_1980# P0 a_9570_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X468 a_15320_100# N a_15140_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X469 a_4160_1500# P1 a_3980_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X470 P1 P2 a_7410_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X471 a_16590_100# N a_16410_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X472 a_8130_3380# N a_7950_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X473 a_19290_3380# X a_19110_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X474 a_14780_100# N a_14600_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X475 a_11730_1980# P0 a_11550_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X476 a_19110_1500# P1 a_18930_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X477 a_5960_1500# P1 a_5780_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X478 a_n340_3380# a_n620_3280# a_n520_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X479 VSSA Y a_12440_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X480 a_9930_3380# Y a_9750_3380# VSSA sky130_fd_pr__nfet_01v8 ad=4e+11p pd=2.8e+06u as=0p ps=0u w=1e+06u l=500000u
X481 a_10110_3380# Y a_9930_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X482 a_7770_3380# N P1 VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X483 a_12080_100# Y a_11900_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X484 VDDA a_21350_1400# a_22170_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X485 a_18750_1500# P1 a_18570_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X486 a_2720_1980# P1 a_2540_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X487 a_4160_100# X a_3980_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X488 a_740_1980# P1 a_560_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X489 a_20190_1500# P2 a_20010_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X490 a_16590_1500# P2 a_16410_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X491 VSSA Y a_11730_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X492 a_1100_3380# Z a_920_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=4e+11p ps=2.8e+06u w=1e+06u l=500000u
X493 a_21990_1500# a_21350_1400# a_21350_1400# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X494 a_15510_1980# P1 a_15330_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X495 VDDA P1 a_9560_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X496 N P2 a_13170_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X497 Z X a_1280_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X498 a_7580_1500# P2 a_7400_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X499 a_11190_1980# P2 a_11010_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X500 a_2900_3380# Z a_2720_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X501 a_920_3380# Z a_740_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X502 VDDA P1 a_20730_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X503 a_19470_100# Z a_19290_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X504 a_11720_1500# P2 a_11540_1500# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X505 a_9390_3380# Y a_9210_3380# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X506 a_20370_100# Z a_20190_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X507 a_12990_1980# P2 a_12810_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X508 a_4340_1980# P2 a_4160_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X509 a_n340_100# a_n620_70# a_n520_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X510 a_2180_1980# P2 a_2000_1980# VDDA sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X511 a_17310_100# N a_17130_100# VSSA sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
.ends

