magic
tech sky130A
timestamp 1637985873
<< metal2 >>
rect 4240 12635 4440 12640
rect 4240 12605 4245 12635
rect 4275 12605 4405 12635
rect 4435 12605 4440 12635
rect 4240 12600 4440 12605
rect 4480 12635 4680 12640
rect 4480 12605 4485 12635
rect 4515 12605 4645 12635
rect 4675 12605 4680 12635
rect 4480 12600 4680 12605
rect 4720 12635 5080 12640
rect 4720 12605 4725 12635
rect 4755 12605 4885 12635
rect 4915 12605 5045 12635
rect 5075 12605 5080 12635
rect 4720 12600 5080 12605
rect 5120 12635 5480 12640
rect 5120 12605 5125 12635
rect 5155 12605 5285 12635
rect 5315 12605 5445 12635
rect 5475 12605 5480 12635
rect 5120 12600 5480 12605
rect 5520 12635 5880 12640
rect 5520 12605 5525 12635
rect 5555 12605 5685 12635
rect 5715 12605 5845 12635
rect 5875 12605 5880 12635
rect 5520 12600 5880 12605
rect 5920 12635 6120 12640
rect 5920 12605 5925 12635
rect 5955 12605 6085 12635
rect 6115 12605 6120 12635
rect 5920 12600 6120 12605
rect 6160 12635 6360 12640
rect 6160 12605 6165 12635
rect 6195 12605 6325 12635
rect 6355 12605 6360 12635
rect 6160 12600 6360 12605
rect 4240 12555 4440 12560
rect 4240 12525 4245 12555
rect 4275 12525 4405 12555
rect 4435 12525 4440 12555
rect 4240 12520 4440 12525
rect 4480 12555 4680 12560
rect 4480 12525 4485 12555
rect 4515 12525 4645 12555
rect 4675 12525 4680 12555
rect 4480 12520 4680 12525
rect 4720 12555 5080 12560
rect 4720 12525 4725 12555
rect 4755 12525 4885 12555
rect 4915 12525 5045 12555
rect 5075 12525 5080 12555
rect 4720 12520 5080 12525
rect 5120 12555 5480 12560
rect 5120 12525 5125 12555
rect 5155 12525 5285 12555
rect 5315 12525 5445 12555
rect 5475 12525 5480 12555
rect 5120 12520 5480 12525
rect 5520 12555 5880 12560
rect 5520 12525 5525 12555
rect 5555 12525 5685 12555
rect 5715 12525 5845 12555
rect 5875 12525 5880 12555
rect 5520 12520 5880 12525
rect 5920 12555 6120 12560
rect 5920 12525 5925 12555
rect 5955 12525 6085 12555
rect 6115 12525 6120 12555
rect 5920 12520 6120 12525
rect 6160 12555 6360 12560
rect 6160 12525 6165 12555
rect 6195 12525 6325 12555
rect 6355 12525 6360 12555
rect 6160 12520 6360 12525
rect 4240 12475 4440 12480
rect 4240 12445 4245 12475
rect 4275 12445 4405 12475
rect 4435 12445 4440 12475
rect 4240 12440 4440 12445
rect 4480 12475 4680 12480
rect 4480 12445 4485 12475
rect 4515 12445 4645 12475
rect 4675 12445 4680 12475
rect 4480 12440 4680 12445
rect 4720 12475 5080 12480
rect 4720 12445 4725 12475
rect 4755 12445 4885 12475
rect 4915 12445 5045 12475
rect 5075 12445 5080 12475
rect 4720 12440 5080 12445
rect 5120 12475 5480 12480
rect 5120 12445 5125 12475
rect 5155 12445 5285 12475
rect 5315 12445 5445 12475
rect 5475 12445 5480 12475
rect 5120 12440 5480 12445
rect 5520 12475 5880 12480
rect 5520 12445 5525 12475
rect 5555 12445 5685 12475
rect 5715 12445 5845 12475
rect 5875 12445 5880 12475
rect 5520 12440 5880 12445
rect 5920 12475 6120 12480
rect 5920 12445 5925 12475
rect 5955 12445 6085 12475
rect 6115 12445 6120 12475
rect 5920 12440 6120 12445
rect 6160 12475 6360 12480
rect 6160 12445 6165 12475
rect 6195 12445 6325 12475
rect 6355 12445 6360 12475
rect 6160 12440 6360 12445
rect 4240 12395 4440 12400
rect 4240 12365 4245 12395
rect 4275 12365 4405 12395
rect 4435 12365 4440 12395
rect 4240 12360 4440 12365
rect 4480 12395 4680 12400
rect 4480 12365 4485 12395
rect 4515 12365 4645 12395
rect 4675 12365 4680 12395
rect 4480 12360 4680 12365
rect 4720 12395 5080 12400
rect 4720 12365 4725 12395
rect 4755 12365 4885 12395
rect 4915 12365 5045 12395
rect 5075 12365 5080 12395
rect 4720 12360 5080 12365
rect 5120 12395 5480 12400
rect 5120 12365 5125 12395
rect 5155 12365 5285 12395
rect 5315 12365 5445 12395
rect 5475 12365 5480 12395
rect 5120 12360 5480 12365
rect 5520 12395 5880 12400
rect 5520 12365 5525 12395
rect 5555 12365 5685 12395
rect 5715 12365 5845 12395
rect 5875 12365 5880 12395
rect 5520 12360 5880 12365
rect 5920 12395 6120 12400
rect 5920 12365 5925 12395
rect 5955 12365 6085 12395
rect 6115 12365 6120 12395
rect 5920 12360 6120 12365
rect 6160 12395 6360 12400
rect 6160 12365 6165 12395
rect 6195 12365 6325 12395
rect 6355 12365 6360 12395
rect 6160 12360 6360 12365
rect 4240 12315 4440 12320
rect 4240 12285 4245 12315
rect 4275 12285 4405 12315
rect 4435 12285 4440 12315
rect 4240 12280 4440 12285
rect 4480 12315 4680 12320
rect 4480 12285 4485 12315
rect 4515 12285 4645 12315
rect 4675 12285 4680 12315
rect 4480 12280 4680 12285
rect 4720 12315 5080 12320
rect 4720 12285 4725 12315
rect 4755 12285 4885 12315
rect 4915 12285 5045 12315
rect 5075 12285 5080 12315
rect 4720 12280 5080 12285
rect 5120 12315 5480 12320
rect 5120 12285 5125 12315
rect 5155 12285 5285 12315
rect 5315 12285 5445 12315
rect 5475 12285 5480 12315
rect 5120 12280 5480 12285
rect 5520 12315 5880 12320
rect 5520 12285 5525 12315
rect 5555 12285 5685 12315
rect 5715 12285 5845 12315
rect 5875 12285 5880 12315
rect 5520 12280 5880 12285
rect 5920 12315 6120 12320
rect 5920 12285 5925 12315
rect 5955 12285 6085 12315
rect 6115 12285 6120 12315
rect 5920 12280 6120 12285
rect 6160 12315 6360 12320
rect 6160 12285 6165 12315
rect 6195 12285 6325 12315
rect 6355 12285 6360 12315
rect 6160 12280 6360 12285
rect 4240 12235 4440 12240
rect 4240 12205 4245 12235
rect 4275 12205 4405 12235
rect 4435 12205 4440 12235
rect 4240 12200 4440 12205
rect 4480 12235 4680 12240
rect 4480 12205 4485 12235
rect 4515 12205 4645 12235
rect 4675 12205 4680 12235
rect 4480 12200 4680 12205
rect 4720 12235 5080 12240
rect 4720 12205 4725 12235
rect 4755 12205 4885 12235
rect 4915 12205 5045 12235
rect 5075 12205 5080 12235
rect 4720 12200 5080 12205
rect 5120 12235 5480 12240
rect 5120 12205 5125 12235
rect 5155 12205 5285 12235
rect 5315 12205 5445 12235
rect 5475 12205 5480 12235
rect 5120 12200 5480 12205
rect 5520 12235 5880 12240
rect 5520 12205 5525 12235
rect 5555 12205 5685 12235
rect 5715 12205 5845 12235
rect 5875 12205 5880 12235
rect 5520 12200 5880 12205
rect 5920 12235 6120 12240
rect 5920 12205 5925 12235
rect 5955 12205 6085 12235
rect 6115 12205 6120 12235
rect 5920 12200 6120 12205
rect 6160 12235 6360 12240
rect 6160 12205 6165 12235
rect 6195 12205 6325 12235
rect 6355 12205 6360 12235
rect 6160 12200 6360 12205
rect 4240 12155 4440 12160
rect 4240 12125 4245 12155
rect 4275 12125 4405 12155
rect 4435 12125 4440 12155
rect 4240 12120 4440 12125
rect 4480 12155 4680 12160
rect 4480 12125 4485 12155
rect 4515 12125 4645 12155
rect 4675 12125 4680 12155
rect 4480 12120 4680 12125
rect 4720 12155 5080 12160
rect 4720 12125 4725 12155
rect 4755 12125 4885 12155
rect 4915 12125 5045 12155
rect 5075 12125 5080 12155
rect 4720 12120 5080 12125
rect 5120 12155 5480 12160
rect 5120 12125 5125 12155
rect 5155 12125 5285 12155
rect 5315 12125 5445 12155
rect 5475 12125 5480 12155
rect 5120 12120 5480 12125
rect 5520 12155 5880 12160
rect 5520 12125 5525 12155
rect 5555 12125 5685 12155
rect 5715 12125 5845 12155
rect 5875 12125 5880 12155
rect 5520 12120 5880 12125
rect 5920 12155 6120 12160
rect 5920 12125 5925 12155
rect 5955 12125 6085 12155
rect 6115 12125 6120 12155
rect 5920 12120 6120 12125
rect 6160 12155 6360 12160
rect 6160 12125 6165 12155
rect 6195 12125 6325 12155
rect 6355 12125 6360 12155
rect 6160 12120 6360 12125
rect 4200 12075 6400 12080
rect 4200 12045 4485 12075
rect 4515 12045 4645 12075
rect 4675 12045 6400 12075
rect 4200 12040 6400 12045
rect 4200 11995 6400 12000
rect 4200 11965 4565 11995
rect 4595 11965 6400 11995
rect 4200 11960 6400 11965
rect 4200 11915 6400 11920
rect 4200 11885 4485 11915
rect 4515 11885 4645 11915
rect 4675 11885 6400 11915
rect 4200 11880 6400 11885
rect 4240 11835 4440 11840
rect 4240 11805 4245 11835
rect 4275 11805 4405 11835
rect 4435 11805 4440 11835
rect 4240 11800 4440 11805
rect 4480 11835 4680 11840
rect 4480 11805 4485 11835
rect 4515 11805 4645 11835
rect 4675 11805 4680 11835
rect 4480 11800 4680 11805
rect 4720 11835 5080 11840
rect 4720 11805 4725 11835
rect 4755 11805 4885 11835
rect 4915 11805 5045 11835
rect 5075 11805 5080 11835
rect 4720 11800 5080 11805
rect 5120 11835 5480 11840
rect 5120 11805 5125 11835
rect 5155 11805 5285 11835
rect 5315 11805 5445 11835
rect 5475 11805 5480 11835
rect 5120 11800 5480 11805
rect 5520 11835 5880 11840
rect 5520 11805 5525 11835
rect 5555 11805 5685 11835
rect 5715 11805 5845 11835
rect 5875 11805 5880 11835
rect 5520 11800 5880 11805
rect 5920 11835 6120 11840
rect 5920 11805 5925 11835
rect 5955 11805 6085 11835
rect 6115 11805 6120 11835
rect 5920 11800 6120 11805
rect 6160 11835 6360 11840
rect 6160 11805 6165 11835
rect 6195 11805 6325 11835
rect 6355 11805 6360 11835
rect 6160 11800 6360 11805
rect 4240 11755 4440 11760
rect 4240 11725 4245 11755
rect 4275 11725 4405 11755
rect 4435 11725 4440 11755
rect 4240 11720 4440 11725
rect 4480 11755 4680 11760
rect 4480 11725 4485 11755
rect 4515 11725 4645 11755
rect 4675 11725 4680 11755
rect 4480 11720 4680 11725
rect 4720 11755 5080 11760
rect 4720 11725 4725 11755
rect 4755 11725 4885 11755
rect 4915 11725 5045 11755
rect 5075 11725 5080 11755
rect 4720 11720 5080 11725
rect 5120 11755 5480 11760
rect 5120 11725 5125 11755
rect 5155 11725 5285 11755
rect 5315 11725 5445 11755
rect 5475 11725 5480 11755
rect 5120 11720 5480 11725
rect 5520 11755 5880 11760
rect 5520 11725 5525 11755
rect 5555 11725 5685 11755
rect 5715 11725 5845 11755
rect 5875 11725 5880 11755
rect 5520 11720 5880 11725
rect 5920 11755 6120 11760
rect 5920 11725 5925 11755
rect 5955 11725 6085 11755
rect 6115 11725 6120 11755
rect 5920 11720 6120 11725
rect 6160 11755 6360 11760
rect 6160 11725 6165 11755
rect 6195 11725 6325 11755
rect 6355 11725 6360 11755
rect 6160 11720 6360 11725
rect 4240 11675 4440 11680
rect 4240 11645 4245 11675
rect 4275 11645 4405 11675
rect 4435 11645 4440 11675
rect 4240 11640 4440 11645
rect 4480 11675 4680 11680
rect 4480 11645 4485 11675
rect 4515 11645 4645 11675
rect 4675 11645 4680 11675
rect 4480 11640 4680 11645
rect 4720 11675 5080 11680
rect 4720 11645 4725 11675
rect 4755 11645 4885 11675
rect 4915 11645 5045 11675
rect 5075 11645 5080 11675
rect 4720 11640 5080 11645
rect 5120 11675 5480 11680
rect 5120 11645 5125 11675
rect 5155 11645 5285 11675
rect 5315 11645 5445 11675
rect 5475 11645 5480 11675
rect 5120 11640 5480 11645
rect 5520 11675 5880 11680
rect 5520 11645 5525 11675
rect 5555 11645 5685 11675
rect 5715 11645 5845 11675
rect 5875 11645 5880 11675
rect 5520 11640 5880 11645
rect 5920 11675 6120 11680
rect 5920 11645 5925 11675
rect 5955 11645 6085 11675
rect 6115 11645 6120 11675
rect 5920 11640 6120 11645
rect 6160 11675 6360 11680
rect 6160 11645 6165 11675
rect 6195 11645 6325 11675
rect 6355 11645 6360 11675
rect 6160 11640 6360 11645
rect 4240 11595 4440 11600
rect 4240 11565 4245 11595
rect 4275 11565 4405 11595
rect 4435 11565 4440 11595
rect 4240 11560 4440 11565
rect 4480 11595 4680 11600
rect 4480 11565 4485 11595
rect 4515 11565 4645 11595
rect 4675 11565 4680 11595
rect 4480 11560 4680 11565
rect 4720 11595 5080 11600
rect 4720 11565 4725 11595
rect 4755 11565 4885 11595
rect 4915 11565 5045 11595
rect 5075 11565 5080 11595
rect 4720 11560 5080 11565
rect 5120 11595 5480 11600
rect 5120 11565 5125 11595
rect 5155 11565 5285 11595
rect 5315 11565 5445 11595
rect 5475 11565 5480 11595
rect 5120 11560 5480 11565
rect 5520 11595 5880 11600
rect 5520 11565 5525 11595
rect 5555 11565 5685 11595
rect 5715 11565 5845 11595
rect 5875 11565 5880 11595
rect 5520 11560 5880 11565
rect 5920 11595 6120 11600
rect 5920 11565 5925 11595
rect 5955 11565 6085 11595
rect 6115 11565 6120 11595
rect 5920 11560 6120 11565
rect 6160 11595 6360 11600
rect 6160 11565 6165 11595
rect 6195 11565 6325 11595
rect 6355 11565 6360 11595
rect 6160 11560 6360 11565
rect 4240 11515 4440 11520
rect 4240 11485 4245 11515
rect 4275 11485 4405 11515
rect 4435 11485 4440 11515
rect 4240 11480 4440 11485
rect 4480 11515 4680 11520
rect 4480 11485 4485 11515
rect 4515 11485 4645 11515
rect 4675 11485 4680 11515
rect 4480 11480 4680 11485
rect 4720 11515 5080 11520
rect 4720 11485 4725 11515
rect 4755 11485 4885 11515
rect 4915 11485 5045 11515
rect 5075 11485 5080 11515
rect 4720 11480 5080 11485
rect 5120 11515 5480 11520
rect 5120 11485 5125 11515
rect 5155 11485 5285 11515
rect 5315 11485 5445 11515
rect 5475 11485 5480 11515
rect 5120 11480 5480 11485
rect 5520 11515 5880 11520
rect 5520 11485 5525 11515
rect 5555 11485 5685 11515
rect 5715 11485 5845 11515
rect 5875 11485 5880 11515
rect 5520 11480 5880 11485
rect 5920 11515 6120 11520
rect 5920 11485 5925 11515
rect 5955 11485 6085 11515
rect 6115 11485 6120 11515
rect 5920 11480 6120 11485
rect 6160 11515 6360 11520
rect 6160 11485 6165 11515
rect 6195 11485 6325 11515
rect 6355 11485 6360 11515
rect 6160 11480 6360 11485
rect 4240 11435 4440 11440
rect 4240 11405 4245 11435
rect 4275 11405 4405 11435
rect 4435 11405 4440 11435
rect 4240 11400 4440 11405
rect 4480 11435 4680 11440
rect 4480 11405 4485 11435
rect 4515 11405 4645 11435
rect 4675 11405 4680 11435
rect 4480 11400 4680 11405
rect 4720 11435 5080 11440
rect 4720 11405 4725 11435
rect 4755 11405 4885 11435
rect 4915 11405 5045 11435
rect 5075 11405 5080 11435
rect 4720 11400 5080 11405
rect 5120 11435 5480 11440
rect 5120 11405 5125 11435
rect 5155 11405 5285 11435
rect 5315 11405 5445 11435
rect 5475 11405 5480 11435
rect 5120 11400 5480 11405
rect 5520 11435 5880 11440
rect 5520 11405 5525 11435
rect 5555 11405 5685 11435
rect 5715 11405 5845 11435
rect 5875 11405 5880 11435
rect 5520 11400 5880 11405
rect 5920 11435 6120 11440
rect 5920 11405 5925 11435
rect 5955 11405 6085 11435
rect 6115 11405 6120 11435
rect 5920 11400 6120 11405
rect 6160 11435 6360 11440
rect 6160 11405 6165 11435
rect 6195 11405 6325 11435
rect 6355 11405 6360 11435
rect 6160 11400 6360 11405
rect 4200 11315 6400 11320
rect 4200 11285 5525 11315
rect 5555 11285 5685 11315
rect 5715 11285 6400 11315
rect 4200 11280 6400 11285
rect 4200 11235 6400 11240
rect 4200 11205 5605 11235
rect 5635 11205 6400 11235
rect 4200 11200 6400 11205
rect 4200 11155 6400 11160
rect 4200 11125 5045 11155
rect 5075 11125 5525 11155
rect 5555 11125 5685 11155
rect 5715 11125 6400 11155
rect 4200 11120 6400 11125
rect 4200 11075 6400 11080
rect 4200 11045 5125 11075
rect 5155 11045 5285 11075
rect 5315 11045 5445 11075
rect 5475 11045 6400 11075
rect 4200 11040 6400 11045
rect 4200 10995 6400 11000
rect 4200 10965 5045 10995
rect 5075 10965 5525 10995
rect 5555 10965 6400 10995
rect 4200 10960 6400 10965
rect 4240 10875 4440 10880
rect 4240 10845 4245 10875
rect 4275 10845 4405 10875
rect 4435 10845 4440 10875
rect 4240 10840 4440 10845
rect 4480 10875 4680 10880
rect 4480 10845 4485 10875
rect 4515 10845 4645 10875
rect 4675 10845 4680 10875
rect 4480 10840 4680 10845
rect 4720 10875 5080 10880
rect 4720 10845 4725 10875
rect 4755 10845 4885 10875
rect 4915 10845 5045 10875
rect 5075 10845 5080 10875
rect 4720 10840 5080 10845
rect 5120 10875 5480 10880
rect 5120 10845 5125 10875
rect 5155 10845 5285 10875
rect 5315 10845 5445 10875
rect 5475 10845 5480 10875
rect 5120 10840 5480 10845
rect 5520 10875 5880 10880
rect 5520 10845 5525 10875
rect 5555 10845 5685 10875
rect 5715 10845 5845 10875
rect 5875 10845 5880 10875
rect 5520 10840 5880 10845
rect 5920 10875 6120 10880
rect 5920 10845 5925 10875
rect 5955 10845 6085 10875
rect 6115 10845 6120 10875
rect 5920 10840 6120 10845
rect 6160 10875 6360 10880
rect 6160 10845 6165 10875
rect 6195 10845 6325 10875
rect 6355 10845 6360 10875
rect 6160 10840 6360 10845
rect 4240 10795 4440 10800
rect 4240 10765 4245 10795
rect 4275 10765 4405 10795
rect 4435 10765 4440 10795
rect 4240 10760 4440 10765
rect 4480 10795 4680 10800
rect 4480 10765 4485 10795
rect 4515 10765 4645 10795
rect 4675 10765 4680 10795
rect 4480 10760 4680 10765
rect 4720 10795 5080 10800
rect 4720 10765 4725 10795
rect 4755 10765 4885 10795
rect 4915 10765 5045 10795
rect 5075 10765 5080 10795
rect 4720 10760 5080 10765
rect 5120 10795 5480 10800
rect 5120 10765 5125 10795
rect 5155 10765 5285 10795
rect 5315 10765 5445 10795
rect 5475 10765 5480 10795
rect 5120 10760 5480 10765
rect 5520 10795 5880 10800
rect 5520 10765 5525 10795
rect 5555 10765 5685 10795
rect 5715 10765 5845 10795
rect 5875 10765 5880 10795
rect 5520 10760 5880 10765
rect 5920 10795 6120 10800
rect 5920 10765 5925 10795
rect 5955 10765 6085 10795
rect 6115 10765 6120 10795
rect 5920 10760 6120 10765
rect 6160 10795 6360 10800
rect 6160 10765 6165 10795
rect 6195 10765 6325 10795
rect 6355 10765 6360 10795
rect 6160 10760 6360 10765
rect 4240 10715 4440 10720
rect 4240 10685 4245 10715
rect 4275 10685 4405 10715
rect 4435 10685 4440 10715
rect 4240 10680 4440 10685
rect 4480 10715 4680 10720
rect 4480 10685 4485 10715
rect 4515 10685 4645 10715
rect 4675 10685 4680 10715
rect 4480 10680 4680 10685
rect 4720 10715 5080 10720
rect 4720 10685 4725 10715
rect 4755 10685 4885 10715
rect 4915 10685 5045 10715
rect 5075 10685 5080 10715
rect 4720 10680 5080 10685
rect 5120 10715 5480 10720
rect 5120 10685 5125 10715
rect 5155 10685 5285 10715
rect 5315 10685 5445 10715
rect 5475 10685 5480 10715
rect 5120 10680 5480 10685
rect 5520 10715 5880 10720
rect 5520 10685 5525 10715
rect 5555 10685 5685 10715
rect 5715 10685 5845 10715
rect 5875 10685 5880 10715
rect 5520 10680 5880 10685
rect 5920 10715 6120 10720
rect 5920 10685 5925 10715
rect 5955 10685 6085 10715
rect 6115 10685 6120 10715
rect 5920 10680 6120 10685
rect 6160 10715 6360 10720
rect 6160 10685 6165 10715
rect 6195 10685 6325 10715
rect 6355 10685 6360 10715
rect 6160 10680 6360 10685
rect 4240 10635 4440 10640
rect 4240 10605 4245 10635
rect 4275 10605 4405 10635
rect 4435 10605 4440 10635
rect 4240 10600 4440 10605
rect 4480 10635 4680 10640
rect 4480 10605 4485 10635
rect 4515 10605 4645 10635
rect 4675 10605 4680 10635
rect 4480 10600 4680 10605
rect 4720 10635 5080 10640
rect 4720 10605 4725 10635
rect 4755 10605 4885 10635
rect 4915 10605 5045 10635
rect 5075 10605 5080 10635
rect 4720 10600 5080 10605
rect 5120 10635 5480 10640
rect 5120 10605 5125 10635
rect 5155 10605 5285 10635
rect 5315 10605 5445 10635
rect 5475 10605 5480 10635
rect 5120 10600 5480 10605
rect 5520 10635 5880 10640
rect 5520 10605 5525 10635
rect 5555 10605 5685 10635
rect 5715 10605 5845 10635
rect 5875 10605 5880 10635
rect 5520 10600 5880 10605
rect 5920 10635 6120 10640
rect 5920 10605 5925 10635
rect 5955 10605 6085 10635
rect 6115 10605 6120 10635
rect 5920 10600 6120 10605
rect 6160 10635 6360 10640
rect 6160 10605 6165 10635
rect 6195 10605 6325 10635
rect 6355 10605 6360 10635
rect 6160 10600 6360 10605
rect 4240 10555 4440 10560
rect 4240 10525 4245 10555
rect 4275 10525 4405 10555
rect 4435 10525 4440 10555
rect 4240 10520 4440 10525
rect 4480 10555 4680 10560
rect 4480 10525 4485 10555
rect 4515 10525 4645 10555
rect 4675 10525 4680 10555
rect 4480 10520 4680 10525
rect 4720 10555 5080 10560
rect 4720 10525 4725 10555
rect 4755 10525 4885 10555
rect 4915 10525 5045 10555
rect 5075 10525 5080 10555
rect 4720 10520 5080 10525
rect 5120 10555 5480 10560
rect 5120 10525 5125 10555
rect 5155 10525 5285 10555
rect 5315 10525 5445 10555
rect 5475 10525 5480 10555
rect 5120 10520 5480 10525
rect 5520 10555 5880 10560
rect 5520 10525 5525 10555
rect 5555 10525 5685 10555
rect 5715 10525 5845 10555
rect 5875 10525 5880 10555
rect 5520 10520 5880 10525
rect 5920 10555 6120 10560
rect 5920 10525 5925 10555
rect 5955 10525 6085 10555
rect 6115 10525 6120 10555
rect 5920 10520 6120 10525
rect 6160 10555 6360 10560
rect 6160 10525 6165 10555
rect 6195 10525 6325 10555
rect 6355 10525 6360 10555
rect 6160 10520 6360 10525
rect 4240 10475 4440 10480
rect 4240 10445 4245 10475
rect 4275 10445 4405 10475
rect 4435 10445 4440 10475
rect 4240 10440 4440 10445
rect 4480 10475 4680 10480
rect 4480 10445 4485 10475
rect 4515 10445 4645 10475
rect 4675 10445 4680 10475
rect 4480 10440 4680 10445
rect 4720 10475 5080 10480
rect 4720 10445 4725 10475
rect 4755 10445 4885 10475
rect 4915 10445 5045 10475
rect 5075 10445 5080 10475
rect 4720 10440 5080 10445
rect 5120 10475 5480 10480
rect 5120 10445 5125 10475
rect 5155 10445 5285 10475
rect 5315 10445 5445 10475
rect 5475 10445 5480 10475
rect 5120 10440 5480 10445
rect 5520 10475 5880 10480
rect 5520 10445 5525 10475
rect 5555 10445 5685 10475
rect 5715 10445 5845 10475
rect 5875 10445 5880 10475
rect 5520 10440 5880 10445
rect 5920 10475 6120 10480
rect 5920 10445 5925 10475
rect 5955 10445 6085 10475
rect 6115 10445 6120 10475
rect 5920 10440 6120 10445
rect 6160 10475 6360 10480
rect 6160 10445 6165 10475
rect 6195 10445 6325 10475
rect 6355 10445 6360 10475
rect 6160 10440 6360 10445
rect 4240 10395 4440 10400
rect 4240 10365 4245 10395
rect 4275 10365 4405 10395
rect 4435 10365 4440 10395
rect 4240 10360 4440 10365
rect 4480 10395 4680 10400
rect 4480 10365 4485 10395
rect 4515 10365 4645 10395
rect 4675 10365 4680 10395
rect 4480 10360 4680 10365
rect 4720 10395 5080 10400
rect 4720 10365 4725 10395
rect 4755 10365 4885 10395
rect 4915 10365 5045 10395
rect 5075 10365 5080 10395
rect 4720 10360 5080 10365
rect 5120 10395 5480 10400
rect 5120 10365 5125 10395
rect 5155 10365 5285 10395
rect 5315 10365 5445 10395
rect 5475 10365 5480 10395
rect 5120 10360 5480 10365
rect 5520 10395 5880 10400
rect 5520 10365 5525 10395
rect 5555 10365 5685 10395
rect 5715 10365 5845 10395
rect 5875 10365 5880 10395
rect 5520 10360 5880 10365
rect 5920 10395 6120 10400
rect 5920 10365 5925 10395
rect 5955 10365 6085 10395
rect 6115 10365 6120 10395
rect 5920 10360 6120 10365
rect 6160 10395 6360 10400
rect 6160 10365 6165 10395
rect 6195 10365 6325 10395
rect 6355 10365 6360 10395
rect 6160 10360 6360 10365
rect 4240 10315 4440 10320
rect 4240 10285 4245 10315
rect 4275 10285 4405 10315
rect 4435 10285 4440 10315
rect 4240 10280 4440 10285
rect 4480 10315 4680 10320
rect 4480 10285 4485 10315
rect 4515 10285 4645 10315
rect 4675 10285 4680 10315
rect 4480 10280 4680 10285
rect 4720 10315 5080 10320
rect 4720 10285 4725 10315
rect 4755 10285 4885 10315
rect 4915 10285 5045 10315
rect 5075 10285 5080 10315
rect 4720 10280 5080 10285
rect 5120 10315 5480 10320
rect 5120 10285 5125 10315
rect 5155 10285 5285 10315
rect 5315 10285 5445 10315
rect 5475 10285 5480 10315
rect 5120 10280 5480 10285
rect 5520 10315 5880 10320
rect 5520 10285 5525 10315
rect 5555 10285 5685 10315
rect 5715 10285 5845 10315
rect 5875 10285 5880 10315
rect 5520 10280 5880 10285
rect 5920 10315 6120 10320
rect 5920 10285 5925 10315
rect 5955 10285 6085 10315
rect 6115 10285 6120 10315
rect 5920 10280 6120 10285
rect 6160 10315 6360 10320
rect 6160 10285 6165 10315
rect 6195 10285 6325 10315
rect 6355 10285 6360 10315
rect 6160 10280 6360 10285
rect 4240 10235 4440 10240
rect 4240 10205 4245 10235
rect 4275 10205 4405 10235
rect 4435 10205 4440 10235
rect 4240 10200 4440 10205
rect 4480 10235 4680 10240
rect 4480 10205 4485 10235
rect 4515 10205 4645 10235
rect 4675 10205 4680 10235
rect 4480 10200 4680 10205
rect 4720 10235 5080 10240
rect 4720 10205 4725 10235
rect 4755 10205 4885 10235
rect 4915 10205 5045 10235
rect 5075 10205 5080 10235
rect 4720 10200 5080 10205
rect 5120 10235 5480 10240
rect 5120 10205 5125 10235
rect 5155 10205 5285 10235
rect 5315 10205 5445 10235
rect 5475 10205 5480 10235
rect 5120 10200 5480 10205
rect 5520 10235 5880 10240
rect 5520 10205 5525 10235
rect 5555 10205 5685 10235
rect 5715 10205 5845 10235
rect 5875 10205 5880 10235
rect 5520 10200 5880 10205
rect 5920 10235 6120 10240
rect 5920 10205 5925 10235
rect 5955 10205 6085 10235
rect 6115 10205 6120 10235
rect 5920 10200 6120 10205
rect 6160 10235 6360 10240
rect 6160 10205 6165 10235
rect 6195 10205 6325 10235
rect 6355 10205 6360 10235
rect 6160 10200 6360 10205
rect 4240 10155 4440 10160
rect 4240 10125 4245 10155
rect 4275 10125 4405 10155
rect 4435 10125 4440 10155
rect 4240 10120 4440 10125
rect 4480 10155 4680 10160
rect 4480 10125 4485 10155
rect 4515 10125 4645 10155
rect 4675 10125 4680 10155
rect 4480 10120 4680 10125
rect 4720 10155 5080 10160
rect 4720 10125 4725 10155
rect 4755 10125 4885 10155
rect 4915 10125 5045 10155
rect 5075 10125 5080 10155
rect 4720 10120 5080 10125
rect 5120 10155 5480 10160
rect 5120 10125 5125 10155
rect 5155 10125 5285 10155
rect 5315 10125 5445 10155
rect 5475 10125 5480 10155
rect 5120 10120 5480 10125
rect 5520 10155 5880 10160
rect 5520 10125 5525 10155
rect 5555 10125 5685 10155
rect 5715 10125 5845 10155
rect 5875 10125 5880 10155
rect 5520 10120 5880 10125
rect 5920 10155 6120 10160
rect 5920 10125 5925 10155
rect 5955 10125 6085 10155
rect 6115 10125 6120 10155
rect 5920 10120 6120 10125
rect 6160 10155 6360 10160
rect 6160 10125 6165 10155
rect 6195 10125 6325 10155
rect 6355 10125 6360 10155
rect 6160 10120 6360 10125
rect 4240 10075 4440 10080
rect 4240 10045 4245 10075
rect 4275 10045 4405 10075
rect 4435 10045 4440 10075
rect 4240 10040 4440 10045
rect 4480 10075 4680 10080
rect 4480 10045 4485 10075
rect 4515 10045 4645 10075
rect 4675 10045 4680 10075
rect 4480 10040 4680 10045
rect 4720 10075 5080 10080
rect 4720 10045 4725 10075
rect 4755 10045 4885 10075
rect 4915 10045 5045 10075
rect 5075 10045 5080 10075
rect 4720 10040 5080 10045
rect 5120 10075 5480 10080
rect 5120 10045 5125 10075
rect 5155 10045 5285 10075
rect 5315 10045 5445 10075
rect 5475 10045 5480 10075
rect 5120 10040 5480 10045
rect 5520 10075 5880 10080
rect 5520 10045 5525 10075
rect 5555 10045 5685 10075
rect 5715 10045 5845 10075
rect 5875 10045 5880 10075
rect 5520 10040 5880 10045
rect 5920 10075 6120 10080
rect 5920 10045 5925 10075
rect 5955 10045 6085 10075
rect 6115 10045 6120 10075
rect 5920 10040 6120 10045
rect 6160 10075 6360 10080
rect 6160 10045 6165 10075
rect 6195 10045 6325 10075
rect 6355 10045 6360 10075
rect 6160 10040 6360 10045
rect 4240 9995 4440 10000
rect 4240 9965 4245 9995
rect 4275 9965 4405 9995
rect 4435 9965 4440 9995
rect 4240 9960 4440 9965
rect 4480 9995 4680 10000
rect 4480 9965 4485 9995
rect 4515 9965 4645 9995
rect 4675 9965 4680 9995
rect 4480 9960 4680 9965
rect 4720 9995 5080 10000
rect 4720 9965 4725 9995
rect 4755 9965 4885 9995
rect 4915 9965 5045 9995
rect 5075 9965 5080 9995
rect 4720 9960 5080 9965
rect 5120 9995 5480 10000
rect 5120 9965 5125 9995
rect 5155 9965 5285 9995
rect 5315 9965 5445 9995
rect 5475 9965 5480 9995
rect 5120 9960 5480 9965
rect 5520 9995 5880 10000
rect 5520 9965 5525 9995
rect 5555 9965 5685 9995
rect 5715 9965 5845 9995
rect 5875 9965 5880 9995
rect 5520 9960 5880 9965
rect 5920 9995 6120 10000
rect 5920 9965 5925 9995
rect 5955 9965 6085 9995
rect 6115 9965 6120 9995
rect 5920 9960 6120 9965
rect 6160 9995 6360 10000
rect 6160 9965 6165 9995
rect 6195 9965 6325 9995
rect 6355 9965 6360 9995
rect 6160 9960 6360 9965
rect 4240 9915 4440 9920
rect 4240 9885 4245 9915
rect 4275 9885 4405 9915
rect 4435 9885 4440 9915
rect 4240 9880 4440 9885
rect 4480 9915 4680 9920
rect 4480 9885 4485 9915
rect 4515 9885 4645 9915
rect 4675 9885 4680 9915
rect 4480 9880 4680 9885
rect 4720 9915 5080 9920
rect 4720 9885 4725 9915
rect 4755 9885 4885 9915
rect 4915 9885 5045 9915
rect 5075 9885 5080 9915
rect 4720 9880 5080 9885
rect 5120 9915 5480 9920
rect 5120 9885 5125 9915
rect 5155 9885 5285 9915
rect 5315 9885 5445 9915
rect 5475 9885 5480 9915
rect 5120 9880 5480 9885
rect 5520 9915 5880 9920
rect 5520 9885 5525 9915
rect 5555 9885 5685 9915
rect 5715 9885 5845 9915
rect 5875 9885 5880 9915
rect 5520 9880 5880 9885
rect 5920 9915 6120 9920
rect 5920 9885 5925 9915
rect 5955 9885 6085 9915
rect 6115 9885 6120 9915
rect 5920 9880 6120 9885
rect 6160 9915 6360 9920
rect 6160 9885 6165 9915
rect 6195 9885 6325 9915
rect 6355 9885 6360 9915
rect 6160 9880 6360 9885
rect 4240 9835 4440 9840
rect 4240 9805 4245 9835
rect 4275 9805 4405 9835
rect 4435 9805 4440 9835
rect 4240 9800 4440 9805
rect 4480 9835 4680 9840
rect 4480 9805 4485 9835
rect 4515 9805 4645 9835
rect 4675 9805 4680 9835
rect 4480 9800 4680 9805
rect 4720 9835 5080 9840
rect 4720 9805 4725 9835
rect 4755 9805 4885 9835
rect 4915 9805 5045 9835
rect 5075 9805 5080 9835
rect 4720 9800 5080 9805
rect 5120 9835 5480 9840
rect 5120 9805 5125 9835
rect 5155 9805 5285 9835
rect 5315 9805 5445 9835
rect 5475 9805 5480 9835
rect 5120 9800 5480 9805
rect 5520 9835 5880 9840
rect 5520 9805 5525 9835
rect 5555 9805 5685 9835
rect 5715 9805 5845 9835
rect 5875 9805 5880 9835
rect 5520 9800 5880 9805
rect 5920 9835 6120 9840
rect 5920 9805 5925 9835
rect 5955 9805 6085 9835
rect 6115 9805 6120 9835
rect 5920 9800 6120 9805
rect 6160 9835 6360 9840
rect 6160 9805 6165 9835
rect 6195 9805 6325 9835
rect 6355 9805 6360 9835
rect 6160 9800 6360 9805
rect 4240 9755 4440 9760
rect 4240 9725 4245 9755
rect 4275 9725 4405 9755
rect 4435 9725 4440 9755
rect 4240 9720 4440 9725
rect 4480 9755 4680 9760
rect 4480 9725 4485 9755
rect 4515 9725 4645 9755
rect 4675 9725 4680 9755
rect 4480 9720 4680 9725
rect 4720 9755 5080 9760
rect 4720 9725 4725 9755
rect 4755 9725 4885 9755
rect 4915 9725 5045 9755
rect 5075 9725 5080 9755
rect 4720 9720 5080 9725
rect 5120 9755 5480 9760
rect 5120 9725 5125 9755
rect 5155 9725 5285 9755
rect 5315 9725 5445 9755
rect 5475 9725 5480 9755
rect 5120 9720 5480 9725
rect 5520 9755 5880 9760
rect 5520 9725 5525 9755
rect 5555 9725 5685 9755
rect 5715 9725 5845 9755
rect 5875 9725 5880 9755
rect 5520 9720 5880 9725
rect 5920 9755 6120 9760
rect 5920 9725 5925 9755
rect 5955 9725 6085 9755
rect 6115 9725 6120 9755
rect 5920 9720 6120 9725
rect 6160 9755 6360 9760
rect 6160 9725 6165 9755
rect 6195 9725 6325 9755
rect 6355 9725 6360 9755
rect 6160 9720 6360 9725
rect 4240 9635 6360 9640
rect 4240 9605 4485 9635
rect 4515 9605 4645 9635
rect 4675 9605 6360 9635
rect 4240 9600 6360 9605
rect 4200 9555 6400 9560
rect 4200 9525 4565 9555
rect 4595 9525 6400 9555
rect 4200 9520 6400 9525
rect 4240 9475 6360 9480
rect 4240 9445 4485 9475
rect 4515 9445 4645 9475
rect 4675 9445 6360 9475
rect 4240 9440 6360 9445
rect 4240 9355 4440 9360
rect 4240 9325 4245 9355
rect 4275 9325 4405 9355
rect 4435 9325 4440 9355
rect 4240 9320 4440 9325
rect 4480 9355 4680 9360
rect 4480 9325 4485 9355
rect 4515 9325 4645 9355
rect 4675 9325 4680 9355
rect 4480 9320 4680 9325
rect 4720 9355 5080 9360
rect 4720 9325 4725 9355
rect 4755 9325 4885 9355
rect 4915 9325 5045 9355
rect 5075 9325 5080 9355
rect 4720 9320 5080 9325
rect 5120 9355 5480 9360
rect 5120 9325 5125 9355
rect 5155 9325 5285 9355
rect 5315 9325 5445 9355
rect 5475 9325 5480 9355
rect 5120 9320 5480 9325
rect 5520 9355 5880 9360
rect 5520 9325 5525 9355
rect 5555 9325 5685 9355
rect 5715 9325 5845 9355
rect 5875 9325 5880 9355
rect 5520 9320 5880 9325
rect 5920 9355 6120 9360
rect 5920 9325 5925 9355
rect 5955 9325 6085 9355
rect 6115 9325 6120 9355
rect 5920 9320 6120 9325
rect 6160 9355 6360 9360
rect 6160 9325 6165 9355
rect 6195 9325 6325 9355
rect 6355 9325 6360 9355
rect 6160 9320 6360 9325
rect 4240 9275 4440 9280
rect 4240 9245 4245 9275
rect 4275 9245 4405 9275
rect 4435 9245 4440 9275
rect 4240 9240 4440 9245
rect 4480 9275 4680 9280
rect 4480 9245 4485 9275
rect 4515 9245 4645 9275
rect 4675 9245 4680 9275
rect 4480 9240 4680 9245
rect 4720 9275 5080 9280
rect 4720 9245 4725 9275
rect 4755 9245 4885 9275
rect 4915 9245 5045 9275
rect 5075 9245 5080 9275
rect 4720 9240 5080 9245
rect 5120 9275 5480 9280
rect 5120 9245 5125 9275
rect 5155 9245 5285 9275
rect 5315 9245 5445 9275
rect 5475 9245 5480 9275
rect 5120 9240 5480 9245
rect 5520 9275 5880 9280
rect 5520 9245 5525 9275
rect 5555 9245 5685 9275
rect 5715 9245 5845 9275
rect 5875 9245 5880 9275
rect 5520 9240 5880 9245
rect 5920 9275 6120 9280
rect 5920 9245 5925 9275
rect 5955 9245 6085 9275
rect 6115 9245 6120 9275
rect 5920 9240 6120 9245
rect 6160 9275 6360 9280
rect 6160 9245 6165 9275
rect 6195 9245 6325 9275
rect 6355 9245 6360 9275
rect 6160 9240 6360 9245
rect 4240 9195 4440 9200
rect 4240 9165 4245 9195
rect 4275 9165 4405 9195
rect 4435 9165 4440 9195
rect 4240 9160 4440 9165
rect 4480 9195 4680 9200
rect 4480 9165 4485 9195
rect 4515 9165 4645 9195
rect 4675 9165 4680 9195
rect 4480 9160 4680 9165
rect 4720 9195 5080 9200
rect 4720 9165 4725 9195
rect 4755 9165 4885 9195
rect 4915 9165 5045 9195
rect 5075 9165 5080 9195
rect 4720 9160 5080 9165
rect 5120 9195 5480 9200
rect 5120 9165 5125 9195
rect 5155 9165 5285 9195
rect 5315 9165 5445 9195
rect 5475 9165 5480 9195
rect 5120 9160 5480 9165
rect 5520 9195 5880 9200
rect 5520 9165 5525 9195
rect 5555 9165 5685 9195
rect 5715 9165 5845 9195
rect 5875 9165 5880 9195
rect 5520 9160 5880 9165
rect 5920 9195 6120 9200
rect 5920 9165 5925 9195
rect 5955 9165 6085 9195
rect 6115 9165 6120 9195
rect 5920 9160 6120 9165
rect 6160 9195 6360 9200
rect 6160 9165 6165 9195
rect 6195 9165 6325 9195
rect 6355 9165 6360 9195
rect 6160 9160 6360 9165
rect 4240 9115 6360 9120
rect 4240 9085 5125 9115
rect 5155 9085 5285 9115
rect 5315 9085 5445 9115
rect 5475 9085 6360 9115
rect 4240 9080 6360 9085
rect 4200 9035 6400 9040
rect 4200 9005 5365 9035
rect 5395 9005 6400 9035
rect 4200 9000 6400 9005
rect 4240 8955 6360 8960
rect 4240 8925 5125 8955
rect 5155 8925 5285 8955
rect 5315 8925 5445 8955
rect 5475 8925 6360 8955
rect 4240 8920 6360 8925
rect 4240 8875 4440 8880
rect 4240 8845 4245 8875
rect 4275 8845 4405 8875
rect 4435 8845 4440 8875
rect 4240 8840 4440 8845
rect 4480 8875 4680 8880
rect 4480 8845 4485 8875
rect 4515 8845 4645 8875
rect 4675 8845 4680 8875
rect 4480 8840 4680 8845
rect 4720 8875 5080 8880
rect 4720 8845 4725 8875
rect 4755 8845 4885 8875
rect 4915 8845 5045 8875
rect 5075 8845 5080 8875
rect 4720 8840 5080 8845
rect 5120 8875 5480 8880
rect 5120 8845 5125 8875
rect 5155 8845 5285 8875
rect 5315 8845 5445 8875
rect 5475 8845 5480 8875
rect 5120 8840 5480 8845
rect 5520 8875 5880 8880
rect 5520 8845 5525 8875
rect 5555 8845 5685 8875
rect 5715 8845 5845 8875
rect 5875 8845 5880 8875
rect 5520 8840 5880 8845
rect 5920 8875 6120 8880
rect 5920 8845 5925 8875
rect 5955 8845 6085 8875
rect 6115 8845 6120 8875
rect 5920 8840 6120 8845
rect 6160 8875 6360 8880
rect 6160 8845 6165 8875
rect 6195 8845 6325 8875
rect 6355 8845 6360 8875
rect 6160 8840 6360 8845
rect 4240 8795 4440 8800
rect 4240 8765 4245 8795
rect 4275 8765 4405 8795
rect 4435 8765 4440 8795
rect 4240 8760 4440 8765
rect 4480 8795 4680 8800
rect 4480 8765 4485 8795
rect 4515 8765 4645 8795
rect 4675 8765 4680 8795
rect 4480 8760 4680 8765
rect 4720 8795 5080 8800
rect 4720 8765 4725 8795
rect 4755 8765 4885 8795
rect 4915 8765 5045 8795
rect 5075 8765 5080 8795
rect 4720 8760 5080 8765
rect 5120 8795 5480 8800
rect 5120 8765 5125 8795
rect 5155 8765 5285 8795
rect 5315 8765 5445 8795
rect 5475 8765 5480 8795
rect 5120 8760 5480 8765
rect 5520 8795 5880 8800
rect 5520 8765 5525 8795
rect 5555 8765 5685 8795
rect 5715 8765 5845 8795
rect 5875 8765 5880 8795
rect 5520 8760 5880 8765
rect 5920 8795 6120 8800
rect 5920 8765 5925 8795
rect 5955 8765 6085 8795
rect 6115 8765 6120 8795
rect 5920 8760 6120 8765
rect 6160 8795 6360 8800
rect 6160 8765 6165 8795
rect 6195 8765 6325 8795
rect 6355 8765 6360 8795
rect 6160 8760 6360 8765
rect 4240 8715 4440 8720
rect 4240 8685 4245 8715
rect 4275 8685 4405 8715
rect 4435 8685 4440 8715
rect 4240 8680 4440 8685
rect 4480 8715 4680 8720
rect 4480 8685 4485 8715
rect 4515 8685 4645 8715
rect 4675 8685 4680 8715
rect 4480 8680 4680 8685
rect 4720 8715 5080 8720
rect 4720 8685 4725 8715
rect 4755 8685 4885 8715
rect 4915 8685 5045 8715
rect 5075 8685 5080 8715
rect 4720 8680 5080 8685
rect 5120 8715 5480 8720
rect 5120 8685 5125 8715
rect 5155 8685 5285 8715
rect 5315 8685 5445 8715
rect 5475 8685 5480 8715
rect 5120 8680 5480 8685
rect 5520 8715 5880 8720
rect 5520 8685 5525 8715
rect 5555 8685 5685 8715
rect 5715 8685 5845 8715
rect 5875 8685 5880 8715
rect 5520 8680 5880 8685
rect 5920 8715 6120 8720
rect 5920 8685 5925 8715
rect 5955 8685 6085 8715
rect 6115 8685 6120 8715
rect 5920 8680 6120 8685
rect 6160 8715 6360 8720
rect 6160 8685 6165 8715
rect 6195 8685 6325 8715
rect 6355 8685 6360 8715
rect 6160 8680 6360 8685
rect 4240 8635 4440 8640
rect 4240 8605 4245 8635
rect 4275 8605 4405 8635
rect 4435 8605 4440 8635
rect 4240 8600 4440 8605
rect 4480 8635 4680 8640
rect 4480 8605 4485 8635
rect 4515 8605 4645 8635
rect 4675 8605 4680 8635
rect 4480 8600 4680 8605
rect 4720 8635 5080 8640
rect 4720 8605 4725 8635
rect 4755 8605 4885 8635
rect 4915 8605 5045 8635
rect 5075 8605 5080 8635
rect 4720 8600 5080 8605
rect 5120 8635 5480 8640
rect 5120 8605 5125 8635
rect 5155 8605 5285 8635
rect 5315 8605 5445 8635
rect 5475 8605 5480 8635
rect 5120 8600 5480 8605
rect 5520 8635 5880 8640
rect 5520 8605 5525 8635
rect 5555 8605 5685 8635
rect 5715 8605 5845 8635
rect 5875 8605 5880 8635
rect 5520 8600 5880 8605
rect 5920 8635 6120 8640
rect 5920 8605 5925 8635
rect 5955 8605 6085 8635
rect 6115 8605 6120 8635
rect 5920 8600 6120 8605
rect 6160 8635 6360 8640
rect 6160 8605 6165 8635
rect 6195 8605 6325 8635
rect 6355 8605 6360 8635
rect 6160 8600 6360 8605
rect 4240 8555 4440 8560
rect 4240 8525 4245 8555
rect 4275 8525 4405 8555
rect 4435 8525 4440 8555
rect 4240 8520 4440 8525
rect 4480 8555 4680 8560
rect 4480 8525 4485 8555
rect 4515 8525 4645 8555
rect 4675 8525 4680 8555
rect 4480 8520 4680 8525
rect 4720 8555 5080 8560
rect 4720 8525 4725 8555
rect 4755 8525 4885 8555
rect 4915 8525 5045 8555
rect 5075 8525 5080 8555
rect 4720 8520 5080 8525
rect 5120 8555 5480 8560
rect 5120 8525 5125 8555
rect 5155 8525 5285 8555
rect 5315 8525 5445 8555
rect 5475 8525 5480 8555
rect 5120 8520 5480 8525
rect 5520 8555 5880 8560
rect 5520 8525 5525 8555
rect 5555 8525 5685 8555
rect 5715 8525 5845 8555
rect 5875 8525 5880 8555
rect 5520 8520 5880 8525
rect 5920 8555 6120 8560
rect 5920 8525 5925 8555
rect 5955 8525 6085 8555
rect 6115 8525 6120 8555
rect 5920 8520 6120 8525
rect 6160 8555 6360 8560
rect 6160 8525 6165 8555
rect 6195 8525 6325 8555
rect 6355 8525 6360 8555
rect 6160 8520 6360 8525
rect 4240 8475 6360 8480
rect 4240 8445 4885 8475
rect 4915 8445 5045 8475
rect 5075 8445 5685 8475
rect 5715 8445 5845 8475
rect 5875 8445 6360 8475
rect 4240 8440 6360 8445
rect 4200 8395 5000 8400
rect 4200 8365 4965 8395
rect 4995 8365 5000 8395
rect 4200 8360 5000 8365
rect 5760 8395 6400 8400
rect 5760 8365 5765 8395
rect 5795 8365 6400 8395
rect 5760 8360 6400 8365
rect 4240 8315 6360 8320
rect 4240 8285 4885 8315
rect 4915 8285 5045 8315
rect 5075 8285 5525 8315
rect 5555 8285 5685 8315
rect 5715 8285 5845 8315
rect 5875 8285 6360 8315
rect 4240 8280 6360 8285
rect 4200 8235 6400 8240
rect 4200 8205 5605 8235
rect 5635 8205 6400 8235
rect 4200 8200 6400 8205
rect 4240 8155 6360 8160
rect 4240 8125 5525 8155
rect 5555 8125 5685 8155
rect 5715 8125 6360 8155
rect 4240 8120 6360 8125
rect 4240 8075 6360 8080
rect 4240 8045 5045 8075
rect 5075 8045 5525 8075
rect 5555 8045 6360 8075
rect 4240 8040 6360 8045
rect 4240 7995 6360 8000
rect 4240 7965 5125 7995
rect 5155 7965 5285 7995
rect 5315 7965 5445 7995
rect 5475 7965 6360 7995
rect 4240 7960 6360 7965
rect 4200 7915 6400 7920
rect 4200 7885 5205 7915
rect 5235 7885 6400 7915
rect 4200 7880 6400 7885
rect 4240 7835 6360 7840
rect 4240 7805 5125 7835
rect 5155 7805 5285 7835
rect 5315 7805 5445 7835
rect 5475 7805 6360 7835
rect 4240 7800 6360 7805
rect 4240 7755 6360 7760
rect 4240 7725 5045 7755
rect 5075 7725 5525 7755
rect 5555 7725 6360 7755
rect 4240 7720 6360 7725
rect 4240 7635 4440 7640
rect 4240 7605 4245 7635
rect 4275 7605 4405 7635
rect 4435 7605 4440 7635
rect 4240 7600 4440 7605
rect 4480 7635 4680 7640
rect 4480 7605 4485 7635
rect 4515 7605 4645 7635
rect 4675 7605 4680 7635
rect 4480 7600 4680 7605
rect 4720 7635 5080 7640
rect 4720 7605 4725 7635
rect 4755 7605 4885 7635
rect 4915 7605 5045 7635
rect 5075 7605 5080 7635
rect 4720 7600 5080 7605
rect 5120 7635 5480 7640
rect 5120 7605 5125 7635
rect 5155 7605 5285 7635
rect 5315 7605 5445 7635
rect 5475 7605 5480 7635
rect 5120 7600 5480 7605
rect 5520 7635 5880 7640
rect 5520 7605 5525 7635
rect 5555 7605 5685 7635
rect 5715 7605 5845 7635
rect 5875 7605 5880 7635
rect 5520 7600 5880 7605
rect 5920 7635 6120 7640
rect 5920 7605 5925 7635
rect 5955 7605 6085 7635
rect 6115 7605 6120 7635
rect 5920 7600 6120 7605
rect 6160 7635 6360 7640
rect 6160 7605 6165 7635
rect 6195 7605 6325 7635
rect 6355 7605 6360 7635
rect 6160 7600 6360 7605
rect 4240 7555 4440 7560
rect 4240 7525 4245 7555
rect 4275 7525 4405 7555
rect 4435 7525 4440 7555
rect 4240 7520 4440 7525
rect 4480 7555 4680 7560
rect 4480 7525 4485 7555
rect 4515 7525 4645 7555
rect 4675 7525 4680 7555
rect 4480 7520 4680 7525
rect 4720 7555 5080 7560
rect 4720 7525 4725 7555
rect 4755 7525 4885 7555
rect 4915 7525 5045 7555
rect 5075 7525 5080 7555
rect 4720 7520 5080 7525
rect 5120 7555 5480 7560
rect 5120 7525 5125 7555
rect 5155 7525 5285 7555
rect 5315 7525 5445 7555
rect 5475 7525 5480 7555
rect 5120 7520 5480 7525
rect 5520 7555 5880 7560
rect 5520 7525 5525 7555
rect 5555 7525 5685 7555
rect 5715 7525 5845 7555
rect 5875 7525 5880 7555
rect 5520 7520 5880 7525
rect 5920 7555 6120 7560
rect 5920 7525 5925 7555
rect 5955 7525 6085 7555
rect 6115 7525 6120 7555
rect 5920 7520 6120 7525
rect 6160 7555 6360 7560
rect 6160 7525 6165 7555
rect 6195 7525 6325 7555
rect 6355 7525 6360 7555
rect 6160 7520 6360 7525
rect 4240 7475 4440 7480
rect 4240 7445 4245 7475
rect 4275 7445 4405 7475
rect 4435 7445 4440 7475
rect 4240 7440 4440 7445
rect 4480 7475 4680 7480
rect 4480 7445 4485 7475
rect 4515 7445 4645 7475
rect 4675 7445 4680 7475
rect 4480 7440 4680 7445
rect 4720 7475 5080 7480
rect 4720 7445 4725 7475
rect 4755 7445 4885 7475
rect 4915 7445 5045 7475
rect 5075 7445 5080 7475
rect 4720 7440 5080 7445
rect 5120 7475 5480 7480
rect 5120 7445 5125 7475
rect 5155 7445 5285 7475
rect 5315 7445 5445 7475
rect 5475 7445 5480 7475
rect 5120 7440 5480 7445
rect 5520 7475 5880 7480
rect 5520 7445 5525 7475
rect 5555 7445 5685 7475
rect 5715 7445 5845 7475
rect 5875 7445 5880 7475
rect 5520 7440 5880 7445
rect 5920 7475 6120 7480
rect 5920 7445 5925 7475
rect 5955 7445 6085 7475
rect 6115 7445 6120 7475
rect 5920 7440 6120 7445
rect 6160 7475 6360 7480
rect 6160 7445 6165 7475
rect 6195 7445 6325 7475
rect 6355 7445 6360 7475
rect 6160 7440 6360 7445
rect 4240 7395 4440 7400
rect 4240 7365 4245 7395
rect 4275 7365 4405 7395
rect 4435 7365 4440 7395
rect 4240 7360 4440 7365
rect 4480 7395 4680 7400
rect 4480 7365 4485 7395
rect 4515 7365 4645 7395
rect 4675 7365 4680 7395
rect 4480 7360 4680 7365
rect 4720 7395 5080 7400
rect 4720 7365 4725 7395
rect 4755 7365 4885 7395
rect 4915 7365 5045 7395
rect 5075 7365 5080 7395
rect 4720 7360 5080 7365
rect 5120 7395 5480 7400
rect 5120 7365 5125 7395
rect 5155 7365 5285 7395
rect 5315 7365 5445 7395
rect 5475 7365 5480 7395
rect 5120 7360 5480 7365
rect 5520 7395 5880 7400
rect 5520 7365 5525 7395
rect 5555 7365 5685 7395
rect 5715 7365 5845 7395
rect 5875 7365 5880 7395
rect 5520 7360 5880 7365
rect 5920 7395 6120 7400
rect 5920 7365 5925 7395
rect 5955 7365 6085 7395
rect 6115 7365 6120 7395
rect 5920 7360 6120 7365
rect 6160 7395 6360 7400
rect 6160 7365 6165 7395
rect 6195 7365 6325 7395
rect 6355 7365 6360 7395
rect 6160 7360 6360 7365
rect 4240 7315 4440 7320
rect 4240 7285 4245 7315
rect 4275 7285 4405 7315
rect 4435 7285 4440 7315
rect 4240 7280 4440 7285
rect 4480 7315 4680 7320
rect 4480 7285 4485 7315
rect 4515 7285 4645 7315
rect 4675 7285 4680 7315
rect 4480 7280 4680 7285
rect 4720 7315 5080 7320
rect 4720 7285 4725 7315
rect 4755 7285 4885 7315
rect 4915 7285 5045 7315
rect 5075 7285 5080 7315
rect 4720 7280 5080 7285
rect 5120 7315 5480 7320
rect 5120 7285 5125 7315
rect 5155 7285 5285 7315
rect 5315 7285 5445 7315
rect 5475 7285 5480 7315
rect 5120 7280 5480 7285
rect 5520 7315 5880 7320
rect 5520 7285 5525 7315
rect 5555 7285 5685 7315
rect 5715 7285 5845 7315
rect 5875 7285 5880 7315
rect 5520 7280 5880 7285
rect 5920 7315 6120 7320
rect 5920 7285 5925 7315
rect 5955 7285 6085 7315
rect 6115 7285 6120 7315
rect 5920 7280 6120 7285
rect 6160 7315 6360 7320
rect 6160 7285 6165 7315
rect 6195 7285 6325 7315
rect 6355 7285 6360 7315
rect 6160 7280 6360 7285
rect 4240 7235 4440 7240
rect 4240 7205 4245 7235
rect 4275 7205 4405 7235
rect 4435 7205 4440 7235
rect 4240 7200 4440 7205
rect 4480 7235 4680 7240
rect 4480 7205 4485 7235
rect 4515 7205 4645 7235
rect 4675 7205 4680 7235
rect 4480 7200 4680 7205
rect 4720 7235 5080 7240
rect 4720 7205 4725 7235
rect 4755 7205 4885 7235
rect 4915 7205 5045 7235
rect 5075 7205 5080 7235
rect 4720 7200 5080 7205
rect 5120 7235 5480 7240
rect 5120 7205 5125 7235
rect 5155 7205 5285 7235
rect 5315 7205 5445 7235
rect 5475 7205 5480 7235
rect 5120 7200 5480 7205
rect 5520 7235 5880 7240
rect 5520 7205 5525 7235
rect 5555 7205 5685 7235
rect 5715 7205 5845 7235
rect 5875 7205 5880 7235
rect 5520 7200 5880 7205
rect 5920 7235 6120 7240
rect 5920 7205 5925 7235
rect 5955 7205 6085 7235
rect 6115 7205 6120 7235
rect 5920 7200 6120 7205
rect 6160 7235 6360 7240
rect 6160 7205 6165 7235
rect 6195 7205 6325 7235
rect 6355 7205 6360 7235
rect 6160 7200 6360 7205
rect 4240 7155 4440 7160
rect 4240 7125 4245 7155
rect 4275 7125 4405 7155
rect 4435 7125 4440 7155
rect 4240 7120 4440 7125
rect 4480 7155 4680 7160
rect 4480 7125 4485 7155
rect 4515 7125 4645 7155
rect 4675 7125 4680 7155
rect 4480 7120 4680 7125
rect 4720 7155 5080 7160
rect 4720 7125 4725 7155
rect 4755 7125 4885 7155
rect 4915 7125 5045 7155
rect 5075 7125 5080 7155
rect 4720 7120 5080 7125
rect 5120 7155 5480 7160
rect 5120 7125 5125 7155
rect 5155 7125 5285 7155
rect 5315 7125 5445 7155
rect 5475 7125 5480 7155
rect 5120 7120 5480 7125
rect 5520 7155 5880 7160
rect 5520 7125 5525 7155
rect 5555 7125 5685 7155
rect 5715 7125 5845 7155
rect 5875 7125 5880 7155
rect 5520 7120 5880 7125
rect 5920 7155 6120 7160
rect 5920 7125 5925 7155
rect 5955 7125 6085 7155
rect 6115 7125 6120 7155
rect 5920 7120 6120 7125
rect 6160 7155 6360 7160
rect 6160 7125 6165 7155
rect 6195 7125 6325 7155
rect 6355 7125 6360 7155
rect 6160 7120 6360 7125
rect 4240 7075 4440 7080
rect 4240 7045 4245 7075
rect 4275 7045 4405 7075
rect 4435 7045 4440 7075
rect 4240 7040 4440 7045
rect 4480 7075 4680 7080
rect 4480 7045 4485 7075
rect 4515 7045 4645 7075
rect 4675 7045 4680 7075
rect 4480 7040 4680 7045
rect 4720 7075 5080 7080
rect 4720 7045 4725 7075
rect 4755 7045 4885 7075
rect 4915 7045 5045 7075
rect 5075 7045 5080 7075
rect 4720 7040 5080 7045
rect 5120 7075 5480 7080
rect 5120 7045 5125 7075
rect 5155 7045 5285 7075
rect 5315 7045 5445 7075
rect 5475 7045 5480 7075
rect 5120 7040 5480 7045
rect 5520 7075 5880 7080
rect 5520 7045 5525 7075
rect 5555 7045 5685 7075
rect 5715 7045 5845 7075
rect 5875 7045 5880 7075
rect 5520 7040 5880 7045
rect 5920 7075 6120 7080
rect 5920 7045 5925 7075
rect 5955 7045 6085 7075
rect 6115 7045 6120 7075
rect 5920 7040 6120 7045
rect 6160 7075 6360 7080
rect 6160 7045 6165 7075
rect 6195 7045 6325 7075
rect 6355 7045 6360 7075
rect 6160 7040 6360 7045
rect 4200 6995 6400 7000
rect 4200 6965 4485 6995
rect 4515 6965 4645 6995
rect 4675 6965 6400 6995
rect 4200 6960 6400 6965
rect 4200 6915 6400 6920
rect 4200 6885 4565 6915
rect 4595 6885 6400 6915
rect 4200 6880 6400 6885
rect 4200 6835 6400 6840
rect 4200 6805 4485 6835
rect 4515 6805 4645 6835
rect 4675 6805 6400 6835
rect 4200 6800 6400 6805
rect 4240 6755 4440 6760
rect 4240 6725 4245 6755
rect 4275 6725 4405 6755
rect 4435 6725 4440 6755
rect 4240 6720 4440 6725
rect 4480 6755 4680 6760
rect 4480 6725 4485 6755
rect 4515 6725 4645 6755
rect 4675 6725 4680 6755
rect 4480 6720 4680 6725
rect 4720 6755 5080 6760
rect 4720 6725 4725 6755
rect 4755 6725 4885 6755
rect 4915 6725 5045 6755
rect 5075 6725 5080 6755
rect 4720 6720 5080 6725
rect 5120 6755 5480 6760
rect 5120 6725 5125 6755
rect 5155 6725 5285 6755
rect 5315 6725 5445 6755
rect 5475 6725 5480 6755
rect 5120 6720 5480 6725
rect 5520 6755 5880 6760
rect 5520 6725 5525 6755
rect 5555 6725 5685 6755
rect 5715 6725 5845 6755
rect 5875 6725 5880 6755
rect 5520 6720 5880 6725
rect 5920 6755 6120 6760
rect 5920 6725 5925 6755
rect 5955 6725 6085 6755
rect 6115 6725 6120 6755
rect 5920 6720 6120 6725
rect 6160 6755 6360 6760
rect 6160 6725 6165 6755
rect 6195 6725 6325 6755
rect 6355 6725 6360 6755
rect 6160 6720 6360 6725
rect 4240 6675 4440 6680
rect 4240 6645 4245 6675
rect 4275 6645 4405 6675
rect 4435 6645 4440 6675
rect 4240 6640 4440 6645
rect 4480 6675 4680 6680
rect 4480 6645 4485 6675
rect 4515 6645 4645 6675
rect 4675 6645 4680 6675
rect 4480 6640 4680 6645
rect 4720 6675 5080 6680
rect 4720 6645 4725 6675
rect 4755 6645 4885 6675
rect 4915 6645 5045 6675
rect 5075 6645 5080 6675
rect 4720 6640 5080 6645
rect 5120 6675 5480 6680
rect 5120 6645 5125 6675
rect 5155 6645 5285 6675
rect 5315 6645 5445 6675
rect 5475 6645 5480 6675
rect 5120 6640 5480 6645
rect 5520 6675 5880 6680
rect 5520 6645 5525 6675
rect 5555 6645 5685 6675
rect 5715 6645 5845 6675
rect 5875 6645 5880 6675
rect 5520 6640 5880 6645
rect 5920 6675 6120 6680
rect 5920 6645 5925 6675
rect 5955 6645 6085 6675
rect 6115 6645 6120 6675
rect 5920 6640 6120 6645
rect 6160 6675 6360 6680
rect 6160 6645 6165 6675
rect 6195 6645 6325 6675
rect 6355 6645 6360 6675
rect 6160 6640 6360 6645
rect 4240 6595 4440 6600
rect 4240 6565 4245 6595
rect 4275 6565 4405 6595
rect 4435 6565 4440 6595
rect 4240 6560 4440 6565
rect 4480 6595 4680 6600
rect 4480 6565 4485 6595
rect 4515 6565 4645 6595
rect 4675 6565 4680 6595
rect 4480 6560 4680 6565
rect 4720 6595 5080 6600
rect 4720 6565 4725 6595
rect 4755 6565 4885 6595
rect 4915 6565 5045 6595
rect 5075 6565 5080 6595
rect 4720 6560 5080 6565
rect 5120 6595 5480 6600
rect 5120 6565 5125 6595
rect 5155 6565 5285 6595
rect 5315 6565 5445 6595
rect 5475 6565 5480 6595
rect 5120 6560 5480 6565
rect 5520 6595 5880 6600
rect 5520 6565 5525 6595
rect 5555 6565 5685 6595
rect 5715 6565 5845 6595
rect 5875 6565 5880 6595
rect 5520 6560 5880 6565
rect 5920 6595 6120 6600
rect 5920 6565 5925 6595
rect 5955 6565 6085 6595
rect 6115 6565 6120 6595
rect 5920 6560 6120 6565
rect 6160 6595 6360 6600
rect 6160 6565 6165 6595
rect 6195 6565 6325 6595
rect 6355 6565 6360 6595
rect 6160 6560 6360 6565
rect 4240 6515 4440 6520
rect 4240 6485 4245 6515
rect 4275 6485 4405 6515
rect 4435 6485 4440 6515
rect 4240 6480 4440 6485
rect 4480 6515 4680 6520
rect 4480 6485 4485 6515
rect 4515 6485 4645 6515
rect 4675 6485 4680 6515
rect 4480 6480 4680 6485
rect 4720 6515 5080 6520
rect 4720 6485 4725 6515
rect 4755 6485 4885 6515
rect 4915 6485 5045 6515
rect 5075 6485 5080 6515
rect 4720 6480 5080 6485
rect 5120 6515 5480 6520
rect 5120 6485 5125 6515
rect 5155 6485 5285 6515
rect 5315 6485 5445 6515
rect 5475 6485 5480 6515
rect 5120 6480 5480 6485
rect 5520 6515 5880 6520
rect 5520 6485 5525 6515
rect 5555 6485 5685 6515
rect 5715 6485 5845 6515
rect 5875 6485 5880 6515
rect 5520 6480 5880 6485
rect 5920 6515 6120 6520
rect 5920 6485 5925 6515
rect 5955 6485 6085 6515
rect 6115 6485 6120 6515
rect 5920 6480 6120 6485
rect 6160 6515 6360 6520
rect 6160 6485 6165 6515
rect 6195 6485 6325 6515
rect 6355 6485 6360 6515
rect 6160 6480 6360 6485
rect 4240 6435 4440 6440
rect 4240 6405 4245 6435
rect 4275 6405 4405 6435
rect 4435 6405 4440 6435
rect 4240 6400 4440 6405
rect 4480 6435 4680 6440
rect 4480 6405 4485 6435
rect 4515 6405 4645 6435
rect 4675 6405 4680 6435
rect 4480 6400 4680 6405
rect 4720 6435 5080 6440
rect 4720 6405 4725 6435
rect 4755 6405 4885 6435
rect 4915 6405 5045 6435
rect 5075 6405 5080 6435
rect 4720 6400 5080 6405
rect 5120 6435 5480 6440
rect 5120 6405 5125 6435
rect 5155 6405 5285 6435
rect 5315 6405 5445 6435
rect 5475 6405 5480 6435
rect 5120 6400 5480 6405
rect 5520 6435 5880 6440
rect 5520 6405 5525 6435
rect 5555 6405 5685 6435
rect 5715 6405 5845 6435
rect 5875 6405 5880 6435
rect 5520 6400 5880 6405
rect 5920 6435 6120 6440
rect 5920 6405 5925 6435
rect 5955 6405 6085 6435
rect 6115 6405 6120 6435
rect 5920 6400 6120 6405
rect 6160 6435 6360 6440
rect 6160 6405 6165 6435
rect 6195 6405 6325 6435
rect 6355 6405 6360 6435
rect 6160 6400 6360 6405
rect 4240 6355 4440 6360
rect 4240 6325 4245 6355
rect 4275 6325 4405 6355
rect 4435 6325 4440 6355
rect 4240 6320 4440 6325
rect 4480 6355 4680 6360
rect 4480 6325 4485 6355
rect 4515 6325 4645 6355
rect 4675 6325 4680 6355
rect 4480 6320 4680 6325
rect 4720 6355 5080 6360
rect 4720 6325 4725 6355
rect 4755 6325 4885 6355
rect 4915 6325 5045 6355
rect 5075 6325 5080 6355
rect 4720 6320 5080 6325
rect 5120 6355 5480 6360
rect 5120 6325 5125 6355
rect 5155 6325 5285 6355
rect 5315 6325 5445 6355
rect 5475 6325 5480 6355
rect 5120 6320 5480 6325
rect 5520 6355 5880 6360
rect 5520 6325 5525 6355
rect 5555 6325 5685 6355
rect 5715 6325 5845 6355
rect 5875 6325 5880 6355
rect 5520 6320 5880 6325
rect 5920 6355 6120 6360
rect 5920 6325 5925 6355
rect 5955 6325 6085 6355
rect 6115 6325 6120 6355
rect 5920 6320 6120 6325
rect 6160 6355 6360 6360
rect 6160 6325 6165 6355
rect 6195 6325 6325 6355
rect 6355 6325 6360 6355
rect 6160 6320 6360 6325
rect 4240 6235 6360 6240
rect 4240 6205 4725 6235
rect 4755 6205 4885 6235
rect 4915 6205 5045 6235
rect 5075 6205 6360 6235
rect 4240 6200 6360 6205
rect 4200 6155 4840 6160
rect 4200 6125 4805 6155
rect 4835 6125 4840 6155
rect 4200 6120 4840 6125
rect 4960 6155 6400 6160
rect 4960 6125 4965 6155
rect 4995 6125 6400 6155
rect 4960 6120 6400 6125
rect 4240 6075 6360 6080
rect 4240 6045 4725 6075
rect 4755 6045 4885 6075
rect 4915 6045 5045 6075
rect 5075 6045 6360 6075
rect 4240 6040 6360 6045
rect 4200 5995 6400 6000
rect 4200 5965 4965 5995
rect 4995 5965 6400 5995
rect 4200 5960 6400 5965
rect 4240 5915 6360 5920
rect 4240 5885 4725 5915
rect 4755 5885 4885 5915
rect 4915 5885 5045 5915
rect 5075 5885 6360 5915
rect 4240 5880 6360 5885
rect 4240 5795 4440 5800
rect 4240 5765 4245 5795
rect 4275 5765 4405 5795
rect 4435 5765 4440 5795
rect 4240 5760 4440 5765
rect 4480 5795 4680 5800
rect 4480 5765 4485 5795
rect 4515 5765 4645 5795
rect 4675 5765 4680 5795
rect 4480 5760 4680 5765
rect 4720 5795 5080 5800
rect 4720 5765 4725 5795
rect 4755 5765 4885 5795
rect 4915 5765 5045 5795
rect 5075 5765 5080 5795
rect 4720 5760 5080 5765
rect 5120 5795 5480 5800
rect 5120 5765 5125 5795
rect 5155 5765 5285 5795
rect 5315 5765 5445 5795
rect 5475 5765 5480 5795
rect 5120 5760 5480 5765
rect 5520 5795 5880 5800
rect 5520 5765 5525 5795
rect 5555 5765 5685 5795
rect 5715 5765 5845 5795
rect 5875 5765 5880 5795
rect 5520 5760 5880 5765
rect 5920 5795 6120 5800
rect 5920 5765 5925 5795
rect 5955 5765 6085 5795
rect 6115 5765 6120 5795
rect 5920 5760 6120 5765
rect 6160 5795 6360 5800
rect 6160 5765 6165 5795
rect 6195 5765 6325 5795
rect 6355 5765 6360 5795
rect 6160 5760 6360 5765
rect 4240 5715 4440 5720
rect 4240 5685 4245 5715
rect 4275 5685 4405 5715
rect 4435 5685 4440 5715
rect 4240 5680 4440 5685
rect 4480 5715 4680 5720
rect 4480 5685 4485 5715
rect 4515 5685 4645 5715
rect 4675 5685 4680 5715
rect 4480 5680 4680 5685
rect 4720 5715 5080 5720
rect 4720 5685 4725 5715
rect 4755 5685 4885 5715
rect 4915 5685 5045 5715
rect 5075 5685 5080 5715
rect 4720 5680 5080 5685
rect 5120 5715 5480 5720
rect 5120 5685 5125 5715
rect 5155 5685 5285 5715
rect 5315 5685 5445 5715
rect 5475 5685 5480 5715
rect 5120 5680 5480 5685
rect 5520 5715 5880 5720
rect 5520 5685 5525 5715
rect 5555 5685 5685 5715
rect 5715 5685 5845 5715
rect 5875 5685 5880 5715
rect 5520 5680 5880 5685
rect 5920 5715 6120 5720
rect 5920 5685 5925 5715
rect 5955 5685 6085 5715
rect 6115 5685 6120 5715
rect 5920 5680 6120 5685
rect 6160 5715 6360 5720
rect 6160 5685 6165 5715
rect 6195 5685 6325 5715
rect 6355 5685 6360 5715
rect 6160 5680 6360 5685
rect 4240 5635 4440 5640
rect 4240 5605 4245 5635
rect 4275 5605 4405 5635
rect 4435 5605 4440 5635
rect 4240 5600 4440 5605
rect 4480 5635 4680 5640
rect 4480 5605 4485 5635
rect 4515 5605 4645 5635
rect 4675 5605 4680 5635
rect 4480 5600 4680 5605
rect 4720 5635 5080 5640
rect 4720 5605 4725 5635
rect 4755 5605 4885 5635
rect 4915 5605 5045 5635
rect 5075 5605 5080 5635
rect 4720 5600 5080 5605
rect 5120 5635 5480 5640
rect 5120 5605 5125 5635
rect 5155 5605 5285 5635
rect 5315 5605 5445 5635
rect 5475 5605 5480 5635
rect 5120 5600 5480 5605
rect 5520 5635 5880 5640
rect 5520 5605 5525 5635
rect 5555 5605 5685 5635
rect 5715 5605 5845 5635
rect 5875 5605 5880 5635
rect 5520 5600 5880 5605
rect 5920 5635 6120 5640
rect 5920 5605 5925 5635
rect 5955 5605 6085 5635
rect 6115 5605 6120 5635
rect 5920 5600 6120 5605
rect 6160 5635 6360 5640
rect 6160 5605 6165 5635
rect 6195 5605 6325 5635
rect 6355 5605 6360 5635
rect 6160 5600 6360 5605
rect 4240 5555 4440 5560
rect 4240 5525 4245 5555
rect 4275 5525 4405 5555
rect 4435 5525 4440 5555
rect 4240 5520 4440 5525
rect 4480 5555 4680 5560
rect 4480 5525 4485 5555
rect 4515 5525 4645 5555
rect 4675 5525 4680 5555
rect 4480 5520 4680 5525
rect 4720 5555 5080 5560
rect 4720 5525 4725 5555
rect 4755 5525 4885 5555
rect 4915 5525 5045 5555
rect 5075 5525 5080 5555
rect 4720 5520 5080 5525
rect 5120 5555 5480 5560
rect 5120 5525 5125 5555
rect 5155 5525 5285 5555
rect 5315 5525 5445 5555
rect 5475 5525 5480 5555
rect 5120 5520 5480 5525
rect 5520 5555 5880 5560
rect 5520 5525 5525 5555
rect 5555 5525 5685 5555
rect 5715 5525 5845 5555
rect 5875 5525 5880 5555
rect 5520 5520 5880 5525
rect 5920 5555 6120 5560
rect 5920 5525 5925 5555
rect 5955 5525 6085 5555
rect 6115 5525 6120 5555
rect 5920 5520 6120 5525
rect 6160 5555 6360 5560
rect 6160 5525 6165 5555
rect 6195 5525 6325 5555
rect 6355 5525 6360 5555
rect 6160 5520 6360 5525
rect 4240 5475 4440 5480
rect 4240 5445 4245 5475
rect 4275 5445 4405 5475
rect 4435 5445 4440 5475
rect 4240 5440 4440 5445
rect 4480 5475 4680 5480
rect 4480 5445 4485 5475
rect 4515 5445 4645 5475
rect 4675 5445 4680 5475
rect 4480 5440 4680 5445
rect 4720 5475 5080 5480
rect 4720 5445 4725 5475
rect 4755 5445 4885 5475
rect 4915 5445 5045 5475
rect 5075 5445 5080 5475
rect 4720 5440 5080 5445
rect 5120 5475 5480 5480
rect 5120 5445 5125 5475
rect 5155 5445 5285 5475
rect 5315 5445 5445 5475
rect 5475 5445 5480 5475
rect 5120 5440 5480 5445
rect 5520 5475 5880 5480
rect 5520 5445 5525 5475
rect 5555 5445 5685 5475
rect 5715 5445 5845 5475
rect 5875 5445 5880 5475
rect 5520 5440 5880 5445
rect 5920 5475 6120 5480
rect 5920 5445 5925 5475
rect 5955 5445 6085 5475
rect 6115 5445 6120 5475
rect 5920 5440 6120 5445
rect 6160 5475 6360 5480
rect 6160 5445 6165 5475
rect 6195 5445 6325 5475
rect 6355 5445 6360 5475
rect 6160 5440 6360 5445
rect 4240 5395 4440 5400
rect 4240 5365 4245 5395
rect 4275 5365 4405 5395
rect 4435 5365 4440 5395
rect 4240 5360 4440 5365
rect 4480 5395 4680 5400
rect 4480 5365 4485 5395
rect 4515 5365 4645 5395
rect 4675 5365 4680 5395
rect 4480 5360 4680 5365
rect 4720 5395 5080 5400
rect 4720 5365 4725 5395
rect 4755 5365 4885 5395
rect 4915 5365 5045 5395
rect 5075 5365 5080 5395
rect 4720 5360 5080 5365
rect 5120 5395 5480 5400
rect 5120 5365 5125 5395
rect 5155 5365 5285 5395
rect 5315 5365 5445 5395
rect 5475 5365 5480 5395
rect 5120 5360 5480 5365
rect 5520 5395 5880 5400
rect 5520 5365 5525 5395
rect 5555 5365 5685 5395
rect 5715 5365 5845 5395
rect 5875 5365 5880 5395
rect 5520 5360 5880 5365
rect 5920 5395 6120 5400
rect 5920 5365 5925 5395
rect 5955 5365 6085 5395
rect 6115 5365 6120 5395
rect 5920 5360 6120 5365
rect 6160 5395 6360 5400
rect 6160 5365 6165 5395
rect 6195 5365 6325 5395
rect 6355 5365 6360 5395
rect 6160 5360 6360 5365
rect 4240 5315 4440 5320
rect 4240 5285 4245 5315
rect 4275 5285 4405 5315
rect 4435 5285 4440 5315
rect 4240 5280 4440 5285
rect 4480 5315 4680 5320
rect 4480 5285 4485 5315
rect 4515 5285 4645 5315
rect 4675 5285 4680 5315
rect 4480 5280 4680 5285
rect 4720 5315 5080 5320
rect 4720 5285 4725 5315
rect 4755 5285 4885 5315
rect 4915 5285 5045 5315
rect 5075 5285 5080 5315
rect 4720 5280 5080 5285
rect 5120 5315 5480 5320
rect 5120 5285 5125 5315
rect 5155 5285 5285 5315
rect 5315 5285 5445 5315
rect 5475 5285 5480 5315
rect 5120 5280 5480 5285
rect 5520 5315 5880 5320
rect 5520 5285 5525 5315
rect 5555 5285 5685 5315
rect 5715 5285 5845 5315
rect 5875 5285 5880 5315
rect 5520 5280 5880 5285
rect 5920 5315 6120 5320
rect 5920 5285 5925 5315
rect 5955 5285 6085 5315
rect 6115 5285 6120 5315
rect 5920 5280 6120 5285
rect 6160 5315 6360 5320
rect 6160 5285 6165 5315
rect 6195 5285 6325 5315
rect 6355 5285 6360 5315
rect 6160 5280 6360 5285
rect 4240 5235 4440 5240
rect 4240 5205 4245 5235
rect 4275 5205 4405 5235
rect 4435 5205 4440 5235
rect 4240 5200 4440 5205
rect 4480 5235 4680 5240
rect 4480 5205 4485 5235
rect 4515 5205 4645 5235
rect 4675 5205 4680 5235
rect 4480 5200 4680 5205
rect 4720 5235 5080 5240
rect 4720 5205 4725 5235
rect 4755 5205 4885 5235
rect 4915 5205 5045 5235
rect 5075 5205 5080 5235
rect 4720 5200 5080 5205
rect 5120 5235 5480 5240
rect 5120 5205 5125 5235
rect 5155 5205 5285 5235
rect 5315 5205 5445 5235
rect 5475 5205 5480 5235
rect 5120 5200 5480 5205
rect 5520 5235 5880 5240
rect 5520 5205 5525 5235
rect 5555 5205 5685 5235
rect 5715 5205 5845 5235
rect 5875 5205 5880 5235
rect 5520 5200 5880 5205
rect 5920 5235 6120 5240
rect 5920 5205 5925 5235
rect 5955 5205 6085 5235
rect 6115 5205 6120 5235
rect 5920 5200 6120 5205
rect 6160 5235 6360 5240
rect 6160 5205 6165 5235
rect 6195 5205 6325 5235
rect 6355 5205 6360 5235
rect 6160 5200 6360 5205
rect 4240 5155 4440 5160
rect 4240 5125 4245 5155
rect 4275 5125 4405 5155
rect 4435 5125 4440 5155
rect 4240 5120 4440 5125
rect 4480 5155 4680 5160
rect 4480 5125 4485 5155
rect 4515 5125 4645 5155
rect 4675 5125 4680 5155
rect 4480 5120 4680 5125
rect 4720 5155 5080 5160
rect 4720 5125 4725 5155
rect 4755 5125 4885 5155
rect 4915 5125 5045 5155
rect 5075 5125 5080 5155
rect 4720 5120 5080 5125
rect 5120 5155 5480 5160
rect 5120 5125 5125 5155
rect 5155 5125 5285 5155
rect 5315 5125 5445 5155
rect 5475 5125 5480 5155
rect 5120 5120 5480 5125
rect 5520 5155 5880 5160
rect 5520 5125 5525 5155
rect 5555 5125 5685 5155
rect 5715 5125 5845 5155
rect 5875 5125 5880 5155
rect 5520 5120 5880 5125
rect 5920 5155 6120 5160
rect 5920 5125 5925 5155
rect 5955 5125 6085 5155
rect 6115 5125 6120 5155
rect 5920 5120 6120 5125
rect 6160 5155 6360 5160
rect 6160 5125 6165 5155
rect 6195 5125 6325 5155
rect 6355 5125 6360 5155
rect 6160 5120 6360 5125
rect 4240 5075 4440 5080
rect 4240 5045 4245 5075
rect 4275 5045 4405 5075
rect 4435 5045 4440 5075
rect 4240 5040 4440 5045
rect 4480 5075 4680 5080
rect 4480 5045 4485 5075
rect 4515 5045 4645 5075
rect 4675 5045 4680 5075
rect 4480 5040 4680 5045
rect 4720 5075 5080 5080
rect 4720 5045 4725 5075
rect 4755 5045 4885 5075
rect 4915 5045 5045 5075
rect 5075 5045 5080 5075
rect 4720 5040 5080 5045
rect 5120 5075 5480 5080
rect 5120 5045 5125 5075
rect 5155 5045 5285 5075
rect 5315 5045 5445 5075
rect 5475 5045 5480 5075
rect 5120 5040 5480 5045
rect 5520 5075 5880 5080
rect 5520 5045 5525 5075
rect 5555 5045 5685 5075
rect 5715 5045 5845 5075
rect 5875 5045 5880 5075
rect 5520 5040 5880 5045
rect 5920 5075 6120 5080
rect 5920 5045 5925 5075
rect 5955 5045 6085 5075
rect 6115 5045 6120 5075
rect 5920 5040 6120 5045
rect 6160 5075 6360 5080
rect 6160 5045 6165 5075
rect 6195 5045 6325 5075
rect 6355 5045 6360 5075
rect 6160 5040 6360 5045
rect 4240 4995 4440 5000
rect 4240 4965 4245 4995
rect 4275 4965 4405 4995
rect 4435 4965 4440 4995
rect 4240 4960 4440 4965
rect 4480 4995 4680 5000
rect 4480 4965 4485 4995
rect 4515 4965 4645 4995
rect 4675 4965 4680 4995
rect 4480 4960 4680 4965
rect 4720 4995 5080 5000
rect 4720 4965 4725 4995
rect 4755 4965 4885 4995
rect 4915 4965 5045 4995
rect 5075 4965 5080 4995
rect 4720 4960 5080 4965
rect 5120 4995 5480 5000
rect 5120 4965 5125 4995
rect 5155 4965 5285 4995
rect 5315 4965 5445 4995
rect 5475 4965 5480 4995
rect 5120 4960 5480 4965
rect 5520 4995 5880 5000
rect 5520 4965 5525 4995
rect 5555 4965 5685 4995
rect 5715 4965 5845 4995
rect 5875 4965 5880 4995
rect 5520 4960 5880 4965
rect 5920 4995 6120 5000
rect 5920 4965 5925 4995
rect 5955 4965 6085 4995
rect 6115 4965 6120 4995
rect 5920 4960 6120 4965
rect 6160 4995 6360 5000
rect 6160 4965 6165 4995
rect 6195 4965 6325 4995
rect 6355 4965 6360 4995
rect 6160 4960 6360 4965
rect 4240 4915 6360 4920
rect 4240 4885 5925 4915
rect 5955 4885 6085 4915
rect 6115 4885 6360 4915
rect 4240 4880 6360 4885
rect 4200 4835 6400 4840
rect 4200 4805 6005 4835
rect 6035 4805 6400 4835
rect 4200 4800 6400 4805
rect 4240 4755 6360 4760
rect 4240 4725 5925 4755
rect 5955 4725 6085 4755
rect 6115 4725 6360 4755
rect 4240 4720 6360 4725
rect 4240 4675 6360 4680
rect 4240 4645 6165 4675
rect 6195 4645 6325 4675
rect 6355 4645 6360 4675
rect 4240 4640 6360 4645
rect 4200 4595 6400 4600
rect 4200 4565 6245 4595
rect 6275 4565 6400 4595
rect 4200 4560 6400 4565
rect 4240 4515 6360 4520
rect 4240 4485 6165 4515
rect 6195 4485 6325 4515
rect 6355 4485 6360 4515
rect 4240 4480 6360 4485
rect 4240 4435 4440 4440
rect 4240 4405 4245 4435
rect 4275 4405 4405 4435
rect 4435 4405 4440 4435
rect 4240 4400 4440 4405
rect 4480 4435 4680 4440
rect 4480 4405 4485 4435
rect 4515 4405 4645 4435
rect 4675 4405 4680 4435
rect 4480 4400 4680 4405
rect 4720 4435 5080 4440
rect 4720 4405 4725 4435
rect 4755 4405 4885 4435
rect 4915 4405 5045 4435
rect 5075 4405 5080 4435
rect 4720 4400 5080 4405
rect 5120 4435 5480 4440
rect 5120 4405 5125 4435
rect 5155 4405 5285 4435
rect 5315 4405 5445 4435
rect 5475 4405 5480 4435
rect 5120 4400 5480 4405
rect 5520 4435 5880 4440
rect 5520 4405 5525 4435
rect 5555 4405 5685 4435
rect 5715 4405 5845 4435
rect 5875 4405 5880 4435
rect 5520 4400 5880 4405
rect 5920 4435 6120 4440
rect 5920 4405 5925 4435
rect 5955 4405 6085 4435
rect 6115 4405 6120 4435
rect 5920 4400 6120 4405
rect 6160 4435 6360 4440
rect 6160 4405 6165 4435
rect 6195 4405 6325 4435
rect 6355 4405 6360 4435
rect 6160 4400 6360 4405
rect 4240 4355 4440 4360
rect 4240 4325 4245 4355
rect 4275 4325 4405 4355
rect 4435 4325 4440 4355
rect 4240 4320 4440 4325
rect 4480 4355 4680 4360
rect 4480 4325 4485 4355
rect 4515 4325 4645 4355
rect 4675 4325 4680 4355
rect 4480 4320 4680 4325
rect 4720 4355 5080 4360
rect 4720 4325 4725 4355
rect 4755 4325 4885 4355
rect 4915 4325 5045 4355
rect 5075 4325 5080 4355
rect 4720 4320 5080 4325
rect 5120 4355 5480 4360
rect 5120 4325 5125 4355
rect 5155 4325 5285 4355
rect 5315 4325 5445 4355
rect 5475 4325 5480 4355
rect 5120 4320 5480 4325
rect 5520 4355 5880 4360
rect 5520 4325 5525 4355
rect 5555 4325 5685 4355
rect 5715 4325 5845 4355
rect 5875 4325 5880 4355
rect 5520 4320 5880 4325
rect 5920 4355 6120 4360
rect 5920 4325 5925 4355
rect 5955 4325 6085 4355
rect 6115 4325 6120 4355
rect 5920 4320 6120 4325
rect 6160 4355 6360 4360
rect 6160 4325 6165 4355
rect 6195 4325 6325 4355
rect 6355 4325 6360 4355
rect 6160 4320 6360 4325
rect 4240 4275 4440 4280
rect 4240 4245 4245 4275
rect 4275 4245 4405 4275
rect 4435 4245 4440 4275
rect 4240 4240 4440 4245
rect 4480 4275 4680 4280
rect 4480 4245 4485 4275
rect 4515 4245 4645 4275
rect 4675 4245 4680 4275
rect 4480 4240 4680 4245
rect 4720 4275 5080 4280
rect 4720 4245 4725 4275
rect 4755 4245 4885 4275
rect 4915 4245 5045 4275
rect 5075 4245 5080 4275
rect 4720 4240 5080 4245
rect 5120 4275 5480 4280
rect 5120 4245 5125 4275
rect 5155 4245 5285 4275
rect 5315 4245 5445 4275
rect 5475 4245 5480 4275
rect 5120 4240 5480 4245
rect 5520 4275 5880 4280
rect 5520 4245 5525 4275
rect 5555 4245 5685 4275
rect 5715 4245 5845 4275
rect 5875 4245 5880 4275
rect 5520 4240 5880 4245
rect 5920 4275 6120 4280
rect 5920 4245 5925 4275
rect 5955 4245 6085 4275
rect 6115 4245 6120 4275
rect 5920 4240 6120 4245
rect 6160 4275 6360 4280
rect 6160 4245 6165 4275
rect 6195 4245 6325 4275
rect 6355 4245 6360 4275
rect 6160 4240 6360 4245
rect 4240 4195 4440 4200
rect 4240 4165 4245 4195
rect 4275 4165 4405 4195
rect 4435 4165 4440 4195
rect 4240 4160 4440 4165
rect 4480 4195 4680 4200
rect 4480 4165 4485 4195
rect 4515 4165 4645 4195
rect 4675 4165 4680 4195
rect 4480 4160 4680 4165
rect 4720 4195 5080 4200
rect 4720 4165 4725 4195
rect 4755 4165 4885 4195
rect 4915 4165 5045 4195
rect 5075 4165 5080 4195
rect 4720 4160 5080 4165
rect 5120 4195 5480 4200
rect 5120 4165 5125 4195
rect 5155 4165 5285 4195
rect 5315 4165 5445 4195
rect 5475 4165 5480 4195
rect 5120 4160 5480 4165
rect 5520 4195 5880 4200
rect 5520 4165 5525 4195
rect 5555 4165 5685 4195
rect 5715 4165 5845 4195
rect 5875 4165 5880 4195
rect 5520 4160 5880 4165
rect 5920 4195 6120 4200
rect 5920 4165 5925 4195
rect 5955 4165 6085 4195
rect 6115 4165 6120 4195
rect 5920 4160 6120 4165
rect 6160 4195 6360 4200
rect 6160 4165 6165 4195
rect 6195 4165 6325 4195
rect 6355 4165 6360 4195
rect 6160 4160 6360 4165
rect 4240 4115 4440 4120
rect 4240 4085 4245 4115
rect 4275 4085 4405 4115
rect 4435 4085 4440 4115
rect 4240 4080 4440 4085
rect 4480 4115 4680 4120
rect 4480 4085 4485 4115
rect 4515 4085 4645 4115
rect 4675 4085 4680 4115
rect 4480 4080 4680 4085
rect 4720 4115 5080 4120
rect 4720 4085 4725 4115
rect 4755 4085 4885 4115
rect 4915 4085 5045 4115
rect 5075 4085 5080 4115
rect 4720 4080 5080 4085
rect 5120 4115 5480 4120
rect 5120 4085 5125 4115
rect 5155 4085 5285 4115
rect 5315 4085 5445 4115
rect 5475 4085 5480 4115
rect 5120 4080 5480 4085
rect 5520 4115 5880 4120
rect 5520 4085 5525 4115
rect 5555 4085 5685 4115
rect 5715 4085 5845 4115
rect 5875 4085 5880 4115
rect 5520 4080 5880 4085
rect 5920 4115 6120 4120
rect 5920 4085 5925 4115
rect 5955 4085 6085 4115
rect 6115 4085 6120 4115
rect 5920 4080 6120 4085
rect 6160 4115 6360 4120
rect 6160 4085 6165 4115
rect 6195 4085 6325 4115
rect 6355 4085 6360 4115
rect 6160 4080 6360 4085
rect 4240 4035 4440 4040
rect 4240 4005 4245 4035
rect 4275 4005 4405 4035
rect 4435 4005 4440 4035
rect 4240 4000 4440 4005
rect 4480 4035 4680 4040
rect 4480 4005 4485 4035
rect 4515 4005 4645 4035
rect 4675 4005 4680 4035
rect 4480 4000 4680 4005
rect 4720 4035 5080 4040
rect 4720 4005 4725 4035
rect 4755 4005 4885 4035
rect 4915 4005 5045 4035
rect 5075 4005 5080 4035
rect 4720 4000 5080 4005
rect 5120 4035 5480 4040
rect 5120 4005 5125 4035
rect 5155 4005 5285 4035
rect 5315 4005 5445 4035
rect 5475 4005 5480 4035
rect 5120 4000 5480 4005
rect 5520 4035 5880 4040
rect 5520 4005 5525 4035
rect 5555 4005 5685 4035
rect 5715 4005 5845 4035
rect 5875 4005 5880 4035
rect 5520 4000 5880 4005
rect 5920 4035 6120 4040
rect 5920 4005 5925 4035
rect 5955 4005 6085 4035
rect 6115 4005 6120 4035
rect 5920 4000 6120 4005
rect 6160 4035 6360 4040
rect 6160 4005 6165 4035
rect 6195 4005 6325 4035
rect 6355 4005 6360 4035
rect 6160 4000 6360 4005
rect 4240 3955 4440 3960
rect 4240 3925 4245 3955
rect 4275 3925 4405 3955
rect 4435 3925 4440 3955
rect 4240 3920 4440 3925
rect 4480 3955 4680 3960
rect 4480 3925 4485 3955
rect 4515 3925 4645 3955
rect 4675 3925 4680 3955
rect 4480 3920 4680 3925
rect 4720 3955 5080 3960
rect 4720 3925 4725 3955
rect 4755 3925 4885 3955
rect 4915 3925 5045 3955
rect 5075 3925 5080 3955
rect 4720 3920 5080 3925
rect 5120 3955 5480 3960
rect 5120 3925 5125 3955
rect 5155 3925 5285 3955
rect 5315 3925 5445 3955
rect 5475 3925 5480 3955
rect 5120 3920 5480 3925
rect 5520 3955 5880 3960
rect 5520 3925 5525 3955
rect 5555 3925 5685 3955
rect 5715 3925 5845 3955
rect 5875 3925 5880 3955
rect 5520 3920 5880 3925
rect 5920 3955 6120 3960
rect 5920 3925 5925 3955
rect 5955 3925 6085 3955
rect 6115 3925 6120 3955
rect 5920 3920 6120 3925
rect 6160 3955 6360 3960
rect 6160 3925 6165 3955
rect 6195 3925 6325 3955
rect 6355 3925 6360 3955
rect 6160 3920 6360 3925
rect 4240 3875 6360 3880
rect 4240 3845 4245 3875
rect 4275 3845 4405 3875
rect 4435 3845 6360 3875
rect 4240 3840 6360 3845
rect 4200 3795 6400 3800
rect 4200 3765 4325 3795
rect 4355 3765 6400 3795
rect 4200 3760 6400 3765
rect 4240 3715 6360 3720
rect 4240 3685 4245 3715
rect 4275 3685 4405 3715
rect 4435 3685 6360 3715
rect 4240 3680 6360 3685
rect 4240 3635 6360 3640
rect 4240 3605 4485 3635
rect 4515 3605 4645 3635
rect 4675 3605 6360 3635
rect 4240 3600 6360 3605
rect 4200 3555 6400 3560
rect 4200 3525 4565 3555
rect 4595 3525 6400 3555
rect 4200 3520 6400 3525
rect 4240 3475 6360 3480
rect 4240 3445 4485 3475
rect 4515 3445 4645 3475
rect 4675 3445 6360 3475
rect 4240 3440 6360 3445
rect 4240 3395 6360 3400
rect 4240 3365 5925 3395
rect 5955 3365 6085 3395
rect 6115 3365 6360 3395
rect 4240 3360 6360 3365
rect 4200 3315 6400 3320
rect 4200 3285 6005 3315
rect 6035 3285 6400 3315
rect 4200 3280 6400 3285
rect 4240 3235 6360 3240
rect 4240 3205 5925 3235
rect 5955 3205 6085 3235
rect 6115 3205 6360 3235
rect 4240 3200 6360 3205
rect 4240 3155 4440 3160
rect 4240 3125 4245 3155
rect 4275 3125 4405 3155
rect 4435 3125 4440 3155
rect 4240 3120 4440 3125
rect 4480 3155 4680 3160
rect 4480 3125 4485 3155
rect 4515 3125 4645 3155
rect 4675 3125 4680 3155
rect 4480 3120 4680 3125
rect 4720 3155 5080 3160
rect 4720 3125 4725 3155
rect 4755 3125 4885 3155
rect 4915 3125 5045 3155
rect 5075 3125 5080 3155
rect 4720 3120 5080 3125
rect 5120 3155 5480 3160
rect 5120 3125 5125 3155
rect 5155 3125 5285 3155
rect 5315 3125 5445 3155
rect 5475 3125 5480 3155
rect 5120 3120 5480 3125
rect 5520 3155 5880 3160
rect 5520 3125 5525 3155
rect 5555 3125 5685 3155
rect 5715 3125 5845 3155
rect 5875 3125 5880 3155
rect 5520 3120 5880 3125
rect 5920 3155 6120 3160
rect 5920 3125 5925 3155
rect 5955 3125 6085 3155
rect 6115 3125 6120 3155
rect 5920 3120 6120 3125
rect 6160 3155 6360 3160
rect 6160 3125 6165 3155
rect 6195 3125 6325 3155
rect 6355 3125 6360 3155
rect 6160 3120 6360 3125
rect 4240 3075 4440 3080
rect 4240 3045 4245 3075
rect 4275 3045 4405 3075
rect 4435 3045 4440 3075
rect 4240 3040 4440 3045
rect 4480 3075 4680 3080
rect 4480 3045 4485 3075
rect 4515 3045 4645 3075
rect 4675 3045 4680 3075
rect 4480 3040 4680 3045
rect 4720 3075 5080 3080
rect 4720 3045 4725 3075
rect 4755 3045 4885 3075
rect 4915 3045 5045 3075
rect 5075 3045 5080 3075
rect 4720 3040 5080 3045
rect 5120 3075 5480 3080
rect 5120 3045 5125 3075
rect 5155 3045 5285 3075
rect 5315 3045 5445 3075
rect 5475 3045 5480 3075
rect 5120 3040 5480 3045
rect 5520 3075 5880 3080
rect 5520 3045 5525 3075
rect 5555 3045 5685 3075
rect 5715 3045 5845 3075
rect 5875 3045 5880 3075
rect 5520 3040 5880 3045
rect 5920 3075 6120 3080
rect 5920 3045 5925 3075
rect 5955 3045 6085 3075
rect 6115 3045 6120 3075
rect 5920 3040 6120 3045
rect 6160 3075 6360 3080
rect 6160 3045 6165 3075
rect 6195 3045 6325 3075
rect 6355 3045 6360 3075
rect 6160 3040 6360 3045
rect 4240 2995 4440 3000
rect 4240 2965 4245 2995
rect 4275 2965 4405 2995
rect 4435 2965 4440 2995
rect 4240 2960 4440 2965
rect 4480 2995 4680 3000
rect 4480 2965 4485 2995
rect 4515 2965 4645 2995
rect 4675 2965 4680 2995
rect 4480 2960 4680 2965
rect 4720 2995 5080 3000
rect 4720 2965 4725 2995
rect 4755 2965 4885 2995
rect 4915 2965 5045 2995
rect 5075 2965 5080 2995
rect 4720 2960 5080 2965
rect 5120 2995 5480 3000
rect 5120 2965 5125 2995
rect 5155 2965 5285 2995
rect 5315 2965 5445 2995
rect 5475 2965 5480 2995
rect 5120 2960 5480 2965
rect 5520 2995 5880 3000
rect 5520 2965 5525 2995
rect 5555 2965 5685 2995
rect 5715 2965 5845 2995
rect 5875 2965 5880 2995
rect 5520 2960 5880 2965
rect 5920 2995 6120 3000
rect 5920 2965 5925 2995
rect 5955 2965 6085 2995
rect 6115 2965 6120 2995
rect 5920 2960 6120 2965
rect 6160 2995 6360 3000
rect 6160 2965 6165 2995
rect 6195 2965 6325 2995
rect 6355 2965 6360 2995
rect 6160 2960 6360 2965
rect 4240 2915 4440 2920
rect 4240 2885 4245 2915
rect 4275 2885 4405 2915
rect 4435 2885 4440 2915
rect 4240 2880 4440 2885
rect 4480 2915 4680 2920
rect 4480 2885 4485 2915
rect 4515 2885 4645 2915
rect 4675 2885 4680 2915
rect 4480 2880 4680 2885
rect 4720 2915 5080 2920
rect 4720 2885 4725 2915
rect 4755 2885 4885 2915
rect 4915 2885 5045 2915
rect 5075 2885 5080 2915
rect 4720 2880 5080 2885
rect 5120 2915 5480 2920
rect 5120 2885 5125 2915
rect 5155 2885 5285 2915
rect 5315 2885 5445 2915
rect 5475 2885 5480 2915
rect 5120 2880 5480 2885
rect 5520 2915 5880 2920
rect 5520 2885 5525 2915
rect 5555 2885 5685 2915
rect 5715 2885 5845 2915
rect 5875 2885 5880 2915
rect 5520 2880 5880 2885
rect 5920 2915 6120 2920
rect 5920 2885 5925 2915
rect 5955 2885 6085 2915
rect 6115 2885 6120 2915
rect 5920 2880 6120 2885
rect 6160 2915 6360 2920
rect 6160 2885 6165 2915
rect 6195 2885 6325 2915
rect 6355 2885 6360 2915
rect 6160 2880 6360 2885
rect 4240 2835 4440 2840
rect 4240 2805 4245 2835
rect 4275 2805 4405 2835
rect 4435 2805 4440 2835
rect 4240 2800 4440 2805
rect 4480 2835 4680 2840
rect 4480 2805 4485 2835
rect 4515 2805 4645 2835
rect 4675 2805 4680 2835
rect 4480 2800 4680 2805
rect 4720 2835 5080 2840
rect 4720 2805 4725 2835
rect 4755 2805 4885 2835
rect 4915 2805 5045 2835
rect 5075 2805 5080 2835
rect 4720 2800 5080 2805
rect 5120 2835 5480 2840
rect 5120 2805 5125 2835
rect 5155 2805 5285 2835
rect 5315 2805 5445 2835
rect 5475 2805 5480 2835
rect 5120 2800 5480 2805
rect 5520 2835 5880 2840
rect 5520 2805 5525 2835
rect 5555 2805 5685 2835
rect 5715 2805 5845 2835
rect 5875 2805 5880 2835
rect 5520 2800 5880 2805
rect 5920 2835 6120 2840
rect 5920 2805 5925 2835
rect 5955 2805 6085 2835
rect 6115 2805 6120 2835
rect 5920 2800 6120 2805
rect 6160 2835 6360 2840
rect 6160 2805 6165 2835
rect 6195 2805 6325 2835
rect 6355 2805 6360 2835
rect 6160 2800 6360 2805
rect 4240 2755 4440 2760
rect 4240 2725 4245 2755
rect 4275 2725 4405 2755
rect 4435 2725 4440 2755
rect 4240 2720 4440 2725
rect 4480 2755 4680 2760
rect 4480 2725 4485 2755
rect 4515 2725 4645 2755
rect 4675 2725 4680 2755
rect 4480 2720 4680 2725
rect 4720 2755 5080 2760
rect 4720 2725 4725 2755
rect 4755 2725 4885 2755
rect 4915 2725 5045 2755
rect 5075 2725 5080 2755
rect 4720 2720 5080 2725
rect 5120 2755 5480 2760
rect 5120 2725 5125 2755
rect 5155 2725 5285 2755
rect 5315 2725 5445 2755
rect 5475 2725 5480 2755
rect 5120 2720 5480 2725
rect 5520 2755 5880 2760
rect 5520 2725 5525 2755
rect 5555 2725 5685 2755
rect 5715 2725 5845 2755
rect 5875 2725 5880 2755
rect 5520 2720 5880 2725
rect 5920 2755 6120 2760
rect 5920 2725 5925 2755
rect 5955 2725 6085 2755
rect 6115 2725 6120 2755
rect 5920 2720 6120 2725
rect 6160 2755 6360 2760
rect 6160 2725 6165 2755
rect 6195 2725 6325 2755
rect 6355 2725 6360 2755
rect 6160 2720 6360 2725
rect 4240 2675 4440 2680
rect 4240 2645 4245 2675
rect 4275 2645 4405 2675
rect 4435 2645 4440 2675
rect 4240 2640 4440 2645
rect 4480 2675 4680 2680
rect 4480 2645 4485 2675
rect 4515 2645 4645 2675
rect 4675 2645 4680 2675
rect 4480 2640 4680 2645
rect 4720 2675 5080 2680
rect 4720 2645 4725 2675
rect 4755 2645 4885 2675
rect 4915 2645 5045 2675
rect 5075 2645 5080 2675
rect 4720 2640 5080 2645
rect 5120 2675 5480 2680
rect 5120 2645 5125 2675
rect 5155 2645 5285 2675
rect 5315 2645 5445 2675
rect 5475 2645 5480 2675
rect 5120 2640 5480 2645
rect 5520 2675 5880 2680
rect 5520 2645 5525 2675
rect 5555 2645 5685 2675
rect 5715 2645 5845 2675
rect 5875 2645 5880 2675
rect 5520 2640 5880 2645
rect 5920 2675 6120 2680
rect 5920 2645 5925 2675
rect 5955 2645 6085 2675
rect 6115 2645 6120 2675
rect 5920 2640 6120 2645
rect 6160 2675 6360 2680
rect 6160 2645 6165 2675
rect 6195 2645 6325 2675
rect 6355 2645 6360 2675
rect 6160 2640 6360 2645
rect 4240 2595 4440 2600
rect 4240 2565 4245 2595
rect 4275 2565 4405 2595
rect 4435 2565 4440 2595
rect 4240 2560 4440 2565
rect 4480 2595 4680 2600
rect 4480 2565 4485 2595
rect 4515 2565 4645 2595
rect 4675 2565 4680 2595
rect 4480 2560 4680 2565
rect 4720 2595 5080 2600
rect 4720 2565 4725 2595
rect 4755 2565 4885 2595
rect 4915 2565 5045 2595
rect 5075 2565 5080 2595
rect 4720 2560 5080 2565
rect 5120 2595 5480 2600
rect 5120 2565 5125 2595
rect 5155 2565 5285 2595
rect 5315 2565 5445 2595
rect 5475 2565 5480 2595
rect 5120 2560 5480 2565
rect 5520 2595 5880 2600
rect 5520 2565 5525 2595
rect 5555 2565 5685 2595
rect 5715 2565 5845 2595
rect 5875 2565 5880 2595
rect 5520 2560 5880 2565
rect 5920 2595 6120 2600
rect 5920 2565 5925 2595
rect 5955 2565 6085 2595
rect 6115 2565 6120 2595
rect 5920 2560 6120 2565
rect 6160 2595 6360 2600
rect 6160 2565 6165 2595
rect 6195 2565 6325 2595
rect 6355 2565 6360 2595
rect 6160 2560 6360 2565
rect 4240 2515 4440 2520
rect 4240 2485 4245 2515
rect 4275 2485 4405 2515
rect 4435 2485 4440 2515
rect 4240 2480 4440 2485
rect 4480 2515 4680 2520
rect 4480 2485 4485 2515
rect 4515 2485 4645 2515
rect 4675 2485 4680 2515
rect 4480 2480 4680 2485
rect 4720 2515 5080 2520
rect 4720 2485 4725 2515
rect 4755 2485 4885 2515
rect 4915 2485 5045 2515
rect 5075 2485 5080 2515
rect 4720 2480 5080 2485
rect 5120 2515 5480 2520
rect 5120 2485 5125 2515
rect 5155 2485 5285 2515
rect 5315 2485 5445 2515
rect 5475 2485 5480 2515
rect 5120 2480 5480 2485
rect 5520 2515 5880 2520
rect 5520 2485 5525 2515
rect 5555 2485 5685 2515
rect 5715 2485 5845 2515
rect 5875 2485 5880 2515
rect 5520 2480 5880 2485
rect 5920 2515 6120 2520
rect 5920 2485 5925 2515
rect 5955 2485 6085 2515
rect 6115 2485 6120 2515
rect 5920 2480 6120 2485
rect 6160 2515 6360 2520
rect 6160 2485 6165 2515
rect 6195 2485 6325 2515
rect 6355 2485 6360 2515
rect 6160 2480 6360 2485
rect 4240 2435 4440 2440
rect 4240 2405 4245 2435
rect 4275 2405 4405 2435
rect 4435 2405 4440 2435
rect 4240 2400 4440 2405
rect 4480 2435 4680 2440
rect 4480 2405 4485 2435
rect 4515 2405 4645 2435
rect 4675 2405 4680 2435
rect 4480 2400 4680 2405
rect 4720 2435 5080 2440
rect 4720 2405 4725 2435
rect 4755 2405 4885 2435
rect 4915 2405 5045 2435
rect 5075 2405 5080 2435
rect 4720 2400 5080 2405
rect 5120 2435 5480 2440
rect 5120 2405 5125 2435
rect 5155 2405 5285 2435
rect 5315 2405 5445 2435
rect 5475 2405 5480 2435
rect 5120 2400 5480 2405
rect 5520 2435 5880 2440
rect 5520 2405 5525 2435
rect 5555 2405 5685 2435
rect 5715 2405 5845 2435
rect 5875 2405 5880 2435
rect 5520 2400 5880 2405
rect 5920 2435 6120 2440
rect 5920 2405 5925 2435
rect 5955 2405 6085 2435
rect 6115 2405 6120 2435
rect 5920 2400 6120 2405
rect 6160 2435 6360 2440
rect 6160 2405 6165 2435
rect 6195 2405 6325 2435
rect 6355 2405 6360 2435
rect 6160 2400 6360 2405
rect 4240 2355 4440 2360
rect 4240 2325 4245 2355
rect 4275 2325 4405 2355
rect 4435 2325 4440 2355
rect 4240 2320 4440 2325
rect 4480 2355 4680 2360
rect 4480 2325 4485 2355
rect 4515 2325 4645 2355
rect 4675 2325 4680 2355
rect 4480 2320 4680 2325
rect 4720 2355 5080 2360
rect 4720 2325 4725 2355
rect 4755 2325 4885 2355
rect 4915 2325 5045 2355
rect 5075 2325 5080 2355
rect 4720 2320 5080 2325
rect 5120 2355 5480 2360
rect 5120 2325 5125 2355
rect 5155 2325 5285 2355
rect 5315 2325 5445 2355
rect 5475 2325 5480 2355
rect 5120 2320 5480 2325
rect 5520 2355 5880 2360
rect 5520 2325 5525 2355
rect 5555 2325 5685 2355
rect 5715 2325 5845 2355
rect 5875 2325 5880 2355
rect 5520 2320 5880 2325
rect 5920 2355 6120 2360
rect 5920 2325 5925 2355
rect 5955 2325 6085 2355
rect 6115 2325 6120 2355
rect 5920 2320 6120 2325
rect 6160 2355 6360 2360
rect 6160 2325 6165 2355
rect 6195 2325 6325 2355
rect 6355 2325 6360 2355
rect 6160 2320 6360 2325
rect 4240 2275 4440 2280
rect 4240 2245 4245 2275
rect 4275 2245 4405 2275
rect 4435 2245 4440 2275
rect 4240 2240 4440 2245
rect 4480 2275 4680 2280
rect 4480 2245 4485 2275
rect 4515 2245 4645 2275
rect 4675 2245 4680 2275
rect 4480 2240 4680 2245
rect 4720 2275 5080 2280
rect 4720 2245 4725 2275
rect 4755 2245 4885 2275
rect 4915 2245 5045 2275
rect 5075 2245 5080 2275
rect 4720 2240 5080 2245
rect 5120 2275 5480 2280
rect 5120 2245 5125 2275
rect 5155 2245 5285 2275
rect 5315 2245 5445 2275
rect 5475 2245 5480 2275
rect 5120 2240 5480 2245
rect 5520 2275 5880 2280
rect 5520 2245 5525 2275
rect 5555 2245 5685 2275
rect 5715 2245 5845 2275
rect 5875 2245 5880 2275
rect 5520 2240 5880 2245
rect 5920 2275 6120 2280
rect 5920 2245 5925 2275
rect 5955 2245 6085 2275
rect 6115 2245 6120 2275
rect 5920 2240 6120 2245
rect 6160 2275 6360 2280
rect 6160 2245 6165 2275
rect 6195 2245 6325 2275
rect 6355 2245 6360 2275
rect 6160 2240 6360 2245
rect 4240 2195 4440 2200
rect 4240 2165 4245 2195
rect 4275 2165 4405 2195
rect 4435 2165 4440 2195
rect 4240 2160 4440 2165
rect 4480 2195 4680 2200
rect 4480 2165 4485 2195
rect 4515 2165 4645 2195
rect 4675 2165 4680 2195
rect 4480 2160 4680 2165
rect 4720 2195 5080 2200
rect 4720 2165 4725 2195
rect 4755 2165 4885 2195
rect 4915 2165 5045 2195
rect 5075 2165 5080 2195
rect 4720 2160 5080 2165
rect 5120 2195 5480 2200
rect 5120 2165 5125 2195
rect 5155 2165 5285 2195
rect 5315 2165 5445 2195
rect 5475 2165 5480 2195
rect 5120 2160 5480 2165
rect 5520 2195 5880 2200
rect 5520 2165 5525 2195
rect 5555 2165 5685 2195
rect 5715 2165 5845 2195
rect 5875 2165 5880 2195
rect 5520 2160 5880 2165
rect 5920 2195 6120 2200
rect 5920 2165 5925 2195
rect 5955 2165 6085 2195
rect 6115 2165 6120 2195
rect 5920 2160 6120 2165
rect 6160 2195 6360 2200
rect 6160 2165 6165 2195
rect 6195 2165 6325 2195
rect 6355 2165 6360 2195
rect 6160 2160 6360 2165
rect 4240 2115 4440 2120
rect 4240 2085 4245 2115
rect 4275 2085 4405 2115
rect 4435 2085 4440 2115
rect 4240 2080 4440 2085
rect 4480 2115 4680 2120
rect 4480 2085 4485 2115
rect 4515 2085 4645 2115
rect 4675 2085 4680 2115
rect 4480 2080 4680 2085
rect 4720 2115 5080 2120
rect 4720 2085 4725 2115
rect 4755 2085 4885 2115
rect 4915 2085 5045 2115
rect 5075 2085 5080 2115
rect 4720 2080 5080 2085
rect 5120 2115 5480 2120
rect 5120 2085 5125 2115
rect 5155 2085 5285 2115
rect 5315 2085 5445 2115
rect 5475 2085 5480 2115
rect 5120 2080 5480 2085
rect 5520 2115 5880 2120
rect 5520 2085 5525 2115
rect 5555 2085 5685 2115
rect 5715 2085 5845 2115
rect 5875 2085 5880 2115
rect 5520 2080 5880 2085
rect 5920 2115 6120 2120
rect 5920 2085 5925 2115
rect 5955 2085 6085 2115
rect 6115 2085 6120 2115
rect 5920 2080 6120 2085
rect 6160 2115 6360 2120
rect 6160 2085 6165 2115
rect 6195 2085 6325 2115
rect 6355 2085 6360 2115
rect 6160 2080 6360 2085
rect 4240 2035 4440 2040
rect 4240 2005 4245 2035
rect 4275 2005 4405 2035
rect 4435 2005 4440 2035
rect 4240 2000 4440 2005
rect 4480 2035 4680 2040
rect 4480 2005 4485 2035
rect 4515 2005 4645 2035
rect 4675 2005 4680 2035
rect 4480 2000 4680 2005
rect 4720 2035 5080 2040
rect 4720 2005 4725 2035
rect 4755 2005 4885 2035
rect 4915 2005 5045 2035
rect 5075 2005 5080 2035
rect 4720 2000 5080 2005
rect 5120 2035 5480 2040
rect 5120 2005 5125 2035
rect 5155 2005 5285 2035
rect 5315 2005 5445 2035
rect 5475 2005 5480 2035
rect 5120 2000 5480 2005
rect 5520 2035 5880 2040
rect 5520 2005 5525 2035
rect 5555 2005 5685 2035
rect 5715 2005 5845 2035
rect 5875 2005 5880 2035
rect 5520 2000 5880 2005
rect 5920 2035 6120 2040
rect 5920 2005 5925 2035
rect 5955 2005 6085 2035
rect 6115 2005 6120 2035
rect 5920 2000 6120 2005
rect 6160 2035 6360 2040
rect 6160 2005 6165 2035
rect 6195 2005 6325 2035
rect 6355 2005 6360 2035
rect 6160 2000 6360 2005
rect 4240 1915 6360 1920
rect 4240 1885 4485 1915
rect 4515 1885 4645 1915
rect 4675 1885 6360 1915
rect 4240 1880 6360 1885
rect 4200 1835 6400 1840
rect 4200 1805 4565 1835
rect 4595 1805 6400 1835
rect 4200 1800 6400 1805
rect 4240 1755 6360 1760
rect 4240 1725 4485 1755
rect 4515 1725 4645 1755
rect 4675 1725 6360 1755
rect 4240 1720 6360 1725
rect 4240 1635 4440 1640
rect 4240 1605 4245 1635
rect 4275 1605 4405 1635
rect 4435 1605 4440 1635
rect 4240 1600 4440 1605
rect 4480 1635 4680 1640
rect 4480 1605 4485 1635
rect 4515 1605 4645 1635
rect 4675 1605 4680 1635
rect 4480 1600 4680 1605
rect 4720 1635 5080 1640
rect 4720 1605 4725 1635
rect 4755 1605 4885 1635
rect 4915 1605 5045 1635
rect 5075 1605 5080 1635
rect 4720 1600 5080 1605
rect 5120 1635 5480 1640
rect 5120 1605 5125 1635
rect 5155 1605 5285 1635
rect 5315 1605 5445 1635
rect 5475 1605 5480 1635
rect 5120 1600 5480 1605
rect 5520 1635 5880 1640
rect 5520 1605 5525 1635
rect 5555 1605 5685 1635
rect 5715 1605 5845 1635
rect 5875 1605 5880 1635
rect 5520 1600 5880 1605
rect 5920 1635 6120 1640
rect 5920 1605 5925 1635
rect 5955 1605 6085 1635
rect 6115 1605 6120 1635
rect 5920 1600 6120 1605
rect 6160 1635 6360 1640
rect 6160 1605 6165 1635
rect 6195 1605 6325 1635
rect 6355 1605 6360 1635
rect 6160 1600 6360 1605
rect 4240 1555 4440 1560
rect 4240 1525 4245 1555
rect 4275 1525 4405 1555
rect 4435 1525 4440 1555
rect 4240 1520 4440 1525
rect 4480 1555 4680 1560
rect 4480 1525 4485 1555
rect 4515 1525 4645 1555
rect 4675 1525 4680 1555
rect 4480 1520 4680 1525
rect 4720 1555 5080 1560
rect 4720 1525 4725 1555
rect 4755 1525 4885 1555
rect 4915 1525 5045 1555
rect 5075 1525 5080 1555
rect 4720 1520 5080 1525
rect 5120 1555 5480 1560
rect 5120 1525 5125 1555
rect 5155 1525 5285 1555
rect 5315 1525 5445 1555
rect 5475 1525 5480 1555
rect 5120 1520 5480 1525
rect 5520 1555 5880 1560
rect 5520 1525 5525 1555
rect 5555 1525 5685 1555
rect 5715 1525 5845 1555
rect 5875 1525 5880 1555
rect 5520 1520 5880 1525
rect 5920 1555 6120 1560
rect 5920 1525 5925 1555
rect 5955 1525 6085 1555
rect 6115 1525 6120 1555
rect 5920 1520 6120 1525
rect 6160 1555 6360 1560
rect 6160 1525 6165 1555
rect 6195 1525 6325 1555
rect 6355 1525 6360 1555
rect 6160 1520 6360 1525
rect 4240 1475 4440 1480
rect 4240 1445 4245 1475
rect 4275 1445 4405 1475
rect 4435 1445 4440 1475
rect 4240 1440 4440 1445
rect 4480 1475 4680 1480
rect 4480 1445 4485 1475
rect 4515 1445 4645 1475
rect 4675 1445 4680 1475
rect 4480 1440 4680 1445
rect 4720 1475 5080 1480
rect 4720 1445 4725 1475
rect 4755 1445 4885 1475
rect 4915 1445 5045 1475
rect 5075 1445 5080 1475
rect 4720 1440 5080 1445
rect 5120 1475 5480 1480
rect 5120 1445 5125 1475
rect 5155 1445 5285 1475
rect 5315 1445 5445 1475
rect 5475 1445 5480 1475
rect 5120 1440 5480 1445
rect 5520 1475 5880 1480
rect 5520 1445 5525 1475
rect 5555 1445 5685 1475
rect 5715 1445 5845 1475
rect 5875 1445 5880 1475
rect 5520 1440 5880 1445
rect 5920 1475 6120 1480
rect 5920 1445 5925 1475
rect 5955 1445 6085 1475
rect 6115 1445 6120 1475
rect 5920 1440 6120 1445
rect 6160 1475 6360 1480
rect 6160 1445 6165 1475
rect 6195 1445 6325 1475
rect 6355 1445 6360 1475
rect 6160 1440 6360 1445
rect 4240 1395 4440 1400
rect 4240 1365 4245 1395
rect 4275 1365 4405 1395
rect 4435 1365 4440 1395
rect 4240 1360 4440 1365
rect 4480 1395 4680 1400
rect 4480 1365 4485 1395
rect 4515 1365 4645 1395
rect 4675 1365 4680 1395
rect 4480 1360 4680 1365
rect 4720 1395 5080 1400
rect 4720 1365 4725 1395
rect 4755 1365 4885 1395
rect 4915 1365 5045 1395
rect 5075 1365 5080 1395
rect 4720 1360 5080 1365
rect 5120 1395 5480 1400
rect 5120 1365 5125 1395
rect 5155 1365 5285 1395
rect 5315 1365 5445 1395
rect 5475 1365 5480 1395
rect 5120 1360 5480 1365
rect 5520 1395 5880 1400
rect 5520 1365 5525 1395
rect 5555 1365 5685 1395
rect 5715 1365 5845 1395
rect 5875 1365 5880 1395
rect 5520 1360 5880 1365
rect 5920 1395 6120 1400
rect 5920 1365 5925 1395
rect 5955 1365 6085 1395
rect 6115 1365 6120 1395
rect 5920 1360 6120 1365
rect 6160 1395 6360 1400
rect 6160 1365 6165 1395
rect 6195 1365 6325 1395
rect 6355 1365 6360 1395
rect 6160 1360 6360 1365
rect 4240 1315 4440 1320
rect 4240 1285 4245 1315
rect 4275 1285 4405 1315
rect 4435 1285 4440 1315
rect 4240 1280 4440 1285
rect 4480 1315 4680 1320
rect 4480 1285 4485 1315
rect 4515 1285 4645 1315
rect 4675 1285 4680 1315
rect 4480 1280 4680 1285
rect 4720 1315 5080 1320
rect 4720 1285 4725 1315
rect 4755 1285 4885 1315
rect 4915 1285 5045 1315
rect 5075 1285 5080 1315
rect 4720 1280 5080 1285
rect 5120 1315 5480 1320
rect 5120 1285 5125 1315
rect 5155 1285 5285 1315
rect 5315 1285 5445 1315
rect 5475 1285 5480 1315
rect 5120 1280 5480 1285
rect 5520 1315 5880 1320
rect 5520 1285 5525 1315
rect 5555 1285 5685 1315
rect 5715 1285 5845 1315
rect 5875 1285 5880 1315
rect 5520 1280 5880 1285
rect 5920 1315 6120 1320
rect 5920 1285 5925 1315
rect 5955 1285 6085 1315
rect 6115 1285 6120 1315
rect 5920 1280 6120 1285
rect 6160 1315 6360 1320
rect 6160 1285 6165 1315
rect 6195 1285 6325 1315
rect 6355 1285 6360 1315
rect 6160 1280 6360 1285
rect 4240 1235 4440 1240
rect 4240 1205 4245 1235
rect 4275 1205 4405 1235
rect 4435 1205 4440 1235
rect 4240 1200 4440 1205
rect 4480 1235 4680 1240
rect 4480 1205 4485 1235
rect 4515 1205 4645 1235
rect 4675 1205 4680 1235
rect 4480 1200 4680 1205
rect 4720 1235 5080 1240
rect 4720 1205 4725 1235
rect 4755 1205 4885 1235
rect 4915 1205 5045 1235
rect 5075 1205 5080 1235
rect 4720 1200 5080 1205
rect 5120 1235 5480 1240
rect 5120 1205 5125 1235
rect 5155 1205 5285 1235
rect 5315 1205 5445 1235
rect 5475 1205 5480 1235
rect 5120 1200 5480 1205
rect 5520 1235 5880 1240
rect 5520 1205 5525 1235
rect 5555 1205 5685 1235
rect 5715 1205 5845 1235
rect 5875 1205 5880 1235
rect 5520 1200 5880 1205
rect 5920 1235 6120 1240
rect 5920 1205 5925 1235
rect 5955 1205 6085 1235
rect 6115 1205 6120 1235
rect 5920 1200 6120 1205
rect 6160 1235 6360 1240
rect 6160 1205 6165 1235
rect 6195 1205 6325 1235
rect 6355 1205 6360 1235
rect 6160 1200 6360 1205
rect 4240 1155 4440 1160
rect 4240 1125 4245 1155
rect 4275 1125 4405 1155
rect 4435 1125 4440 1155
rect 4240 1120 4440 1125
rect 4480 1155 4680 1160
rect 4480 1125 4485 1155
rect 4515 1125 4645 1155
rect 4675 1125 4680 1155
rect 4480 1120 4680 1125
rect 4720 1155 5080 1160
rect 4720 1125 4725 1155
rect 4755 1125 4885 1155
rect 4915 1125 5045 1155
rect 5075 1125 5080 1155
rect 4720 1120 5080 1125
rect 5120 1155 5480 1160
rect 5120 1125 5125 1155
rect 5155 1125 5285 1155
rect 5315 1125 5445 1155
rect 5475 1125 5480 1155
rect 5120 1120 5480 1125
rect 5520 1155 5880 1160
rect 5520 1125 5525 1155
rect 5555 1125 5685 1155
rect 5715 1125 5845 1155
rect 5875 1125 5880 1155
rect 5520 1120 5880 1125
rect 5920 1155 6120 1160
rect 5920 1125 5925 1155
rect 5955 1125 6085 1155
rect 6115 1125 6120 1155
rect 5920 1120 6120 1125
rect 6160 1155 6360 1160
rect 6160 1125 6165 1155
rect 6195 1125 6325 1155
rect 6355 1125 6360 1155
rect 6160 1120 6360 1125
rect 4240 1075 4440 1080
rect 4240 1045 4245 1075
rect 4275 1045 4405 1075
rect 4435 1045 4440 1075
rect 4240 1040 4440 1045
rect 4480 1075 4680 1080
rect 4480 1045 4485 1075
rect 4515 1045 4645 1075
rect 4675 1045 4680 1075
rect 4480 1040 4680 1045
rect 4720 1075 5080 1080
rect 4720 1045 4725 1075
rect 4755 1045 4885 1075
rect 4915 1045 5045 1075
rect 5075 1045 5080 1075
rect 4720 1040 5080 1045
rect 5120 1075 5480 1080
rect 5120 1045 5125 1075
rect 5155 1045 5285 1075
rect 5315 1045 5445 1075
rect 5475 1045 5480 1075
rect 5120 1040 5480 1045
rect 5520 1075 5880 1080
rect 5520 1045 5525 1075
rect 5555 1045 5685 1075
rect 5715 1045 5845 1075
rect 5875 1045 5880 1075
rect 5520 1040 5880 1045
rect 5920 1075 6120 1080
rect 5920 1045 5925 1075
rect 5955 1045 6085 1075
rect 6115 1045 6120 1075
rect 5920 1040 6120 1045
rect 6160 1075 6360 1080
rect 6160 1045 6165 1075
rect 6195 1045 6325 1075
rect 6355 1045 6360 1075
rect 6160 1040 6360 1045
rect 4240 995 6360 1000
rect 4240 965 6165 995
rect 6195 965 6325 995
rect 6355 965 6360 995
rect 4240 960 6360 965
rect 4200 915 6400 920
rect 4200 885 6245 915
rect 6275 885 6400 915
rect 4200 880 6400 885
rect 4240 835 6360 840
rect 4240 805 6165 835
rect 6195 805 6325 835
rect 6355 805 6360 835
rect 4240 800 6360 805
rect 4240 755 4440 760
rect 4240 725 4245 755
rect 4275 725 4405 755
rect 4435 725 4440 755
rect 4240 720 4440 725
rect 4480 755 4680 760
rect 4480 725 4485 755
rect 4515 725 4645 755
rect 4675 725 4680 755
rect 4480 720 4680 725
rect 4720 755 5080 760
rect 4720 725 4725 755
rect 4755 725 4885 755
rect 4915 725 5045 755
rect 5075 725 5080 755
rect 4720 720 5080 725
rect 5120 755 5480 760
rect 5120 725 5125 755
rect 5155 725 5285 755
rect 5315 725 5445 755
rect 5475 725 5480 755
rect 5120 720 5480 725
rect 5520 755 5880 760
rect 5520 725 5525 755
rect 5555 725 5685 755
rect 5715 725 5845 755
rect 5875 725 5880 755
rect 5520 720 5880 725
rect 5920 755 6120 760
rect 5920 725 5925 755
rect 5955 725 6085 755
rect 6115 725 6120 755
rect 5920 720 6120 725
rect 6160 755 6360 760
rect 6160 725 6165 755
rect 6195 725 6325 755
rect 6355 725 6360 755
rect 6160 720 6360 725
rect 4240 675 4440 680
rect 4240 645 4245 675
rect 4275 645 4405 675
rect 4435 645 4440 675
rect 4240 640 4440 645
rect 4480 675 4680 680
rect 4480 645 4485 675
rect 4515 645 4645 675
rect 4675 645 4680 675
rect 4480 640 4680 645
rect 4720 675 5080 680
rect 4720 645 4725 675
rect 4755 645 4885 675
rect 4915 645 5045 675
rect 5075 645 5080 675
rect 4720 640 5080 645
rect 5120 675 5480 680
rect 5120 645 5125 675
rect 5155 645 5285 675
rect 5315 645 5445 675
rect 5475 645 5480 675
rect 5120 640 5480 645
rect 5520 675 5880 680
rect 5520 645 5525 675
rect 5555 645 5685 675
rect 5715 645 5845 675
rect 5875 645 5880 675
rect 5520 640 5880 645
rect 5920 675 6120 680
rect 5920 645 5925 675
rect 5955 645 6085 675
rect 6115 645 6120 675
rect 5920 640 6120 645
rect 6160 675 6360 680
rect 6160 645 6165 675
rect 6195 645 6325 675
rect 6355 645 6360 675
rect 6160 640 6360 645
rect 4240 595 4440 600
rect 4240 565 4245 595
rect 4275 565 4405 595
rect 4435 565 4440 595
rect 4240 560 4440 565
rect 4480 595 4680 600
rect 4480 565 4485 595
rect 4515 565 4645 595
rect 4675 565 4680 595
rect 4480 560 4680 565
rect 4720 595 5080 600
rect 4720 565 4725 595
rect 4755 565 4885 595
rect 4915 565 5045 595
rect 5075 565 5080 595
rect 4720 560 5080 565
rect 5120 595 5480 600
rect 5120 565 5125 595
rect 5155 565 5285 595
rect 5315 565 5445 595
rect 5475 565 5480 595
rect 5120 560 5480 565
rect 5520 595 5880 600
rect 5520 565 5525 595
rect 5555 565 5685 595
rect 5715 565 5845 595
rect 5875 565 5880 595
rect 5520 560 5880 565
rect 5920 595 6120 600
rect 5920 565 5925 595
rect 5955 565 6085 595
rect 6115 565 6120 595
rect 5920 560 6120 565
rect 6160 595 6360 600
rect 6160 565 6165 595
rect 6195 565 6325 595
rect 6355 565 6360 595
rect 6160 560 6360 565
rect 4240 475 6360 480
rect 4240 445 4245 475
rect 4275 445 4405 475
rect 4435 445 6360 475
rect 4240 440 6360 445
rect 4200 395 6400 400
rect 4200 365 4325 395
rect 4355 365 6400 395
rect 4200 360 6400 365
rect 4240 315 6360 320
rect 4240 285 4245 315
rect 4275 285 4405 315
rect 4435 285 6360 315
rect 4240 280 6360 285
rect 4240 195 4440 200
rect 4240 165 4245 195
rect 4275 165 4405 195
rect 4435 165 4440 195
rect 4240 160 4440 165
rect 4480 195 4680 200
rect 4480 165 4485 195
rect 4515 165 4645 195
rect 4675 165 4680 195
rect 4480 160 4680 165
rect 4720 195 5080 200
rect 4720 165 4725 195
rect 4755 165 4885 195
rect 4915 165 5045 195
rect 5075 165 5080 195
rect 4720 160 5080 165
rect 5120 195 5480 200
rect 5120 165 5125 195
rect 5155 165 5285 195
rect 5315 165 5445 195
rect 5475 165 5480 195
rect 5120 160 5480 165
rect 5520 195 5880 200
rect 5520 165 5525 195
rect 5555 165 5685 195
rect 5715 165 5845 195
rect 5875 165 5880 195
rect 5520 160 5880 165
rect 5920 195 6120 200
rect 5920 165 5925 195
rect 5955 165 6085 195
rect 6115 165 6120 195
rect 5920 160 6120 165
rect 6160 195 6360 200
rect 6160 165 6165 195
rect 6195 165 6325 195
rect 6355 165 6360 195
rect 6160 160 6360 165
rect 4240 115 4440 120
rect 4240 85 4245 115
rect 4275 85 4405 115
rect 4435 85 4440 115
rect 4240 80 4440 85
rect 4480 115 4680 120
rect 4480 85 4485 115
rect 4515 85 4645 115
rect 4675 85 4680 115
rect 4480 80 4680 85
rect 4720 115 5080 120
rect 4720 85 4725 115
rect 4755 85 4885 115
rect 4915 85 5045 115
rect 5075 85 5080 115
rect 4720 80 5080 85
rect 5120 115 5480 120
rect 5120 85 5125 115
rect 5155 85 5285 115
rect 5315 85 5445 115
rect 5475 85 5480 115
rect 5120 80 5480 85
rect 5520 115 5880 120
rect 5520 85 5525 115
rect 5555 85 5685 115
rect 5715 85 5845 115
rect 5875 85 5880 115
rect 5520 80 5880 85
rect 5920 115 6120 120
rect 5920 85 5925 115
rect 5955 85 6085 115
rect 6115 85 6120 115
rect 5920 80 6120 85
rect 6160 115 6360 120
rect 6160 85 6165 115
rect 6195 85 6325 115
rect 6355 85 6360 115
rect 6160 80 6360 85
rect 4240 35 4440 40
rect 4240 5 4245 35
rect 4275 5 4405 35
rect 4435 5 4440 35
rect 4240 0 4440 5
rect 4480 35 4680 40
rect 4480 5 4485 35
rect 4515 5 4645 35
rect 4675 5 4680 35
rect 4480 0 4680 5
rect 4720 35 5080 40
rect 4720 5 4725 35
rect 4755 5 4885 35
rect 4915 5 5045 35
rect 5075 5 5080 35
rect 4720 0 5080 5
rect 5120 35 5480 40
rect 5120 5 5125 35
rect 5155 5 5285 35
rect 5315 5 5445 35
rect 5475 5 5480 35
rect 5120 0 5480 5
rect 5520 35 5880 40
rect 5520 5 5525 35
rect 5555 5 5685 35
rect 5715 5 5845 35
rect 5875 5 5880 35
rect 5520 0 5880 5
rect 5920 35 6120 40
rect 5920 5 5925 35
rect 5955 5 6085 35
rect 6115 5 6120 35
rect 5920 0 6120 5
rect 6160 35 6360 40
rect 6160 5 6165 35
rect 6195 5 6325 35
rect 6355 5 6360 35
rect 6160 0 6360 5
<< via2 >>
rect 4245 12605 4275 12635
rect 4405 12605 4435 12635
rect 4485 12605 4515 12635
rect 4645 12605 4675 12635
rect 4725 12605 4755 12635
rect 4885 12605 4915 12635
rect 5045 12605 5075 12635
rect 5125 12605 5155 12635
rect 5285 12605 5315 12635
rect 5445 12605 5475 12635
rect 5525 12605 5555 12635
rect 5685 12605 5715 12635
rect 5845 12605 5875 12635
rect 5925 12605 5955 12635
rect 6085 12605 6115 12635
rect 6165 12605 6195 12635
rect 6325 12605 6355 12635
rect 4245 12525 4275 12555
rect 4405 12525 4435 12555
rect 4485 12525 4515 12555
rect 4645 12525 4675 12555
rect 4725 12525 4755 12555
rect 4885 12525 4915 12555
rect 5045 12525 5075 12555
rect 5125 12525 5155 12555
rect 5285 12525 5315 12555
rect 5445 12525 5475 12555
rect 5525 12525 5555 12555
rect 5685 12525 5715 12555
rect 5845 12525 5875 12555
rect 5925 12525 5955 12555
rect 6085 12525 6115 12555
rect 6165 12525 6195 12555
rect 6325 12525 6355 12555
rect 4245 12445 4275 12475
rect 4405 12445 4435 12475
rect 4485 12445 4515 12475
rect 4645 12445 4675 12475
rect 4725 12445 4755 12475
rect 4885 12445 4915 12475
rect 5045 12445 5075 12475
rect 5125 12445 5155 12475
rect 5285 12445 5315 12475
rect 5445 12445 5475 12475
rect 5525 12445 5555 12475
rect 5685 12445 5715 12475
rect 5845 12445 5875 12475
rect 5925 12445 5955 12475
rect 6085 12445 6115 12475
rect 6165 12445 6195 12475
rect 6325 12445 6355 12475
rect 4245 12365 4275 12395
rect 4405 12365 4435 12395
rect 4485 12365 4515 12395
rect 4645 12365 4675 12395
rect 4725 12365 4755 12395
rect 4885 12365 4915 12395
rect 5045 12365 5075 12395
rect 5125 12365 5155 12395
rect 5285 12365 5315 12395
rect 5445 12365 5475 12395
rect 5525 12365 5555 12395
rect 5685 12365 5715 12395
rect 5845 12365 5875 12395
rect 5925 12365 5955 12395
rect 6085 12365 6115 12395
rect 6165 12365 6195 12395
rect 6325 12365 6355 12395
rect 4245 12285 4275 12315
rect 4405 12285 4435 12315
rect 4485 12285 4515 12315
rect 4645 12285 4675 12315
rect 4725 12285 4755 12315
rect 4885 12285 4915 12315
rect 5045 12285 5075 12315
rect 5125 12285 5155 12315
rect 5285 12285 5315 12315
rect 5445 12285 5475 12315
rect 5525 12285 5555 12315
rect 5685 12285 5715 12315
rect 5845 12285 5875 12315
rect 5925 12285 5955 12315
rect 6085 12285 6115 12315
rect 6165 12285 6195 12315
rect 6325 12285 6355 12315
rect 4245 12205 4275 12235
rect 4405 12205 4435 12235
rect 4485 12205 4515 12235
rect 4645 12205 4675 12235
rect 4725 12205 4755 12235
rect 4885 12205 4915 12235
rect 5045 12205 5075 12235
rect 5125 12205 5155 12235
rect 5285 12205 5315 12235
rect 5445 12205 5475 12235
rect 5525 12205 5555 12235
rect 5685 12205 5715 12235
rect 5845 12205 5875 12235
rect 5925 12205 5955 12235
rect 6085 12205 6115 12235
rect 6165 12205 6195 12235
rect 6325 12205 6355 12235
rect 4245 12125 4275 12155
rect 4405 12125 4435 12155
rect 4485 12125 4515 12155
rect 4645 12125 4675 12155
rect 4725 12125 4755 12155
rect 4885 12125 4915 12155
rect 5045 12125 5075 12155
rect 5125 12125 5155 12155
rect 5285 12125 5315 12155
rect 5445 12125 5475 12155
rect 5525 12125 5555 12155
rect 5685 12125 5715 12155
rect 5845 12125 5875 12155
rect 5925 12125 5955 12155
rect 6085 12125 6115 12155
rect 6165 12125 6195 12155
rect 6325 12125 6355 12155
rect 4485 12045 4515 12075
rect 4645 12045 4675 12075
rect 4565 11965 4595 11995
rect 4485 11885 4515 11915
rect 4645 11885 4675 11915
rect 4245 11805 4275 11835
rect 4405 11805 4435 11835
rect 4485 11805 4515 11835
rect 4645 11805 4675 11835
rect 4725 11805 4755 11835
rect 4885 11805 4915 11835
rect 5045 11805 5075 11835
rect 5125 11805 5155 11835
rect 5285 11805 5315 11835
rect 5445 11805 5475 11835
rect 5525 11805 5555 11835
rect 5685 11805 5715 11835
rect 5845 11805 5875 11835
rect 5925 11805 5955 11835
rect 6085 11805 6115 11835
rect 6165 11805 6195 11835
rect 6325 11805 6355 11835
rect 4245 11725 4275 11755
rect 4405 11725 4435 11755
rect 4485 11725 4515 11755
rect 4645 11725 4675 11755
rect 4725 11725 4755 11755
rect 4885 11725 4915 11755
rect 5045 11725 5075 11755
rect 5125 11725 5155 11755
rect 5285 11725 5315 11755
rect 5445 11725 5475 11755
rect 5525 11725 5555 11755
rect 5685 11725 5715 11755
rect 5845 11725 5875 11755
rect 5925 11725 5955 11755
rect 6085 11725 6115 11755
rect 6165 11725 6195 11755
rect 6325 11725 6355 11755
rect 4245 11645 4275 11675
rect 4405 11645 4435 11675
rect 4485 11645 4515 11675
rect 4645 11645 4675 11675
rect 4725 11645 4755 11675
rect 4885 11645 4915 11675
rect 5045 11645 5075 11675
rect 5125 11645 5155 11675
rect 5285 11645 5315 11675
rect 5445 11645 5475 11675
rect 5525 11645 5555 11675
rect 5685 11645 5715 11675
rect 5845 11645 5875 11675
rect 5925 11645 5955 11675
rect 6085 11645 6115 11675
rect 6165 11645 6195 11675
rect 6325 11645 6355 11675
rect 4245 11565 4275 11595
rect 4405 11565 4435 11595
rect 4485 11565 4515 11595
rect 4645 11565 4675 11595
rect 4725 11565 4755 11595
rect 4885 11565 4915 11595
rect 5045 11565 5075 11595
rect 5125 11565 5155 11595
rect 5285 11565 5315 11595
rect 5445 11565 5475 11595
rect 5525 11565 5555 11595
rect 5685 11565 5715 11595
rect 5845 11565 5875 11595
rect 5925 11565 5955 11595
rect 6085 11565 6115 11595
rect 6165 11565 6195 11595
rect 6325 11565 6355 11595
rect 4245 11485 4275 11515
rect 4405 11485 4435 11515
rect 4485 11485 4515 11515
rect 4645 11485 4675 11515
rect 4725 11485 4755 11515
rect 4885 11485 4915 11515
rect 5045 11485 5075 11515
rect 5125 11485 5155 11515
rect 5285 11485 5315 11515
rect 5445 11485 5475 11515
rect 5525 11485 5555 11515
rect 5685 11485 5715 11515
rect 5845 11485 5875 11515
rect 5925 11485 5955 11515
rect 6085 11485 6115 11515
rect 6165 11485 6195 11515
rect 6325 11485 6355 11515
rect 4245 11405 4275 11435
rect 4405 11405 4435 11435
rect 4485 11405 4515 11435
rect 4645 11405 4675 11435
rect 4725 11405 4755 11435
rect 4885 11405 4915 11435
rect 5045 11405 5075 11435
rect 5125 11405 5155 11435
rect 5285 11405 5315 11435
rect 5445 11405 5475 11435
rect 5525 11405 5555 11435
rect 5685 11405 5715 11435
rect 5845 11405 5875 11435
rect 5925 11405 5955 11435
rect 6085 11405 6115 11435
rect 6165 11405 6195 11435
rect 6325 11405 6355 11435
rect 5525 11285 5555 11315
rect 5685 11285 5715 11315
rect 5605 11205 5635 11235
rect 5045 11125 5075 11155
rect 5525 11125 5555 11155
rect 5685 11125 5715 11155
rect 5125 11045 5155 11075
rect 5285 11045 5315 11075
rect 5445 11045 5475 11075
rect 5045 10965 5075 10995
rect 5525 10965 5555 10995
rect 4245 10845 4275 10875
rect 4405 10845 4435 10875
rect 4485 10845 4515 10875
rect 4645 10845 4675 10875
rect 4725 10845 4755 10875
rect 4885 10845 4915 10875
rect 5045 10845 5075 10875
rect 5125 10845 5155 10875
rect 5285 10845 5315 10875
rect 5445 10845 5475 10875
rect 5525 10845 5555 10875
rect 5685 10845 5715 10875
rect 5845 10845 5875 10875
rect 5925 10845 5955 10875
rect 6085 10845 6115 10875
rect 6165 10845 6195 10875
rect 6325 10845 6355 10875
rect 4245 10765 4275 10795
rect 4405 10765 4435 10795
rect 4485 10765 4515 10795
rect 4645 10765 4675 10795
rect 4725 10765 4755 10795
rect 4885 10765 4915 10795
rect 5045 10765 5075 10795
rect 5125 10765 5155 10795
rect 5285 10765 5315 10795
rect 5445 10765 5475 10795
rect 5525 10765 5555 10795
rect 5685 10765 5715 10795
rect 5845 10765 5875 10795
rect 5925 10765 5955 10795
rect 6085 10765 6115 10795
rect 6165 10765 6195 10795
rect 6325 10765 6355 10795
rect 4245 10685 4275 10715
rect 4405 10685 4435 10715
rect 4485 10685 4515 10715
rect 4645 10685 4675 10715
rect 4725 10685 4755 10715
rect 4885 10685 4915 10715
rect 5045 10685 5075 10715
rect 5125 10685 5155 10715
rect 5285 10685 5315 10715
rect 5445 10685 5475 10715
rect 5525 10685 5555 10715
rect 5685 10685 5715 10715
rect 5845 10685 5875 10715
rect 5925 10685 5955 10715
rect 6085 10685 6115 10715
rect 6165 10685 6195 10715
rect 6325 10685 6355 10715
rect 4245 10605 4275 10635
rect 4405 10605 4435 10635
rect 4485 10605 4515 10635
rect 4645 10605 4675 10635
rect 4725 10605 4755 10635
rect 4885 10605 4915 10635
rect 5045 10605 5075 10635
rect 5125 10605 5155 10635
rect 5285 10605 5315 10635
rect 5445 10605 5475 10635
rect 5525 10605 5555 10635
rect 5685 10605 5715 10635
rect 5845 10605 5875 10635
rect 5925 10605 5955 10635
rect 6085 10605 6115 10635
rect 6165 10605 6195 10635
rect 6325 10605 6355 10635
rect 4245 10525 4275 10555
rect 4405 10525 4435 10555
rect 4485 10525 4515 10555
rect 4645 10525 4675 10555
rect 4725 10525 4755 10555
rect 4885 10525 4915 10555
rect 5045 10525 5075 10555
rect 5125 10525 5155 10555
rect 5285 10525 5315 10555
rect 5445 10525 5475 10555
rect 5525 10525 5555 10555
rect 5685 10525 5715 10555
rect 5845 10525 5875 10555
rect 5925 10525 5955 10555
rect 6085 10525 6115 10555
rect 6165 10525 6195 10555
rect 6325 10525 6355 10555
rect 4245 10445 4275 10475
rect 4405 10445 4435 10475
rect 4485 10445 4515 10475
rect 4645 10445 4675 10475
rect 4725 10445 4755 10475
rect 4885 10445 4915 10475
rect 5045 10445 5075 10475
rect 5125 10445 5155 10475
rect 5285 10445 5315 10475
rect 5445 10445 5475 10475
rect 5525 10445 5555 10475
rect 5685 10445 5715 10475
rect 5845 10445 5875 10475
rect 5925 10445 5955 10475
rect 6085 10445 6115 10475
rect 6165 10445 6195 10475
rect 6325 10445 6355 10475
rect 4245 10365 4275 10395
rect 4405 10365 4435 10395
rect 4485 10365 4515 10395
rect 4645 10365 4675 10395
rect 4725 10365 4755 10395
rect 4885 10365 4915 10395
rect 5045 10365 5075 10395
rect 5125 10365 5155 10395
rect 5285 10365 5315 10395
rect 5445 10365 5475 10395
rect 5525 10365 5555 10395
rect 5685 10365 5715 10395
rect 5845 10365 5875 10395
rect 5925 10365 5955 10395
rect 6085 10365 6115 10395
rect 6165 10365 6195 10395
rect 6325 10365 6355 10395
rect 4245 10285 4275 10315
rect 4405 10285 4435 10315
rect 4485 10285 4515 10315
rect 4645 10285 4675 10315
rect 4725 10285 4755 10315
rect 4885 10285 4915 10315
rect 5045 10285 5075 10315
rect 5125 10285 5155 10315
rect 5285 10285 5315 10315
rect 5445 10285 5475 10315
rect 5525 10285 5555 10315
rect 5685 10285 5715 10315
rect 5845 10285 5875 10315
rect 5925 10285 5955 10315
rect 6085 10285 6115 10315
rect 6165 10285 6195 10315
rect 6325 10285 6355 10315
rect 4245 10205 4275 10235
rect 4405 10205 4435 10235
rect 4485 10205 4515 10235
rect 4645 10205 4675 10235
rect 4725 10205 4755 10235
rect 4885 10205 4915 10235
rect 5045 10205 5075 10235
rect 5125 10205 5155 10235
rect 5285 10205 5315 10235
rect 5445 10205 5475 10235
rect 5525 10205 5555 10235
rect 5685 10205 5715 10235
rect 5845 10205 5875 10235
rect 5925 10205 5955 10235
rect 6085 10205 6115 10235
rect 6165 10205 6195 10235
rect 6325 10205 6355 10235
rect 4245 10125 4275 10155
rect 4405 10125 4435 10155
rect 4485 10125 4515 10155
rect 4645 10125 4675 10155
rect 4725 10125 4755 10155
rect 4885 10125 4915 10155
rect 5045 10125 5075 10155
rect 5125 10125 5155 10155
rect 5285 10125 5315 10155
rect 5445 10125 5475 10155
rect 5525 10125 5555 10155
rect 5685 10125 5715 10155
rect 5845 10125 5875 10155
rect 5925 10125 5955 10155
rect 6085 10125 6115 10155
rect 6165 10125 6195 10155
rect 6325 10125 6355 10155
rect 4245 10045 4275 10075
rect 4405 10045 4435 10075
rect 4485 10045 4515 10075
rect 4645 10045 4675 10075
rect 4725 10045 4755 10075
rect 4885 10045 4915 10075
rect 5045 10045 5075 10075
rect 5125 10045 5155 10075
rect 5285 10045 5315 10075
rect 5445 10045 5475 10075
rect 5525 10045 5555 10075
rect 5685 10045 5715 10075
rect 5845 10045 5875 10075
rect 5925 10045 5955 10075
rect 6085 10045 6115 10075
rect 6165 10045 6195 10075
rect 6325 10045 6355 10075
rect 4245 9965 4275 9995
rect 4405 9965 4435 9995
rect 4485 9965 4515 9995
rect 4645 9965 4675 9995
rect 4725 9965 4755 9995
rect 4885 9965 4915 9995
rect 5045 9965 5075 9995
rect 5125 9965 5155 9995
rect 5285 9965 5315 9995
rect 5445 9965 5475 9995
rect 5525 9965 5555 9995
rect 5685 9965 5715 9995
rect 5845 9965 5875 9995
rect 5925 9965 5955 9995
rect 6085 9965 6115 9995
rect 6165 9965 6195 9995
rect 6325 9965 6355 9995
rect 4245 9885 4275 9915
rect 4405 9885 4435 9915
rect 4485 9885 4515 9915
rect 4645 9885 4675 9915
rect 4725 9885 4755 9915
rect 4885 9885 4915 9915
rect 5045 9885 5075 9915
rect 5125 9885 5155 9915
rect 5285 9885 5315 9915
rect 5445 9885 5475 9915
rect 5525 9885 5555 9915
rect 5685 9885 5715 9915
rect 5845 9885 5875 9915
rect 5925 9885 5955 9915
rect 6085 9885 6115 9915
rect 6165 9885 6195 9915
rect 6325 9885 6355 9915
rect 4245 9805 4275 9835
rect 4405 9805 4435 9835
rect 4485 9805 4515 9835
rect 4645 9805 4675 9835
rect 4725 9805 4755 9835
rect 4885 9805 4915 9835
rect 5045 9805 5075 9835
rect 5125 9805 5155 9835
rect 5285 9805 5315 9835
rect 5445 9805 5475 9835
rect 5525 9805 5555 9835
rect 5685 9805 5715 9835
rect 5845 9805 5875 9835
rect 5925 9805 5955 9835
rect 6085 9805 6115 9835
rect 6165 9805 6195 9835
rect 6325 9805 6355 9835
rect 4245 9725 4275 9755
rect 4405 9725 4435 9755
rect 4485 9725 4515 9755
rect 4645 9725 4675 9755
rect 4725 9725 4755 9755
rect 4885 9725 4915 9755
rect 5045 9725 5075 9755
rect 5125 9725 5155 9755
rect 5285 9725 5315 9755
rect 5445 9725 5475 9755
rect 5525 9725 5555 9755
rect 5685 9725 5715 9755
rect 5845 9725 5875 9755
rect 5925 9725 5955 9755
rect 6085 9725 6115 9755
rect 6165 9725 6195 9755
rect 6325 9725 6355 9755
rect 4485 9605 4515 9635
rect 4645 9605 4675 9635
rect 4565 9525 4595 9555
rect 4485 9445 4515 9475
rect 4645 9445 4675 9475
rect 4245 9325 4275 9355
rect 4405 9325 4435 9355
rect 4485 9325 4515 9355
rect 4645 9325 4675 9355
rect 4725 9325 4755 9355
rect 4885 9325 4915 9355
rect 5045 9325 5075 9355
rect 5125 9325 5155 9355
rect 5285 9325 5315 9355
rect 5445 9325 5475 9355
rect 5525 9325 5555 9355
rect 5685 9325 5715 9355
rect 5845 9325 5875 9355
rect 5925 9325 5955 9355
rect 6085 9325 6115 9355
rect 6165 9325 6195 9355
rect 6325 9325 6355 9355
rect 4245 9245 4275 9275
rect 4405 9245 4435 9275
rect 4485 9245 4515 9275
rect 4645 9245 4675 9275
rect 4725 9245 4755 9275
rect 4885 9245 4915 9275
rect 5045 9245 5075 9275
rect 5125 9245 5155 9275
rect 5285 9245 5315 9275
rect 5445 9245 5475 9275
rect 5525 9245 5555 9275
rect 5685 9245 5715 9275
rect 5845 9245 5875 9275
rect 5925 9245 5955 9275
rect 6085 9245 6115 9275
rect 6165 9245 6195 9275
rect 6325 9245 6355 9275
rect 4245 9165 4275 9195
rect 4405 9165 4435 9195
rect 4485 9165 4515 9195
rect 4645 9165 4675 9195
rect 4725 9165 4755 9195
rect 4885 9165 4915 9195
rect 5045 9165 5075 9195
rect 5125 9165 5155 9195
rect 5285 9165 5315 9195
rect 5445 9165 5475 9195
rect 5525 9165 5555 9195
rect 5685 9165 5715 9195
rect 5845 9165 5875 9195
rect 5925 9165 5955 9195
rect 6085 9165 6115 9195
rect 6165 9165 6195 9195
rect 6325 9165 6355 9195
rect 5125 9085 5155 9115
rect 5285 9085 5315 9115
rect 5445 9085 5475 9115
rect 5365 9005 5395 9035
rect 5125 8925 5155 8955
rect 5285 8925 5315 8955
rect 5445 8925 5475 8955
rect 4245 8845 4275 8875
rect 4405 8845 4435 8875
rect 4485 8845 4515 8875
rect 4645 8845 4675 8875
rect 4725 8845 4755 8875
rect 4885 8845 4915 8875
rect 5045 8845 5075 8875
rect 5125 8845 5155 8875
rect 5285 8845 5315 8875
rect 5445 8845 5475 8875
rect 5525 8845 5555 8875
rect 5685 8845 5715 8875
rect 5845 8845 5875 8875
rect 5925 8845 5955 8875
rect 6085 8845 6115 8875
rect 6165 8845 6195 8875
rect 6325 8845 6355 8875
rect 4245 8765 4275 8795
rect 4405 8765 4435 8795
rect 4485 8765 4515 8795
rect 4645 8765 4675 8795
rect 4725 8765 4755 8795
rect 4885 8765 4915 8795
rect 5045 8765 5075 8795
rect 5125 8765 5155 8795
rect 5285 8765 5315 8795
rect 5445 8765 5475 8795
rect 5525 8765 5555 8795
rect 5685 8765 5715 8795
rect 5845 8765 5875 8795
rect 5925 8765 5955 8795
rect 6085 8765 6115 8795
rect 6165 8765 6195 8795
rect 6325 8765 6355 8795
rect 4245 8685 4275 8715
rect 4405 8685 4435 8715
rect 4485 8685 4515 8715
rect 4645 8685 4675 8715
rect 4725 8685 4755 8715
rect 4885 8685 4915 8715
rect 5045 8685 5075 8715
rect 5125 8685 5155 8715
rect 5285 8685 5315 8715
rect 5445 8685 5475 8715
rect 5525 8685 5555 8715
rect 5685 8685 5715 8715
rect 5845 8685 5875 8715
rect 5925 8685 5955 8715
rect 6085 8685 6115 8715
rect 6165 8685 6195 8715
rect 6325 8685 6355 8715
rect 4245 8605 4275 8635
rect 4405 8605 4435 8635
rect 4485 8605 4515 8635
rect 4645 8605 4675 8635
rect 4725 8605 4755 8635
rect 4885 8605 4915 8635
rect 5045 8605 5075 8635
rect 5125 8605 5155 8635
rect 5285 8605 5315 8635
rect 5445 8605 5475 8635
rect 5525 8605 5555 8635
rect 5685 8605 5715 8635
rect 5845 8605 5875 8635
rect 5925 8605 5955 8635
rect 6085 8605 6115 8635
rect 6165 8605 6195 8635
rect 6325 8605 6355 8635
rect 4245 8525 4275 8555
rect 4405 8525 4435 8555
rect 4485 8525 4515 8555
rect 4645 8525 4675 8555
rect 4725 8525 4755 8555
rect 4885 8525 4915 8555
rect 5045 8525 5075 8555
rect 5125 8525 5155 8555
rect 5285 8525 5315 8555
rect 5445 8525 5475 8555
rect 5525 8525 5555 8555
rect 5685 8525 5715 8555
rect 5845 8525 5875 8555
rect 5925 8525 5955 8555
rect 6085 8525 6115 8555
rect 6165 8525 6195 8555
rect 6325 8525 6355 8555
rect 4885 8445 4915 8475
rect 5045 8445 5075 8475
rect 5685 8445 5715 8475
rect 5845 8445 5875 8475
rect 4965 8365 4995 8395
rect 5765 8365 5795 8395
rect 4885 8285 4915 8315
rect 5045 8285 5075 8315
rect 5525 8285 5555 8315
rect 5685 8285 5715 8315
rect 5845 8285 5875 8315
rect 5605 8205 5635 8235
rect 5525 8125 5555 8155
rect 5685 8125 5715 8155
rect 5045 8045 5075 8075
rect 5525 8045 5555 8075
rect 5125 7965 5155 7995
rect 5285 7965 5315 7995
rect 5445 7965 5475 7995
rect 5205 7885 5235 7915
rect 5125 7805 5155 7835
rect 5285 7805 5315 7835
rect 5445 7805 5475 7835
rect 5045 7725 5075 7755
rect 5525 7725 5555 7755
rect 4245 7605 4275 7635
rect 4405 7605 4435 7635
rect 4485 7605 4515 7635
rect 4645 7605 4675 7635
rect 4725 7605 4755 7635
rect 4885 7605 4915 7635
rect 5045 7605 5075 7635
rect 5125 7605 5155 7635
rect 5285 7605 5315 7635
rect 5445 7605 5475 7635
rect 5525 7605 5555 7635
rect 5685 7605 5715 7635
rect 5845 7605 5875 7635
rect 5925 7605 5955 7635
rect 6085 7605 6115 7635
rect 6165 7605 6195 7635
rect 6325 7605 6355 7635
rect 4245 7525 4275 7555
rect 4405 7525 4435 7555
rect 4485 7525 4515 7555
rect 4645 7525 4675 7555
rect 4725 7525 4755 7555
rect 4885 7525 4915 7555
rect 5045 7525 5075 7555
rect 5125 7525 5155 7555
rect 5285 7525 5315 7555
rect 5445 7525 5475 7555
rect 5525 7525 5555 7555
rect 5685 7525 5715 7555
rect 5845 7525 5875 7555
rect 5925 7525 5955 7555
rect 6085 7525 6115 7555
rect 6165 7525 6195 7555
rect 6325 7525 6355 7555
rect 4245 7445 4275 7475
rect 4405 7445 4435 7475
rect 4485 7445 4515 7475
rect 4645 7445 4675 7475
rect 4725 7445 4755 7475
rect 4885 7445 4915 7475
rect 5045 7445 5075 7475
rect 5125 7445 5155 7475
rect 5285 7445 5315 7475
rect 5445 7445 5475 7475
rect 5525 7445 5555 7475
rect 5685 7445 5715 7475
rect 5845 7445 5875 7475
rect 5925 7445 5955 7475
rect 6085 7445 6115 7475
rect 6165 7445 6195 7475
rect 6325 7445 6355 7475
rect 4245 7365 4275 7395
rect 4405 7365 4435 7395
rect 4485 7365 4515 7395
rect 4645 7365 4675 7395
rect 4725 7365 4755 7395
rect 4885 7365 4915 7395
rect 5045 7365 5075 7395
rect 5125 7365 5155 7395
rect 5285 7365 5315 7395
rect 5445 7365 5475 7395
rect 5525 7365 5555 7395
rect 5685 7365 5715 7395
rect 5845 7365 5875 7395
rect 5925 7365 5955 7395
rect 6085 7365 6115 7395
rect 6165 7365 6195 7395
rect 6325 7365 6355 7395
rect 4245 7285 4275 7315
rect 4405 7285 4435 7315
rect 4485 7285 4515 7315
rect 4645 7285 4675 7315
rect 4725 7285 4755 7315
rect 4885 7285 4915 7315
rect 5045 7285 5075 7315
rect 5125 7285 5155 7315
rect 5285 7285 5315 7315
rect 5445 7285 5475 7315
rect 5525 7285 5555 7315
rect 5685 7285 5715 7315
rect 5845 7285 5875 7315
rect 5925 7285 5955 7315
rect 6085 7285 6115 7315
rect 6165 7285 6195 7315
rect 6325 7285 6355 7315
rect 4245 7205 4275 7235
rect 4405 7205 4435 7235
rect 4485 7205 4515 7235
rect 4645 7205 4675 7235
rect 4725 7205 4755 7235
rect 4885 7205 4915 7235
rect 5045 7205 5075 7235
rect 5125 7205 5155 7235
rect 5285 7205 5315 7235
rect 5445 7205 5475 7235
rect 5525 7205 5555 7235
rect 5685 7205 5715 7235
rect 5845 7205 5875 7235
rect 5925 7205 5955 7235
rect 6085 7205 6115 7235
rect 6165 7205 6195 7235
rect 6325 7205 6355 7235
rect 4245 7125 4275 7155
rect 4405 7125 4435 7155
rect 4485 7125 4515 7155
rect 4645 7125 4675 7155
rect 4725 7125 4755 7155
rect 4885 7125 4915 7155
rect 5045 7125 5075 7155
rect 5125 7125 5155 7155
rect 5285 7125 5315 7155
rect 5445 7125 5475 7155
rect 5525 7125 5555 7155
rect 5685 7125 5715 7155
rect 5845 7125 5875 7155
rect 5925 7125 5955 7155
rect 6085 7125 6115 7155
rect 6165 7125 6195 7155
rect 6325 7125 6355 7155
rect 4245 7045 4275 7075
rect 4405 7045 4435 7075
rect 4485 7045 4515 7075
rect 4645 7045 4675 7075
rect 4725 7045 4755 7075
rect 4885 7045 4915 7075
rect 5045 7045 5075 7075
rect 5125 7045 5155 7075
rect 5285 7045 5315 7075
rect 5445 7045 5475 7075
rect 5525 7045 5555 7075
rect 5685 7045 5715 7075
rect 5845 7045 5875 7075
rect 5925 7045 5955 7075
rect 6085 7045 6115 7075
rect 6165 7045 6195 7075
rect 6325 7045 6355 7075
rect 4485 6965 4515 6995
rect 4645 6965 4675 6995
rect 4565 6885 4595 6915
rect 4485 6805 4515 6835
rect 4645 6805 4675 6835
rect 4245 6725 4275 6755
rect 4405 6725 4435 6755
rect 4485 6725 4515 6755
rect 4645 6725 4675 6755
rect 4725 6725 4755 6755
rect 4885 6725 4915 6755
rect 5045 6725 5075 6755
rect 5125 6725 5155 6755
rect 5285 6725 5315 6755
rect 5445 6725 5475 6755
rect 5525 6725 5555 6755
rect 5685 6725 5715 6755
rect 5845 6725 5875 6755
rect 5925 6725 5955 6755
rect 6085 6725 6115 6755
rect 6165 6725 6195 6755
rect 6325 6725 6355 6755
rect 4245 6645 4275 6675
rect 4405 6645 4435 6675
rect 4485 6645 4515 6675
rect 4645 6645 4675 6675
rect 4725 6645 4755 6675
rect 4885 6645 4915 6675
rect 5045 6645 5075 6675
rect 5125 6645 5155 6675
rect 5285 6645 5315 6675
rect 5445 6645 5475 6675
rect 5525 6645 5555 6675
rect 5685 6645 5715 6675
rect 5845 6645 5875 6675
rect 5925 6645 5955 6675
rect 6085 6645 6115 6675
rect 6165 6645 6195 6675
rect 6325 6645 6355 6675
rect 4245 6565 4275 6595
rect 4405 6565 4435 6595
rect 4485 6565 4515 6595
rect 4645 6565 4675 6595
rect 4725 6565 4755 6595
rect 4885 6565 4915 6595
rect 5045 6565 5075 6595
rect 5125 6565 5155 6595
rect 5285 6565 5315 6595
rect 5445 6565 5475 6595
rect 5525 6565 5555 6595
rect 5685 6565 5715 6595
rect 5845 6565 5875 6595
rect 5925 6565 5955 6595
rect 6085 6565 6115 6595
rect 6165 6565 6195 6595
rect 6325 6565 6355 6595
rect 4245 6485 4275 6515
rect 4405 6485 4435 6515
rect 4485 6485 4515 6515
rect 4645 6485 4675 6515
rect 4725 6485 4755 6515
rect 4885 6485 4915 6515
rect 5045 6485 5075 6515
rect 5125 6485 5155 6515
rect 5285 6485 5315 6515
rect 5445 6485 5475 6515
rect 5525 6485 5555 6515
rect 5685 6485 5715 6515
rect 5845 6485 5875 6515
rect 5925 6485 5955 6515
rect 6085 6485 6115 6515
rect 6165 6485 6195 6515
rect 6325 6485 6355 6515
rect 4245 6405 4275 6435
rect 4405 6405 4435 6435
rect 4485 6405 4515 6435
rect 4645 6405 4675 6435
rect 4725 6405 4755 6435
rect 4885 6405 4915 6435
rect 5045 6405 5075 6435
rect 5125 6405 5155 6435
rect 5285 6405 5315 6435
rect 5445 6405 5475 6435
rect 5525 6405 5555 6435
rect 5685 6405 5715 6435
rect 5845 6405 5875 6435
rect 5925 6405 5955 6435
rect 6085 6405 6115 6435
rect 6165 6405 6195 6435
rect 6325 6405 6355 6435
rect 4245 6325 4275 6355
rect 4405 6325 4435 6355
rect 4485 6325 4515 6355
rect 4645 6325 4675 6355
rect 4725 6325 4755 6355
rect 4885 6325 4915 6355
rect 5045 6325 5075 6355
rect 5125 6325 5155 6355
rect 5285 6325 5315 6355
rect 5445 6325 5475 6355
rect 5525 6325 5555 6355
rect 5685 6325 5715 6355
rect 5845 6325 5875 6355
rect 5925 6325 5955 6355
rect 6085 6325 6115 6355
rect 6165 6325 6195 6355
rect 6325 6325 6355 6355
rect 4725 6205 4755 6235
rect 4885 6205 4915 6235
rect 5045 6205 5075 6235
rect 4805 6125 4835 6155
rect 4965 6125 4995 6155
rect 4725 6045 4755 6075
rect 4885 6045 4915 6075
rect 5045 6045 5075 6075
rect 4965 5965 4995 5995
rect 4725 5885 4755 5915
rect 4885 5885 4915 5915
rect 5045 5885 5075 5915
rect 4245 5765 4275 5795
rect 4405 5765 4435 5795
rect 4485 5765 4515 5795
rect 4645 5765 4675 5795
rect 4725 5765 4755 5795
rect 4885 5765 4915 5795
rect 5045 5765 5075 5795
rect 5125 5765 5155 5795
rect 5285 5765 5315 5795
rect 5445 5765 5475 5795
rect 5525 5765 5555 5795
rect 5685 5765 5715 5795
rect 5845 5765 5875 5795
rect 5925 5765 5955 5795
rect 6085 5765 6115 5795
rect 6165 5765 6195 5795
rect 6325 5765 6355 5795
rect 4245 5685 4275 5715
rect 4405 5685 4435 5715
rect 4485 5685 4515 5715
rect 4645 5685 4675 5715
rect 4725 5685 4755 5715
rect 4885 5685 4915 5715
rect 5045 5685 5075 5715
rect 5125 5685 5155 5715
rect 5285 5685 5315 5715
rect 5445 5685 5475 5715
rect 5525 5685 5555 5715
rect 5685 5685 5715 5715
rect 5845 5685 5875 5715
rect 5925 5685 5955 5715
rect 6085 5685 6115 5715
rect 6165 5685 6195 5715
rect 6325 5685 6355 5715
rect 4245 5605 4275 5635
rect 4405 5605 4435 5635
rect 4485 5605 4515 5635
rect 4645 5605 4675 5635
rect 4725 5605 4755 5635
rect 4885 5605 4915 5635
rect 5045 5605 5075 5635
rect 5125 5605 5155 5635
rect 5285 5605 5315 5635
rect 5445 5605 5475 5635
rect 5525 5605 5555 5635
rect 5685 5605 5715 5635
rect 5845 5605 5875 5635
rect 5925 5605 5955 5635
rect 6085 5605 6115 5635
rect 6165 5605 6195 5635
rect 6325 5605 6355 5635
rect 4245 5525 4275 5555
rect 4405 5525 4435 5555
rect 4485 5525 4515 5555
rect 4645 5525 4675 5555
rect 4725 5525 4755 5555
rect 4885 5525 4915 5555
rect 5045 5525 5075 5555
rect 5125 5525 5155 5555
rect 5285 5525 5315 5555
rect 5445 5525 5475 5555
rect 5525 5525 5555 5555
rect 5685 5525 5715 5555
rect 5845 5525 5875 5555
rect 5925 5525 5955 5555
rect 6085 5525 6115 5555
rect 6165 5525 6195 5555
rect 6325 5525 6355 5555
rect 4245 5445 4275 5475
rect 4405 5445 4435 5475
rect 4485 5445 4515 5475
rect 4645 5445 4675 5475
rect 4725 5445 4755 5475
rect 4885 5445 4915 5475
rect 5045 5445 5075 5475
rect 5125 5445 5155 5475
rect 5285 5445 5315 5475
rect 5445 5445 5475 5475
rect 5525 5445 5555 5475
rect 5685 5445 5715 5475
rect 5845 5445 5875 5475
rect 5925 5445 5955 5475
rect 6085 5445 6115 5475
rect 6165 5445 6195 5475
rect 6325 5445 6355 5475
rect 4245 5365 4275 5395
rect 4405 5365 4435 5395
rect 4485 5365 4515 5395
rect 4645 5365 4675 5395
rect 4725 5365 4755 5395
rect 4885 5365 4915 5395
rect 5045 5365 5075 5395
rect 5125 5365 5155 5395
rect 5285 5365 5315 5395
rect 5445 5365 5475 5395
rect 5525 5365 5555 5395
rect 5685 5365 5715 5395
rect 5845 5365 5875 5395
rect 5925 5365 5955 5395
rect 6085 5365 6115 5395
rect 6165 5365 6195 5395
rect 6325 5365 6355 5395
rect 4245 5285 4275 5315
rect 4405 5285 4435 5315
rect 4485 5285 4515 5315
rect 4645 5285 4675 5315
rect 4725 5285 4755 5315
rect 4885 5285 4915 5315
rect 5045 5285 5075 5315
rect 5125 5285 5155 5315
rect 5285 5285 5315 5315
rect 5445 5285 5475 5315
rect 5525 5285 5555 5315
rect 5685 5285 5715 5315
rect 5845 5285 5875 5315
rect 5925 5285 5955 5315
rect 6085 5285 6115 5315
rect 6165 5285 6195 5315
rect 6325 5285 6355 5315
rect 4245 5205 4275 5235
rect 4405 5205 4435 5235
rect 4485 5205 4515 5235
rect 4645 5205 4675 5235
rect 4725 5205 4755 5235
rect 4885 5205 4915 5235
rect 5045 5205 5075 5235
rect 5125 5205 5155 5235
rect 5285 5205 5315 5235
rect 5445 5205 5475 5235
rect 5525 5205 5555 5235
rect 5685 5205 5715 5235
rect 5845 5205 5875 5235
rect 5925 5205 5955 5235
rect 6085 5205 6115 5235
rect 6165 5205 6195 5235
rect 6325 5205 6355 5235
rect 4245 5125 4275 5155
rect 4405 5125 4435 5155
rect 4485 5125 4515 5155
rect 4645 5125 4675 5155
rect 4725 5125 4755 5155
rect 4885 5125 4915 5155
rect 5045 5125 5075 5155
rect 5125 5125 5155 5155
rect 5285 5125 5315 5155
rect 5445 5125 5475 5155
rect 5525 5125 5555 5155
rect 5685 5125 5715 5155
rect 5845 5125 5875 5155
rect 5925 5125 5955 5155
rect 6085 5125 6115 5155
rect 6165 5125 6195 5155
rect 6325 5125 6355 5155
rect 4245 5045 4275 5075
rect 4405 5045 4435 5075
rect 4485 5045 4515 5075
rect 4645 5045 4675 5075
rect 4725 5045 4755 5075
rect 4885 5045 4915 5075
rect 5045 5045 5075 5075
rect 5125 5045 5155 5075
rect 5285 5045 5315 5075
rect 5445 5045 5475 5075
rect 5525 5045 5555 5075
rect 5685 5045 5715 5075
rect 5845 5045 5875 5075
rect 5925 5045 5955 5075
rect 6085 5045 6115 5075
rect 6165 5045 6195 5075
rect 6325 5045 6355 5075
rect 4245 4965 4275 4995
rect 4405 4965 4435 4995
rect 4485 4965 4515 4995
rect 4645 4965 4675 4995
rect 4725 4965 4755 4995
rect 4885 4965 4915 4995
rect 5045 4965 5075 4995
rect 5125 4965 5155 4995
rect 5285 4965 5315 4995
rect 5445 4965 5475 4995
rect 5525 4965 5555 4995
rect 5685 4965 5715 4995
rect 5845 4965 5875 4995
rect 5925 4965 5955 4995
rect 6085 4965 6115 4995
rect 6165 4965 6195 4995
rect 6325 4965 6355 4995
rect 5925 4885 5955 4915
rect 6085 4885 6115 4915
rect 6005 4805 6035 4835
rect 5925 4725 5955 4755
rect 6085 4725 6115 4755
rect 6165 4645 6195 4675
rect 6325 4645 6355 4675
rect 6245 4565 6275 4595
rect 6165 4485 6195 4515
rect 6325 4485 6355 4515
rect 4245 4405 4275 4435
rect 4405 4405 4435 4435
rect 4485 4405 4515 4435
rect 4645 4405 4675 4435
rect 4725 4405 4755 4435
rect 4885 4405 4915 4435
rect 5045 4405 5075 4435
rect 5125 4405 5155 4435
rect 5285 4405 5315 4435
rect 5445 4405 5475 4435
rect 5525 4405 5555 4435
rect 5685 4405 5715 4435
rect 5845 4405 5875 4435
rect 5925 4405 5955 4435
rect 6085 4405 6115 4435
rect 6165 4405 6195 4435
rect 6325 4405 6355 4435
rect 4245 4325 4275 4355
rect 4405 4325 4435 4355
rect 4485 4325 4515 4355
rect 4645 4325 4675 4355
rect 4725 4325 4755 4355
rect 4885 4325 4915 4355
rect 5045 4325 5075 4355
rect 5125 4325 5155 4355
rect 5285 4325 5315 4355
rect 5445 4325 5475 4355
rect 5525 4325 5555 4355
rect 5685 4325 5715 4355
rect 5845 4325 5875 4355
rect 5925 4325 5955 4355
rect 6085 4325 6115 4355
rect 6165 4325 6195 4355
rect 6325 4325 6355 4355
rect 4245 4245 4275 4275
rect 4405 4245 4435 4275
rect 4485 4245 4515 4275
rect 4645 4245 4675 4275
rect 4725 4245 4755 4275
rect 4885 4245 4915 4275
rect 5045 4245 5075 4275
rect 5125 4245 5155 4275
rect 5285 4245 5315 4275
rect 5445 4245 5475 4275
rect 5525 4245 5555 4275
rect 5685 4245 5715 4275
rect 5845 4245 5875 4275
rect 5925 4245 5955 4275
rect 6085 4245 6115 4275
rect 6165 4245 6195 4275
rect 6325 4245 6355 4275
rect 4245 4165 4275 4195
rect 4405 4165 4435 4195
rect 4485 4165 4515 4195
rect 4645 4165 4675 4195
rect 4725 4165 4755 4195
rect 4885 4165 4915 4195
rect 5045 4165 5075 4195
rect 5125 4165 5155 4195
rect 5285 4165 5315 4195
rect 5445 4165 5475 4195
rect 5525 4165 5555 4195
rect 5685 4165 5715 4195
rect 5845 4165 5875 4195
rect 5925 4165 5955 4195
rect 6085 4165 6115 4195
rect 6165 4165 6195 4195
rect 6325 4165 6355 4195
rect 4245 4085 4275 4115
rect 4405 4085 4435 4115
rect 4485 4085 4515 4115
rect 4645 4085 4675 4115
rect 4725 4085 4755 4115
rect 4885 4085 4915 4115
rect 5045 4085 5075 4115
rect 5125 4085 5155 4115
rect 5285 4085 5315 4115
rect 5445 4085 5475 4115
rect 5525 4085 5555 4115
rect 5685 4085 5715 4115
rect 5845 4085 5875 4115
rect 5925 4085 5955 4115
rect 6085 4085 6115 4115
rect 6165 4085 6195 4115
rect 6325 4085 6355 4115
rect 4245 4005 4275 4035
rect 4405 4005 4435 4035
rect 4485 4005 4515 4035
rect 4645 4005 4675 4035
rect 4725 4005 4755 4035
rect 4885 4005 4915 4035
rect 5045 4005 5075 4035
rect 5125 4005 5155 4035
rect 5285 4005 5315 4035
rect 5445 4005 5475 4035
rect 5525 4005 5555 4035
rect 5685 4005 5715 4035
rect 5845 4005 5875 4035
rect 5925 4005 5955 4035
rect 6085 4005 6115 4035
rect 6165 4005 6195 4035
rect 6325 4005 6355 4035
rect 4245 3925 4275 3955
rect 4405 3925 4435 3955
rect 4485 3925 4515 3955
rect 4645 3925 4675 3955
rect 4725 3925 4755 3955
rect 4885 3925 4915 3955
rect 5045 3925 5075 3955
rect 5125 3925 5155 3955
rect 5285 3925 5315 3955
rect 5445 3925 5475 3955
rect 5525 3925 5555 3955
rect 5685 3925 5715 3955
rect 5845 3925 5875 3955
rect 5925 3925 5955 3955
rect 6085 3925 6115 3955
rect 6165 3925 6195 3955
rect 6325 3925 6355 3955
rect 4245 3845 4275 3875
rect 4405 3845 4435 3875
rect 4325 3765 4355 3795
rect 4245 3685 4275 3715
rect 4405 3685 4435 3715
rect 4485 3605 4515 3635
rect 4645 3605 4675 3635
rect 4565 3525 4595 3555
rect 4485 3445 4515 3475
rect 4645 3445 4675 3475
rect 5925 3365 5955 3395
rect 6085 3365 6115 3395
rect 6005 3285 6035 3315
rect 5925 3205 5955 3235
rect 6085 3205 6115 3235
rect 4245 3125 4275 3155
rect 4405 3125 4435 3155
rect 4485 3125 4515 3155
rect 4645 3125 4675 3155
rect 4725 3125 4755 3155
rect 4885 3125 4915 3155
rect 5045 3125 5075 3155
rect 5125 3125 5155 3155
rect 5285 3125 5315 3155
rect 5445 3125 5475 3155
rect 5525 3125 5555 3155
rect 5685 3125 5715 3155
rect 5845 3125 5875 3155
rect 5925 3125 5955 3155
rect 6085 3125 6115 3155
rect 6165 3125 6195 3155
rect 6325 3125 6355 3155
rect 4245 3045 4275 3075
rect 4405 3045 4435 3075
rect 4485 3045 4515 3075
rect 4645 3045 4675 3075
rect 4725 3045 4755 3075
rect 4885 3045 4915 3075
rect 5045 3045 5075 3075
rect 5125 3045 5155 3075
rect 5285 3045 5315 3075
rect 5445 3045 5475 3075
rect 5525 3045 5555 3075
rect 5685 3045 5715 3075
rect 5845 3045 5875 3075
rect 5925 3045 5955 3075
rect 6085 3045 6115 3075
rect 6165 3045 6195 3075
rect 6325 3045 6355 3075
rect 4245 2965 4275 2995
rect 4405 2965 4435 2995
rect 4485 2965 4515 2995
rect 4645 2965 4675 2995
rect 4725 2965 4755 2995
rect 4885 2965 4915 2995
rect 5045 2965 5075 2995
rect 5125 2965 5155 2995
rect 5285 2965 5315 2995
rect 5445 2965 5475 2995
rect 5525 2965 5555 2995
rect 5685 2965 5715 2995
rect 5845 2965 5875 2995
rect 5925 2965 5955 2995
rect 6085 2965 6115 2995
rect 6165 2965 6195 2995
rect 6325 2965 6355 2995
rect 4245 2885 4275 2915
rect 4405 2885 4435 2915
rect 4485 2885 4515 2915
rect 4645 2885 4675 2915
rect 4725 2885 4755 2915
rect 4885 2885 4915 2915
rect 5045 2885 5075 2915
rect 5125 2885 5155 2915
rect 5285 2885 5315 2915
rect 5445 2885 5475 2915
rect 5525 2885 5555 2915
rect 5685 2885 5715 2915
rect 5845 2885 5875 2915
rect 5925 2885 5955 2915
rect 6085 2885 6115 2915
rect 6165 2885 6195 2915
rect 6325 2885 6355 2915
rect 4245 2805 4275 2835
rect 4405 2805 4435 2835
rect 4485 2805 4515 2835
rect 4645 2805 4675 2835
rect 4725 2805 4755 2835
rect 4885 2805 4915 2835
rect 5045 2805 5075 2835
rect 5125 2805 5155 2835
rect 5285 2805 5315 2835
rect 5445 2805 5475 2835
rect 5525 2805 5555 2835
rect 5685 2805 5715 2835
rect 5845 2805 5875 2835
rect 5925 2805 5955 2835
rect 6085 2805 6115 2835
rect 6165 2805 6195 2835
rect 6325 2805 6355 2835
rect 4245 2725 4275 2755
rect 4405 2725 4435 2755
rect 4485 2725 4515 2755
rect 4645 2725 4675 2755
rect 4725 2725 4755 2755
rect 4885 2725 4915 2755
rect 5045 2725 5075 2755
rect 5125 2725 5155 2755
rect 5285 2725 5315 2755
rect 5445 2725 5475 2755
rect 5525 2725 5555 2755
rect 5685 2725 5715 2755
rect 5845 2725 5875 2755
rect 5925 2725 5955 2755
rect 6085 2725 6115 2755
rect 6165 2725 6195 2755
rect 6325 2725 6355 2755
rect 4245 2645 4275 2675
rect 4405 2645 4435 2675
rect 4485 2645 4515 2675
rect 4645 2645 4675 2675
rect 4725 2645 4755 2675
rect 4885 2645 4915 2675
rect 5045 2645 5075 2675
rect 5125 2645 5155 2675
rect 5285 2645 5315 2675
rect 5445 2645 5475 2675
rect 5525 2645 5555 2675
rect 5685 2645 5715 2675
rect 5845 2645 5875 2675
rect 5925 2645 5955 2675
rect 6085 2645 6115 2675
rect 6165 2645 6195 2675
rect 6325 2645 6355 2675
rect 4245 2565 4275 2595
rect 4405 2565 4435 2595
rect 4485 2565 4515 2595
rect 4645 2565 4675 2595
rect 4725 2565 4755 2595
rect 4885 2565 4915 2595
rect 5045 2565 5075 2595
rect 5125 2565 5155 2595
rect 5285 2565 5315 2595
rect 5445 2565 5475 2595
rect 5525 2565 5555 2595
rect 5685 2565 5715 2595
rect 5845 2565 5875 2595
rect 5925 2565 5955 2595
rect 6085 2565 6115 2595
rect 6165 2565 6195 2595
rect 6325 2565 6355 2595
rect 4245 2485 4275 2515
rect 4405 2485 4435 2515
rect 4485 2485 4515 2515
rect 4645 2485 4675 2515
rect 4725 2485 4755 2515
rect 4885 2485 4915 2515
rect 5045 2485 5075 2515
rect 5125 2485 5155 2515
rect 5285 2485 5315 2515
rect 5445 2485 5475 2515
rect 5525 2485 5555 2515
rect 5685 2485 5715 2515
rect 5845 2485 5875 2515
rect 5925 2485 5955 2515
rect 6085 2485 6115 2515
rect 6165 2485 6195 2515
rect 6325 2485 6355 2515
rect 4245 2405 4275 2435
rect 4405 2405 4435 2435
rect 4485 2405 4515 2435
rect 4645 2405 4675 2435
rect 4725 2405 4755 2435
rect 4885 2405 4915 2435
rect 5045 2405 5075 2435
rect 5125 2405 5155 2435
rect 5285 2405 5315 2435
rect 5445 2405 5475 2435
rect 5525 2405 5555 2435
rect 5685 2405 5715 2435
rect 5845 2405 5875 2435
rect 5925 2405 5955 2435
rect 6085 2405 6115 2435
rect 6165 2405 6195 2435
rect 6325 2405 6355 2435
rect 4245 2325 4275 2355
rect 4405 2325 4435 2355
rect 4485 2325 4515 2355
rect 4645 2325 4675 2355
rect 4725 2325 4755 2355
rect 4885 2325 4915 2355
rect 5045 2325 5075 2355
rect 5125 2325 5155 2355
rect 5285 2325 5315 2355
rect 5445 2325 5475 2355
rect 5525 2325 5555 2355
rect 5685 2325 5715 2355
rect 5845 2325 5875 2355
rect 5925 2325 5955 2355
rect 6085 2325 6115 2355
rect 6165 2325 6195 2355
rect 6325 2325 6355 2355
rect 4245 2245 4275 2275
rect 4405 2245 4435 2275
rect 4485 2245 4515 2275
rect 4645 2245 4675 2275
rect 4725 2245 4755 2275
rect 4885 2245 4915 2275
rect 5045 2245 5075 2275
rect 5125 2245 5155 2275
rect 5285 2245 5315 2275
rect 5445 2245 5475 2275
rect 5525 2245 5555 2275
rect 5685 2245 5715 2275
rect 5845 2245 5875 2275
rect 5925 2245 5955 2275
rect 6085 2245 6115 2275
rect 6165 2245 6195 2275
rect 6325 2245 6355 2275
rect 4245 2165 4275 2195
rect 4405 2165 4435 2195
rect 4485 2165 4515 2195
rect 4645 2165 4675 2195
rect 4725 2165 4755 2195
rect 4885 2165 4915 2195
rect 5045 2165 5075 2195
rect 5125 2165 5155 2195
rect 5285 2165 5315 2195
rect 5445 2165 5475 2195
rect 5525 2165 5555 2195
rect 5685 2165 5715 2195
rect 5845 2165 5875 2195
rect 5925 2165 5955 2195
rect 6085 2165 6115 2195
rect 6165 2165 6195 2195
rect 6325 2165 6355 2195
rect 4245 2085 4275 2115
rect 4405 2085 4435 2115
rect 4485 2085 4515 2115
rect 4645 2085 4675 2115
rect 4725 2085 4755 2115
rect 4885 2085 4915 2115
rect 5045 2085 5075 2115
rect 5125 2085 5155 2115
rect 5285 2085 5315 2115
rect 5445 2085 5475 2115
rect 5525 2085 5555 2115
rect 5685 2085 5715 2115
rect 5845 2085 5875 2115
rect 5925 2085 5955 2115
rect 6085 2085 6115 2115
rect 6165 2085 6195 2115
rect 6325 2085 6355 2115
rect 4245 2005 4275 2035
rect 4405 2005 4435 2035
rect 4485 2005 4515 2035
rect 4645 2005 4675 2035
rect 4725 2005 4755 2035
rect 4885 2005 4915 2035
rect 5045 2005 5075 2035
rect 5125 2005 5155 2035
rect 5285 2005 5315 2035
rect 5445 2005 5475 2035
rect 5525 2005 5555 2035
rect 5685 2005 5715 2035
rect 5845 2005 5875 2035
rect 5925 2005 5955 2035
rect 6085 2005 6115 2035
rect 6165 2005 6195 2035
rect 6325 2005 6355 2035
rect 4485 1885 4515 1915
rect 4645 1885 4675 1915
rect 4565 1805 4595 1835
rect 4485 1725 4515 1755
rect 4645 1725 4675 1755
rect 4245 1605 4275 1635
rect 4405 1605 4435 1635
rect 4485 1605 4515 1635
rect 4645 1605 4675 1635
rect 4725 1605 4755 1635
rect 4885 1605 4915 1635
rect 5045 1605 5075 1635
rect 5125 1605 5155 1635
rect 5285 1605 5315 1635
rect 5445 1605 5475 1635
rect 5525 1605 5555 1635
rect 5685 1605 5715 1635
rect 5845 1605 5875 1635
rect 5925 1605 5955 1635
rect 6085 1605 6115 1635
rect 6165 1605 6195 1635
rect 6325 1605 6355 1635
rect 4245 1525 4275 1555
rect 4405 1525 4435 1555
rect 4485 1525 4515 1555
rect 4645 1525 4675 1555
rect 4725 1525 4755 1555
rect 4885 1525 4915 1555
rect 5045 1525 5075 1555
rect 5125 1525 5155 1555
rect 5285 1525 5315 1555
rect 5445 1525 5475 1555
rect 5525 1525 5555 1555
rect 5685 1525 5715 1555
rect 5845 1525 5875 1555
rect 5925 1525 5955 1555
rect 6085 1525 6115 1555
rect 6165 1525 6195 1555
rect 6325 1525 6355 1555
rect 4245 1445 4275 1475
rect 4405 1445 4435 1475
rect 4485 1445 4515 1475
rect 4645 1445 4675 1475
rect 4725 1445 4755 1475
rect 4885 1445 4915 1475
rect 5045 1445 5075 1475
rect 5125 1445 5155 1475
rect 5285 1445 5315 1475
rect 5445 1445 5475 1475
rect 5525 1445 5555 1475
rect 5685 1445 5715 1475
rect 5845 1445 5875 1475
rect 5925 1445 5955 1475
rect 6085 1445 6115 1475
rect 6165 1445 6195 1475
rect 6325 1445 6355 1475
rect 4245 1365 4275 1395
rect 4405 1365 4435 1395
rect 4485 1365 4515 1395
rect 4645 1365 4675 1395
rect 4725 1365 4755 1395
rect 4885 1365 4915 1395
rect 5045 1365 5075 1395
rect 5125 1365 5155 1395
rect 5285 1365 5315 1395
rect 5445 1365 5475 1395
rect 5525 1365 5555 1395
rect 5685 1365 5715 1395
rect 5845 1365 5875 1395
rect 5925 1365 5955 1395
rect 6085 1365 6115 1395
rect 6165 1365 6195 1395
rect 6325 1365 6355 1395
rect 4245 1285 4275 1315
rect 4405 1285 4435 1315
rect 4485 1285 4515 1315
rect 4645 1285 4675 1315
rect 4725 1285 4755 1315
rect 4885 1285 4915 1315
rect 5045 1285 5075 1315
rect 5125 1285 5155 1315
rect 5285 1285 5315 1315
rect 5445 1285 5475 1315
rect 5525 1285 5555 1315
rect 5685 1285 5715 1315
rect 5845 1285 5875 1315
rect 5925 1285 5955 1315
rect 6085 1285 6115 1315
rect 6165 1285 6195 1315
rect 6325 1285 6355 1315
rect 4245 1205 4275 1235
rect 4405 1205 4435 1235
rect 4485 1205 4515 1235
rect 4645 1205 4675 1235
rect 4725 1205 4755 1235
rect 4885 1205 4915 1235
rect 5045 1205 5075 1235
rect 5125 1205 5155 1235
rect 5285 1205 5315 1235
rect 5445 1205 5475 1235
rect 5525 1205 5555 1235
rect 5685 1205 5715 1235
rect 5845 1205 5875 1235
rect 5925 1205 5955 1235
rect 6085 1205 6115 1235
rect 6165 1205 6195 1235
rect 6325 1205 6355 1235
rect 4245 1125 4275 1155
rect 4405 1125 4435 1155
rect 4485 1125 4515 1155
rect 4645 1125 4675 1155
rect 4725 1125 4755 1155
rect 4885 1125 4915 1155
rect 5045 1125 5075 1155
rect 5125 1125 5155 1155
rect 5285 1125 5315 1155
rect 5445 1125 5475 1155
rect 5525 1125 5555 1155
rect 5685 1125 5715 1155
rect 5845 1125 5875 1155
rect 5925 1125 5955 1155
rect 6085 1125 6115 1155
rect 6165 1125 6195 1155
rect 6325 1125 6355 1155
rect 4245 1045 4275 1075
rect 4405 1045 4435 1075
rect 4485 1045 4515 1075
rect 4645 1045 4675 1075
rect 4725 1045 4755 1075
rect 4885 1045 4915 1075
rect 5045 1045 5075 1075
rect 5125 1045 5155 1075
rect 5285 1045 5315 1075
rect 5445 1045 5475 1075
rect 5525 1045 5555 1075
rect 5685 1045 5715 1075
rect 5845 1045 5875 1075
rect 5925 1045 5955 1075
rect 6085 1045 6115 1075
rect 6165 1045 6195 1075
rect 6325 1045 6355 1075
rect 6165 965 6195 995
rect 6325 965 6355 995
rect 6245 885 6275 915
rect 6165 805 6195 835
rect 6325 805 6355 835
rect 4245 725 4275 755
rect 4405 725 4435 755
rect 4485 725 4515 755
rect 4645 725 4675 755
rect 4725 725 4755 755
rect 4885 725 4915 755
rect 5045 725 5075 755
rect 5125 725 5155 755
rect 5285 725 5315 755
rect 5445 725 5475 755
rect 5525 725 5555 755
rect 5685 725 5715 755
rect 5845 725 5875 755
rect 5925 725 5955 755
rect 6085 725 6115 755
rect 6165 725 6195 755
rect 6325 725 6355 755
rect 4245 645 4275 675
rect 4405 645 4435 675
rect 4485 645 4515 675
rect 4645 645 4675 675
rect 4725 645 4755 675
rect 4885 645 4915 675
rect 5045 645 5075 675
rect 5125 645 5155 675
rect 5285 645 5315 675
rect 5445 645 5475 675
rect 5525 645 5555 675
rect 5685 645 5715 675
rect 5845 645 5875 675
rect 5925 645 5955 675
rect 6085 645 6115 675
rect 6165 645 6195 675
rect 6325 645 6355 675
rect 4245 565 4275 595
rect 4405 565 4435 595
rect 4485 565 4515 595
rect 4645 565 4675 595
rect 4725 565 4755 595
rect 4885 565 4915 595
rect 5045 565 5075 595
rect 5125 565 5155 595
rect 5285 565 5315 595
rect 5445 565 5475 595
rect 5525 565 5555 595
rect 5685 565 5715 595
rect 5845 565 5875 595
rect 5925 565 5955 595
rect 6085 565 6115 595
rect 6165 565 6195 595
rect 6325 565 6355 595
rect 4245 445 4275 475
rect 4405 445 4435 475
rect 4325 365 4355 395
rect 4245 285 4275 315
rect 4405 285 4435 315
rect 4245 165 4275 195
rect 4405 165 4435 195
rect 4485 165 4515 195
rect 4645 165 4675 195
rect 4725 165 4755 195
rect 4885 165 4915 195
rect 5045 165 5075 195
rect 5125 165 5155 195
rect 5285 165 5315 195
rect 5445 165 5475 195
rect 5525 165 5555 195
rect 5685 165 5715 195
rect 5845 165 5875 195
rect 5925 165 5955 195
rect 6085 165 6115 195
rect 6165 165 6195 195
rect 6325 165 6355 195
rect 4245 85 4275 115
rect 4405 85 4435 115
rect 4485 85 4515 115
rect 4645 85 4675 115
rect 4725 85 4755 115
rect 4885 85 4915 115
rect 5045 85 5075 115
rect 5125 85 5155 115
rect 5285 85 5315 115
rect 5445 85 5475 115
rect 5525 85 5555 115
rect 5685 85 5715 115
rect 5845 85 5875 115
rect 5925 85 5955 115
rect 6085 85 6115 115
rect 6165 85 6195 115
rect 6325 85 6355 115
rect 4245 5 4275 35
rect 4405 5 4435 35
rect 4485 5 4515 35
rect 4645 5 4675 35
rect 4725 5 4755 35
rect 4885 5 4915 35
rect 5045 5 5075 35
rect 5125 5 5155 35
rect 5285 5 5315 35
rect 5445 5 5475 35
rect 5525 5 5555 35
rect 5685 5 5715 35
rect 5845 5 5875 35
rect 5925 5 5955 35
rect 6085 5 6115 35
rect 6165 5 6195 35
rect 6325 5 6355 35
<< metal3 >>
rect 0 16916 40 16920
rect 0 16884 4 16916
rect 36 16884 40 16916
rect 0 15476 40 16884
rect 0 15444 4 15476
rect 36 15444 40 15476
rect 0 14036 40 15444
rect 0 14004 4 14036
rect 36 14004 40 14036
rect 0 13716 40 14004
rect 80 16836 120 16920
rect 80 16804 84 16836
rect 116 16804 120 16836
rect 80 15556 120 16804
rect 80 15524 84 15556
rect 116 15524 120 15556
rect 80 13956 120 15524
rect 80 13924 84 13956
rect 116 13924 120 13956
rect 80 13796 120 13924
rect 80 13764 84 13796
rect 116 13764 120 13796
rect 80 13760 120 13764
rect 160 16756 200 16920
rect 160 16724 164 16756
rect 196 16724 200 16756
rect 160 13876 200 16724
rect 160 13844 164 13876
rect 196 13844 200 13876
rect 160 13760 200 13844
rect 240 16836 280 16920
rect 240 16804 244 16836
rect 276 16804 280 16836
rect 240 15556 280 16804
rect 240 15524 244 15556
rect 276 15524 280 15556
rect 240 13956 280 15524
rect 240 13924 244 13956
rect 276 13924 280 13956
rect 240 13796 280 13924
rect 240 13764 244 13796
rect 276 13764 280 13796
rect 240 13760 280 13764
rect 320 16916 360 16920
rect 320 16884 324 16916
rect 356 16884 360 16916
rect 320 15476 360 16884
rect 10240 16916 10280 16920
rect 10240 16884 10244 16916
rect 10276 16884 10280 16916
rect 400 16836 440 16840
rect 400 16804 404 16836
rect 436 16804 440 16836
rect 400 15556 440 16804
rect 10160 16836 10200 16840
rect 10160 16804 10164 16836
rect 10196 16804 10200 16836
rect 480 16756 520 16760
rect 480 16724 484 16756
rect 516 16724 520 16756
rect 480 16680 520 16724
rect 1520 16756 1560 16760
rect 1520 16724 1524 16756
rect 1556 16724 1560 16756
rect 1520 16680 1560 16724
rect 480 15600 1560 16680
rect 1600 16756 1640 16760
rect 1600 16724 1604 16756
rect 1636 16724 1640 16756
rect 1600 16680 1640 16724
rect 2640 16756 2680 16760
rect 2640 16724 2644 16756
rect 2676 16724 2680 16756
rect 2640 16680 2680 16724
rect 1600 15600 2680 16680
rect 2720 16756 2760 16760
rect 2720 16724 2724 16756
rect 2756 16724 2760 16756
rect 2720 16680 2760 16724
rect 3760 16756 3800 16760
rect 3760 16724 3764 16756
rect 3796 16724 3800 16756
rect 3760 16680 3800 16724
rect 2720 15600 3800 16680
rect 3840 16756 3880 16760
rect 3840 16724 3844 16756
rect 3876 16724 3880 16756
rect 3840 16680 3880 16724
rect 4880 16756 4920 16760
rect 4880 16724 4884 16756
rect 4916 16724 4920 16756
rect 4880 16680 4920 16724
rect 3840 15600 4920 16680
rect 5680 16756 5720 16760
rect 5680 16724 5684 16756
rect 5716 16724 5720 16756
rect 5680 16680 5720 16724
rect 6720 16756 6760 16760
rect 6720 16724 6724 16756
rect 6756 16724 6760 16756
rect 6720 16680 6760 16724
rect 5680 15600 6760 16680
rect 6800 16756 6840 16760
rect 6800 16724 6804 16756
rect 6836 16724 6840 16756
rect 6800 16680 6840 16724
rect 7840 16756 7880 16760
rect 7840 16724 7844 16756
rect 7876 16724 7880 16756
rect 7840 16680 7880 16724
rect 6800 15600 7880 16680
rect 7920 16756 7960 16760
rect 7920 16724 7924 16756
rect 7956 16724 7960 16756
rect 7920 16680 7960 16724
rect 8960 16756 9000 16760
rect 8960 16724 8964 16756
rect 8996 16724 9000 16756
rect 8960 16680 9000 16724
rect 7920 15600 9000 16680
rect 9040 16756 9080 16760
rect 9040 16724 9044 16756
rect 9076 16724 9080 16756
rect 9040 16680 9080 16724
rect 10080 16756 10120 16760
rect 10080 16724 10084 16756
rect 10116 16724 10120 16756
rect 10080 16680 10120 16724
rect 9040 15600 10120 16680
rect 400 15524 404 15556
rect 436 15524 440 15556
rect 400 15520 440 15524
rect 10160 15556 10200 16804
rect 10160 15524 10164 15556
rect 10196 15524 10200 15556
rect 10160 15520 10200 15524
rect 320 15444 324 15476
rect 356 15444 360 15476
rect 320 14036 360 15444
rect 10240 15476 10280 16884
rect 10240 15444 10244 15476
rect 10276 15444 10280 15476
rect 400 15396 440 15400
rect 400 15364 404 15396
rect 436 15364 440 15396
rect 400 14116 440 15364
rect 4960 15396 5000 15400
rect 4960 15364 4964 15396
rect 4996 15364 5000 15396
rect 480 15316 520 15320
rect 480 15284 484 15316
rect 516 15284 520 15316
rect 480 15240 520 15284
rect 1520 15316 1560 15320
rect 1520 15284 1524 15316
rect 1556 15284 1560 15316
rect 1520 15240 1560 15284
rect 480 14160 1560 15240
rect 1600 15316 1640 15320
rect 1600 15284 1604 15316
rect 1636 15284 1640 15316
rect 1600 15240 1640 15284
rect 2640 15316 2680 15320
rect 2640 15284 2644 15316
rect 2676 15284 2680 15316
rect 2640 15240 2680 15284
rect 1600 14160 2680 15240
rect 2720 15316 2760 15320
rect 2720 15284 2724 15316
rect 2756 15284 2760 15316
rect 2720 15240 2760 15284
rect 3760 15316 3800 15320
rect 3760 15284 3764 15316
rect 3796 15284 3800 15316
rect 3760 15240 3800 15284
rect 2720 14160 3800 15240
rect 3840 15316 3880 15320
rect 3840 15284 3844 15316
rect 3876 15284 3880 15316
rect 3840 15240 3880 15284
rect 4880 15316 4920 15320
rect 4880 15284 4884 15316
rect 4916 15284 4920 15316
rect 4880 15240 4920 15284
rect 3840 14160 4920 15240
rect 400 14084 404 14116
rect 436 14084 440 14116
rect 400 14080 440 14084
rect 4960 14116 5000 15364
rect 4960 14084 4964 14116
rect 4996 14084 5000 14116
rect 4960 14080 5000 14084
rect 320 14004 324 14036
rect 356 14004 360 14036
rect 0 13684 4 13716
rect 36 13684 40 13716
rect 0 13680 40 13684
rect 320 13716 360 14004
rect 5040 14036 5080 15400
rect 5040 14004 5044 14036
rect 5076 14004 5080 14036
rect 320 13684 324 13716
rect 356 13684 360 13716
rect 320 13680 360 13684
rect 4480 13956 4520 13960
rect 4480 13924 4484 13956
rect 4516 13924 4520 13956
rect 4480 13796 4520 13924
rect 4480 13764 4484 13796
rect 4516 13764 4520 13796
rect 4240 13636 4280 13640
rect 4240 13444 4244 13636
rect 4276 13444 4280 13636
rect 4240 12636 4280 13444
rect 4400 13636 4440 13640
rect 4400 13444 4404 13636
rect 4436 13444 4440 13636
rect 4240 12604 4244 12636
rect 4276 12604 4280 12636
rect 4240 12556 4280 12604
rect 4240 12524 4244 12556
rect 4276 12524 4280 12556
rect 4240 12476 4280 12524
rect 4240 12444 4244 12476
rect 4276 12444 4280 12476
rect 4240 12396 4280 12444
rect 4240 12364 4244 12396
rect 4276 12364 4280 12396
rect 4240 12316 4280 12364
rect 4240 12284 4244 12316
rect 4276 12284 4280 12316
rect 4240 12236 4280 12284
rect 4240 12204 4244 12236
rect 4276 12204 4280 12236
rect 4240 12156 4280 12204
rect 4240 12124 4244 12156
rect 4276 12124 4280 12156
rect 4240 11836 4280 12124
rect 4240 11804 4244 11836
rect 4276 11804 4280 11836
rect 4240 11756 4280 11804
rect 4240 11724 4244 11756
rect 4276 11724 4280 11756
rect 4240 11676 4280 11724
rect 4240 11644 4244 11676
rect 4276 11644 4280 11676
rect 4240 11596 4280 11644
rect 4240 11564 4244 11596
rect 4276 11564 4280 11596
rect 4240 11516 4280 11564
rect 4240 11484 4244 11516
rect 4276 11484 4280 11516
rect 4240 11436 4280 11484
rect 4240 11404 4244 11436
rect 4276 11404 4280 11436
rect 4240 10876 4280 11404
rect 4240 10844 4244 10876
rect 4276 10844 4280 10876
rect 4240 10796 4280 10844
rect 4240 10764 4244 10796
rect 4276 10764 4280 10796
rect 4240 10716 4280 10764
rect 4240 10684 4244 10716
rect 4276 10684 4280 10716
rect 4240 10636 4280 10684
rect 4240 10604 4244 10636
rect 4276 10604 4280 10636
rect 4240 10556 4280 10604
rect 4240 10524 4244 10556
rect 4276 10524 4280 10556
rect 4240 10476 4280 10524
rect 4240 10444 4244 10476
rect 4276 10444 4280 10476
rect 4240 10396 4280 10444
rect 4240 10364 4244 10396
rect 4276 10364 4280 10396
rect 4240 10316 4280 10364
rect 4240 10284 4244 10316
rect 4276 10284 4280 10316
rect 4240 10236 4280 10284
rect 4240 10204 4244 10236
rect 4276 10204 4280 10236
rect 4240 10156 4280 10204
rect 4240 10124 4244 10156
rect 4276 10124 4280 10156
rect 4240 10076 4280 10124
rect 4240 10044 4244 10076
rect 4276 10044 4280 10076
rect 4240 9996 4280 10044
rect 4240 9964 4244 9996
rect 4276 9964 4280 9996
rect 4240 9916 4280 9964
rect 4240 9884 4244 9916
rect 4276 9884 4280 9916
rect 4240 9836 4280 9884
rect 4240 9804 4244 9836
rect 4276 9804 4280 9836
rect 4240 9756 4280 9804
rect 4240 9724 4244 9756
rect 4276 9724 4280 9756
rect 4240 9356 4280 9724
rect 4240 9324 4244 9356
rect 4276 9324 4280 9356
rect 4240 9276 4280 9324
rect 4240 9244 4244 9276
rect 4276 9244 4280 9276
rect 4240 9196 4280 9244
rect 4240 9164 4244 9196
rect 4276 9164 4280 9196
rect 4240 8876 4280 9164
rect 4240 8844 4244 8876
rect 4276 8844 4280 8876
rect 4240 8796 4280 8844
rect 4240 8764 4244 8796
rect 4276 8764 4280 8796
rect 4240 8716 4280 8764
rect 4240 8684 4244 8716
rect 4276 8684 4280 8716
rect 4240 8636 4280 8684
rect 4240 8604 4244 8636
rect 4276 8604 4280 8636
rect 4240 8556 4280 8604
rect 4240 8524 4244 8556
rect 4276 8524 4280 8556
rect 4240 7636 4280 8524
rect 4240 7604 4244 7636
rect 4276 7604 4280 7636
rect 4240 7556 4280 7604
rect 4240 7524 4244 7556
rect 4276 7524 4280 7556
rect 4240 7476 4280 7524
rect 4240 7444 4244 7476
rect 4276 7444 4280 7476
rect 4240 7396 4280 7444
rect 4240 7364 4244 7396
rect 4276 7364 4280 7396
rect 4240 7316 4280 7364
rect 4240 7284 4244 7316
rect 4276 7284 4280 7316
rect 4240 7236 4280 7284
rect 4240 7204 4244 7236
rect 4276 7204 4280 7236
rect 4240 7156 4280 7204
rect 4240 7124 4244 7156
rect 4276 7124 4280 7156
rect 4240 7076 4280 7124
rect 4240 7044 4244 7076
rect 4276 7044 4280 7076
rect 4240 6756 4280 7044
rect 4240 6724 4244 6756
rect 4276 6724 4280 6756
rect 4240 6676 4280 6724
rect 4240 6644 4244 6676
rect 4276 6644 4280 6676
rect 4240 6596 4280 6644
rect 4240 6564 4244 6596
rect 4276 6564 4280 6596
rect 4240 6516 4280 6564
rect 4240 6484 4244 6516
rect 4276 6484 4280 6516
rect 4240 6436 4280 6484
rect 4240 6404 4244 6436
rect 4276 6404 4280 6436
rect 4240 6356 4280 6404
rect 4240 6324 4244 6356
rect 4276 6324 4280 6356
rect 4240 5796 4280 6324
rect 4240 5764 4244 5796
rect 4276 5764 4280 5796
rect 4240 5716 4280 5764
rect 4240 5684 4244 5716
rect 4276 5684 4280 5716
rect 4240 5636 4280 5684
rect 4240 5604 4244 5636
rect 4276 5604 4280 5636
rect 4240 5556 4280 5604
rect 4240 5524 4244 5556
rect 4276 5524 4280 5556
rect 4240 5476 4280 5524
rect 4240 5444 4244 5476
rect 4276 5444 4280 5476
rect 4240 5396 4280 5444
rect 4240 5364 4244 5396
rect 4276 5364 4280 5396
rect 4240 5316 4280 5364
rect 4240 5284 4244 5316
rect 4276 5284 4280 5316
rect 4240 5236 4280 5284
rect 4240 5204 4244 5236
rect 4276 5204 4280 5236
rect 4240 5156 4280 5204
rect 4240 5124 4244 5156
rect 4276 5124 4280 5156
rect 4240 5076 4280 5124
rect 4240 5044 4244 5076
rect 4276 5044 4280 5076
rect 4240 4996 4280 5044
rect 4240 4964 4244 4996
rect 4276 4964 4280 4996
rect 4240 4436 4280 4964
rect 4240 4404 4244 4436
rect 4276 4404 4280 4436
rect 4240 4356 4280 4404
rect 4240 4324 4244 4356
rect 4276 4324 4280 4356
rect 4240 4276 4280 4324
rect 4240 4244 4244 4276
rect 4276 4244 4280 4276
rect 4240 4196 4280 4244
rect 4240 4164 4244 4196
rect 4276 4164 4280 4196
rect 4240 4116 4280 4164
rect 4240 4084 4244 4116
rect 4276 4084 4280 4116
rect 4240 4036 4280 4084
rect 4240 4004 4244 4036
rect 4276 4004 4280 4036
rect 4240 3956 4280 4004
rect 4240 3924 4244 3956
rect 4276 3924 4280 3956
rect 4240 3875 4280 3924
rect 4240 3845 4245 3875
rect 4275 3845 4280 3875
rect 4240 3715 4280 3845
rect 4240 3685 4245 3715
rect 4275 3685 4280 3715
rect 4240 3156 4280 3685
rect 4240 3124 4244 3156
rect 4276 3124 4280 3156
rect 4240 3076 4280 3124
rect 4240 3044 4244 3076
rect 4276 3044 4280 3076
rect 4240 2996 4280 3044
rect 4240 2964 4244 2996
rect 4276 2964 4280 2996
rect 4240 2916 4280 2964
rect 4240 2884 4244 2916
rect 4276 2884 4280 2916
rect 4240 2836 4280 2884
rect 4240 2804 4244 2836
rect 4276 2804 4280 2836
rect 4240 2756 4280 2804
rect 4240 2724 4244 2756
rect 4276 2724 4280 2756
rect 4240 2676 4280 2724
rect 4240 2644 4244 2676
rect 4276 2644 4280 2676
rect 4240 2596 4280 2644
rect 4240 2564 4244 2596
rect 4276 2564 4280 2596
rect 4240 2516 4280 2564
rect 4240 2484 4244 2516
rect 4276 2484 4280 2516
rect 4240 2436 4280 2484
rect 4240 2404 4244 2436
rect 4276 2404 4280 2436
rect 4240 2356 4280 2404
rect 4240 2324 4244 2356
rect 4276 2324 4280 2356
rect 4240 2276 4280 2324
rect 4240 2244 4244 2276
rect 4276 2244 4280 2276
rect 4240 2196 4280 2244
rect 4240 2164 4244 2196
rect 4276 2164 4280 2196
rect 4240 2116 4280 2164
rect 4240 2084 4244 2116
rect 4276 2084 4280 2116
rect 4240 2036 4280 2084
rect 4240 2004 4244 2036
rect 4276 2004 4280 2036
rect 4240 1636 4280 2004
rect 4240 1604 4244 1636
rect 4276 1604 4280 1636
rect 4240 1556 4280 1604
rect 4240 1524 4244 1556
rect 4276 1524 4280 1556
rect 4240 1476 4280 1524
rect 4240 1444 4244 1476
rect 4276 1444 4280 1476
rect 4240 1396 4280 1444
rect 4240 1364 4244 1396
rect 4276 1364 4280 1396
rect 4240 1316 4280 1364
rect 4240 1284 4244 1316
rect 4276 1284 4280 1316
rect 4240 1236 4280 1284
rect 4240 1204 4244 1236
rect 4276 1204 4280 1236
rect 4240 1156 4280 1204
rect 4240 1124 4244 1156
rect 4276 1124 4280 1156
rect 4240 1076 4280 1124
rect 4240 1044 4244 1076
rect 4276 1044 4280 1076
rect 4240 756 4280 1044
rect 4240 724 4244 756
rect 4276 724 4280 756
rect 4240 676 4280 724
rect 4240 644 4244 676
rect 4276 644 4280 676
rect 4240 596 4280 644
rect 4240 564 4244 596
rect 4276 564 4280 596
rect 4240 475 4280 564
rect 4240 445 4245 475
rect 4275 445 4280 475
rect 4240 315 4280 445
rect 4240 285 4245 315
rect 4275 285 4280 315
rect 4240 196 4280 285
rect 4240 164 4244 196
rect 4276 164 4280 196
rect 4240 116 4280 164
rect 4240 84 4244 116
rect 4276 84 4280 116
rect 4240 36 4280 84
rect 4240 4 4244 36
rect 4276 4 4280 36
rect 4240 -40 4280 4
rect 4320 3795 4360 12680
rect 4320 3765 4325 3795
rect 4355 3765 4360 3795
rect 4320 395 4360 3765
rect 4320 365 4325 395
rect 4355 365 4360 395
rect 4320 -40 4360 365
rect 4400 12636 4440 13444
rect 4400 12604 4404 12636
rect 4436 12604 4440 12636
rect 4400 12556 4440 12604
rect 4400 12524 4404 12556
rect 4436 12524 4440 12556
rect 4400 12476 4440 12524
rect 4400 12444 4404 12476
rect 4436 12444 4440 12476
rect 4400 12396 4440 12444
rect 4400 12364 4404 12396
rect 4436 12364 4440 12396
rect 4400 12316 4440 12364
rect 4400 12284 4404 12316
rect 4436 12284 4440 12316
rect 4400 12236 4440 12284
rect 4400 12204 4404 12236
rect 4436 12204 4440 12236
rect 4400 12156 4440 12204
rect 4400 12124 4404 12156
rect 4436 12124 4440 12156
rect 4400 11836 4440 12124
rect 4400 11804 4404 11836
rect 4436 11804 4440 11836
rect 4400 11756 4440 11804
rect 4400 11724 4404 11756
rect 4436 11724 4440 11756
rect 4400 11676 4440 11724
rect 4400 11644 4404 11676
rect 4436 11644 4440 11676
rect 4400 11596 4440 11644
rect 4400 11564 4404 11596
rect 4436 11564 4440 11596
rect 4400 11516 4440 11564
rect 4400 11484 4404 11516
rect 4436 11484 4440 11516
rect 4400 11436 4440 11484
rect 4400 11404 4404 11436
rect 4436 11404 4440 11436
rect 4400 10876 4440 11404
rect 4400 10844 4404 10876
rect 4436 10844 4440 10876
rect 4400 10796 4440 10844
rect 4400 10764 4404 10796
rect 4436 10764 4440 10796
rect 4400 10716 4440 10764
rect 4400 10684 4404 10716
rect 4436 10684 4440 10716
rect 4400 10636 4440 10684
rect 4400 10604 4404 10636
rect 4436 10604 4440 10636
rect 4400 10556 4440 10604
rect 4400 10524 4404 10556
rect 4436 10524 4440 10556
rect 4400 10476 4440 10524
rect 4400 10444 4404 10476
rect 4436 10444 4440 10476
rect 4400 10396 4440 10444
rect 4400 10364 4404 10396
rect 4436 10364 4440 10396
rect 4400 10316 4440 10364
rect 4400 10284 4404 10316
rect 4436 10284 4440 10316
rect 4400 10236 4440 10284
rect 4400 10204 4404 10236
rect 4436 10204 4440 10236
rect 4400 10156 4440 10204
rect 4400 10124 4404 10156
rect 4436 10124 4440 10156
rect 4400 10076 4440 10124
rect 4400 10044 4404 10076
rect 4436 10044 4440 10076
rect 4400 9996 4440 10044
rect 4400 9964 4404 9996
rect 4436 9964 4440 9996
rect 4400 9916 4440 9964
rect 4400 9884 4404 9916
rect 4436 9884 4440 9916
rect 4400 9836 4440 9884
rect 4400 9804 4404 9836
rect 4436 9804 4440 9836
rect 4400 9756 4440 9804
rect 4400 9724 4404 9756
rect 4436 9724 4440 9756
rect 4400 9356 4440 9724
rect 4400 9324 4404 9356
rect 4436 9324 4440 9356
rect 4400 9276 4440 9324
rect 4400 9244 4404 9276
rect 4436 9244 4440 9276
rect 4400 9196 4440 9244
rect 4400 9164 4404 9196
rect 4436 9164 4440 9196
rect 4400 8876 4440 9164
rect 4400 8844 4404 8876
rect 4436 8844 4440 8876
rect 4400 8796 4440 8844
rect 4400 8764 4404 8796
rect 4436 8764 4440 8796
rect 4400 8716 4440 8764
rect 4400 8684 4404 8716
rect 4436 8684 4440 8716
rect 4400 8636 4440 8684
rect 4400 8604 4404 8636
rect 4436 8604 4440 8636
rect 4400 8556 4440 8604
rect 4400 8524 4404 8556
rect 4436 8524 4440 8556
rect 4400 7636 4440 8524
rect 4400 7604 4404 7636
rect 4436 7604 4440 7636
rect 4400 7556 4440 7604
rect 4400 7524 4404 7556
rect 4436 7524 4440 7556
rect 4400 7476 4440 7524
rect 4400 7444 4404 7476
rect 4436 7444 4440 7476
rect 4400 7396 4440 7444
rect 4400 7364 4404 7396
rect 4436 7364 4440 7396
rect 4400 7316 4440 7364
rect 4400 7284 4404 7316
rect 4436 7284 4440 7316
rect 4400 7236 4440 7284
rect 4400 7204 4404 7236
rect 4436 7204 4440 7236
rect 4400 7156 4440 7204
rect 4400 7124 4404 7156
rect 4436 7124 4440 7156
rect 4400 7076 4440 7124
rect 4400 7044 4404 7076
rect 4436 7044 4440 7076
rect 4400 6756 4440 7044
rect 4400 6724 4404 6756
rect 4436 6724 4440 6756
rect 4400 6676 4440 6724
rect 4400 6644 4404 6676
rect 4436 6644 4440 6676
rect 4400 6596 4440 6644
rect 4400 6564 4404 6596
rect 4436 6564 4440 6596
rect 4400 6516 4440 6564
rect 4400 6484 4404 6516
rect 4436 6484 4440 6516
rect 4400 6436 4440 6484
rect 4400 6404 4404 6436
rect 4436 6404 4440 6436
rect 4400 6356 4440 6404
rect 4400 6324 4404 6356
rect 4436 6324 4440 6356
rect 4400 5796 4440 6324
rect 4400 5764 4404 5796
rect 4436 5764 4440 5796
rect 4400 5716 4440 5764
rect 4400 5684 4404 5716
rect 4436 5684 4440 5716
rect 4400 5636 4440 5684
rect 4400 5604 4404 5636
rect 4436 5604 4440 5636
rect 4400 5556 4440 5604
rect 4400 5524 4404 5556
rect 4436 5524 4440 5556
rect 4400 5476 4440 5524
rect 4400 5444 4404 5476
rect 4436 5444 4440 5476
rect 4400 5396 4440 5444
rect 4400 5364 4404 5396
rect 4436 5364 4440 5396
rect 4400 5316 4440 5364
rect 4400 5284 4404 5316
rect 4436 5284 4440 5316
rect 4400 5236 4440 5284
rect 4400 5204 4404 5236
rect 4436 5204 4440 5236
rect 4400 5156 4440 5204
rect 4400 5124 4404 5156
rect 4436 5124 4440 5156
rect 4400 5076 4440 5124
rect 4400 5044 4404 5076
rect 4436 5044 4440 5076
rect 4400 4996 4440 5044
rect 4400 4964 4404 4996
rect 4436 4964 4440 4996
rect 4400 4436 4440 4964
rect 4400 4404 4404 4436
rect 4436 4404 4440 4436
rect 4400 4356 4440 4404
rect 4400 4324 4404 4356
rect 4436 4324 4440 4356
rect 4400 4276 4440 4324
rect 4400 4244 4404 4276
rect 4436 4244 4440 4276
rect 4400 4196 4440 4244
rect 4400 4164 4404 4196
rect 4436 4164 4440 4196
rect 4400 4116 4440 4164
rect 4400 4084 4404 4116
rect 4436 4084 4440 4116
rect 4400 4036 4440 4084
rect 4400 4004 4404 4036
rect 4436 4004 4440 4036
rect 4400 3956 4440 4004
rect 4400 3924 4404 3956
rect 4436 3924 4440 3956
rect 4400 3875 4440 3924
rect 4400 3845 4405 3875
rect 4435 3845 4440 3875
rect 4400 3715 4440 3845
rect 4400 3685 4405 3715
rect 4435 3685 4440 3715
rect 4400 3156 4440 3685
rect 4400 3124 4404 3156
rect 4436 3124 4440 3156
rect 4400 3076 4440 3124
rect 4400 3044 4404 3076
rect 4436 3044 4440 3076
rect 4400 2996 4440 3044
rect 4400 2964 4404 2996
rect 4436 2964 4440 2996
rect 4400 2916 4440 2964
rect 4400 2884 4404 2916
rect 4436 2884 4440 2916
rect 4400 2836 4440 2884
rect 4400 2804 4404 2836
rect 4436 2804 4440 2836
rect 4400 2756 4440 2804
rect 4400 2724 4404 2756
rect 4436 2724 4440 2756
rect 4400 2676 4440 2724
rect 4400 2644 4404 2676
rect 4436 2644 4440 2676
rect 4400 2596 4440 2644
rect 4400 2564 4404 2596
rect 4436 2564 4440 2596
rect 4400 2516 4440 2564
rect 4400 2484 4404 2516
rect 4436 2484 4440 2516
rect 4400 2436 4440 2484
rect 4400 2404 4404 2436
rect 4436 2404 4440 2436
rect 4400 2356 4440 2404
rect 4400 2324 4404 2356
rect 4436 2324 4440 2356
rect 4400 2276 4440 2324
rect 4400 2244 4404 2276
rect 4436 2244 4440 2276
rect 4400 2196 4440 2244
rect 4400 2164 4404 2196
rect 4436 2164 4440 2196
rect 4400 2116 4440 2164
rect 4400 2084 4404 2116
rect 4436 2084 4440 2116
rect 4400 2036 4440 2084
rect 4400 2004 4404 2036
rect 4436 2004 4440 2036
rect 4400 1636 4440 2004
rect 4400 1604 4404 1636
rect 4436 1604 4440 1636
rect 4400 1556 4440 1604
rect 4400 1524 4404 1556
rect 4436 1524 4440 1556
rect 4400 1476 4440 1524
rect 4400 1444 4404 1476
rect 4436 1444 4440 1476
rect 4400 1396 4440 1444
rect 4400 1364 4404 1396
rect 4436 1364 4440 1396
rect 4400 1316 4440 1364
rect 4400 1284 4404 1316
rect 4436 1284 4440 1316
rect 4400 1236 4440 1284
rect 4400 1204 4404 1236
rect 4436 1204 4440 1236
rect 4400 1156 4440 1204
rect 4400 1124 4404 1156
rect 4436 1124 4440 1156
rect 4400 1076 4440 1124
rect 4400 1044 4404 1076
rect 4436 1044 4440 1076
rect 4400 756 4440 1044
rect 4400 724 4404 756
rect 4436 724 4440 756
rect 4400 676 4440 724
rect 4400 644 4404 676
rect 4436 644 4440 676
rect 4400 596 4440 644
rect 4400 564 4404 596
rect 4436 564 4440 596
rect 4400 475 4440 564
rect 4400 445 4405 475
rect 4435 445 4440 475
rect 4400 315 4440 445
rect 4400 285 4405 315
rect 4435 285 4440 315
rect 4400 196 4440 285
rect 4400 164 4404 196
rect 4436 164 4440 196
rect 4400 116 4440 164
rect 4400 84 4404 116
rect 4436 84 4440 116
rect 4400 36 4440 84
rect 4400 4 4404 36
rect 4436 4 4440 36
rect 4400 -40 4440 4
rect 4480 13156 4520 13764
rect 4480 12964 4484 13156
rect 4516 12964 4520 13156
rect 4480 12636 4520 12964
rect 4480 12604 4484 12636
rect 4516 12604 4520 12636
rect 4480 12556 4520 12604
rect 4480 12524 4484 12556
rect 4516 12524 4520 12556
rect 4480 12476 4520 12524
rect 4480 12444 4484 12476
rect 4516 12444 4520 12476
rect 4480 12396 4520 12444
rect 4480 12364 4484 12396
rect 4516 12364 4520 12396
rect 4480 12316 4520 12364
rect 4480 12284 4484 12316
rect 4516 12284 4520 12316
rect 4480 12236 4520 12284
rect 4480 12204 4484 12236
rect 4516 12204 4520 12236
rect 4480 12156 4520 12204
rect 4480 12124 4484 12156
rect 4516 12124 4520 12156
rect 4480 12075 4520 12124
rect 4480 12045 4485 12075
rect 4515 12045 4520 12075
rect 4480 11915 4520 12045
rect 4480 11885 4485 11915
rect 4515 11885 4520 11915
rect 4480 11836 4520 11885
rect 4480 11804 4484 11836
rect 4516 11804 4520 11836
rect 4480 11756 4520 11804
rect 4480 11724 4484 11756
rect 4516 11724 4520 11756
rect 4480 11676 4520 11724
rect 4480 11644 4484 11676
rect 4516 11644 4520 11676
rect 4480 11596 4520 11644
rect 4480 11564 4484 11596
rect 4516 11564 4520 11596
rect 4480 11516 4520 11564
rect 4480 11484 4484 11516
rect 4516 11484 4520 11516
rect 4480 11436 4520 11484
rect 4480 11404 4484 11436
rect 4516 11404 4520 11436
rect 4480 10876 4520 11404
rect 4480 10844 4484 10876
rect 4516 10844 4520 10876
rect 4480 10796 4520 10844
rect 4480 10764 4484 10796
rect 4516 10764 4520 10796
rect 4480 10716 4520 10764
rect 4480 10684 4484 10716
rect 4516 10684 4520 10716
rect 4480 10636 4520 10684
rect 4480 10604 4484 10636
rect 4516 10604 4520 10636
rect 4480 10556 4520 10604
rect 4480 10524 4484 10556
rect 4516 10524 4520 10556
rect 4480 10476 4520 10524
rect 4480 10444 4484 10476
rect 4516 10444 4520 10476
rect 4480 10396 4520 10444
rect 4480 10364 4484 10396
rect 4516 10364 4520 10396
rect 4480 10316 4520 10364
rect 4480 10284 4484 10316
rect 4516 10284 4520 10316
rect 4480 10236 4520 10284
rect 4480 10204 4484 10236
rect 4516 10204 4520 10236
rect 4480 10156 4520 10204
rect 4480 10124 4484 10156
rect 4516 10124 4520 10156
rect 4480 10076 4520 10124
rect 4480 10044 4484 10076
rect 4516 10044 4520 10076
rect 4480 9996 4520 10044
rect 4480 9964 4484 9996
rect 4516 9964 4520 9996
rect 4480 9916 4520 9964
rect 4480 9884 4484 9916
rect 4516 9884 4520 9916
rect 4480 9836 4520 9884
rect 4480 9804 4484 9836
rect 4516 9804 4520 9836
rect 4480 9756 4520 9804
rect 4480 9724 4484 9756
rect 4516 9724 4520 9756
rect 4480 9635 4520 9724
rect 4480 9605 4485 9635
rect 4515 9605 4520 9635
rect 4480 9475 4520 9605
rect 4480 9445 4485 9475
rect 4515 9445 4520 9475
rect 4480 9356 4520 9445
rect 4480 9324 4484 9356
rect 4516 9324 4520 9356
rect 4480 9276 4520 9324
rect 4480 9244 4484 9276
rect 4516 9244 4520 9276
rect 4480 9196 4520 9244
rect 4480 9164 4484 9196
rect 4516 9164 4520 9196
rect 4480 8876 4520 9164
rect 4480 8844 4484 8876
rect 4516 8844 4520 8876
rect 4480 8796 4520 8844
rect 4480 8764 4484 8796
rect 4516 8764 4520 8796
rect 4480 8716 4520 8764
rect 4480 8684 4484 8716
rect 4516 8684 4520 8716
rect 4480 8636 4520 8684
rect 4480 8604 4484 8636
rect 4516 8604 4520 8636
rect 4480 8556 4520 8604
rect 4480 8524 4484 8556
rect 4516 8524 4520 8556
rect 4480 7636 4520 8524
rect 4480 7604 4484 7636
rect 4516 7604 4520 7636
rect 4480 7556 4520 7604
rect 4480 7524 4484 7556
rect 4516 7524 4520 7556
rect 4480 7476 4520 7524
rect 4480 7444 4484 7476
rect 4516 7444 4520 7476
rect 4480 7396 4520 7444
rect 4480 7364 4484 7396
rect 4516 7364 4520 7396
rect 4480 7316 4520 7364
rect 4480 7284 4484 7316
rect 4516 7284 4520 7316
rect 4480 7236 4520 7284
rect 4480 7204 4484 7236
rect 4516 7204 4520 7236
rect 4480 7156 4520 7204
rect 4480 7124 4484 7156
rect 4516 7124 4520 7156
rect 4480 7076 4520 7124
rect 4480 7044 4484 7076
rect 4516 7044 4520 7076
rect 4480 6995 4520 7044
rect 4480 6965 4485 6995
rect 4515 6965 4520 6995
rect 4480 6835 4520 6965
rect 4480 6805 4485 6835
rect 4515 6805 4520 6835
rect 4480 6756 4520 6805
rect 4480 6724 4484 6756
rect 4516 6724 4520 6756
rect 4480 6676 4520 6724
rect 4480 6644 4484 6676
rect 4516 6644 4520 6676
rect 4480 6596 4520 6644
rect 4480 6564 4484 6596
rect 4516 6564 4520 6596
rect 4480 6516 4520 6564
rect 4480 6484 4484 6516
rect 4516 6484 4520 6516
rect 4480 6436 4520 6484
rect 4480 6404 4484 6436
rect 4516 6404 4520 6436
rect 4480 6356 4520 6404
rect 4480 6324 4484 6356
rect 4516 6324 4520 6356
rect 4480 5796 4520 6324
rect 4480 5764 4484 5796
rect 4516 5764 4520 5796
rect 4480 5716 4520 5764
rect 4480 5684 4484 5716
rect 4516 5684 4520 5716
rect 4480 5636 4520 5684
rect 4480 5604 4484 5636
rect 4516 5604 4520 5636
rect 4480 5556 4520 5604
rect 4480 5524 4484 5556
rect 4516 5524 4520 5556
rect 4480 5476 4520 5524
rect 4480 5444 4484 5476
rect 4516 5444 4520 5476
rect 4480 5396 4520 5444
rect 4480 5364 4484 5396
rect 4516 5364 4520 5396
rect 4480 5316 4520 5364
rect 4480 5284 4484 5316
rect 4516 5284 4520 5316
rect 4480 5236 4520 5284
rect 4480 5204 4484 5236
rect 4516 5204 4520 5236
rect 4480 5156 4520 5204
rect 4480 5124 4484 5156
rect 4516 5124 4520 5156
rect 4480 5076 4520 5124
rect 4480 5044 4484 5076
rect 4516 5044 4520 5076
rect 4480 4996 4520 5044
rect 4480 4964 4484 4996
rect 4516 4964 4520 4996
rect 4480 4436 4520 4964
rect 4480 4404 4484 4436
rect 4516 4404 4520 4436
rect 4480 4356 4520 4404
rect 4480 4324 4484 4356
rect 4516 4324 4520 4356
rect 4480 4276 4520 4324
rect 4480 4244 4484 4276
rect 4516 4244 4520 4276
rect 4480 4196 4520 4244
rect 4480 4164 4484 4196
rect 4516 4164 4520 4196
rect 4480 4116 4520 4164
rect 4480 4084 4484 4116
rect 4516 4084 4520 4116
rect 4480 4036 4520 4084
rect 4480 4004 4484 4036
rect 4516 4004 4520 4036
rect 4480 3956 4520 4004
rect 4480 3924 4484 3956
rect 4516 3924 4520 3956
rect 4480 3635 4520 3924
rect 4480 3605 4485 3635
rect 4515 3605 4520 3635
rect 4480 3475 4520 3605
rect 4480 3445 4485 3475
rect 4515 3445 4520 3475
rect 4480 3156 4520 3445
rect 4480 3124 4484 3156
rect 4516 3124 4520 3156
rect 4480 3076 4520 3124
rect 4480 3044 4484 3076
rect 4516 3044 4520 3076
rect 4480 2996 4520 3044
rect 4480 2964 4484 2996
rect 4516 2964 4520 2996
rect 4480 2916 4520 2964
rect 4480 2884 4484 2916
rect 4516 2884 4520 2916
rect 4480 2836 4520 2884
rect 4480 2804 4484 2836
rect 4516 2804 4520 2836
rect 4480 2756 4520 2804
rect 4480 2724 4484 2756
rect 4516 2724 4520 2756
rect 4480 2676 4520 2724
rect 4480 2644 4484 2676
rect 4516 2644 4520 2676
rect 4480 2596 4520 2644
rect 4480 2564 4484 2596
rect 4516 2564 4520 2596
rect 4480 2516 4520 2564
rect 4480 2484 4484 2516
rect 4516 2484 4520 2516
rect 4480 2436 4520 2484
rect 4480 2404 4484 2436
rect 4516 2404 4520 2436
rect 4480 2356 4520 2404
rect 4480 2324 4484 2356
rect 4516 2324 4520 2356
rect 4480 2276 4520 2324
rect 4480 2244 4484 2276
rect 4516 2244 4520 2276
rect 4480 2196 4520 2244
rect 4480 2164 4484 2196
rect 4516 2164 4520 2196
rect 4480 2116 4520 2164
rect 4480 2084 4484 2116
rect 4516 2084 4520 2116
rect 4480 2036 4520 2084
rect 4480 2004 4484 2036
rect 4516 2004 4520 2036
rect 4480 1915 4520 2004
rect 4480 1885 4485 1915
rect 4515 1885 4520 1915
rect 4480 1755 4520 1885
rect 4480 1725 4485 1755
rect 4515 1725 4520 1755
rect 4480 1636 4520 1725
rect 4480 1604 4484 1636
rect 4516 1604 4520 1636
rect 4480 1556 4520 1604
rect 4480 1524 4484 1556
rect 4516 1524 4520 1556
rect 4480 1476 4520 1524
rect 4480 1444 4484 1476
rect 4516 1444 4520 1476
rect 4480 1396 4520 1444
rect 4480 1364 4484 1396
rect 4516 1364 4520 1396
rect 4480 1316 4520 1364
rect 4480 1284 4484 1316
rect 4516 1284 4520 1316
rect 4480 1236 4520 1284
rect 4480 1204 4484 1236
rect 4516 1204 4520 1236
rect 4480 1156 4520 1204
rect 4480 1124 4484 1156
rect 4516 1124 4520 1156
rect 4480 1076 4520 1124
rect 4480 1044 4484 1076
rect 4516 1044 4520 1076
rect 4480 756 4520 1044
rect 4480 724 4484 756
rect 4516 724 4520 756
rect 4480 676 4520 724
rect 4480 644 4484 676
rect 4516 644 4520 676
rect 4480 596 4520 644
rect 4480 564 4484 596
rect 4516 564 4520 596
rect 4480 196 4520 564
rect 4480 164 4484 196
rect 4516 164 4520 196
rect 4480 116 4520 164
rect 4480 84 4484 116
rect 4516 84 4520 116
rect 4480 36 4520 84
rect 4480 4 4484 36
rect 4516 4 4520 36
rect 4480 -40 4520 4
rect 4560 13876 4600 13960
rect 4560 13844 4564 13876
rect 4596 13844 4600 13876
rect 4560 11995 4600 13844
rect 4560 11965 4565 11995
rect 4595 11965 4600 11995
rect 4560 9555 4600 11965
rect 4560 9525 4565 9555
rect 4595 9525 4600 9555
rect 4560 6915 4600 9525
rect 4560 6885 4565 6915
rect 4595 6885 4600 6915
rect 4560 3555 4600 6885
rect 4560 3525 4565 3555
rect 4595 3525 4600 3555
rect 4560 1835 4600 3525
rect 4560 1805 4565 1835
rect 4595 1805 4600 1835
rect 4560 -40 4600 1805
rect 4640 13956 4680 13960
rect 4640 13924 4644 13956
rect 4676 13924 4680 13956
rect 4640 13796 4680 13924
rect 4640 13764 4644 13796
rect 4676 13764 4680 13796
rect 4640 13156 4680 13764
rect 5040 13716 5080 14004
rect 5040 13684 5044 13716
rect 5076 13684 5080 13716
rect 4640 12964 4644 13156
rect 4676 12964 4680 13156
rect 4640 12636 4680 12964
rect 4640 12604 4644 12636
rect 4676 12604 4680 12636
rect 4640 12556 4680 12604
rect 4640 12524 4644 12556
rect 4676 12524 4680 12556
rect 4640 12476 4680 12524
rect 4640 12444 4644 12476
rect 4676 12444 4680 12476
rect 4640 12396 4680 12444
rect 4640 12364 4644 12396
rect 4676 12364 4680 12396
rect 4640 12316 4680 12364
rect 4640 12284 4644 12316
rect 4676 12284 4680 12316
rect 4640 12236 4680 12284
rect 4640 12204 4644 12236
rect 4676 12204 4680 12236
rect 4640 12156 4680 12204
rect 4640 12124 4644 12156
rect 4676 12124 4680 12156
rect 4640 12075 4680 12124
rect 4640 12045 4645 12075
rect 4675 12045 4680 12075
rect 4640 11915 4680 12045
rect 4640 11885 4645 11915
rect 4675 11885 4680 11915
rect 4640 11836 4680 11885
rect 4640 11804 4644 11836
rect 4676 11804 4680 11836
rect 4640 11756 4680 11804
rect 4640 11724 4644 11756
rect 4676 11724 4680 11756
rect 4640 11676 4680 11724
rect 4640 11644 4644 11676
rect 4676 11644 4680 11676
rect 4640 11596 4680 11644
rect 4640 11564 4644 11596
rect 4676 11564 4680 11596
rect 4640 11516 4680 11564
rect 4640 11484 4644 11516
rect 4676 11484 4680 11516
rect 4640 11436 4680 11484
rect 4640 11404 4644 11436
rect 4676 11404 4680 11436
rect 4640 10876 4680 11404
rect 4640 10844 4644 10876
rect 4676 10844 4680 10876
rect 4640 10796 4680 10844
rect 4640 10764 4644 10796
rect 4676 10764 4680 10796
rect 4640 10716 4680 10764
rect 4640 10684 4644 10716
rect 4676 10684 4680 10716
rect 4640 10636 4680 10684
rect 4640 10604 4644 10636
rect 4676 10604 4680 10636
rect 4640 10556 4680 10604
rect 4640 10524 4644 10556
rect 4676 10524 4680 10556
rect 4640 10476 4680 10524
rect 4640 10444 4644 10476
rect 4676 10444 4680 10476
rect 4640 10396 4680 10444
rect 4640 10364 4644 10396
rect 4676 10364 4680 10396
rect 4640 10316 4680 10364
rect 4640 10284 4644 10316
rect 4676 10284 4680 10316
rect 4640 10236 4680 10284
rect 4640 10204 4644 10236
rect 4676 10204 4680 10236
rect 4640 10156 4680 10204
rect 4640 10124 4644 10156
rect 4676 10124 4680 10156
rect 4640 10076 4680 10124
rect 4640 10044 4644 10076
rect 4676 10044 4680 10076
rect 4640 9996 4680 10044
rect 4640 9964 4644 9996
rect 4676 9964 4680 9996
rect 4640 9916 4680 9964
rect 4640 9884 4644 9916
rect 4676 9884 4680 9916
rect 4640 9836 4680 9884
rect 4640 9804 4644 9836
rect 4676 9804 4680 9836
rect 4640 9756 4680 9804
rect 4640 9724 4644 9756
rect 4676 9724 4680 9756
rect 4640 9635 4680 9724
rect 4640 9605 4645 9635
rect 4675 9605 4680 9635
rect 4640 9475 4680 9605
rect 4640 9445 4645 9475
rect 4675 9445 4680 9475
rect 4640 9356 4680 9445
rect 4640 9324 4644 9356
rect 4676 9324 4680 9356
rect 4640 9276 4680 9324
rect 4640 9244 4644 9276
rect 4676 9244 4680 9276
rect 4640 9196 4680 9244
rect 4640 9164 4644 9196
rect 4676 9164 4680 9196
rect 4640 8876 4680 9164
rect 4640 8844 4644 8876
rect 4676 8844 4680 8876
rect 4640 8796 4680 8844
rect 4640 8764 4644 8796
rect 4676 8764 4680 8796
rect 4640 8716 4680 8764
rect 4640 8684 4644 8716
rect 4676 8684 4680 8716
rect 4640 8636 4680 8684
rect 4640 8604 4644 8636
rect 4676 8604 4680 8636
rect 4640 8556 4680 8604
rect 4640 8524 4644 8556
rect 4676 8524 4680 8556
rect 4640 7636 4680 8524
rect 4640 7604 4644 7636
rect 4676 7604 4680 7636
rect 4640 7556 4680 7604
rect 4640 7524 4644 7556
rect 4676 7524 4680 7556
rect 4640 7476 4680 7524
rect 4640 7444 4644 7476
rect 4676 7444 4680 7476
rect 4640 7396 4680 7444
rect 4640 7364 4644 7396
rect 4676 7364 4680 7396
rect 4640 7316 4680 7364
rect 4640 7284 4644 7316
rect 4676 7284 4680 7316
rect 4640 7236 4680 7284
rect 4640 7204 4644 7236
rect 4676 7204 4680 7236
rect 4640 7156 4680 7204
rect 4640 7124 4644 7156
rect 4676 7124 4680 7156
rect 4640 7076 4680 7124
rect 4640 7044 4644 7076
rect 4676 7044 4680 7076
rect 4640 6995 4680 7044
rect 4640 6965 4645 6995
rect 4675 6965 4680 6995
rect 4640 6835 4680 6965
rect 4640 6805 4645 6835
rect 4675 6805 4680 6835
rect 4640 6756 4680 6805
rect 4640 6724 4644 6756
rect 4676 6724 4680 6756
rect 4640 6676 4680 6724
rect 4640 6644 4644 6676
rect 4676 6644 4680 6676
rect 4640 6596 4680 6644
rect 4640 6564 4644 6596
rect 4676 6564 4680 6596
rect 4640 6516 4680 6564
rect 4640 6484 4644 6516
rect 4676 6484 4680 6516
rect 4640 6436 4680 6484
rect 4640 6404 4644 6436
rect 4676 6404 4680 6436
rect 4640 6356 4680 6404
rect 4640 6324 4644 6356
rect 4676 6324 4680 6356
rect 4640 5796 4680 6324
rect 4640 5764 4644 5796
rect 4676 5764 4680 5796
rect 4640 5716 4680 5764
rect 4640 5684 4644 5716
rect 4676 5684 4680 5716
rect 4640 5636 4680 5684
rect 4640 5604 4644 5636
rect 4676 5604 4680 5636
rect 4640 5556 4680 5604
rect 4640 5524 4644 5556
rect 4676 5524 4680 5556
rect 4640 5476 4680 5524
rect 4640 5444 4644 5476
rect 4676 5444 4680 5476
rect 4640 5396 4680 5444
rect 4640 5364 4644 5396
rect 4676 5364 4680 5396
rect 4640 5316 4680 5364
rect 4640 5284 4644 5316
rect 4676 5284 4680 5316
rect 4640 5236 4680 5284
rect 4640 5204 4644 5236
rect 4676 5204 4680 5236
rect 4640 5156 4680 5204
rect 4640 5124 4644 5156
rect 4676 5124 4680 5156
rect 4640 5076 4680 5124
rect 4640 5044 4644 5076
rect 4676 5044 4680 5076
rect 4640 4996 4680 5044
rect 4640 4964 4644 4996
rect 4676 4964 4680 4996
rect 4640 4436 4680 4964
rect 4640 4404 4644 4436
rect 4676 4404 4680 4436
rect 4640 4356 4680 4404
rect 4640 4324 4644 4356
rect 4676 4324 4680 4356
rect 4640 4276 4680 4324
rect 4640 4244 4644 4276
rect 4676 4244 4680 4276
rect 4640 4196 4680 4244
rect 4640 4164 4644 4196
rect 4676 4164 4680 4196
rect 4640 4116 4680 4164
rect 4640 4084 4644 4116
rect 4676 4084 4680 4116
rect 4640 4036 4680 4084
rect 4640 4004 4644 4036
rect 4676 4004 4680 4036
rect 4640 3956 4680 4004
rect 4640 3924 4644 3956
rect 4676 3924 4680 3956
rect 4640 3635 4680 3924
rect 4640 3605 4645 3635
rect 4675 3605 4680 3635
rect 4640 3475 4680 3605
rect 4640 3445 4645 3475
rect 4675 3445 4680 3475
rect 4640 3156 4680 3445
rect 4640 3124 4644 3156
rect 4676 3124 4680 3156
rect 4640 3076 4680 3124
rect 4640 3044 4644 3076
rect 4676 3044 4680 3076
rect 4640 2996 4680 3044
rect 4640 2964 4644 2996
rect 4676 2964 4680 2996
rect 4640 2916 4680 2964
rect 4640 2884 4644 2916
rect 4676 2884 4680 2916
rect 4640 2836 4680 2884
rect 4640 2804 4644 2836
rect 4676 2804 4680 2836
rect 4640 2756 4680 2804
rect 4640 2724 4644 2756
rect 4676 2724 4680 2756
rect 4640 2676 4680 2724
rect 4640 2644 4644 2676
rect 4676 2644 4680 2676
rect 4640 2596 4680 2644
rect 4640 2564 4644 2596
rect 4676 2564 4680 2596
rect 4640 2516 4680 2564
rect 4640 2484 4644 2516
rect 4676 2484 4680 2516
rect 4640 2436 4680 2484
rect 4640 2404 4644 2436
rect 4676 2404 4680 2436
rect 4640 2356 4680 2404
rect 4640 2324 4644 2356
rect 4676 2324 4680 2356
rect 4640 2276 4680 2324
rect 4640 2244 4644 2276
rect 4676 2244 4680 2276
rect 4640 2196 4680 2244
rect 4640 2164 4644 2196
rect 4676 2164 4680 2196
rect 4640 2116 4680 2164
rect 4640 2084 4644 2116
rect 4676 2084 4680 2116
rect 4640 2036 4680 2084
rect 4640 2004 4644 2036
rect 4676 2004 4680 2036
rect 4640 1915 4680 2004
rect 4640 1885 4645 1915
rect 4675 1885 4680 1915
rect 4640 1755 4680 1885
rect 4640 1725 4645 1755
rect 4675 1725 4680 1755
rect 4640 1636 4680 1725
rect 4640 1604 4644 1636
rect 4676 1604 4680 1636
rect 4640 1556 4680 1604
rect 4640 1524 4644 1556
rect 4676 1524 4680 1556
rect 4640 1476 4680 1524
rect 4640 1444 4644 1476
rect 4676 1444 4680 1476
rect 4640 1396 4680 1444
rect 4640 1364 4644 1396
rect 4676 1364 4680 1396
rect 4640 1316 4680 1364
rect 4640 1284 4644 1316
rect 4676 1284 4680 1316
rect 4640 1236 4680 1284
rect 4640 1204 4644 1236
rect 4676 1204 4680 1236
rect 4640 1156 4680 1204
rect 4640 1124 4644 1156
rect 4676 1124 4680 1156
rect 4640 1076 4680 1124
rect 4640 1044 4644 1076
rect 4676 1044 4680 1076
rect 4640 756 4680 1044
rect 4640 724 4644 756
rect 4676 724 4680 756
rect 4640 676 4680 724
rect 4640 644 4644 676
rect 4676 644 4680 676
rect 4640 596 4680 644
rect 4640 564 4644 596
rect 4676 564 4680 596
rect 4640 196 4680 564
rect 4640 164 4644 196
rect 4676 164 4680 196
rect 4640 116 4680 164
rect 4640 84 4644 116
rect 4676 84 4680 116
rect 4640 36 4680 84
rect 4640 4 4644 36
rect 4676 4 4680 36
rect 4640 -40 4680 4
rect 4720 13396 4760 13400
rect 4720 13204 4724 13396
rect 4756 13204 4760 13396
rect 4720 12636 4760 13204
rect 4880 13396 4920 13400
rect 4880 13204 4884 13396
rect 4916 13204 4920 13396
rect 4720 12604 4724 12636
rect 4756 12604 4760 12636
rect 4720 12556 4760 12604
rect 4720 12524 4724 12556
rect 4756 12524 4760 12556
rect 4720 12476 4760 12524
rect 4720 12444 4724 12476
rect 4756 12444 4760 12476
rect 4720 12396 4760 12444
rect 4720 12364 4724 12396
rect 4756 12364 4760 12396
rect 4720 12316 4760 12364
rect 4720 12284 4724 12316
rect 4756 12284 4760 12316
rect 4720 12236 4760 12284
rect 4720 12204 4724 12236
rect 4756 12204 4760 12236
rect 4720 12156 4760 12204
rect 4720 12124 4724 12156
rect 4756 12124 4760 12156
rect 4720 11836 4760 12124
rect 4720 11804 4724 11836
rect 4756 11804 4760 11836
rect 4720 11756 4760 11804
rect 4720 11724 4724 11756
rect 4756 11724 4760 11756
rect 4720 11676 4760 11724
rect 4720 11644 4724 11676
rect 4756 11644 4760 11676
rect 4720 11596 4760 11644
rect 4720 11564 4724 11596
rect 4756 11564 4760 11596
rect 4720 11516 4760 11564
rect 4720 11484 4724 11516
rect 4756 11484 4760 11516
rect 4720 11436 4760 11484
rect 4720 11404 4724 11436
rect 4756 11404 4760 11436
rect 4720 10876 4760 11404
rect 4720 10844 4724 10876
rect 4756 10844 4760 10876
rect 4720 10796 4760 10844
rect 4720 10764 4724 10796
rect 4756 10764 4760 10796
rect 4720 10716 4760 10764
rect 4720 10684 4724 10716
rect 4756 10684 4760 10716
rect 4720 10636 4760 10684
rect 4720 10604 4724 10636
rect 4756 10604 4760 10636
rect 4720 10556 4760 10604
rect 4720 10524 4724 10556
rect 4756 10524 4760 10556
rect 4720 10476 4760 10524
rect 4720 10444 4724 10476
rect 4756 10444 4760 10476
rect 4720 10396 4760 10444
rect 4720 10364 4724 10396
rect 4756 10364 4760 10396
rect 4720 10316 4760 10364
rect 4720 10284 4724 10316
rect 4756 10284 4760 10316
rect 4720 10236 4760 10284
rect 4720 10204 4724 10236
rect 4756 10204 4760 10236
rect 4720 10156 4760 10204
rect 4720 10124 4724 10156
rect 4756 10124 4760 10156
rect 4720 10076 4760 10124
rect 4720 10044 4724 10076
rect 4756 10044 4760 10076
rect 4720 9996 4760 10044
rect 4720 9964 4724 9996
rect 4756 9964 4760 9996
rect 4720 9916 4760 9964
rect 4720 9884 4724 9916
rect 4756 9884 4760 9916
rect 4720 9836 4760 9884
rect 4720 9804 4724 9836
rect 4756 9804 4760 9836
rect 4720 9756 4760 9804
rect 4720 9724 4724 9756
rect 4756 9724 4760 9756
rect 4720 9356 4760 9724
rect 4720 9324 4724 9356
rect 4756 9324 4760 9356
rect 4720 9276 4760 9324
rect 4720 9244 4724 9276
rect 4756 9244 4760 9276
rect 4720 9196 4760 9244
rect 4720 9164 4724 9196
rect 4756 9164 4760 9196
rect 4720 8876 4760 9164
rect 4720 8844 4724 8876
rect 4756 8844 4760 8876
rect 4720 8796 4760 8844
rect 4720 8764 4724 8796
rect 4756 8764 4760 8796
rect 4720 8716 4760 8764
rect 4720 8684 4724 8716
rect 4756 8684 4760 8716
rect 4720 8636 4760 8684
rect 4720 8604 4724 8636
rect 4756 8604 4760 8636
rect 4720 8556 4760 8604
rect 4720 8524 4724 8556
rect 4756 8524 4760 8556
rect 4720 7636 4760 8524
rect 4720 7604 4724 7636
rect 4756 7604 4760 7636
rect 4720 7556 4760 7604
rect 4720 7524 4724 7556
rect 4756 7524 4760 7556
rect 4720 7476 4760 7524
rect 4720 7444 4724 7476
rect 4756 7444 4760 7476
rect 4720 7396 4760 7444
rect 4720 7364 4724 7396
rect 4756 7364 4760 7396
rect 4720 7316 4760 7364
rect 4720 7284 4724 7316
rect 4756 7284 4760 7316
rect 4720 7236 4760 7284
rect 4720 7204 4724 7236
rect 4756 7204 4760 7236
rect 4720 7156 4760 7204
rect 4720 7124 4724 7156
rect 4756 7124 4760 7156
rect 4720 7076 4760 7124
rect 4720 7044 4724 7076
rect 4756 7044 4760 7076
rect 4720 6756 4760 7044
rect 4720 6724 4724 6756
rect 4756 6724 4760 6756
rect 4720 6676 4760 6724
rect 4720 6644 4724 6676
rect 4756 6644 4760 6676
rect 4720 6596 4760 6644
rect 4720 6564 4724 6596
rect 4756 6564 4760 6596
rect 4720 6516 4760 6564
rect 4720 6484 4724 6516
rect 4756 6484 4760 6516
rect 4720 6436 4760 6484
rect 4720 6404 4724 6436
rect 4756 6404 4760 6436
rect 4720 6356 4760 6404
rect 4720 6324 4724 6356
rect 4756 6324 4760 6356
rect 4720 6235 4760 6324
rect 4720 6205 4725 6235
rect 4755 6205 4760 6235
rect 4720 6075 4760 6205
rect 4720 6045 4725 6075
rect 4755 6045 4760 6075
rect 4720 5915 4760 6045
rect 4720 5885 4725 5915
rect 4755 5885 4760 5915
rect 4720 5796 4760 5885
rect 4720 5764 4724 5796
rect 4756 5764 4760 5796
rect 4720 5716 4760 5764
rect 4720 5684 4724 5716
rect 4756 5684 4760 5716
rect 4720 5636 4760 5684
rect 4720 5604 4724 5636
rect 4756 5604 4760 5636
rect 4720 5556 4760 5604
rect 4720 5524 4724 5556
rect 4756 5524 4760 5556
rect 4720 5476 4760 5524
rect 4720 5444 4724 5476
rect 4756 5444 4760 5476
rect 4720 5396 4760 5444
rect 4720 5364 4724 5396
rect 4756 5364 4760 5396
rect 4720 5316 4760 5364
rect 4720 5284 4724 5316
rect 4756 5284 4760 5316
rect 4720 5236 4760 5284
rect 4720 5204 4724 5236
rect 4756 5204 4760 5236
rect 4720 5156 4760 5204
rect 4720 5124 4724 5156
rect 4756 5124 4760 5156
rect 4720 5076 4760 5124
rect 4720 5044 4724 5076
rect 4756 5044 4760 5076
rect 4720 4996 4760 5044
rect 4720 4964 4724 4996
rect 4756 4964 4760 4996
rect 4720 4436 4760 4964
rect 4720 4404 4724 4436
rect 4756 4404 4760 4436
rect 4720 4356 4760 4404
rect 4720 4324 4724 4356
rect 4756 4324 4760 4356
rect 4720 4276 4760 4324
rect 4720 4244 4724 4276
rect 4756 4244 4760 4276
rect 4720 4196 4760 4244
rect 4720 4164 4724 4196
rect 4756 4164 4760 4196
rect 4720 4116 4760 4164
rect 4720 4084 4724 4116
rect 4756 4084 4760 4116
rect 4720 4036 4760 4084
rect 4720 4004 4724 4036
rect 4756 4004 4760 4036
rect 4720 3956 4760 4004
rect 4720 3924 4724 3956
rect 4756 3924 4760 3956
rect 4720 3156 4760 3924
rect 4720 3124 4724 3156
rect 4756 3124 4760 3156
rect 4720 3076 4760 3124
rect 4720 3044 4724 3076
rect 4756 3044 4760 3076
rect 4720 2996 4760 3044
rect 4720 2964 4724 2996
rect 4756 2964 4760 2996
rect 4720 2916 4760 2964
rect 4720 2884 4724 2916
rect 4756 2884 4760 2916
rect 4720 2836 4760 2884
rect 4720 2804 4724 2836
rect 4756 2804 4760 2836
rect 4720 2756 4760 2804
rect 4720 2724 4724 2756
rect 4756 2724 4760 2756
rect 4720 2676 4760 2724
rect 4720 2644 4724 2676
rect 4756 2644 4760 2676
rect 4720 2596 4760 2644
rect 4720 2564 4724 2596
rect 4756 2564 4760 2596
rect 4720 2516 4760 2564
rect 4720 2484 4724 2516
rect 4756 2484 4760 2516
rect 4720 2436 4760 2484
rect 4720 2404 4724 2436
rect 4756 2404 4760 2436
rect 4720 2356 4760 2404
rect 4720 2324 4724 2356
rect 4756 2324 4760 2356
rect 4720 2276 4760 2324
rect 4720 2244 4724 2276
rect 4756 2244 4760 2276
rect 4720 2196 4760 2244
rect 4720 2164 4724 2196
rect 4756 2164 4760 2196
rect 4720 2116 4760 2164
rect 4720 2084 4724 2116
rect 4756 2084 4760 2116
rect 4720 2036 4760 2084
rect 4720 2004 4724 2036
rect 4756 2004 4760 2036
rect 4720 1636 4760 2004
rect 4720 1604 4724 1636
rect 4756 1604 4760 1636
rect 4720 1556 4760 1604
rect 4720 1524 4724 1556
rect 4756 1524 4760 1556
rect 4720 1476 4760 1524
rect 4720 1444 4724 1476
rect 4756 1444 4760 1476
rect 4720 1396 4760 1444
rect 4720 1364 4724 1396
rect 4756 1364 4760 1396
rect 4720 1316 4760 1364
rect 4720 1284 4724 1316
rect 4756 1284 4760 1316
rect 4720 1236 4760 1284
rect 4720 1204 4724 1236
rect 4756 1204 4760 1236
rect 4720 1156 4760 1204
rect 4720 1124 4724 1156
rect 4756 1124 4760 1156
rect 4720 1076 4760 1124
rect 4720 1044 4724 1076
rect 4756 1044 4760 1076
rect 4720 756 4760 1044
rect 4720 724 4724 756
rect 4756 724 4760 756
rect 4720 676 4760 724
rect 4720 644 4724 676
rect 4756 644 4760 676
rect 4720 596 4760 644
rect 4720 564 4724 596
rect 4756 564 4760 596
rect 4720 196 4760 564
rect 4720 164 4724 196
rect 4756 164 4760 196
rect 4720 116 4760 164
rect 4720 84 4724 116
rect 4756 84 4760 116
rect 4720 36 4760 84
rect 4720 4 4724 36
rect 4756 4 4760 36
rect 4720 -40 4760 4
rect 4800 6155 4840 12680
rect 4800 6125 4805 6155
rect 4835 6125 4840 6155
rect 4800 -40 4840 6125
rect 4880 12636 4920 13204
rect 5040 13396 5080 13684
rect 5040 13204 5044 13396
rect 5076 13204 5080 13396
rect 4880 12604 4884 12636
rect 4916 12604 4920 12636
rect 4880 12556 4920 12604
rect 4880 12524 4884 12556
rect 4916 12524 4920 12556
rect 4880 12476 4920 12524
rect 4880 12444 4884 12476
rect 4916 12444 4920 12476
rect 4880 12396 4920 12444
rect 4880 12364 4884 12396
rect 4916 12364 4920 12396
rect 4880 12316 4920 12364
rect 4880 12284 4884 12316
rect 4916 12284 4920 12316
rect 4880 12236 4920 12284
rect 4880 12204 4884 12236
rect 4916 12204 4920 12236
rect 4880 12156 4920 12204
rect 4880 12124 4884 12156
rect 4916 12124 4920 12156
rect 4880 11836 4920 12124
rect 4880 11804 4884 11836
rect 4916 11804 4920 11836
rect 4880 11756 4920 11804
rect 4880 11724 4884 11756
rect 4916 11724 4920 11756
rect 4880 11676 4920 11724
rect 4880 11644 4884 11676
rect 4916 11644 4920 11676
rect 4880 11596 4920 11644
rect 4880 11564 4884 11596
rect 4916 11564 4920 11596
rect 4880 11516 4920 11564
rect 4880 11484 4884 11516
rect 4916 11484 4920 11516
rect 4880 11436 4920 11484
rect 4880 11404 4884 11436
rect 4916 11404 4920 11436
rect 4880 10876 4920 11404
rect 4880 10844 4884 10876
rect 4916 10844 4920 10876
rect 4880 10796 4920 10844
rect 4880 10764 4884 10796
rect 4916 10764 4920 10796
rect 4880 10716 4920 10764
rect 4880 10684 4884 10716
rect 4916 10684 4920 10716
rect 4880 10636 4920 10684
rect 4880 10604 4884 10636
rect 4916 10604 4920 10636
rect 4880 10556 4920 10604
rect 4880 10524 4884 10556
rect 4916 10524 4920 10556
rect 4880 10476 4920 10524
rect 4880 10444 4884 10476
rect 4916 10444 4920 10476
rect 4880 10396 4920 10444
rect 4880 10364 4884 10396
rect 4916 10364 4920 10396
rect 4880 10316 4920 10364
rect 4880 10284 4884 10316
rect 4916 10284 4920 10316
rect 4880 10236 4920 10284
rect 4880 10204 4884 10236
rect 4916 10204 4920 10236
rect 4880 10156 4920 10204
rect 4880 10124 4884 10156
rect 4916 10124 4920 10156
rect 4880 10076 4920 10124
rect 4880 10044 4884 10076
rect 4916 10044 4920 10076
rect 4880 9996 4920 10044
rect 4880 9964 4884 9996
rect 4916 9964 4920 9996
rect 4880 9916 4920 9964
rect 4880 9884 4884 9916
rect 4916 9884 4920 9916
rect 4880 9836 4920 9884
rect 4880 9804 4884 9836
rect 4916 9804 4920 9836
rect 4880 9756 4920 9804
rect 4880 9724 4884 9756
rect 4916 9724 4920 9756
rect 4880 9356 4920 9724
rect 4880 9324 4884 9356
rect 4916 9324 4920 9356
rect 4880 9276 4920 9324
rect 4880 9244 4884 9276
rect 4916 9244 4920 9276
rect 4880 9196 4920 9244
rect 4880 9164 4884 9196
rect 4916 9164 4920 9196
rect 4880 8876 4920 9164
rect 4880 8844 4884 8876
rect 4916 8844 4920 8876
rect 4880 8796 4920 8844
rect 4880 8764 4884 8796
rect 4916 8764 4920 8796
rect 4880 8716 4920 8764
rect 4880 8684 4884 8716
rect 4916 8684 4920 8716
rect 4880 8636 4920 8684
rect 4880 8604 4884 8636
rect 4916 8604 4920 8636
rect 4880 8556 4920 8604
rect 4880 8524 4884 8556
rect 4916 8524 4920 8556
rect 4880 8475 4920 8524
rect 4880 8445 4885 8475
rect 4915 8445 4920 8475
rect 4880 8315 4920 8445
rect 4880 8285 4885 8315
rect 4915 8285 4920 8315
rect 4880 7636 4920 8285
rect 4880 7604 4884 7636
rect 4916 7604 4920 7636
rect 4880 7556 4920 7604
rect 4880 7524 4884 7556
rect 4916 7524 4920 7556
rect 4880 7476 4920 7524
rect 4880 7444 4884 7476
rect 4916 7444 4920 7476
rect 4880 7396 4920 7444
rect 4880 7364 4884 7396
rect 4916 7364 4920 7396
rect 4880 7316 4920 7364
rect 4880 7284 4884 7316
rect 4916 7284 4920 7316
rect 4880 7236 4920 7284
rect 4880 7204 4884 7236
rect 4916 7204 4920 7236
rect 4880 7156 4920 7204
rect 4880 7124 4884 7156
rect 4916 7124 4920 7156
rect 4880 7076 4920 7124
rect 4880 7044 4884 7076
rect 4916 7044 4920 7076
rect 4880 6756 4920 7044
rect 4880 6724 4884 6756
rect 4916 6724 4920 6756
rect 4880 6676 4920 6724
rect 4880 6644 4884 6676
rect 4916 6644 4920 6676
rect 4880 6596 4920 6644
rect 4880 6564 4884 6596
rect 4916 6564 4920 6596
rect 4880 6516 4920 6564
rect 4880 6484 4884 6516
rect 4916 6484 4920 6516
rect 4880 6436 4920 6484
rect 4880 6404 4884 6436
rect 4916 6404 4920 6436
rect 4880 6356 4920 6404
rect 4880 6324 4884 6356
rect 4916 6324 4920 6356
rect 4880 6235 4920 6324
rect 4880 6205 4885 6235
rect 4915 6205 4920 6235
rect 4880 6075 4920 6205
rect 4880 6045 4885 6075
rect 4915 6045 4920 6075
rect 4880 5915 4920 6045
rect 4880 5885 4885 5915
rect 4915 5885 4920 5915
rect 4880 5796 4920 5885
rect 4880 5764 4884 5796
rect 4916 5764 4920 5796
rect 4880 5716 4920 5764
rect 4880 5684 4884 5716
rect 4916 5684 4920 5716
rect 4880 5636 4920 5684
rect 4880 5604 4884 5636
rect 4916 5604 4920 5636
rect 4880 5556 4920 5604
rect 4880 5524 4884 5556
rect 4916 5524 4920 5556
rect 4880 5476 4920 5524
rect 4880 5444 4884 5476
rect 4916 5444 4920 5476
rect 4880 5396 4920 5444
rect 4880 5364 4884 5396
rect 4916 5364 4920 5396
rect 4880 5316 4920 5364
rect 4880 5284 4884 5316
rect 4916 5284 4920 5316
rect 4880 5236 4920 5284
rect 4880 5204 4884 5236
rect 4916 5204 4920 5236
rect 4880 5156 4920 5204
rect 4880 5124 4884 5156
rect 4916 5124 4920 5156
rect 4880 5076 4920 5124
rect 4880 5044 4884 5076
rect 4916 5044 4920 5076
rect 4880 4996 4920 5044
rect 4880 4964 4884 4996
rect 4916 4964 4920 4996
rect 4880 4436 4920 4964
rect 4880 4404 4884 4436
rect 4916 4404 4920 4436
rect 4880 4356 4920 4404
rect 4880 4324 4884 4356
rect 4916 4324 4920 4356
rect 4880 4276 4920 4324
rect 4880 4244 4884 4276
rect 4916 4244 4920 4276
rect 4880 4196 4920 4244
rect 4880 4164 4884 4196
rect 4916 4164 4920 4196
rect 4880 4116 4920 4164
rect 4880 4084 4884 4116
rect 4916 4084 4920 4116
rect 4880 4036 4920 4084
rect 4880 4004 4884 4036
rect 4916 4004 4920 4036
rect 4880 3956 4920 4004
rect 4880 3924 4884 3956
rect 4916 3924 4920 3956
rect 4880 3156 4920 3924
rect 4880 3124 4884 3156
rect 4916 3124 4920 3156
rect 4880 3076 4920 3124
rect 4880 3044 4884 3076
rect 4916 3044 4920 3076
rect 4880 2996 4920 3044
rect 4880 2964 4884 2996
rect 4916 2964 4920 2996
rect 4880 2916 4920 2964
rect 4880 2884 4884 2916
rect 4916 2884 4920 2916
rect 4880 2836 4920 2884
rect 4880 2804 4884 2836
rect 4916 2804 4920 2836
rect 4880 2756 4920 2804
rect 4880 2724 4884 2756
rect 4916 2724 4920 2756
rect 4880 2676 4920 2724
rect 4880 2644 4884 2676
rect 4916 2644 4920 2676
rect 4880 2596 4920 2644
rect 4880 2564 4884 2596
rect 4916 2564 4920 2596
rect 4880 2516 4920 2564
rect 4880 2484 4884 2516
rect 4916 2484 4920 2516
rect 4880 2436 4920 2484
rect 4880 2404 4884 2436
rect 4916 2404 4920 2436
rect 4880 2356 4920 2404
rect 4880 2324 4884 2356
rect 4916 2324 4920 2356
rect 4880 2276 4920 2324
rect 4880 2244 4884 2276
rect 4916 2244 4920 2276
rect 4880 2196 4920 2244
rect 4880 2164 4884 2196
rect 4916 2164 4920 2196
rect 4880 2116 4920 2164
rect 4880 2084 4884 2116
rect 4916 2084 4920 2116
rect 4880 2036 4920 2084
rect 4880 2004 4884 2036
rect 4916 2004 4920 2036
rect 4880 1636 4920 2004
rect 4880 1604 4884 1636
rect 4916 1604 4920 1636
rect 4880 1556 4920 1604
rect 4880 1524 4884 1556
rect 4916 1524 4920 1556
rect 4880 1476 4920 1524
rect 4880 1444 4884 1476
rect 4916 1444 4920 1476
rect 4880 1396 4920 1444
rect 4880 1364 4884 1396
rect 4916 1364 4920 1396
rect 4880 1316 4920 1364
rect 4880 1284 4884 1316
rect 4916 1284 4920 1316
rect 4880 1236 4920 1284
rect 4880 1204 4884 1236
rect 4916 1204 4920 1236
rect 4880 1156 4920 1204
rect 4880 1124 4884 1156
rect 4916 1124 4920 1156
rect 4880 1076 4920 1124
rect 4880 1044 4884 1076
rect 4916 1044 4920 1076
rect 4880 756 4920 1044
rect 4880 724 4884 756
rect 4916 724 4920 756
rect 4880 676 4920 724
rect 4880 644 4884 676
rect 4916 644 4920 676
rect 4880 596 4920 644
rect 4880 564 4884 596
rect 4916 564 4920 596
rect 4880 196 4920 564
rect 4880 164 4884 196
rect 4916 164 4920 196
rect 4880 116 4920 164
rect 4880 84 4884 116
rect 4916 84 4920 116
rect 4880 36 4920 84
rect 4880 4 4884 36
rect 4916 4 4920 36
rect 4880 -40 4920 4
rect 4960 8395 5000 12680
rect 4960 8365 4965 8395
rect 4995 8365 5000 8395
rect 4960 6155 5000 8365
rect 4960 6125 4965 6155
rect 4995 6125 5000 6155
rect 4960 5995 5000 6125
rect 4960 5965 4965 5995
rect 4995 5965 5000 5995
rect 4960 -40 5000 5965
rect 5040 12636 5080 13204
rect 5040 12604 5044 12636
rect 5076 12604 5080 12636
rect 5040 12556 5080 12604
rect 5040 12524 5044 12556
rect 5076 12524 5080 12556
rect 5040 12476 5080 12524
rect 5040 12444 5044 12476
rect 5076 12444 5080 12476
rect 5040 12396 5080 12444
rect 5040 12364 5044 12396
rect 5076 12364 5080 12396
rect 5040 12316 5080 12364
rect 5040 12284 5044 12316
rect 5076 12284 5080 12316
rect 5040 12236 5080 12284
rect 5040 12204 5044 12236
rect 5076 12204 5080 12236
rect 5040 12156 5080 12204
rect 5040 12124 5044 12156
rect 5076 12124 5080 12156
rect 5040 11836 5080 12124
rect 5040 11804 5044 11836
rect 5076 11804 5080 11836
rect 5040 11756 5080 11804
rect 5040 11724 5044 11756
rect 5076 11724 5080 11756
rect 5040 11676 5080 11724
rect 5040 11644 5044 11676
rect 5076 11644 5080 11676
rect 5040 11596 5080 11644
rect 5040 11564 5044 11596
rect 5076 11564 5080 11596
rect 5040 11516 5080 11564
rect 5040 11484 5044 11516
rect 5076 11484 5080 11516
rect 5040 11436 5080 11484
rect 5040 11404 5044 11436
rect 5076 11404 5080 11436
rect 5040 11155 5080 11404
rect 5040 11125 5045 11155
rect 5075 11125 5080 11155
rect 5040 10995 5080 11125
rect 5040 10965 5045 10995
rect 5075 10965 5080 10995
rect 5040 10876 5080 10965
rect 5040 10844 5044 10876
rect 5076 10844 5080 10876
rect 5040 10796 5080 10844
rect 5040 10764 5044 10796
rect 5076 10764 5080 10796
rect 5040 10716 5080 10764
rect 5040 10684 5044 10716
rect 5076 10684 5080 10716
rect 5040 10636 5080 10684
rect 5040 10604 5044 10636
rect 5076 10604 5080 10636
rect 5040 10556 5080 10604
rect 5040 10524 5044 10556
rect 5076 10524 5080 10556
rect 5040 10476 5080 10524
rect 5040 10444 5044 10476
rect 5076 10444 5080 10476
rect 5040 10396 5080 10444
rect 5040 10364 5044 10396
rect 5076 10364 5080 10396
rect 5040 10316 5080 10364
rect 5040 10284 5044 10316
rect 5076 10284 5080 10316
rect 5040 10236 5080 10284
rect 5040 10204 5044 10236
rect 5076 10204 5080 10236
rect 5040 10156 5080 10204
rect 5040 10124 5044 10156
rect 5076 10124 5080 10156
rect 5040 10076 5080 10124
rect 5040 10044 5044 10076
rect 5076 10044 5080 10076
rect 5040 9996 5080 10044
rect 5040 9964 5044 9996
rect 5076 9964 5080 9996
rect 5040 9916 5080 9964
rect 5040 9884 5044 9916
rect 5076 9884 5080 9916
rect 5040 9836 5080 9884
rect 5040 9804 5044 9836
rect 5076 9804 5080 9836
rect 5040 9756 5080 9804
rect 5040 9724 5044 9756
rect 5076 9724 5080 9756
rect 5040 9356 5080 9724
rect 5040 9324 5044 9356
rect 5076 9324 5080 9356
rect 5040 9276 5080 9324
rect 5040 9244 5044 9276
rect 5076 9244 5080 9276
rect 5040 9196 5080 9244
rect 5040 9164 5044 9196
rect 5076 9164 5080 9196
rect 5040 8876 5080 9164
rect 5040 8844 5044 8876
rect 5076 8844 5080 8876
rect 5040 8796 5080 8844
rect 5040 8764 5044 8796
rect 5076 8764 5080 8796
rect 5040 8716 5080 8764
rect 5040 8684 5044 8716
rect 5076 8684 5080 8716
rect 5040 8636 5080 8684
rect 5040 8604 5044 8636
rect 5076 8604 5080 8636
rect 5040 8556 5080 8604
rect 5040 8524 5044 8556
rect 5076 8524 5080 8556
rect 5040 8475 5080 8524
rect 5040 8445 5045 8475
rect 5075 8445 5080 8475
rect 5040 8315 5080 8445
rect 5040 8285 5045 8315
rect 5075 8285 5080 8315
rect 5040 8075 5080 8285
rect 5040 8045 5045 8075
rect 5075 8045 5080 8075
rect 5040 7755 5080 8045
rect 5040 7725 5045 7755
rect 5075 7725 5080 7755
rect 5040 7636 5080 7725
rect 5040 7604 5044 7636
rect 5076 7604 5080 7636
rect 5040 7556 5080 7604
rect 5040 7524 5044 7556
rect 5076 7524 5080 7556
rect 5040 7476 5080 7524
rect 5040 7444 5044 7476
rect 5076 7444 5080 7476
rect 5040 7396 5080 7444
rect 5040 7364 5044 7396
rect 5076 7364 5080 7396
rect 5040 7316 5080 7364
rect 5040 7284 5044 7316
rect 5076 7284 5080 7316
rect 5040 7236 5080 7284
rect 5040 7204 5044 7236
rect 5076 7204 5080 7236
rect 5040 7156 5080 7204
rect 5040 7124 5044 7156
rect 5076 7124 5080 7156
rect 5040 7076 5080 7124
rect 5040 7044 5044 7076
rect 5076 7044 5080 7076
rect 5040 6756 5080 7044
rect 5040 6724 5044 6756
rect 5076 6724 5080 6756
rect 5040 6676 5080 6724
rect 5040 6644 5044 6676
rect 5076 6644 5080 6676
rect 5040 6596 5080 6644
rect 5040 6564 5044 6596
rect 5076 6564 5080 6596
rect 5040 6516 5080 6564
rect 5040 6484 5044 6516
rect 5076 6484 5080 6516
rect 5040 6436 5080 6484
rect 5040 6404 5044 6436
rect 5076 6404 5080 6436
rect 5040 6356 5080 6404
rect 5040 6324 5044 6356
rect 5076 6324 5080 6356
rect 5040 6235 5080 6324
rect 5040 6205 5045 6235
rect 5075 6205 5080 6235
rect 5040 6075 5080 6205
rect 5040 6045 5045 6075
rect 5075 6045 5080 6075
rect 5040 5915 5080 6045
rect 5040 5885 5045 5915
rect 5075 5885 5080 5915
rect 5040 5796 5080 5885
rect 5040 5764 5044 5796
rect 5076 5764 5080 5796
rect 5040 5716 5080 5764
rect 5040 5684 5044 5716
rect 5076 5684 5080 5716
rect 5040 5636 5080 5684
rect 5040 5604 5044 5636
rect 5076 5604 5080 5636
rect 5040 5556 5080 5604
rect 5040 5524 5044 5556
rect 5076 5524 5080 5556
rect 5040 5476 5080 5524
rect 5040 5444 5044 5476
rect 5076 5444 5080 5476
rect 5040 5396 5080 5444
rect 5040 5364 5044 5396
rect 5076 5364 5080 5396
rect 5040 5316 5080 5364
rect 5040 5284 5044 5316
rect 5076 5284 5080 5316
rect 5040 5236 5080 5284
rect 5040 5204 5044 5236
rect 5076 5204 5080 5236
rect 5040 5156 5080 5204
rect 5040 5124 5044 5156
rect 5076 5124 5080 5156
rect 5040 5076 5080 5124
rect 5040 5044 5044 5076
rect 5076 5044 5080 5076
rect 5040 4996 5080 5044
rect 5040 4964 5044 4996
rect 5076 4964 5080 4996
rect 5040 4436 5080 4964
rect 5040 4404 5044 4436
rect 5076 4404 5080 4436
rect 5040 4356 5080 4404
rect 5040 4324 5044 4356
rect 5076 4324 5080 4356
rect 5040 4276 5080 4324
rect 5040 4244 5044 4276
rect 5076 4244 5080 4276
rect 5040 4196 5080 4244
rect 5040 4164 5044 4196
rect 5076 4164 5080 4196
rect 5040 4116 5080 4164
rect 5040 4084 5044 4116
rect 5076 4084 5080 4116
rect 5040 4036 5080 4084
rect 5040 4004 5044 4036
rect 5076 4004 5080 4036
rect 5040 3956 5080 4004
rect 5040 3924 5044 3956
rect 5076 3924 5080 3956
rect 5040 3156 5080 3924
rect 5040 3124 5044 3156
rect 5076 3124 5080 3156
rect 5040 3076 5080 3124
rect 5040 3044 5044 3076
rect 5076 3044 5080 3076
rect 5040 2996 5080 3044
rect 5040 2964 5044 2996
rect 5076 2964 5080 2996
rect 5040 2916 5080 2964
rect 5040 2884 5044 2916
rect 5076 2884 5080 2916
rect 5040 2836 5080 2884
rect 5040 2804 5044 2836
rect 5076 2804 5080 2836
rect 5040 2756 5080 2804
rect 5040 2724 5044 2756
rect 5076 2724 5080 2756
rect 5040 2676 5080 2724
rect 5040 2644 5044 2676
rect 5076 2644 5080 2676
rect 5040 2596 5080 2644
rect 5040 2564 5044 2596
rect 5076 2564 5080 2596
rect 5040 2516 5080 2564
rect 5040 2484 5044 2516
rect 5076 2484 5080 2516
rect 5040 2436 5080 2484
rect 5040 2404 5044 2436
rect 5076 2404 5080 2436
rect 5040 2356 5080 2404
rect 5040 2324 5044 2356
rect 5076 2324 5080 2356
rect 5040 2276 5080 2324
rect 5040 2244 5044 2276
rect 5076 2244 5080 2276
rect 5040 2196 5080 2244
rect 5040 2164 5044 2196
rect 5076 2164 5080 2196
rect 5040 2116 5080 2164
rect 5040 2084 5044 2116
rect 5076 2084 5080 2116
rect 5040 2036 5080 2084
rect 5040 2004 5044 2036
rect 5076 2004 5080 2036
rect 5040 1636 5080 2004
rect 5040 1604 5044 1636
rect 5076 1604 5080 1636
rect 5040 1556 5080 1604
rect 5040 1524 5044 1556
rect 5076 1524 5080 1556
rect 5040 1476 5080 1524
rect 5040 1444 5044 1476
rect 5076 1444 5080 1476
rect 5040 1396 5080 1444
rect 5040 1364 5044 1396
rect 5076 1364 5080 1396
rect 5040 1316 5080 1364
rect 5040 1284 5044 1316
rect 5076 1284 5080 1316
rect 5040 1236 5080 1284
rect 5040 1204 5044 1236
rect 5076 1204 5080 1236
rect 5040 1156 5080 1204
rect 5040 1124 5044 1156
rect 5076 1124 5080 1156
rect 5040 1076 5080 1124
rect 5040 1044 5044 1076
rect 5076 1044 5080 1076
rect 5040 756 5080 1044
rect 5040 724 5044 756
rect 5076 724 5080 756
rect 5040 676 5080 724
rect 5040 644 5044 676
rect 5076 644 5080 676
rect 5040 596 5080 644
rect 5040 564 5044 596
rect 5076 564 5080 596
rect 5040 196 5080 564
rect 5040 164 5044 196
rect 5076 164 5080 196
rect 5040 116 5080 164
rect 5040 84 5044 116
rect 5076 84 5080 116
rect 5040 36 5080 84
rect 5040 4 5044 36
rect 5076 4 5080 36
rect 5040 -40 5080 4
rect 5120 15396 5160 15400
rect 5120 15364 5124 15396
rect 5156 15364 5160 15396
rect 5120 14116 5160 15364
rect 5120 14084 5124 14116
rect 5156 14084 5160 14116
rect 5120 12636 5160 14084
rect 5120 12604 5124 12636
rect 5156 12604 5160 12636
rect 5120 12556 5160 12604
rect 5120 12524 5124 12556
rect 5156 12524 5160 12556
rect 5120 12476 5160 12524
rect 5120 12444 5124 12476
rect 5156 12444 5160 12476
rect 5120 12396 5160 12444
rect 5120 12364 5124 12396
rect 5156 12364 5160 12396
rect 5120 12316 5160 12364
rect 5120 12284 5124 12316
rect 5156 12284 5160 12316
rect 5120 12236 5160 12284
rect 5120 12204 5124 12236
rect 5156 12204 5160 12236
rect 5120 12156 5160 12204
rect 5120 12124 5124 12156
rect 5156 12124 5160 12156
rect 5120 11836 5160 12124
rect 5120 11804 5124 11836
rect 5156 11804 5160 11836
rect 5120 11756 5160 11804
rect 5120 11724 5124 11756
rect 5156 11724 5160 11756
rect 5120 11676 5160 11724
rect 5120 11644 5124 11676
rect 5156 11644 5160 11676
rect 5120 11596 5160 11644
rect 5120 11564 5124 11596
rect 5156 11564 5160 11596
rect 5120 11516 5160 11564
rect 5120 11484 5124 11516
rect 5156 11484 5160 11516
rect 5120 11436 5160 11484
rect 5120 11404 5124 11436
rect 5156 11404 5160 11436
rect 5120 11075 5160 11404
rect 5120 11045 5125 11075
rect 5155 11045 5160 11075
rect 5120 10876 5160 11045
rect 5120 10844 5124 10876
rect 5156 10844 5160 10876
rect 5120 10796 5160 10844
rect 5120 10764 5124 10796
rect 5156 10764 5160 10796
rect 5120 10716 5160 10764
rect 5120 10684 5124 10716
rect 5156 10684 5160 10716
rect 5120 10636 5160 10684
rect 5120 10604 5124 10636
rect 5156 10604 5160 10636
rect 5120 10556 5160 10604
rect 5120 10524 5124 10556
rect 5156 10524 5160 10556
rect 5120 10476 5160 10524
rect 5120 10444 5124 10476
rect 5156 10444 5160 10476
rect 5120 10396 5160 10444
rect 5120 10364 5124 10396
rect 5156 10364 5160 10396
rect 5120 10316 5160 10364
rect 5120 10284 5124 10316
rect 5156 10284 5160 10316
rect 5120 10236 5160 10284
rect 5120 10204 5124 10236
rect 5156 10204 5160 10236
rect 5120 10156 5160 10204
rect 5120 10124 5124 10156
rect 5156 10124 5160 10156
rect 5120 10076 5160 10124
rect 5120 10044 5124 10076
rect 5156 10044 5160 10076
rect 5120 9996 5160 10044
rect 5120 9964 5124 9996
rect 5156 9964 5160 9996
rect 5120 9916 5160 9964
rect 5120 9884 5124 9916
rect 5156 9884 5160 9916
rect 5120 9836 5160 9884
rect 5120 9804 5124 9836
rect 5156 9804 5160 9836
rect 5120 9756 5160 9804
rect 5120 9724 5124 9756
rect 5156 9724 5160 9756
rect 5120 9356 5160 9724
rect 5120 9324 5124 9356
rect 5156 9324 5160 9356
rect 5120 9276 5160 9324
rect 5120 9244 5124 9276
rect 5156 9244 5160 9276
rect 5120 9196 5160 9244
rect 5120 9164 5124 9196
rect 5156 9164 5160 9196
rect 5120 9115 5160 9164
rect 5120 9085 5125 9115
rect 5155 9085 5160 9115
rect 5120 8955 5160 9085
rect 5120 8925 5125 8955
rect 5155 8925 5160 8955
rect 5120 8876 5160 8925
rect 5120 8844 5124 8876
rect 5156 8844 5160 8876
rect 5120 8796 5160 8844
rect 5120 8764 5124 8796
rect 5156 8764 5160 8796
rect 5120 8716 5160 8764
rect 5120 8684 5124 8716
rect 5156 8684 5160 8716
rect 5120 8636 5160 8684
rect 5120 8604 5124 8636
rect 5156 8604 5160 8636
rect 5120 8556 5160 8604
rect 5120 8524 5124 8556
rect 5156 8524 5160 8556
rect 5120 7995 5160 8524
rect 5120 7965 5125 7995
rect 5155 7965 5160 7995
rect 5120 7835 5160 7965
rect 5120 7805 5125 7835
rect 5155 7805 5160 7835
rect 5120 7636 5160 7805
rect 5120 7604 5124 7636
rect 5156 7604 5160 7636
rect 5120 7556 5160 7604
rect 5120 7524 5124 7556
rect 5156 7524 5160 7556
rect 5120 7476 5160 7524
rect 5120 7444 5124 7476
rect 5156 7444 5160 7476
rect 5120 7396 5160 7444
rect 5120 7364 5124 7396
rect 5156 7364 5160 7396
rect 5120 7316 5160 7364
rect 5120 7284 5124 7316
rect 5156 7284 5160 7316
rect 5120 7236 5160 7284
rect 5120 7204 5124 7236
rect 5156 7204 5160 7236
rect 5120 7156 5160 7204
rect 5120 7124 5124 7156
rect 5156 7124 5160 7156
rect 5120 7076 5160 7124
rect 5120 7044 5124 7076
rect 5156 7044 5160 7076
rect 5120 6756 5160 7044
rect 5120 6724 5124 6756
rect 5156 6724 5160 6756
rect 5120 6676 5160 6724
rect 5120 6644 5124 6676
rect 5156 6644 5160 6676
rect 5120 6596 5160 6644
rect 5120 6564 5124 6596
rect 5156 6564 5160 6596
rect 5120 6516 5160 6564
rect 5120 6484 5124 6516
rect 5156 6484 5160 6516
rect 5120 6436 5160 6484
rect 5120 6404 5124 6436
rect 5156 6404 5160 6436
rect 5120 6356 5160 6404
rect 5120 6324 5124 6356
rect 5156 6324 5160 6356
rect 5120 5796 5160 6324
rect 5120 5764 5124 5796
rect 5156 5764 5160 5796
rect 5120 5716 5160 5764
rect 5120 5684 5124 5716
rect 5156 5684 5160 5716
rect 5120 5636 5160 5684
rect 5120 5604 5124 5636
rect 5156 5604 5160 5636
rect 5120 5556 5160 5604
rect 5120 5524 5124 5556
rect 5156 5524 5160 5556
rect 5120 5476 5160 5524
rect 5120 5444 5124 5476
rect 5156 5444 5160 5476
rect 5120 5396 5160 5444
rect 5120 5364 5124 5396
rect 5156 5364 5160 5396
rect 5120 5316 5160 5364
rect 5120 5284 5124 5316
rect 5156 5284 5160 5316
rect 5120 5236 5160 5284
rect 5120 5204 5124 5236
rect 5156 5204 5160 5236
rect 5120 5156 5160 5204
rect 5120 5124 5124 5156
rect 5156 5124 5160 5156
rect 5120 5076 5160 5124
rect 5120 5044 5124 5076
rect 5156 5044 5160 5076
rect 5120 4996 5160 5044
rect 5120 4964 5124 4996
rect 5156 4964 5160 4996
rect 5120 4436 5160 4964
rect 5120 4404 5124 4436
rect 5156 4404 5160 4436
rect 5120 4356 5160 4404
rect 5120 4324 5124 4356
rect 5156 4324 5160 4356
rect 5120 4276 5160 4324
rect 5120 4244 5124 4276
rect 5156 4244 5160 4276
rect 5120 4196 5160 4244
rect 5120 4164 5124 4196
rect 5156 4164 5160 4196
rect 5120 4116 5160 4164
rect 5120 4084 5124 4116
rect 5156 4084 5160 4116
rect 5120 4036 5160 4084
rect 5120 4004 5124 4036
rect 5156 4004 5160 4036
rect 5120 3956 5160 4004
rect 5120 3924 5124 3956
rect 5156 3924 5160 3956
rect 5120 3156 5160 3924
rect 5120 3124 5124 3156
rect 5156 3124 5160 3156
rect 5120 3076 5160 3124
rect 5120 3044 5124 3076
rect 5156 3044 5160 3076
rect 5120 2996 5160 3044
rect 5120 2964 5124 2996
rect 5156 2964 5160 2996
rect 5120 2916 5160 2964
rect 5120 2884 5124 2916
rect 5156 2884 5160 2916
rect 5120 2836 5160 2884
rect 5120 2804 5124 2836
rect 5156 2804 5160 2836
rect 5120 2756 5160 2804
rect 5120 2724 5124 2756
rect 5156 2724 5160 2756
rect 5120 2676 5160 2724
rect 5120 2644 5124 2676
rect 5156 2644 5160 2676
rect 5120 2596 5160 2644
rect 5120 2564 5124 2596
rect 5156 2564 5160 2596
rect 5120 2516 5160 2564
rect 5120 2484 5124 2516
rect 5156 2484 5160 2516
rect 5120 2436 5160 2484
rect 5120 2404 5124 2436
rect 5156 2404 5160 2436
rect 5120 2356 5160 2404
rect 5120 2324 5124 2356
rect 5156 2324 5160 2356
rect 5120 2276 5160 2324
rect 5120 2244 5124 2276
rect 5156 2244 5160 2276
rect 5120 2196 5160 2244
rect 5120 2164 5124 2196
rect 5156 2164 5160 2196
rect 5120 2116 5160 2164
rect 5120 2084 5124 2116
rect 5156 2084 5160 2116
rect 5120 2036 5160 2084
rect 5120 2004 5124 2036
rect 5156 2004 5160 2036
rect 5120 1636 5160 2004
rect 5120 1604 5124 1636
rect 5156 1604 5160 1636
rect 5120 1556 5160 1604
rect 5120 1524 5124 1556
rect 5156 1524 5160 1556
rect 5120 1476 5160 1524
rect 5120 1444 5124 1476
rect 5156 1444 5160 1476
rect 5120 1396 5160 1444
rect 5120 1364 5124 1396
rect 5156 1364 5160 1396
rect 5120 1316 5160 1364
rect 5120 1284 5124 1316
rect 5156 1284 5160 1316
rect 5120 1236 5160 1284
rect 5120 1204 5124 1236
rect 5156 1204 5160 1236
rect 5120 1156 5160 1204
rect 5120 1124 5124 1156
rect 5156 1124 5160 1156
rect 5120 1076 5160 1124
rect 5120 1044 5124 1076
rect 5156 1044 5160 1076
rect 5120 756 5160 1044
rect 5120 724 5124 756
rect 5156 724 5160 756
rect 5120 676 5160 724
rect 5120 644 5124 676
rect 5156 644 5160 676
rect 5120 596 5160 644
rect 5120 564 5124 596
rect 5156 564 5160 596
rect 5120 196 5160 564
rect 5120 164 5124 196
rect 5156 164 5160 196
rect 5120 116 5160 164
rect 5120 84 5124 116
rect 5156 84 5160 116
rect 5120 36 5160 84
rect 5120 4 5124 36
rect 5156 4 5160 36
rect 5120 -40 5160 4
rect 5200 15316 5240 15400
rect 5200 15284 5204 15316
rect 5236 15284 5240 15316
rect 5200 7915 5240 15284
rect 5200 7885 5205 7915
rect 5235 7885 5240 7915
rect 5200 -40 5240 7885
rect 5280 15396 5320 15400
rect 5280 15364 5284 15396
rect 5316 15364 5320 15396
rect 5280 14116 5320 15364
rect 5280 14084 5284 14116
rect 5316 14084 5320 14116
rect 5280 12636 5320 14084
rect 5280 12604 5284 12636
rect 5316 12604 5320 12636
rect 5280 12556 5320 12604
rect 5280 12524 5284 12556
rect 5316 12524 5320 12556
rect 5280 12476 5320 12524
rect 5280 12444 5284 12476
rect 5316 12444 5320 12476
rect 5280 12396 5320 12444
rect 5280 12364 5284 12396
rect 5316 12364 5320 12396
rect 5280 12316 5320 12364
rect 5280 12284 5284 12316
rect 5316 12284 5320 12316
rect 5280 12236 5320 12284
rect 5280 12204 5284 12236
rect 5316 12204 5320 12236
rect 5280 12156 5320 12204
rect 5280 12124 5284 12156
rect 5316 12124 5320 12156
rect 5280 11836 5320 12124
rect 5280 11804 5284 11836
rect 5316 11804 5320 11836
rect 5280 11756 5320 11804
rect 5280 11724 5284 11756
rect 5316 11724 5320 11756
rect 5280 11676 5320 11724
rect 5280 11644 5284 11676
rect 5316 11644 5320 11676
rect 5280 11596 5320 11644
rect 5280 11564 5284 11596
rect 5316 11564 5320 11596
rect 5280 11516 5320 11564
rect 5280 11484 5284 11516
rect 5316 11484 5320 11516
rect 5280 11436 5320 11484
rect 5280 11404 5284 11436
rect 5316 11404 5320 11436
rect 5280 11075 5320 11404
rect 5280 11045 5285 11075
rect 5315 11045 5320 11075
rect 5280 10876 5320 11045
rect 5280 10844 5284 10876
rect 5316 10844 5320 10876
rect 5280 10796 5320 10844
rect 5280 10764 5284 10796
rect 5316 10764 5320 10796
rect 5280 10716 5320 10764
rect 5280 10684 5284 10716
rect 5316 10684 5320 10716
rect 5280 10636 5320 10684
rect 5280 10604 5284 10636
rect 5316 10604 5320 10636
rect 5280 10556 5320 10604
rect 5280 10524 5284 10556
rect 5316 10524 5320 10556
rect 5280 10476 5320 10524
rect 5280 10444 5284 10476
rect 5316 10444 5320 10476
rect 5280 10396 5320 10444
rect 5280 10364 5284 10396
rect 5316 10364 5320 10396
rect 5280 10316 5320 10364
rect 5280 10284 5284 10316
rect 5316 10284 5320 10316
rect 5280 10236 5320 10284
rect 5280 10204 5284 10236
rect 5316 10204 5320 10236
rect 5280 10156 5320 10204
rect 5280 10124 5284 10156
rect 5316 10124 5320 10156
rect 5280 10076 5320 10124
rect 5280 10044 5284 10076
rect 5316 10044 5320 10076
rect 5280 9996 5320 10044
rect 5280 9964 5284 9996
rect 5316 9964 5320 9996
rect 5280 9916 5320 9964
rect 5280 9884 5284 9916
rect 5316 9884 5320 9916
rect 5280 9836 5320 9884
rect 5280 9804 5284 9836
rect 5316 9804 5320 9836
rect 5280 9756 5320 9804
rect 5280 9724 5284 9756
rect 5316 9724 5320 9756
rect 5280 9356 5320 9724
rect 5280 9324 5284 9356
rect 5316 9324 5320 9356
rect 5280 9276 5320 9324
rect 5280 9244 5284 9276
rect 5316 9244 5320 9276
rect 5280 9196 5320 9244
rect 5280 9164 5284 9196
rect 5316 9164 5320 9196
rect 5280 9115 5320 9164
rect 5280 9085 5285 9115
rect 5315 9085 5320 9115
rect 5280 8955 5320 9085
rect 5280 8925 5285 8955
rect 5315 8925 5320 8955
rect 5280 8876 5320 8925
rect 5280 8844 5284 8876
rect 5316 8844 5320 8876
rect 5280 8796 5320 8844
rect 5280 8764 5284 8796
rect 5316 8764 5320 8796
rect 5280 8716 5320 8764
rect 5280 8684 5284 8716
rect 5316 8684 5320 8716
rect 5280 8636 5320 8684
rect 5280 8604 5284 8636
rect 5316 8604 5320 8636
rect 5280 8556 5320 8604
rect 5280 8524 5284 8556
rect 5316 8524 5320 8556
rect 5280 7995 5320 8524
rect 5280 7965 5285 7995
rect 5315 7965 5320 7995
rect 5280 7835 5320 7965
rect 5280 7805 5285 7835
rect 5315 7805 5320 7835
rect 5280 7636 5320 7805
rect 5280 7604 5284 7636
rect 5316 7604 5320 7636
rect 5280 7556 5320 7604
rect 5280 7524 5284 7556
rect 5316 7524 5320 7556
rect 5280 7476 5320 7524
rect 5280 7444 5284 7476
rect 5316 7444 5320 7476
rect 5280 7396 5320 7444
rect 5280 7364 5284 7396
rect 5316 7364 5320 7396
rect 5280 7316 5320 7364
rect 5280 7284 5284 7316
rect 5316 7284 5320 7316
rect 5280 7236 5320 7284
rect 5280 7204 5284 7236
rect 5316 7204 5320 7236
rect 5280 7156 5320 7204
rect 5280 7124 5284 7156
rect 5316 7124 5320 7156
rect 5280 7076 5320 7124
rect 5280 7044 5284 7076
rect 5316 7044 5320 7076
rect 5280 6756 5320 7044
rect 5280 6724 5284 6756
rect 5316 6724 5320 6756
rect 5280 6676 5320 6724
rect 5280 6644 5284 6676
rect 5316 6644 5320 6676
rect 5280 6596 5320 6644
rect 5280 6564 5284 6596
rect 5316 6564 5320 6596
rect 5280 6516 5320 6564
rect 5280 6484 5284 6516
rect 5316 6484 5320 6516
rect 5280 6436 5320 6484
rect 5280 6404 5284 6436
rect 5316 6404 5320 6436
rect 5280 6356 5320 6404
rect 5280 6324 5284 6356
rect 5316 6324 5320 6356
rect 5280 5796 5320 6324
rect 5280 5764 5284 5796
rect 5316 5764 5320 5796
rect 5280 5716 5320 5764
rect 5280 5684 5284 5716
rect 5316 5684 5320 5716
rect 5280 5636 5320 5684
rect 5280 5604 5284 5636
rect 5316 5604 5320 5636
rect 5280 5556 5320 5604
rect 5280 5524 5284 5556
rect 5316 5524 5320 5556
rect 5280 5476 5320 5524
rect 5280 5444 5284 5476
rect 5316 5444 5320 5476
rect 5280 5396 5320 5444
rect 5280 5364 5284 5396
rect 5316 5364 5320 5396
rect 5280 5316 5320 5364
rect 5280 5284 5284 5316
rect 5316 5284 5320 5316
rect 5280 5236 5320 5284
rect 5280 5204 5284 5236
rect 5316 5204 5320 5236
rect 5280 5156 5320 5204
rect 5280 5124 5284 5156
rect 5316 5124 5320 5156
rect 5280 5076 5320 5124
rect 5280 5044 5284 5076
rect 5316 5044 5320 5076
rect 5280 4996 5320 5044
rect 5280 4964 5284 4996
rect 5316 4964 5320 4996
rect 5280 4436 5320 4964
rect 5280 4404 5284 4436
rect 5316 4404 5320 4436
rect 5280 4356 5320 4404
rect 5280 4324 5284 4356
rect 5316 4324 5320 4356
rect 5280 4276 5320 4324
rect 5280 4244 5284 4276
rect 5316 4244 5320 4276
rect 5280 4196 5320 4244
rect 5280 4164 5284 4196
rect 5316 4164 5320 4196
rect 5280 4116 5320 4164
rect 5280 4084 5284 4116
rect 5316 4084 5320 4116
rect 5280 4036 5320 4084
rect 5280 4004 5284 4036
rect 5316 4004 5320 4036
rect 5280 3956 5320 4004
rect 5280 3924 5284 3956
rect 5316 3924 5320 3956
rect 5280 3156 5320 3924
rect 5280 3124 5284 3156
rect 5316 3124 5320 3156
rect 5280 3076 5320 3124
rect 5280 3044 5284 3076
rect 5316 3044 5320 3076
rect 5280 2996 5320 3044
rect 5280 2964 5284 2996
rect 5316 2964 5320 2996
rect 5280 2916 5320 2964
rect 5280 2884 5284 2916
rect 5316 2884 5320 2916
rect 5280 2836 5320 2884
rect 5280 2804 5284 2836
rect 5316 2804 5320 2836
rect 5280 2756 5320 2804
rect 5280 2724 5284 2756
rect 5316 2724 5320 2756
rect 5280 2676 5320 2724
rect 5280 2644 5284 2676
rect 5316 2644 5320 2676
rect 5280 2596 5320 2644
rect 5280 2564 5284 2596
rect 5316 2564 5320 2596
rect 5280 2516 5320 2564
rect 5280 2484 5284 2516
rect 5316 2484 5320 2516
rect 5280 2436 5320 2484
rect 5280 2404 5284 2436
rect 5316 2404 5320 2436
rect 5280 2356 5320 2404
rect 5280 2324 5284 2356
rect 5316 2324 5320 2356
rect 5280 2276 5320 2324
rect 5280 2244 5284 2276
rect 5316 2244 5320 2276
rect 5280 2196 5320 2244
rect 5280 2164 5284 2196
rect 5316 2164 5320 2196
rect 5280 2116 5320 2164
rect 5280 2084 5284 2116
rect 5316 2084 5320 2116
rect 5280 2036 5320 2084
rect 5280 2004 5284 2036
rect 5316 2004 5320 2036
rect 5280 1636 5320 2004
rect 5280 1604 5284 1636
rect 5316 1604 5320 1636
rect 5280 1556 5320 1604
rect 5280 1524 5284 1556
rect 5316 1524 5320 1556
rect 5280 1476 5320 1524
rect 5280 1444 5284 1476
rect 5316 1444 5320 1476
rect 5280 1396 5320 1444
rect 5280 1364 5284 1396
rect 5316 1364 5320 1396
rect 5280 1316 5320 1364
rect 5280 1284 5284 1316
rect 5316 1284 5320 1316
rect 5280 1236 5320 1284
rect 5280 1204 5284 1236
rect 5316 1204 5320 1236
rect 5280 1156 5320 1204
rect 5280 1124 5284 1156
rect 5316 1124 5320 1156
rect 5280 1076 5320 1124
rect 5280 1044 5284 1076
rect 5316 1044 5320 1076
rect 5280 756 5320 1044
rect 5280 724 5284 756
rect 5316 724 5320 756
rect 5280 676 5320 724
rect 5280 644 5284 676
rect 5316 644 5320 676
rect 5280 596 5320 644
rect 5280 564 5284 596
rect 5316 564 5320 596
rect 5280 196 5320 564
rect 5280 164 5284 196
rect 5316 164 5320 196
rect 5280 116 5320 164
rect 5280 84 5284 116
rect 5316 84 5320 116
rect 5280 36 5320 84
rect 5280 4 5284 36
rect 5316 4 5320 36
rect 5280 -40 5320 4
rect 5360 15316 5400 15400
rect 5360 15284 5364 15316
rect 5396 15284 5400 15316
rect 5360 9035 5400 15284
rect 5360 9005 5365 9035
rect 5395 9005 5400 9035
rect 5360 -40 5400 9005
rect 5440 15396 5480 15400
rect 5440 15364 5444 15396
rect 5476 15364 5480 15396
rect 5440 14116 5480 15364
rect 5440 14084 5444 14116
rect 5476 14084 5480 14116
rect 5440 12636 5480 14084
rect 5440 12604 5444 12636
rect 5476 12604 5480 12636
rect 5440 12556 5480 12604
rect 5440 12524 5444 12556
rect 5476 12524 5480 12556
rect 5440 12476 5480 12524
rect 5440 12444 5444 12476
rect 5476 12444 5480 12476
rect 5440 12396 5480 12444
rect 5440 12364 5444 12396
rect 5476 12364 5480 12396
rect 5440 12316 5480 12364
rect 5440 12284 5444 12316
rect 5476 12284 5480 12316
rect 5440 12236 5480 12284
rect 5440 12204 5444 12236
rect 5476 12204 5480 12236
rect 5440 12156 5480 12204
rect 5440 12124 5444 12156
rect 5476 12124 5480 12156
rect 5440 11836 5480 12124
rect 5440 11804 5444 11836
rect 5476 11804 5480 11836
rect 5440 11756 5480 11804
rect 5440 11724 5444 11756
rect 5476 11724 5480 11756
rect 5440 11676 5480 11724
rect 5440 11644 5444 11676
rect 5476 11644 5480 11676
rect 5440 11596 5480 11644
rect 5440 11564 5444 11596
rect 5476 11564 5480 11596
rect 5440 11516 5480 11564
rect 5440 11484 5444 11516
rect 5476 11484 5480 11516
rect 5440 11436 5480 11484
rect 5440 11404 5444 11436
rect 5476 11404 5480 11436
rect 5440 11075 5480 11404
rect 5440 11045 5445 11075
rect 5475 11045 5480 11075
rect 5440 10876 5480 11045
rect 5440 10844 5444 10876
rect 5476 10844 5480 10876
rect 5440 10796 5480 10844
rect 5440 10764 5444 10796
rect 5476 10764 5480 10796
rect 5440 10716 5480 10764
rect 5440 10684 5444 10716
rect 5476 10684 5480 10716
rect 5440 10636 5480 10684
rect 5440 10604 5444 10636
rect 5476 10604 5480 10636
rect 5440 10556 5480 10604
rect 5440 10524 5444 10556
rect 5476 10524 5480 10556
rect 5440 10476 5480 10524
rect 5440 10444 5444 10476
rect 5476 10444 5480 10476
rect 5440 10396 5480 10444
rect 5440 10364 5444 10396
rect 5476 10364 5480 10396
rect 5440 10316 5480 10364
rect 5440 10284 5444 10316
rect 5476 10284 5480 10316
rect 5440 10236 5480 10284
rect 5440 10204 5444 10236
rect 5476 10204 5480 10236
rect 5440 10156 5480 10204
rect 5440 10124 5444 10156
rect 5476 10124 5480 10156
rect 5440 10076 5480 10124
rect 5440 10044 5444 10076
rect 5476 10044 5480 10076
rect 5440 9996 5480 10044
rect 5440 9964 5444 9996
rect 5476 9964 5480 9996
rect 5440 9916 5480 9964
rect 5440 9884 5444 9916
rect 5476 9884 5480 9916
rect 5440 9836 5480 9884
rect 5440 9804 5444 9836
rect 5476 9804 5480 9836
rect 5440 9756 5480 9804
rect 5440 9724 5444 9756
rect 5476 9724 5480 9756
rect 5440 9356 5480 9724
rect 5440 9324 5444 9356
rect 5476 9324 5480 9356
rect 5440 9276 5480 9324
rect 5440 9244 5444 9276
rect 5476 9244 5480 9276
rect 5440 9196 5480 9244
rect 5440 9164 5444 9196
rect 5476 9164 5480 9196
rect 5440 9115 5480 9164
rect 5440 9085 5445 9115
rect 5475 9085 5480 9115
rect 5440 8955 5480 9085
rect 5440 8925 5445 8955
rect 5475 8925 5480 8955
rect 5440 8876 5480 8925
rect 5440 8844 5444 8876
rect 5476 8844 5480 8876
rect 5440 8796 5480 8844
rect 5440 8764 5444 8796
rect 5476 8764 5480 8796
rect 5440 8716 5480 8764
rect 5440 8684 5444 8716
rect 5476 8684 5480 8716
rect 5440 8636 5480 8684
rect 5440 8604 5444 8636
rect 5476 8604 5480 8636
rect 5440 8556 5480 8604
rect 5440 8524 5444 8556
rect 5476 8524 5480 8556
rect 5440 7995 5480 8524
rect 5440 7965 5445 7995
rect 5475 7965 5480 7995
rect 5440 7835 5480 7965
rect 5440 7805 5445 7835
rect 5475 7805 5480 7835
rect 5440 7636 5480 7805
rect 5440 7604 5444 7636
rect 5476 7604 5480 7636
rect 5440 7556 5480 7604
rect 5440 7524 5444 7556
rect 5476 7524 5480 7556
rect 5440 7476 5480 7524
rect 5440 7444 5444 7476
rect 5476 7444 5480 7476
rect 5440 7396 5480 7444
rect 5440 7364 5444 7396
rect 5476 7364 5480 7396
rect 5440 7316 5480 7364
rect 5440 7284 5444 7316
rect 5476 7284 5480 7316
rect 5440 7236 5480 7284
rect 5440 7204 5444 7236
rect 5476 7204 5480 7236
rect 5440 7156 5480 7204
rect 5440 7124 5444 7156
rect 5476 7124 5480 7156
rect 5440 7076 5480 7124
rect 5440 7044 5444 7076
rect 5476 7044 5480 7076
rect 5440 6756 5480 7044
rect 5440 6724 5444 6756
rect 5476 6724 5480 6756
rect 5440 6676 5480 6724
rect 5440 6644 5444 6676
rect 5476 6644 5480 6676
rect 5440 6596 5480 6644
rect 5440 6564 5444 6596
rect 5476 6564 5480 6596
rect 5440 6516 5480 6564
rect 5440 6484 5444 6516
rect 5476 6484 5480 6516
rect 5440 6436 5480 6484
rect 5440 6404 5444 6436
rect 5476 6404 5480 6436
rect 5440 6356 5480 6404
rect 5440 6324 5444 6356
rect 5476 6324 5480 6356
rect 5440 5796 5480 6324
rect 5440 5764 5444 5796
rect 5476 5764 5480 5796
rect 5440 5716 5480 5764
rect 5440 5684 5444 5716
rect 5476 5684 5480 5716
rect 5440 5636 5480 5684
rect 5440 5604 5444 5636
rect 5476 5604 5480 5636
rect 5440 5556 5480 5604
rect 5440 5524 5444 5556
rect 5476 5524 5480 5556
rect 5440 5476 5480 5524
rect 5440 5444 5444 5476
rect 5476 5444 5480 5476
rect 5440 5396 5480 5444
rect 5440 5364 5444 5396
rect 5476 5364 5480 5396
rect 5440 5316 5480 5364
rect 5440 5284 5444 5316
rect 5476 5284 5480 5316
rect 5440 5236 5480 5284
rect 5440 5204 5444 5236
rect 5476 5204 5480 5236
rect 5440 5156 5480 5204
rect 5440 5124 5444 5156
rect 5476 5124 5480 5156
rect 5440 5076 5480 5124
rect 5440 5044 5444 5076
rect 5476 5044 5480 5076
rect 5440 4996 5480 5044
rect 5440 4964 5444 4996
rect 5476 4964 5480 4996
rect 5440 4436 5480 4964
rect 5440 4404 5444 4436
rect 5476 4404 5480 4436
rect 5440 4356 5480 4404
rect 5440 4324 5444 4356
rect 5476 4324 5480 4356
rect 5440 4276 5480 4324
rect 5440 4244 5444 4276
rect 5476 4244 5480 4276
rect 5440 4196 5480 4244
rect 5440 4164 5444 4196
rect 5476 4164 5480 4196
rect 5440 4116 5480 4164
rect 5440 4084 5444 4116
rect 5476 4084 5480 4116
rect 5440 4036 5480 4084
rect 5440 4004 5444 4036
rect 5476 4004 5480 4036
rect 5440 3956 5480 4004
rect 5440 3924 5444 3956
rect 5476 3924 5480 3956
rect 5440 3156 5480 3924
rect 5440 3124 5444 3156
rect 5476 3124 5480 3156
rect 5440 3076 5480 3124
rect 5440 3044 5444 3076
rect 5476 3044 5480 3076
rect 5440 2996 5480 3044
rect 5440 2964 5444 2996
rect 5476 2964 5480 2996
rect 5440 2916 5480 2964
rect 5440 2884 5444 2916
rect 5476 2884 5480 2916
rect 5440 2836 5480 2884
rect 5440 2804 5444 2836
rect 5476 2804 5480 2836
rect 5440 2756 5480 2804
rect 5440 2724 5444 2756
rect 5476 2724 5480 2756
rect 5440 2676 5480 2724
rect 5440 2644 5444 2676
rect 5476 2644 5480 2676
rect 5440 2596 5480 2644
rect 5440 2564 5444 2596
rect 5476 2564 5480 2596
rect 5440 2516 5480 2564
rect 5440 2484 5444 2516
rect 5476 2484 5480 2516
rect 5440 2436 5480 2484
rect 5440 2404 5444 2436
rect 5476 2404 5480 2436
rect 5440 2356 5480 2404
rect 5440 2324 5444 2356
rect 5476 2324 5480 2356
rect 5440 2276 5480 2324
rect 5440 2244 5444 2276
rect 5476 2244 5480 2276
rect 5440 2196 5480 2244
rect 5440 2164 5444 2196
rect 5476 2164 5480 2196
rect 5440 2116 5480 2164
rect 5440 2084 5444 2116
rect 5476 2084 5480 2116
rect 5440 2036 5480 2084
rect 5440 2004 5444 2036
rect 5476 2004 5480 2036
rect 5440 1636 5480 2004
rect 5440 1604 5444 1636
rect 5476 1604 5480 1636
rect 5440 1556 5480 1604
rect 5440 1524 5444 1556
rect 5476 1524 5480 1556
rect 5440 1476 5480 1524
rect 5440 1444 5444 1476
rect 5476 1444 5480 1476
rect 5440 1396 5480 1444
rect 5440 1364 5444 1396
rect 5476 1364 5480 1396
rect 5440 1316 5480 1364
rect 5440 1284 5444 1316
rect 5476 1284 5480 1316
rect 5440 1236 5480 1284
rect 5440 1204 5444 1236
rect 5476 1204 5480 1236
rect 5440 1156 5480 1204
rect 5440 1124 5444 1156
rect 5476 1124 5480 1156
rect 5440 1076 5480 1124
rect 5440 1044 5444 1076
rect 5476 1044 5480 1076
rect 5440 756 5480 1044
rect 5440 724 5444 756
rect 5476 724 5480 756
rect 5440 676 5480 724
rect 5440 644 5444 676
rect 5476 644 5480 676
rect 5440 596 5480 644
rect 5440 564 5444 596
rect 5476 564 5480 596
rect 5440 196 5480 564
rect 5440 164 5444 196
rect 5476 164 5480 196
rect 5440 116 5480 164
rect 5440 84 5444 116
rect 5476 84 5480 116
rect 5440 36 5480 84
rect 5440 4 5444 36
rect 5476 4 5480 36
rect 5440 -40 5480 4
rect 5520 14036 5560 15400
rect 5600 15396 5640 15400
rect 5600 15364 5604 15396
rect 5636 15364 5640 15396
rect 5600 14116 5640 15364
rect 10160 15396 10200 15400
rect 10160 15364 10164 15396
rect 10196 15364 10200 15396
rect 5680 15316 5720 15320
rect 5680 15284 5684 15316
rect 5716 15284 5720 15316
rect 5680 15240 5720 15284
rect 6720 15316 6760 15320
rect 6720 15284 6724 15316
rect 6756 15284 6760 15316
rect 6720 15240 6760 15284
rect 5680 14160 6760 15240
rect 6800 15316 6840 15320
rect 6800 15284 6804 15316
rect 6836 15284 6840 15316
rect 6800 15240 6840 15284
rect 7840 15316 7880 15320
rect 7840 15284 7844 15316
rect 7876 15284 7880 15316
rect 7840 15240 7880 15284
rect 6800 14160 7880 15240
rect 7920 15316 7960 15320
rect 7920 15284 7924 15316
rect 7956 15284 7960 15316
rect 7920 15240 7960 15284
rect 8960 15316 9000 15320
rect 8960 15284 8964 15316
rect 8996 15284 9000 15316
rect 8960 15240 9000 15284
rect 7920 14160 9000 15240
rect 9040 15316 9080 15320
rect 9040 15284 9044 15316
rect 9076 15284 9080 15316
rect 9040 15240 9080 15284
rect 10080 15316 10120 15320
rect 10080 15284 10084 15316
rect 10116 15284 10120 15316
rect 10080 15240 10120 15284
rect 9040 14160 10120 15240
rect 5600 14084 5604 14116
rect 5636 14084 5640 14116
rect 5600 14080 5640 14084
rect 10160 14116 10200 15364
rect 10160 14084 10164 14116
rect 10196 14084 10200 14116
rect 10160 14080 10200 14084
rect 5520 14004 5524 14036
rect 5556 14004 5560 14036
rect 5520 13716 5560 14004
rect 5520 13684 5524 13716
rect 5556 13684 5560 13716
rect 5520 13396 5560 13684
rect 10240 14036 10280 15444
rect 10240 14004 10244 14036
rect 10276 14004 10280 14036
rect 10240 13716 10280 14004
rect 10320 16836 10360 16920
rect 10320 16804 10324 16836
rect 10356 16804 10360 16836
rect 10320 15556 10360 16804
rect 10320 15524 10324 15556
rect 10356 15524 10360 15556
rect 10320 13956 10360 15524
rect 10320 13924 10324 13956
rect 10356 13924 10360 13956
rect 10320 13796 10360 13924
rect 10320 13764 10324 13796
rect 10356 13764 10360 13796
rect 10320 13760 10360 13764
rect 10400 16756 10440 16920
rect 10400 16724 10404 16756
rect 10436 16724 10440 16756
rect 10400 13876 10440 16724
rect 10400 13844 10404 13876
rect 10436 13844 10440 13876
rect 10400 13760 10440 13844
rect 10480 16836 10520 16920
rect 10480 16804 10484 16836
rect 10516 16804 10520 16836
rect 10480 15556 10520 16804
rect 10480 15524 10484 15556
rect 10516 15524 10520 15556
rect 10480 13956 10520 15524
rect 10480 13924 10484 13956
rect 10516 13924 10520 13956
rect 10480 13796 10520 13924
rect 10480 13764 10484 13796
rect 10516 13764 10520 13796
rect 10480 13760 10520 13764
rect 10560 16916 10600 16920
rect 10560 16884 10564 16916
rect 10596 16884 10600 16916
rect 10560 15476 10600 16884
rect 10560 15444 10564 15476
rect 10596 15444 10600 15476
rect 10560 14036 10600 15444
rect 10560 14004 10564 14036
rect 10596 14004 10600 14036
rect 10240 13684 10244 13716
rect 10276 13684 10280 13716
rect 10240 13680 10280 13684
rect 10560 13716 10600 14004
rect 10560 13684 10564 13716
rect 10596 13684 10600 13716
rect 10560 13680 10600 13684
rect 5520 13204 5524 13396
rect 5556 13204 5560 13396
rect 5520 12636 5560 13204
rect 5680 13396 5720 13400
rect 5680 13204 5684 13396
rect 5716 13204 5720 13396
rect 5520 12604 5524 12636
rect 5556 12604 5560 12636
rect 5520 12556 5560 12604
rect 5520 12524 5524 12556
rect 5556 12524 5560 12556
rect 5520 12476 5560 12524
rect 5520 12444 5524 12476
rect 5556 12444 5560 12476
rect 5520 12396 5560 12444
rect 5520 12364 5524 12396
rect 5556 12364 5560 12396
rect 5520 12316 5560 12364
rect 5520 12284 5524 12316
rect 5556 12284 5560 12316
rect 5520 12236 5560 12284
rect 5520 12204 5524 12236
rect 5556 12204 5560 12236
rect 5520 12156 5560 12204
rect 5520 12124 5524 12156
rect 5556 12124 5560 12156
rect 5520 11836 5560 12124
rect 5520 11804 5524 11836
rect 5556 11804 5560 11836
rect 5520 11756 5560 11804
rect 5520 11724 5524 11756
rect 5556 11724 5560 11756
rect 5520 11676 5560 11724
rect 5520 11644 5524 11676
rect 5556 11644 5560 11676
rect 5520 11596 5560 11644
rect 5520 11564 5524 11596
rect 5556 11564 5560 11596
rect 5520 11516 5560 11564
rect 5520 11484 5524 11516
rect 5556 11484 5560 11516
rect 5520 11436 5560 11484
rect 5520 11404 5524 11436
rect 5556 11404 5560 11436
rect 5520 11315 5560 11404
rect 5520 11285 5525 11315
rect 5555 11285 5560 11315
rect 5520 11155 5560 11285
rect 5520 11125 5525 11155
rect 5555 11125 5560 11155
rect 5520 10995 5560 11125
rect 5520 10965 5525 10995
rect 5555 10965 5560 10995
rect 5520 10876 5560 10965
rect 5520 10844 5524 10876
rect 5556 10844 5560 10876
rect 5520 10796 5560 10844
rect 5520 10764 5524 10796
rect 5556 10764 5560 10796
rect 5520 10716 5560 10764
rect 5520 10684 5524 10716
rect 5556 10684 5560 10716
rect 5520 10636 5560 10684
rect 5520 10604 5524 10636
rect 5556 10604 5560 10636
rect 5520 10556 5560 10604
rect 5520 10524 5524 10556
rect 5556 10524 5560 10556
rect 5520 10476 5560 10524
rect 5520 10444 5524 10476
rect 5556 10444 5560 10476
rect 5520 10396 5560 10444
rect 5520 10364 5524 10396
rect 5556 10364 5560 10396
rect 5520 10316 5560 10364
rect 5520 10284 5524 10316
rect 5556 10284 5560 10316
rect 5520 10236 5560 10284
rect 5520 10204 5524 10236
rect 5556 10204 5560 10236
rect 5520 10156 5560 10204
rect 5520 10124 5524 10156
rect 5556 10124 5560 10156
rect 5520 10076 5560 10124
rect 5520 10044 5524 10076
rect 5556 10044 5560 10076
rect 5520 9996 5560 10044
rect 5520 9964 5524 9996
rect 5556 9964 5560 9996
rect 5520 9916 5560 9964
rect 5520 9884 5524 9916
rect 5556 9884 5560 9916
rect 5520 9836 5560 9884
rect 5520 9804 5524 9836
rect 5556 9804 5560 9836
rect 5520 9756 5560 9804
rect 5520 9724 5524 9756
rect 5556 9724 5560 9756
rect 5520 9356 5560 9724
rect 5520 9324 5524 9356
rect 5556 9324 5560 9356
rect 5520 9276 5560 9324
rect 5520 9244 5524 9276
rect 5556 9244 5560 9276
rect 5520 9196 5560 9244
rect 5520 9164 5524 9196
rect 5556 9164 5560 9196
rect 5520 8876 5560 9164
rect 5520 8844 5524 8876
rect 5556 8844 5560 8876
rect 5520 8796 5560 8844
rect 5520 8764 5524 8796
rect 5556 8764 5560 8796
rect 5520 8716 5560 8764
rect 5520 8684 5524 8716
rect 5556 8684 5560 8716
rect 5520 8636 5560 8684
rect 5520 8604 5524 8636
rect 5556 8604 5560 8636
rect 5520 8556 5560 8604
rect 5520 8524 5524 8556
rect 5556 8524 5560 8556
rect 5520 8315 5560 8524
rect 5520 8285 5525 8315
rect 5555 8285 5560 8315
rect 5520 8155 5560 8285
rect 5520 8125 5525 8155
rect 5555 8125 5560 8155
rect 5520 8075 5560 8125
rect 5520 8045 5525 8075
rect 5555 8045 5560 8075
rect 5520 7755 5560 8045
rect 5520 7725 5525 7755
rect 5555 7725 5560 7755
rect 5520 7636 5560 7725
rect 5520 7604 5524 7636
rect 5556 7604 5560 7636
rect 5520 7556 5560 7604
rect 5520 7524 5524 7556
rect 5556 7524 5560 7556
rect 5520 7476 5560 7524
rect 5520 7444 5524 7476
rect 5556 7444 5560 7476
rect 5520 7396 5560 7444
rect 5520 7364 5524 7396
rect 5556 7364 5560 7396
rect 5520 7316 5560 7364
rect 5520 7284 5524 7316
rect 5556 7284 5560 7316
rect 5520 7236 5560 7284
rect 5520 7204 5524 7236
rect 5556 7204 5560 7236
rect 5520 7156 5560 7204
rect 5520 7124 5524 7156
rect 5556 7124 5560 7156
rect 5520 7076 5560 7124
rect 5520 7044 5524 7076
rect 5556 7044 5560 7076
rect 5520 6756 5560 7044
rect 5520 6724 5524 6756
rect 5556 6724 5560 6756
rect 5520 6676 5560 6724
rect 5520 6644 5524 6676
rect 5556 6644 5560 6676
rect 5520 6596 5560 6644
rect 5520 6564 5524 6596
rect 5556 6564 5560 6596
rect 5520 6516 5560 6564
rect 5520 6484 5524 6516
rect 5556 6484 5560 6516
rect 5520 6436 5560 6484
rect 5520 6404 5524 6436
rect 5556 6404 5560 6436
rect 5520 6356 5560 6404
rect 5520 6324 5524 6356
rect 5556 6324 5560 6356
rect 5520 5796 5560 6324
rect 5520 5764 5524 5796
rect 5556 5764 5560 5796
rect 5520 5716 5560 5764
rect 5520 5684 5524 5716
rect 5556 5684 5560 5716
rect 5520 5636 5560 5684
rect 5520 5604 5524 5636
rect 5556 5604 5560 5636
rect 5520 5556 5560 5604
rect 5520 5524 5524 5556
rect 5556 5524 5560 5556
rect 5520 5476 5560 5524
rect 5520 5444 5524 5476
rect 5556 5444 5560 5476
rect 5520 5396 5560 5444
rect 5520 5364 5524 5396
rect 5556 5364 5560 5396
rect 5520 5316 5560 5364
rect 5520 5284 5524 5316
rect 5556 5284 5560 5316
rect 5520 5236 5560 5284
rect 5520 5204 5524 5236
rect 5556 5204 5560 5236
rect 5520 5156 5560 5204
rect 5520 5124 5524 5156
rect 5556 5124 5560 5156
rect 5520 5076 5560 5124
rect 5520 5044 5524 5076
rect 5556 5044 5560 5076
rect 5520 4996 5560 5044
rect 5520 4964 5524 4996
rect 5556 4964 5560 4996
rect 5520 4436 5560 4964
rect 5520 4404 5524 4436
rect 5556 4404 5560 4436
rect 5520 4356 5560 4404
rect 5520 4324 5524 4356
rect 5556 4324 5560 4356
rect 5520 4276 5560 4324
rect 5520 4244 5524 4276
rect 5556 4244 5560 4276
rect 5520 4196 5560 4244
rect 5520 4164 5524 4196
rect 5556 4164 5560 4196
rect 5520 4116 5560 4164
rect 5520 4084 5524 4116
rect 5556 4084 5560 4116
rect 5520 4036 5560 4084
rect 5520 4004 5524 4036
rect 5556 4004 5560 4036
rect 5520 3956 5560 4004
rect 5520 3924 5524 3956
rect 5556 3924 5560 3956
rect 5520 3156 5560 3924
rect 5520 3124 5524 3156
rect 5556 3124 5560 3156
rect 5520 3076 5560 3124
rect 5520 3044 5524 3076
rect 5556 3044 5560 3076
rect 5520 2996 5560 3044
rect 5520 2964 5524 2996
rect 5556 2964 5560 2996
rect 5520 2916 5560 2964
rect 5520 2884 5524 2916
rect 5556 2884 5560 2916
rect 5520 2836 5560 2884
rect 5520 2804 5524 2836
rect 5556 2804 5560 2836
rect 5520 2756 5560 2804
rect 5520 2724 5524 2756
rect 5556 2724 5560 2756
rect 5520 2676 5560 2724
rect 5520 2644 5524 2676
rect 5556 2644 5560 2676
rect 5520 2596 5560 2644
rect 5520 2564 5524 2596
rect 5556 2564 5560 2596
rect 5520 2516 5560 2564
rect 5520 2484 5524 2516
rect 5556 2484 5560 2516
rect 5520 2436 5560 2484
rect 5520 2404 5524 2436
rect 5556 2404 5560 2436
rect 5520 2356 5560 2404
rect 5520 2324 5524 2356
rect 5556 2324 5560 2356
rect 5520 2276 5560 2324
rect 5520 2244 5524 2276
rect 5556 2244 5560 2276
rect 5520 2196 5560 2244
rect 5520 2164 5524 2196
rect 5556 2164 5560 2196
rect 5520 2116 5560 2164
rect 5520 2084 5524 2116
rect 5556 2084 5560 2116
rect 5520 2036 5560 2084
rect 5520 2004 5524 2036
rect 5556 2004 5560 2036
rect 5520 1636 5560 2004
rect 5520 1604 5524 1636
rect 5556 1604 5560 1636
rect 5520 1556 5560 1604
rect 5520 1524 5524 1556
rect 5556 1524 5560 1556
rect 5520 1476 5560 1524
rect 5520 1444 5524 1476
rect 5556 1444 5560 1476
rect 5520 1396 5560 1444
rect 5520 1364 5524 1396
rect 5556 1364 5560 1396
rect 5520 1316 5560 1364
rect 5520 1284 5524 1316
rect 5556 1284 5560 1316
rect 5520 1236 5560 1284
rect 5520 1204 5524 1236
rect 5556 1204 5560 1236
rect 5520 1156 5560 1204
rect 5520 1124 5524 1156
rect 5556 1124 5560 1156
rect 5520 1076 5560 1124
rect 5520 1044 5524 1076
rect 5556 1044 5560 1076
rect 5520 756 5560 1044
rect 5520 724 5524 756
rect 5556 724 5560 756
rect 5520 676 5560 724
rect 5520 644 5524 676
rect 5556 644 5560 676
rect 5520 596 5560 644
rect 5520 564 5524 596
rect 5556 564 5560 596
rect 5520 196 5560 564
rect 5520 164 5524 196
rect 5556 164 5560 196
rect 5520 116 5560 164
rect 5520 84 5524 116
rect 5556 84 5560 116
rect 5520 36 5560 84
rect 5520 4 5524 36
rect 5556 4 5560 36
rect 5520 -40 5560 4
rect 5600 11235 5640 12680
rect 5600 11205 5605 11235
rect 5635 11205 5640 11235
rect 5600 8235 5640 11205
rect 5600 8205 5605 8235
rect 5635 8205 5640 8235
rect 5600 -40 5640 8205
rect 5680 12636 5720 13204
rect 5840 13396 5880 13400
rect 5840 13204 5844 13396
rect 5876 13204 5880 13396
rect 5680 12604 5684 12636
rect 5716 12604 5720 12636
rect 5680 12556 5720 12604
rect 5680 12524 5684 12556
rect 5716 12524 5720 12556
rect 5680 12476 5720 12524
rect 5680 12444 5684 12476
rect 5716 12444 5720 12476
rect 5680 12396 5720 12444
rect 5680 12364 5684 12396
rect 5716 12364 5720 12396
rect 5680 12316 5720 12364
rect 5680 12284 5684 12316
rect 5716 12284 5720 12316
rect 5680 12236 5720 12284
rect 5680 12204 5684 12236
rect 5716 12204 5720 12236
rect 5680 12156 5720 12204
rect 5680 12124 5684 12156
rect 5716 12124 5720 12156
rect 5680 11836 5720 12124
rect 5680 11804 5684 11836
rect 5716 11804 5720 11836
rect 5680 11756 5720 11804
rect 5680 11724 5684 11756
rect 5716 11724 5720 11756
rect 5680 11676 5720 11724
rect 5680 11644 5684 11676
rect 5716 11644 5720 11676
rect 5680 11596 5720 11644
rect 5680 11564 5684 11596
rect 5716 11564 5720 11596
rect 5680 11516 5720 11564
rect 5680 11484 5684 11516
rect 5716 11484 5720 11516
rect 5680 11436 5720 11484
rect 5680 11404 5684 11436
rect 5716 11404 5720 11436
rect 5680 11315 5720 11404
rect 5680 11285 5685 11315
rect 5715 11285 5720 11315
rect 5680 11155 5720 11285
rect 5680 11125 5685 11155
rect 5715 11125 5720 11155
rect 5680 10876 5720 11125
rect 5680 10844 5684 10876
rect 5716 10844 5720 10876
rect 5680 10796 5720 10844
rect 5680 10764 5684 10796
rect 5716 10764 5720 10796
rect 5680 10716 5720 10764
rect 5680 10684 5684 10716
rect 5716 10684 5720 10716
rect 5680 10636 5720 10684
rect 5680 10604 5684 10636
rect 5716 10604 5720 10636
rect 5680 10556 5720 10604
rect 5680 10524 5684 10556
rect 5716 10524 5720 10556
rect 5680 10476 5720 10524
rect 5680 10444 5684 10476
rect 5716 10444 5720 10476
rect 5680 10396 5720 10444
rect 5680 10364 5684 10396
rect 5716 10364 5720 10396
rect 5680 10316 5720 10364
rect 5680 10284 5684 10316
rect 5716 10284 5720 10316
rect 5680 10236 5720 10284
rect 5680 10204 5684 10236
rect 5716 10204 5720 10236
rect 5680 10156 5720 10204
rect 5680 10124 5684 10156
rect 5716 10124 5720 10156
rect 5680 10076 5720 10124
rect 5680 10044 5684 10076
rect 5716 10044 5720 10076
rect 5680 9996 5720 10044
rect 5680 9964 5684 9996
rect 5716 9964 5720 9996
rect 5680 9916 5720 9964
rect 5680 9884 5684 9916
rect 5716 9884 5720 9916
rect 5680 9836 5720 9884
rect 5680 9804 5684 9836
rect 5716 9804 5720 9836
rect 5680 9756 5720 9804
rect 5680 9724 5684 9756
rect 5716 9724 5720 9756
rect 5680 9356 5720 9724
rect 5680 9324 5684 9356
rect 5716 9324 5720 9356
rect 5680 9276 5720 9324
rect 5680 9244 5684 9276
rect 5716 9244 5720 9276
rect 5680 9196 5720 9244
rect 5680 9164 5684 9196
rect 5716 9164 5720 9196
rect 5680 8876 5720 9164
rect 5680 8844 5684 8876
rect 5716 8844 5720 8876
rect 5680 8796 5720 8844
rect 5680 8764 5684 8796
rect 5716 8764 5720 8796
rect 5680 8716 5720 8764
rect 5680 8684 5684 8716
rect 5716 8684 5720 8716
rect 5680 8636 5720 8684
rect 5680 8604 5684 8636
rect 5716 8604 5720 8636
rect 5680 8556 5720 8604
rect 5680 8524 5684 8556
rect 5716 8524 5720 8556
rect 5680 8475 5720 8524
rect 5680 8445 5685 8475
rect 5715 8445 5720 8475
rect 5680 8315 5720 8445
rect 5680 8285 5685 8315
rect 5715 8285 5720 8315
rect 5680 8155 5720 8285
rect 5680 8125 5685 8155
rect 5715 8125 5720 8155
rect 5680 7636 5720 8125
rect 5680 7604 5684 7636
rect 5716 7604 5720 7636
rect 5680 7556 5720 7604
rect 5680 7524 5684 7556
rect 5716 7524 5720 7556
rect 5680 7476 5720 7524
rect 5680 7444 5684 7476
rect 5716 7444 5720 7476
rect 5680 7396 5720 7444
rect 5680 7364 5684 7396
rect 5716 7364 5720 7396
rect 5680 7316 5720 7364
rect 5680 7284 5684 7316
rect 5716 7284 5720 7316
rect 5680 7236 5720 7284
rect 5680 7204 5684 7236
rect 5716 7204 5720 7236
rect 5680 7156 5720 7204
rect 5680 7124 5684 7156
rect 5716 7124 5720 7156
rect 5680 7076 5720 7124
rect 5680 7044 5684 7076
rect 5716 7044 5720 7076
rect 5680 6756 5720 7044
rect 5680 6724 5684 6756
rect 5716 6724 5720 6756
rect 5680 6676 5720 6724
rect 5680 6644 5684 6676
rect 5716 6644 5720 6676
rect 5680 6596 5720 6644
rect 5680 6564 5684 6596
rect 5716 6564 5720 6596
rect 5680 6516 5720 6564
rect 5680 6484 5684 6516
rect 5716 6484 5720 6516
rect 5680 6436 5720 6484
rect 5680 6404 5684 6436
rect 5716 6404 5720 6436
rect 5680 6356 5720 6404
rect 5680 6324 5684 6356
rect 5716 6324 5720 6356
rect 5680 5796 5720 6324
rect 5680 5764 5684 5796
rect 5716 5764 5720 5796
rect 5680 5716 5720 5764
rect 5680 5684 5684 5716
rect 5716 5684 5720 5716
rect 5680 5636 5720 5684
rect 5680 5604 5684 5636
rect 5716 5604 5720 5636
rect 5680 5556 5720 5604
rect 5680 5524 5684 5556
rect 5716 5524 5720 5556
rect 5680 5476 5720 5524
rect 5680 5444 5684 5476
rect 5716 5444 5720 5476
rect 5680 5396 5720 5444
rect 5680 5364 5684 5396
rect 5716 5364 5720 5396
rect 5680 5316 5720 5364
rect 5680 5284 5684 5316
rect 5716 5284 5720 5316
rect 5680 5236 5720 5284
rect 5680 5204 5684 5236
rect 5716 5204 5720 5236
rect 5680 5156 5720 5204
rect 5680 5124 5684 5156
rect 5716 5124 5720 5156
rect 5680 5076 5720 5124
rect 5680 5044 5684 5076
rect 5716 5044 5720 5076
rect 5680 4996 5720 5044
rect 5680 4964 5684 4996
rect 5716 4964 5720 4996
rect 5680 4436 5720 4964
rect 5680 4404 5684 4436
rect 5716 4404 5720 4436
rect 5680 4356 5720 4404
rect 5680 4324 5684 4356
rect 5716 4324 5720 4356
rect 5680 4276 5720 4324
rect 5680 4244 5684 4276
rect 5716 4244 5720 4276
rect 5680 4196 5720 4244
rect 5680 4164 5684 4196
rect 5716 4164 5720 4196
rect 5680 4116 5720 4164
rect 5680 4084 5684 4116
rect 5716 4084 5720 4116
rect 5680 4036 5720 4084
rect 5680 4004 5684 4036
rect 5716 4004 5720 4036
rect 5680 3956 5720 4004
rect 5680 3924 5684 3956
rect 5716 3924 5720 3956
rect 5680 3156 5720 3924
rect 5680 3124 5684 3156
rect 5716 3124 5720 3156
rect 5680 3076 5720 3124
rect 5680 3044 5684 3076
rect 5716 3044 5720 3076
rect 5680 2996 5720 3044
rect 5680 2964 5684 2996
rect 5716 2964 5720 2996
rect 5680 2916 5720 2964
rect 5680 2884 5684 2916
rect 5716 2884 5720 2916
rect 5680 2836 5720 2884
rect 5680 2804 5684 2836
rect 5716 2804 5720 2836
rect 5680 2756 5720 2804
rect 5680 2724 5684 2756
rect 5716 2724 5720 2756
rect 5680 2676 5720 2724
rect 5680 2644 5684 2676
rect 5716 2644 5720 2676
rect 5680 2596 5720 2644
rect 5680 2564 5684 2596
rect 5716 2564 5720 2596
rect 5680 2516 5720 2564
rect 5680 2484 5684 2516
rect 5716 2484 5720 2516
rect 5680 2436 5720 2484
rect 5680 2404 5684 2436
rect 5716 2404 5720 2436
rect 5680 2356 5720 2404
rect 5680 2324 5684 2356
rect 5716 2324 5720 2356
rect 5680 2276 5720 2324
rect 5680 2244 5684 2276
rect 5716 2244 5720 2276
rect 5680 2196 5720 2244
rect 5680 2164 5684 2196
rect 5716 2164 5720 2196
rect 5680 2116 5720 2164
rect 5680 2084 5684 2116
rect 5716 2084 5720 2116
rect 5680 2036 5720 2084
rect 5680 2004 5684 2036
rect 5716 2004 5720 2036
rect 5680 1636 5720 2004
rect 5680 1604 5684 1636
rect 5716 1604 5720 1636
rect 5680 1556 5720 1604
rect 5680 1524 5684 1556
rect 5716 1524 5720 1556
rect 5680 1476 5720 1524
rect 5680 1444 5684 1476
rect 5716 1444 5720 1476
rect 5680 1396 5720 1444
rect 5680 1364 5684 1396
rect 5716 1364 5720 1396
rect 5680 1316 5720 1364
rect 5680 1284 5684 1316
rect 5716 1284 5720 1316
rect 5680 1236 5720 1284
rect 5680 1204 5684 1236
rect 5716 1204 5720 1236
rect 5680 1156 5720 1204
rect 5680 1124 5684 1156
rect 5716 1124 5720 1156
rect 5680 1076 5720 1124
rect 5680 1044 5684 1076
rect 5716 1044 5720 1076
rect 5680 756 5720 1044
rect 5680 724 5684 756
rect 5716 724 5720 756
rect 5680 676 5720 724
rect 5680 644 5684 676
rect 5716 644 5720 676
rect 5680 596 5720 644
rect 5680 564 5684 596
rect 5716 564 5720 596
rect 5680 196 5720 564
rect 5680 164 5684 196
rect 5716 164 5720 196
rect 5680 116 5720 164
rect 5680 84 5684 116
rect 5716 84 5720 116
rect 5680 36 5720 84
rect 5680 4 5684 36
rect 5716 4 5720 36
rect 5680 -40 5720 4
rect 5760 8395 5800 12680
rect 5760 8365 5765 8395
rect 5795 8365 5800 8395
rect 5760 -40 5800 8365
rect 5840 12636 5880 13204
rect 6160 13396 6200 13400
rect 6160 13204 6164 13396
rect 6196 13204 6200 13396
rect 5840 12604 5844 12636
rect 5876 12604 5880 12636
rect 5840 12556 5880 12604
rect 5840 12524 5844 12556
rect 5876 12524 5880 12556
rect 5840 12476 5880 12524
rect 5840 12444 5844 12476
rect 5876 12444 5880 12476
rect 5840 12396 5880 12444
rect 5840 12364 5844 12396
rect 5876 12364 5880 12396
rect 5840 12316 5880 12364
rect 5840 12284 5844 12316
rect 5876 12284 5880 12316
rect 5840 12236 5880 12284
rect 5840 12204 5844 12236
rect 5876 12204 5880 12236
rect 5840 12156 5880 12204
rect 5840 12124 5844 12156
rect 5876 12124 5880 12156
rect 5840 11836 5880 12124
rect 5840 11804 5844 11836
rect 5876 11804 5880 11836
rect 5840 11756 5880 11804
rect 5840 11724 5844 11756
rect 5876 11724 5880 11756
rect 5840 11676 5880 11724
rect 5840 11644 5844 11676
rect 5876 11644 5880 11676
rect 5840 11596 5880 11644
rect 5840 11564 5844 11596
rect 5876 11564 5880 11596
rect 5840 11516 5880 11564
rect 5840 11484 5844 11516
rect 5876 11484 5880 11516
rect 5840 11436 5880 11484
rect 5840 11404 5844 11436
rect 5876 11404 5880 11436
rect 5840 10876 5880 11404
rect 5840 10844 5844 10876
rect 5876 10844 5880 10876
rect 5840 10796 5880 10844
rect 5840 10764 5844 10796
rect 5876 10764 5880 10796
rect 5840 10716 5880 10764
rect 5840 10684 5844 10716
rect 5876 10684 5880 10716
rect 5840 10636 5880 10684
rect 5840 10604 5844 10636
rect 5876 10604 5880 10636
rect 5840 10556 5880 10604
rect 5840 10524 5844 10556
rect 5876 10524 5880 10556
rect 5840 10476 5880 10524
rect 5840 10444 5844 10476
rect 5876 10444 5880 10476
rect 5840 10396 5880 10444
rect 5840 10364 5844 10396
rect 5876 10364 5880 10396
rect 5840 10316 5880 10364
rect 5840 10284 5844 10316
rect 5876 10284 5880 10316
rect 5840 10236 5880 10284
rect 5840 10204 5844 10236
rect 5876 10204 5880 10236
rect 5840 10156 5880 10204
rect 5840 10124 5844 10156
rect 5876 10124 5880 10156
rect 5840 10076 5880 10124
rect 5840 10044 5844 10076
rect 5876 10044 5880 10076
rect 5840 9996 5880 10044
rect 5840 9964 5844 9996
rect 5876 9964 5880 9996
rect 5840 9916 5880 9964
rect 5840 9884 5844 9916
rect 5876 9884 5880 9916
rect 5840 9836 5880 9884
rect 5840 9804 5844 9836
rect 5876 9804 5880 9836
rect 5840 9756 5880 9804
rect 5840 9724 5844 9756
rect 5876 9724 5880 9756
rect 5840 9356 5880 9724
rect 5840 9324 5844 9356
rect 5876 9324 5880 9356
rect 5840 9276 5880 9324
rect 5840 9244 5844 9276
rect 5876 9244 5880 9276
rect 5840 9196 5880 9244
rect 5840 9164 5844 9196
rect 5876 9164 5880 9196
rect 5840 8876 5880 9164
rect 5840 8844 5844 8876
rect 5876 8844 5880 8876
rect 5840 8796 5880 8844
rect 5840 8764 5844 8796
rect 5876 8764 5880 8796
rect 5840 8716 5880 8764
rect 5840 8684 5844 8716
rect 5876 8684 5880 8716
rect 5840 8636 5880 8684
rect 5840 8604 5844 8636
rect 5876 8604 5880 8636
rect 5840 8556 5880 8604
rect 5840 8524 5844 8556
rect 5876 8524 5880 8556
rect 5840 8475 5880 8524
rect 5840 8445 5845 8475
rect 5875 8445 5880 8475
rect 5840 8315 5880 8445
rect 5840 8285 5845 8315
rect 5875 8285 5880 8315
rect 5840 7636 5880 8285
rect 5840 7604 5844 7636
rect 5876 7604 5880 7636
rect 5840 7556 5880 7604
rect 5840 7524 5844 7556
rect 5876 7524 5880 7556
rect 5840 7476 5880 7524
rect 5840 7444 5844 7476
rect 5876 7444 5880 7476
rect 5840 7396 5880 7444
rect 5840 7364 5844 7396
rect 5876 7364 5880 7396
rect 5840 7316 5880 7364
rect 5840 7284 5844 7316
rect 5876 7284 5880 7316
rect 5840 7236 5880 7284
rect 5840 7204 5844 7236
rect 5876 7204 5880 7236
rect 5840 7156 5880 7204
rect 5840 7124 5844 7156
rect 5876 7124 5880 7156
rect 5840 7076 5880 7124
rect 5840 7044 5844 7076
rect 5876 7044 5880 7076
rect 5840 6756 5880 7044
rect 5840 6724 5844 6756
rect 5876 6724 5880 6756
rect 5840 6676 5880 6724
rect 5840 6644 5844 6676
rect 5876 6644 5880 6676
rect 5840 6596 5880 6644
rect 5840 6564 5844 6596
rect 5876 6564 5880 6596
rect 5840 6516 5880 6564
rect 5840 6484 5844 6516
rect 5876 6484 5880 6516
rect 5840 6436 5880 6484
rect 5840 6404 5844 6436
rect 5876 6404 5880 6436
rect 5840 6356 5880 6404
rect 5840 6324 5844 6356
rect 5876 6324 5880 6356
rect 5840 5796 5880 6324
rect 5840 5764 5844 5796
rect 5876 5764 5880 5796
rect 5840 5716 5880 5764
rect 5840 5684 5844 5716
rect 5876 5684 5880 5716
rect 5840 5636 5880 5684
rect 5840 5604 5844 5636
rect 5876 5604 5880 5636
rect 5840 5556 5880 5604
rect 5840 5524 5844 5556
rect 5876 5524 5880 5556
rect 5840 5476 5880 5524
rect 5840 5444 5844 5476
rect 5876 5444 5880 5476
rect 5840 5396 5880 5444
rect 5840 5364 5844 5396
rect 5876 5364 5880 5396
rect 5840 5316 5880 5364
rect 5840 5284 5844 5316
rect 5876 5284 5880 5316
rect 5840 5236 5880 5284
rect 5840 5204 5844 5236
rect 5876 5204 5880 5236
rect 5840 5156 5880 5204
rect 5840 5124 5844 5156
rect 5876 5124 5880 5156
rect 5840 5076 5880 5124
rect 5840 5044 5844 5076
rect 5876 5044 5880 5076
rect 5840 4996 5880 5044
rect 5840 4964 5844 4996
rect 5876 4964 5880 4996
rect 5840 4436 5880 4964
rect 5840 4404 5844 4436
rect 5876 4404 5880 4436
rect 5840 4356 5880 4404
rect 5840 4324 5844 4356
rect 5876 4324 5880 4356
rect 5840 4276 5880 4324
rect 5840 4244 5844 4276
rect 5876 4244 5880 4276
rect 5840 4196 5880 4244
rect 5840 4164 5844 4196
rect 5876 4164 5880 4196
rect 5840 4116 5880 4164
rect 5840 4084 5844 4116
rect 5876 4084 5880 4116
rect 5840 4036 5880 4084
rect 5840 4004 5844 4036
rect 5876 4004 5880 4036
rect 5840 3956 5880 4004
rect 5840 3924 5844 3956
rect 5876 3924 5880 3956
rect 5840 3156 5880 3924
rect 5840 3124 5844 3156
rect 5876 3124 5880 3156
rect 5840 3076 5880 3124
rect 5840 3044 5844 3076
rect 5876 3044 5880 3076
rect 5840 2996 5880 3044
rect 5840 2964 5844 2996
rect 5876 2964 5880 2996
rect 5840 2916 5880 2964
rect 5840 2884 5844 2916
rect 5876 2884 5880 2916
rect 5840 2836 5880 2884
rect 5840 2804 5844 2836
rect 5876 2804 5880 2836
rect 5840 2756 5880 2804
rect 5840 2724 5844 2756
rect 5876 2724 5880 2756
rect 5840 2676 5880 2724
rect 5840 2644 5844 2676
rect 5876 2644 5880 2676
rect 5840 2596 5880 2644
rect 5840 2564 5844 2596
rect 5876 2564 5880 2596
rect 5840 2516 5880 2564
rect 5840 2484 5844 2516
rect 5876 2484 5880 2516
rect 5840 2436 5880 2484
rect 5840 2404 5844 2436
rect 5876 2404 5880 2436
rect 5840 2356 5880 2404
rect 5840 2324 5844 2356
rect 5876 2324 5880 2356
rect 5840 2276 5880 2324
rect 5840 2244 5844 2276
rect 5876 2244 5880 2276
rect 5840 2196 5880 2244
rect 5840 2164 5844 2196
rect 5876 2164 5880 2196
rect 5840 2116 5880 2164
rect 5840 2084 5844 2116
rect 5876 2084 5880 2116
rect 5840 2036 5880 2084
rect 5840 2004 5844 2036
rect 5876 2004 5880 2036
rect 5840 1636 5880 2004
rect 5840 1604 5844 1636
rect 5876 1604 5880 1636
rect 5840 1556 5880 1604
rect 5840 1524 5844 1556
rect 5876 1524 5880 1556
rect 5840 1476 5880 1524
rect 5840 1444 5844 1476
rect 5876 1444 5880 1476
rect 5840 1396 5880 1444
rect 5840 1364 5844 1396
rect 5876 1364 5880 1396
rect 5840 1316 5880 1364
rect 5840 1284 5844 1316
rect 5876 1284 5880 1316
rect 5840 1236 5880 1284
rect 5840 1204 5844 1236
rect 5876 1204 5880 1236
rect 5840 1156 5880 1204
rect 5840 1124 5844 1156
rect 5876 1124 5880 1156
rect 5840 1076 5880 1124
rect 5840 1044 5844 1076
rect 5876 1044 5880 1076
rect 5840 756 5880 1044
rect 5840 724 5844 756
rect 5876 724 5880 756
rect 5840 676 5880 724
rect 5840 644 5844 676
rect 5876 644 5880 676
rect 5840 596 5880 644
rect 5840 564 5844 596
rect 5876 564 5880 596
rect 5840 196 5880 564
rect 5840 164 5844 196
rect 5876 164 5880 196
rect 5840 116 5880 164
rect 5840 84 5844 116
rect 5876 84 5880 116
rect 5840 36 5880 84
rect 5840 4 5844 36
rect 5876 4 5880 36
rect 5840 -40 5880 4
rect 5920 12916 5960 12920
rect 5920 12724 5924 12916
rect 5956 12724 5960 12916
rect 5920 12636 5960 12724
rect 6080 12916 6120 12920
rect 6080 12724 6084 12916
rect 6116 12724 6120 12916
rect 5920 12604 5924 12636
rect 5956 12604 5960 12636
rect 5920 12556 5960 12604
rect 5920 12524 5924 12556
rect 5956 12524 5960 12556
rect 5920 12476 5960 12524
rect 5920 12444 5924 12476
rect 5956 12444 5960 12476
rect 5920 12396 5960 12444
rect 5920 12364 5924 12396
rect 5956 12364 5960 12396
rect 5920 12316 5960 12364
rect 5920 12284 5924 12316
rect 5956 12284 5960 12316
rect 5920 12236 5960 12284
rect 5920 12204 5924 12236
rect 5956 12204 5960 12236
rect 5920 12156 5960 12204
rect 5920 12124 5924 12156
rect 5956 12124 5960 12156
rect 5920 11836 5960 12124
rect 5920 11804 5924 11836
rect 5956 11804 5960 11836
rect 5920 11756 5960 11804
rect 5920 11724 5924 11756
rect 5956 11724 5960 11756
rect 5920 11676 5960 11724
rect 5920 11644 5924 11676
rect 5956 11644 5960 11676
rect 5920 11596 5960 11644
rect 5920 11564 5924 11596
rect 5956 11564 5960 11596
rect 5920 11516 5960 11564
rect 5920 11484 5924 11516
rect 5956 11484 5960 11516
rect 5920 11436 5960 11484
rect 5920 11404 5924 11436
rect 5956 11404 5960 11436
rect 5920 10876 5960 11404
rect 5920 10844 5924 10876
rect 5956 10844 5960 10876
rect 5920 10796 5960 10844
rect 5920 10764 5924 10796
rect 5956 10764 5960 10796
rect 5920 10716 5960 10764
rect 5920 10684 5924 10716
rect 5956 10684 5960 10716
rect 5920 10636 5960 10684
rect 5920 10604 5924 10636
rect 5956 10604 5960 10636
rect 5920 10556 5960 10604
rect 5920 10524 5924 10556
rect 5956 10524 5960 10556
rect 5920 10476 5960 10524
rect 5920 10444 5924 10476
rect 5956 10444 5960 10476
rect 5920 10396 5960 10444
rect 5920 10364 5924 10396
rect 5956 10364 5960 10396
rect 5920 10316 5960 10364
rect 5920 10284 5924 10316
rect 5956 10284 5960 10316
rect 5920 10236 5960 10284
rect 5920 10204 5924 10236
rect 5956 10204 5960 10236
rect 5920 10156 5960 10204
rect 5920 10124 5924 10156
rect 5956 10124 5960 10156
rect 5920 10076 5960 10124
rect 5920 10044 5924 10076
rect 5956 10044 5960 10076
rect 5920 9996 5960 10044
rect 5920 9964 5924 9996
rect 5956 9964 5960 9996
rect 5920 9916 5960 9964
rect 5920 9884 5924 9916
rect 5956 9884 5960 9916
rect 5920 9836 5960 9884
rect 5920 9804 5924 9836
rect 5956 9804 5960 9836
rect 5920 9756 5960 9804
rect 5920 9724 5924 9756
rect 5956 9724 5960 9756
rect 5920 9356 5960 9724
rect 5920 9324 5924 9356
rect 5956 9324 5960 9356
rect 5920 9276 5960 9324
rect 5920 9244 5924 9276
rect 5956 9244 5960 9276
rect 5920 9196 5960 9244
rect 5920 9164 5924 9196
rect 5956 9164 5960 9196
rect 5920 8876 5960 9164
rect 5920 8844 5924 8876
rect 5956 8844 5960 8876
rect 5920 8796 5960 8844
rect 5920 8764 5924 8796
rect 5956 8764 5960 8796
rect 5920 8716 5960 8764
rect 5920 8684 5924 8716
rect 5956 8684 5960 8716
rect 5920 8636 5960 8684
rect 5920 8604 5924 8636
rect 5956 8604 5960 8636
rect 5920 8556 5960 8604
rect 5920 8524 5924 8556
rect 5956 8524 5960 8556
rect 5920 7636 5960 8524
rect 5920 7604 5924 7636
rect 5956 7604 5960 7636
rect 5920 7556 5960 7604
rect 5920 7524 5924 7556
rect 5956 7524 5960 7556
rect 5920 7476 5960 7524
rect 5920 7444 5924 7476
rect 5956 7444 5960 7476
rect 5920 7396 5960 7444
rect 5920 7364 5924 7396
rect 5956 7364 5960 7396
rect 5920 7316 5960 7364
rect 5920 7284 5924 7316
rect 5956 7284 5960 7316
rect 5920 7236 5960 7284
rect 5920 7204 5924 7236
rect 5956 7204 5960 7236
rect 5920 7156 5960 7204
rect 5920 7124 5924 7156
rect 5956 7124 5960 7156
rect 5920 7076 5960 7124
rect 5920 7044 5924 7076
rect 5956 7044 5960 7076
rect 5920 6756 5960 7044
rect 5920 6724 5924 6756
rect 5956 6724 5960 6756
rect 5920 6676 5960 6724
rect 5920 6644 5924 6676
rect 5956 6644 5960 6676
rect 5920 6596 5960 6644
rect 5920 6564 5924 6596
rect 5956 6564 5960 6596
rect 5920 6516 5960 6564
rect 5920 6484 5924 6516
rect 5956 6484 5960 6516
rect 5920 6436 5960 6484
rect 5920 6404 5924 6436
rect 5956 6404 5960 6436
rect 5920 6356 5960 6404
rect 5920 6324 5924 6356
rect 5956 6324 5960 6356
rect 5920 5796 5960 6324
rect 5920 5764 5924 5796
rect 5956 5764 5960 5796
rect 5920 5716 5960 5764
rect 5920 5684 5924 5716
rect 5956 5684 5960 5716
rect 5920 5636 5960 5684
rect 5920 5604 5924 5636
rect 5956 5604 5960 5636
rect 5920 5556 5960 5604
rect 5920 5524 5924 5556
rect 5956 5524 5960 5556
rect 5920 5476 5960 5524
rect 5920 5444 5924 5476
rect 5956 5444 5960 5476
rect 5920 5396 5960 5444
rect 5920 5364 5924 5396
rect 5956 5364 5960 5396
rect 5920 5316 5960 5364
rect 5920 5284 5924 5316
rect 5956 5284 5960 5316
rect 5920 5236 5960 5284
rect 5920 5204 5924 5236
rect 5956 5204 5960 5236
rect 5920 5156 5960 5204
rect 5920 5124 5924 5156
rect 5956 5124 5960 5156
rect 5920 5076 5960 5124
rect 5920 5044 5924 5076
rect 5956 5044 5960 5076
rect 5920 4996 5960 5044
rect 5920 4964 5924 4996
rect 5956 4964 5960 4996
rect 5920 4915 5960 4964
rect 5920 4885 5925 4915
rect 5955 4885 5960 4915
rect 5920 4755 5960 4885
rect 5920 4725 5925 4755
rect 5955 4725 5960 4755
rect 5920 4436 5960 4725
rect 5920 4404 5924 4436
rect 5956 4404 5960 4436
rect 5920 4356 5960 4404
rect 5920 4324 5924 4356
rect 5956 4324 5960 4356
rect 5920 4276 5960 4324
rect 5920 4244 5924 4276
rect 5956 4244 5960 4276
rect 5920 4196 5960 4244
rect 5920 4164 5924 4196
rect 5956 4164 5960 4196
rect 5920 4116 5960 4164
rect 5920 4084 5924 4116
rect 5956 4084 5960 4116
rect 5920 4036 5960 4084
rect 5920 4004 5924 4036
rect 5956 4004 5960 4036
rect 5920 3956 5960 4004
rect 5920 3924 5924 3956
rect 5956 3924 5960 3956
rect 5920 3395 5960 3924
rect 5920 3365 5925 3395
rect 5955 3365 5960 3395
rect 5920 3235 5960 3365
rect 5920 3205 5925 3235
rect 5955 3205 5960 3235
rect 5920 3156 5960 3205
rect 5920 3124 5924 3156
rect 5956 3124 5960 3156
rect 5920 3076 5960 3124
rect 5920 3044 5924 3076
rect 5956 3044 5960 3076
rect 5920 2996 5960 3044
rect 5920 2964 5924 2996
rect 5956 2964 5960 2996
rect 5920 2916 5960 2964
rect 5920 2884 5924 2916
rect 5956 2884 5960 2916
rect 5920 2836 5960 2884
rect 5920 2804 5924 2836
rect 5956 2804 5960 2836
rect 5920 2756 5960 2804
rect 5920 2724 5924 2756
rect 5956 2724 5960 2756
rect 5920 2676 5960 2724
rect 5920 2644 5924 2676
rect 5956 2644 5960 2676
rect 5920 2596 5960 2644
rect 5920 2564 5924 2596
rect 5956 2564 5960 2596
rect 5920 2516 5960 2564
rect 5920 2484 5924 2516
rect 5956 2484 5960 2516
rect 5920 2436 5960 2484
rect 5920 2404 5924 2436
rect 5956 2404 5960 2436
rect 5920 2356 5960 2404
rect 5920 2324 5924 2356
rect 5956 2324 5960 2356
rect 5920 2276 5960 2324
rect 5920 2244 5924 2276
rect 5956 2244 5960 2276
rect 5920 2196 5960 2244
rect 5920 2164 5924 2196
rect 5956 2164 5960 2196
rect 5920 2116 5960 2164
rect 5920 2084 5924 2116
rect 5956 2084 5960 2116
rect 5920 2036 5960 2084
rect 5920 2004 5924 2036
rect 5956 2004 5960 2036
rect 5920 1636 5960 2004
rect 5920 1604 5924 1636
rect 5956 1604 5960 1636
rect 5920 1556 5960 1604
rect 5920 1524 5924 1556
rect 5956 1524 5960 1556
rect 5920 1476 5960 1524
rect 5920 1444 5924 1476
rect 5956 1444 5960 1476
rect 5920 1396 5960 1444
rect 5920 1364 5924 1396
rect 5956 1364 5960 1396
rect 5920 1316 5960 1364
rect 5920 1284 5924 1316
rect 5956 1284 5960 1316
rect 5920 1236 5960 1284
rect 5920 1204 5924 1236
rect 5956 1204 5960 1236
rect 5920 1156 5960 1204
rect 5920 1124 5924 1156
rect 5956 1124 5960 1156
rect 5920 1076 5960 1124
rect 5920 1044 5924 1076
rect 5956 1044 5960 1076
rect 5920 756 5960 1044
rect 5920 724 5924 756
rect 5956 724 5960 756
rect 5920 676 5960 724
rect 5920 644 5924 676
rect 5956 644 5960 676
rect 5920 596 5960 644
rect 5920 564 5924 596
rect 5956 564 5960 596
rect 5920 196 5960 564
rect 5920 164 5924 196
rect 5956 164 5960 196
rect 5920 116 5960 164
rect 5920 84 5924 116
rect 5956 84 5960 116
rect 5920 36 5960 84
rect 5920 4 5924 36
rect 5956 4 5960 36
rect 5920 -40 5960 4
rect 6000 4835 6040 12680
rect 6000 4805 6005 4835
rect 6035 4805 6040 4835
rect 6000 3315 6040 4805
rect 6000 3285 6005 3315
rect 6035 3285 6040 3315
rect 6000 -40 6040 3285
rect 6080 12636 6120 12724
rect 6080 12604 6084 12636
rect 6116 12604 6120 12636
rect 6080 12556 6120 12604
rect 6080 12524 6084 12556
rect 6116 12524 6120 12556
rect 6080 12476 6120 12524
rect 6080 12444 6084 12476
rect 6116 12444 6120 12476
rect 6080 12396 6120 12444
rect 6080 12364 6084 12396
rect 6116 12364 6120 12396
rect 6080 12316 6120 12364
rect 6080 12284 6084 12316
rect 6116 12284 6120 12316
rect 6080 12236 6120 12284
rect 6080 12204 6084 12236
rect 6116 12204 6120 12236
rect 6080 12156 6120 12204
rect 6080 12124 6084 12156
rect 6116 12124 6120 12156
rect 6080 11836 6120 12124
rect 6080 11804 6084 11836
rect 6116 11804 6120 11836
rect 6080 11756 6120 11804
rect 6080 11724 6084 11756
rect 6116 11724 6120 11756
rect 6080 11676 6120 11724
rect 6080 11644 6084 11676
rect 6116 11644 6120 11676
rect 6080 11596 6120 11644
rect 6080 11564 6084 11596
rect 6116 11564 6120 11596
rect 6080 11516 6120 11564
rect 6080 11484 6084 11516
rect 6116 11484 6120 11516
rect 6080 11436 6120 11484
rect 6080 11404 6084 11436
rect 6116 11404 6120 11436
rect 6080 10876 6120 11404
rect 6080 10844 6084 10876
rect 6116 10844 6120 10876
rect 6080 10796 6120 10844
rect 6080 10764 6084 10796
rect 6116 10764 6120 10796
rect 6080 10716 6120 10764
rect 6080 10684 6084 10716
rect 6116 10684 6120 10716
rect 6080 10636 6120 10684
rect 6080 10604 6084 10636
rect 6116 10604 6120 10636
rect 6080 10556 6120 10604
rect 6080 10524 6084 10556
rect 6116 10524 6120 10556
rect 6080 10476 6120 10524
rect 6080 10444 6084 10476
rect 6116 10444 6120 10476
rect 6080 10396 6120 10444
rect 6080 10364 6084 10396
rect 6116 10364 6120 10396
rect 6080 10316 6120 10364
rect 6080 10284 6084 10316
rect 6116 10284 6120 10316
rect 6080 10236 6120 10284
rect 6080 10204 6084 10236
rect 6116 10204 6120 10236
rect 6080 10156 6120 10204
rect 6080 10124 6084 10156
rect 6116 10124 6120 10156
rect 6080 10076 6120 10124
rect 6080 10044 6084 10076
rect 6116 10044 6120 10076
rect 6080 9996 6120 10044
rect 6080 9964 6084 9996
rect 6116 9964 6120 9996
rect 6080 9916 6120 9964
rect 6080 9884 6084 9916
rect 6116 9884 6120 9916
rect 6080 9836 6120 9884
rect 6080 9804 6084 9836
rect 6116 9804 6120 9836
rect 6080 9756 6120 9804
rect 6080 9724 6084 9756
rect 6116 9724 6120 9756
rect 6080 9356 6120 9724
rect 6080 9324 6084 9356
rect 6116 9324 6120 9356
rect 6080 9276 6120 9324
rect 6080 9244 6084 9276
rect 6116 9244 6120 9276
rect 6080 9196 6120 9244
rect 6080 9164 6084 9196
rect 6116 9164 6120 9196
rect 6080 8876 6120 9164
rect 6080 8844 6084 8876
rect 6116 8844 6120 8876
rect 6080 8796 6120 8844
rect 6080 8764 6084 8796
rect 6116 8764 6120 8796
rect 6080 8716 6120 8764
rect 6080 8684 6084 8716
rect 6116 8684 6120 8716
rect 6080 8636 6120 8684
rect 6080 8604 6084 8636
rect 6116 8604 6120 8636
rect 6080 8556 6120 8604
rect 6080 8524 6084 8556
rect 6116 8524 6120 8556
rect 6080 7636 6120 8524
rect 6080 7604 6084 7636
rect 6116 7604 6120 7636
rect 6080 7556 6120 7604
rect 6080 7524 6084 7556
rect 6116 7524 6120 7556
rect 6080 7476 6120 7524
rect 6080 7444 6084 7476
rect 6116 7444 6120 7476
rect 6080 7396 6120 7444
rect 6080 7364 6084 7396
rect 6116 7364 6120 7396
rect 6080 7316 6120 7364
rect 6080 7284 6084 7316
rect 6116 7284 6120 7316
rect 6080 7236 6120 7284
rect 6080 7204 6084 7236
rect 6116 7204 6120 7236
rect 6080 7156 6120 7204
rect 6080 7124 6084 7156
rect 6116 7124 6120 7156
rect 6080 7076 6120 7124
rect 6080 7044 6084 7076
rect 6116 7044 6120 7076
rect 6080 6756 6120 7044
rect 6080 6724 6084 6756
rect 6116 6724 6120 6756
rect 6080 6676 6120 6724
rect 6080 6644 6084 6676
rect 6116 6644 6120 6676
rect 6080 6596 6120 6644
rect 6080 6564 6084 6596
rect 6116 6564 6120 6596
rect 6080 6516 6120 6564
rect 6080 6484 6084 6516
rect 6116 6484 6120 6516
rect 6080 6436 6120 6484
rect 6080 6404 6084 6436
rect 6116 6404 6120 6436
rect 6080 6356 6120 6404
rect 6080 6324 6084 6356
rect 6116 6324 6120 6356
rect 6080 5796 6120 6324
rect 6080 5764 6084 5796
rect 6116 5764 6120 5796
rect 6080 5716 6120 5764
rect 6080 5684 6084 5716
rect 6116 5684 6120 5716
rect 6080 5636 6120 5684
rect 6080 5604 6084 5636
rect 6116 5604 6120 5636
rect 6080 5556 6120 5604
rect 6080 5524 6084 5556
rect 6116 5524 6120 5556
rect 6080 5476 6120 5524
rect 6080 5444 6084 5476
rect 6116 5444 6120 5476
rect 6080 5396 6120 5444
rect 6080 5364 6084 5396
rect 6116 5364 6120 5396
rect 6080 5316 6120 5364
rect 6080 5284 6084 5316
rect 6116 5284 6120 5316
rect 6080 5236 6120 5284
rect 6080 5204 6084 5236
rect 6116 5204 6120 5236
rect 6080 5156 6120 5204
rect 6080 5124 6084 5156
rect 6116 5124 6120 5156
rect 6080 5076 6120 5124
rect 6080 5044 6084 5076
rect 6116 5044 6120 5076
rect 6080 4996 6120 5044
rect 6080 4964 6084 4996
rect 6116 4964 6120 4996
rect 6080 4915 6120 4964
rect 6080 4885 6085 4915
rect 6115 4885 6120 4915
rect 6080 4755 6120 4885
rect 6080 4725 6085 4755
rect 6115 4725 6120 4755
rect 6080 4436 6120 4725
rect 6080 4404 6084 4436
rect 6116 4404 6120 4436
rect 6080 4356 6120 4404
rect 6080 4324 6084 4356
rect 6116 4324 6120 4356
rect 6080 4276 6120 4324
rect 6080 4244 6084 4276
rect 6116 4244 6120 4276
rect 6080 4196 6120 4244
rect 6080 4164 6084 4196
rect 6116 4164 6120 4196
rect 6080 4116 6120 4164
rect 6080 4084 6084 4116
rect 6116 4084 6120 4116
rect 6080 4036 6120 4084
rect 6080 4004 6084 4036
rect 6116 4004 6120 4036
rect 6080 3956 6120 4004
rect 6080 3924 6084 3956
rect 6116 3924 6120 3956
rect 6080 3395 6120 3924
rect 6080 3365 6085 3395
rect 6115 3365 6120 3395
rect 6080 3235 6120 3365
rect 6080 3205 6085 3235
rect 6115 3205 6120 3235
rect 6080 3156 6120 3205
rect 6080 3124 6084 3156
rect 6116 3124 6120 3156
rect 6080 3076 6120 3124
rect 6080 3044 6084 3076
rect 6116 3044 6120 3076
rect 6080 2996 6120 3044
rect 6080 2964 6084 2996
rect 6116 2964 6120 2996
rect 6080 2916 6120 2964
rect 6080 2884 6084 2916
rect 6116 2884 6120 2916
rect 6080 2836 6120 2884
rect 6080 2804 6084 2836
rect 6116 2804 6120 2836
rect 6080 2756 6120 2804
rect 6080 2724 6084 2756
rect 6116 2724 6120 2756
rect 6080 2676 6120 2724
rect 6080 2644 6084 2676
rect 6116 2644 6120 2676
rect 6080 2596 6120 2644
rect 6080 2564 6084 2596
rect 6116 2564 6120 2596
rect 6080 2516 6120 2564
rect 6080 2484 6084 2516
rect 6116 2484 6120 2516
rect 6080 2436 6120 2484
rect 6080 2404 6084 2436
rect 6116 2404 6120 2436
rect 6080 2356 6120 2404
rect 6080 2324 6084 2356
rect 6116 2324 6120 2356
rect 6080 2276 6120 2324
rect 6080 2244 6084 2276
rect 6116 2244 6120 2276
rect 6080 2196 6120 2244
rect 6080 2164 6084 2196
rect 6116 2164 6120 2196
rect 6080 2116 6120 2164
rect 6080 2084 6084 2116
rect 6116 2084 6120 2116
rect 6080 2036 6120 2084
rect 6080 2004 6084 2036
rect 6116 2004 6120 2036
rect 6080 1636 6120 2004
rect 6080 1604 6084 1636
rect 6116 1604 6120 1636
rect 6080 1556 6120 1604
rect 6080 1524 6084 1556
rect 6116 1524 6120 1556
rect 6080 1476 6120 1524
rect 6080 1444 6084 1476
rect 6116 1444 6120 1476
rect 6080 1396 6120 1444
rect 6080 1364 6084 1396
rect 6116 1364 6120 1396
rect 6080 1316 6120 1364
rect 6080 1284 6084 1316
rect 6116 1284 6120 1316
rect 6080 1236 6120 1284
rect 6080 1204 6084 1236
rect 6116 1204 6120 1236
rect 6080 1156 6120 1204
rect 6080 1124 6084 1156
rect 6116 1124 6120 1156
rect 6080 1076 6120 1124
rect 6080 1044 6084 1076
rect 6116 1044 6120 1076
rect 6080 756 6120 1044
rect 6080 724 6084 756
rect 6116 724 6120 756
rect 6080 676 6120 724
rect 6080 644 6084 676
rect 6116 644 6120 676
rect 6080 596 6120 644
rect 6080 564 6084 596
rect 6116 564 6120 596
rect 6080 196 6120 564
rect 6080 164 6084 196
rect 6116 164 6120 196
rect 6080 116 6120 164
rect 6080 84 6084 116
rect 6116 84 6120 116
rect 6080 36 6120 84
rect 6080 4 6084 36
rect 6116 4 6120 36
rect 6080 -40 6120 4
rect 6160 12636 6200 13204
rect 6320 13396 6360 13400
rect 6320 13204 6324 13396
rect 6356 13204 6360 13396
rect 6160 12604 6164 12636
rect 6196 12604 6200 12636
rect 6160 12556 6200 12604
rect 6160 12524 6164 12556
rect 6196 12524 6200 12556
rect 6160 12476 6200 12524
rect 6160 12444 6164 12476
rect 6196 12444 6200 12476
rect 6160 12396 6200 12444
rect 6160 12364 6164 12396
rect 6196 12364 6200 12396
rect 6160 12316 6200 12364
rect 6160 12284 6164 12316
rect 6196 12284 6200 12316
rect 6160 12236 6200 12284
rect 6160 12204 6164 12236
rect 6196 12204 6200 12236
rect 6160 12156 6200 12204
rect 6160 12124 6164 12156
rect 6196 12124 6200 12156
rect 6160 11836 6200 12124
rect 6160 11804 6164 11836
rect 6196 11804 6200 11836
rect 6160 11756 6200 11804
rect 6160 11724 6164 11756
rect 6196 11724 6200 11756
rect 6160 11676 6200 11724
rect 6160 11644 6164 11676
rect 6196 11644 6200 11676
rect 6160 11596 6200 11644
rect 6160 11564 6164 11596
rect 6196 11564 6200 11596
rect 6160 11516 6200 11564
rect 6160 11484 6164 11516
rect 6196 11484 6200 11516
rect 6160 11436 6200 11484
rect 6160 11404 6164 11436
rect 6196 11404 6200 11436
rect 6160 10876 6200 11404
rect 6160 10844 6164 10876
rect 6196 10844 6200 10876
rect 6160 10796 6200 10844
rect 6160 10764 6164 10796
rect 6196 10764 6200 10796
rect 6160 10716 6200 10764
rect 6160 10684 6164 10716
rect 6196 10684 6200 10716
rect 6160 10636 6200 10684
rect 6160 10604 6164 10636
rect 6196 10604 6200 10636
rect 6160 10556 6200 10604
rect 6160 10524 6164 10556
rect 6196 10524 6200 10556
rect 6160 10476 6200 10524
rect 6160 10444 6164 10476
rect 6196 10444 6200 10476
rect 6160 10396 6200 10444
rect 6160 10364 6164 10396
rect 6196 10364 6200 10396
rect 6160 10316 6200 10364
rect 6160 10284 6164 10316
rect 6196 10284 6200 10316
rect 6160 10236 6200 10284
rect 6160 10204 6164 10236
rect 6196 10204 6200 10236
rect 6160 10156 6200 10204
rect 6160 10124 6164 10156
rect 6196 10124 6200 10156
rect 6160 10076 6200 10124
rect 6160 10044 6164 10076
rect 6196 10044 6200 10076
rect 6160 9996 6200 10044
rect 6160 9964 6164 9996
rect 6196 9964 6200 9996
rect 6160 9916 6200 9964
rect 6160 9884 6164 9916
rect 6196 9884 6200 9916
rect 6160 9836 6200 9884
rect 6160 9804 6164 9836
rect 6196 9804 6200 9836
rect 6160 9756 6200 9804
rect 6160 9724 6164 9756
rect 6196 9724 6200 9756
rect 6160 9356 6200 9724
rect 6160 9324 6164 9356
rect 6196 9324 6200 9356
rect 6160 9276 6200 9324
rect 6160 9244 6164 9276
rect 6196 9244 6200 9276
rect 6160 9196 6200 9244
rect 6160 9164 6164 9196
rect 6196 9164 6200 9196
rect 6160 8876 6200 9164
rect 6160 8844 6164 8876
rect 6196 8844 6200 8876
rect 6160 8796 6200 8844
rect 6160 8764 6164 8796
rect 6196 8764 6200 8796
rect 6160 8716 6200 8764
rect 6160 8684 6164 8716
rect 6196 8684 6200 8716
rect 6160 8636 6200 8684
rect 6160 8604 6164 8636
rect 6196 8604 6200 8636
rect 6160 8556 6200 8604
rect 6160 8524 6164 8556
rect 6196 8524 6200 8556
rect 6160 7636 6200 8524
rect 6160 7604 6164 7636
rect 6196 7604 6200 7636
rect 6160 7556 6200 7604
rect 6160 7524 6164 7556
rect 6196 7524 6200 7556
rect 6160 7476 6200 7524
rect 6160 7444 6164 7476
rect 6196 7444 6200 7476
rect 6160 7396 6200 7444
rect 6160 7364 6164 7396
rect 6196 7364 6200 7396
rect 6160 7316 6200 7364
rect 6160 7284 6164 7316
rect 6196 7284 6200 7316
rect 6160 7236 6200 7284
rect 6160 7204 6164 7236
rect 6196 7204 6200 7236
rect 6160 7156 6200 7204
rect 6160 7124 6164 7156
rect 6196 7124 6200 7156
rect 6160 7076 6200 7124
rect 6160 7044 6164 7076
rect 6196 7044 6200 7076
rect 6160 6756 6200 7044
rect 6160 6724 6164 6756
rect 6196 6724 6200 6756
rect 6160 6676 6200 6724
rect 6160 6644 6164 6676
rect 6196 6644 6200 6676
rect 6160 6596 6200 6644
rect 6160 6564 6164 6596
rect 6196 6564 6200 6596
rect 6160 6516 6200 6564
rect 6160 6484 6164 6516
rect 6196 6484 6200 6516
rect 6160 6436 6200 6484
rect 6160 6404 6164 6436
rect 6196 6404 6200 6436
rect 6160 6356 6200 6404
rect 6160 6324 6164 6356
rect 6196 6324 6200 6356
rect 6160 5796 6200 6324
rect 6160 5764 6164 5796
rect 6196 5764 6200 5796
rect 6160 5716 6200 5764
rect 6160 5684 6164 5716
rect 6196 5684 6200 5716
rect 6160 5636 6200 5684
rect 6160 5604 6164 5636
rect 6196 5604 6200 5636
rect 6160 5556 6200 5604
rect 6160 5524 6164 5556
rect 6196 5524 6200 5556
rect 6160 5476 6200 5524
rect 6160 5444 6164 5476
rect 6196 5444 6200 5476
rect 6160 5396 6200 5444
rect 6160 5364 6164 5396
rect 6196 5364 6200 5396
rect 6160 5316 6200 5364
rect 6160 5284 6164 5316
rect 6196 5284 6200 5316
rect 6160 5236 6200 5284
rect 6160 5204 6164 5236
rect 6196 5204 6200 5236
rect 6160 5156 6200 5204
rect 6160 5124 6164 5156
rect 6196 5124 6200 5156
rect 6160 5076 6200 5124
rect 6160 5044 6164 5076
rect 6196 5044 6200 5076
rect 6160 4996 6200 5044
rect 6160 4964 6164 4996
rect 6196 4964 6200 4996
rect 6160 4675 6200 4964
rect 6160 4645 6165 4675
rect 6195 4645 6200 4675
rect 6160 4515 6200 4645
rect 6160 4485 6165 4515
rect 6195 4485 6200 4515
rect 6160 4436 6200 4485
rect 6160 4404 6164 4436
rect 6196 4404 6200 4436
rect 6160 4356 6200 4404
rect 6160 4324 6164 4356
rect 6196 4324 6200 4356
rect 6160 4276 6200 4324
rect 6160 4244 6164 4276
rect 6196 4244 6200 4276
rect 6160 4196 6200 4244
rect 6160 4164 6164 4196
rect 6196 4164 6200 4196
rect 6160 4116 6200 4164
rect 6160 4084 6164 4116
rect 6196 4084 6200 4116
rect 6160 4036 6200 4084
rect 6160 4004 6164 4036
rect 6196 4004 6200 4036
rect 6160 3956 6200 4004
rect 6160 3924 6164 3956
rect 6196 3924 6200 3956
rect 6160 3156 6200 3924
rect 6160 3124 6164 3156
rect 6196 3124 6200 3156
rect 6160 3076 6200 3124
rect 6160 3044 6164 3076
rect 6196 3044 6200 3076
rect 6160 2996 6200 3044
rect 6160 2964 6164 2996
rect 6196 2964 6200 2996
rect 6160 2916 6200 2964
rect 6160 2884 6164 2916
rect 6196 2884 6200 2916
rect 6160 2836 6200 2884
rect 6160 2804 6164 2836
rect 6196 2804 6200 2836
rect 6160 2756 6200 2804
rect 6160 2724 6164 2756
rect 6196 2724 6200 2756
rect 6160 2676 6200 2724
rect 6160 2644 6164 2676
rect 6196 2644 6200 2676
rect 6160 2596 6200 2644
rect 6160 2564 6164 2596
rect 6196 2564 6200 2596
rect 6160 2516 6200 2564
rect 6160 2484 6164 2516
rect 6196 2484 6200 2516
rect 6160 2436 6200 2484
rect 6160 2404 6164 2436
rect 6196 2404 6200 2436
rect 6160 2356 6200 2404
rect 6160 2324 6164 2356
rect 6196 2324 6200 2356
rect 6160 2276 6200 2324
rect 6160 2244 6164 2276
rect 6196 2244 6200 2276
rect 6160 2196 6200 2244
rect 6160 2164 6164 2196
rect 6196 2164 6200 2196
rect 6160 2116 6200 2164
rect 6160 2084 6164 2116
rect 6196 2084 6200 2116
rect 6160 2036 6200 2084
rect 6160 2004 6164 2036
rect 6196 2004 6200 2036
rect 6160 1636 6200 2004
rect 6160 1604 6164 1636
rect 6196 1604 6200 1636
rect 6160 1556 6200 1604
rect 6160 1524 6164 1556
rect 6196 1524 6200 1556
rect 6160 1476 6200 1524
rect 6160 1444 6164 1476
rect 6196 1444 6200 1476
rect 6160 1396 6200 1444
rect 6160 1364 6164 1396
rect 6196 1364 6200 1396
rect 6160 1316 6200 1364
rect 6160 1284 6164 1316
rect 6196 1284 6200 1316
rect 6160 1236 6200 1284
rect 6160 1204 6164 1236
rect 6196 1204 6200 1236
rect 6160 1156 6200 1204
rect 6160 1124 6164 1156
rect 6196 1124 6200 1156
rect 6160 1076 6200 1124
rect 6160 1044 6164 1076
rect 6196 1044 6200 1076
rect 6160 995 6200 1044
rect 6160 965 6165 995
rect 6195 965 6200 995
rect 6160 835 6200 965
rect 6160 805 6165 835
rect 6195 805 6200 835
rect 6160 756 6200 805
rect 6160 724 6164 756
rect 6196 724 6200 756
rect 6160 676 6200 724
rect 6160 644 6164 676
rect 6196 644 6200 676
rect 6160 596 6200 644
rect 6160 564 6164 596
rect 6196 564 6200 596
rect 6160 196 6200 564
rect 6160 164 6164 196
rect 6196 164 6200 196
rect 6160 116 6200 164
rect 6160 84 6164 116
rect 6196 84 6200 116
rect 6160 36 6200 84
rect 6160 4 6164 36
rect 6196 4 6200 36
rect 6160 -40 6200 4
rect 6240 4595 6280 12680
rect 6240 4565 6245 4595
rect 6275 4565 6280 4595
rect 6240 915 6280 4565
rect 6240 885 6245 915
rect 6275 885 6280 915
rect 6240 -40 6280 885
rect 6320 12636 6360 13204
rect 6320 12604 6324 12636
rect 6356 12604 6360 12636
rect 6320 12556 6360 12604
rect 6320 12524 6324 12556
rect 6356 12524 6360 12556
rect 6320 12476 6360 12524
rect 6320 12444 6324 12476
rect 6356 12444 6360 12476
rect 6320 12396 6360 12444
rect 6320 12364 6324 12396
rect 6356 12364 6360 12396
rect 6320 12316 6360 12364
rect 6320 12284 6324 12316
rect 6356 12284 6360 12316
rect 6320 12236 6360 12284
rect 6320 12204 6324 12236
rect 6356 12204 6360 12236
rect 6320 12156 6360 12204
rect 6320 12124 6324 12156
rect 6356 12124 6360 12156
rect 6320 11836 6360 12124
rect 6320 11804 6324 11836
rect 6356 11804 6360 11836
rect 6320 11756 6360 11804
rect 6320 11724 6324 11756
rect 6356 11724 6360 11756
rect 6320 11676 6360 11724
rect 6320 11644 6324 11676
rect 6356 11644 6360 11676
rect 6320 11596 6360 11644
rect 6320 11564 6324 11596
rect 6356 11564 6360 11596
rect 6320 11516 6360 11564
rect 6320 11484 6324 11516
rect 6356 11484 6360 11516
rect 6320 11436 6360 11484
rect 6320 11404 6324 11436
rect 6356 11404 6360 11436
rect 6320 10876 6360 11404
rect 6320 10844 6324 10876
rect 6356 10844 6360 10876
rect 6320 10796 6360 10844
rect 6320 10764 6324 10796
rect 6356 10764 6360 10796
rect 6320 10716 6360 10764
rect 6320 10684 6324 10716
rect 6356 10684 6360 10716
rect 6320 10636 6360 10684
rect 6320 10604 6324 10636
rect 6356 10604 6360 10636
rect 6320 10556 6360 10604
rect 6320 10524 6324 10556
rect 6356 10524 6360 10556
rect 6320 10476 6360 10524
rect 6320 10444 6324 10476
rect 6356 10444 6360 10476
rect 6320 10396 6360 10444
rect 6320 10364 6324 10396
rect 6356 10364 6360 10396
rect 6320 10316 6360 10364
rect 6320 10284 6324 10316
rect 6356 10284 6360 10316
rect 6320 10236 6360 10284
rect 6320 10204 6324 10236
rect 6356 10204 6360 10236
rect 6320 10156 6360 10204
rect 6320 10124 6324 10156
rect 6356 10124 6360 10156
rect 6320 10076 6360 10124
rect 6320 10044 6324 10076
rect 6356 10044 6360 10076
rect 6320 9996 6360 10044
rect 6320 9964 6324 9996
rect 6356 9964 6360 9996
rect 6320 9916 6360 9964
rect 6320 9884 6324 9916
rect 6356 9884 6360 9916
rect 6320 9836 6360 9884
rect 6320 9804 6324 9836
rect 6356 9804 6360 9836
rect 6320 9756 6360 9804
rect 6320 9724 6324 9756
rect 6356 9724 6360 9756
rect 6320 9356 6360 9724
rect 6320 9324 6324 9356
rect 6356 9324 6360 9356
rect 6320 9276 6360 9324
rect 6320 9244 6324 9276
rect 6356 9244 6360 9276
rect 6320 9196 6360 9244
rect 6320 9164 6324 9196
rect 6356 9164 6360 9196
rect 6320 8876 6360 9164
rect 6320 8844 6324 8876
rect 6356 8844 6360 8876
rect 6320 8796 6360 8844
rect 6320 8764 6324 8796
rect 6356 8764 6360 8796
rect 6320 8716 6360 8764
rect 6320 8684 6324 8716
rect 6356 8684 6360 8716
rect 6320 8636 6360 8684
rect 6320 8604 6324 8636
rect 6356 8604 6360 8636
rect 6320 8556 6360 8604
rect 6320 8524 6324 8556
rect 6356 8524 6360 8556
rect 6320 7636 6360 8524
rect 6320 7604 6324 7636
rect 6356 7604 6360 7636
rect 6320 7556 6360 7604
rect 6320 7524 6324 7556
rect 6356 7524 6360 7556
rect 6320 7476 6360 7524
rect 6320 7444 6324 7476
rect 6356 7444 6360 7476
rect 6320 7396 6360 7444
rect 6320 7364 6324 7396
rect 6356 7364 6360 7396
rect 6320 7316 6360 7364
rect 6320 7284 6324 7316
rect 6356 7284 6360 7316
rect 6320 7236 6360 7284
rect 6320 7204 6324 7236
rect 6356 7204 6360 7236
rect 6320 7156 6360 7204
rect 6320 7124 6324 7156
rect 6356 7124 6360 7156
rect 6320 7076 6360 7124
rect 6320 7044 6324 7076
rect 6356 7044 6360 7076
rect 6320 6756 6360 7044
rect 6320 6724 6324 6756
rect 6356 6724 6360 6756
rect 6320 6676 6360 6724
rect 6320 6644 6324 6676
rect 6356 6644 6360 6676
rect 6320 6596 6360 6644
rect 6320 6564 6324 6596
rect 6356 6564 6360 6596
rect 6320 6516 6360 6564
rect 6320 6484 6324 6516
rect 6356 6484 6360 6516
rect 6320 6436 6360 6484
rect 6320 6404 6324 6436
rect 6356 6404 6360 6436
rect 6320 6356 6360 6404
rect 6320 6324 6324 6356
rect 6356 6324 6360 6356
rect 6320 5796 6360 6324
rect 6320 5764 6324 5796
rect 6356 5764 6360 5796
rect 6320 5716 6360 5764
rect 6320 5684 6324 5716
rect 6356 5684 6360 5716
rect 6320 5636 6360 5684
rect 6320 5604 6324 5636
rect 6356 5604 6360 5636
rect 6320 5556 6360 5604
rect 6320 5524 6324 5556
rect 6356 5524 6360 5556
rect 6320 5476 6360 5524
rect 6320 5444 6324 5476
rect 6356 5444 6360 5476
rect 6320 5396 6360 5444
rect 6320 5364 6324 5396
rect 6356 5364 6360 5396
rect 6320 5316 6360 5364
rect 6320 5284 6324 5316
rect 6356 5284 6360 5316
rect 6320 5236 6360 5284
rect 6320 5204 6324 5236
rect 6356 5204 6360 5236
rect 6320 5156 6360 5204
rect 6320 5124 6324 5156
rect 6356 5124 6360 5156
rect 6320 5076 6360 5124
rect 6320 5044 6324 5076
rect 6356 5044 6360 5076
rect 6320 4996 6360 5044
rect 6320 4964 6324 4996
rect 6356 4964 6360 4996
rect 6320 4675 6360 4964
rect 6320 4645 6325 4675
rect 6355 4645 6360 4675
rect 6320 4515 6360 4645
rect 6320 4485 6325 4515
rect 6355 4485 6360 4515
rect 6320 4436 6360 4485
rect 6320 4404 6324 4436
rect 6356 4404 6360 4436
rect 6320 4356 6360 4404
rect 6320 4324 6324 4356
rect 6356 4324 6360 4356
rect 6320 4276 6360 4324
rect 6320 4244 6324 4276
rect 6356 4244 6360 4276
rect 6320 4196 6360 4244
rect 6320 4164 6324 4196
rect 6356 4164 6360 4196
rect 6320 4116 6360 4164
rect 6320 4084 6324 4116
rect 6356 4084 6360 4116
rect 6320 4036 6360 4084
rect 6320 4004 6324 4036
rect 6356 4004 6360 4036
rect 6320 3956 6360 4004
rect 6320 3924 6324 3956
rect 6356 3924 6360 3956
rect 6320 3156 6360 3924
rect 6320 3124 6324 3156
rect 6356 3124 6360 3156
rect 6320 3076 6360 3124
rect 6320 3044 6324 3076
rect 6356 3044 6360 3076
rect 6320 2996 6360 3044
rect 6320 2964 6324 2996
rect 6356 2964 6360 2996
rect 6320 2916 6360 2964
rect 6320 2884 6324 2916
rect 6356 2884 6360 2916
rect 6320 2836 6360 2884
rect 6320 2804 6324 2836
rect 6356 2804 6360 2836
rect 6320 2756 6360 2804
rect 6320 2724 6324 2756
rect 6356 2724 6360 2756
rect 6320 2676 6360 2724
rect 6320 2644 6324 2676
rect 6356 2644 6360 2676
rect 6320 2596 6360 2644
rect 6320 2564 6324 2596
rect 6356 2564 6360 2596
rect 6320 2516 6360 2564
rect 6320 2484 6324 2516
rect 6356 2484 6360 2516
rect 6320 2436 6360 2484
rect 6320 2404 6324 2436
rect 6356 2404 6360 2436
rect 6320 2356 6360 2404
rect 6320 2324 6324 2356
rect 6356 2324 6360 2356
rect 6320 2276 6360 2324
rect 6320 2244 6324 2276
rect 6356 2244 6360 2276
rect 6320 2196 6360 2244
rect 6320 2164 6324 2196
rect 6356 2164 6360 2196
rect 6320 2116 6360 2164
rect 6320 2084 6324 2116
rect 6356 2084 6360 2116
rect 6320 2036 6360 2084
rect 6320 2004 6324 2036
rect 6356 2004 6360 2036
rect 6320 1636 6360 2004
rect 6320 1604 6324 1636
rect 6356 1604 6360 1636
rect 6320 1556 6360 1604
rect 6320 1524 6324 1556
rect 6356 1524 6360 1556
rect 6320 1476 6360 1524
rect 6320 1444 6324 1476
rect 6356 1444 6360 1476
rect 6320 1396 6360 1444
rect 6320 1364 6324 1396
rect 6356 1364 6360 1396
rect 6320 1316 6360 1364
rect 6320 1284 6324 1316
rect 6356 1284 6360 1316
rect 6320 1236 6360 1284
rect 6320 1204 6324 1236
rect 6356 1204 6360 1236
rect 6320 1156 6360 1204
rect 6320 1124 6324 1156
rect 6356 1124 6360 1156
rect 6320 1076 6360 1124
rect 6320 1044 6324 1076
rect 6356 1044 6360 1076
rect 6320 995 6360 1044
rect 6320 965 6325 995
rect 6355 965 6360 995
rect 6320 835 6360 965
rect 6320 805 6325 835
rect 6355 805 6360 835
rect 6320 756 6360 805
rect 6320 724 6324 756
rect 6356 724 6360 756
rect 6320 676 6360 724
rect 6320 644 6324 676
rect 6356 644 6360 676
rect 6320 596 6360 644
rect 6320 564 6324 596
rect 6356 564 6360 596
rect 6320 196 6360 564
rect 6320 164 6324 196
rect 6356 164 6360 196
rect 6320 116 6360 164
rect 6320 84 6324 116
rect 6356 84 6360 116
rect 6320 36 6360 84
rect 6320 4 6324 36
rect 6356 4 6360 36
rect 6320 -40 6360 4
<< via3 >>
rect 4 16884 36 16916
rect 4 15444 36 15476
rect 4 14004 36 14036
rect 84 16804 116 16836
rect 84 15524 116 15556
rect 84 13924 116 13956
rect 84 13764 116 13796
rect 164 16724 196 16756
rect 164 13844 196 13876
rect 244 16804 276 16836
rect 244 15524 276 15556
rect 244 13924 276 13956
rect 244 13764 276 13796
rect 324 16884 356 16916
rect 10244 16884 10276 16916
rect 404 16804 436 16836
rect 10164 16804 10196 16836
rect 484 16724 516 16756
rect 1524 16724 1556 16756
rect 1604 16724 1636 16756
rect 2644 16724 2676 16756
rect 2724 16724 2756 16756
rect 3764 16724 3796 16756
rect 3844 16724 3876 16756
rect 4884 16724 4916 16756
rect 5684 16724 5716 16756
rect 6724 16724 6756 16756
rect 6804 16724 6836 16756
rect 7844 16724 7876 16756
rect 7924 16724 7956 16756
rect 8964 16724 8996 16756
rect 9044 16724 9076 16756
rect 10084 16724 10116 16756
rect 404 15524 436 15556
rect 10164 15524 10196 15556
rect 324 15444 356 15476
rect 10244 15444 10276 15476
rect 404 15364 436 15396
rect 4964 15364 4996 15396
rect 484 15284 516 15316
rect 1524 15284 1556 15316
rect 1604 15284 1636 15316
rect 2644 15284 2676 15316
rect 2724 15284 2756 15316
rect 3764 15284 3796 15316
rect 3844 15284 3876 15316
rect 4884 15284 4916 15316
rect 404 14084 436 14116
rect 4964 14084 4996 14116
rect 324 14004 356 14036
rect 4 13684 36 13716
rect 5044 14004 5076 14036
rect 324 13684 356 13716
rect 4484 13924 4516 13956
rect 4484 13764 4516 13796
rect 4244 13444 4276 13636
rect 4404 13444 4436 13636
rect 4244 12635 4276 12636
rect 4244 12605 4245 12635
rect 4245 12605 4275 12635
rect 4275 12605 4276 12635
rect 4244 12604 4276 12605
rect 4244 12555 4276 12556
rect 4244 12525 4245 12555
rect 4245 12525 4275 12555
rect 4275 12525 4276 12555
rect 4244 12524 4276 12525
rect 4244 12475 4276 12476
rect 4244 12445 4245 12475
rect 4245 12445 4275 12475
rect 4275 12445 4276 12475
rect 4244 12444 4276 12445
rect 4244 12395 4276 12396
rect 4244 12365 4245 12395
rect 4245 12365 4275 12395
rect 4275 12365 4276 12395
rect 4244 12364 4276 12365
rect 4244 12315 4276 12316
rect 4244 12285 4245 12315
rect 4245 12285 4275 12315
rect 4275 12285 4276 12315
rect 4244 12284 4276 12285
rect 4244 12235 4276 12236
rect 4244 12205 4245 12235
rect 4245 12205 4275 12235
rect 4275 12205 4276 12235
rect 4244 12204 4276 12205
rect 4244 12155 4276 12156
rect 4244 12125 4245 12155
rect 4245 12125 4275 12155
rect 4275 12125 4276 12155
rect 4244 12124 4276 12125
rect 4244 11835 4276 11836
rect 4244 11805 4245 11835
rect 4245 11805 4275 11835
rect 4275 11805 4276 11835
rect 4244 11804 4276 11805
rect 4244 11755 4276 11756
rect 4244 11725 4245 11755
rect 4245 11725 4275 11755
rect 4275 11725 4276 11755
rect 4244 11724 4276 11725
rect 4244 11675 4276 11676
rect 4244 11645 4245 11675
rect 4245 11645 4275 11675
rect 4275 11645 4276 11675
rect 4244 11644 4276 11645
rect 4244 11595 4276 11596
rect 4244 11565 4245 11595
rect 4245 11565 4275 11595
rect 4275 11565 4276 11595
rect 4244 11564 4276 11565
rect 4244 11515 4276 11516
rect 4244 11485 4245 11515
rect 4245 11485 4275 11515
rect 4275 11485 4276 11515
rect 4244 11484 4276 11485
rect 4244 11435 4276 11436
rect 4244 11405 4245 11435
rect 4245 11405 4275 11435
rect 4275 11405 4276 11435
rect 4244 11404 4276 11405
rect 4244 10875 4276 10876
rect 4244 10845 4245 10875
rect 4245 10845 4275 10875
rect 4275 10845 4276 10875
rect 4244 10844 4276 10845
rect 4244 10795 4276 10796
rect 4244 10765 4245 10795
rect 4245 10765 4275 10795
rect 4275 10765 4276 10795
rect 4244 10764 4276 10765
rect 4244 10715 4276 10716
rect 4244 10685 4245 10715
rect 4245 10685 4275 10715
rect 4275 10685 4276 10715
rect 4244 10684 4276 10685
rect 4244 10635 4276 10636
rect 4244 10605 4245 10635
rect 4245 10605 4275 10635
rect 4275 10605 4276 10635
rect 4244 10604 4276 10605
rect 4244 10555 4276 10556
rect 4244 10525 4245 10555
rect 4245 10525 4275 10555
rect 4275 10525 4276 10555
rect 4244 10524 4276 10525
rect 4244 10475 4276 10476
rect 4244 10445 4245 10475
rect 4245 10445 4275 10475
rect 4275 10445 4276 10475
rect 4244 10444 4276 10445
rect 4244 10395 4276 10396
rect 4244 10365 4245 10395
rect 4245 10365 4275 10395
rect 4275 10365 4276 10395
rect 4244 10364 4276 10365
rect 4244 10315 4276 10316
rect 4244 10285 4245 10315
rect 4245 10285 4275 10315
rect 4275 10285 4276 10315
rect 4244 10284 4276 10285
rect 4244 10235 4276 10236
rect 4244 10205 4245 10235
rect 4245 10205 4275 10235
rect 4275 10205 4276 10235
rect 4244 10204 4276 10205
rect 4244 10155 4276 10156
rect 4244 10125 4245 10155
rect 4245 10125 4275 10155
rect 4275 10125 4276 10155
rect 4244 10124 4276 10125
rect 4244 10075 4276 10076
rect 4244 10045 4245 10075
rect 4245 10045 4275 10075
rect 4275 10045 4276 10075
rect 4244 10044 4276 10045
rect 4244 9995 4276 9996
rect 4244 9965 4245 9995
rect 4245 9965 4275 9995
rect 4275 9965 4276 9995
rect 4244 9964 4276 9965
rect 4244 9915 4276 9916
rect 4244 9885 4245 9915
rect 4245 9885 4275 9915
rect 4275 9885 4276 9915
rect 4244 9884 4276 9885
rect 4244 9835 4276 9836
rect 4244 9805 4245 9835
rect 4245 9805 4275 9835
rect 4275 9805 4276 9835
rect 4244 9804 4276 9805
rect 4244 9755 4276 9756
rect 4244 9725 4245 9755
rect 4245 9725 4275 9755
rect 4275 9725 4276 9755
rect 4244 9724 4276 9725
rect 4244 9355 4276 9356
rect 4244 9325 4245 9355
rect 4245 9325 4275 9355
rect 4275 9325 4276 9355
rect 4244 9324 4276 9325
rect 4244 9275 4276 9276
rect 4244 9245 4245 9275
rect 4245 9245 4275 9275
rect 4275 9245 4276 9275
rect 4244 9244 4276 9245
rect 4244 9195 4276 9196
rect 4244 9165 4245 9195
rect 4245 9165 4275 9195
rect 4275 9165 4276 9195
rect 4244 9164 4276 9165
rect 4244 8875 4276 8876
rect 4244 8845 4245 8875
rect 4245 8845 4275 8875
rect 4275 8845 4276 8875
rect 4244 8844 4276 8845
rect 4244 8795 4276 8796
rect 4244 8765 4245 8795
rect 4245 8765 4275 8795
rect 4275 8765 4276 8795
rect 4244 8764 4276 8765
rect 4244 8715 4276 8716
rect 4244 8685 4245 8715
rect 4245 8685 4275 8715
rect 4275 8685 4276 8715
rect 4244 8684 4276 8685
rect 4244 8635 4276 8636
rect 4244 8605 4245 8635
rect 4245 8605 4275 8635
rect 4275 8605 4276 8635
rect 4244 8604 4276 8605
rect 4244 8555 4276 8556
rect 4244 8525 4245 8555
rect 4245 8525 4275 8555
rect 4275 8525 4276 8555
rect 4244 8524 4276 8525
rect 4244 7635 4276 7636
rect 4244 7605 4245 7635
rect 4245 7605 4275 7635
rect 4275 7605 4276 7635
rect 4244 7604 4276 7605
rect 4244 7555 4276 7556
rect 4244 7525 4245 7555
rect 4245 7525 4275 7555
rect 4275 7525 4276 7555
rect 4244 7524 4276 7525
rect 4244 7475 4276 7476
rect 4244 7445 4245 7475
rect 4245 7445 4275 7475
rect 4275 7445 4276 7475
rect 4244 7444 4276 7445
rect 4244 7395 4276 7396
rect 4244 7365 4245 7395
rect 4245 7365 4275 7395
rect 4275 7365 4276 7395
rect 4244 7364 4276 7365
rect 4244 7315 4276 7316
rect 4244 7285 4245 7315
rect 4245 7285 4275 7315
rect 4275 7285 4276 7315
rect 4244 7284 4276 7285
rect 4244 7235 4276 7236
rect 4244 7205 4245 7235
rect 4245 7205 4275 7235
rect 4275 7205 4276 7235
rect 4244 7204 4276 7205
rect 4244 7155 4276 7156
rect 4244 7125 4245 7155
rect 4245 7125 4275 7155
rect 4275 7125 4276 7155
rect 4244 7124 4276 7125
rect 4244 7075 4276 7076
rect 4244 7045 4245 7075
rect 4245 7045 4275 7075
rect 4275 7045 4276 7075
rect 4244 7044 4276 7045
rect 4244 6755 4276 6756
rect 4244 6725 4245 6755
rect 4245 6725 4275 6755
rect 4275 6725 4276 6755
rect 4244 6724 4276 6725
rect 4244 6675 4276 6676
rect 4244 6645 4245 6675
rect 4245 6645 4275 6675
rect 4275 6645 4276 6675
rect 4244 6644 4276 6645
rect 4244 6595 4276 6596
rect 4244 6565 4245 6595
rect 4245 6565 4275 6595
rect 4275 6565 4276 6595
rect 4244 6564 4276 6565
rect 4244 6515 4276 6516
rect 4244 6485 4245 6515
rect 4245 6485 4275 6515
rect 4275 6485 4276 6515
rect 4244 6484 4276 6485
rect 4244 6435 4276 6436
rect 4244 6405 4245 6435
rect 4245 6405 4275 6435
rect 4275 6405 4276 6435
rect 4244 6404 4276 6405
rect 4244 6355 4276 6356
rect 4244 6325 4245 6355
rect 4245 6325 4275 6355
rect 4275 6325 4276 6355
rect 4244 6324 4276 6325
rect 4244 5795 4276 5796
rect 4244 5765 4245 5795
rect 4245 5765 4275 5795
rect 4275 5765 4276 5795
rect 4244 5764 4276 5765
rect 4244 5715 4276 5716
rect 4244 5685 4245 5715
rect 4245 5685 4275 5715
rect 4275 5685 4276 5715
rect 4244 5684 4276 5685
rect 4244 5635 4276 5636
rect 4244 5605 4245 5635
rect 4245 5605 4275 5635
rect 4275 5605 4276 5635
rect 4244 5604 4276 5605
rect 4244 5555 4276 5556
rect 4244 5525 4245 5555
rect 4245 5525 4275 5555
rect 4275 5525 4276 5555
rect 4244 5524 4276 5525
rect 4244 5475 4276 5476
rect 4244 5445 4245 5475
rect 4245 5445 4275 5475
rect 4275 5445 4276 5475
rect 4244 5444 4276 5445
rect 4244 5395 4276 5396
rect 4244 5365 4245 5395
rect 4245 5365 4275 5395
rect 4275 5365 4276 5395
rect 4244 5364 4276 5365
rect 4244 5315 4276 5316
rect 4244 5285 4245 5315
rect 4245 5285 4275 5315
rect 4275 5285 4276 5315
rect 4244 5284 4276 5285
rect 4244 5235 4276 5236
rect 4244 5205 4245 5235
rect 4245 5205 4275 5235
rect 4275 5205 4276 5235
rect 4244 5204 4276 5205
rect 4244 5155 4276 5156
rect 4244 5125 4245 5155
rect 4245 5125 4275 5155
rect 4275 5125 4276 5155
rect 4244 5124 4276 5125
rect 4244 5075 4276 5076
rect 4244 5045 4245 5075
rect 4245 5045 4275 5075
rect 4275 5045 4276 5075
rect 4244 5044 4276 5045
rect 4244 4995 4276 4996
rect 4244 4965 4245 4995
rect 4245 4965 4275 4995
rect 4275 4965 4276 4995
rect 4244 4964 4276 4965
rect 4244 4435 4276 4436
rect 4244 4405 4245 4435
rect 4245 4405 4275 4435
rect 4275 4405 4276 4435
rect 4244 4404 4276 4405
rect 4244 4355 4276 4356
rect 4244 4325 4245 4355
rect 4245 4325 4275 4355
rect 4275 4325 4276 4355
rect 4244 4324 4276 4325
rect 4244 4275 4276 4276
rect 4244 4245 4245 4275
rect 4245 4245 4275 4275
rect 4275 4245 4276 4275
rect 4244 4244 4276 4245
rect 4244 4195 4276 4196
rect 4244 4165 4245 4195
rect 4245 4165 4275 4195
rect 4275 4165 4276 4195
rect 4244 4164 4276 4165
rect 4244 4115 4276 4116
rect 4244 4085 4245 4115
rect 4245 4085 4275 4115
rect 4275 4085 4276 4115
rect 4244 4084 4276 4085
rect 4244 4035 4276 4036
rect 4244 4005 4245 4035
rect 4245 4005 4275 4035
rect 4275 4005 4276 4035
rect 4244 4004 4276 4005
rect 4244 3955 4276 3956
rect 4244 3925 4245 3955
rect 4245 3925 4275 3955
rect 4275 3925 4276 3955
rect 4244 3924 4276 3925
rect 4244 3155 4276 3156
rect 4244 3125 4245 3155
rect 4245 3125 4275 3155
rect 4275 3125 4276 3155
rect 4244 3124 4276 3125
rect 4244 3075 4276 3076
rect 4244 3045 4245 3075
rect 4245 3045 4275 3075
rect 4275 3045 4276 3075
rect 4244 3044 4276 3045
rect 4244 2995 4276 2996
rect 4244 2965 4245 2995
rect 4245 2965 4275 2995
rect 4275 2965 4276 2995
rect 4244 2964 4276 2965
rect 4244 2915 4276 2916
rect 4244 2885 4245 2915
rect 4245 2885 4275 2915
rect 4275 2885 4276 2915
rect 4244 2884 4276 2885
rect 4244 2835 4276 2836
rect 4244 2805 4245 2835
rect 4245 2805 4275 2835
rect 4275 2805 4276 2835
rect 4244 2804 4276 2805
rect 4244 2755 4276 2756
rect 4244 2725 4245 2755
rect 4245 2725 4275 2755
rect 4275 2725 4276 2755
rect 4244 2724 4276 2725
rect 4244 2675 4276 2676
rect 4244 2645 4245 2675
rect 4245 2645 4275 2675
rect 4275 2645 4276 2675
rect 4244 2644 4276 2645
rect 4244 2595 4276 2596
rect 4244 2565 4245 2595
rect 4245 2565 4275 2595
rect 4275 2565 4276 2595
rect 4244 2564 4276 2565
rect 4244 2515 4276 2516
rect 4244 2485 4245 2515
rect 4245 2485 4275 2515
rect 4275 2485 4276 2515
rect 4244 2484 4276 2485
rect 4244 2435 4276 2436
rect 4244 2405 4245 2435
rect 4245 2405 4275 2435
rect 4275 2405 4276 2435
rect 4244 2404 4276 2405
rect 4244 2355 4276 2356
rect 4244 2325 4245 2355
rect 4245 2325 4275 2355
rect 4275 2325 4276 2355
rect 4244 2324 4276 2325
rect 4244 2275 4276 2276
rect 4244 2245 4245 2275
rect 4245 2245 4275 2275
rect 4275 2245 4276 2275
rect 4244 2244 4276 2245
rect 4244 2195 4276 2196
rect 4244 2165 4245 2195
rect 4245 2165 4275 2195
rect 4275 2165 4276 2195
rect 4244 2164 4276 2165
rect 4244 2115 4276 2116
rect 4244 2085 4245 2115
rect 4245 2085 4275 2115
rect 4275 2085 4276 2115
rect 4244 2084 4276 2085
rect 4244 2035 4276 2036
rect 4244 2005 4245 2035
rect 4245 2005 4275 2035
rect 4275 2005 4276 2035
rect 4244 2004 4276 2005
rect 4244 1635 4276 1636
rect 4244 1605 4245 1635
rect 4245 1605 4275 1635
rect 4275 1605 4276 1635
rect 4244 1604 4276 1605
rect 4244 1555 4276 1556
rect 4244 1525 4245 1555
rect 4245 1525 4275 1555
rect 4275 1525 4276 1555
rect 4244 1524 4276 1525
rect 4244 1475 4276 1476
rect 4244 1445 4245 1475
rect 4245 1445 4275 1475
rect 4275 1445 4276 1475
rect 4244 1444 4276 1445
rect 4244 1395 4276 1396
rect 4244 1365 4245 1395
rect 4245 1365 4275 1395
rect 4275 1365 4276 1395
rect 4244 1364 4276 1365
rect 4244 1315 4276 1316
rect 4244 1285 4245 1315
rect 4245 1285 4275 1315
rect 4275 1285 4276 1315
rect 4244 1284 4276 1285
rect 4244 1235 4276 1236
rect 4244 1205 4245 1235
rect 4245 1205 4275 1235
rect 4275 1205 4276 1235
rect 4244 1204 4276 1205
rect 4244 1155 4276 1156
rect 4244 1125 4245 1155
rect 4245 1125 4275 1155
rect 4275 1125 4276 1155
rect 4244 1124 4276 1125
rect 4244 1075 4276 1076
rect 4244 1045 4245 1075
rect 4245 1045 4275 1075
rect 4275 1045 4276 1075
rect 4244 1044 4276 1045
rect 4244 755 4276 756
rect 4244 725 4245 755
rect 4245 725 4275 755
rect 4275 725 4276 755
rect 4244 724 4276 725
rect 4244 675 4276 676
rect 4244 645 4245 675
rect 4245 645 4275 675
rect 4275 645 4276 675
rect 4244 644 4276 645
rect 4244 595 4276 596
rect 4244 565 4245 595
rect 4245 565 4275 595
rect 4275 565 4276 595
rect 4244 564 4276 565
rect 4244 195 4276 196
rect 4244 165 4245 195
rect 4245 165 4275 195
rect 4275 165 4276 195
rect 4244 164 4276 165
rect 4244 115 4276 116
rect 4244 85 4245 115
rect 4245 85 4275 115
rect 4275 85 4276 115
rect 4244 84 4276 85
rect 4244 35 4276 36
rect 4244 5 4245 35
rect 4245 5 4275 35
rect 4275 5 4276 35
rect 4244 4 4276 5
rect 4404 12635 4436 12636
rect 4404 12605 4405 12635
rect 4405 12605 4435 12635
rect 4435 12605 4436 12635
rect 4404 12604 4436 12605
rect 4404 12555 4436 12556
rect 4404 12525 4405 12555
rect 4405 12525 4435 12555
rect 4435 12525 4436 12555
rect 4404 12524 4436 12525
rect 4404 12475 4436 12476
rect 4404 12445 4405 12475
rect 4405 12445 4435 12475
rect 4435 12445 4436 12475
rect 4404 12444 4436 12445
rect 4404 12395 4436 12396
rect 4404 12365 4405 12395
rect 4405 12365 4435 12395
rect 4435 12365 4436 12395
rect 4404 12364 4436 12365
rect 4404 12315 4436 12316
rect 4404 12285 4405 12315
rect 4405 12285 4435 12315
rect 4435 12285 4436 12315
rect 4404 12284 4436 12285
rect 4404 12235 4436 12236
rect 4404 12205 4405 12235
rect 4405 12205 4435 12235
rect 4435 12205 4436 12235
rect 4404 12204 4436 12205
rect 4404 12155 4436 12156
rect 4404 12125 4405 12155
rect 4405 12125 4435 12155
rect 4435 12125 4436 12155
rect 4404 12124 4436 12125
rect 4404 11835 4436 11836
rect 4404 11805 4405 11835
rect 4405 11805 4435 11835
rect 4435 11805 4436 11835
rect 4404 11804 4436 11805
rect 4404 11755 4436 11756
rect 4404 11725 4405 11755
rect 4405 11725 4435 11755
rect 4435 11725 4436 11755
rect 4404 11724 4436 11725
rect 4404 11675 4436 11676
rect 4404 11645 4405 11675
rect 4405 11645 4435 11675
rect 4435 11645 4436 11675
rect 4404 11644 4436 11645
rect 4404 11595 4436 11596
rect 4404 11565 4405 11595
rect 4405 11565 4435 11595
rect 4435 11565 4436 11595
rect 4404 11564 4436 11565
rect 4404 11515 4436 11516
rect 4404 11485 4405 11515
rect 4405 11485 4435 11515
rect 4435 11485 4436 11515
rect 4404 11484 4436 11485
rect 4404 11435 4436 11436
rect 4404 11405 4405 11435
rect 4405 11405 4435 11435
rect 4435 11405 4436 11435
rect 4404 11404 4436 11405
rect 4404 10875 4436 10876
rect 4404 10845 4405 10875
rect 4405 10845 4435 10875
rect 4435 10845 4436 10875
rect 4404 10844 4436 10845
rect 4404 10795 4436 10796
rect 4404 10765 4405 10795
rect 4405 10765 4435 10795
rect 4435 10765 4436 10795
rect 4404 10764 4436 10765
rect 4404 10715 4436 10716
rect 4404 10685 4405 10715
rect 4405 10685 4435 10715
rect 4435 10685 4436 10715
rect 4404 10684 4436 10685
rect 4404 10635 4436 10636
rect 4404 10605 4405 10635
rect 4405 10605 4435 10635
rect 4435 10605 4436 10635
rect 4404 10604 4436 10605
rect 4404 10555 4436 10556
rect 4404 10525 4405 10555
rect 4405 10525 4435 10555
rect 4435 10525 4436 10555
rect 4404 10524 4436 10525
rect 4404 10475 4436 10476
rect 4404 10445 4405 10475
rect 4405 10445 4435 10475
rect 4435 10445 4436 10475
rect 4404 10444 4436 10445
rect 4404 10395 4436 10396
rect 4404 10365 4405 10395
rect 4405 10365 4435 10395
rect 4435 10365 4436 10395
rect 4404 10364 4436 10365
rect 4404 10315 4436 10316
rect 4404 10285 4405 10315
rect 4405 10285 4435 10315
rect 4435 10285 4436 10315
rect 4404 10284 4436 10285
rect 4404 10235 4436 10236
rect 4404 10205 4405 10235
rect 4405 10205 4435 10235
rect 4435 10205 4436 10235
rect 4404 10204 4436 10205
rect 4404 10155 4436 10156
rect 4404 10125 4405 10155
rect 4405 10125 4435 10155
rect 4435 10125 4436 10155
rect 4404 10124 4436 10125
rect 4404 10075 4436 10076
rect 4404 10045 4405 10075
rect 4405 10045 4435 10075
rect 4435 10045 4436 10075
rect 4404 10044 4436 10045
rect 4404 9995 4436 9996
rect 4404 9965 4405 9995
rect 4405 9965 4435 9995
rect 4435 9965 4436 9995
rect 4404 9964 4436 9965
rect 4404 9915 4436 9916
rect 4404 9885 4405 9915
rect 4405 9885 4435 9915
rect 4435 9885 4436 9915
rect 4404 9884 4436 9885
rect 4404 9835 4436 9836
rect 4404 9805 4405 9835
rect 4405 9805 4435 9835
rect 4435 9805 4436 9835
rect 4404 9804 4436 9805
rect 4404 9755 4436 9756
rect 4404 9725 4405 9755
rect 4405 9725 4435 9755
rect 4435 9725 4436 9755
rect 4404 9724 4436 9725
rect 4404 9355 4436 9356
rect 4404 9325 4405 9355
rect 4405 9325 4435 9355
rect 4435 9325 4436 9355
rect 4404 9324 4436 9325
rect 4404 9275 4436 9276
rect 4404 9245 4405 9275
rect 4405 9245 4435 9275
rect 4435 9245 4436 9275
rect 4404 9244 4436 9245
rect 4404 9195 4436 9196
rect 4404 9165 4405 9195
rect 4405 9165 4435 9195
rect 4435 9165 4436 9195
rect 4404 9164 4436 9165
rect 4404 8875 4436 8876
rect 4404 8845 4405 8875
rect 4405 8845 4435 8875
rect 4435 8845 4436 8875
rect 4404 8844 4436 8845
rect 4404 8795 4436 8796
rect 4404 8765 4405 8795
rect 4405 8765 4435 8795
rect 4435 8765 4436 8795
rect 4404 8764 4436 8765
rect 4404 8715 4436 8716
rect 4404 8685 4405 8715
rect 4405 8685 4435 8715
rect 4435 8685 4436 8715
rect 4404 8684 4436 8685
rect 4404 8635 4436 8636
rect 4404 8605 4405 8635
rect 4405 8605 4435 8635
rect 4435 8605 4436 8635
rect 4404 8604 4436 8605
rect 4404 8555 4436 8556
rect 4404 8525 4405 8555
rect 4405 8525 4435 8555
rect 4435 8525 4436 8555
rect 4404 8524 4436 8525
rect 4404 7635 4436 7636
rect 4404 7605 4405 7635
rect 4405 7605 4435 7635
rect 4435 7605 4436 7635
rect 4404 7604 4436 7605
rect 4404 7555 4436 7556
rect 4404 7525 4405 7555
rect 4405 7525 4435 7555
rect 4435 7525 4436 7555
rect 4404 7524 4436 7525
rect 4404 7475 4436 7476
rect 4404 7445 4405 7475
rect 4405 7445 4435 7475
rect 4435 7445 4436 7475
rect 4404 7444 4436 7445
rect 4404 7395 4436 7396
rect 4404 7365 4405 7395
rect 4405 7365 4435 7395
rect 4435 7365 4436 7395
rect 4404 7364 4436 7365
rect 4404 7315 4436 7316
rect 4404 7285 4405 7315
rect 4405 7285 4435 7315
rect 4435 7285 4436 7315
rect 4404 7284 4436 7285
rect 4404 7235 4436 7236
rect 4404 7205 4405 7235
rect 4405 7205 4435 7235
rect 4435 7205 4436 7235
rect 4404 7204 4436 7205
rect 4404 7155 4436 7156
rect 4404 7125 4405 7155
rect 4405 7125 4435 7155
rect 4435 7125 4436 7155
rect 4404 7124 4436 7125
rect 4404 7075 4436 7076
rect 4404 7045 4405 7075
rect 4405 7045 4435 7075
rect 4435 7045 4436 7075
rect 4404 7044 4436 7045
rect 4404 6755 4436 6756
rect 4404 6725 4405 6755
rect 4405 6725 4435 6755
rect 4435 6725 4436 6755
rect 4404 6724 4436 6725
rect 4404 6675 4436 6676
rect 4404 6645 4405 6675
rect 4405 6645 4435 6675
rect 4435 6645 4436 6675
rect 4404 6644 4436 6645
rect 4404 6595 4436 6596
rect 4404 6565 4405 6595
rect 4405 6565 4435 6595
rect 4435 6565 4436 6595
rect 4404 6564 4436 6565
rect 4404 6515 4436 6516
rect 4404 6485 4405 6515
rect 4405 6485 4435 6515
rect 4435 6485 4436 6515
rect 4404 6484 4436 6485
rect 4404 6435 4436 6436
rect 4404 6405 4405 6435
rect 4405 6405 4435 6435
rect 4435 6405 4436 6435
rect 4404 6404 4436 6405
rect 4404 6355 4436 6356
rect 4404 6325 4405 6355
rect 4405 6325 4435 6355
rect 4435 6325 4436 6355
rect 4404 6324 4436 6325
rect 4404 5795 4436 5796
rect 4404 5765 4405 5795
rect 4405 5765 4435 5795
rect 4435 5765 4436 5795
rect 4404 5764 4436 5765
rect 4404 5715 4436 5716
rect 4404 5685 4405 5715
rect 4405 5685 4435 5715
rect 4435 5685 4436 5715
rect 4404 5684 4436 5685
rect 4404 5635 4436 5636
rect 4404 5605 4405 5635
rect 4405 5605 4435 5635
rect 4435 5605 4436 5635
rect 4404 5604 4436 5605
rect 4404 5555 4436 5556
rect 4404 5525 4405 5555
rect 4405 5525 4435 5555
rect 4435 5525 4436 5555
rect 4404 5524 4436 5525
rect 4404 5475 4436 5476
rect 4404 5445 4405 5475
rect 4405 5445 4435 5475
rect 4435 5445 4436 5475
rect 4404 5444 4436 5445
rect 4404 5395 4436 5396
rect 4404 5365 4405 5395
rect 4405 5365 4435 5395
rect 4435 5365 4436 5395
rect 4404 5364 4436 5365
rect 4404 5315 4436 5316
rect 4404 5285 4405 5315
rect 4405 5285 4435 5315
rect 4435 5285 4436 5315
rect 4404 5284 4436 5285
rect 4404 5235 4436 5236
rect 4404 5205 4405 5235
rect 4405 5205 4435 5235
rect 4435 5205 4436 5235
rect 4404 5204 4436 5205
rect 4404 5155 4436 5156
rect 4404 5125 4405 5155
rect 4405 5125 4435 5155
rect 4435 5125 4436 5155
rect 4404 5124 4436 5125
rect 4404 5075 4436 5076
rect 4404 5045 4405 5075
rect 4405 5045 4435 5075
rect 4435 5045 4436 5075
rect 4404 5044 4436 5045
rect 4404 4995 4436 4996
rect 4404 4965 4405 4995
rect 4405 4965 4435 4995
rect 4435 4965 4436 4995
rect 4404 4964 4436 4965
rect 4404 4435 4436 4436
rect 4404 4405 4405 4435
rect 4405 4405 4435 4435
rect 4435 4405 4436 4435
rect 4404 4404 4436 4405
rect 4404 4355 4436 4356
rect 4404 4325 4405 4355
rect 4405 4325 4435 4355
rect 4435 4325 4436 4355
rect 4404 4324 4436 4325
rect 4404 4275 4436 4276
rect 4404 4245 4405 4275
rect 4405 4245 4435 4275
rect 4435 4245 4436 4275
rect 4404 4244 4436 4245
rect 4404 4195 4436 4196
rect 4404 4165 4405 4195
rect 4405 4165 4435 4195
rect 4435 4165 4436 4195
rect 4404 4164 4436 4165
rect 4404 4115 4436 4116
rect 4404 4085 4405 4115
rect 4405 4085 4435 4115
rect 4435 4085 4436 4115
rect 4404 4084 4436 4085
rect 4404 4035 4436 4036
rect 4404 4005 4405 4035
rect 4405 4005 4435 4035
rect 4435 4005 4436 4035
rect 4404 4004 4436 4005
rect 4404 3955 4436 3956
rect 4404 3925 4405 3955
rect 4405 3925 4435 3955
rect 4435 3925 4436 3955
rect 4404 3924 4436 3925
rect 4404 3155 4436 3156
rect 4404 3125 4405 3155
rect 4405 3125 4435 3155
rect 4435 3125 4436 3155
rect 4404 3124 4436 3125
rect 4404 3075 4436 3076
rect 4404 3045 4405 3075
rect 4405 3045 4435 3075
rect 4435 3045 4436 3075
rect 4404 3044 4436 3045
rect 4404 2995 4436 2996
rect 4404 2965 4405 2995
rect 4405 2965 4435 2995
rect 4435 2965 4436 2995
rect 4404 2964 4436 2965
rect 4404 2915 4436 2916
rect 4404 2885 4405 2915
rect 4405 2885 4435 2915
rect 4435 2885 4436 2915
rect 4404 2884 4436 2885
rect 4404 2835 4436 2836
rect 4404 2805 4405 2835
rect 4405 2805 4435 2835
rect 4435 2805 4436 2835
rect 4404 2804 4436 2805
rect 4404 2755 4436 2756
rect 4404 2725 4405 2755
rect 4405 2725 4435 2755
rect 4435 2725 4436 2755
rect 4404 2724 4436 2725
rect 4404 2675 4436 2676
rect 4404 2645 4405 2675
rect 4405 2645 4435 2675
rect 4435 2645 4436 2675
rect 4404 2644 4436 2645
rect 4404 2595 4436 2596
rect 4404 2565 4405 2595
rect 4405 2565 4435 2595
rect 4435 2565 4436 2595
rect 4404 2564 4436 2565
rect 4404 2515 4436 2516
rect 4404 2485 4405 2515
rect 4405 2485 4435 2515
rect 4435 2485 4436 2515
rect 4404 2484 4436 2485
rect 4404 2435 4436 2436
rect 4404 2405 4405 2435
rect 4405 2405 4435 2435
rect 4435 2405 4436 2435
rect 4404 2404 4436 2405
rect 4404 2355 4436 2356
rect 4404 2325 4405 2355
rect 4405 2325 4435 2355
rect 4435 2325 4436 2355
rect 4404 2324 4436 2325
rect 4404 2275 4436 2276
rect 4404 2245 4405 2275
rect 4405 2245 4435 2275
rect 4435 2245 4436 2275
rect 4404 2244 4436 2245
rect 4404 2195 4436 2196
rect 4404 2165 4405 2195
rect 4405 2165 4435 2195
rect 4435 2165 4436 2195
rect 4404 2164 4436 2165
rect 4404 2115 4436 2116
rect 4404 2085 4405 2115
rect 4405 2085 4435 2115
rect 4435 2085 4436 2115
rect 4404 2084 4436 2085
rect 4404 2035 4436 2036
rect 4404 2005 4405 2035
rect 4405 2005 4435 2035
rect 4435 2005 4436 2035
rect 4404 2004 4436 2005
rect 4404 1635 4436 1636
rect 4404 1605 4405 1635
rect 4405 1605 4435 1635
rect 4435 1605 4436 1635
rect 4404 1604 4436 1605
rect 4404 1555 4436 1556
rect 4404 1525 4405 1555
rect 4405 1525 4435 1555
rect 4435 1525 4436 1555
rect 4404 1524 4436 1525
rect 4404 1475 4436 1476
rect 4404 1445 4405 1475
rect 4405 1445 4435 1475
rect 4435 1445 4436 1475
rect 4404 1444 4436 1445
rect 4404 1395 4436 1396
rect 4404 1365 4405 1395
rect 4405 1365 4435 1395
rect 4435 1365 4436 1395
rect 4404 1364 4436 1365
rect 4404 1315 4436 1316
rect 4404 1285 4405 1315
rect 4405 1285 4435 1315
rect 4435 1285 4436 1315
rect 4404 1284 4436 1285
rect 4404 1235 4436 1236
rect 4404 1205 4405 1235
rect 4405 1205 4435 1235
rect 4435 1205 4436 1235
rect 4404 1204 4436 1205
rect 4404 1155 4436 1156
rect 4404 1125 4405 1155
rect 4405 1125 4435 1155
rect 4435 1125 4436 1155
rect 4404 1124 4436 1125
rect 4404 1075 4436 1076
rect 4404 1045 4405 1075
rect 4405 1045 4435 1075
rect 4435 1045 4436 1075
rect 4404 1044 4436 1045
rect 4404 755 4436 756
rect 4404 725 4405 755
rect 4405 725 4435 755
rect 4435 725 4436 755
rect 4404 724 4436 725
rect 4404 675 4436 676
rect 4404 645 4405 675
rect 4405 645 4435 675
rect 4435 645 4436 675
rect 4404 644 4436 645
rect 4404 595 4436 596
rect 4404 565 4405 595
rect 4405 565 4435 595
rect 4435 565 4436 595
rect 4404 564 4436 565
rect 4404 195 4436 196
rect 4404 165 4405 195
rect 4405 165 4435 195
rect 4435 165 4436 195
rect 4404 164 4436 165
rect 4404 115 4436 116
rect 4404 85 4405 115
rect 4405 85 4435 115
rect 4435 85 4436 115
rect 4404 84 4436 85
rect 4404 35 4436 36
rect 4404 5 4405 35
rect 4405 5 4435 35
rect 4435 5 4436 35
rect 4404 4 4436 5
rect 4484 12964 4516 13156
rect 4484 12635 4516 12636
rect 4484 12605 4485 12635
rect 4485 12605 4515 12635
rect 4515 12605 4516 12635
rect 4484 12604 4516 12605
rect 4484 12555 4516 12556
rect 4484 12525 4485 12555
rect 4485 12525 4515 12555
rect 4515 12525 4516 12555
rect 4484 12524 4516 12525
rect 4484 12475 4516 12476
rect 4484 12445 4485 12475
rect 4485 12445 4515 12475
rect 4515 12445 4516 12475
rect 4484 12444 4516 12445
rect 4484 12395 4516 12396
rect 4484 12365 4485 12395
rect 4485 12365 4515 12395
rect 4515 12365 4516 12395
rect 4484 12364 4516 12365
rect 4484 12315 4516 12316
rect 4484 12285 4485 12315
rect 4485 12285 4515 12315
rect 4515 12285 4516 12315
rect 4484 12284 4516 12285
rect 4484 12235 4516 12236
rect 4484 12205 4485 12235
rect 4485 12205 4515 12235
rect 4515 12205 4516 12235
rect 4484 12204 4516 12205
rect 4484 12155 4516 12156
rect 4484 12125 4485 12155
rect 4485 12125 4515 12155
rect 4515 12125 4516 12155
rect 4484 12124 4516 12125
rect 4484 11835 4516 11836
rect 4484 11805 4485 11835
rect 4485 11805 4515 11835
rect 4515 11805 4516 11835
rect 4484 11804 4516 11805
rect 4484 11755 4516 11756
rect 4484 11725 4485 11755
rect 4485 11725 4515 11755
rect 4515 11725 4516 11755
rect 4484 11724 4516 11725
rect 4484 11675 4516 11676
rect 4484 11645 4485 11675
rect 4485 11645 4515 11675
rect 4515 11645 4516 11675
rect 4484 11644 4516 11645
rect 4484 11595 4516 11596
rect 4484 11565 4485 11595
rect 4485 11565 4515 11595
rect 4515 11565 4516 11595
rect 4484 11564 4516 11565
rect 4484 11515 4516 11516
rect 4484 11485 4485 11515
rect 4485 11485 4515 11515
rect 4515 11485 4516 11515
rect 4484 11484 4516 11485
rect 4484 11435 4516 11436
rect 4484 11405 4485 11435
rect 4485 11405 4515 11435
rect 4515 11405 4516 11435
rect 4484 11404 4516 11405
rect 4484 10875 4516 10876
rect 4484 10845 4485 10875
rect 4485 10845 4515 10875
rect 4515 10845 4516 10875
rect 4484 10844 4516 10845
rect 4484 10795 4516 10796
rect 4484 10765 4485 10795
rect 4485 10765 4515 10795
rect 4515 10765 4516 10795
rect 4484 10764 4516 10765
rect 4484 10715 4516 10716
rect 4484 10685 4485 10715
rect 4485 10685 4515 10715
rect 4515 10685 4516 10715
rect 4484 10684 4516 10685
rect 4484 10635 4516 10636
rect 4484 10605 4485 10635
rect 4485 10605 4515 10635
rect 4515 10605 4516 10635
rect 4484 10604 4516 10605
rect 4484 10555 4516 10556
rect 4484 10525 4485 10555
rect 4485 10525 4515 10555
rect 4515 10525 4516 10555
rect 4484 10524 4516 10525
rect 4484 10475 4516 10476
rect 4484 10445 4485 10475
rect 4485 10445 4515 10475
rect 4515 10445 4516 10475
rect 4484 10444 4516 10445
rect 4484 10395 4516 10396
rect 4484 10365 4485 10395
rect 4485 10365 4515 10395
rect 4515 10365 4516 10395
rect 4484 10364 4516 10365
rect 4484 10315 4516 10316
rect 4484 10285 4485 10315
rect 4485 10285 4515 10315
rect 4515 10285 4516 10315
rect 4484 10284 4516 10285
rect 4484 10235 4516 10236
rect 4484 10205 4485 10235
rect 4485 10205 4515 10235
rect 4515 10205 4516 10235
rect 4484 10204 4516 10205
rect 4484 10155 4516 10156
rect 4484 10125 4485 10155
rect 4485 10125 4515 10155
rect 4515 10125 4516 10155
rect 4484 10124 4516 10125
rect 4484 10075 4516 10076
rect 4484 10045 4485 10075
rect 4485 10045 4515 10075
rect 4515 10045 4516 10075
rect 4484 10044 4516 10045
rect 4484 9995 4516 9996
rect 4484 9965 4485 9995
rect 4485 9965 4515 9995
rect 4515 9965 4516 9995
rect 4484 9964 4516 9965
rect 4484 9915 4516 9916
rect 4484 9885 4485 9915
rect 4485 9885 4515 9915
rect 4515 9885 4516 9915
rect 4484 9884 4516 9885
rect 4484 9835 4516 9836
rect 4484 9805 4485 9835
rect 4485 9805 4515 9835
rect 4515 9805 4516 9835
rect 4484 9804 4516 9805
rect 4484 9755 4516 9756
rect 4484 9725 4485 9755
rect 4485 9725 4515 9755
rect 4515 9725 4516 9755
rect 4484 9724 4516 9725
rect 4484 9355 4516 9356
rect 4484 9325 4485 9355
rect 4485 9325 4515 9355
rect 4515 9325 4516 9355
rect 4484 9324 4516 9325
rect 4484 9275 4516 9276
rect 4484 9245 4485 9275
rect 4485 9245 4515 9275
rect 4515 9245 4516 9275
rect 4484 9244 4516 9245
rect 4484 9195 4516 9196
rect 4484 9165 4485 9195
rect 4485 9165 4515 9195
rect 4515 9165 4516 9195
rect 4484 9164 4516 9165
rect 4484 8875 4516 8876
rect 4484 8845 4485 8875
rect 4485 8845 4515 8875
rect 4515 8845 4516 8875
rect 4484 8844 4516 8845
rect 4484 8795 4516 8796
rect 4484 8765 4485 8795
rect 4485 8765 4515 8795
rect 4515 8765 4516 8795
rect 4484 8764 4516 8765
rect 4484 8715 4516 8716
rect 4484 8685 4485 8715
rect 4485 8685 4515 8715
rect 4515 8685 4516 8715
rect 4484 8684 4516 8685
rect 4484 8635 4516 8636
rect 4484 8605 4485 8635
rect 4485 8605 4515 8635
rect 4515 8605 4516 8635
rect 4484 8604 4516 8605
rect 4484 8555 4516 8556
rect 4484 8525 4485 8555
rect 4485 8525 4515 8555
rect 4515 8525 4516 8555
rect 4484 8524 4516 8525
rect 4484 7635 4516 7636
rect 4484 7605 4485 7635
rect 4485 7605 4515 7635
rect 4515 7605 4516 7635
rect 4484 7604 4516 7605
rect 4484 7555 4516 7556
rect 4484 7525 4485 7555
rect 4485 7525 4515 7555
rect 4515 7525 4516 7555
rect 4484 7524 4516 7525
rect 4484 7475 4516 7476
rect 4484 7445 4485 7475
rect 4485 7445 4515 7475
rect 4515 7445 4516 7475
rect 4484 7444 4516 7445
rect 4484 7395 4516 7396
rect 4484 7365 4485 7395
rect 4485 7365 4515 7395
rect 4515 7365 4516 7395
rect 4484 7364 4516 7365
rect 4484 7315 4516 7316
rect 4484 7285 4485 7315
rect 4485 7285 4515 7315
rect 4515 7285 4516 7315
rect 4484 7284 4516 7285
rect 4484 7235 4516 7236
rect 4484 7205 4485 7235
rect 4485 7205 4515 7235
rect 4515 7205 4516 7235
rect 4484 7204 4516 7205
rect 4484 7155 4516 7156
rect 4484 7125 4485 7155
rect 4485 7125 4515 7155
rect 4515 7125 4516 7155
rect 4484 7124 4516 7125
rect 4484 7075 4516 7076
rect 4484 7045 4485 7075
rect 4485 7045 4515 7075
rect 4515 7045 4516 7075
rect 4484 7044 4516 7045
rect 4484 6755 4516 6756
rect 4484 6725 4485 6755
rect 4485 6725 4515 6755
rect 4515 6725 4516 6755
rect 4484 6724 4516 6725
rect 4484 6675 4516 6676
rect 4484 6645 4485 6675
rect 4485 6645 4515 6675
rect 4515 6645 4516 6675
rect 4484 6644 4516 6645
rect 4484 6595 4516 6596
rect 4484 6565 4485 6595
rect 4485 6565 4515 6595
rect 4515 6565 4516 6595
rect 4484 6564 4516 6565
rect 4484 6515 4516 6516
rect 4484 6485 4485 6515
rect 4485 6485 4515 6515
rect 4515 6485 4516 6515
rect 4484 6484 4516 6485
rect 4484 6435 4516 6436
rect 4484 6405 4485 6435
rect 4485 6405 4515 6435
rect 4515 6405 4516 6435
rect 4484 6404 4516 6405
rect 4484 6355 4516 6356
rect 4484 6325 4485 6355
rect 4485 6325 4515 6355
rect 4515 6325 4516 6355
rect 4484 6324 4516 6325
rect 4484 5795 4516 5796
rect 4484 5765 4485 5795
rect 4485 5765 4515 5795
rect 4515 5765 4516 5795
rect 4484 5764 4516 5765
rect 4484 5715 4516 5716
rect 4484 5685 4485 5715
rect 4485 5685 4515 5715
rect 4515 5685 4516 5715
rect 4484 5684 4516 5685
rect 4484 5635 4516 5636
rect 4484 5605 4485 5635
rect 4485 5605 4515 5635
rect 4515 5605 4516 5635
rect 4484 5604 4516 5605
rect 4484 5555 4516 5556
rect 4484 5525 4485 5555
rect 4485 5525 4515 5555
rect 4515 5525 4516 5555
rect 4484 5524 4516 5525
rect 4484 5475 4516 5476
rect 4484 5445 4485 5475
rect 4485 5445 4515 5475
rect 4515 5445 4516 5475
rect 4484 5444 4516 5445
rect 4484 5395 4516 5396
rect 4484 5365 4485 5395
rect 4485 5365 4515 5395
rect 4515 5365 4516 5395
rect 4484 5364 4516 5365
rect 4484 5315 4516 5316
rect 4484 5285 4485 5315
rect 4485 5285 4515 5315
rect 4515 5285 4516 5315
rect 4484 5284 4516 5285
rect 4484 5235 4516 5236
rect 4484 5205 4485 5235
rect 4485 5205 4515 5235
rect 4515 5205 4516 5235
rect 4484 5204 4516 5205
rect 4484 5155 4516 5156
rect 4484 5125 4485 5155
rect 4485 5125 4515 5155
rect 4515 5125 4516 5155
rect 4484 5124 4516 5125
rect 4484 5075 4516 5076
rect 4484 5045 4485 5075
rect 4485 5045 4515 5075
rect 4515 5045 4516 5075
rect 4484 5044 4516 5045
rect 4484 4995 4516 4996
rect 4484 4965 4485 4995
rect 4485 4965 4515 4995
rect 4515 4965 4516 4995
rect 4484 4964 4516 4965
rect 4484 4435 4516 4436
rect 4484 4405 4485 4435
rect 4485 4405 4515 4435
rect 4515 4405 4516 4435
rect 4484 4404 4516 4405
rect 4484 4355 4516 4356
rect 4484 4325 4485 4355
rect 4485 4325 4515 4355
rect 4515 4325 4516 4355
rect 4484 4324 4516 4325
rect 4484 4275 4516 4276
rect 4484 4245 4485 4275
rect 4485 4245 4515 4275
rect 4515 4245 4516 4275
rect 4484 4244 4516 4245
rect 4484 4195 4516 4196
rect 4484 4165 4485 4195
rect 4485 4165 4515 4195
rect 4515 4165 4516 4195
rect 4484 4164 4516 4165
rect 4484 4115 4516 4116
rect 4484 4085 4485 4115
rect 4485 4085 4515 4115
rect 4515 4085 4516 4115
rect 4484 4084 4516 4085
rect 4484 4035 4516 4036
rect 4484 4005 4485 4035
rect 4485 4005 4515 4035
rect 4515 4005 4516 4035
rect 4484 4004 4516 4005
rect 4484 3955 4516 3956
rect 4484 3925 4485 3955
rect 4485 3925 4515 3955
rect 4515 3925 4516 3955
rect 4484 3924 4516 3925
rect 4484 3155 4516 3156
rect 4484 3125 4485 3155
rect 4485 3125 4515 3155
rect 4515 3125 4516 3155
rect 4484 3124 4516 3125
rect 4484 3075 4516 3076
rect 4484 3045 4485 3075
rect 4485 3045 4515 3075
rect 4515 3045 4516 3075
rect 4484 3044 4516 3045
rect 4484 2995 4516 2996
rect 4484 2965 4485 2995
rect 4485 2965 4515 2995
rect 4515 2965 4516 2995
rect 4484 2964 4516 2965
rect 4484 2915 4516 2916
rect 4484 2885 4485 2915
rect 4485 2885 4515 2915
rect 4515 2885 4516 2915
rect 4484 2884 4516 2885
rect 4484 2835 4516 2836
rect 4484 2805 4485 2835
rect 4485 2805 4515 2835
rect 4515 2805 4516 2835
rect 4484 2804 4516 2805
rect 4484 2755 4516 2756
rect 4484 2725 4485 2755
rect 4485 2725 4515 2755
rect 4515 2725 4516 2755
rect 4484 2724 4516 2725
rect 4484 2675 4516 2676
rect 4484 2645 4485 2675
rect 4485 2645 4515 2675
rect 4515 2645 4516 2675
rect 4484 2644 4516 2645
rect 4484 2595 4516 2596
rect 4484 2565 4485 2595
rect 4485 2565 4515 2595
rect 4515 2565 4516 2595
rect 4484 2564 4516 2565
rect 4484 2515 4516 2516
rect 4484 2485 4485 2515
rect 4485 2485 4515 2515
rect 4515 2485 4516 2515
rect 4484 2484 4516 2485
rect 4484 2435 4516 2436
rect 4484 2405 4485 2435
rect 4485 2405 4515 2435
rect 4515 2405 4516 2435
rect 4484 2404 4516 2405
rect 4484 2355 4516 2356
rect 4484 2325 4485 2355
rect 4485 2325 4515 2355
rect 4515 2325 4516 2355
rect 4484 2324 4516 2325
rect 4484 2275 4516 2276
rect 4484 2245 4485 2275
rect 4485 2245 4515 2275
rect 4515 2245 4516 2275
rect 4484 2244 4516 2245
rect 4484 2195 4516 2196
rect 4484 2165 4485 2195
rect 4485 2165 4515 2195
rect 4515 2165 4516 2195
rect 4484 2164 4516 2165
rect 4484 2115 4516 2116
rect 4484 2085 4485 2115
rect 4485 2085 4515 2115
rect 4515 2085 4516 2115
rect 4484 2084 4516 2085
rect 4484 2035 4516 2036
rect 4484 2005 4485 2035
rect 4485 2005 4515 2035
rect 4515 2005 4516 2035
rect 4484 2004 4516 2005
rect 4484 1635 4516 1636
rect 4484 1605 4485 1635
rect 4485 1605 4515 1635
rect 4515 1605 4516 1635
rect 4484 1604 4516 1605
rect 4484 1555 4516 1556
rect 4484 1525 4485 1555
rect 4485 1525 4515 1555
rect 4515 1525 4516 1555
rect 4484 1524 4516 1525
rect 4484 1475 4516 1476
rect 4484 1445 4485 1475
rect 4485 1445 4515 1475
rect 4515 1445 4516 1475
rect 4484 1444 4516 1445
rect 4484 1395 4516 1396
rect 4484 1365 4485 1395
rect 4485 1365 4515 1395
rect 4515 1365 4516 1395
rect 4484 1364 4516 1365
rect 4484 1315 4516 1316
rect 4484 1285 4485 1315
rect 4485 1285 4515 1315
rect 4515 1285 4516 1315
rect 4484 1284 4516 1285
rect 4484 1235 4516 1236
rect 4484 1205 4485 1235
rect 4485 1205 4515 1235
rect 4515 1205 4516 1235
rect 4484 1204 4516 1205
rect 4484 1155 4516 1156
rect 4484 1125 4485 1155
rect 4485 1125 4515 1155
rect 4515 1125 4516 1155
rect 4484 1124 4516 1125
rect 4484 1075 4516 1076
rect 4484 1045 4485 1075
rect 4485 1045 4515 1075
rect 4515 1045 4516 1075
rect 4484 1044 4516 1045
rect 4484 755 4516 756
rect 4484 725 4485 755
rect 4485 725 4515 755
rect 4515 725 4516 755
rect 4484 724 4516 725
rect 4484 675 4516 676
rect 4484 645 4485 675
rect 4485 645 4515 675
rect 4515 645 4516 675
rect 4484 644 4516 645
rect 4484 595 4516 596
rect 4484 565 4485 595
rect 4485 565 4515 595
rect 4515 565 4516 595
rect 4484 564 4516 565
rect 4484 195 4516 196
rect 4484 165 4485 195
rect 4485 165 4515 195
rect 4515 165 4516 195
rect 4484 164 4516 165
rect 4484 115 4516 116
rect 4484 85 4485 115
rect 4485 85 4515 115
rect 4515 85 4516 115
rect 4484 84 4516 85
rect 4484 35 4516 36
rect 4484 5 4485 35
rect 4485 5 4515 35
rect 4515 5 4516 35
rect 4484 4 4516 5
rect 4564 13844 4596 13876
rect 4644 13924 4676 13956
rect 4644 13764 4676 13796
rect 5044 13684 5076 13716
rect 4644 12964 4676 13156
rect 4644 12635 4676 12636
rect 4644 12605 4645 12635
rect 4645 12605 4675 12635
rect 4675 12605 4676 12635
rect 4644 12604 4676 12605
rect 4644 12555 4676 12556
rect 4644 12525 4645 12555
rect 4645 12525 4675 12555
rect 4675 12525 4676 12555
rect 4644 12524 4676 12525
rect 4644 12475 4676 12476
rect 4644 12445 4645 12475
rect 4645 12445 4675 12475
rect 4675 12445 4676 12475
rect 4644 12444 4676 12445
rect 4644 12395 4676 12396
rect 4644 12365 4645 12395
rect 4645 12365 4675 12395
rect 4675 12365 4676 12395
rect 4644 12364 4676 12365
rect 4644 12315 4676 12316
rect 4644 12285 4645 12315
rect 4645 12285 4675 12315
rect 4675 12285 4676 12315
rect 4644 12284 4676 12285
rect 4644 12235 4676 12236
rect 4644 12205 4645 12235
rect 4645 12205 4675 12235
rect 4675 12205 4676 12235
rect 4644 12204 4676 12205
rect 4644 12155 4676 12156
rect 4644 12125 4645 12155
rect 4645 12125 4675 12155
rect 4675 12125 4676 12155
rect 4644 12124 4676 12125
rect 4644 11835 4676 11836
rect 4644 11805 4645 11835
rect 4645 11805 4675 11835
rect 4675 11805 4676 11835
rect 4644 11804 4676 11805
rect 4644 11755 4676 11756
rect 4644 11725 4645 11755
rect 4645 11725 4675 11755
rect 4675 11725 4676 11755
rect 4644 11724 4676 11725
rect 4644 11675 4676 11676
rect 4644 11645 4645 11675
rect 4645 11645 4675 11675
rect 4675 11645 4676 11675
rect 4644 11644 4676 11645
rect 4644 11595 4676 11596
rect 4644 11565 4645 11595
rect 4645 11565 4675 11595
rect 4675 11565 4676 11595
rect 4644 11564 4676 11565
rect 4644 11515 4676 11516
rect 4644 11485 4645 11515
rect 4645 11485 4675 11515
rect 4675 11485 4676 11515
rect 4644 11484 4676 11485
rect 4644 11435 4676 11436
rect 4644 11405 4645 11435
rect 4645 11405 4675 11435
rect 4675 11405 4676 11435
rect 4644 11404 4676 11405
rect 4644 10875 4676 10876
rect 4644 10845 4645 10875
rect 4645 10845 4675 10875
rect 4675 10845 4676 10875
rect 4644 10844 4676 10845
rect 4644 10795 4676 10796
rect 4644 10765 4645 10795
rect 4645 10765 4675 10795
rect 4675 10765 4676 10795
rect 4644 10764 4676 10765
rect 4644 10715 4676 10716
rect 4644 10685 4645 10715
rect 4645 10685 4675 10715
rect 4675 10685 4676 10715
rect 4644 10684 4676 10685
rect 4644 10635 4676 10636
rect 4644 10605 4645 10635
rect 4645 10605 4675 10635
rect 4675 10605 4676 10635
rect 4644 10604 4676 10605
rect 4644 10555 4676 10556
rect 4644 10525 4645 10555
rect 4645 10525 4675 10555
rect 4675 10525 4676 10555
rect 4644 10524 4676 10525
rect 4644 10475 4676 10476
rect 4644 10445 4645 10475
rect 4645 10445 4675 10475
rect 4675 10445 4676 10475
rect 4644 10444 4676 10445
rect 4644 10395 4676 10396
rect 4644 10365 4645 10395
rect 4645 10365 4675 10395
rect 4675 10365 4676 10395
rect 4644 10364 4676 10365
rect 4644 10315 4676 10316
rect 4644 10285 4645 10315
rect 4645 10285 4675 10315
rect 4675 10285 4676 10315
rect 4644 10284 4676 10285
rect 4644 10235 4676 10236
rect 4644 10205 4645 10235
rect 4645 10205 4675 10235
rect 4675 10205 4676 10235
rect 4644 10204 4676 10205
rect 4644 10155 4676 10156
rect 4644 10125 4645 10155
rect 4645 10125 4675 10155
rect 4675 10125 4676 10155
rect 4644 10124 4676 10125
rect 4644 10075 4676 10076
rect 4644 10045 4645 10075
rect 4645 10045 4675 10075
rect 4675 10045 4676 10075
rect 4644 10044 4676 10045
rect 4644 9995 4676 9996
rect 4644 9965 4645 9995
rect 4645 9965 4675 9995
rect 4675 9965 4676 9995
rect 4644 9964 4676 9965
rect 4644 9915 4676 9916
rect 4644 9885 4645 9915
rect 4645 9885 4675 9915
rect 4675 9885 4676 9915
rect 4644 9884 4676 9885
rect 4644 9835 4676 9836
rect 4644 9805 4645 9835
rect 4645 9805 4675 9835
rect 4675 9805 4676 9835
rect 4644 9804 4676 9805
rect 4644 9755 4676 9756
rect 4644 9725 4645 9755
rect 4645 9725 4675 9755
rect 4675 9725 4676 9755
rect 4644 9724 4676 9725
rect 4644 9355 4676 9356
rect 4644 9325 4645 9355
rect 4645 9325 4675 9355
rect 4675 9325 4676 9355
rect 4644 9324 4676 9325
rect 4644 9275 4676 9276
rect 4644 9245 4645 9275
rect 4645 9245 4675 9275
rect 4675 9245 4676 9275
rect 4644 9244 4676 9245
rect 4644 9195 4676 9196
rect 4644 9165 4645 9195
rect 4645 9165 4675 9195
rect 4675 9165 4676 9195
rect 4644 9164 4676 9165
rect 4644 8875 4676 8876
rect 4644 8845 4645 8875
rect 4645 8845 4675 8875
rect 4675 8845 4676 8875
rect 4644 8844 4676 8845
rect 4644 8795 4676 8796
rect 4644 8765 4645 8795
rect 4645 8765 4675 8795
rect 4675 8765 4676 8795
rect 4644 8764 4676 8765
rect 4644 8715 4676 8716
rect 4644 8685 4645 8715
rect 4645 8685 4675 8715
rect 4675 8685 4676 8715
rect 4644 8684 4676 8685
rect 4644 8635 4676 8636
rect 4644 8605 4645 8635
rect 4645 8605 4675 8635
rect 4675 8605 4676 8635
rect 4644 8604 4676 8605
rect 4644 8555 4676 8556
rect 4644 8525 4645 8555
rect 4645 8525 4675 8555
rect 4675 8525 4676 8555
rect 4644 8524 4676 8525
rect 4644 7635 4676 7636
rect 4644 7605 4645 7635
rect 4645 7605 4675 7635
rect 4675 7605 4676 7635
rect 4644 7604 4676 7605
rect 4644 7555 4676 7556
rect 4644 7525 4645 7555
rect 4645 7525 4675 7555
rect 4675 7525 4676 7555
rect 4644 7524 4676 7525
rect 4644 7475 4676 7476
rect 4644 7445 4645 7475
rect 4645 7445 4675 7475
rect 4675 7445 4676 7475
rect 4644 7444 4676 7445
rect 4644 7395 4676 7396
rect 4644 7365 4645 7395
rect 4645 7365 4675 7395
rect 4675 7365 4676 7395
rect 4644 7364 4676 7365
rect 4644 7315 4676 7316
rect 4644 7285 4645 7315
rect 4645 7285 4675 7315
rect 4675 7285 4676 7315
rect 4644 7284 4676 7285
rect 4644 7235 4676 7236
rect 4644 7205 4645 7235
rect 4645 7205 4675 7235
rect 4675 7205 4676 7235
rect 4644 7204 4676 7205
rect 4644 7155 4676 7156
rect 4644 7125 4645 7155
rect 4645 7125 4675 7155
rect 4675 7125 4676 7155
rect 4644 7124 4676 7125
rect 4644 7075 4676 7076
rect 4644 7045 4645 7075
rect 4645 7045 4675 7075
rect 4675 7045 4676 7075
rect 4644 7044 4676 7045
rect 4644 6755 4676 6756
rect 4644 6725 4645 6755
rect 4645 6725 4675 6755
rect 4675 6725 4676 6755
rect 4644 6724 4676 6725
rect 4644 6675 4676 6676
rect 4644 6645 4645 6675
rect 4645 6645 4675 6675
rect 4675 6645 4676 6675
rect 4644 6644 4676 6645
rect 4644 6595 4676 6596
rect 4644 6565 4645 6595
rect 4645 6565 4675 6595
rect 4675 6565 4676 6595
rect 4644 6564 4676 6565
rect 4644 6515 4676 6516
rect 4644 6485 4645 6515
rect 4645 6485 4675 6515
rect 4675 6485 4676 6515
rect 4644 6484 4676 6485
rect 4644 6435 4676 6436
rect 4644 6405 4645 6435
rect 4645 6405 4675 6435
rect 4675 6405 4676 6435
rect 4644 6404 4676 6405
rect 4644 6355 4676 6356
rect 4644 6325 4645 6355
rect 4645 6325 4675 6355
rect 4675 6325 4676 6355
rect 4644 6324 4676 6325
rect 4644 5795 4676 5796
rect 4644 5765 4645 5795
rect 4645 5765 4675 5795
rect 4675 5765 4676 5795
rect 4644 5764 4676 5765
rect 4644 5715 4676 5716
rect 4644 5685 4645 5715
rect 4645 5685 4675 5715
rect 4675 5685 4676 5715
rect 4644 5684 4676 5685
rect 4644 5635 4676 5636
rect 4644 5605 4645 5635
rect 4645 5605 4675 5635
rect 4675 5605 4676 5635
rect 4644 5604 4676 5605
rect 4644 5555 4676 5556
rect 4644 5525 4645 5555
rect 4645 5525 4675 5555
rect 4675 5525 4676 5555
rect 4644 5524 4676 5525
rect 4644 5475 4676 5476
rect 4644 5445 4645 5475
rect 4645 5445 4675 5475
rect 4675 5445 4676 5475
rect 4644 5444 4676 5445
rect 4644 5395 4676 5396
rect 4644 5365 4645 5395
rect 4645 5365 4675 5395
rect 4675 5365 4676 5395
rect 4644 5364 4676 5365
rect 4644 5315 4676 5316
rect 4644 5285 4645 5315
rect 4645 5285 4675 5315
rect 4675 5285 4676 5315
rect 4644 5284 4676 5285
rect 4644 5235 4676 5236
rect 4644 5205 4645 5235
rect 4645 5205 4675 5235
rect 4675 5205 4676 5235
rect 4644 5204 4676 5205
rect 4644 5155 4676 5156
rect 4644 5125 4645 5155
rect 4645 5125 4675 5155
rect 4675 5125 4676 5155
rect 4644 5124 4676 5125
rect 4644 5075 4676 5076
rect 4644 5045 4645 5075
rect 4645 5045 4675 5075
rect 4675 5045 4676 5075
rect 4644 5044 4676 5045
rect 4644 4995 4676 4996
rect 4644 4965 4645 4995
rect 4645 4965 4675 4995
rect 4675 4965 4676 4995
rect 4644 4964 4676 4965
rect 4644 4435 4676 4436
rect 4644 4405 4645 4435
rect 4645 4405 4675 4435
rect 4675 4405 4676 4435
rect 4644 4404 4676 4405
rect 4644 4355 4676 4356
rect 4644 4325 4645 4355
rect 4645 4325 4675 4355
rect 4675 4325 4676 4355
rect 4644 4324 4676 4325
rect 4644 4275 4676 4276
rect 4644 4245 4645 4275
rect 4645 4245 4675 4275
rect 4675 4245 4676 4275
rect 4644 4244 4676 4245
rect 4644 4195 4676 4196
rect 4644 4165 4645 4195
rect 4645 4165 4675 4195
rect 4675 4165 4676 4195
rect 4644 4164 4676 4165
rect 4644 4115 4676 4116
rect 4644 4085 4645 4115
rect 4645 4085 4675 4115
rect 4675 4085 4676 4115
rect 4644 4084 4676 4085
rect 4644 4035 4676 4036
rect 4644 4005 4645 4035
rect 4645 4005 4675 4035
rect 4675 4005 4676 4035
rect 4644 4004 4676 4005
rect 4644 3955 4676 3956
rect 4644 3925 4645 3955
rect 4645 3925 4675 3955
rect 4675 3925 4676 3955
rect 4644 3924 4676 3925
rect 4644 3155 4676 3156
rect 4644 3125 4645 3155
rect 4645 3125 4675 3155
rect 4675 3125 4676 3155
rect 4644 3124 4676 3125
rect 4644 3075 4676 3076
rect 4644 3045 4645 3075
rect 4645 3045 4675 3075
rect 4675 3045 4676 3075
rect 4644 3044 4676 3045
rect 4644 2995 4676 2996
rect 4644 2965 4645 2995
rect 4645 2965 4675 2995
rect 4675 2965 4676 2995
rect 4644 2964 4676 2965
rect 4644 2915 4676 2916
rect 4644 2885 4645 2915
rect 4645 2885 4675 2915
rect 4675 2885 4676 2915
rect 4644 2884 4676 2885
rect 4644 2835 4676 2836
rect 4644 2805 4645 2835
rect 4645 2805 4675 2835
rect 4675 2805 4676 2835
rect 4644 2804 4676 2805
rect 4644 2755 4676 2756
rect 4644 2725 4645 2755
rect 4645 2725 4675 2755
rect 4675 2725 4676 2755
rect 4644 2724 4676 2725
rect 4644 2675 4676 2676
rect 4644 2645 4645 2675
rect 4645 2645 4675 2675
rect 4675 2645 4676 2675
rect 4644 2644 4676 2645
rect 4644 2595 4676 2596
rect 4644 2565 4645 2595
rect 4645 2565 4675 2595
rect 4675 2565 4676 2595
rect 4644 2564 4676 2565
rect 4644 2515 4676 2516
rect 4644 2485 4645 2515
rect 4645 2485 4675 2515
rect 4675 2485 4676 2515
rect 4644 2484 4676 2485
rect 4644 2435 4676 2436
rect 4644 2405 4645 2435
rect 4645 2405 4675 2435
rect 4675 2405 4676 2435
rect 4644 2404 4676 2405
rect 4644 2355 4676 2356
rect 4644 2325 4645 2355
rect 4645 2325 4675 2355
rect 4675 2325 4676 2355
rect 4644 2324 4676 2325
rect 4644 2275 4676 2276
rect 4644 2245 4645 2275
rect 4645 2245 4675 2275
rect 4675 2245 4676 2275
rect 4644 2244 4676 2245
rect 4644 2195 4676 2196
rect 4644 2165 4645 2195
rect 4645 2165 4675 2195
rect 4675 2165 4676 2195
rect 4644 2164 4676 2165
rect 4644 2115 4676 2116
rect 4644 2085 4645 2115
rect 4645 2085 4675 2115
rect 4675 2085 4676 2115
rect 4644 2084 4676 2085
rect 4644 2035 4676 2036
rect 4644 2005 4645 2035
rect 4645 2005 4675 2035
rect 4675 2005 4676 2035
rect 4644 2004 4676 2005
rect 4644 1635 4676 1636
rect 4644 1605 4645 1635
rect 4645 1605 4675 1635
rect 4675 1605 4676 1635
rect 4644 1604 4676 1605
rect 4644 1555 4676 1556
rect 4644 1525 4645 1555
rect 4645 1525 4675 1555
rect 4675 1525 4676 1555
rect 4644 1524 4676 1525
rect 4644 1475 4676 1476
rect 4644 1445 4645 1475
rect 4645 1445 4675 1475
rect 4675 1445 4676 1475
rect 4644 1444 4676 1445
rect 4644 1395 4676 1396
rect 4644 1365 4645 1395
rect 4645 1365 4675 1395
rect 4675 1365 4676 1395
rect 4644 1364 4676 1365
rect 4644 1315 4676 1316
rect 4644 1285 4645 1315
rect 4645 1285 4675 1315
rect 4675 1285 4676 1315
rect 4644 1284 4676 1285
rect 4644 1235 4676 1236
rect 4644 1205 4645 1235
rect 4645 1205 4675 1235
rect 4675 1205 4676 1235
rect 4644 1204 4676 1205
rect 4644 1155 4676 1156
rect 4644 1125 4645 1155
rect 4645 1125 4675 1155
rect 4675 1125 4676 1155
rect 4644 1124 4676 1125
rect 4644 1075 4676 1076
rect 4644 1045 4645 1075
rect 4645 1045 4675 1075
rect 4675 1045 4676 1075
rect 4644 1044 4676 1045
rect 4644 755 4676 756
rect 4644 725 4645 755
rect 4645 725 4675 755
rect 4675 725 4676 755
rect 4644 724 4676 725
rect 4644 675 4676 676
rect 4644 645 4645 675
rect 4645 645 4675 675
rect 4675 645 4676 675
rect 4644 644 4676 645
rect 4644 595 4676 596
rect 4644 565 4645 595
rect 4645 565 4675 595
rect 4675 565 4676 595
rect 4644 564 4676 565
rect 4644 195 4676 196
rect 4644 165 4645 195
rect 4645 165 4675 195
rect 4675 165 4676 195
rect 4644 164 4676 165
rect 4644 115 4676 116
rect 4644 85 4645 115
rect 4645 85 4675 115
rect 4675 85 4676 115
rect 4644 84 4676 85
rect 4644 35 4676 36
rect 4644 5 4645 35
rect 4645 5 4675 35
rect 4675 5 4676 35
rect 4644 4 4676 5
rect 4724 13204 4756 13396
rect 4884 13204 4916 13396
rect 4724 12635 4756 12636
rect 4724 12605 4725 12635
rect 4725 12605 4755 12635
rect 4755 12605 4756 12635
rect 4724 12604 4756 12605
rect 4724 12555 4756 12556
rect 4724 12525 4725 12555
rect 4725 12525 4755 12555
rect 4755 12525 4756 12555
rect 4724 12524 4756 12525
rect 4724 12475 4756 12476
rect 4724 12445 4725 12475
rect 4725 12445 4755 12475
rect 4755 12445 4756 12475
rect 4724 12444 4756 12445
rect 4724 12395 4756 12396
rect 4724 12365 4725 12395
rect 4725 12365 4755 12395
rect 4755 12365 4756 12395
rect 4724 12364 4756 12365
rect 4724 12315 4756 12316
rect 4724 12285 4725 12315
rect 4725 12285 4755 12315
rect 4755 12285 4756 12315
rect 4724 12284 4756 12285
rect 4724 12235 4756 12236
rect 4724 12205 4725 12235
rect 4725 12205 4755 12235
rect 4755 12205 4756 12235
rect 4724 12204 4756 12205
rect 4724 12155 4756 12156
rect 4724 12125 4725 12155
rect 4725 12125 4755 12155
rect 4755 12125 4756 12155
rect 4724 12124 4756 12125
rect 4724 11835 4756 11836
rect 4724 11805 4725 11835
rect 4725 11805 4755 11835
rect 4755 11805 4756 11835
rect 4724 11804 4756 11805
rect 4724 11755 4756 11756
rect 4724 11725 4725 11755
rect 4725 11725 4755 11755
rect 4755 11725 4756 11755
rect 4724 11724 4756 11725
rect 4724 11675 4756 11676
rect 4724 11645 4725 11675
rect 4725 11645 4755 11675
rect 4755 11645 4756 11675
rect 4724 11644 4756 11645
rect 4724 11595 4756 11596
rect 4724 11565 4725 11595
rect 4725 11565 4755 11595
rect 4755 11565 4756 11595
rect 4724 11564 4756 11565
rect 4724 11515 4756 11516
rect 4724 11485 4725 11515
rect 4725 11485 4755 11515
rect 4755 11485 4756 11515
rect 4724 11484 4756 11485
rect 4724 11435 4756 11436
rect 4724 11405 4725 11435
rect 4725 11405 4755 11435
rect 4755 11405 4756 11435
rect 4724 11404 4756 11405
rect 4724 10875 4756 10876
rect 4724 10845 4725 10875
rect 4725 10845 4755 10875
rect 4755 10845 4756 10875
rect 4724 10844 4756 10845
rect 4724 10795 4756 10796
rect 4724 10765 4725 10795
rect 4725 10765 4755 10795
rect 4755 10765 4756 10795
rect 4724 10764 4756 10765
rect 4724 10715 4756 10716
rect 4724 10685 4725 10715
rect 4725 10685 4755 10715
rect 4755 10685 4756 10715
rect 4724 10684 4756 10685
rect 4724 10635 4756 10636
rect 4724 10605 4725 10635
rect 4725 10605 4755 10635
rect 4755 10605 4756 10635
rect 4724 10604 4756 10605
rect 4724 10555 4756 10556
rect 4724 10525 4725 10555
rect 4725 10525 4755 10555
rect 4755 10525 4756 10555
rect 4724 10524 4756 10525
rect 4724 10475 4756 10476
rect 4724 10445 4725 10475
rect 4725 10445 4755 10475
rect 4755 10445 4756 10475
rect 4724 10444 4756 10445
rect 4724 10395 4756 10396
rect 4724 10365 4725 10395
rect 4725 10365 4755 10395
rect 4755 10365 4756 10395
rect 4724 10364 4756 10365
rect 4724 10315 4756 10316
rect 4724 10285 4725 10315
rect 4725 10285 4755 10315
rect 4755 10285 4756 10315
rect 4724 10284 4756 10285
rect 4724 10235 4756 10236
rect 4724 10205 4725 10235
rect 4725 10205 4755 10235
rect 4755 10205 4756 10235
rect 4724 10204 4756 10205
rect 4724 10155 4756 10156
rect 4724 10125 4725 10155
rect 4725 10125 4755 10155
rect 4755 10125 4756 10155
rect 4724 10124 4756 10125
rect 4724 10075 4756 10076
rect 4724 10045 4725 10075
rect 4725 10045 4755 10075
rect 4755 10045 4756 10075
rect 4724 10044 4756 10045
rect 4724 9995 4756 9996
rect 4724 9965 4725 9995
rect 4725 9965 4755 9995
rect 4755 9965 4756 9995
rect 4724 9964 4756 9965
rect 4724 9915 4756 9916
rect 4724 9885 4725 9915
rect 4725 9885 4755 9915
rect 4755 9885 4756 9915
rect 4724 9884 4756 9885
rect 4724 9835 4756 9836
rect 4724 9805 4725 9835
rect 4725 9805 4755 9835
rect 4755 9805 4756 9835
rect 4724 9804 4756 9805
rect 4724 9755 4756 9756
rect 4724 9725 4725 9755
rect 4725 9725 4755 9755
rect 4755 9725 4756 9755
rect 4724 9724 4756 9725
rect 4724 9355 4756 9356
rect 4724 9325 4725 9355
rect 4725 9325 4755 9355
rect 4755 9325 4756 9355
rect 4724 9324 4756 9325
rect 4724 9275 4756 9276
rect 4724 9245 4725 9275
rect 4725 9245 4755 9275
rect 4755 9245 4756 9275
rect 4724 9244 4756 9245
rect 4724 9195 4756 9196
rect 4724 9165 4725 9195
rect 4725 9165 4755 9195
rect 4755 9165 4756 9195
rect 4724 9164 4756 9165
rect 4724 8875 4756 8876
rect 4724 8845 4725 8875
rect 4725 8845 4755 8875
rect 4755 8845 4756 8875
rect 4724 8844 4756 8845
rect 4724 8795 4756 8796
rect 4724 8765 4725 8795
rect 4725 8765 4755 8795
rect 4755 8765 4756 8795
rect 4724 8764 4756 8765
rect 4724 8715 4756 8716
rect 4724 8685 4725 8715
rect 4725 8685 4755 8715
rect 4755 8685 4756 8715
rect 4724 8684 4756 8685
rect 4724 8635 4756 8636
rect 4724 8605 4725 8635
rect 4725 8605 4755 8635
rect 4755 8605 4756 8635
rect 4724 8604 4756 8605
rect 4724 8555 4756 8556
rect 4724 8525 4725 8555
rect 4725 8525 4755 8555
rect 4755 8525 4756 8555
rect 4724 8524 4756 8525
rect 4724 7635 4756 7636
rect 4724 7605 4725 7635
rect 4725 7605 4755 7635
rect 4755 7605 4756 7635
rect 4724 7604 4756 7605
rect 4724 7555 4756 7556
rect 4724 7525 4725 7555
rect 4725 7525 4755 7555
rect 4755 7525 4756 7555
rect 4724 7524 4756 7525
rect 4724 7475 4756 7476
rect 4724 7445 4725 7475
rect 4725 7445 4755 7475
rect 4755 7445 4756 7475
rect 4724 7444 4756 7445
rect 4724 7395 4756 7396
rect 4724 7365 4725 7395
rect 4725 7365 4755 7395
rect 4755 7365 4756 7395
rect 4724 7364 4756 7365
rect 4724 7315 4756 7316
rect 4724 7285 4725 7315
rect 4725 7285 4755 7315
rect 4755 7285 4756 7315
rect 4724 7284 4756 7285
rect 4724 7235 4756 7236
rect 4724 7205 4725 7235
rect 4725 7205 4755 7235
rect 4755 7205 4756 7235
rect 4724 7204 4756 7205
rect 4724 7155 4756 7156
rect 4724 7125 4725 7155
rect 4725 7125 4755 7155
rect 4755 7125 4756 7155
rect 4724 7124 4756 7125
rect 4724 7075 4756 7076
rect 4724 7045 4725 7075
rect 4725 7045 4755 7075
rect 4755 7045 4756 7075
rect 4724 7044 4756 7045
rect 4724 6755 4756 6756
rect 4724 6725 4725 6755
rect 4725 6725 4755 6755
rect 4755 6725 4756 6755
rect 4724 6724 4756 6725
rect 4724 6675 4756 6676
rect 4724 6645 4725 6675
rect 4725 6645 4755 6675
rect 4755 6645 4756 6675
rect 4724 6644 4756 6645
rect 4724 6595 4756 6596
rect 4724 6565 4725 6595
rect 4725 6565 4755 6595
rect 4755 6565 4756 6595
rect 4724 6564 4756 6565
rect 4724 6515 4756 6516
rect 4724 6485 4725 6515
rect 4725 6485 4755 6515
rect 4755 6485 4756 6515
rect 4724 6484 4756 6485
rect 4724 6435 4756 6436
rect 4724 6405 4725 6435
rect 4725 6405 4755 6435
rect 4755 6405 4756 6435
rect 4724 6404 4756 6405
rect 4724 6355 4756 6356
rect 4724 6325 4725 6355
rect 4725 6325 4755 6355
rect 4755 6325 4756 6355
rect 4724 6324 4756 6325
rect 4724 5795 4756 5796
rect 4724 5765 4725 5795
rect 4725 5765 4755 5795
rect 4755 5765 4756 5795
rect 4724 5764 4756 5765
rect 4724 5715 4756 5716
rect 4724 5685 4725 5715
rect 4725 5685 4755 5715
rect 4755 5685 4756 5715
rect 4724 5684 4756 5685
rect 4724 5635 4756 5636
rect 4724 5605 4725 5635
rect 4725 5605 4755 5635
rect 4755 5605 4756 5635
rect 4724 5604 4756 5605
rect 4724 5555 4756 5556
rect 4724 5525 4725 5555
rect 4725 5525 4755 5555
rect 4755 5525 4756 5555
rect 4724 5524 4756 5525
rect 4724 5475 4756 5476
rect 4724 5445 4725 5475
rect 4725 5445 4755 5475
rect 4755 5445 4756 5475
rect 4724 5444 4756 5445
rect 4724 5395 4756 5396
rect 4724 5365 4725 5395
rect 4725 5365 4755 5395
rect 4755 5365 4756 5395
rect 4724 5364 4756 5365
rect 4724 5315 4756 5316
rect 4724 5285 4725 5315
rect 4725 5285 4755 5315
rect 4755 5285 4756 5315
rect 4724 5284 4756 5285
rect 4724 5235 4756 5236
rect 4724 5205 4725 5235
rect 4725 5205 4755 5235
rect 4755 5205 4756 5235
rect 4724 5204 4756 5205
rect 4724 5155 4756 5156
rect 4724 5125 4725 5155
rect 4725 5125 4755 5155
rect 4755 5125 4756 5155
rect 4724 5124 4756 5125
rect 4724 5075 4756 5076
rect 4724 5045 4725 5075
rect 4725 5045 4755 5075
rect 4755 5045 4756 5075
rect 4724 5044 4756 5045
rect 4724 4995 4756 4996
rect 4724 4965 4725 4995
rect 4725 4965 4755 4995
rect 4755 4965 4756 4995
rect 4724 4964 4756 4965
rect 4724 4435 4756 4436
rect 4724 4405 4725 4435
rect 4725 4405 4755 4435
rect 4755 4405 4756 4435
rect 4724 4404 4756 4405
rect 4724 4355 4756 4356
rect 4724 4325 4725 4355
rect 4725 4325 4755 4355
rect 4755 4325 4756 4355
rect 4724 4324 4756 4325
rect 4724 4275 4756 4276
rect 4724 4245 4725 4275
rect 4725 4245 4755 4275
rect 4755 4245 4756 4275
rect 4724 4244 4756 4245
rect 4724 4195 4756 4196
rect 4724 4165 4725 4195
rect 4725 4165 4755 4195
rect 4755 4165 4756 4195
rect 4724 4164 4756 4165
rect 4724 4115 4756 4116
rect 4724 4085 4725 4115
rect 4725 4085 4755 4115
rect 4755 4085 4756 4115
rect 4724 4084 4756 4085
rect 4724 4035 4756 4036
rect 4724 4005 4725 4035
rect 4725 4005 4755 4035
rect 4755 4005 4756 4035
rect 4724 4004 4756 4005
rect 4724 3955 4756 3956
rect 4724 3925 4725 3955
rect 4725 3925 4755 3955
rect 4755 3925 4756 3955
rect 4724 3924 4756 3925
rect 4724 3155 4756 3156
rect 4724 3125 4725 3155
rect 4725 3125 4755 3155
rect 4755 3125 4756 3155
rect 4724 3124 4756 3125
rect 4724 3075 4756 3076
rect 4724 3045 4725 3075
rect 4725 3045 4755 3075
rect 4755 3045 4756 3075
rect 4724 3044 4756 3045
rect 4724 2995 4756 2996
rect 4724 2965 4725 2995
rect 4725 2965 4755 2995
rect 4755 2965 4756 2995
rect 4724 2964 4756 2965
rect 4724 2915 4756 2916
rect 4724 2885 4725 2915
rect 4725 2885 4755 2915
rect 4755 2885 4756 2915
rect 4724 2884 4756 2885
rect 4724 2835 4756 2836
rect 4724 2805 4725 2835
rect 4725 2805 4755 2835
rect 4755 2805 4756 2835
rect 4724 2804 4756 2805
rect 4724 2755 4756 2756
rect 4724 2725 4725 2755
rect 4725 2725 4755 2755
rect 4755 2725 4756 2755
rect 4724 2724 4756 2725
rect 4724 2675 4756 2676
rect 4724 2645 4725 2675
rect 4725 2645 4755 2675
rect 4755 2645 4756 2675
rect 4724 2644 4756 2645
rect 4724 2595 4756 2596
rect 4724 2565 4725 2595
rect 4725 2565 4755 2595
rect 4755 2565 4756 2595
rect 4724 2564 4756 2565
rect 4724 2515 4756 2516
rect 4724 2485 4725 2515
rect 4725 2485 4755 2515
rect 4755 2485 4756 2515
rect 4724 2484 4756 2485
rect 4724 2435 4756 2436
rect 4724 2405 4725 2435
rect 4725 2405 4755 2435
rect 4755 2405 4756 2435
rect 4724 2404 4756 2405
rect 4724 2355 4756 2356
rect 4724 2325 4725 2355
rect 4725 2325 4755 2355
rect 4755 2325 4756 2355
rect 4724 2324 4756 2325
rect 4724 2275 4756 2276
rect 4724 2245 4725 2275
rect 4725 2245 4755 2275
rect 4755 2245 4756 2275
rect 4724 2244 4756 2245
rect 4724 2195 4756 2196
rect 4724 2165 4725 2195
rect 4725 2165 4755 2195
rect 4755 2165 4756 2195
rect 4724 2164 4756 2165
rect 4724 2115 4756 2116
rect 4724 2085 4725 2115
rect 4725 2085 4755 2115
rect 4755 2085 4756 2115
rect 4724 2084 4756 2085
rect 4724 2035 4756 2036
rect 4724 2005 4725 2035
rect 4725 2005 4755 2035
rect 4755 2005 4756 2035
rect 4724 2004 4756 2005
rect 4724 1635 4756 1636
rect 4724 1605 4725 1635
rect 4725 1605 4755 1635
rect 4755 1605 4756 1635
rect 4724 1604 4756 1605
rect 4724 1555 4756 1556
rect 4724 1525 4725 1555
rect 4725 1525 4755 1555
rect 4755 1525 4756 1555
rect 4724 1524 4756 1525
rect 4724 1475 4756 1476
rect 4724 1445 4725 1475
rect 4725 1445 4755 1475
rect 4755 1445 4756 1475
rect 4724 1444 4756 1445
rect 4724 1395 4756 1396
rect 4724 1365 4725 1395
rect 4725 1365 4755 1395
rect 4755 1365 4756 1395
rect 4724 1364 4756 1365
rect 4724 1315 4756 1316
rect 4724 1285 4725 1315
rect 4725 1285 4755 1315
rect 4755 1285 4756 1315
rect 4724 1284 4756 1285
rect 4724 1235 4756 1236
rect 4724 1205 4725 1235
rect 4725 1205 4755 1235
rect 4755 1205 4756 1235
rect 4724 1204 4756 1205
rect 4724 1155 4756 1156
rect 4724 1125 4725 1155
rect 4725 1125 4755 1155
rect 4755 1125 4756 1155
rect 4724 1124 4756 1125
rect 4724 1075 4756 1076
rect 4724 1045 4725 1075
rect 4725 1045 4755 1075
rect 4755 1045 4756 1075
rect 4724 1044 4756 1045
rect 4724 755 4756 756
rect 4724 725 4725 755
rect 4725 725 4755 755
rect 4755 725 4756 755
rect 4724 724 4756 725
rect 4724 675 4756 676
rect 4724 645 4725 675
rect 4725 645 4755 675
rect 4755 645 4756 675
rect 4724 644 4756 645
rect 4724 595 4756 596
rect 4724 565 4725 595
rect 4725 565 4755 595
rect 4755 565 4756 595
rect 4724 564 4756 565
rect 4724 195 4756 196
rect 4724 165 4725 195
rect 4725 165 4755 195
rect 4755 165 4756 195
rect 4724 164 4756 165
rect 4724 115 4756 116
rect 4724 85 4725 115
rect 4725 85 4755 115
rect 4755 85 4756 115
rect 4724 84 4756 85
rect 4724 35 4756 36
rect 4724 5 4725 35
rect 4725 5 4755 35
rect 4755 5 4756 35
rect 4724 4 4756 5
rect 5044 13204 5076 13396
rect 4884 12635 4916 12636
rect 4884 12605 4885 12635
rect 4885 12605 4915 12635
rect 4915 12605 4916 12635
rect 4884 12604 4916 12605
rect 4884 12555 4916 12556
rect 4884 12525 4885 12555
rect 4885 12525 4915 12555
rect 4915 12525 4916 12555
rect 4884 12524 4916 12525
rect 4884 12475 4916 12476
rect 4884 12445 4885 12475
rect 4885 12445 4915 12475
rect 4915 12445 4916 12475
rect 4884 12444 4916 12445
rect 4884 12395 4916 12396
rect 4884 12365 4885 12395
rect 4885 12365 4915 12395
rect 4915 12365 4916 12395
rect 4884 12364 4916 12365
rect 4884 12315 4916 12316
rect 4884 12285 4885 12315
rect 4885 12285 4915 12315
rect 4915 12285 4916 12315
rect 4884 12284 4916 12285
rect 4884 12235 4916 12236
rect 4884 12205 4885 12235
rect 4885 12205 4915 12235
rect 4915 12205 4916 12235
rect 4884 12204 4916 12205
rect 4884 12155 4916 12156
rect 4884 12125 4885 12155
rect 4885 12125 4915 12155
rect 4915 12125 4916 12155
rect 4884 12124 4916 12125
rect 4884 11835 4916 11836
rect 4884 11805 4885 11835
rect 4885 11805 4915 11835
rect 4915 11805 4916 11835
rect 4884 11804 4916 11805
rect 4884 11755 4916 11756
rect 4884 11725 4885 11755
rect 4885 11725 4915 11755
rect 4915 11725 4916 11755
rect 4884 11724 4916 11725
rect 4884 11675 4916 11676
rect 4884 11645 4885 11675
rect 4885 11645 4915 11675
rect 4915 11645 4916 11675
rect 4884 11644 4916 11645
rect 4884 11595 4916 11596
rect 4884 11565 4885 11595
rect 4885 11565 4915 11595
rect 4915 11565 4916 11595
rect 4884 11564 4916 11565
rect 4884 11515 4916 11516
rect 4884 11485 4885 11515
rect 4885 11485 4915 11515
rect 4915 11485 4916 11515
rect 4884 11484 4916 11485
rect 4884 11435 4916 11436
rect 4884 11405 4885 11435
rect 4885 11405 4915 11435
rect 4915 11405 4916 11435
rect 4884 11404 4916 11405
rect 4884 10875 4916 10876
rect 4884 10845 4885 10875
rect 4885 10845 4915 10875
rect 4915 10845 4916 10875
rect 4884 10844 4916 10845
rect 4884 10795 4916 10796
rect 4884 10765 4885 10795
rect 4885 10765 4915 10795
rect 4915 10765 4916 10795
rect 4884 10764 4916 10765
rect 4884 10715 4916 10716
rect 4884 10685 4885 10715
rect 4885 10685 4915 10715
rect 4915 10685 4916 10715
rect 4884 10684 4916 10685
rect 4884 10635 4916 10636
rect 4884 10605 4885 10635
rect 4885 10605 4915 10635
rect 4915 10605 4916 10635
rect 4884 10604 4916 10605
rect 4884 10555 4916 10556
rect 4884 10525 4885 10555
rect 4885 10525 4915 10555
rect 4915 10525 4916 10555
rect 4884 10524 4916 10525
rect 4884 10475 4916 10476
rect 4884 10445 4885 10475
rect 4885 10445 4915 10475
rect 4915 10445 4916 10475
rect 4884 10444 4916 10445
rect 4884 10395 4916 10396
rect 4884 10365 4885 10395
rect 4885 10365 4915 10395
rect 4915 10365 4916 10395
rect 4884 10364 4916 10365
rect 4884 10315 4916 10316
rect 4884 10285 4885 10315
rect 4885 10285 4915 10315
rect 4915 10285 4916 10315
rect 4884 10284 4916 10285
rect 4884 10235 4916 10236
rect 4884 10205 4885 10235
rect 4885 10205 4915 10235
rect 4915 10205 4916 10235
rect 4884 10204 4916 10205
rect 4884 10155 4916 10156
rect 4884 10125 4885 10155
rect 4885 10125 4915 10155
rect 4915 10125 4916 10155
rect 4884 10124 4916 10125
rect 4884 10075 4916 10076
rect 4884 10045 4885 10075
rect 4885 10045 4915 10075
rect 4915 10045 4916 10075
rect 4884 10044 4916 10045
rect 4884 9995 4916 9996
rect 4884 9965 4885 9995
rect 4885 9965 4915 9995
rect 4915 9965 4916 9995
rect 4884 9964 4916 9965
rect 4884 9915 4916 9916
rect 4884 9885 4885 9915
rect 4885 9885 4915 9915
rect 4915 9885 4916 9915
rect 4884 9884 4916 9885
rect 4884 9835 4916 9836
rect 4884 9805 4885 9835
rect 4885 9805 4915 9835
rect 4915 9805 4916 9835
rect 4884 9804 4916 9805
rect 4884 9755 4916 9756
rect 4884 9725 4885 9755
rect 4885 9725 4915 9755
rect 4915 9725 4916 9755
rect 4884 9724 4916 9725
rect 4884 9355 4916 9356
rect 4884 9325 4885 9355
rect 4885 9325 4915 9355
rect 4915 9325 4916 9355
rect 4884 9324 4916 9325
rect 4884 9275 4916 9276
rect 4884 9245 4885 9275
rect 4885 9245 4915 9275
rect 4915 9245 4916 9275
rect 4884 9244 4916 9245
rect 4884 9195 4916 9196
rect 4884 9165 4885 9195
rect 4885 9165 4915 9195
rect 4915 9165 4916 9195
rect 4884 9164 4916 9165
rect 4884 8875 4916 8876
rect 4884 8845 4885 8875
rect 4885 8845 4915 8875
rect 4915 8845 4916 8875
rect 4884 8844 4916 8845
rect 4884 8795 4916 8796
rect 4884 8765 4885 8795
rect 4885 8765 4915 8795
rect 4915 8765 4916 8795
rect 4884 8764 4916 8765
rect 4884 8715 4916 8716
rect 4884 8685 4885 8715
rect 4885 8685 4915 8715
rect 4915 8685 4916 8715
rect 4884 8684 4916 8685
rect 4884 8635 4916 8636
rect 4884 8605 4885 8635
rect 4885 8605 4915 8635
rect 4915 8605 4916 8635
rect 4884 8604 4916 8605
rect 4884 8555 4916 8556
rect 4884 8525 4885 8555
rect 4885 8525 4915 8555
rect 4915 8525 4916 8555
rect 4884 8524 4916 8525
rect 4884 7635 4916 7636
rect 4884 7605 4885 7635
rect 4885 7605 4915 7635
rect 4915 7605 4916 7635
rect 4884 7604 4916 7605
rect 4884 7555 4916 7556
rect 4884 7525 4885 7555
rect 4885 7525 4915 7555
rect 4915 7525 4916 7555
rect 4884 7524 4916 7525
rect 4884 7475 4916 7476
rect 4884 7445 4885 7475
rect 4885 7445 4915 7475
rect 4915 7445 4916 7475
rect 4884 7444 4916 7445
rect 4884 7395 4916 7396
rect 4884 7365 4885 7395
rect 4885 7365 4915 7395
rect 4915 7365 4916 7395
rect 4884 7364 4916 7365
rect 4884 7315 4916 7316
rect 4884 7285 4885 7315
rect 4885 7285 4915 7315
rect 4915 7285 4916 7315
rect 4884 7284 4916 7285
rect 4884 7235 4916 7236
rect 4884 7205 4885 7235
rect 4885 7205 4915 7235
rect 4915 7205 4916 7235
rect 4884 7204 4916 7205
rect 4884 7155 4916 7156
rect 4884 7125 4885 7155
rect 4885 7125 4915 7155
rect 4915 7125 4916 7155
rect 4884 7124 4916 7125
rect 4884 7075 4916 7076
rect 4884 7045 4885 7075
rect 4885 7045 4915 7075
rect 4915 7045 4916 7075
rect 4884 7044 4916 7045
rect 4884 6755 4916 6756
rect 4884 6725 4885 6755
rect 4885 6725 4915 6755
rect 4915 6725 4916 6755
rect 4884 6724 4916 6725
rect 4884 6675 4916 6676
rect 4884 6645 4885 6675
rect 4885 6645 4915 6675
rect 4915 6645 4916 6675
rect 4884 6644 4916 6645
rect 4884 6595 4916 6596
rect 4884 6565 4885 6595
rect 4885 6565 4915 6595
rect 4915 6565 4916 6595
rect 4884 6564 4916 6565
rect 4884 6515 4916 6516
rect 4884 6485 4885 6515
rect 4885 6485 4915 6515
rect 4915 6485 4916 6515
rect 4884 6484 4916 6485
rect 4884 6435 4916 6436
rect 4884 6405 4885 6435
rect 4885 6405 4915 6435
rect 4915 6405 4916 6435
rect 4884 6404 4916 6405
rect 4884 6355 4916 6356
rect 4884 6325 4885 6355
rect 4885 6325 4915 6355
rect 4915 6325 4916 6355
rect 4884 6324 4916 6325
rect 4884 5795 4916 5796
rect 4884 5765 4885 5795
rect 4885 5765 4915 5795
rect 4915 5765 4916 5795
rect 4884 5764 4916 5765
rect 4884 5715 4916 5716
rect 4884 5685 4885 5715
rect 4885 5685 4915 5715
rect 4915 5685 4916 5715
rect 4884 5684 4916 5685
rect 4884 5635 4916 5636
rect 4884 5605 4885 5635
rect 4885 5605 4915 5635
rect 4915 5605 4916 5635
rect 4884 5604 4916 5605
rect 4884 5555 4916 5556
rect 4884 5525 4885 5555
rect 4885 5525 4915 5555
rect 4915 5525 4916 5555
rect 4884 5524 4916 5525
rect 4884 5475 4916 5476
rect 4884 5445 4885 5475
rect 4885 5445 4915 5475
rect 4915 5445 4916 5475
rect 4884 5444 4916 5445
rect 4884 5395 4916 5396
rect 4884 5365 4885 5395
rect 4885 5365 4915 5395
rect 4915 5365 4916 5395
rect 4884 5364 4916 5365
rect 4884 5315 4916 5316
rect 4884 5285 4885 5315
rect 4885 5285 4915 5315
rect 4915 5285 4916 5315
rect 4884 5284 4916 5285
rect 4884 5235 4916 5236
rect 4884 5205 4885 5235
rect 4885 5205 4915 5235
rect 4915 5205 4916 5235
rect 4884 5204 4916 5205
rect 4884 5155 4916 5156
rect 4884 5125 4885 5155
rect 4885 5125 4915 5155
rect 4915 5125 4916 5155
rect 4884 5124 4916 5125
rect 4884 5075 4916 5076
rect 4884 5045 4885 5075
rect 4885 5045 4915 5075
rect 4915 5045 4916 5075
rect 4884 5044 4916 5045
rect 4884 4995 4916 4996
rect 4884 4965 4885 4995
rect 4885 4965 4915 4995
rect 4915 4965 4916 4995
rect 4884 4964 4916 4965
rect 4884 4435 4916 4436
rect 4884 4405 4885 4435
rect 4885 4405 4915 4435
rect 4915 4405 4916 4435
rect 4884 4404 4916 4405
rect 4884 4355 4916 4356
rect 4884 4325 4885 4355
rect 4885 4325 4915 4355
rect 4915 4325 4916 4355
rect 4884 4324 4916 4325
rect 4884 4275 4916 4276
rect 4884 4245 4885 4275
rect 4885 4245 4915 4275
rect 4915 4245 4916 4275
rect 4884 4244 4916 4245
rect 4884 4195 4916 4196
rect 4884 4165 4885 4195
rect 4885 4165 4915 4195
rect 4915 4165 4916 4195
rect 4884 4164 4916 4165
rect 4884 4115 4916 4116
rect 4884 4085 4885 4115
rect 4885 4085 4915 4115
rect 4915 4085 4916 4115
rect 4884 4084 4916 4085
rect 4884 4035 4916 4036
rect 4884 4005 4885 4035
rect 4885 4005 4915 4035
rect 4915 4005 4916 4035
rect 4884 4004 4916 4005
rect 4884 3955 4916 3956
rect 4884 3925 4885 3955
rect 4885 3925 4915 3955
rect 4915 3925 4916 3955
rect 4884 3924 4916 3925
rect 4884 3155 4916 3156
rect 4884 3125 4885 3155
rect 4885 3125 4915 3155
rect 4915 3125 4916 3155
rect 4884 3124 4916 3125
rect 4884 3075 4916 3076
rect 4884 3045 4885 3075
rect 4885 3045 4915 3075
rect 4915 3045 4916 3075
rect 4884 3044 4916 3045
rect 4884 2995 4916 2996
rect 4884 2965 4885 2995
rect 4885 2965 4915 2995
rect 4915 2965 4916 2995
rect 4884 2964 4916 2965
rect 4884 2915 4916 2916
rect 4884 2885 4885 2915
rect 4885 2885 4915 2915
rect 4915 2885 4916 2915
rect 4884 2884 4916 2885
rect 4884 2835 4916 2836
rect 4884 2805 4885 2835
rect 4885 2805 4915 2835
rect 4915 2805 4916 2835
rect 4884 2804 4916 2805
rect 4884 2755 4916 2756
rect 4884 2725 4885 2755
rect 4885 2725 4915 2755
rect 4915 2725 4916 2755
rect 4884 2724 4916 2725
rect 4884 2675 4916 2676
rect 4884 2645 4885 2675
rect 4885 2645 4915 2675
rect 4915 2645 4916 2675
rect 4884 2644 4916 2645
rect 4884 2595 4916 2596
rect 4884 2565 4885 2595
rect 4885 2565 4915 2595
rect 4915 2565 4916 2595
rect 4884 2564 4916 2565
rect 4884 2515 4916 2516
rect 4884 2485 4885 2515
rect 4885 2485 4915 2515
rect 4915 2485 4916 2515
rect 4884 2484 4916 2485
rect 4884 2435 4916 2436
rect 4884 2405 4885 2435
rect 4885 2405 4915 2435
rect 4915 2405 4916 2435
rect 4884 2404 4916 2405
rect 4884 2355 4916 2356
rect 4884 2325 4885 2355
rect 4885 2325 4915 2355
rect 4915 2325 4916 2355
rect 4884 2324 4916 2325
rect 4884 2275 4916 2276
rect 4884 2245 4885 2275
rect 4885 2245 4915 2275
rect 4915 2245 4916 2275
rect 4884 2244 4916 2245
rect 4884 2195 4916 2196
rect 4884 2165 4885 2195
rect 4885 2165 4915 2195
rect 4915 2165 4916 2195
rect 4884 2164 4916 2165
rect 4884 2115 4916 2116
rect 4884 2085 4885 2115
rect 4885 2085 4915 2115
rect 4915 2085 4916 2115
rect 4884 2084 4916 2085
rect 4884 2035 4916 2036
rect 4884 2005 4885 2035
rect 4885 2005 4915 2035
rect 4915 2005 4916 2035
rect 4884 2004 4916 2005
rect 4884 1635 4916 1636
rect 4884 1605 4885 1635
rect 4885 1605 4915 1635
rect 4915 1605 4916 1635
rect 4884 1604 4916 1605
rect 4884 1555 4916 1556
rect 4884 1525 4885 1555
rect 4885 1525 4915 1555
rect 4915 1525 4916 1555
rect 4884 1524 4916 1525
rect 4884 1475 4916 1476
rect 4884 1445 4885 1475
rect 4885 1445 4915 1475
rect 4915 1445 4916 1475
rect 4884 1444 4916 1445
rect 4884 1395 4916 1396
rect 4884 1365 4885 1395
rect 4885 1365 4915 1395
rect 4915 1365 4916 1395
rect 4884 1364 4916 1365
rect 4884 1315 4916 1316
rect 4884 1285 4885 1315
rect 4885 1285 4915 1315
rect 4915 1285 4916 1315
rect 4884 1284 4916 1285
rect 4884 1235 4916 1236
rect 4884 1205 4885 1235
rect 4885 1205 4915 1235
rect 4915 1205 4916 1235
rect 4884 1204 4916 1205
rect 4884 1155 4916 1156
rect 4884 1125 4885 1155
rect 4885 1125 4915 1155
rect 4915 1125 4916 1155
rect 4884 1124 4916 1125
rect 4884 1075 4916 1076
rect 4884 1045 4885 1075
rect 4885 1045 4915 1075
rect 4915 1045 4916 1075
rect 4884 1044 4916 1045
rect 4884 755 4916 756
rect 4884 725 4885 755
rect 4885 725 4915 755
rect 4915 725 4916 755
rect 4884 724 4916 725
rect 4884 675 4916 676
rect 4884 645 4885 675
rect 4885 645 4915 675
rect 4915 645 4916 675
rect 4884 644 4916 645
rect 4884 595 4916 596
rect 4884 565 4885 595
rect 4885 565 4915 595
rect 4915 565 4916 595
rect 4884 564 4916 565
rect 4884 195 4916 196
rect 4884 165 4885 195
rect 4885 165 4915 195
rect 4915 165 4916 195
rect 4884 164 4916 165
rect 4884 115 4916 116
rect 4884 85 4885 115
rect 4885 85 4915 115
rect 4915 85 4916 115
rect 4884 84 4916 85
rect 4884 35 4916 36
rect 4884 5 4885 35
rect 4885 5 4915 35
rect 4915 5 4916 35
rect 4884 4 4916 5
rect 5044 12635 5076 12636
rect 5044 12605 5045 12635
rect 5045 12605 5075 12635
rect 5075 12605 5076 12635
rect 5044 12604 5076 12605
rect 5044 12555 5076 12556
rect 5044 12525 5045 12555
rect 5045 12525 5075 12555
rect 5075 12525 5076 12555
rect 5044 12524 5076 12525
rect 5044 12475 5076 12476
rect 5044 12445 5045 12475
rect 5045 12445 5075 12475
rect 5075 12445 5076 12475
rect 5044 12444 5076 12445
rect 5044 12395 5076 12396
rect 5044 12365 5045 12395
rect 5045 12365 5075 12395
rect 5075 12365 5076 12395
rect 5044 12364 5076 12365
rect 5044 12315 5076 12316
rect 5044 12285 5045 12315
rect 5045 12285 5075 12315
rect 5075 12285 5076 12315
rect 5044 12284 5076 12285
rect 5044 12235 5076 12236
rect 5044 12205 5045 12235
rect 5045 12205 5075 12235
rect 5075 12205 5076 12235
rect 5044 12204 5076 12205
rect 5044 12155 5076 12156
rect 5044 12125 5045 12155
rect 5045 12125 5075 12155
rect 5075 12125 5076 12155
rect 5044 12124 5076 12125
rect 5044 11835 5076 11836
rect 5044 11805 5045 11835
rect 5045 11805 5075 11835
rect 5075 11805 5076 11835
rect 5044 11804 5076 11805
rect 5044 11755 5076 11756
rect 5044 11725 5045 11755
rect 5045 11725 5075 11755
rect 5075 11725 5076 11755
rect 5044 11724 5076 11725
rect 5044 11675 5076 11676
rect 5044 11645 5045 11675
rect 5045 11645 5075 11675
rect 5075 11645 5076 11675
rect 5044 11644 5076 11645
rect 5044 11595 5076 11596
rect 5044 11565 5045 11595
rect 5045 11565 5075 11595
rect 5075 11565 5076 11595
rect 5044 11564 5076 11565
rect 5044 11515 5076 11516
rect 5044 11485 5045 11515
rect 5045 11485 5075 11515
rect 5075 11485 5076 11515
rect 5044 11484 5076 11485
rect 5044 11435 5076 11436
rect 5044 11405 5045 11435
rect 5045 11405 5075 11435
rect 5075 11405 5076 11435
rect 5044 11404 5076 11405
rect 5044 10875 5076 10876
rect 5044 10845 5045 10875
rect 5045 10845 5075 10875
rect 5075 10845 5076 10875
rect 5044 10844 5076 10845
rect 5044 10795 5076 10796
rect 5044 10765 5045 10795
rect 5045 10765 5075 10795
rect 5075 10765 5076 10795
rect 5044 10764 5076 10765
rect 5044 10715 5076 10716
rect 5044 10685 5045 10715
rect 5045 10685 5075 10715
rect 5075 10685 5076 10715
rect 5044 10684 5076 10685
rect 5044 10635 5076 10636
rect 5044 10605 5045 10635
rect 5045 10605 5075 10635
rect 5075 10605 5076 10635
rect 5044 10604 5076 10605
rect 5044 10555 5076 10556
rect 5044 10525 5045 10555
rect 5045 10525 5075 10555
rect 5075 10525 5076 10555
rect 5044 10524 5076 10525
rect 5044 10475 5076 10476
rect 5044 10445 5045 10475
rect 5045 10445 5075 10475
rect 5075 10445 5076 10475
rect 5044 10444 5076 10445
rect 5044 10395 5076 10396
rect 5044 10365 5045 10395
rect 5045 10365 5075 10395
rect 5075 10365 5076 10395
rect 5044 10364 5076 10365
rect 5044 10315 5076 10316
rect 5044 10285 5045 10315
rect 5045 10285 5075 10315
rect 5075 10285 5076 10315
rect 5044 10284 5076 10285
rect 5044 10235 5076 10236
rect 5044 10205 5045 10235
rect 5045 10205 5075 10235
rect 5075 10205 5076 10235
rect 5044 10204 5076 10205
rect 5044 10155 5076 10156
rect 5044 10125 5045 10155
rect 5045 10125 5075 10155
rect 5075 10125 5076 10155
rect 5044 10124 5076 10125
rect 5044 10075 5076 10076
rect 5044 10045 5045 10075
rect 5045 10045 5075 10075
rect 5075 10045 5076 10075
rect 5044 10044 5076 10045
rect 5044 9995 5076 9996
rect 5044 9965 5045 9995
rect 5045 9965 5075 9995
rect 5075 9965 5076 9995
rect 5044 9964 5076 9965
rect 5044 9915 5076 9916
rect 5044 9885 5045 9915
rect 5045 9885 5075 9915
rect 5075 9885 5076 9915
rect 5044 9884 5076 9885
rect 5044 9835 5076 9836
rect 5044 9805 5045 9835
rect 5045 9805 5075 9835
rect 5075 9805 5076 9835
rect 5044 9804 5076 9805
rect 5044 9755 5076 9756
rect 5044 9725 5045 9755
rect 5045 9725 5075 9755
rect 5075 9725 5076 9755
rect 5044 9724 5076 9725
rect 5044 9355 5076 9356
rect 5044 9325 5045 9355
rect 5045 9325 5075 9355
rect 5075 9325 5076 9355
rect 5044 9324 5076 9325
rect 5044 9275 5076 9276
rect 5044 9245 5045 9275
rect 5045 9245 5075 9275
rect 5075 9245 5076 9275
rect 5044 9244 5076 9245
rect 5044 9195 5076 9196
rect 5044 9165 5045 9195
rect 5045 9165 5075 9195
rect 5075 9165 5076 9195
rect 5044 9164 5076 9165
rect 5044 8875 5076 8876
rect 5044 8845 5045 8875
rect 5045 8845 5075 8875
rect 5075 8845 5076 8875
rect 5044 8844 5076 8845
rect 5044 8795 5076 8796
rect 5044 8765 5045 8795
rect 5045 8765 5075 8795
rect 5075 8765 5076 8795
rect 5044 8764 5076 8765
rect 5044 8715 5076 8716
rect 5044 8685 5045 8715
rect 5045 8685 5075 8715
rect 5075 8685 5076 8715
rect 5044 8684 5076 8685
rect 5044 8635 5076 8636
rect 5044 8605 5045 8635
rect 5045 8605 5075 8635
rect 5075 8605 5076 8635
rect 5044 8604 5076 8605
rect 5044 8555 5076 8556
rect 5044 8525 5045 8555
rect 5045 8525 5075 8555
rect 5075 8525 5076 8555
rect 5044 8524 5076 8525
rect 5044 7635 5076 7636
rect 5044 7605 5045 7635
rect 5045 7605 5075 7635
rect 5075 7605 5076 7635
rect 5044 7604 5076 7605
rect 5044 7555 5076 7556
rect 5044 7525 5045 7555
rect 5045 7525 5075 7555
rect 5075 7525 5076 7555
rect 5044 7524 5076 7525
rect 5044 7475 5076 7476
rect 5044 7445 5045 7475
rect 5045 7445 5075 7475
rect 5075 7445 5076 7475
rect 5044 7444 5076 7445
rect 5044 7395 5076 7396
rect 5044 7365 5045 7395
rect 5045 7365 5075 7395
rect 5075 7365 5076 7395
rect 5044 7364 5076 7365
rect 5044 7315 5076 7316
rect 5044 7285 5045 7315
rect 5045 7285 5075 7315
rect 5075 7285 5076 7315
rect 5044 7284 5076 7285
rect 5044 7235 5076 7236
rect 5044 7205 5045 7235
rect 5045 7205 5075 7235
rect 5075 7205 5076 7235
rect 5044 7204 5076 7205
rect 5044 7155 5076 7156
rect 5044 7125 5045 7155
rect 5045 7125 5075 7155
rect 5075 7125 5076 7155
rect 5044 7124 5076 7125
rect 5044 7075 5076 7076
rect 5044 7045 5045 7075
rect 5045 7045 5075 7075
rect 5075 7045 5076 7075
rect 5044 7044 5076 7045
rect 5044 6755 5076 6756
rect 5044 6725 5045 6755
rect 5045 6725 5075 6755
rect 5075 6725 5076 6755
rect 5044 6724 5076 6725
rect 5044 6675 5076 6676
rect 5044 6645 5045 6675
rect 5045 6645 5075 6675
rect 5075 6645 5076 6675
rect 5044 6644 5076 6645
rect 5044 6595 5076 6596
rect 5044 6565 5045 6595
rect 5045 6565 5075 6595
rect 5075 6565 5076 6595
rect 5044 6564 5076 6565
rect 5044 6515 5076 6516
rect 5044 6485 5045 6515
rect 5045 6485 5075 6515
rect 5075 6485 5076 6515
rect 5044 6484 5076 6485
rect 5044 6435 5076 6436
rect 5044 6405 5045 6435
rect 5045 6405 5075 6435
rect 5075 6405 5076 6435
rect 5044 6404 5076 6405
rect 5044 6355 5076 6356
rect 5044 6325 5045 6355
rect 5045 6325 5075 6355
rect 5075 6325 5076 6355
rect 5044 6324 5076 6325
rect 5044 5795 5076 5796
rect 5044 5765 5045 5795
rect 5045 5765 5075 5795
rect 5075 5765 5076 5795
rect 5044 5764 5076 5765
rect 5044 5715 5076 5716
rect 5044 5685 5045 5715
rect 5045 5685 5075 5715
rect 5075 5685 5076 5715
rect 5044 5684 5076 5685
rect 5044 5635 5076 5636
rect 5044 5605 5045 5635
rect 5045 5605 5075 5635
rect 5075 5605 5076 5635
rect 5044 5604 5076 5605
rect 5044 5555 5076 5556
rect 5044 5525 5045 5555
rect 5045 5525 5075 5555
rect 5075 5525 5076 5555
rect 5044 5524 5076 5525
rect 5044 5475 5076 5476
rect 5044 5445 5045 5475
rect 5045 5445 5075 5475
rect 5075 5445 5076 5475
rect 5044 5444 5076 5445
rect 5044 5395 5076 5396
rect 5044 5365 5045 5395
rect 5045 5365 5075 5395
rect 5075 5365 5076 5395
rect 5044 5364 5076 5365
rect 5044 5315 5076 5316
rect 5044 5285 5045 5315
rect 5045 5285 5075 5315
rect 5075 5285 5076 5315
rect 5044 5284 5076 5285
rect 5044 5235 5076 5236
rect 5044 5205 5045 5235
rect 5045 5205 5075 5235
rect 5075 5205 5076 5235
rect 5044 5204 5076 5205
rect 5044 5155 5076 5156
rect 5044 5125 5045 5155
rect 5045 5125 5075 5155
rect 5075 5125 5076 5155
rect 5044 5124 5076 5125
rect 5044 5075 5076 5076
rect 5044 5045 5045 5075
rect 5045 5045 5075 5075
rect 5075 5045 5076 5075
rect 5044 5044 5076 5045
rect 5044 4995 5076 4996
rect 5044 4965 5045 4995
rect 5045 4965 5075 4995
rect 5075 4965 5076 4995
rect 5044 4964 5076 4965
rect 5044 4435 5076 4436
rect 5044 4405 5045 4435
rect 5045 4405 5075 4435
rect 5075 4405 5076 4435
rect 5044 4404 5076 4405
rect 5044 4355 5076 4356
rect 5044 4325 5045 4355
rect 5045 4325 5075 4355
rect 5075 4325 5076 4355
rect 5044 4324 5076 4325
rect 5044 4275 5076 4276
rect 5044 4245 5045 4275
rect 5045 4245 5075 4275
rect 5075 4245 5076 4275
rect 5044 4244 5076 4245
rect 5044 4195 5076 4196
rect 5044 4165 5045 4195
rect 5045 4165 5075 4195
rect 5075 4165 5076 4195
rect 5044 4164 5076 4165
rect 5044 4115 5076 4116
rect 5044 4085 5045 4115
rect 5045 4085 5075 4115
rect 5075 4085 5076 4115
rect 5044 4084 5076 4085
rect 5044 4035 5076 4036
rect 5044 4005 5045 4035
rect 5045 4005 5075 4035
rect 5075 4005 5076 4035
rect 5044 4004 5076 4005
rect 5044 3955 5076 3956
rect 5044 3925 5045 3955
rect 5045 3925 5075 3955
rect 5075 3925 5076 3955
rect 5044 3924 5076 3925
rect 5044 3155 5076 3156
rect 5044 3125 5045 3155
rect 5045 3125 5075 3155
rect 5075 3125 5076 3155
rect 5044 3124 5076 3125
rect 5044 3075 5076 3076
rect 5044 3045 5045 3075
rect 5045 3045 5075 3075
rect 5075 3045 5076 3075
rect 5044 3044 5076 3045
rect 5044 2995 5076 2996
rect 5044 2965 5045 2995
rect 5045 2965 5075 2995
rect 5075 2965 5076 2995
rect 5044 2964 5076 2965
rect 5044 2915 5076 2916
rect 5044 2885 5045 2915
rect 5045 2885 5075 2915
rect 5075 2885 5076 2915
rect 5044 2884 5076 2885
rect 5044 2835 5076 2836
rect 5044 2805 5045 2835
rect 5045 2805 5075 2835
rect 5075 2805 5076 2835
rect 5044 2804 5076 2805
rect 5044 2755 5076 2756
rect 5044 2725 5045 2755
rect 5045 2725 5075 2755
rect 5075 2725 5076 2755
rect 5044 2724 5076 2725
rect 5044 2675 5076 2676
rect 5044 2645 5045 2675
rect 5045 2645 5075 2675
rect 5075 2645 5076 2675
rect 5044 2644 5076 2645
rect 5044 2595 5076 2596
rect 5044 2565 5045 2595
rect 5045 2565 5075 2595
rect 5075 2565 5076 2595
rect 5044 2564 5076 2565
rect 5044 2515 5076 2516
rect 5044 2485 5045 2515
rect 5045 2485 5075 2515
rect 5075 2485 5076 2515
rect 5044 2484 5076 2485
rect 5044 2435 5076 2436
rect 5044 2405 5045 2435
rect 5045 2405 5075 2435
rect 5075 2405 5076 2435
rect 5044 2404 5076 2405
rect 5044 2355 5076 2356
rect 5044 2325 5045 2355
rect 5045 2325 5075 2355
rect 5075 2325 5076 2355
rect 5044 2324 5076 2325
rect 5044 2275 5076 2276
rect 5044 2245 5045 2275
rect 5045 2245 5075 2275
rect 5075 2245 5076 2275
rect 5044 2244 5076 2245
rect 5044 2195 5076 2196
rect 5044 2165 5045 2195
rect 5045 2165 5075 2195
rect 5075 2165 5076 2195
rect 5044 2164 5076 2165
rect 5044 2115 5076 2116
rect 5044 2085 5045 2115
rect 5045 2085 5075 2115
rect 5075 2085 5076 2115
rect 5044 2084 5076 2085
rect 5044 2035 5076 2036
rect 5044 2005 5045 2035
rect 5045 2005 5075 2035
rect 5075 2005 5076 2035
rect 5044 2004 5076 2005
rect 5044 1635 5076 1636
rect 5044 1605 5045 1635
rect 5045 1605 5075 1635
rect 5075 1605 5076 1635
rect 5044 1604 5076 1605
rect 5044 1555 5076 1556
rect 5044 1525 5045 1555
rect 5045 1525 5075 1555
rect 5075 1525 5076 1555
rect 5044 1524 5076 1525
rect 5044 1475 5076 1476
rect 5044 1445 5045 1475
rect 5045 1445 5075 1475
rect 5075 1445 5076 1475
rect 5044 1444 5076 1445
rect 5044 1395 5076 1396
rect 5044 1365 5045 1395
rect 5045 1365 5075 1395
rect 5075 1365 5076 1395
rect 5044 1364 5076 1365
rect 5044 1315 5076 1316
rect 5044 1285 5045 1315
rect 5045 1285 5075 1315
rect 5075 1285 5076 1315
rect 5044 1284 5076 1285
rect 5044 1235 5076 1236
rect 5044 1205 5045 1235
rect 5045 1205 5075 1235
rect 5075 1205 5076 1235
rect 5044 1204 5076 1205
rect 5044 1155 5076 1156
rect 5044 1125 5045 1155
rect 5045 1125 5075 1155
rect 5075 1125 5076 1155
rect 5044 1124 5076 1125
rect 5044 1075 5076 1076
rect 5044 1045 5045 1075
rect 5045 1045 5075 1075
rect 5075 1045 5076 1075
rect 5044 1044 5076 1045
rect 5044 755 5076 756
rect 5044 725 5045 755
rect 5045 725 5075 755
rect 5075 725 5076 755
rect 5044 724 5076 725
rect 5044 675 5076 676
rect 5044 645 5045 675
rect 5045 645 5075 675
rect 5075 645 5076 675
rect 5044 644 5076 645
rect 5044 595 5076 596
rect 5044 565 5045 595
rect 5045 565 5075 595
rect 5075 565 5076 595
rect 5044 564 5076 565
rect 5044 195 5076 196
rect 5044 165 5045 195
rect 5045 165 5075 195
rect 5075 165 5076 195
rect 5044 164 5076 165
rect 5044 115 5076 116
rect 5044 85 5045 115
rect 5045 85 5075 115
rect 5075 85 5076 115
rect 5044 84 5076 85
rect 5044 35 5076 36
rect 5044 5 5045 35
rect 5045 5 5075 35
rect 5075 5 5076 35
rect 5044 4 5076 5
rect 5124 15364 5156 15396
rect 5124 14084 5156 14116
rect 5124 12635 5156 12636
rect 5124 12605 5125 12635
rect 5125 12605 5155 12635
rect 5155 12605 5156 12635
rect 5124 12604 5156 12605
rect 5124 12555 5156 12556
rect 5124 12525 5125 12555
rect 5125 12525 5155 12555
rect 5155 12525 5156 12555
rect 5124 12524 5156 12525
rect 5124 12475 5156 12476
rect 5124 12445 5125 12475
rect 5125 12445 5155 12475
rect 5155 12445 5156 12475
rect 5124 12444 5156 12445
rect 5124 12395 5156 12396
rect 5124 12365 5125 12395
rect 5125 12365 5155 12395
rect 5155 12365 5156 12395
rect 5124 12364 5156 12365
rect 5124 12315 5156 12316
rect 5124 12285 5125 12315
rect 5125 12285 5155 12315
rect 5155 12285 5156 12315
rect 5124 12284 5156 12285
rect 5124 12235 5156 12236
rect 5124 12205 5125 12235
rect 5125 12205 5155 12235
rect 5155 12205 5156 12235
rect 5124 12204 5156 12205
rect 5124 12155 5156 12156
rect 5124 12125 5125 12155
rect 5125 12125 5155 12155
rect 5155 12125 5156 12155
rect 5124 12124 5156 12125
rect 5124 11835 5156 11836
rect 5124 11805 5125 11835
rect 5125 11805 5155 11835
rect 5155 11805 5156 11835
rect 5124 11804 5156 11805
rect 5124 11755 5156 11756
rect 5124 11725 5125 11755
rect 5125 11725 5155 11755
rect 5155 11725 5156 11755
rect 5124 11724 5156 11725
rect 5124 11675 5156 11676
rect 5124 11645 5125 11675
rect 5125 11645 5155 11675
rect 5155 11645 5156 11675
rect 5124 11644 5156 11645
rect 5124 11595 5156 11596
rect 5124 11565 5125 11595
rect 5125 11565 5155 11595
rect 5155 11565 5156 11595
rect 5124 11564 5156 11565
rect 5124 11515 5156 11516
rect 5124 11485 5125 11515
rect 5125 11485 5155 11515
rect 5155 11485 5156 11515
rect 5124 11484 5156 11485
rect 5124 11435 5156 11436
rect 5124 11405 5125 11435
rect 5125 11405 5155 11435
rect 5155 11405 5156 11435
rect 5124 11404 5156 11405
rect 5124 10875 5156 10876
rect 5124 10845 5125 10875
rect 5125 10845 5155 10875
rect 5155 10845 5156 10875
rect 5124 10844 5156 10845
rect 5124 10795 5156 10796
rect 5124 10765 5125 10795
rect 5125 10765 5155 10795
rect 5155 10765 5156 10795
rect 5124 10764 5156 10765
rect 5124 10715 5156 10716
rect 5124 10685 5125 10715
rect 5125 10685 5155 10715
rect 5155 10685 5156 10715
rect 5124 10684 5156 10685
rect 5124 10635 5156 10636
rect 5124 10605 5125 10635
rect 5125 10605 5155 10635
rect 5155 10605 5156 10635
rect 5124 10604 5156 10605
rect 5124 10555 5156 10556
rect 5124 10525 5125 10555
rect 5125 10525 5155 10555
rect 5155 10525 5156 10555
rect 5124 10524 5156 10525
rect 5124 10475 5156 10476
rect 5124 10445 5125 10475
rect 5125 10445 5155 10475
rect 5155 10445 5156 10475
rect 5124 10444 5156 10445
rect 5124 10395 5156 10396
rect 5124 10365 5125 10395
rect 5125 10365 5155 10395
rect 5155 10365 5156 10395
rect 5124 10364 5156 10365
rect 5124 10315 5156 10316
rect 5124 10285 5125 10315
rect 5125 10285 5155 10315
rect 5155 10285 5156 10315
rect 5124 10284 5156 10285
rect 5124 10235 5156 10236
rect 5124 10205 5125 10235
rect 5125 10205 5155 10235
rect 5155 10205 5156 10235
rect 5124 10204 5156 10205
rect 5124 10155 5156 10156
rect 5124 10125 5125 10155
rect 5125 10125 5155 10155
rect 5155 10125 5156 10155
rect 5124 10124 5156 10125
rect 5124 10075 5156 10076
rect 5124 10045 5125 10075
rect 5125 10045 5155 10075
rect 5155 10045 5156 10075
rect 5124 10044 5156 10045
rect 5124 9995 5156 9996
rect 5124 9965 5125 9995
rect 5125 9965 5155 9995
rect 5155 9965 5156 9995
rect 5124 9964 5156 9965
rect 5124 9915 5156 9916
rect 5124 9885 5125 9915
rect 5125 9885 5155 9915
rect 5155 9885 5156 9915
rect 5124 9884 5156 9885
rect 5124 9835 5156 9836
rect 5124 9805 5125 9835
rect 5125 9805 5155 9835
rect 5155 9805 5156 9835
rect 5124 9804 5156 9805
rect 5124 9755 5156 9756
rect 5124 9725 5125 9755
rect 5125 9725 5155 9755
rect 5155 9725 5156 9755
rect 5124 9724 5156 9725
rect 5124 9355 5156 9356
rect 5124 9325 5125 9355
rect 5125 9325 5155 9355
rect 5155 9325 5156 9355
rect 5124 9324 5156 9325
rect 5124 9275 5156 9276
rect 5124 9245 5125 9275
rect 5125 9245 5155 9275
rect 5155 9245 5156 9275
rect 5124 9244 5156 9245
rect 5124 9195 5156 9196
rect 5124 9165 5125 9195
rect 5125 9165 5155 9195
rect 5155 9165 5156 9195
rect 5124 9164 5156 9165
rect 5124 8875 5156 8876
rect 5124 8845 5125 8875
rect 5125 8845 5155 8875
rect 5155 8845 5156 8875
rect 5124 8844 5156 8845
rect 5124 8795 5156 8796
rect 5124 8765 5125 8795
rect 5125 8765 5155 8795
rect 5155 8765 5156 8795
rect 5124 8764 5156 8765
rect 5124 8715 5156 8716
rect 5124 8685 5125 8715
rect 5125 8685 5155 8715
rect 5155 8685 5156 8715
rect 5124 8684 5156 8685
rect 5124 8635 5156 8636
rect 5124 8605 5125 8635
rect 5125 8605 5155 8635
rect 5155 8605 5156 8635
rect 5124 8604 5156 8605
rect 5124 8555 5156 8556
rect 5124 8525 5125 8555
rect 5125 8525 5155 8555
rect 5155 8525 5156 8555
rect 5124 8524 5156 8525
rect 5124 7635 5156 7636
rect 5124 7605 5125 7635
rect 5125 7605 5155 7635
rect 5155 7605 5156 7635
rect 5124 7604 5156 7605
rect 5124 7555 5156 7556
rect 5124 7525 5125 7555
rect 5125 7525 5155 7555
rect 5155 7525 5156 7555
rect 5124 7524 5156 7525
rect 5124 7475 5156 7476
rect 5124 7445 5125 7475
rect 5125 7445 5155 7475
rect 5155 7445 5156 7475
rect 5124 7444 5156 7445
rect 5124 7395 5156 7396
rect 5124 7365 5125 7395
rect 5125 7365 5155 7395
rect 5155 7365 5156 7395
rect 5124 7364 5156 7365
rect 5124 7315 5156 7316
rect 5124 7285 5125 7315
rect 5125 7285 5155 7315
rect 5155 7285 5156 7315
rect 5124 7284 5156 7285
rect 5124 7235 5156 7236
rect 5124 7205 5125 7235
rect 5125 7205 5155 7235
rect 5155 7205 5156 7235
rect 5124 7204 5156 7205
rect 5124 7155 5156 7156
rect 5124 7125 5125 7155
rect 5125 7125 5155 7155
rect 5155 7125 5156 7155
rect 5124 7124 5156 7125
rect 5124 7075 5156 7076
rect 5124 7045 5125 7075
rect 5125 7045 5155 7075
rect 5155 7045 5156 7075
rect 5124 7044 5156 7045
rect 5124 6755 5156 6756
rect 5124 6725 5125 6755
rect 5125 6725 5155 6755
rect 5155 6725 5156 6755
rect 5124 6724 5156 6725
rect 5124 6675 5156 6676
rect 5124 6645 5125 6675
rect 5125 6645 5155 6675
rect 5155 6645 5156 6675
rect 5124 6644 5156 6645
rect 5124 6595 5156 6596
rect 5124 6565 5125 6595
rect 5125 6565 5155 6595
rect 5155 6565 5156 6595
rect 5124 6564 5156 6565
rect 5124 6515 5156 6516
rect 5124 6485 5125 6515
rect 5125 6485 5155 6515
rect 5155 6485 5156 6515
rect 5124 6484 5156 6485
rect 5124 6435 5156 6436
rect 5124 6405 5125 6435
rect 5125 6405 5155 6435
rect 5155 6405 5156 6435
rect 5124 6404 5156 6405
rect 5124 6355 5156 6356
rect 5124 6325 5125 6355
rect 5125 6325 5155 6355
rect 5155 6325 5156 6355
rect 5124 6324 5156 6325
rect 5124 5795 5156 5796
rect 5124 5765 5125 5795
rect 5125 5765 5155 5795
rect 5155 5765 5156 5795
rect 5124 5764 5156 5765
rect 5124 5715 5156 5716
rect 5124 5685 5125 5715
rect 5125 5685 5155 5715
rect 5155 5685 5156 5715
rect 5124 5684 5156 5685
rect 5124 5635 5156 5636
rect 5124 5605 5125 5635
rect 5125 5605 5155 5635
rect 5155 5605 5156 5635
rect 5124 5604 5156 5605
rect 5124 5555 5156 5556
rect 5124 5525 5125 5555
rect 5125 5525 5155 5555
rect 5155 5525 5156 5555
rect 5124 5524 5156 5525
rect 5124 5475 5156 5476
rect 5124 5445 5125 5475
rect 5125 5445 5155 5475
rect 5155 5445 5156 5475
rect 5124 5444 5156 5445
rect 5124 5395 5156 5396
rect 5124 5365 5125 5395
rect 5125 5365 5155 5395
rect 5155 5365 5156 5395
rect 5124 5364 5156 5365
rect 5124 5315 5156 5316
rect 5124 5285 5125 5315
rect 5125 5285 5155 5315
rect 5155 5285 5156 5315
rect 5124 5284 5156 5285
rect 5124 5235 5156 5236
rect 5124 5205 5125 5235
rect 5125 5205 5155 5235
rect 5155 5205 5156 5235
rect 5124 5204 5156 5205
rect 5124 5155 5156 5156
rect 5124 5125 5125 5155
rect 5125 5125 5155 5155
rect 5155 5125 5156 5155
rect 5124 5124 5156 5125
rect 5124 5075 5156 5076
rect 5124 5045 5125 5075
rect 5125 5045 5155 5075
rect 5155 5045 5156 5075
rect 5124 5044 5156 5045
rect 5124 4995 5156 4996
rect 5124 4965 5125 4995
rect 5125 4965 5155 4995
rect 5155 4965 5156 4995
rect 5124 4964 5156 4965
rect 5124 4435 5156 4436
rect 5124 4405 5125 4435
rect 5125 4405 5155 4435
rect 5155 4405 5156 4435
rect 5124 4404 5156 4405
rect 5124 4355 5156 4356
rect 5124 4325 5125 4355
rect 5125 4325 5155 4355
rect 5155 4325 5156 4355
rect 5124 4324 5156 4325
rect 5124 4275 5156 4276
rect 5124 4245 5125 4275
rect 5125 4245 5155 4275
rect 5155 4245 5156 4275
rect 5124 4244 5156 4245
rect 5124 4195 5156 4196
rect 5124 4165 5125 4195
rect 5125 4165 5155 4195
rect 5155 4165 5156 4195
rect 5124 4164 5156 4165
rect 5124 4115 5156 4116
rect 5124 4085 5125 4115
rect 5125 4085 5155 4115
rect 5155 4085 5156 4115
rect 5124 4084 5156 4085
rect 5124 4035 5156 4036
rect 5124 4005 5125 4035
rect 5125 4005 5155 4035
rect 5155 4005 5156 4035
rect 5124 4004 5156 4005
rect 5124 3955 5156 3956
rect 5124 3925 5125 3955
rect 5125 3925 5155 3955
rect 5155 3925 5156 3955
rect 5124 3924 5156 3925
rect 5124 3155 5156 3156
rect 5124 3125 5125 3155
rect 5125 3125 5155 3155
rect 5155 3125 5156 3155
rect 5124 3124 5156 3125
rect 5124 3075 5156 3076
rect 5124 3045 5125 3075
rect 5125 3045 5155 3075
rect 5155 3045 5156 3075
rect 5124 3044 5156 3045
rect 5124 2995 5156 2996
rect 5124 2965 5125 2995
rect 5125 2965 5155 2995
rect 5155 2965 5156 2995
rect 5124 2964 5156 2965
rect 5124 2915 5156 2916
rect 5124 2885 5125 2915
rect 5125 2885 5155 2915
rect 5155 2885 5156 2915
rect 5124 2884 5156 2885
rect 5124 2835 5156 2836
rect 5124 2805 5125 2835
rect 5125 2805 5155 2835
rect 5155 2805 5156 2835
rect 5124 2804 5156 2805
rect 5124 2755 5156 2756
rect 5124 2725 5125 2755
rect 5125 2725 5155 2755
rect 5155 2725 5156 2755
rect 5124 2724 5156 2725
rect 5124 2675 5156 2676
rect 5124 2645 5125 2675
rect 5125 2645 5155 2675
rect 5155 2645 5156 2675
rect 5124 2644 5156 2645
rect 5124 2595 5156 2596
rect 5124 2565 5125 2595
rect 5125 2565 5155 2595
rect 5155 2565 5156 2595
rect 5124 2564 5156 2565
rect 5124 2515 5156 2516
rect 5124 2485 5125 2515
rect 5125 2485 5155 2515
rect 5155 2485 5156 2515
rect 5124 2484 5156 2485
rect 5124 2435 5156 2436
rect 5124 2405 5125 2435
rect 5125 2405 5155 2435
rect 5155 2405 5156 2435
rect 5124 2404 5156 2405
rect 5124 2355 5156 2356
rect 5124 2325 5125 2355
rect 5125 2325 5155 2355
rect 5155 2325 5156 2355
rect 5124 2324 5156 2325
rect 5124 2275 5156 2276
rect 5124 2245 5125 2275
rect 5125 2245 5155 2275
rect 5155 2245 5156 2275
rect 5124 2244 5156 2245
rect 5124 2195 5156 2196
rect 5124 2165 5125 2195
rect 5125 2165 5155 2195
rect 5155 2165 5156 2195
rect 5124 2164 5156 2165
rect 5124 2115 5156 2116
rect 5124 2085 5125 2115
rect 5125 2085 5155 2115
rect 5155 2085 5156 2115
rect 5124 2084 5156 2085
rect 5124 2035 5156 2036
rect 5124 2005 5125 2035
rect 5125 2005 5155 2035
rect 5155 2005 5156 2035
rect 5124 2004 5156 2005
rect 5124 1635 5156 1636
rect 5124 1605 5125 1635
rect 5125 1605 5155 1635
rect 5155 1605 5156 1635
rect 5124 1604 5156 1605
rect 5124 1555 5156 1556
rect 5124 1525 5125 1555
rect 5125 1525 5155 1555
rect 5155 1525 5156 1555
rect 5124 1524 5156 1525
rect 5124 1475 5156 1476
rect 5124 1445 5125 1475
rect 5125 1445 5155 1475
rect 5155 1445 5156 1475
rect 5124 1444 5156 1445
rect 5124 1395 5156 1396
rect 5124 1365 5125 1395
rect 5125 1365 5155 1395
rect 5155 1365 5156 1395
rect 5124 1364 5156 1365
rect 5124 1315 5156 1316
rect 5124 1285 5125 1315
rect 5125 1285 5155 1315
rect 5155 1285 5156 1315
rect 5124 1284 5156 1285
rect 5124 1235 5156 1236
rect 5124 1205 5125 1235
rect 5125 1205 5155 1235
rect 5155 1205 5156 1235
rect 5124 1204 5156 1205
rect 5124 1155 5156 1156
rect 5124 1125 5125 1155
rect 5125 1125 5155 1155
rect 5155 1125 5156 1155
rect 5124 1124 5156 1125
rect 5124 1075 5156 1076
rect 5124 1045 5125 1075
rect 5125 1045 5155 1075
rect 5155 1045 5156 1075
rect 5124 1044 5156 1045
rect 5124 755 5156 756
rect 5124 725 5125 755
rect 5125 725 5155 755
rect 5155 725 5156 755
rect 5124 724 5156 725
rect 5124 675 5156 676
rect 5124 645 5125 675
rect 5125 645 5155 675
rect 5155 645 5156 675
rect 5124 644 5156 645
rect 5124 595 5156 596
rect 5124 565 5125 595
rect 5125 565 5155 595
rect 5155 565 5156 595
rect 5124 564 5156 565
rect 5124 195 5156 196
rect 5124 165 5125 195
rect 5125 165 5155 195
rect 5155 165 5156 195
rect 5124 164 5156 165
rect 5124 115 5156 116
rect 5124 85 5125 115
rect 5125 85 5155 115
rect 5155 85 5156 115
rect 5124 84 5156 85
rect 5124 35 5156 36
rect 5124 5 5125 35
rect 5125 5 5155 35
rect 5155 5 5156 35
rect 5124 4 5156 5
rect 5204 15284 5236 15316
rect 5284 15364 5316 15396
rect 5284 14084 5316 14116
rect 5284 12635 5316 12636
rect 5284 12605 5285 12635
rect 5285 12605 5315 12635
rect 5315 12605 5316 12635
rect 5284 12604 5316 12605
rect 5284 12555 5316 12556
rect 5284 12525 5285 12555
rect 5285 12525 5315 12555
rect 5315 12525 5316 12555
rect 5284 12524 5316 12525
rect 5284 12475 5316 12476
rect 5284 12445 5285 12475
rect 5285 12445 5315 12475
rect 5315 12445 5316 12475
rect 5284 12444 5316 12445
rect 5284 12395 5316 12396
rect 5284 12365 5285 12395
rect 5285 12365 5315 12395
rect 5315 12365 5316 12395
rect 5284 12364 5316 12365
rect 5284 12315 5316 12316
rect 5284 12285 5285 12315
rect 5285 12285 5315 12315
rect 5315 12285 5316 12315
rect 5284 12284 5316 12285
rect 5284 12235 5316 12236
rect 5284 12205 5285 12235
rect 5285 12205 5315 12235
rect 5315 12205 5316 12235
rect 5284 12204 5316 12205
rect 5284 12155 5316 12156
rect 5284 12125 5285 12155
rect 5285 12125 5315 12155
rect 5315 12125 5316 12155
rect 5284 12124 5316 12125
rect 5284 11835 5316 11836
rect 5284 11805 5285 11835
rect 5285 11805 5315 11835
rect 5315 11805 5316 11835
rect 5284 11804 5316 11805
rect 5284 11755 5316 11756
rect 5284 11725 5285 11755
rect 5285 11725 5315 11755
rect 5315 11725 5316 11755
rect 5284 11724 5316 11725
rect 5284 11675 5316 11676
rect 5284 11645 5285 11675
rect 5285 11645 5315 11675
rect 5315 11645 5316 11675
rect 5284 11644 5316 11645
rect 5284 11595 5316 11596
rect 5284 11565 5285 11595
rect 5285 11565 5315 11595
rect 5315 11565 5316 11595
rect 5284 11564 5316 11565
rect 5284 11515 5316 11516
rect 5284 11485 5285 11515
rect 5285 11485 5315 11515
rect 5315 11485 5316 11515
rect 5284 11484 5316 11485
rect 5284 11435 5316 11436
rect 5284 11405 5285 11435
rect 5285 11405 5315 11435
rect 5315 11405 5316 11435
rect 5284 11404 5316 11405
rect 5284 10875 5316 10876
rect 5284 10845 5285 10875
rect 5285 10845 5315 10875
rect 5315 10845 5316 10875
rect 5284 10844 5316 10845
rect 5284 10795 5316 10796
rect 5284 10765 5285 10795
rect 5285 10765 5315 10795
rect 5315 10765 5316 10795
rect 5284 10764 5316 10765
rect 5284 10715 5316 10716
rect 5284 10685 5285 10715
rect 5285 10685 5315 10715
rect 5315 10685 5316 10715
rect 5284 10684 5316 10685
rect 5284 10635 5316 10636
rect 5284 10605 5285 10635
rect 5285 10605 5315 10635
rect 5315 10605 5316 10635
rect 5284 10604 5316 10605
rect 5284 10555 5316 10556
rect 5284 10525 5285 10555
rect 5285 10525 5315 10555
rect 5315 10525 5316 10555
rect 5284 10524 5316 10525
rect 5284 10475 5316 10476
rect 5284 10445 5285 10475
rect 5285 10445 5315 10475
rect 5315 10445 5316 10475
rect 5284 10444 5316 10445
rect 5284 10395 5316 10396
rect 5284 10365 5285 10395
rect 5285 10365 5315 10395
rect 5315 10365 5316 10395
rect 5284 10364 5316 10365
rect 5284 10315 5316 10316
rect 5284 10285 5285 10315
rect 5285 10285 5315 10315
rect 5315 10285 5316 10315
rect 5284 10284 5316 10285
rect 5284 10235 5316 10236
rect 5284 10205 5285 10235
rect 5285 10205 5315 10235
rect 5315 10205 5316 10235
rect 5284 10204 5316 10205
rect 5284 10155 5316 10156
rect 5284 10125 5285 10155
rect 5285 10125 5315 10155
rect 5315 10125 5316 10155
rect 5284 10124 5316 10125
rect 5284 10075 5316 10076
rect 5284 10045 5285 10075
rect 5285 10045 5315 10075
rect 5315 10045 5316 10075
rect 5284 10044 5316 10045
rect 5284 9995 5316 9996
rect 5284 9965 5285 9995
rect 5285 9965 5315 9995
rect 5315 9965 5316 9995
rect 5284 9964 5316 9965
rect 5284 9915 5316 9916
rect 5284 9885 5285 9915
rect 5285 9885 5315 9915
rect 5315 9885 5316 9915
rect 5284 9884 5316 9885
rect 5284 9835 5316 9836
rect 5284 9805 5285 9835
rect 5285 9805 5315 9835
rect 5315 9805 5316 9835
rect 5284 9804 5316 9805
rect 5284 9755 5316 9756
rect 5284 9725 5285 9755
rect 5285 9725 5315 9755
rect 5315 9725 5316 9755
rect 5284 9724 5316 9725
rect 5284 9355 5316 9356
rect 5284 9325 5285 9355
rect 5285 9325 5315 9355
rect 5315 9325 5316 9355
rect 5284 9324 5316 9325
rect 5284 9275 5316 9276
rect 5284 9245 5285 9275
rect 5285 9245 5315 9275
rect 5315 9245 5316 9275
rect 5284 9244 5316 9245
rect 5284 9195 5316 9196
rect 5284 9165 5285 9195
rect 5285 9165 5315 9195
rect 5315 9165 5316 9195
rect 5284 9164 5316 9165
rect 5284 8875 5316 8876
rect 5284 8845 5285 8875
rect 5285 8845 5315 8875
rect 5315 8845 5316 8875
rect 5284 8844 5316 8845
rect 5284 8795 5316 8796
rect 5284 8765 5285 8795
rect 5285 8765 5315 8795
rect 5315 8765 5316 8795
rect 5284 8764 5316 8765
rect 5284 8715 5316 8716
rect 5284 8685 5285 8715
rect 5285 8685 5315 8715
rect 5315 8685 5316 8715
rect 5284 8684 5316 8685
rect 5284 8635 5316 8636
rect 5284 8605 5285 8635
rect 5285 8605 5315 8635
rect 5315 8605 5316 8635
rect 5284 8604 5316 8605
rect 5284 8555 5316 8556
rect 5284 8525 5285 8555
rect 5285 8525 5315 8555
rect 5315 8525 5316 8555
rect 5284 8524 5316 8525
rect 5284 7635 5316 7636
rect 5284 7605 5285 7635
rect 5285 7605 5315 7635
rect 5315 7605 5316 7635
rect 5284 7604 5316 7605
rect 5284 7555 5316 7556
rect 5284 7525 5285 7555
rect 5285 7525 5315 7555
rect 5315 7525 5316 7555
rect 5284 7524 5316 7525
rect 5284 7475 5316 7476
rect 5284 7445 5285 7475
rect 5285 7445 5315 7475
rect 5315 7445 5316 7475
rect 5284 7444 5316 7445
rect 5284 7395 5316 7396
rect 5284 7365 5285 7395
rect 5285 7365 5315 7395
rect 5315 7365 5316 7395
rect 5284 7364 5316 7365
rect 5284 7315 5316 7316
rect 5284 7285 5285 7315
rect 5285 7285 5315 7315
rect 5315 7285 5316 7315
rect 5284 7284 5316 7285
rect 5284 7235 5316 7236
rect 5284 7205 5285 7235
rect 5285 7205 5315 7235
rect 5315 7205 5316 7235
rect 5284 7204 5316 7205
rect 5284 7155 5316 7156
rect 5284 7125 5285 7155
rect 5285 7125 5315 7155
rect 5315 7125 5316 7155
rect 5284 7124 5316 7125
rect 5284 7075 5316 7076
rect 5284 7045 5285 7075
rect 5285 7045 5315 7075
rect 5315 7045 5316 7075
rect 5284 7044 5316 7045
rect 5284 6755 5316 6756
rect 5284 6725 5285 6755
rect 5285 6725 5315 6755
rect 5315 6725 5316 6755
rect 5284 6724 5316 6725
rect 5284 6675 5316 6676
rect 5284 6645 5285 6675
rect 5285 6645 5315 6675
rect 5315 6645 5316 6675
rect 5284 6644 5316 6645
rect 5284 6595 5316 6596
rect 5284 6565 5285 6595
rect 5285 6565 5315 6595
rect 5315 6565 5316 6595
rect 5284 6564 5316 6565
rect 5284 6515 5316 6516
rect 5284 6485 5285 6515
rect 5285 6485 5315 6515
rect 5315 6485 5316 6515
rect 5284 6484 5316 6485
rect 5284 6435 5316 6436
rect 5284 6405 5285 6435
rect 5285 6405 5315 6435
rect 5315 6405 5316 6435
rect 5284 6404 5316 6405
rect 5284 6355 5316 6356
rect 5284 6325 5285 6355
rect 5285 6325 5315 6355
rect 5315 6325 5316 6355
rect 5284 6324 5316 6325
rect 5284 5795 5316 5796
rect 5284 5765 5285 5795
rect 5285 5765 5315 5795
rect 5315 5765 5316 5795
rect 5284 5764 5316 5765
rect 5284 5715 5316 5716
rect 5284 5685 5285 5715
rect 5285 5685 5315 5715
rect 5315 5685 5316 5715
rect 5284 5684 5316 5685
rect 5284 5635 5316 5636
rect 5284 5605 5285 5635
rect 5285 5605 5315 5635
rect 5315 5605 5316 5635
rect 5284 5604 5316 5605
rect 5284 5555 5316 5556
rect 5284 5525 5285 5555
rect 5285 5525 5315 5555
rect 5315 5525 5316 5555
rect 5284 5524 5316 5525
rect 5284 5475 5316 5476
rect 5284 5445 5285 5475
rect 5285 5445 5315 5475
rect 5315 5445 5316 5475
rect 5284 5444 5316 5445
rect 5284 5395 5316 5396
rect 5284 5365 5285 5395
rect 5285 5365 5315 5395
rect 5315 5365 5316 5395
rect 5284 5364 5316 5365
rect 5284 5315 5316 5316
rect 5284 5285 5285 5315
rect 5285 5285 5315 5315
rect 5315 5285 5316 5315
rect 5284 5284 5316 5285
rect 5284 5235 5316 5236
rect 5284 5205 5285 5235
rect 5285 5205 5315 5235
rect 5315 5205 5316 5235
rect 5284 5204 5316 5205
rect 5284 5155 5316 5156
rect 5284 5125 5285 5155
rect 5285 5125 5315 5155
rect 5315 5125 5316 5155
rect 5284 5124 5316 5125
rect 5284 5075 5316 5076
rect 5284 5045 5285 5075
rect 5285 5045 5315 5075
rect 5315 5045 5316 5075
rect 5284 5044 5316 5045
rect 5284 4995 5316 4996
rect 5284 4965 5285 4995
rect 5285 4965 5315 4995
rect 5315 4965 5316 4995
rect 5284 4964 5316 4965
rect 5284 4435 5316 4436
rect 5284 4405 5285 4435
rect 5285 4405 5315 4435
rect 5315 4405 5316 4435
rect 5284 4404 5316 4405
rect 5284 4355 5316 4356
rect 5284 4325 5285 4355
rect 5285 4325 5315 4355
rect 5315 4325 5316 4355
rect 5284 4324 5316 4325
rect 5284 4275 5316 4276
rect 5284 4245 5285 4275
rect 5285 4245 5315 4275
rect 5315 4245 5316 4275
rect 5284 4244 5316 4245
rect 5284 4195 5316 4196
rect 5284 4165 5285 4195
rect 5285 4165 5315 4195
rect 5315 4165 5316 4195
rect 5284 4164 5316 4165
rect 5284 4115 5316 4116
rect 5284 4085 5285 4115
rect 5285 4085 5315 4115
rect 5315 4085 5316 4115
rect 5284 4084 5316 4085
rect 5284 4035 5316 4036
rect 5284 4005 5285 4035
rect 5285 4005 5315 4035
rect 5315 4005 5316 4035
rect 5284 4004 5316 4005
rect 5284 3955 5316 3956
rect 5284 3925 5285 3955
rect 5285 3925 5315 3955
rect 5315 3925 5316 3955
rect 5284 3924 5316 3925
rect 5284 3155 5316 3156
rect 5284 3125 5285 3155
rect 5285 3125 5315 3155
rect 5315 3125 5316 3155
rect 5284 3124 5316 3125
rect 5284 3075 5316 3076
rect 5284 3045 5285 3075
rect 5285 3045 5315 3075
rect 5315 3045 5316 3075
rect 5284 3044 5316 3045
rect 5284 2995 5316 2996
rect 5284 2965 5285 2995
rect 5285 2965 5315 2995
rect 5315 2965 5316 2995
rect 5284 2964 5316 2965
rect 5284 2915 5316 2916
rect 5284 2885 5285 2915
rect 5285 2885 5315 2915
rect 5315 2885 5316 2915
rect 5284 2884 5316 2885
rect 5284 2835 5316 2836
rect 5284 2805 5285 2835
rect 5285 2805 5315 2835
rect 5315 2805 5316 2835
rect 5284 2804 5316 2805
rect 5284 2755 5316 2756
rect 5284 2725 5285 2755
rect 5285 2725 5315 2755
rect 5315 2725 5316 2755
rect 5284 2724 5316 2725
rect 5284 2675 5316 2676
rect 5284 2645 5285 2675
rect 5285 2645 5315 2675
rect 5315 2645 5316 2675
rect 5284 2644 5316 2645
rect 5284 2595 5316 2596
rect 5284 2565 5285 2595
rect 5285 2565 5315 2595
rect 5315 2565 5316 2595
rect 5284 2564 5316 2565
rect 5284 2515 5316 2516
rect 5284 2485 5285 2515
rect 5285 2485 5315 2515
rect 5315 2485 5316 2515
rect 5284 2484 5316 2485
rect 5284 2435 5316 2436
rect 5284 2405 5285 2435
rect 5285 2405 5315 2435
rect 5315 2405 5316 2435
rect 5284 2404 5316 2405
rect 5284 2355 5316 2356
rect 5284 2325 5285 2355
rect 5285 2325 5315 2355
rect 5315 2325 5316 2355
rect 5284 2324 5316 2325
rect 5284 2275 5316 2276
rect 5284 2245 5285 2275
rect 5285 2245 5315 2275
rect 5315 2245 5316 2275
rect 5284 2244 5316 2245
rect 5284 2195 5316 2196
rect 5284 2165 5285 2195
rect 5285 2165 5315 2195
rect 5315 2165 5316 2195
rect 5284 2164 5316 2165
rect 5284 2115 5316 2116
rect 5284 2085 5285 2115
rect 5285 2085 5315 2115
rect 5315 2085 5316 2115
rect 5284 2084 5316 2085
rect 5284 2035 5316 2036
rect 5284 2005 5285 2035
rect 5285 2005 5315 2035
rect 5315 2005 5316 2035
rect 5284 2004 5316 2005
rect 5284 1635 5316 1636
rect 5284 1605 5285 1635
rect 5285 1605 5315 1635
rect 5315 1605 5316 1635
rect 5284 1604 5316 1605
rect 5284 1555 5316 1556
rect 5284 1525 5285 1555
rect 5285 1525 5315 1555
rect 5315 1525 5316 1555
rect 5284 1524 5316 1525
rect 5284 1475 5316 1476
rect 5284 1445 5285 1475
rect 5285 1445 5315 1475
rect 5315 1445 5316 1475
rect 5284 1444 5316 1445
rect 5284 1395 5316 1396
rect 5284 1365 5285 1395
rect 5285 1365 5315 1395
rect 5315 1365 5316 1395
rect 5284 1364 5316 1365
rect 5284 1315 5316 1316
rect 5284 1285 5285 1315
rect 5285 1285 5315 1315
rect 5315 1285 5316 1315
rect 5284 1284 5316 1285
rect 5284 1235 5316 1236
rect 5284 1205 5285 1235
rect 5285 1205 5315 1235
rect 5315 1205 5316 1235
rect 5284 1204 5316 1205
rect 5284 1155 5316 1156
rect 5284 1125 5285 1155
rect 5285 1125 5315 1155
rect 5315 1125 5316 1155
rect 5284 1124 5316 1125
rect 5284 1075 5316 1076
rect 5284 1045 5285 1075
rect 5285 1045 5315 1075
rect 5315 1045 5316 1075
rect 5284 1044 5316 1045
rect 5284 755 5316 756
rect 5284 725 5285 755
rect 5285 725 5315 755
rect 5315 725 5316 755
rect 5284 724 5316 725
rect 5284 675 5316 676
rect 5284 645 5285 675
rect 5285 645 5315 675
rect 5315 645 5316 675
rect 5284 644 5316 645
rect 5284 595 5316 596
rect 5284 565 5285 595
rect 5285 565 5315 595
rect 5315 565 5316 595
rect 5284 564 5316 565
rect 5284 195 5316 196
rect 5284 165 5285 195
rect 5285 165 5315 195
rect 5315 165 5316 195
rect 5284 164 5316 165
rect 5284 115 5316 116
rect 5284 85 5285 115
rect 5285 85 5315 115
rect 5315 85 5316 115
rect 5284 84 5316 85
rect 5284 35 5316 36
rect 5284 5 5285 35
rect 5285 5 5315 35
rect 5315 5 5316 35
rect 5284 4 5316 5
rect 5364 15284 5396 15316
rect 5444 15364 5476 15396
rect 5444 14084 5476 14116
rect 5444 12635 5476 12636
rect 5444 12605 5445 12635
rect 5445 12605 5475 12635
rect 5475 12605 5476 12635
rect 5444 12604 5476 12605
rect 5444 12555 5476 12556
rect 5444 12525 5445 12555
rect 5445 12525 5475 12555
rect 5475 12525 5476 12555
rect 5444 12524 5476 12525
rect 5444 12475 5476 12476
rect 5444 12445 5445 12475
rect 5445 12445 5475 12475
rect 5475 12445 5476 12475
rect 5444 12444 5476 12445
rect 5444 12395 5476 12396
rect 5444 12365 5445 12395
rect 5445 12365 5475 12395
rect 5475 12365 5476 12395
rect 5444 12364 5476 12365
rect 5444 12315 5476 12316
rect 5444 12285 5445 12315
rect 5445 12285 5475 12315
rect 5475 12285 5476 12315
rect 5444 12284 5476 12285
rect 5444 12235 5476 12236
rect 5444 12205 5445 12235
rect 5445 12205 5475 12235
rect 5475 12205 5476 12235
rect 5444 12204 5476 12205
rect 5444 12155 5476 12156
rect 5444 12125 5445 12155
rect 5445 12125 5475 12155
rect 5475 12125 5476 12155
rect 5444 12124 5476 12125
rect 5444 11835 5476 11836
rect 5444 11805 5445 11835
rect 5445 11805 5475 11835
rect 5475 11805 5476 11835
rect 5444 11804 5476 11805
rect 5444 11755 5476 11756
rect 5444 11725 5445 11755
rect 5445 11725 5475 11755
rect 5475 11725 5476 11755
rect 5444 11724 5476 11725
rect 5444 11675 5476 11676
rect 5444 11645 5445 11675
rect 5445 11645 5475 11675
rect 5475 11645 5476 11675
rect 5444 11644 5476 11645
rect 5444 11595 5476 11596
rect 5444 11565 5445 11595
rect 5445 11565 5475 11595
rect 5475 11565 5476 11595
rect 5444 11564 5476 11565
rect 5444 11515 5476 11516
rect 5444 11485 5445 11515
rect 5445 11485 5475 11515
rect 5475 11485 5476 11515
rect 5444 11484 5476 11485
rect 5444 11435 5476 11436
rect 5444 11405 5445 11435
rect 5445 11405 5475 11435
rect 5475 11405 5476 11435
rect 5444 11404 5476 11405
rect 5444 10875 5476 10876
rect 5444 10845 5445 10875
rect 5445 10845 5475 10875
rect 5475 10845 5476 10875
rect 5444 10844 5476 10845
rect 5444 10795 5476 10796
rect 5444 10765 5445 10795
rect 5445 10765 5475 10795
rect 5475 10765 5476 10795
rect 5444 10764 5476 10765
rect 5444 10715 5476 10716
rect 5444 10685 5445 10715
rect 5445 10685 5475 10715
rect 5475 10685 5476 10715
rect 5444 10684 5476 10685
rect 5444 10635 5476 10636
rect 5444 10605 5445 10635
rect 5445 10605 5475 10635
rect 5475 10605 5476 10635
rect 5444 10604 5476 10605
rect 5444 10555 5476 10556
rect 5444 10525 5445 10555
rect 5445 10525 5475 10555
rect 5475 10525 5476 10555
rect 5444 10524 5476 10525
rect 5444 10475 5476 10476
rect 5444 10445 5445 10475
rect 5445 10445 5475 10475
rect 5475 10445 5476 10475
rect 5444 10444 5476 10445
rect 5444 10395 5476 10396
rect 5444 10365 5445 10395
rect 5445 10365 5475 10395
rect 5475 10365 5476 10395
rect 5444 10364 5476 10365
rect 5444 10315 5476 10316
rect 5444 10285 5445 10315
rect 5445 10285 5475 10315
rect 5475 10285 5476 10315
rect 5444 10284 5476 10285
rect 5444 10235 5476 10236
rect 5444 10205 5445 10235
rect 5445 10205 5475 10235
rect 5475 10205 5476 10235
rect 5444 10204 5476 10205
rect 5444 10155 5476 10156
rect 5444 10125 5445 10155
rect 5445 10125 5475 10155
rect 5475 10125 5476 10155
rect 5444 10124 5476 10125
rect 5444 10075 5476 10076
rect 5444 10045 5445 10075
rect 5445 10045 5475 10075
rect 5475 10045 5476 10075
rect 5444 10044 5476 10045
rect 5444 9995 5476 9996
rect 5444 9965 5445 9995
rect 5445 9965 5475 9995
rect 5475 9965 5476 9995
rect 5444 9964 5476 9965
rect 5444 9915 5476 9916
rect 5444 9885 5445 9915
rect 5445 9885 5475 9915
rect 5475 9885 5476 9915
rect 5444 9884 5476 9885
rect 5444 9835 5476 9836
rect 5444 9805 5445 9835
rect 5445 9805 5475 9835
rect 5475 9805 5476 9835
rect 5444 9804 5476 9805
rect 5444 9755 5476 9756
rect 5444 9725 5445 9755
rect 5445 9725 5475 9755
rect 5475 9725 5476 9755
rect 5444 9724 5476 9725
rect 5444 9355 5476 9356
rect 5444 9325 5445 9355
rect 5445 9325 5475 9355
rect 5475 9325 5476 9355
rect 5444 9324 5476 9325
rect 5444 9275 5476 9276
rect 5444 9245 5445 9275
rect 5445 9245 5475 9275
rect 5475 9245 5476 9275
rect 5444 9244 5476 9245
rect 5444 9195 5476 9196
rect 5444 9165 5445 9195
rect 5445 9165 5475 9195
rect 5475 9165 5476 9195
rect 5444 9164 5476 9165
rect 5444 8875 5476 8876
rect 5444 8845 5445 8875
rect 5445 8845 5475 8875
rect 5475 8845 5476 8875
rect 5444 8844 5476 8845
rect 5444 8795 5476 8796
rect 5444 8765 5445 8795
rect 5445 8765 5475 8795
rect 5475 8765 5476 8795
rect 5444 8764 5476 8765
rect 5444 8715 5476 8716
rect 5444 8685 5445 8715
rect 5445 8685 5475 8715
rect 5475 8685 5476 8715
rect 5444 8684 5476 8685
rect 5444 8635 5476 8636
rect 5444 8605 5445 8635
rect 5445 8605 5475 8635
rect 5475 8605 5476 8635
rect 5444 8604 5476 8605
rect 5444 8555 5476 8556
rect 5444 8525 5445 8555
rect 5445 8525 5475 8555
rect 5475 8525 5476 8555
rect 5444 8524 5476 8525
rect 5444 7635 5476 7636
rect 5444 7605 5445 7635
rect 5445 7605 5475 7635
rect 5475 7605 5476 7635
rect 5444 7604 5476 7605
rect 5444 7555 5476 7556
rect 5444 7525 5445 7555
rect 5445 7525 5475 7555
rect 5475 7525 5476 7555
rect 5444 7524 5476 7525
rect 5444 7475 5476 7476
rect 5444 7445 5445 7475
rect 5445 7445 5475 7475
rect 5475 7445 5476 7475
rect 5444 7444 5476 7445
rect 5444 7395 5476 7396
rect 5444 7365 5445 7395
rect 5445 7365 5475 7395
rect 5475 7365 5476 7395
rect 5444 7364 5476 7365
rect 5444 7315 5476 7316
rect 5444 7285 5445 7315
rect 5445 7285 5475 7315
rect 5475 7285 5476 7315
rect 5444 7284 5476 7285
rect 5444 7235 5476 7236
rect 5444 7205 5445 7235
rect 5445 7205 5475 7235
rect 5475 7205 5476 7235
rect 5444 7204 5476 7205
rect 5444 7155 5476 7156
rect 5444 7125 5445 7155
rect 5445 7125 5475 7155
rect 5475 7125 5476 7155
rect 5444 7124 5476 7125
rect 5444 7075 5476 7076
rect 5444 7045 5445 7075
rect 5445 7045 5475 7075
rect 5475 7045 5476 7075
rect 5444 7044 5476 7045
rect 5444 6755 5476 6756
rect 5444 6725 5445 6755
rect 5445 6725 5475 6755
rect 5475 6725 5476 6755
rect 5444 6724 5476 6725
rect 5444 6675 5476 6676
rect 5444 6645 5445 6675
rect 5445 6645 5475 6675
rect 5475 6645 5476 6675
rect 5444 6644 5476 6645
rect 5444 6595 5476 6596
rect 5444 6565 5445 6595
rect 5445 6565 5475 6595
rect 5475 6565 5476 6595
rect 5444 6564 5476 6565
rect 5444 6515 5476 6516
rect 5444 6485 5445 6515
rect 5445 6485 5475 6515
rect 5475 6485 5476 6515
rect 5444 6484 5476 6485
rect 5444 6435 5476 6436
rect 5444 6405 5445 6435
rect 5445 6405 5475 6435
rect 5475 6405 5476 6435
rect 5444 6404 5476 6405
rect 5444 6355 5476 6356
rect 5444 6325 5445 6355
rect 5445 6325 5475 6355
rect 5475 6325 5476 6355
rect 5444 6324 5476 6325
rect 5444 5795 5476 5796
rect 5444 5765 5445 5795
rect 5445 5765 5475 5795
rect 5475 5765 5476 5795
rect 5444 5764 5476 5765
rect 5444 5715 5476 5716
rect 5444 5685 5445 5715
rect 5445 5685 5475 5715
rect 5475 5685 5476 5715
rect 5444 5684 5476 5685
rect 5444 5635 5476 5636
rect 5444 5605 5445 5635
rect 5445 5605 5475 5635
rect 5475 5605 5476 5635
rect 5444 5604 5476 5605
rect 5444 5555 5476 5556
rect 5444 5525 5445 5555
rect 5445 5525 5475 5555
rect 5475 5525 5476 5555
rect 5444 5524 5476 5525
rect 5444 5475 5476 5476
rect 5444 5445 5445 5475
rect 5445 5445 5475 5475
rect 5475 5445 5476 5475
rect 5444 5444 5476 5445
rect 5444 5395 5476 5396
rect 5444 5365 5445 5395
rect 5445 5365 5475 5395
rect 5475 5365 5476 5395
rect 5444 5364 5476 5365
rect 5444 5315 5476 5316
rect 5444 5285 5445 5315
rect 5445 5285 5475 5315
rect 5475 5285 5476 5315
rect 5444 5284 5476 5285
rect 5444 5235 5476 5236
rect 5444 5205 5445 5235
rect 5445 5205 5475 5235
rect 5475 5205 5476 5235
rect 5444 5204 5476 5205
rect 5444 5155 5476 5156
rect 5444 5125 5445 5155
rect 5445 5125 5475 5155
rect 5475 5125 5476 5155
rect 5444 5124 5476 5125
rect 5444 5075 5476 5076
rect 5444 5045 5445 5075
rect 5445 5045 5475 5075
rect 5475 5045 5476 5075
rect 5444 5044 5476 5045
rect 5444 4995 5476 4996
rect 5444 4965 5445 4995
rect 5445 4965 5475 4995
rect 5475 4965 5476 4995
rect 5444 4964 5476 4965
rect 5444 4435 5476 4436
rect 5444 4405 5445 4435
rect 5445 4405 5475 4435
rect 5475 4405 5476 4435
rect 5444 4404 5476 4405
rect 5444 4355 5476 4356
rect 5444 4325 5445 4355
rect 5445 4325 5475 4355
rect 5475 4325 5476 4355
rect 5444 4324 5476 4325
rect 5444 4275 5476 4276
rect 5444 4245 5445 4275
rect 5445 4245 5475 4275
rect 5475 4245 5476 4275
rect 5444 4244 5476 4245
rect 5444 4195 5476 4196
rect 5444 4165 5445 4195
rect 5445 4165 5475 4195
rect 5475 4165 5476 4195
rect 5444 4164 5476 4165
rect 5444 4115 5476 4116
rect 5444 4085 5445 4115
rect 5445 4085 5475 4115
rect 5475 4085 5476 4115
rect 5444 4084 5476 4085
rect 5444 4035 5476 4036
rect 5444 4005 5445 4035
rect 5445 4005 5475 4035
rect 5475 4005 5476 4035
rect 5444 4004 5476 4005
rect 5444 3955 5476 3956
rect 5444 3925 5445 3955
rect 5445 3925 5475 3955
rect 5475 3925 5476 3955
rect 5444 3924 5476 3925
rect 5444 3155 5476 3156
rect 5444 3125 5445 3155
rect 5445 3125 5475 3155
rect 5475 3125 5476 3155
rect 5444 3124 5476 3125
rect 5444 3075 5476 3076
rect 5444 3045 5445 3075
rect 5445 3045 5475 3075
rect 5475 3045 5476 3075
rect 5444 3044 5476 3045
rect 5444 2995 5476 2996
rect 5444 2965 5445 2995
rect 5445 2965 5475 2995
rect 5475 2965 5476 2995
rect 5444 2964 5476 2965
rect 5444 2915 5476 2916
rect 5444 2885 5445 2915
rect 5445 2885 5475 2915
rect 5475 2885 5476 2915
rect 5444 2884 5476 2885
rect 5444 2835 5476 2836
rect 5444 2805 5445 2835
rect 5445 2805 5475 2835
rect 5475 2805 5476 2835
rect 5444 2804 5476 2805
rect 5444 2755 5476 2756
rect 5444 2725 5445 2755
rect 5445 2725 5475 2755
rect 5475 2725 5476 2755
rect 5444 2724 5476 2725
rect 5444 2675 5476 2676
rect 5444 2645 5445 2675
rect 5445 2645 5475 2675
rect 5475 2645 5476 2675
rect 5444 2644 5476 2645
rect 5444 2595 5476 2596
rect 5444 2565 5445 2595
rect 5445 2565 5475 2595
rect 5475 2565 5476 2595
rect 5444 2564 5476 2565
rect 5444 2515 5476 2516
rect 5444 2485 5445 2515
rect 5445 2485 5475 2515
rect 5475 2485 5476 2515
rect 5444 2484 5476 2485
rect 5444 2435 5476 2436
rect 5444 2405 5445 2435
rect 5445 2405 5475 2435
rect 5475 2405 5476 2435
rect 5444 2404 5476 2405
rect 5444 2355 5476 2356
rect 5444 2325 5445 2355
rect 5445 2325 5475 2355
rect 5475 2325 5476 2355
rect 5444 2324 5476 2325
rect 5444 2275 5476 2276
rect 5444 2245 5445 2275
rect 5445 2245 5475 2275
rect 5475 2245 5476 2275
rect 5444 2244 5476 2245
rect 5444 2195 5476 2196
rect 5444 2165 5445 2195
rect 5445 2165 5475 2195
rect 5475 2165 5476 2195
rect 5444 2164 5476 2165
rect 5444 2115 5476 2116
rect 5444 2085 5445 2115
rect 5445 2085 5475 2115
rect 5475 2085 5476 2115
rect 5444 2084 5476 2085
rect 5444 2035 5476 2036
rect 5444 2005 5445 2035
rect 5445 2005 5475 2035
rect 5475 2005 5476 2035
rect 5444 2004 5476 2005
rect 5444 1635 5476 1636
rect 5444 1605 5445 1635
rect 5445 1605 5475 1635
rect 5475 1605 5476 1635
rect 5444 1604 5476 1605
rect 5444 1555 5476 1556
rect 5444 1525 5445 1555
rect 5445 1525 5475 1555
rect 5475 1525 5476 1555
rect 5444 1524 5476 1525
rect 5444 1475 5476 1476
rect 5444 1445 5445 1475
rect 5445 1445 5475 1475
rect 5475 1445 5476 1475
rect 5444 1444 5476 1445
rect 5444 1395 5476 1396
rect 5444 1365 5445 1395
rect 5445 1365 5475 1395
rect 5475 1365 5476 1395
rect 5444 1364 5476 1365
rect 5444 1315 5476 1316
rect 5444 1285 5445 1315
rect 5445 1285 5475 1315
rect 5475 1285 5476 1315
rect 5444 1284 5476 1285
rect 5444 1235 5476 1236
rect 5444 1205 5445 1235
rect 5445 1205 5475 1235
rect 5475 1205 5476 1235
rect 5444 1204 5476 1205
rect 5444 1155 5476 1156
rect 5444 1125 5445 1155
rect 5445 1125 5475 1155
rect 5475 1125 5476 1155
rect 5444 1124 5476 1125
rect 5444 1075 5476 1076
rect 5444 1045 5445 1075
rect 5445 1045 5475 1075
rect 5475 1045 5476 1075
rect 5444 1044 5476 1045
rect 5444 755 5476 756
rect 5444 725 5445 755
rect 5445 725 5475 755
rect 5475 725 5476 755
rect 5444 724 5476 725
rect 5444 675 5476 676
rect 5444 645 5445 675
rect 5445 645 5475 675
rect 5475 645 5476 675
rect 5444 644 5476 645
rect 5444 595 5476 596
rect 5444 565 5445 595
rect 5445 565 5475 595
rect 5475 565 5476 595
rect 5444 564 5476 565
rect 5444 195 5476 196
rect 5444 165 5445 195
rect 5445 165 5475 195
rect 5475 165 5476 195
rect 5444 164 5476 165
rect 5444 115 5476 116
rect 5444 85 5445 115
rect 5445 85 5475 115
rect 5475 85 5476 115
rect 5444 84 5476 85
rect 5444 35 5476 36
rect 5444 5 5445 35
rect 5445 5 5475 35
rect 5475 5 5476 35
rect 5444 4 5476 5
rect 5604 15364 5636 15396
rect 10164 15364 10196 15396
rect 5684 15284 5716 15316
rect 6724 15284 6756 15316
rect 6804 15284 6836 15316
rect 7844 15284 7876 15316
rect 7924 15284 7956 15316
rect 8964 15284 8996 15316
rect 9044 15284 9076 15316
rect 10084 15284 10116 15316
rect 5604 14084 5636 14116
rect 10164 14084 10196 14116
rect 5524 14004 5556 14036
rect 5524 13684 5556 13716
rect 10244 14004 10276 14036
rect 10324 16804 10356 16836
rect 10324 15524 10356 15556
rect 10324 13924 10356 13956
rect 10324 13764 10356 13796
rect 10404 16724 10436 16756
rect 10404 13844 10436 13876
rect 10484 16804 10516 16836
rect 10484 15524 10516 15556
rect 10484 13924 10516 13956
rect 10484 13764 10516 13796
rect 10564 16884 10596 16916
rect 10564 15444 10596 15476
rect 10564 14004 10596 14036
rect 10244 13684 10276 13716
rect 10564 13684 10596 13716
rect 5524 13204 5556 13396
rect 5684 13204 5716 13396
rect 5524 12635 5556 12636
rect 5524 12605 5525 12635
rect 5525 12605 5555 12635
rect 5555 12605 5556 12635
rect 5524 12604 5556 12605
rect 5524 12555 5556 12556
rect 5524 12525 5525 12555
rect 5525 12525 5555 12555
rect 5555 12525 5556 12555
rect 5524 12524 5556 12525
rect 5524 12475 5556 12476
rect 5524 12445 5525 12475
rect 5525 12445 5555 12475
rect 5555 12445 5556 12475
rect 5524 12444 5556 12445
rect 5524 12395 5556 12396
rect 5524 12365 5525 12395
rect 5525 12365 5555 12395
rect 5555 12365 5556 12395
rect 5524 12364 5556 12365
rect 5524 12315 5556 12316
rect 5524 12285 5525 12315
rect 5525 12285 5555 12315
rect 5555 12285 5556 12315
rect 5524 12284 5556 12285
rect 5524 12235 5556 12236
rect 5524 12205 5525 12235
rect 5525 12205 5555 12235
rect 5555 12205 5556 12235
rect 5524 12204 5556 12205
rect 5524 12155 5556 12156
rect 5524 12125 5525 12155
rect 5525 12125 5555 12155
rect 5555 12125 5556 12155
rect 5524 12124 5556 12125
rect 5524 11835 5556 11836
rect 5524 11805 5525 11835
rect 5525 11805 5555 11835
rect 5555 11805 5556 11835
rect 5524 11804 5556 11805
rect 5524 11755 5556 11756
rect 5524 11725 5525 11755
rect 5525 11725 5555 11755
rect 5555 11725 5556 11755
rect 5524 11724 5556 11725
rect 5524 11675 5556 11676
rect 5524 11645 5525 11675
rect 5525 11645 5555 11675
rect 5555 11645 5556 11675
rect 5524 11644 5556 11645
rect 5524 11595 5556 11596
rect 5524 11565 5525 11595
rect 5525 11565 5555 11595
rect 5555 11565 5556 11595
rect 5524 11564 5556 11565
rect 5524 11515 5556 11516
rect 5524 11485 5525 11515
rect 5525 11485 5555 11515
rect 5555 11485 5556 11515
rect 5524 11484 5556 11485
rect 5524 11435 5556 11436
rect 5524 11405 5525 11435
rect 5525 11405 5555 11435
rect 5555 11405 5556 11435
rect 5524 11404 5556 11405
rect 5524 10875 5556 10876
rect 5524 10845 5525 10875
rect 5525 10845 5555 10875
rect 5555 10845 5556 10875
rect 5524 10844 5556 10845
rect 5524 10795 5556 10796
rect 5524 10765 5525 10795
rect 5525 10765 5555 10795
rect 5555 10765 5556 10795
rect 5524 10764 5556 10765
rect 5524 10715 5556 10716
rect 5524 10685 5525 10715
rect 5525 10685 5555 10715
rect 5555 10685 5556 10715
rect 5524 10684 5556 10685
rect 5524 10635 5556 10636
rect 5524 10605 5525 10635
rect 5525 10605 5555 10635
rect 5555 10605 5556 10635
rect 5524 10604 5556 10605
rect 5524 10555 5556 10556
rect 5524 10525 5525 10555
rect 5525 10525 5555 10555
rect 5555 10525 5556 10555
rect 5524 10524 5556 10525
rect 5524 10475 5556 10476
rect 5524 10445 5525 10475
rect 5525 10445 5555 10475
rect 5555 10445 5556 10475
rect 5524 10444 5556 10445
rect 5524 10395 5556 10396
rect 5524 10365 5525 10395
rect 5525 10365 5555 10395
rect 5555 10365 5556 10395
rect 5524 10364 5556 10365
rect 5524 10315 5556 10316
rect 5524 10285 5525 10315
rect 5525 10285 5555 10315
rect 5555 10285 5556 10315
rect 5524 10284 5556 10285
rect 5524 10235 5556 10236
rect 5524 10205 5525 10235
rect 5525 10205 5555 10235
rect 5555 10205 5556 10235
rect 5524 10204 5556 10205
rect 5524 10155 5556 10156
rect 5524 10125 5525 10155
rect 5525 10125 5555 10155
rect 5555 10125 5556 10155
rect 5524 10124 5556 10125
rect 5524 10075 5556 10076
rect 5524 10045 5525 10075
rect 5525 10045 5555 10075
rect 5555 10045 5556 10075
rect 5524 10044 5556 10045
rect 5524 9995 5556 9996
rect 5524 9965 5525 9995
rect 5525 9965 5555 9995
rect 5555 9965 5556 9995
rect 5524 9964 5556 9965
rect 5524 9915 5556 9916
rect 5524 9885 5525 9915
rect 5525 9885 5555 9915
rect 5555 9885 5556 9915
rect 5524 9884 5556 9885
rect 5524 9835 5556 9836
rect 5524 9805 5525 9835
rect 5525 9805 5555 9835
rect 5555 9805 5556 9835
rect 5524 9804 5556 9805
rect 5524 9755 5556 9756
rect 5524 9725 5525 9755
rect 5525 9725 5555 9755
rect 5555 9725 5556 9755
rect 5524 9724 5556 9725
rect 5524 9355 5556 9356
rect 5524 9325 5525 9355
rect 5525 9325 5555 9355
rect 5555 9325 5556 9355
rect 5524 9324 5556 9325
rect 5524 9275 5556 9276
rect 5524 9245 5525 9275
rect 5525 9245 5555 9275
rect 5555 9245 5556 9275
rect 5524 9244 5556 9245
rect 5524 9195 5556 9196
rect 5524 9165 5525 9195
rect 5525 9165 5555 9195
rect 5555 9165 5556 9195
rect 5524 9164 5556 9165
rect 5524 8875 5556 8876
rect 5524 8845 5525 8875
rect 5525 8845 5555 8875
rect 5555 8845 5556 8875
rect 5524 8844 5556 8845
rect 5524 8795 5556 8796
rect 5524 8765 5525 8795
rect 5525 8765 5555 8795
rect 5555 8765 5556 8795
rect 5524 8764 5556 8765
rect 5524 8715 5556 8716
rect 5524 8685 5525 8715
rect 5525 8685 5555 8715
rect 5555 8685 5556 8715
rect 5524 8684 5556 8685
rect 5524 8635 5556 8636
rect 5524 8605 5525 8635
rect 5525 8605 5555 8635
rect 5555 8605 5556 8635
rect 5524 8604 5556 8605
rect 5524 8555 5556 8556
rect 5524 8525 5525 8555
rect 5525 8525 5555 8555
rect 5555 8525 5556 8555
rect 5524 8524 5556 8525
rect 5524 7635 5556 7636
rect 5524 7605 5525 7635
rect 5525 7605 5555 7635
rect 5555 7605 5556 7635
rect 5524 7604 5556 7605
rect 5524 7555 5556 7556
rect 5524 7525 5525 7555
rect 5525 7525 5555 7555
rect 5555 7525 5556 7555
rect 5524 7524 5556 7525
rect 5524 7475 5556 7476
rect 5524 7445 5525 7475
rect 5525 7445 5555 7475
rect 5555 7445 5556 7475
rect 5524 7444 5556 7445
rect 5524 7395 5556 7396
rect 5524 7365 5525 7395
rect 5525 7365 5555 7395
rect 5555 7365 5556 7395
rect 5524 7364 5556 7365
rect 5524 7315 5556 7316
rect 5524 7285 5525 7315
rect 5525 7285 5555 7315
rect 5555 7285 5556 7315
rect 5524 7284 5556 7285
rect 5524 7235 5556 7236
rect 5524 7205 5525 7235
rect 5525 7205 5555 7235
rect 5555 7205 5556 7235
rect 5524 7204 5556 7205
rect 5524 7155 5556 7156
rect 5524 7125 5525 7155
rect 5525 7125 5555 7155
rect 5555 7125 5556 7155
rect 5524 7124 5556 7125
rect 5524 7075 5556 7076
rect 5524 7045 5525 7075
rect 5525 7045 5555 7075
rect 5555 7045 5556 7075
rect 5524 7044 5556 7045
rect 5524 6755 5556 6756
rect 5524 6725 5525 6755
rect 5525 6725 5555 6755
rect 5555 6725 5556 6755
rect 5524 6724 5556 6725
rect 5524 6675 5556 6676
rect 5524 6645 5525 6675
rect 5525 6645 5555 6675
rect 5555 6645 5556 6675
rect 5524 6644 5556 6645
rect 5524 6595 5556 6596
rect 5524 6565 5525 6595
rect 5525 6565 5555 6595
rect 5555 6565 5556 6595
rect 5524 6564 5556 6565
rect 5524 6515 5556 6516
rect 5524 6485 5525 6515
rect 5525 6485 5555 6515
rect 5555 6485 5556 6515
rect 5524 6484 5556 6485
rect 5524 6435 5556 6436
rect 5524 6405 5525 6435
rect 5525 6405 5555 6435
rect 5555 6405 5556 6435
rect 5524 6404 5556 6405
rect 5524 6355 5556 6356
rect 5524 6325 5525 6355
rect 5525 6325 5555 6355
rect 5555 6325 5556 6355
rect 5524 6324 5556 6325
rect 5524 5795 5556 5796
rect 5524 5765 5525 5795
rect 5525 5765 5555 5795
rect 5555 5765 5556 5795
rect 5524 5764 5556 5765
rect 5524 5715 5556 5716
rect 5524 5685 5525 5715
rect 5525 5685 5555 5715
rect 5555 5685 5556 5715
rect 5524 5684 5556 5685
rect 5524 5635 5556 5636
rect 5524 5605 5525 5635
rect 5525 5605 5555 5635
rect 5555 5605 5556 5635
rect 5524 5604 5556 5605
rect 5524 5555 5556 5556
rect 5524 5525 5525 5555
rect 5525 5525 5555 5555
rect 5555 5525 5556 5555
rect 5524 5524 5556 5525
rect 5524 5475 5556 5476
rect 5524 5445 5525 5475
rect 5525 5445 5555 5475
rect 5555 5445 5556 5475
rect 5524 5444 5556 5445
rect 5524 5395 5556 5396
rect 5524 5365 5525 5395
rect 5525 5365 5555 5395
rect 5555 5365 5556 5395
rect 5524 5364 5556 5365
rect 5524 5315 5556 5316
rect 5524 5285 5525 5315
rect 5525 5285 5555 5315
rect 5555 5285 5556 5315
rect 5524 5284 5556 5285
rect 5524 5235 5556 5236
rect 5524 5205 5525 5235
rect 5525 5205 5555 5235
rect 5555 5205 5556 5235
rect 5524 5204 5556 5205
rect 5524 5155 5556 5156
rect 5524 5125 5525 5155
rect 5525 5125 5555 5155
rect 5555 5125 5556 5155
rect 5524 5124 5556 5125
rect 5524 5075 5556 5076
rect 5524 5045 5525 5075
rect 5525 5045 5555 5075
rect 5555 5045 5556 5075
rect 5524 5044 5556 5045
rect 5524 4995 5556 4996
rect 5524 4965 5525 4995
rect 5525 4965 5555 4995
rect 5555 4965 5556 4995
rect 5524 4964 5556 4965
rect 5524 4435 5556 4436
rect 5524 4405 5525 4435
rect 5525 4405 5555 4435
rect 5555 4405 5556 4435
rect 5524 4404 5556 4405
rect 5524 4355 5556 4356
rect 5524 4325 5525 4355
rect 5525 4325 5555 4355
rect 5555 4325 5556 4355
rect 5524 4324 5556 4325
rect 5524 4275 5556 4276
rect 5524 4245 5525 4275
rect 5525 4245 5555 4275
rect 5555 4245 5556 4275
rect 5524 4244 5556 4245
rect 5524 4195 5556 4196
rect 5524 4165 5525 4195
rect 5525 4165 5555 4195
rect 5555 4165 5556 4195
rect 5524 4164 5556 4165
rect 5524 4115 5556 4116
rect 5524 4085 5525 4115
rect 5525 4085 5555 4115
rect 5555 4085 5556 4115
rect 5524 4084 5556 4085
rect 5524 4035 5556 4036
rect 5524 4005 5525 4035
rect 5525 4005 5555 4035
rect 5555 4005 5556 4035
rect 5524 4004 5556 4005
rect 5524 3955 5556 3956
rect 5524 3925 5525 3955
rect 5525 3925 5555 3955
rect 5555 3925 5556 3955
rect 5524 3924 5556 3925
rect 5524 3155 5556 3156
rect 5524 3125 5525 3155
rect 5525 3125 5555 3155
rect 5555 3125 5556 3155
rect 5524 3124 5556 3125
rect 5524 3075 5556 3076
rect 5524 3045 5525 3075
rect 5525 3045 5555 3075
rect 5555 3045 5556 3075
rect 5524 3044 5556 3045
rect 5524 2995 5556 2996
rect 5524 2965 5525 2995
rect 5525 2965 5555 2995
rect 5555 2965 5556 2995
rect 5524 2964 5556 2965
rect 5524 2915 5556 2916
rect 5524 2885 5525 2915
rect 5525 2885 5555 2915
rect 5555 2885 5556 2915
rect 5524 2884 5556 2885
rect 5524 2835 5556 2836
rect 5524 2805 5525 2835
rect 5525 2805 5555 2835
rect 5555 2805 5556 2835
rect 5524 2804 5556 2805
rect 5524 2755 5556 2756
rect 5524 2725 5525 2755
rect 5525 2725 5555 2755
rect 5555 2725 5556 2755
rect 5524 2724 5556 2725
rect 5524 2675 5556 2676
rect 5524 2645 5525 2675
rect 5525 2645 5555 2675
rect 5555 2645 5556 2675
rect 5524 2644 5556 2645
rect 5524 2595 5556 2596
rect 5524 2565 5525 2595
rect 5525 2565 5555 2595
rect 5555 2565 5556 2595
rect 5524 2564 5556 2565
rect 5524 2515 5556 2516
rect 5524 2485 5525 2515
rect 5525 2485 5555 2515
rect 5555 2485 5556 2515
rect 5524 2484 5556 2485
rect 5524 2435 5556 2436
rect 5524 2405 5525 2435
rect 5525 2405 5555 2435
rect 5555 2405 5556 2435
rect 5524 2404 5556 2405
rect 5524 2355 5556 2356
rect 5524 2325 5525 2355
rect 5525 2325 5555 2355
rect 5555 2325 5556 2355
rect 5524 2324 5556 2325
rect 5524 2275 5556 2276
rect 5524 2245 5525 2275
rect 5525 2245 5555 2275
rect 5555 2245 5556 2275
rect 5524 2244 5556 2245
rect 5524 2195 5556 2196
rect 5524 2165 5525 2195
rect 5525 2165 5555 2195
rect 5555 2165 5556 2195
rect 5524 2164 5556 2165
rect 5524 2115 5556 2116
rect 5524 2085 5525 2115
rect 5525 2085 5555 2115
rect 5555 2085 5556 2115
rect 5524 2084 5556 2085
rect 5524 2035 5556 2036
rect 5524 2005 5525 2035
rect 5525 2005 5555 2035
rect 5555 2005 5556 2035
rect 5524 2004 5556 2005
rect 5524 1635 5556 1636
rect 5524 1605 5525 1635
rect 5525 1605 5555 1635
rect 5555 1605 5556 1635
rect 5524 1604 5556 1605
rect 5524 1555 5556 1556
rect 5524 1525 5525 1555
rect 5525 1525 5555 1555
rect 5555 1525 5556 1555
rect 5524 1524 5556 1525
rect 5524 1475 5556 1476
rect 5524 1445 5525 1475
rect 5525 1445 5555 1475
rect 5555 1445 5556 1475
rect 5524 1444 5556 1445
rect 5524 1395 5556 1396
rect 5524 1365 5525 1395
rect 5525 1365 5555 1395
rect 5555 1365 5556 1395
rect 5524 1364 5556 1365
rect 5524 1315 5556 1316
rect 5524 1285 5525 1315
rect 5525 1285 5555 1315
rect 5555 1285 5556 1315
rect 5524 1284 5556 1285
rect 5524 1235 5556 1236
rect 5524 1205 5525 1235
rect 5525 1205 5555 1235
rect 5555 1205 5556 1235
rect 5524 1204 5556 1205
rect 5524 1155 5556 1156
rect 5524 1125 5525 1155
rect 5525 1125 5555 1155
rect 5555 1125 5556 1155
rect 5524 1124 5556 1125
rect 5524 1075 5556 1076
rect 5524 1045 5525 1075
rect 5525 1045 5555 1075
rect 5555 1045 5556 1075
rect 5524 1044 5556 1045
rect 5524 755 5556 756
rect 5524 725 5525 755
rect 5525 725 5555 755
rect 5555 725 5556 755
rect 5524 724 5556 725
rect 5524 675 5556 676
rect 5524 645 5525 675
rect 5525 645 5555 675
rect 5555 645 5556 675
rect 5524 644 5556 645
rect 5524 595 5556 596
rect 5524 565 5525 595
rect 5525 565 5555 595
rect 5555 565 5556 595
rect 5524 564 5556 565
rect 5524 195 5556 196
rect 5524 165 5525 195
rect 5525 165 5555 195
rect 5555 165 5556 195
rect 5524 164 5556 165
rect 5524 115 5556 116
rect 5524 85 5525 115
rect 5525 85 5555 115
rect 5555 85 5556 115
rect 5524 84 5556 85
rect 5524 35 5556 36
rect 5524 5 5525 35
rect 5525 5 5555 35
rect 5555 5 5556 35
rect 5524 4 5556 5
rect 5844 13204 5876 13396
rect 5684 12635 5716 12636
rect 5684 12605 5685 12635
rect 5685 12605 5715 12635
rect 5715 12605 5716 12635
rect 5684 12604 5716 12605
rect 5684 12555 5716 12556
rect 5684 12525 5685 12555
rect 5685 12525 5715 12555
rect 5715 12525 5716 12555
rect 5684 12524 5716 12525
rect 5684 12475 5716 12476
rect 5684 12445 5685 12475
rect 5685 12445 5715 12475
rect 5715 12445 5716 12475
rect 5684 12444 5716 12445
rect 5684 12395 5716 12396
rect 5684 12365 5685 12395
rect 5685 12365 5715 12395
rect 5715 12365 5716 12395
rect 5684 12364 5716 12365
rect 5684 12315 5716 12316
rect 5684 12285 5685 12315
rect 5685 12285 5715 12315
rect 5715 12285 5716 12315
rect 5684 12284 5716 12285
rect 5684 12235 5716 12236
rect 5684 12205 5685 12235
rect 5685 12205 5715 12235
rect 5715 12205 5716 12235
rect 5684 12204 5716 12205
rect 5684 12155 5716 12156
rect 5684 12125 5685 12155
rect 5685 12125 5715 12155
rect 5715 12125 5716 12155
rect 5684 12124 5716 12125
rect 5684 11835 5716 11836
rect 5684 11805 5685 11835
rect 5685 11805 5715 11835
rect 5715 11805 5716 11835
rect 5684 11804 5716 11805
rect 5684 11755 5716 11756
rect 5684 11725 5685 11755
rect 5685 11725 5715 11755
rect 5715 11725 5716 11755
rect 5684 11724 5716 11725
rect 5684 11675 5716 11676
rect 5684 11645 5685 11675
rect 5685 11645 5715 11675
rect 5715 11645 5716 11675
rect 5684 11644 5716 11645
rect 5684 11595 5716 11596
rect 5684 11565 5685 11595
rect 5685 11565 5715 11595
rect 5715 11565 5716 11595
rect 5684 11564 5716 11565
rect 5684 11515 5716 11516
rect 5684 11485 5685 11515
rect 5685 11485 5715 11515
rect 5715 11485 5716 11515
rect 5684 11484 5716 11485
rect 5684 11435 5716 11436
rect 5684 11405 5685 11435
rect 5685 11405 5715 11435
rect 5715 11405 5716 11435
rect 5684 11404 5716 11405
rect 5684 10875 5716 10876
rect 5684 10845 5685 10875
rect 5685 10845 5715 10875
rect 5715 10845 5716 10875
rect 5684 10844 5716 10845
rect 5684 10795 5716 10796
rect 5684 10765 5685 10795
rect 5685 10765 5715 10795
rect 5715 10765 5716 10795
rect 5684 10764 5716 10765
rect 5684 10715 5716 10716
rect 5684 10685 5685 10715
rect 5685 10685 5715 10715
rect 5715 10685 5716 10715
rect 5684 10684 5716 10685
rect 5684 10635 5716 10636
rect 5684 10605 5685 10635
rect 5685 10605 5715 10635
rect 5715 10605 5716 10635
rect 5684 10604 5716 10605
rect 5684 10555 5716 10556
rect 5684 10525 5685 10555
rect 5685 10525 5715 10555
rect 5715 10525 5716 10555
rect 5684 10524 5716 10525
rect 5684 10475 5716 10476
rect 5684 10445 5685 10475
rect 5685 10445 5715 10475
rect 5715 10445 5716 10475
rect 5684 10444 5716 10445
rect 5684 10395 5716 10396
rect 5684 10365 5685 10395
rect 5685 10365 5715 10395
rect 5715 10365 5716 10395
rect 5684 10364 5716 10365
rect 5684 10315 5716 10316
rect 5684 10285 5685 10315
rect 5685 10285 5715 10315
rect 5715 10285 5716 10315
rect 5684 10284 5716 10285
rect 5684 10235 5716 10236
rect 5684 10205 5685 10235
rect 5685 10205 5715 10235
rect 5715 10205 5716 10235
rect 5684 10204 5716 10205
rect 5684 10155 5716 10156
rect 5684 10125 5685 10155
rect 5685 10125 5715 10155
rect 5715 10125 5716 10155
rect 5684 10124 5716 10125
rect 5684 10075 5716 10076
rect 5684 10045 5685 10075
rect 5685 10045 5715 10075
rect 5715 10045 5716 10075
rect 5684 10044 5716 10045
rect 5684 9995 5716 9996
rect 5684 9965 5685 9995
rect 5685 9965 5715 9995
rect 5715 9965 5716 9995
rect 5684 9964 5716 9965
rect 5684 9915 5716 9916
rect 5684 9885 5685 9915
rect 5685 9885 5715 9915
rect 5715 9885 5716 9915
rect 5684 9884 5716 9885
rect 5684 9835 5716 9836
rect 5684 9805 5685 9835
rect 5685 9805 5715 9835
rect 5715 9805 5716 9835
rect 5684 9804 5716 9805
rect 5684 9755 5716 9756
rect 5684 9725 5685 9755
rect 5685 9725 5715 9755
rect 5715 9725 5716 9755
rect 5684 9724 5716 9725
rect 5684 9355 5716 9356
rect 5684 9325 5685 9355
rect 5685 9325 5715 9355
rect 5715 9325 5716 9355
rect 5684 9324 5716 9325
rect 5684 9275 5716 9276
rect 5684 9245 5685 9275
rect 5685 9245 5715 9275
rect 5715 9245 5716 9275
rect 5684 9244 5716 9245
rect 5684 9195 5716 9196
rect 5684 9165 5685 9195
rect 5685 9165 5715 9195
rect 5715 9165 5716 9195
rect 5684 9164 5716 9165
rect 5684 8875 5716 8876
rect 5684 8845 5685 8875
rect 5685 8845 5715 8875
rect 5715 8845 5716 8875
rect 5684 8844 5716 8845
rect 5684 8795 5716 8796
rect 5684 8765 5685 8795
rect 5685 8765 5715 8795
rect 5715 8765 5716 8795
rect 5684 8764 5716 8765
rect 5684 8715 5716 8716
rect 5684 8685 5685 8715
rect 5685 8685 5715 8715
rect 5715 8685 5716 8715
rect 5684 8684 5716 8685
rect 5684 8635 5716 8636
rect 5684 8605 5685 8635
rect 5685 8605 5715 8635
rect 5715 8605 5716 8635
rect 5684 8604 5716 8605
rect 5684 8555 5716 8556
rect 5684 8525 5685 8555
rect 5685 8525 5715 8555
rect 5715 8525 5716 8555
rect 5684 8524 5716 8525
rect 5684 7635 5716 7636
rect 5684 7605 5685 7635
rect 5685 7605 5715 7635
rect 5715 7605 5716 7635
rect 5684 7604 5716 7605
rect 5684 7555 5716 7556
rect 5684 7525 5685 7555
rect 5685 7525 5715 7555
rect 5715 7525 5716 7555
rect 5684 7524 5716 7525
rect 5684 7475 5716 7476
rect 5684 7445 5685 7475
rect 5685 7445 5715 7475
rect 5715 7445 5716 7475
rect 5684 7444 5716 7445
rect 5684 7395 5716 7396
rect 5684 7365 5685 7395
rect 5685 7365 5715 7395
rect 5715 7365 5716 7395
rect 5684 7364 5716 7365
rect 5684 7315 5716 7316
rect 5684 7285 5685 7315
rect 5685 7285 5715 7315
rect 5715 7285 5716 7315
rect 5684 7284 5716 7285
rect 5684 7235 5716 7236
rect 5684 7205 5685 7235
rect 5685 7205 5715 7235
rect 5715 7205 5716 7235
rect 5684 7204 5716 7205
rect 5684 7155 5716 7156
rect 5684 7125 5685 7155
rect 5685 7125 5715 7155
rect 5715 7125 5716 7155
rect 5684 7124 5716 7125
rect 5684 7075 5716 7076
rect 5684 7045 5685 7075
rect 5685 7045 5715 7075
rect 5715 7045 5716 7075
rect 5684 7044 5716 7045
rect 5684 6755 5716 6756
rect 5684 6725 5685 6755
rect 5685 6725 5715 6755
rect 5715 6725 5716 6755
rect 5684 6724 5716 6725
rect 5684 6675 5716 6676
rect 5684 6645 5685 6675
rect 5685 6645 5715 6675
rect 5715 6645 5716 6675
rect 5684 6644 5716 6645
rect 5684 6595 5716 6596
rect 5684 6565 5685 6595
rect 5685 6565 5715 6595
rect 5715 6565 5716 6595
rect 5684 6564 5716 6565
rect 5684 6515 5716 6516
rect 5684 6485 5685 6515
rect 5685 6485 5715 6515
rect 5715 6485 5716 6515
rect 5684 6484 5716 6485
rect 5684 6435 5716 6436
rect 5684 6405 5685 6435
rect 5685 6405 5715 6435
rect 5715 6405 5716 6435
rect 5684 6404 5716 6405
rect 5684 6355 5716 6356
rect 5684 6325 5685 6355
rect 5685 6325 5715 6355
rect 5715 6325 5716 6355
rect 5684 6324 5716 6325
rect 5684 5795 5716 5796
rect 5684 5765 5685 5795
rect 5685 5765 5715 5795
rect 5715 5765 5716 5795
rect 5684 5764 5716 5765
rect 5684 5715 5716 5716
rect 5684 5685 5685 5715
rect 5685 5685 5715 5715
rect 5715 5685 5716 5715
rect 5684 5684 5716 5685
rect 5684 5635 5716 5636
rect 5684 5605 5685 5635
rect 5685 5605 5715 5635
rect 5715 5605 5716 5635
rect 5684 5604 5716 5605
rect 5684 5555 5716 5556
rect 5684 5525 5685 5555
rect 5685 5525 5715 5555
rect 5715 5525 5716 5555
rect 5684 5524 5716 5525
rect 5684 5475 5716 5476
rect 5684 5445 5685 5475
rect 5685 5445 5715 5475
rect 5715 5445 5716 5475
rect 5684 5444 5716 5445
rect 5684 5395 5716 5396
rect 5684 5365 5685 5395
rect 5685 5365 5715 5395
rect 5715 5365 5716 5395
rect 5684 5364 5716 5365
rect 5684 5315 5716 5316
rect 5684 5285 5685 5315
rect 5685 5285 5715 5315
rect 5715 5285 5716 5315
rect 5684 5284 5716 5285
rect 5684 5235 5716 5236
rect 5684 5205 5685 5235
rect 5685 5205 5715 5235
rect 5715 5205 5716 5235
rect 5684 5204 5716 5205
rect 5684 5155 5716 5156
rect 5684 5125 5685 5155
rect 5685 5125 5715 5155
rect 5715 5125 5716 5155
rect 5684 5124 5716 5125
rect 5684 5075 5716 5076
rect 5684 5045 5685 5075
rect 5685 5045 5715 5075
rect 5715 5045 5716 5075
rect 5684 5044 5716 5045
rect 5684 4995 5716 4996
rect 5684 4965 5685 4995
rect 5685 4965 5715 4995
rect 5715 4965 5716 4995
rect 5684 4964 5716 4965
rect 5684 4435 5716 4436
rect 5684 4405 5685 4435
rect 5685 4405 5715 4435
rect 5715 4405 5716 4435
rect 5684 4404 5716 4405
rect 5684 4355 5716 4356
rect 5684 4325 5685 4355
rect 5685 4325 5715 4355
rect 5715 4325 5716 4355
rect 5684 4324 5716 4325
rect 5684 4275 5716 4276
rect 5684 4245 5685 4275
rect 5685 4245 5715 4275
rect 5715 4245 5716 4275
rect 5684 4244 5716 4245
rect 5684 4195 5716 4196
rect 5684 4165 5685 4195
rect 5685 4165 5715 4195
rect 5715 4165 5716 4195
rect 5684 4164 5716 4165
rect 5684 4115 5716 4116
rect 5684 4085 5685 4115
rect 5685 4085 5715 4115
rect 5715 4085 5716 4115
rect 5684 4084 5716 4085
rect 5684 4035 5716 4036
rect 5684 4005 5685 4035
rect 5685 4005 5715 4035
rect 5715 4005 5716 4035
rect 5684 4004 5716 4005
rect 5684 3955 5716 3956
rect 5684 3925 5685 3955
rect 5685 3925 5715 3955
rect 5715 3925 5716 3955
rect 5684 3924 5716 3925
rect 5684 3155 5716 3156
rect 5684 3125 5685 3155
rect 5685 3125 5715 3155
rect 5715 3125 5716 3155
rect 5684 3124 5716 3125
rect 5684 3075 5716 3076
rect 5684 3045 5685 3075
rect 5685 3045 5715 3075
rect 5715 3045 5716 3075
rect 5684 3044 5716 3045
rect 5684 2995 5716 2996
rect 5684 2965 5685 2995
rect 5685 2965 5715 2995
rect 5715 2965 5716 2995
rect 5684 2964 5716 2965
rect 5684 2915 5716 2916
rect 5684 2885 5685 2915
rect 5685 2885 5715 2915
rect 5715 2885 5716 2915
rect 5684 2884 5716 2885
rect 5684 2835 5716 2836
rect 5684 2805 5685 2835
rect 5685 2805 5715 2835
rect 5715 2805 5716 2835
rect 5684 2804 5716 2805
rect 5684 2755 5716 2756
rect 5684 2725 5685 2755
rect 5685 2725 5715 2755
rect 5715 2725 5716 2755
rect 5684 2724 5716 2725
rect 5684 2675 5716 2676
rect 5684 2645 5685 2675
rect 5685 2645 5715 2675
rect 5715 2645 5716 2675
rect 5684 2644 5716 2645
rect 5684 2595 5716 2596
rect 5684 2565 5685 2595
rect 5685 2565 5715 2595
rect 5715 2565 5716 2595
rect 5684 2564 5716 2565
rect 5684 2515 5716 2516
rect 5684 2485 5685 2515
rect 5685 2485 5715 2515
rect 5715 2485 5716 2515
rect 5684 2484 5716 2485
rect 5684 2435 5716 2436
rect 5684 2405 5685 2435
rect 5685 2405 5715 2435
rect 5715 2405 5716 2435
rect 5684 2404 5716 2405
rect 5684 2355 5716 2356
rect 5684 2325 5685 2355
rect 5685 2325 5715 2355
rect 5715 2325 5716 2355
rect 5684 2324 5716 2325
rect 5684 2275 5716 2276
rect 5684 2245 5685 2275
rect 5685 2245 5715 2275
rect 5715 2245 5716 2275
rect 5684 2244 5716 2245
rect 5684 2195 5716 2196
rect 5684 2165 5685 2195
rect 5685 2165 5715 2195
rect 5715 2165 5716 2195
rect 5684 2164 5716 2165
rect 5684 2115 5716 2116
rect 5684 2085 5685 2115
rect 5685 2085 5715 2115
rect 5715 2085 5716 2115
rect 5684 2084 5716 2085
rect 5684 2035 5716 2036
rect 5684 2005 5685 2035
rect 5685 2005 5715 2035
rect 5715 2005 5716 2035
rect 5684 2004 5716 2005
rect 5684 1635 5716 1636
rect 5684 1605 5685 1635
rect 5685 1605 5715 1635
rect 5715 1605 5716 1635
rect 5684 1604 5716 1605
rect 5684 1555 5716 1556
rect 5684 1525 5685 1555
rect 5685 1525 5715 1555
rect 5715 1525 5716 1555
rect 5684 1524 5716 1525
rect 5684 1475 5716 1476
rect 5684 1445 5685 1475
rect 5685 1445 5715 1475
rect 5715 1445 5716 1475
rect 5684 1444 5716 1445
rect 5684 1395 5716 1396
rect 5684 1365 5685 1395
rect 5685 1365 5715 1395
rect 5715 1365 5716 1395
rect 5684 1364 5716 1365
rect 5684 1315 5716 1316
rect 5684 1285 5685 1315
rect 5685 1285 5715 1315
rect 5715 1285 5716 1315
rect 5684 1284 5716 1285
rect 5684 1235 5716 1236
rect 5684 1205 5685 1235
rect 5685 1205 5715 1235
rect 5715 1205 5716 1235
rect 5684 1204 5716 1205
rect 5684 1155 5716 1156
rect 5684 1125 5685 1155
rect 5685 1125 5715 1155
rect 5715 1125 5716 1155
rect 5684 1124 5716 1125
rect 5684 1075 5716 1076
rect 5684 1045 5685 1075
rect 5685 1045 5715 1075
rect 5715 1045 5716 1075
rect 5684 1044 5716 1045
rect 5684 755 5716 756
rect 5684 725 5685 755
rect 5685 725 5715 755
rect 5715 725 5716 755
rect 5684 724 5716 725
rect 5684 675 5716 676
rect 5684 645 5685 675
rect 5685 645 5715 675
rect 5715 645 5716 675
rect 5684 644 5716 645
rect 5684 595 5716 596
rect 5684 565 5685 595
rect 5685 565 5715 595
rect 5715 565 5716 595
rect 5684 564 5716 565
rect 5684 195 5716 196
rect 5684 165 5685 195
rect 5685 165 5715 195
rect 5715 165 5716 195
rect 5684 164 5716 165
rect 5684 115 5716 116
rect 5684 85 5685 115
rect 5685 85 5715 115
rect 5715 85 5716 115
rect 5684 84 5716 85
rect 5684 35 5716 36
rect 5684 5 5685 35
rect 5685 5 5715 35
rect 5715 5 5716 35
rect 5684 4 5716 5
rect 6164 13204 6196 13396
rect 5844 12635 5876 12636
rect 5844 12605 5845 12635
rect 5845 12605 5875 12635
rect 5875 12605 5876 12635
rect 5844 12604 5876 12605
rect 5844 12555 5876 12556
rect 5844 12525 5845 12555
rect 5845 12525 5875 12555
rect 5875 12525 5876 12555
rect 5844 12524 5876 12525
rect 5844 12475 5876 12476
rect 5844 12445 5845 12475
rect 5845 12445 5875 12475
rect 5875 12445 5876 12475
rect 5844 12444 5876 12445
rect 5844 12395 5876 12396
rect 5844 12365 5845 12395
rect 5845 12365 5875 12395
rect 5875 12365 5876 12395
rect 5844 12364 5876 12365
rect 5844 12315 5876 12316
rect 5844 12285 5845 12315
rect 5845 12285 5875 12315
rect 5875 12285 5876 12315
rect 5844 12284 5876 12285
rect 5844 12235 5876 12236
rect 5844 12205 5845 12235
rect 5845 12205 5875 12235
rect 5875 12205 5876 12235
rect 5844 12204 5876 12205
rect 5844 12155 5876 12156
rect 5844 12125 5845 12155
rect 5845 12125 5875 12155
rect 5875 12125 5876 12155
rect 5844 12124 5876 12125
rect 5844 11835 5876 11836
rect 5844 11805 5845 11835
rect 5845 11805 5875 11835
rect 5875 11805 5876 11835
rect 5844 11804 5876 11805
rect 5844 11755 5876 11756
rect 5844 11725 5845 11755
rect 5845 11725 5875 11755
rect 5875 11725 5876 11755
rect 5844 11724 5876 11725
rect 5844 11675 5876 11676
rect 5844 11645 5845 11675
rect 5845 11645 5875 11675
rect 5875 11645 5876 11675
rect 5844 11644 5876 11645
rect 5844 11595 5876 11596
rect 5844 11565 5845 11595
rect 5845 11565 5875 11595
rect 5875 11565 5876 11595
rect 5844 11564 5876 11565
rect 5844 11515 5876 11516
rect 5844 11485 5845 11515
rect 5845 11485 5875 11515
rect 5875 11485 5876 11515
rect 5844 11484 5876 11485
rect 5844 11435 5876 11436
rect 5844 11405 5845 11435
rect 5845 11405 5875 11435
rect 5875 11405 5876 11435
rect 5844 11404 5876 11405
rect 5844 10875 5876 10876
rect 5844 10845 5845 10875
rect 5845 10845 5875 10875
rect 5875 10845 5876 10875
rect 5844 10844 5876 10845
rect 5844 10795 5876 10796
rect 5844 10765 5845 10795
rect 5845 10765 5875 10795
rect 5875 10765 5876 10795
rect 5844 10764 5876 10765
rect 5844 10715 5876 10716
rect 5844 10685 5845 10715
rect 5845 10685 5875 10715
rect 5875 10685 5876 10715
rect 5844 10684 5876 10685
rect 5844 10635 5876 10636
rect 5844 10605 5845 10635
rect 5845 10605 5875 10635
rect 5875 10605 5876 10635
rect 5844 10604 5876 10605
rect 5844 10555 5876 10556
rect 5844 10525 5845 10555
rect 5845 10525 5875 10555
rect 5875 10525 5876 10555
rect 5844 10524 5876 10525
rect 5844 10475 5876 10476
rect 5844 10445 5845 10475
rect 5845 10445 5875 10475
rect 5875 10445 5876 10475
rect 5844 10444 5876 10445
rect 5844 10395 5876 10396
rect 5844 10365 5845 10395
rect 5845 10365 5875 10395
rect 5875 10365 5876 10395
rect 5844 10364 5876 10365
rect 5844 10315 5876 10316
rect 5844 10285 5845 10315
rect 5845 10285 5875 10315
rect 5875 10285 5876 10315
rect 5844 10284 5876 10285
rect 5844 10235 5876 10236
rect 5844 10205 5845 10235
rect 5845 10205 5875 10235
rect 5875 10205 5876 10235
rect 5844 10204 5876 10205
rect 5844 10155 5876 10156
rect 5844 10125 5845 10155
rect 5845 10125 5875 10155
rect 5875 10125 5876 10155
rect 5844 10124 5876 10125
rect 5844 10075 5876 10076
rect 5844 10045 5845 10075
rect 5845 10045 5875 10075
rect 5875 10045 5876 10075
rect 5844 10044 5876 10045
rect 5844 9995 5876 9996
rect 5844 9965 5845 9995
rect 5845 9965 5875 9995
rect 5875 9965 5876 9995
rect 5844 9964 5876 9965
rect 5844 9915 5876 9916
rect 5844 9885 5845 9915
rect 5845 9885 5875 9915
rect 5875 9885 5876 9915
rect 5844 9884 5876 9885
rect 5844 9835 5876 9836
rect 5844 9805 5845 9835
rect 5845 9805 5875 9835
rect 5875 9805 5876 9835
rect 5844 9804 5876 9805
rect 5844 9755 5876 9756
rect 5844 9725 5845 9755
rect 5845 9725 5875 9755
rect 5875 9725 5876 9755
rect 5844 9724 5876 9725
rect 5844 9355 5876 9356
rect 5844 9325 5845 9355
rect 5845 9325 5875 9355
rect 5875 9325 5876 9355
rect 5844 9324 5876 9325
rect 5844 9275 5876 9276
rect 5844 9245 5845 9275
rect 5845 9245 5875 9275
rect 5875 9245 5876 9275
rect 5844 9244 5876 9245
rect 5844 9195 5876 9196
rect 5844 9165 5845 9195
rect 5845 9165 5875 9195
rect 5875 9165 5876 9195
rect 5844 9164 5876 9165
rect 5844 8875 5876 8876
rect 5844 8845 5845 8875
rect 5845 8845 5875 8875
rect 5875 8845 5876 8875
rect 5844 8844 5876 8845
rect 5844 8795 5876 8796
rect 5844 8765 5845 8795
rect 5845 8765 5875 8795
rect 5875 8765 5876 8795
rect 5844 8764 5876 8765
rect 5844 8715 5876 8716
rect 5844 8685 5845 8715
rect 5845 8685 5875 8715
rect 5875 8685 5876 8715
rect 5844 8684 5876 8685
rect 5844 8635 5876 8636
rect 5844 8605 5845 8635
rect 5845 8605 5875 8635
rect 5875 8605 5876 8635
rect 5844 8604 5876 8605
rect 5844 8555 5876 8556
rect 5844 8525 5845 8555
rect 5845 8525 5875 8555
rect 5875 8525 5876 8555
rect 5844 8524 5876 8525
rect 5844 7635 5876 7636
rect 5844 7605 5845 7635
rect 5845 7605 5875 7635
rect 5875 7605 5876 7635
rect 5844 7604 5876 7605
rect 5844 7555 5876 7556
rect 5844 7525 5845 7555
rect 5845 7525 5875 7555
rect 5875 7525 5876 7555
rect 5844 7524 5876 7525
rect 5844 7475 5876 7476
rect 5844 7445 5845 7475
rect 5845 7445 5875 7475
rect 5875 7445 5876 7475
rect 5844 7444 5876 7445
rect 5844 7395 5876 7396
rect 5844 7365 5845 7395
rect 5845 7365 5875 7395
rect 5875 7365 5876 7395
rect 5844 7364 5876 7365
rect 5844 7315 5876 7316
rect 5844 7285 5845 7315
rect 5845 7285 5875 7315
rect 5875 7285 5876 7315
rect 5844 7284 5876 7285
rect 5844 7235 5876 7236
rect 5844 7205 5845 7235
rect 5845 7205 5875 7235
rect 5875 7205 5876 7235
rect 5844 7204 5876 7205
rect 5844 7155 5876 7156
rect 5844 7125 5845 7155
rect 5845 7125 5875 7155
rect 5875 7125 5876 7155
rect 5844 7124 5876 7125
rect 5844 7075 5876 7076
rect 5844 7045 5845 7075
rect 5845 7045 5875 7075
rect 5875 7045 5876 7075
rect 5844 7044 5876 7045
rect 5844 6755 5876 6756
rect 5844 6725 5845 6755
rect 5845 6725 5875 6755
rect 5875 6725 5876 6755
rect 5844 6724 5876 6725
rect 5844 6675 5876 6676
rect 5844 6645 5845 6675
rect 5845 6645 5875 6675
rect 5875 6645 5876 6675
rect 5844 6644 5876 6645
rect 5844 6595 5876 6596
rect 5844 6565 5845 6595
rect 5845 6565 5875 6595
rect 5875 6565 5876 6595
rect 5844 6564 5876 6565
rect 5844 6515 5876 6516
rect 5844 6485 5845 6515
rect 5845 6485 5875 6515
rect 5875 6485 5876 6515
rect 5844 6484 5876 6485
rect 5844 6435 5876 6436
rect 5844 6405 5845 6435
rect 5845 6405 5875 6435
rect 5875 6405 5876 6435
rect 5844 6404 5876 6405
rect 5844 6355 5876 6356
rect 5844 6325 5845 6355
rect 5845 6325 5875 6355
rect 5875 6325 5876 6355
rect 5844 6324 5876 6325
rect 5844 5795 5876 5796
rect 5844 5765 5845 5795
rect 5845 5765 5875 5795
rect 5875 5765 5876 5795
rect 5844 5764 5876 5765
rect 5844 5715 5876 5716
rect 5844 5685 5845 5715
rect 5845 5685 5875 5715
rect 5875 5685 5876 5715
rect 5844 5684 5876 5685
rect 5844 5635 5876 5636
rect 5844 5605 5845 5635
rect 5845 5605 5875 5635
rect 5875 5605 5876 5635
rect 5844 5604 5876 5605
rect 5844 5555 5876 5556
rect 5844 5525 5845 5555
rect 5845 5525 5875 5555
rect 5875 5525 5876 5555
rect 5844 5524 5876 5525
rect 5844 5475 5876 5476
rect 5844 5445 5845 5475
rect 5845 5445 5875 5475
rect 5875 5445 5876 5475
rect 5844 5444 5876 5445
rect 5844 5395 5876 5396
rect 5844 5365 5845 5395
rect 5845 5365 5875 5395
rect 5875 5365 5876 5395
rect 5844 5364 5876 5365
rect 5844 5315 5876 5316
rect 5844 5285 5845 5315
rect 5845 5285 5875 5315
rect 5875 5285 5876 5315
rect 5844 5284 5876 5285
rect 5844 5235 5876 5236
rect 5844 5205 5845 5235
rect 5845 5205 5875 5235
rect 5875 5205 5876 5235
rect 5844 5204 5876 5205
rect 5844 5155 5876 5156
rect 5844 5125 5845 5155
rect 5845 5125 5875 5155
rect 5875 5125 5876 5155
rect 5844 5124 5876 5125
rect 5844 5075 5876 5076
rect 5844 5045 5845 5075
rect 5845 5045 5875 5075
rect 5875 5045 5876 5075
rect 5844 5044 5876 5045
rect 5844 4995 5876 4996
rect 5844 4965 5845 4995
rect 5845 4965 5875 4995
rect 5875 4965 5876 4995
rect 5844 4964 5876 4965
rect 5844 4435 5876 4436
rect 5844 4405 5845 4435
rect 5845 4405 5875 4435
rect 5875 4405 5876 4435
rect 5844 4404 5876 4405
rect 5844 4355 5876 4356
rect 5844 4325 5845 4355
rect 5845 4325 5875 4355
rect 5875 4325 5876 4355
rect 5844 4324 5876 4325
rect 5844 4275 5876 4276
rect 5844 4245 5845 4275
rect 5845 4245 5875 4275
rect 5875 4245 5876 4275
rect 5844 4244 5876 4245
rect 5844 4195 5876 4196
rect 5844 4165 5845 4195
rect 5845 4165 5875 4195
rect 5875 4165 5876 4195
rect 5844 4164 5876 4165
rect 5844 4115 5876 4116
rect 5844 4085 5845 4115
rect 5845 4085 5875 4115
rect 5875 4085 5876 4115
rect 5844 4084 5876 4085
rect 5844 4035 5876 4036
rect 5844 4005 5845 4035
rect 5845 4005 5875 4035
rect 5875 4005 5876 4035
rect 5844 4004 5876 4005
rect 5844 3955 5876 3956
rect 5844 3925 5845 3955
rect 5845 3925 5875 3955
rect 5875 3925 5876 3955
rect 5844 3924 5876 3925
rect 5844 3155 5876 3156
rect 5844 3125 5845 3155
rect 5845 3125 5875 3155
rect 5875 3125 5876 3155
rect 5844 3124 5876 3125
rect 5844 3075 5876 3076
rect 5844 3045 5845 3075
rect 5845 3045 5875 3075
rect 5875 3045 5876 3075
rect 5844 3044 5876 3045
rect 5844 2995 5876 2996
rect 5844 2965 5845 2995
rect 5845 2965 5875 2995
rect 5875 2965 5876 2995
rect 5844 2964 5876 2965
rect 5844 2915 5876 2916
rect 5844 2885 5845 2915
rect 5845 2885 5875 2915
rect 5875 2885 5876 2915
rect 5844 2884 5876 2885
rect 5844 2835 5876 2836
rect 5844 2805 5845 2835
rect 5845 2805 5875 2835
rect 5875 2805 5876 2835
rect 5844 2804 5876 2805
rect 5844 2755 5876 2756
rect 5844 2725 5845 2755
rect 5845 2725 5875 2755
rect 5875 2725 5876 2755
rect 5844 2724 5876 2725
rect 5844 2675 5876 2676
rect 5844 2645 5845 2675
rect 5845 2645 5875 2675
rect 5875 2645 5876 2675
rect 5844 2644 5876 2645
rect 5844 2595 5876 2596
rect 5844 2565 5845 2595
rect 5845 2565 5875 2595
rect 5875 2565 5876 2595
rect 5844 2564 5876 2565
rect 5844 2515 5876 2516
rect 5844 2485 5845 2515
rect 5845 2485 5875 2515
rect 5875 2485 5876 2515
rect 5844 2484 5876 2485
rect 5844 2435 5876 2436
rect 5844 2405 5845 2435
rect 5845 2405 5875 2435
rect 5875 2405 5876 2435
rect 5844 2404 5876 2405
rect 5844 2355 5876 2356
rect 5844 2325 5845 2355
rect 5845 2325 5875 2355
rect 5875 2325 5876 2355
rect 5844 2324 5876 2325
rect 5844 2275 5876 2276
rect 5844 2245 5845 2275
rect 5845 2245 5875 2275
rect 5875 2245 5876 2275
rect 5844 2244 5876 2245
rect 5844 2195 5876 2196
rect 5844 2165 5845 2195
rect 5845 2165 5875 2195
rect 5875 2165 5876 2195
rect 5844 2164 5876 2165
rect 5844 2115 5876 2116
rect 5844 2085 5845 2115
rect 5845 2085 5875 2115
rect 5875 2085 5876 2115
rect 5844 2084 5876 2085
rect 5844 2035 5876 2036
rect 5844 2005 5845 2035
rect 5845 2005 5875 2035
rect 5875 2005 5876 2035
rect 5844 2004 5876 2005
rect 5844 1635 5876 1636
rect 5844 1605 5845 1635
rect 5845 1605 5875 1635
rect 5875 1605 5876 1635
rect 5844 1604 5876 1605
rect 5844 1555 5876 1556
rect 5844 1525 5845 1555
rect 5845 1525 5875 1555
rect 5875 1525 5876 1555
rect 5844 1524 5876 1525
rect 5844 1475 5876 1476
rect 5844 1445 5845 1475
rect 5845 1445 5875 1475
rect 5875 1445 5876 1475
rect 5844 1444 5876 1445
rect 5844 1395 5876 1396
rect 5844 1365 5845 1395
rect 5845 1365 5875 1395
rect 5875 1365 5876 1395
rect 5844 1364 5876 1365
rect 5844 1315 5876 1316
rect 5844 1285 5845 1315
rect 5845 1285 5875 1315
rect 5875 1285 5876 1315
rect 5844 1284 5876 1285
rect 5844 1235 5876 1236
rect 5844 1205 5845 1235
rect 5845 1205 5875 1235
rect 5875 1205 5876 1235
rect 5844 1204 5876 1205
rect 5844 1155 5876 1156
rect 5844 1125 5845 1155
rect 5845 1125 5875 1155
rect 5875 1125 5876 1155
rect 5844 1124 5876 1125
rect 5844 1075 5876 1076
rect 5844 1045 5845 1075
rect 5845 1045 5875 1075
rect 5875 1045 5876 1075
rect 5844 1044 5876 1045
rect 5844 755 5876 756
rect 5844 725 5845 755
rect 5845 725 5875 755
rect 5875 725 5876 755
rect 5844 724 5876 725
rect 5844 675 5876 676
rect 5844 645 5845 675
rect 5845 645 5875 675
rect 5875 645 5876 675
rect 5844 644 5876 645
rect 5844 595 5876 596
rect 5844 565 5845 595
rect 5845 565 5875 595
rect 5875 565 5876 595
rect 5844 564 5876 565
rect 5844 195 5876 196
rect 5844 165 5845 195
rect 5845 165 5875 195
rect 5875 165 5876 195
rect 5844 164 5876 165
rect 5844 115 5876 116
rect 5844 85 5845 115
rect 5845 85 5875 115
rect 5875 85 5876 115
rect 5844 84 5876 85
rect 5844 35 5876 36
rect 5844 5 5845 35
rect 5845 5 5875 35
rect 5875 5 5876 35
rect 5844 4 5876 5
rect 5924 12724 5956 12916
rect 6084 12724 6116 12916
rect 5924 12635 5956 12636
rect 5924 12605 5925 12635
rect 5925 12605 5955 12635
rect 5955 12605 5956 12635
rect 5924 12604 5956 12605
rect 5924 12555 5956 12556
rect 5924 12525 5925 12555
rect 5925 12525 5955 12555
rect 5955 12525 5956 12555
rect 5924 12524 5956 12525
rect 5924 12475 5956 12476
rect 5924 12445 5925 12475
rect 5925 12445 5955 12475
rect 5955 12445 5956 12475
rect 5924 12444 5956 12445
rect 5924 12395 5956 12396
rect 5924 12365 5925 12395
rect 5925 12365 5955 12395
rect 5955 12365 5956 12395
rect 5924 12364 5956 12365
rect 5924 12315 5956 12316
rect 5924 12285 5925 12315
rect 5925 12285 5955 12315
rect 5955 12285 5956 12315
rect 5924 12284 5956 12285
rect 5924 12235 5956 12236
rect 5924 12205 5925 12235
rect 5925 12205 5955 12235
rect 5955 12205 5956 12235
rect 5924 12204 5956 12205
rect 5924 12155 5956 12156
rect 5924 12125 5925 12155
rect 5925 12125 5955 12155
rect 5955 12125 5956 12155
rect 5924 12124 5956 12125
rect 5924 11835 5956 11836
rect 5924 11805 5925 11835
rect 5925 11805 5955 11835
rect 5955 11805 5956 11835
rect 5924 11804 5956 11805
rect 5924 11755 5956 11756
rect 5924 11725 5925 11755
rect 5925 11725 5955 11755
rect 5955 11725 5956 11755
rect 5924 11724 5956 11725
rect 5924 11675 5956 11676
rect 5924 11645 5925 11675
rect 5925 11645 5955 11675
rect 5955 11645 5956 11675
rect 5924 11644 5956 11645
rect 5924 11595 5956 11596
rect 5924 11565 5925 11595
rect 5925 11565 5955 11595
rect 5955 11565 5956 11595
rect 5924 11564 5956 11565
rect 5924 11515 5956 11516
rect 5924 11485 5925 11515
rect 5925 11485 5955 11515
rect 5955 11485 5956 11515
rect 5924 11484 5956 11485
rect 5924 11435 5956 11436
rect 5924 11405 5925 11435
rect 5925 11405 5955 11435
rect 5955 11405 5956 11435
rect 5924 11404 5956 11405
rect 5924 10875 5956 10876
rect 5924 10845 5925 10875
rect 5925 10845 5955 10875
rect 5955 10845 5956 10875
rect 5924 10844 5956 10845
rect 5924 10795 5956 10796
rect 5924 10765 5925 10795
rect 5925 10765 5955 10795
rect 5955 10765 5956 10795
rect 5924 10764 5956 10765
rect 5924 10715 5956 10716
rect 5924 10685 5925 10715
rect 5925 10685 5955 10715
rect 5955 10685 5956 10715
rect 5924 10684 5956 10685
rect 5924 10635 5956 10636
rect 5924 10605 5925 10635
rect 5925 10605 5955 10635
rect 5955 10605 5956 10635
rect 5924 10604 5956 10605
rect 5924 10555 5956 10556
rect 5924 10525 5925 10555
rect 5925 10525 5955 10555
rect 5955 10525 5956 10555
rect 5924 10524 5956 10525
rect 5924 10475 5956 10476
rect 5924 10445 5925 10475
rect 5925 10445 5955 10475
rect 5955 10445 5956 10475
rect 5924 10444 5956 10445
rect 5924 10395 5956 10396
rect 5924 10365 5925 10395
rect 5925 10365 5955 10395
rect 5955 10365 5956 10395
rect 5924 10364 5956 10365
rect 5924 10315 5956 10316
rect 5924 10285 5925 10315
rect 5925 10285 5955 10315
rect 5955 10285 5956 10315
rect 5924 10284 5956 10285
rect 5924 10235 5956 10236
rect 5924 10205 5925 10235
rect 5925 10205 5955 10235
rect 5955 10205 5956 10235
rect 5924 10204 5956 10205
rect 5924 10155 5956 10156
rect 5924 10125 5925 10155
rect 5925 10125 5955 10155
rect 5955 10125 5956 10155
rect 5924 10124 5956 10125
rect 5924 10075 5956 10076
rect 5924 10045 5925 10075
rect 5925 10045 5955 10075
rect 5955 10045 5956 10075
rect 5924 10044 5956 10045
rect 5924 9995 5956 9996
rect 5924 9965 5925 9995
rect 5925 9965 5955 9995
rect 5955 9965 5956 9995
rect 5924 9964 5956 9965
rect 5924 9915 5956 9916
rect 5924 9885 5925 9915
rect 5925 9885 5955 9915
rect 5955 9885 5956 9915
rect 5924 9884 5956 9885
rect 5924 9835 5956 9836
rect 5924 9805 5925 9835
rect 5925 9805 5955 9835
rect 5955 9805 5956 9835
rect 5924 9804 5956 9805
rect 5924 9755 5956 9756
rect 5924 9725 5925 9755
rect 5925 9725 5955 9755
rect 5955 9725 5956 9755
rect 5924 9724 5956 9725
rect 5924 9355 5956 9356
rect 5924 9325 5925 9355
rect 5925 9325 5955 9355
rect 5955 9325 5956 9355
rect 5924 9324 5956 9325
rect 5924 9275 5956 9276
rect 5924 9245 5925 9275
rect 5925 9245 5955 9275
rect 5955 9245 5956 9275
rect 5924 9244 5956 9245
rect 5924 9195 5956 9196
rect 5924 9165 5925 9195
rect 5925 9165 5955 9195
rect 5955 9165 5956 9195
rect 5924 9164 5956 9165
rect 5924 8875 5956 8876
rect 5924 8845 5925 8875
rect 5925 8845 5955 8875
rect 5955 8845 5956 8875
rect 5924 8844 5956 8845
rect 5924 8795 5956 8796
rect 5924 8765 5925 8795
rect 5925 8765 5955 8795
rect 5955 8765 5956 8795
rect 5924 8764 5956 8765
rect 5924 8715 5956 8716
rect 5924 8685 5925 8715
rect 5925 8685 5955 8715
rect 5955 8685 5956 8715
rect 5924 8684 5956 8685
rect 5924 8635 5956 8636
rect 5924 8605 5925 8635
rect 5925 8605 5955 8635
rect 5955 8605 5956 8635
rect 5924 8604 5956 8605
rect 5924 8555 5956 8556
rect 5924 8525 5925 8555
rect 5925 8525 5955 8555
rect 5955 8525 5956 8555
rect 5924 8524 5956 8525
rect 5924 7635 5956 7636
rect 5924 7605 5925 7635
rect 5925 7605 5955 7635
rect 5955 7605 5956 7635
rect 5924 7604 5956 7605
rect 5924 7555 5956 7556
rect 5924 7525 5925 7555
rect 5925 7525 5955 7555
rect 5955 7525 5956 7555
rect 5924 7524 5956 7525
rect 5924 7475 5956 7476
rect 5924 7445 5925 7475
rect 5925 7445 5955 7475
rect 5955 7445 5956 7475
rect 5924 7444 5956 7445
rect 5924 7395 5956 7396
rect 5924 7365 5925 7395
rect 5925 7365 5955 7395
rect 5955 7365 5956 7395
rect 5924 7364 5956 7365
rect 5924 7315 5956 7316
rect 5924 7285 5925 7315
rect 5925 7285 5955 7315
rect 5955 7285 5956 7315
rect 5924 7284 5956 7285
rect 5924 7235 5956 7236
rect 5924 7205 5925 7235
rect 5925 7205 5955 7235
rect 5955 7205 5956 7235
rect 5924 7204 5956 7205
rect 5924 7155 5956 7156
rect 5924 7125 5925 7155
rect 5925 7125 5955 7155
rect 5955 7125 5956 7155
rect 5924 7124 5956 7125
rect 5924 7075 5956 7076
rect 5924 7045 5925 7075
rect 5925 7045 5955 7075
rect 5955 7045 5956 7075
rect 5924 7044 5956 7045
rect 5924 6755 5956 6756
rect 5924 6725 5925 6755
rect 5925 6725 5955 6755
rect 5955 6725 5956 6755
rect 5924 6724 5956 6725
rect 5924 6675 5956 6676
rect 5924 6645 5925 6675
rect 5925 6645 5955 6675
rect 5955 6645 5956 6675
rect 5924 6644 5956 6645
rect 5924 6595 5956 6596
rect 5924 6565 5925 6595
rect 5925 6565 5955 6595
rect 5955 6565 5956 6595
rect 5924 6564 5956 6565
rect 5924 6515 5956 6516
rect 5924 6485 5925 6515
rect 5925 6485 5955 6515
rect 5955 6485 5956 6515
rect 5924 6484 5956 6485
rect 5924 6435 5956 6436
rect 5924 6405 5925 6435
rect 5925 6405 5955 6435
rect 5955 6405 5956 6435
rect 5924 6404 5956 6405
rect 5924 6355 5956 6356
rect 5924 6325 5925 6355
rect 5925 6325 5955 6355
rect 5955 6325 5956 6355
rect 5924 6324 5956 6325
rect 5924 5795 5956 5796
rect 5924 5765 5925 5795
rect 5925 5765 5955 5795
rect 5955 5765 5956 5795
rect 5924 5764 5956 5765
rect 5924 5715 5956 5716
rect 5924 5685 5925 5715
rect 5925 5685 5955 5715
rect 5955 5685 5956 5715
rect 5924 5684 5956 5685
rect 5924 5635 5956 5636
rect 5924 5605 5925 5635
rect 5925 5605 5955 5635
rect 5955 5605 5956 5635
rect 5924 5604 5956 5605
rect 5924 5555 5956 5556
rect 5924 5525 5925 5555
rect 5925 5525 5955 5555
rect 5955 5525 5956 5555
rect 5924 5524 5956 5525
rect 5924 5475 5956 5476
rect 5924 5445 5925 5475
rect 5925 5445 5955 5475
rect 5955 5445 5956 5475
rect 5924 5444 5956 5445
rect 5924 5395 5956 5396
rect 5924 5365 5925 5395
rect 5925 5365 5955 5395
rect 5955 5365 5956 5395
rect 5924 5364 5956 5365
rect 5924 5315 5956 5316
rect 5924 5285 5925 5315
rect 5925 5285 5955 5315
rect 5955 5285 5956 5315
rect 5924 5284 5956 5285
rect 5924 5235 5956 5236
rect 5924 5205 5925 5235
rect 5925 5205 5955 5235
rect 5955 5205 5956 5235
rect 5924 5204 5956 5205
rect 5924 5155 5956 5156
rect 5924 5125 5925 5155
rect 5925 5125 5955 5155
rect 5955 5125 5956 5155
rect 5924 5124 5956 5125
rect 5924 5075 5956 5076
rect 5924 5045 5925 5075
rect 5925 5045 5955 5075
rect 5955 5045 5956 5075
rect 5924 5044 5956 5045
rect 5924 4995 5956 4996
rect 5924 4965 5925 4995
rect 5925 4965 5955 4995
rect 5955 4965 5956 4995
rect 5924 4964 5956 4965
rect 5924 4435 5956 4436
rect 5924 4405 5925 4435
rect 5925 4405 5955 4435
rect 5955 4405 5956 4435
rect 5924 4404 5956 4405
rect 5924 4355 5956 4356
rect 5924 4325 5925 4355
rect 5925 4325 5955 4355
rect 5955 4325 5956 4355
rect 5924 4324 5956 4325
rect 5924 4275 5956 4276
rect 5924 4245 5925 4275
rect 5925 4245 5955 4275
rect 5955 4245 5956 4275
rect 5924 4244 5956 4245
rect 5924 4195 5956 4196
rect 5924 4165 5925 4195
rect 5925 4165 5955 4195
rect 5955 4165 5956 4195
rect 5924 4164 5956 4165
rect 5924 4115 5956 4116
rect 5924 4085 5925 4115
rect 5925 4085 5955 4115
rect 5955 4085 5956 4115
rect 5924 4084 5956 4085
rect 5924 4035 5956 4036
rect 5924 4005 5925 4035
rect 5925 4005 5955 4035
rect 5955 4005 5956 4035
rect 5924 4004 5956 4005
rect 5924 3955 5956 3956
rect 5924 3925 5925 3955
rect 5925 3925 5955 3955
rect 5955 3925 5956 3955
rect 5924 3924 5956 3925
rect 5924 3155 5956 3156
rect 5924 3125 5925 3155
rect 5925 3125 5955 3155
rect 5955 3125 5956 3155
rect 5924 3124 5956 3125
rect 5924 3075 5956 3076
rect 5924 3045 5925 3075
rect 5925 3045 5955 3075
rect 5955 3045 5956 3075
rect 5924 3044 5956 3045
rect 5924 2995 5956 2996
rect 5924 2965 5925 2995
rect 5925 2965 5955 2995
rect 5955 2965 5956 2995
rect 5924 2964 5956 2965
rect 5924 2915 5956 2916
rect 5924 2885 5925 2915
rect 5925 2885 5955 2915
rect 5955 2885 5956 2915
rect 5924 2884 5956 2885
rect 5924 2835 5956 2836
rect 5924 2805 5925 2835
rect 5925 2805 5955 2835
rect 5955 2805 5956 2835
rect 5924 2804 5956 2805
rect 5924 2755 5956 2756
rect 5924 2725 5925 2755
rect 5925 2725 5955 2755
rect 5955 2725 5956 2755
rect 5924 2724 5956 2725
rect 5924 2675 5956 2676
rect 5924 2645 5925 2675
rect 5925 2645 5955 2675
rect 5955 2645 5956 2675
rect 5924 2644 5956 2645
rect 5924 2595 5956 2596
rect 5924 2565 5925 2595
rect 5925 2565 5955 2595
rect 5955 2565 5956 2595
rect 5924 2564 5956 2565
rect 5924 2515 5956 2516
rect 5924 2485 5925 2515
rect 5925 2485 5955 2515
rect 5955 2485 5956 2515
rect 5924 2484 5956 2485
rect 5924 2435 5956 2436
rect 5924 2405 5925 2435
rect 5925 2405 5955 2435
rect 5955 2405 5956 2435
rect 5924 2404 5956 2405
rect 5924 2355 5956 2356
rect 5924 2325 5925 2355
rect 5925 2325 5955 2355
rect 5955 2325 5956 2355
rect 5924 2324 5956 2325
rect 5924 2275 5956 2276
rect 5924 2245 5925 2275
rect 5925 2245 5955 2275
rect 5955 2245 5956 2275
rect 5924 2244 5956 2245
rect 5924 2195 5956 2196
rect 5924 2165 5925 2195
rect 5925 2165 5955 2195
rect 5955 2165 5956 2195
rect 5924 2164 5956 2165
rect 5924 2115 5956 2116
rect 5924 2085 5925 2115
rect 5925 2085 5955 2115
rect 5955 2085 5956 2115
rect 5924 2084 5956 2085
rect 5924 2035 5956 2036
rect 5924 2005 5925 2035
rect 5925 2005 5955 2035
rect 5955 2005 5956 2035
rect 5924 2004 5956 2005
rect 5924 1635 5956 1636
rect 5924 1605 5925 1635
rect 5925 1605 5955 1635
rect 5955 1605 5956 1635
rect 5924 1604 5956 1605
rect 5924 1555 5956 1556
rect 5924 1525 5925 1555
rect 5925 1525 5955 1555
rect 5955 1525 5956 1555
rect 5924 1524 5956 1525
rect 5924 1475 5956 1476
rect 5924 1445 5925 1475
rect 5925 1445 5955 1475
rect 5955 1445 5956 1475
rect 5924 1444 5956 1445
rect 5924 1395 5956 1396
rect 5924 1365 5925 1395
rect 5925 1365 5955 1395
rect 5955 1365 5956 1395
rect 5924 1364 5956 1365
rect 5924 1315 5956 1316
rect 5924 1285 5925 1315
rect 5925 1285 5955 1315
rect 5955 1285 5956 1315
rect 5924 1284 5956 1285
rect 5924 1235 5956 1236
rect 5924 1205 5925 1235
rect 5925 1205 5955 1235
rect 5955 1205 5956 1235
rect 5924 1204 5956 1205
rect 5924 1155 5956 1156
rect 5924 1125 5925 1155
rect 5925 1125 5955 1155
rect 5955 1125 5956 1155
rect 5924 1124 5956 1125
rect 5924 1075 5956 1076
rect 5924 1045 5925 1075
rect 5925 1045 5955 1075
rect 5955 1045 5956 1075
rect 5924 1044 5956 1045
rect 5924 755 5956 756
rect 5924 725 5925 755
rect 5925 725 5955 755
rect 5955 725 5956 755
rect 5924 724 5956 725
rect 5924 675 5956 676
rect 5924 645 5925 675
rect 5925 645 5955 675
rect 5955 645 5956 675
rect 5924 644 5956 645
rect 5924 595 5956 596
rect 5924 565 5925 595
rect 5925 565 5955 595
rect 5955 565 5956 595
rect 5924 564 5956 565
rect 5924 195 5956 196
rect 5924 165 5925 195
rect 5925 165 5955 195
rect 5955 165 5956 195
rect 5924 164 5956 165
rect 5924 115 5956 116
rect 5924 85 5925 115
rect 5925 85 5955 115
rect 5955 85 5956 115
rect 5924 84 5956 85
rect 5924 35 5956 36
rect 5924 5 5925 35
rect 5925 5 5955 35
rect 5955 5 5956 35
rect 5924 4 5956 5
rect 6084 12635 6116 12636
rect 6084 12605 6085 12635
rect 6085 12605 6115 12635
rect 6115 12605 6116 12635
rect 6084 12604 6116 12605
rect 6084 12555 6116 12556
rect 6084 12525 6085 12555
rect 6085 12525 6115 12555
rect 6115 12525 6116 12555
rect 6084 12524 6116 12525
rect 6084 12475 6116 12476
rect 6084 12445 6085 12475
rect 6085 12445 6115 12475
rect 6115 12445 6116 12475
rect 6084 12444 6116 12445
rect 6084 12395 6116 12396
rect 6084 12365 6085 12395
rect 6085 12365 6115 12395
rect 6115 12365 6116 12395
rect 6084 12364 6116 12365
rect 6084 12315 6116 12316
rect 6084 12285 6085 12315
rect 6085 12285 6115 12315
rect 6115 12285 6116 12315
rect 6084 12284 6116 12285
rect 6084 12235 6116 12236
rect 6084 12205 6085 12235
rect 6085 12205 6115 12235
rect 6115 12205 6116 12235
rect 6084 12204 6116 12205
rect 6084 12155 6116 12156
rect 6084 12125 6085 12155
rect 6085 12125 6115 12155
rect 6115 12125 6116 12155
rect 6084 12124 6116 12125
rect 6084 11835 6116 11836
rect 6084 11805 6085 11835
rect 6085 11805 6115 11835
rect 6115 11805 6116 11835
rect 6084 11804 6116 11805
rect 6084 11755 6116 11756
rect 6084 11725 6085 11755
rect 6085 11725 6115 11755
rect 6115 11725 6116 11755
rect 6084 11724 6116 11725
rect 6084 11675 6116 11676
rect 6084 11645 6085 11675
rect 6085 11645 6115 11675
rect 6115 11645 6116 11675
rect 6084 11644 6116 11645
rect 6084 11595 6116 11596
rect 6084 11565 6085 11595
rect 6085 11565 6115 11595
rect 6115 11565 6116 11595
rect 6084 11564 6116 11565
rect 6084 11515 6116 11516
rect 6084 11485 6085 11515
rect 6085 11485 6115 11515
rect 6115 11485 6116 11515
rect 6084 11484 6116 11485
rect 6084 11435 6116 11436
rect 6084 11405 6085 11435
rect 6085 11405 6115 11435
rect 6115 11405 6116 11435
rect 6084 11404 6116 11405
rect 6084 10875 6116 10876
rect 6084 10845 6085 10875
rect 6085 10845 6115 10875
rect 6115 10845 6116 10875
rect 6084 10844 6116 10845
rect 6084 10795 6116 10796
rect 6084 10765 6085 10795
rect 6085 10765 6115 10795
rect 6115 10765 6116 10795
rect 6084 10764 6116 10765
rect 6084 10715 6116 10716
rect 6084 10685 6085 10715
rect 6085 10685 6115 10715
rect 6115 10685 6116 10715
rect 6084 10684 6116 10685
rect 6084 10635 6116 10636
rect 6084 10605 6085 10635
rect 6085 10605 6115 10635
rect 6115 10605 6116 10635
rect 6084 10604 6116 10605
rect 6084 10555 6116 10556
rect 6084 10525 6085 10555
rect 6085 10525 6115 10555
rect 6115 10525 6116 10555
rect 6084 10524 6116 10525
rect 6084 10475 6116 10476
rect 6084 10445 6085 10475
rect 6085 10445 6115 10475
rect 6115 10445 6116 10475
rect 6084 10444 6116 10445
rect 6084 10395 6116 10396
rect 6084 10365 6085 10395
rect 6085 10365 6115 10395
rect 6115 10365 6116 10395
rect 6084 10364 6116 10365
rect 6084 10315 6116 10316
rect 6084 10285 6085 10315
rect 6085 10285 6115 10315
rect 6115 10285 6116 10315
rect 6084 10284 6116 10285
rect 6084 10235 6116 10236
rect 6084 10205 6085 10235
rect 6085 10205 6115 10235
rect 6115 10205 6116 10235
rect 6084 10204 6116 10205
rect 6084 10155 6116 10156
rect 6084 10125 6085 10155
rect 6085 10125 6115 10155
rect 6115 10125 6116 10155
rect 6084 10124 6116 10125
rect 6084 10075 6116 10076
rect 6084 10045 6085 10075
rect 6085 10045 6115 10075
rect 6115 10045 6116 10075
rect 6084 10044 6116 10045
rect 6084 9995 6116 9996
rect 6084 9965 6085 9995
rect 6085 9965 6115 9995
rect 6115 9965 6116 9995
rect 6084 9964 6116 9965
rect 6084 9915 6116 9916
rect 6084 9885 6085 9915
rect 6085 9885 6115 9915
rect 6115 9885 6116 9915
rect 6084 9884 6116 9885
rect 6084 9835 6116 9836
rect 6084 9805 6085 9835
rect 6085 9805 6115 9835
rect 6115 9805 6116 9835
rect 6084 9804 6116 9805
rect 6084 9755 6116 9756
rect 6084 9725 6085 9755
rect 6085 9725 6115 9755
rect 6115 9725 6116 9755
rect 6084 9724 6116 9725
rect 6084 9355 6116 9356
rect 6084 9325 6085 9355
rect 6085 9325 6115 9355
rect 6115 9325 6116 9355
rect 6084 9324 6116 9325
rect 6084 9275 6116 9276
rect 6084 9245 6085 9275
rect 6085 9245 6115 9275
rect 6115 9245 6116 9275
rect 6084 9244 6116 9245
rect 6084 9195 6116 9196
rect 6084 9165 6085 9195
rect 6085 9165 6115 9195
rect 6115 9165 6116 9195
rect 6084 9164 6116 9165
rect 6084 8875 6116 8876
rect 6084 8845 6085 8875
rect 6085 8845 6115 8875
rect 6115 8845 6116 8875
rect 6084 8844 6116 8845
rect 6084 8795 6116 8796
rect 6084 8765 6085 8795
rect 6085 8765 6115 8795
rect 6115 8765 6116 8795
rect 6084 8764 6116 8765
rect 6084 8715 6116 8716
rect 6084 8685 6085 8715
rect 6085 8685 6115 8715
rect 6115 8685 6116 8715
rect 6084 8684 6116 8685
rect 6084 8635 6116 8636
rect 6084 8605 6085 8635
rect 6085 8605 6115 8635
rect 6115 8605 6116 8635
rect 6084 8604 6116 8605
rect 6084 8555 6116 8556
rect 6084 8525 6085 8555
rect 6085 8525 6115 8555
rect 6115 8525 6116 8555
rect 6084 8524 6116 8525
rect 6084 7635 6116 7636
rect 6084 7605 6085 7635
rect 6085 7605 6115 7635
rect 6115 7605 6116 7635
rect 6084 7604 6116 7605
rect 6084 7555 6116 7556
rect 6084 7525 6085 7555
rect 6085 7525 6115 7555
rect 6115 7525 6116 7555
rect 6084 7524 6116 7525
rect 6084 7475 6116 7476
rect 6084 7445 6085 7475
rect 6085 7445 6115 7475
rect 6115 7445 6116 7475
rect 6084 7444 6116 7445
rect 6084 7395 6116 7396
rect 6084 7365 6085 7395
rect 6085 7365 6115 7395
rect 6115 7365 6116 7395
rect 6084 7364 6116 7365
rect 6084 7315 6116 7316
rect 6084 7285 6085 7315
rect 6085 7285 6115 7315
rect 6115 7285 6116 7315
rect 6084 7284 6116 7285
rect 6084 7235 6116 7236
rect 6084 7205 6085 7235
rect 6085 7205 6115 7235
rect 6115 7205 6116 7235
rect 6084 7204 6116 7205
rect 6084 7155 6116 7156
rect 6084 7125 6085 7155
rect 6085 7125 6115 7155
rect 6115 7125 6116 7155
rect 6084 7124 6116 7125
rect 6084 7075 6116 7076
rect 6084 7045 6085 7075
rect 6085 7045 6115 7075
rect 6115 7045 6116 7075
rect 6084 7044 6116 7045
rect 6084 6755 6116 6756
rect 6084 6725 6085 6755
rect 6085 6725 6115 6755
rect 6115 6725 6116 6755
rect 6084 6724 6116 6725
rect 6084 6675 6116 6676
rect 6084 6645 6085 6675
rect 6085 6645 6115 6675
rect 6115 6645 6116 6675
rect 6084 6644 6116 6645
rect 6084 6595 6116 6596
rect 6084 6565 6085 6595
rect 6085 6565 6115 6595
rect 6115 6565 6116 6595
rect 6084 6564 6116 6565
rect 6084 6515 6116 6516
rect 6084 6485 6085 6515
rect 6085 6485 6115 6515
rect 6115 6485 6116 6515
rect 6084 6484 6116 6485
rect 6084 6435 6116 6436
rect 6084 6405 6085 6435
rect 6085 6405 6115 6435
rect 6115 6405 6116 6435
rect 6084 6404 6116 6405
rect 6084 6355 6116 6356
rect 6084 6325 6085 6355
rect 6085 6325 6115 6355
rect 6115 6325 6116 6355
rect 6084 6324 6116 6325
rect 6084 5795 6116 5796
rect 6084 5765 6085 5795
rect 6085 5765 6115 5795
rect 6115 5765 6116 5795
rect 6084 5764 6116 5765
rect 6084 5715 6116 5716
rect 6084 5685 6085 5715
rect 6085 5685 6115 5715
rect 6115 5685 6116 5715
rect 6084 5684 6116 5685
rect 6084 5635 6116 5636
rect 6084 5605 6085 5635
rect 6085 5605 6115 5635
rect 6115 5605 6116 5635
rect 6084 5604 6116 5605
rect 6084 5555 6116 5556
rect 6084 5525 6085 5555
rect 6085 5525 6115 5555
rect 6115 5525 6116 5555
rect 6084 5524 6116 5525
rect 6084 5475 6116 5476
rect 6084 5445 6085 5475
rect 6085 5445 6115 5475
rect 6115 5445 6116 5475
rect 6084 5444 6116 5445
rect 6084 5395 6116 5396
rect 6084 5365 6085 5395
rect 6085 5365 6115 5395
rect 6115 5365 6116 5395
rect 6084 5364 6116 5365
rect 6084 5315 6116 5316
rect 6084 5285 6085 5315
rect 6085 5285 6115 5315
rect 6115 5285 6116 5315
rect 6084 5284 6116 5285
rect 6084 5235 6116 5236
rect 6084 5205 6085 5235
rect 6085 5205 6115 5235
rect 6115 5205 6116 5235
rect 6084 5204 6116 5205
rect 6084 5155 6116 5156
rect 6084 5125 6085 5155
rect 6085 5125 6115 5155
rect 6115 5125 6116 5155
rect 6084 5124 6116 5125
rect 6084 5075 6116 5076
rect 6084 5045 6085 5075
rect 6085 5045 6115 5075
rect 6115 5045 6116 5075
rect 6084 5044 6116 5045
rect 6084 4995 6116 4996
rect 6084 4965 6085 4995
rect 6085 4965 6115 4995
rect 6115 4965 6116 4995
rect 6084 4964 6116 4965
rect 6084 4435 6116 4436
rect 6084 4405 6085 4435
rect 6085 4405 6115 4435
rect 6115 4405 6116 4435
rect 6084 4404 6116 4405
rect 6084 4355 6116 4356
rect 6084 4325 6085 4355
rect 6085 4325 6115 4355
rect 6115 4325 6116 4355
rect 6084 4324 6116 4325
rect 6084 4275 6116 4276
rect 6084 4245 6085 4275
rect 6085 4245 6115 4275
rect 6115 4245 6116 4275
rect 6084 4244 6116 4245
rect 6084 4195 6116 4196
rect 6084 4165 6085 4195
rect 6085 4165 6115 4195
rect 6115 4165 6116 4195
rect 6084 4164 6116 4165
rect 6084 4115 6116 4116
rect 6084 4085 6085 4115
rect 6085 4085 6115 4115
rect 6115 4085 6116 4115
rect 6084 4084 6116 4085
rect 6084 4035 6116 4036
rect 6084 4005 6085 4035
rect 6085 4005 6115 4035
rect 6115 4005 6116 4035
rect 6084 4004 6116 4005
rect 6084 3955 6116 3956
rect 6084 3925 6085 3955
rect 6085 3925 6115 3955
rect 6115 3925 6116 3955
rect 6084 3924 6116 3925
rect 6084 3155 6116 3156
rect 6084 3125 6085 3155
rect 6085 3125 6115 3155
rect 6115 3125 6116 3155
rect 6084 3124 6116 3125
rect 6084 3075 6116 3076
rect 6084 3045 6085 3075
rect 6085 3045 6115 3075
rect 6115 3045 6116 3075
rect 6084 3044 6116 3045
rect 6084 2995 6116 2996
rect 6084 2965 6085 2995
rect 6085 2965 6115 2995
rect 6115 2965 6116 2995
rect 6084 2964 6116 2965
rect 6084 2915 6116 2916
rect 6084 2885 6085 2915
rect 6085 2885 6115 2915
rect 6115 2885 6116 2915
rect 6084 2884 6116 2885
rect 6084 2835 6116 2836
rect 6084 2805 6085 2835
rect 6085 2805 6115 2835
rect 6115 2805 6116 2835
rect 6084 2804 6116 2805
rect 6084 2755 6116 2756
rect 6084 2725 6085 2755
rect 6085 2725 6115 2755
rect 6115 2725 6116 2755
rect 6084 2724 6116 2725
rect 6084 2675 6116 2676
rect 6084 2645 6085 2675
rect 6085 2645 6115 2675
rect 6115 2645 6116 2675
rect 6084 2644 6116 2645
rect 6084 2595 6116 2596
rect 6084 2565 6085 2595
rect 6085 2565 6115 2595
rect 6115 2565 6116 2595
rect 6084 2564 6116 2565
rect 6084 2515 6116 2516
rect 6084 2485 6085 2515
rect 6085 2485 6115 2515
rect 6115 2485 6116 2515
rect 6084 2484 6116 2485
rect 6084 2435 6116 2436
rect 6084 2405 6085 2435
rect 6085 2405 6115 2435
rect 6115 2405 6116 2435
rect 6084 2404 6116 2405
rect 6084 2355 6116 2356
rect 6084 2325 6085 2355
rect 6085 2325 6115 2355
rect 6115 2325 6116 2355
rect 6084 2324 6116 2325
rect 6084 2275 6116 2276
rect 6084 2245 6085 2275
rect 6085 2245 6115 2275
rect 6115 2245 6116 2275
rect 6084 2244 6116 2245
rect 6084 2195 6116 2196
rect 6084 2165 6085 2195
rect 6085 2165 6115 2195
rect 6115 2165 6116 2195
rect 6084 2164 6116 2165
rect 6084 2115 6116 2116
rect 6084 2085 6085 2115
rect 6085 2085 6115 2115
rect 6115 2085 6116 2115
rect 6084 2084 6116 2085
rect 6084 2035 6116 2036
rect 6084 2005 6085 2035
rect 6085 2005 6115 2035
rect 6115 2005 6116 2035
rect 6084 2004 6116 2005
rect 6084 1635 6116 1636
rect 6084 1605 6085 1635
rect 6085 1605 6115 1635
rect 6115 1605 6116 1635
rect 6084 1604 6116 1605
rect 6084 1555 6116 1556
rect 6084 1525 6085 1555
rect 6085 1525 6115 1555
rect 6115 1525 6116 1555
rect 6084 1524 6116 1525
rect 6084 1475 6116 1476
rect 6084 1445 6085 1475
rect 6085 1445 6115 1475
rect 6115 1445 6116 1475
rect 6084 1444 6116 1445
rect 6084 1395 6116 1396
rect 6084 1365 6085 1395
rect 6085 1365 6115 1395
rect 6115 1365 6116 1395
rect 6084 1364 6116 1365
rect 6084 1315 6116 1316
rect 6084 1285 6085 1315
rect 6085 1285 6115 1315
rect 6115 1285 6116 1315
rect 6084 1284 6116 1285
rect 6084 1235 6116 1236
rect 6084 1205 6085 1235
rect 6085 1205 6115 1235
rect 6115 1205 6116 1235
rect 6084 1204 6116 1205
rect 6084 1155 6116 1156
rect 6084 1125 6085 1155
rect 6085 1125 6115 1155
rect 6115 1125 6116 1155
rect 6084 1124 6116 1125
rect 6084 1075 6116 1076
rect 6084 1045 6085 1075
rect 6085 1045 6115 1075
rect 6115 1045 6116 1075
rect 6084 1044 6116 1045
rect 6084 755 6116 756
rect 6084 725 6085 755
rect 6085 725 6115 755
rect 6115 725 6116 755
rect 6084 724 6116 725
rect 6084 675 6116 676
rect 6084 645 6085 675
rect 6085 645 6115 675
rect 6115 645 6116 675
rect 6084 644 6116 645
rect 6084 595 6116 596
rect 6084 565 6085 595
rect 6085 565 6115 595
rect 6115 565 6116 595
rect 6084 564 6116 565
rect 6084 195 6116 196
rect 6084 165 6085 195
rect 6085 165 6115 195
rect 6115 165 6116 195
rect 6084 164 6116 165
rect 6084 115 6116 116
rect 6084 85 6085 115
rect 6085 85 6115 115
rect 6115 85 6116 115
rect 6084 84 6116 85
rect 6084 35 6116 36
rect 6084 5 6085 35
rect 6085 5 6115 35
rect 6115 5 6116 35
rect 6084 4 6116 5
rect 6324 13204 6356 13396
rect 6164 12635 6196 12636
rect 6164 12605 6165 12635
rect 6165 12605 6195 12635
rect 6195 12605 6196 12635
rect 6164 12604 6196 12605
rect 6164 12555 6196 12556
rect 6164 12525 6165 12555
rect 6165 12525 6195 12555
rect 6195 12525 6196 12555
rect 6164 12524 6196 12525
rect 6164 12475 6196 12476
rect 6164 12445 6165 12475
rect 6165 12445 6195 12475
rect 6195 12445 6196 12475
rect 6164 12444 6196 12445
rect 6164 12395 6196 12396
rect 6164 12365 6165 12395
rect 6165 12365 6195 12395
rect 6195 12365 6196 12395
rect 6164 12364 6196 12365
rect 6164 12315 6196 12316
rect 6164 12285 6165 12315
rect 6165 12285 6195 12315
rect 6195 12285 6196 12315
rect 6164 12284 6196 12285
rect 6164 12235 6196 12236
rect 6164 12205 6165 12235
rect 6165 12205 6195 12235
rect 6195 12205 6196 12235
rect 6164 12204 6196 12205
rect 6164 12155 6196 12156
rect 6164 12125 6165 12155
rect 6165 12125 6195 12155
rect 6195 12125 6196 12155
rect 6164 12124 6196 12125
rect 6164 11835 6196 11836
rect 6164 11805 6165 11835
rect 6165 11805 6195 11835
rect 6195 11805 6196 11835
rect 6164 11804 6196 11805
rect 6164 11755 6196 11756
rect 6164 11725 6165 11755
rect 6165 11725 6195 11755
rect 6195 11725 6196 11755
rect 6164 11724 6196 11725
rect 6164 11675 6196 11676
rect 6164 11645 6165 11675
rect 6165 11645 6195 11675
rect 6195 11645 6196 11675
rect 6164 11644 6196 11645
rect 6164 11595 6196 11596
rect 6164 11565 6165 11595
rect 6165 11565 6195 11595
rect 6195 11565 6196 11595
rect 6164 11564 6196 11565
rect 6164 11515 6196 11516
rect 6164 11485 6165 11515
rect 6165 11485 6195 11515
rect 6195 11485 6196 11515
rect 6164 11484 6196 11485
rect 6164 11435 6196 11436
rect 6164 11405 6165 11435
rect 6165 11405 6195 11435
rect 6195 11405 6196 11435
rect 6164 11404 6196 11405
rect 6164 10875 6196 10876
rect 6164 10845 6165 10875
rect 6165 10845 6195 10875
rect 6195 10845 6196 10875
rect 6164 10844 6196 10845
rect 6164 10795 6196 10796
rect 6164 10765 6165 10795
rect 6165 10765 6195 10795
rect 6195 10765 6196 10795
rect 6164 10764 6196 10765
rect 6164 10715 6196 10716
rect 6164 10685 6165 10715
rect 6165 10685 6195 10715
rect 6195 10685 6196 10715
rect 6164 10684 6196 10685
rect 6164 10635 6196 10636
rect 6164 10605 6165 10635
rect 6165 10605 6195 10635
rect 6195 10605 6196 10635
rect 6164 10604 6196 10605
rect 6164 10555 6196 10556
rect 6164 10525 6165 10555
rect 6165 10525 6195 10555
rect 6195 10525 6196 10555
rect 6164 10524 6196 10525
rect 6164 10475 6196 10476
rect 6164 10445 6165 10475
rect 6165 10445 6195 10475
rect 6195 10445 6196 10475
rect 6164 10444 6196 10445
rect 6164 10395 6196 10396
rect 6164 10365 6165 10395
rect 6165 10365 6195 10395
rect 6195 10365 6196 10395
rect 6164 10364 6196 10365
rect 6164 10315 6196 10316
rect 6164 10285 6165 10315
rect 6165 10285 6195 10315
rect 6195 10285 6196 10315
rect 6164 10284 6196 10285
rect 6164 10235 6196 10236
rect 6164 10205 6165 10235
rect 6165 10205 6195 10235
rect 6195 10205 6196 10235
rect 6164 10204 6196 10205
rect 6164 10155 6196 10156
rect 6164 10125 6165 10155
rect 6165 10125 6195 10155
rect 6195 10125 6196 10155
rect 6164 10124 6196 10125
rect 6164 10075 6196 10076
rect 6164 10045 6165 10075
rect 6165 10045 6195 10075
rect 6195 10045 6196 10075
rect 6164 10044 6196 10045
rect 6164 9995 6196 9996
rect 6164 9965 6165 9995
rect 6165 9965 6195 9995
rect 6195 9965 6196 9995
rect 6164 9964 6196 9965
rect 6164 9915 6196 9916
rect 6164 9885 6165 9915
rect 6165 9885 6195 9915
rect 6195 9885 6196 9915
rect 6164 9884 6196 9885
rect 6164 9835 6196 9836
rect 6164 9805 6165 9835
rect 6165 9805 6195 9835
rect 6195 9805 6196 9835
rect 6164 9804 6196 9805
rect 6164 9755 6196 9756
rect 6164 9725 6165 9755
rect 6165 9725 6195 9755
rect 6195 9725 6196 9755
rect 6164 9724 6196 9725
rect 6164 9355 6196 9356
rect 6164 9325 6165 9355
rect 6165 9325 6195 9355
rect 6195 9325 6196 9355
rect 6164 9324 6196 9325
rect 6164 9275 6196 9276
rect 6164 9245 6165 9275
rect 6165 9245 6195 9275
rect 6195 9245 6196 9275
rect 6164 9244 6196 9245
rect 6164 9195 6196 9196
rect 6164 9165 6165 9195
rect 6165 9165 6195 9195
rect 6195 9165 6196 9195
rect 6164 9164 6196 9165
rect 6164 8875 6196 8876
rect 6164 8845 6165 8875
rect 6165 8845 6195 8875
rect 6195 8845 6196 8875
rect 6164 8844 6196 8845
rect 6164 8795 6196 8796
rect 6164 8765 6165 8795
rect 6165 8765 6195 8795
rect 6195 8765 6196 8795
rect 6164 8764 6196 8765
rect 6164 8715 6196 8716
rect 6164 8685 6165 8715
rect 6165 8685 6195 8715
rect 6195 8685 6196 8715
rect 6164 8684 6196 8685
rect 6164 8635 6196 8636
rect 6164 8605 6165 8635
rect 6165 8605 6195 8635
rect 6195 8605 6196 8635
rect 6164 8604 6196 8605
rect 6164 8555 6196 8556
rect 6164 8525 6165 8555
rect 6165 8525 6195 8555
rect 6195 8525 6196 8555
rect 6164 8524 6196 8525
rect 6164 7635 6196 7636
rect 6164 7605 6165 7635
rect 6165 7605 6195 7635
rect 6195 7605 6196 7635
rect 6164 7604 6196 7605
rect 6164 7555 6196 7556
rect 6164 7525 6165 7555
rect 6165 7525 6195 7555
rect 6195 7525 6196 7555
rect 6164 7524 6196 7525
rect 6164 7475 6196 7476
rect 6164 7445 6165 7475
rect 6165 7445 6195 7475
rect 6195 7445 6196 7475
rect 6164 7444 6196 7445
rect 6164 7395 6196 7396
rect 6164 7365 6165 7395
rect 6165 7365 6195 7395
rect 6195 7365 6196 7395
rect 6164 7364 6196 7365
rect 6164 7315 6196 7316
rect 6164 7285 6165 7315
rect 6165 7285 6195 7315
rect 6195 7285 6196 7315
rect 6164 7284 6196 7285
rect 6164 7235 6196 7236
rect 6164 7205 6165 7235
rect 6165 7205 6195 7235
rect 6195 7205 6196 7235
rect 6164 7204 6196 7205
rect 6164 7155 6196 7156
rect 6164 7125 6165 7155
rect 6165 7125 6195 7155
rect 6195 7125 6196 7155
rect 6164 7124 6196 7125
rect 6164 7075 6196 7076
rect 6164 7045 6165 7075
rect 6165 7045 6195 7075
rect 6195 7045 6196 7075
rect 6164 7044 6196 7045
rect 6164 6755 6196 6756
rect 6164 6725 6165 6755
rect 6165 6725 6195 6755
rect 6195 6725 6196 6755
rect 6164 6724 6196 6725
rect 6164 6675 6196 6676
rect 6164 6645 6165 6675
rect 6165 6645 6195 6675
rect 6195 6645 6196 6675
rect 6164 6644 6196 6645
rect 6164 6595 6196 6596
rect 6164 6565 6165 6595
rect 6165 6565 6195 6595
rect 6195 6565 6196 6595
rect 6164 6564 6196 6565
rect 6164 6515 6196 6516
rect 6164 6485 6165 6515
rect 6165 6485 6195 6515
rect 6195 6485 6196 6515
rect 6164 6484 6196 6485
rect 6164 6435 6196 6436
rect 6164 6405 6165 6435
rect 6165 6405 6195 6435
rect 6195 6405 6196 6435
rect 6164 6404 6196 6405
rect 6164 6355 6196 6356
rect 6164 6325 6165 6355
rect 6165 6325 6195 6355
rect 6195 6325 6196 6355
rect 6164 6324 6196 6325
rect 6164 5795 6196 5796
rect 6164 5765 6165 5795
rect 6165 5765 6195 5795
rect 6195 5765 6196 5795
rect 6164 5764 6196 5765
rect 6164 5715 6196 5716
rect 6164 5685 6165 5715
rect 6165 5685 6195 5715
rect 6195 5685 6196 5715
rect 6164 5684 6196 5685
rect 6164 5635 6196 5636
rect 6164 5605 6165 5635
rect 6165 5605 6195 5635
rect 6195 5605 6196 5635
rect 6164 5604 6196 5605
rect 6164 5555 6196 5556
rect 6164 5525 6165 5555
rect 6165 5525 6195 5555
rect 6195 5525 6196 5555
rect 6164 5524 6196 5525
rect 6164 5475 6196 5476
rect 6164 5445 6165 5475
rect 6165 5445 6195 5475
rect 6195 5445 6196 5475
rect 6164 5444 6196 5445
rect 6164 5395 6196 5396
rect 6164 5365 6165 5395
rect 6165 5365 6195 5395
rect 6195 5365 6196 5395
rect 6164 5364 6196 5365
rect 6164 5315 6196 5316
rect 6164 5285 6165 5315
rect 6165 5285 6195 5315
rect 6195 5285 6196 5315
rect 6164 5284 6196 5285
rect 6164 5235 6196 5236
rect 6164 5205 6165 5235
rect 6165 5205 6195 5235
rect 6195 5205 6196 5235
rect 6164 5204 6196 5205
rect 6164 5155 6196 5156
rect 6164 5125 6165 5155
rect 6165 5125 6195 5155
rect 6195 5125 6196 5155
rect 6164 5124 6196 5125
rect 6164 5075 6196 5076
rect 6164 5045 6165 5075
rect 6165 5045 6195 5075
rect 6195 5045 6196 5075
rect 6164 5044 6196 5045
rect 6164 4995 6196 4996
rect 6164 4965 6165 4995
rect 6165 4965 6195 4995
rect 6195 4965 6196 4995
rect 6164 4964 6196 4965
rect 6164 4435 6196 4436
rect 6164 4405 6165 4435
rect 6165 4405 6195 4435
rect 6195 4405 6196 4435
rect 6164 4404 6196 4405
rect 6164 4355 6196 4356
rect 6164 4325 6165 4355
rect 6165 4325 6195 4355
rect 6195 4325 6196 4355
rect 6164 4324 6196 4325
rect 6164 4275 6196 4276
rect 6164 4245 6165 4275
rect 6165 4245 6195 4275
rect 6195 4245 6196 4275
rect 6164 4244 6196 4245
rect 6164 4195 6196 4196
rect 6164 4165 6165 4195
rect 6165 4165 6195 4195
rect 6195 4165 6196 4195
rect 6164 4164 6196 4165
rect 6164 4115 6196 4116
rect 6164 4085 6165 4115
rect 6165 4085 6195 4115
rect 6195 4085 6196 4115
rect 6164 4084 6196 4085
rect 6164 4035 6196 4036
rect 6164 4005 6165 4035
rect 6165 4005 6195 4035
rect 6195 4005 6196 4035
rect 6164 4004 6196 4005
rect 6164 3955 6196 3956
rect 6164 3925 6165 3955
rect 6165 3925 6195 3955
rect 6195 3925 6196 3955
rect 6164 3924 6196 3925
rect 6164 3155 6196 3156
rect 6164 3125 6165 3155
rect 6165 3125 6195 3155
rect 6195 3125 6196 3155
rect 6164 3124 6196 3125
rect 6164 3075 6196 3076
rect 6164 3045 6165 3075
rect 6165 3045 6195 3075
rect 6195 3045 6196 3075
rect 6164 3044 6196 3045
rect 6164 2995 6196 2996
rect 6164 2965 6165 2995
rect 6165 2965 6195 2995
rect 6195 2965 6196 2995
rect 6164 2964 6196 2965
rect 6164 2915 6196 2916
rect 6164 2885 6165 2915
rect 6165 2885 6195 2915
rect 6195 2885 6196 2915
rect 6164 2884 6196 2885
rect 6164 2835 6196 2836
rect 6164 2805 6165 2835
rect 6165 2805 6195 2835
rect 6195 2805 6196 2835
rect 6164 2804 6196 2805
rect 6164 2755 6196 2756
rect 6164 2725 6165 2755
rect 6165 2725 6195 2755
rect 6195 2725 6196 2755
rect 6164 2724 6196 2725
rect 6164 2675 6196 2676
rect 6164 2645 6165 2675
rect 6165 2645 6195 2675
rect 6195 2645 6196 2675
rect 6164 2644 6196 2645
rect 6164 2595 6196 2596
rect 6164 2565 6165 2595
rect 6165 2565 6195 2595
rect 6195 2565 6196 2595
rect 6164 2564 6196 2565
rect 6164 2515 6196 2516
rect 6164 2485 6165 2515
rect 6165 2485 6195 2515
rect 6195 2485 6196 2515
rect 6164 2484 6196 2485
rect 6164 2435 6196 2436
rect 6164 2405 6165 2435
rect 6165 2405 6195 2435
rect 6195 2405 6196 2435
rect 6164 2404 6196 2405
rect 6164 2355 6196 2356
rect 6164 2325 6165 2355
rect 6165 2325 6195 2355
rect 6195 2325 6196 2355
rect 6164 2324 6196 2325
rect 6164 2275 6196 2276
rect 6164 2245 6165 2275
rect 6165 2245 6195 2275
rect 6195 2245 6196 2275
rect 6164 2244 6196 2245
rect 6164 2195 6196 2196
rect 6164 2165 6165 2195
rect 6165 2165 6195 2195
rect 6195 2165 6196 2195
rect 6164 2164 6196 2165
rect 6164 2115 6196 2116
rect 6164 2085 6165 2115
rect 6165 2085 6195 2115
rect 6195 2085 6196 2115
rect 6164 2084 6196 2085
rect 6164 2035 6196 2036
rect 6164 2005 6165 2035
rect 6165 2005 6195 2035
rect 6195 2005 6196 2035
rect 6164 2004 6196 2005
rect 6164 1635 6196 1636
rect 6164 1605 6165 1635
rect 6165 1605 6195 1635
rect 6195 1605 6196 1635
rect 6164 1604 6196 1605
rect 6164 1555 6196 1556
rect 6164 1525 6165 1555
rect 6165 1525 6195 1555
rect 6195 1525 6196 1555
rect 6164 1524 6196 1525
rect 6164 1475 6196 1476
rect 6164 1445 6165 1475
rect 6165 1445 6195 1475
rect 6195 1445 6196 1475
rect 6164 1444 6196 1445
rect 6164 1395 6196 1396
rect 6164 1365 6165 1395
rect 6165 1365 6195 1395
rect 6195 1365 6196 1395
rect 6164 1364 6196 1365
rect 6164 1315 6196 1316
rect 6164 1285 6165 1315
rect 6165 1285 6195 1315
rect 6195 1285 6196 1315
rect 6164 1284 6196 1285
rect 6164 1235 6196 1236
rect 6164 1205 6165 1235
rect 6165 1205 6195 1235
rect 6195 1205 6196 1235
rect 6164 1204 6196 1205
rect 6164 1155 6196 1156
rect 6164 1125 6165 1155
rect 6165 1125 6195 1155
rect 6195 1125 6196 1155
rect 6164 1124 6196 1125
rect 6164 1075 6196 1076
rect 6164 1045 6165 1075
rect 6165 1045 6195 1075
rect 6195 1045 6196 1075
rect 6164 1044 6196 1045
rect 6164 755 6196 756
rect 6164 725 6165 755
rect 6165 725 6195 755
rect 6195 725 6196 755
rect 6164 724 6196 725
rect 6164 675 6196 676
rect 6164 645 6165 675
rect 6165 645 6195 675
rect 6195 645 6196 675
rect 6164 644 6196 645
rect 6164 595 6196 596
rect 6164 565 6165 595
rect 6165 565 6195 595
rect 6195 565 6196 595
rect 6164 564 6196 565
rect 6164 195 6196 196
rect 6164 165 6165 195
rect 6165 165 6195 195
rect 6195 165 6196 195
rect 6164 164 6196 165
rect 6164 115 6196 116
rect 6164 85 6165 115
rect 6165 85 6195 115
rect 6195 85 6196 115
rect 6164 84 6196 85
rect 6164 35 6196 36
rect 6164 5 6165 35
rect 6165 5 6195 35
rect 6195 5 6196 35
rect 6164 4 6196 5
rect 6324 12635 6356 12636
rect 6324 12605 6325 12635
rect 6325 12605 6355 12635
rect 6355 12605 6356 12635
rect 6324 12604 6356 12605
rect 6324 12555 6356 12556
rect 6324 12525 6325 12555
rect 6325 12525 6355 12555
rect 6355 12525 6356 12555
rect 6324 12524 6356 12525
rect 6324 12475 6356 12476
rect 6324 12445 6325 12475
rect 6325 12445 6355 12475
rect 6355 12445 6356 12475
rect 6324 12444 6356 12445
rect 6324 12395 6356 12396
rect 6324 12365 6325 12395
rect 6325 12365 6355 12395
rect 6355 12365 6356 12395
rect 6324 12364 6356 12365
rect 6324 12315 6356 12316
rect 6324 12285 6325 12315
rect 6325 12285 6355 12315
rect 6355 12285 6356 12315
rect 6324 12284 6356 12285
rect 6324 12235 6356 12236
rect 6324 12205 6325 12235
rect 6325 12205 6355 12235
rect 6355 12205 6356 12235
rect 6324 12204 6356 12205
rect 6324 12155 6356 12156
rect 6324 12125 6325 12155
rect 6325 12125 6355 12155
rect 6355 12125 6356 12155
rect 6324 12124 6356 12125
rect 6324 11835 6356 11836
rect 6324 11805 6325 11835
rect 6325 11805 6355 11835
rect 6355 11805 6356 11835
rect 6324 11804 6356 11805
rect 6324 11755 6356 11756
rect 6324 11725 6325 11755
rect 6325 11725 6355 11755
rect 6355 11725 6356 11755
rect 6324 11724 6356 11725
rect 6324 11675 6356 11676
rect 6324 11645 6325 11675
rect 6325 11645 6355 11675
rect 6355 11645 6356 11675
rect 6324 11644 6356 11645
rect 6324 11595 6356 11596
rect 6324 11565 6325 11595
rect 6325 11565 6355 11595
rect 6355 11565 6356 11595
rect 6324 11564 6356 11565
rect 6324 11515 6356 11516
rect 6324 11485 6325 11515
rect 6325 11485 6355 11515
rect 6355 11485 6356 11515
rect 6324 11484 6356 11485
rect 6324 11435 6356 11436
rect 6324 11405 6325 11435
rect 6325 11405 6355 11435
rect 6355 11405 6356 11435
rect 6324 11404 6356 11405
rect 6324 10875 6356 10876
rect 6324 10845 6325 10875
rect 6325 10845 6355 10875
rect 6355 10845 6356 10875
rect 6324 10844 6356 10845
rect 6324 10795 6356 10796
rect 6324 10765 6325 10795
rect 6325 10765 6355 10795
rect 6355 10765 6356 10795
rect 6324 10764 6356 10765
rect 6324 10715 6356 10716
rect 6324 10685 6325 10715
rect 6325 10685 6355 10715
rect 6355 10685 6356 10715
rect 6324 10684 6356 10685
rect 6324 10635 6356 10636
rect 6324 10605 6325 10635
rect 6325 10605 6355 10635
rect 6355 10605 6356 10635
rect 6324 10604 6356 10605
rect 6324 10555 6356 10556
rect 6324 10525 6325 10555
rect 6325 10525 6355 10555
rect 6355 10525 6356 10555
rect 6324 10524 6356 10525
rect 6324 10475 6356 10476
rect 6324 10445 6325 10475
rect 6325 10445 6355 10475
rect 6355 10445 6356 10475
rect 6324 10444 6356 10445
rect 6324 10395 6356 10396
rect 6324 10365 6325 10395
rect 6325 10365 6355 10395
rect 6355 10365 6356 10395
rect 6324 10364 6356 10365
rect 6324 10315 6356 10316
rect 6324 10285 6325 10315
rect 6325 10285 6355 10315
rect 6355 10285 6356 10315
rect 6324 10284 6356 10285
rect 6324 10235 6356 10236
rect 6324 10205 6325 10235
rect 6325 10205 6355 10235
rect 6355 10205 6356 10235
rect 6324 10204 6356 10205
rect 6324 10155 6356 10156
rect 6324 10125 6325 10155
rect 6325 10125 6355 10155
rect 6355 10125 6356 10155
rect 6324 10124 6356 10125
rect 6324 10075 6356 10076
rect 6324 10045 6325 10075
rect 6325 10045 6355 10075
rect 6355 10045 6356 10075
rect 6324 10044 6356 10045
rect 6324 9995 6356 9996
rect 6324 9965 6325 9995
rect 6325 9965 6355 9995
rect 6355 9965 6356 9995
rect 6324 9964 6356 9965
rect 6324 9915 6356 9916
rect 6324 9885 6325 9915
rect 6325 9885 6355 9915
rect 6355 9885 6356 9915
rect 6324 9884 6356 9885
rect 6324 9835 6356 9836
rect 6324 9805 6325 9835
rect 6325 9805 6355 9835
rect 6355 9805 6356 9835
rect 6324 9804 6356 9805
rect 6324 9755 6356 9756
rect 6324 9725 6325 9755
rect 6325 9725 6355 9755
rect 6355 9725 6356 9755
rect 6324 9724 6356 9725
rect 6324 9355 6356 9356
rect 6324 9325 6325 9355
rect 6325 9325 6355 9355
rect 6355 9325 6356 9355
rect 6324 9324 6356 9325
rect 6324 9275 6356 9276
rect 6324 9245 6325 9275
rect 6325 9245 6355 9275
rect 6355 9245 6356 9275
rect 6324 9244 6356 9245
rect 6324 9195 6356 9196
rect 6324 9165 6325 9195
rect 6325 9165 6355 9195
rect 6355 9165 6356 9195
rect 6324 9164 6356 9165
rect 6324 8875 6356 8876
rect 6324 8845 6325 8875
rect 6325 8845 6355 8875
rect 6355 8845 6356 8875
rect 6324 8844 6356 8845
rect 6324 8795 6356 8796
rect 6324 8765 6325 8795
rect 6325 8765 6355 8795
rect 6355 8765 6356 8795
rect 6324 8764 6356 8765
rect 6324 8715 6356 8716
rect 6324 8685 6325 8715
rect 6325 8685 6355 8715
rect 6355 8685 6356 8715
rect 6324 8684 6356 8685
rect 6324 8635 6356 8636
rect 6324 8605 6325 8635
rect 6325 8605 6355 8635
rect 6355 8605 6356 8635
rect 6324 8604 6356 8605
rect 6324 8555 6356 8556
rect 6324 8525 6325 8555
rect 6325 8525 6355 8555
rect 6355 8525 6356 8555
rect 6324 8524 6356 8525
rect 6324 7635 6356 7636
rect 6324 7605 6325 7635
rect 6325 7605 6355 7635
rect 6355 7605 6356 7635
rect 6324 7604 6356 7605
rect 6324 7555 6356 7556
rect 6324 7525 6325 7555
rect 6325 7525 6355 7555
rect 6355 7525 6356 7555
rect 6324 7524 6356 7525
rect 6324 7475 6356 7476
rect 6324 7445 6325 7475
rect 6325 7445 6355 7475
rect 6355 7445 6356 7475
rect 6324 7444 6356 7445
rect 6324 7395 6356 7396
rect 6324 7365 6325 7395
rect 6325 7365 6355 7395
rect 6355 7365 6356 7395
rect 6324 7364 6356 7365
rect 6324 7315 6356 7316
rect 6324 7285 6325 7315
rect 6325 7285 6355 7315
rect 6355 7285 6356 7315
rect 6324 7284 6356 7285
rect 6324 7235 6356 7236
rect 6324 7205 6325 7235
rect 6325 7205 6355 7235
rect 6355 7205 6356 7235
rect 6324 7204 6356 7205
rect 6324 7155 6356 7156
rect 6324 7125 6325 7155
rect 6325 7125 6355 7155
rect 6355 7125 6356 7155
rect 6324 7124 6356 7125
rect 6324 7075 6356 7076
rect 6324 7045 6325 7075
rect 6325 7045 6355 7075
rect 6355 7045 6356 7075
rect 6324 7044 6356 7045
rect 6324 6755 6356 6756
rect 6324 6725 6325 6755
rect 6325 6725 6355 6755
rect 6355 6725 6356 6755
rect 6324 6724 6356 6725
rect 6324 6675 6356 6676
rect 6324 6645 6325 6675
rect 6325 6645 6355 6675
rect 6355 6645 6356 6675
rect 6324 6644 6356 6645
rect 6324 6595 6356 6596
rect 6324 6565 6325 6595
rect 6325 6565 6355 6595
rect 6355 6565 6356 6595
rect 6324 6564 6356 6565
rect 6324 6515 6356 6516
rect 6324 6485 6325 6515
rect 6325 6485 6355 6515
rect 6355 6485 6356 6515
rect 6324 6484 6356 6485
rect 6324 6435 6356 6436
rect 6324 6405 6325 6435
rect 6325 6405 6355 6435
rect 6355 6405 6356 6435
rect 6324 6404 6356 6405
rect 6324 6355 6356 6356
rect 6324 6325 6325 6355
rect 6325 6325 6355 6355
rect 6355 6325 6356 6355
rect 6324 6324 6356 6325
rect 6324 5795 6356 5796
rect 6324 5765 6325 5795
rect 6325 5765 6355 5795
rect 6355 5765 6356 5795
rect 6324 5764 6356 5765
rect 6324 5715 6356 5716
rect 6324 5685 6325 5715
rect 6325 5685 6355 5715
rect 6355 5685 6356 5715
rect 6324 5684 6356 5685
rect 6324 5635 6356 5636
rect 6324 5605 6325 5635
rect 6325 5605 6355 5635
rect 6355 5605 6356 5635
rect 6324 5604 6356 5605
rect 6324 5555 6356 5556
rect 6324 5525 6325 5555
rect 6325 5525 6355 5555
rect 6355 5525 6356 5555
rect 6324 5524 6356 5525
rect 6324 5475 6356 5476
rect 6324 5445 6325 5475
rect 6325 5445 6355 5475
rect 6355 5445 6356 5475
rect 6324 5444 6356 5445
rect 6324 5395 6356 5396
rect 6324 5365 6325 5395
rect 6325 5365 6355 5395
rect 6355 5365 6356 5395
rect 6324 5364 6356 5365
rect 6324 5315 6356 5316
rect 6324 5285 6325 5315
rect 6325 5285 6355 5315
rect 6355 5285 6356 5315
rect 6324 5284 6356 5285
rect 6324 5235 6356 5236
rect 6324 5205 6325 5235
rect 6325 5205 6355 5235
rect 6355 5205 6356 5235
rect 6324 5204 6356 5205
rect 6324 5155 6356 5156
rect 6324 5125 6325 5155
rect 6325 5125 6355 5155
rect 6355 5125 6356 5155
rect 6324 5124 6356 5125
rect 6324 5075 6356 5076
rect 6324 5045 6325 5075
rect 6325 5045 6355 5075
rect 6355 5045 6356 5075
rect 6324 5044 6356 5045
rect 6324 4995 6356 4996
rect 6324 4965 6325 4995
rect 6325 4965 6355 4995
rect 6355 4965 6356 4995
rect 6324 4964 6356 4965
rect 6324 4435 6356 4436
rect 6324 4405 6325 4435
rect 6325 4405 6355 4435
rect 6355 4405 6356 4435
rect 6324 4404 6356 4405
rect 6324 4355 6356 4356
rect 6324 4325 6325 4355
rect 6325 4325 6355 4355
rect 6355 4325 6356 4355
rect 6324 4324 6356 4325
rect 6324 4275 6356 4276
rect 6324 4245 6325 4275
rect 6325 4245 6355 4275
rect 6355 4245 6356 4275
rect 6324 4244 6356 4245
rect 6324 4195 6356 4196
rect 6324 4165 6325 4195
rect 6325 4165 6355 4195
rect 6355 4165 6356 4195
rect 6324 4164 6356 4165
rect 6324 4115 6356 4116
rect 6324 4085 6325 4115
rect 6325 4085 6355 4115
rect 6355 4085 6356 4115
rect 6324 4084 6356 4085
rect 6324 4035 6356 4036
rect 6324 4005 6325 4035
rect 6325 4005 6355 4035
rect 6355 4005 6356 4035
rect 6324 4004 6356 4005
rect 6324 3955 6356 3956
rect 6324 3925 6325 3955
rect 6325 3925 6355 3955
rect 6355 3925 6356 3955
rect 6324 3924 6356 3925
rect 6324 3155 6356 3156
rect 6324 3125 6325 3155
rect 6325 3125 6355 3155
rect 6355 3125 6356 3155
rect 6324 3124 6356 3125
rect 6324 3075 6356 3076
rect 6324 3045 6325 3075
rect 6325 3045 6355 3075
rect 6355 3045 6356 3075
rect 6324 3044 6356 3045
rect 6324 2995 6356 2996
rect 6324 2965 6325 2995
rect 6325 2965 6355 2995
rect 6355 2965 6356 2995
rect 6324 2964 6356 2965
rect 6324 2915 6356 2916
rect 6324 2885 6325 2915
rect 6325 2885 6355 2915
rect 6355 2885 6356 2915
rect 6324 2884 6356 2885
rect 6324 2835 6356 2836
rect 6324 2805 6325 2835
rect 6325 2805 6355 2835
rect 6355 2805 6356 2835
rect 6324 2804 6356 2805
rect 6324 2755 6356 2756
rect 6324 2725 6325 2755
rect 6325 2725 6355 2755
rect 6355 2725 6356 2755
rect 6324 2724 6356 2725
rect 6324 2675 6356 2676
rect 6324 2645 6325 2675
rect 6325 2645 6355 2675
rect 6355 2645 6356 2675
rect 6324 2644 6356 2645
rect 6324 2595 6356 2596
rect 6324 2565 6325 2595
rect 6325 2565 6355 2595
rect 6355 2565 6356 2595
rect 6324 2564 6356 2565
rect 6324 2515 6356 2516
rect 6324 2485 6325 2515
rect 6325 2485 6355 2515
rect 6355 2485 6356 2515
rect 6324 2484 6356 2485
rect 6324 2435 6356 2436
rect 6324 2405 6325 2435
rect 6325 2405 6355 2435
rect 6355 2405 6356 2435
rect 6324 2404 6356 2405
rect 6324 2355 6356 2356
rect 6324 2325 6325 2355
rect 6325 2325 6355 2355
rect 6355 2325 6356 2355
rect 6324 2324 6356 2325
rect 6324 2275 6356 2276
rect 6324 2245 6325 2275
rect 6325 2245 6355 2275
rect 6355 2245 6356 2275
rect 6324 2244 6356 2245
rect 6324 2195 6356 2196
rect 6324 2165 6325 2195
rect 6325 2165 6355 2195
rect 6355 2165 6356 2195
rect 6324 2164 6356 2165
rect 6324 2115 6356 2116
rect 6324 2085 6325 2115
rect 6325 2085 6355 2115
rect 6355 2085 6356 2115
rect 6324 2084 6356 2085
rect 6324 2035 6356 2036
rect 6324 2005 6325 2035
rect 6325 2005 6355 2035
rect 6355 2005 6356 2035
rect 6324 2004 6356 2005
rect 6324 1635 6356 1636
rect 6324 1605 6325 1635
rect 6325 1605 6355 1635
rect 6355 1605 6356 1635
rect 6324 1604 6356 1605
rect 6324 1555 6356 1556
rect 6324 1525 6325 1555
rect 6325 1525 6355 1555
rect 6355 1525 6356 1555
rect 6324 1524 6356 1525
rect 6324 1475 6356 1476
rect 6324 1445 6325 1475
rect 6325 1445 6355 1475
rect 6355 1445 6356 1475
rect 6324 1444 6356 1445
rect 6324 1395 6356 1396
rect 6324 1365 6325 1395
rect 6325 1365 6355 1395
rect 6355 1365 6356 1395
rect 6324 1364 6356 1365
rect 6324 1315 6356 1316
rect 6324 1285 6325 1315
rect 6325 1285 6355 1315
rect 6355 1285 6356 1315
rect 6324 1284 6356 1285
rect 6324 1235 6356 1236
rect 6324 1205 6325 1235
rect 6325 1205 6355 1235
rect 6355 1205 6356 1235
rect 6324 1204 6356 1205
rect 6324 1155 6356 1156
rect 6324 1125 6325 1155
rect 6325 1125 6355 1155
rect 6355 1125 6356 1155
rect 6324 1124 6356 1125
rect 6324 1075 6356 1076
rect 6324 1045 6325 1075
rect 6325 1045 6355 1075
rect 6355 1045 6356 1075
rect 6324 1044 6356 1045
rect 6324 755 6356 756
rect 6324 725 6325 755
rect 6325 725 6355 755
rect 6355 725 6356 755
rect 6324 724 6356 725
rect 6324 675 6356 676
rect 6324 645 6325 675
rect 6325 645 6355 675
rect 6355 645 6356 675
rect 6324 644 6356 645
rect 6324 595 6356 596
rect 6324 565 6325 595
rect 6325 565 6355 595
rect 6355 565 6356 595
rect 6324 564 6356 565
rect 6324 195 6356 196
rect 6324 165 6325 195
rect 6325 165 6355 195
rect 6355 165 6356 195
rect 6324 164 6356 165
rect 6324 115 6356 116
rect 6324 85 6325 115
rect 6325 85 6355 115
rect 6355 85 6356 115
rect 6324 84 6356 85
rect 6324 35 6356 36
rect 6324 5 6325 35
rect 6325 5 6355 35
rect 6355 5 6356 35
rect 6324 4 6356 5
<< mimcap >>
rect 520 16600 1520 16640
rect 520 15680 560 16600
rect 1480 15680 1520 16600
rect 520 15640 1520 15680
rect 1640 16600 2640 16640
rect 1640 15680 1680 16600
rect 2600 15680 2640 16600
rect 1640 15640 2640 15680
rect 2760 16600 3760 16640
rect 2760 15680 2800 16600
rect 3720 15680 3760 16600
rect 2760 15640 3760 15680
rect 3880 16600 4880 16640
rect 3880 15680 3920 16600
rect 4840 15680 4880 16600
rect 3880 15640 4880 15680
rect 5720 16600 6720 16640
rect 5720 15680 5760 16600
rect 6680 15680 6720 16600
rect 5720 15640 6720 15680
rect 6840 16600 7840 16640
rect 6840 15680 6880 16600
rect 7800 15680 7840 16600
rect 6840 15640 7840 15680
rect 7960 16600 8960 16640
rect 7960 15680 8000 16600
rect 8920 15680 8960 16600
rect 7960 15640 8960 15680
rect 9080 16600 10080 16640
rect 9080 15680 9120 16600
rect 10040 15680 10080 16600
rect 9080 15640 10080 15680
rect 520 15160 1520 15200
rect 520 14240 560 15160
rect 1480 14240 1520 15160
rect 520 14200 1520 14240
rect 1640 15160 2640 15200
rect 1640 14240 1680 15160
rect 2600 14240 2640 15160
rect 1640 14200 2640 14240
rect 2760 15160 3760 15200
rect 2760 14240 2800 15160
rect 3720 14240 3760 15160
rect 2760 14200 3760 14240
rect 3880 15160 4880 15200
rect 3880 14240 3920 15160
rect 4840 14240 4880 15160
rect 3880 14200 4880 14240
rect 5720 15160 6720 15200
rect 5720 14240 5760 15160
rect 6680 14240 6720 15160
rect 5720 14200 6720 14240
rect 6840 15160 7840 15200
rect 6840 14240 6880 15160
rect 7800 14240 7840 15160
rect 6840 14200 7840 14240
rect 7960 15160 8960 15200
rect 7960 14240 8000 15160
rect 8920 14240 8960 15160
rect 7960 14200 8960 14240
rect 9080 15160 10080 15200
rect 9080 14240 9120 15160
rect 10040 14240 10080 15160
rect 9080 14200 10080 14240
<< mimcapcontact >>
rect 560 15680 1480 16600
rect 1680 15680 2600 16600
rect 2800 15680 3720 16600
rect 3920 15680 4840 16600
rect 5760 15680 6680 16600
rect 6880 15680 7800 16600
rect 8000 15680 8920 16600
rect 9120 15680 10040 16600
rect 560 14240 1480 15160
rect 1680 14240 2600 15160
rect 2800 14240 3720 15160
rect 3920 14240 4840 15160
rect 5760 14240 6680 15160
rect 6880 14240 7800 15160
rect 8000 14240 8920 15160
rect 9120 14240 10040 15160
<< metal4 >>
rect 0 16916 10600 16920
rect 0 16884 4 16916
rect 36 16884 324 16916
rect 356 16884 10244 16916
rect 10276 16884 10564 16916
rect 10596 16884 10600 16916
rect 0 16880 10600 16884
rect 0 16836 10600 16840
rect 0 16804 84 16836
rect 116 16804 244 16836
rect 276 16804 404 16836
rect 436 16804 10164 16836
rect 10196 16804 10324 16836
rect 10356 16804 10484 16836
rect 10516 16804 10600 16836
rect 0 16800 10600 16804
rect 80 16756 10520 16760
rect 80 16724 164 16756
rect 196 16724 484 16756
rect 516 16724 1524 16756
rect 1556 16724 1604 16756
rect 1636 16724 2644 16756
rect 2676 16724 2724 16756
rect 2756 16724 3764 16756
rect 3796 16724 3844 16756
rect 3876 16724 4884 16756
rect 4916 16724 5684 16756
rect 5716 16724 6724 16756
rect 6756 16724 6804 16756
rect 6836 16724 7844 16756
rect 7876 16724 7924 16756
rect 7956 16724 8964 16756
rect 8996 16724 9044 16756
rect 9076 16724 10084 16756
rect 10116 16724 10404 16756
rect 10436 16724 10520 16756
rect 80 16720 10520 16724
rect 480 16600 1560 16680
rect 480 15680 560 16600
rect 1480 15680 1560 16600
rect 480 15600 1560 15680
rect 480 15560 520 15600
rect 1520 15560 1560 15600
rect 1600 16600 2680 16680
rect 1600 15680 1680 16600
rect 2600 15680 2680 16600
rect 1600 15600 2680 15680
rect 1600 15560 1640 15600
rect 2640 15560 2680 15600
rect 2720 16600 3800 16680
rect 2720 15680 2800 16600
rect 3720 15680 3800 16600
rect 2720 15600 3800 15680
rect 2720 15560 2760 15600
rect 3760 15560 3800 15600
rect 3840 16600 4920 16680
rect 3840 15680 3920 16600
rect 4840 15680 4920 16600
rect 3840 15600 4920 15680
rect 3840 15560 3880 15600
rect 4880 15560 4920 15600
rect 5680 16600 6760 16680
rect 5680 15680 5760 16600
rect 6680 15680 6760 16600
rect 5680 15600 6760 15680
rect 5680 15560 5720 15600
rect 6720 15560 6760 15600
rect 6800 16600 7880 16680
rect 6800 15680 6880 16600
rect 7800 15680 7880 16600
rect 6800 15600 7880 15680
rect 6800 15560 6840 15600
rect 7840 15560 7880 15600
rect 7920 16600 9000 16680
rect 7920 15680 8000 16600
rect 8920 15680 9000 16600
rect 7920 15600 9000 15680
rect 7920 15560 7960 15600
rect 8960 15560 9000 15600
rect 9040 16600 10120 16680
rect 9040 15680 9120 16600
rect 10040 15680 10120 16600
rect 9040 15600 10120 15680
rect 9040 15560 9080 15600
rect 10080 15560 10120 15600
rect 0 15556 10600 15560
rect 0 15524 84 15556
rect 116 15524 244 15556
rect 276 15524 404 15556
rect 436 15524 10164 15556
rect 10196 15524 10324 15556
rect 10356 15524 10484 15556
rect 10516 15524 10600 15556
rect 0 15520 10600 15524
rect 0 15476 10600 15480
rect 0 15444 4 15476
rect 36 15444 324 15476
rect 356 15444 10244 15476
rect 10276 15444 10564 15476
rect 10596 15444 10600 15476
rect 0 15440 10600 15444
rect 400 15396 10200 15400
rect 400 15364 404 15396
rect 436 15364 4964 15396
rect 4996 15364 5124 15396
rect 5156 15364 5284 15396
rect 5316 15364 5444 15396
rect 5476 15364 5604 15396
rect 5636 15364 10164 15396
rect 10196 15364 10200 15396
rect 400 15360 10200 15364
rect 480 15316 5240 15320
rect 480 15284 484 15316
rect 516 15284 1524 15316
rect 1556 15284 1604 15316
rect 1636 15284 2644 15316
rect 2676 15284 2724 15316
rect 2756 15284 3764 15316
rect 3796 15284 3844 15316
rect 3876 15284 4884 15316
rect 4916 15284 5204 15316
rect 5236 15284 5240 15316
rect 480 15280 5240 15284
rect 5360 15316 10160 15320
rect 5360 15284 5364 15316
rect 5396 15284 5684 15316
rect 5716 15284 6724 15316
rect 6756 15284 6804 15316
rect 6836 15284 7844 15316
rect 7876 15284 7924 15316
rect 7956 15284 8964 15316
rect 8996 15284 9044 15316
rect 9076 15284 10084 15316
rect 10116 15284 10160 15316
rect 5360 15280 10160 15284
rect 480 15160 1560 15240
rect 480 14240 560 15160
rect 1480 14240 1560 15160
rect 480 14160 1560 14240
rect 480 14120 520 14160
rect 1520 14120 1560 14160
rect 1600 15160 2680 15240
rect 1600 14240 1680 15160
rect 2600 14240 2680 15160
rect 1600 14160 2680 14240
rect 1600 14120 1640 14160
rect 2640 14120 2680 14160
rect 2720 15160 3800 15240
rect 2720 14240 2800 15160
rect 3720 14240 3800 15160
rect 2720 14160 3800 14240
rect 2720 14120 2760 14160
rect 3760 14120 3800 14160
rect 3840 15160 4920 15240
rect 3840 14240 3920 15160
rect 4840 14240 4920 15160
rect 3840 14160 4920 14240
rect 3840 14120 3880 14160
rect 4880 14120 4920 14160
rect 5680 15160 6760 15240
rect 5680 14240 5760 15160
rect 6680 14240 6760 15160
rect 5680 14160 6760 14240
rect 5680 14120 5720 14160
rect 6720 14120 6760 14160
rect 6800 15160 7880 15240
rect 6800 14240 6880 15160
rect 7800 14240 7880 15160
rect 6800 14160 7880 14240
rect 6800 14120 6840 14160
rect 7840 14120 7880 14160
rect 7920 15160 9000 15240
rect 7920 14240 8000 15160
rect 8920 14240 9000 15160
rect 7920 14160 9000 14240
rect 7920 14120 7960 14160
rect 8960 14120 9000 14160
rect 9040 15160 10120 15240
rect 9040 14240 9120 15160
rect 10040 14240 10120 15160
rect 9040 14160 10120 14240
rect 9040 14120 9080 14160
rect 10080 14120 10120 14160
rect 400 14116 10200 14120
rect 400 14084 404 14116
rect 436 14084 4964 14116
rect 4996 14084 5124 14116
rect 5156 14084 5284 14116
rect 5316 14084 5444 14116
rect 5476 14084 5604 14116
rect 5636 14084 10164 14116
rect 10196 14084 10200 14116
rect 400 14080 10200 14084
rect 0 14036 10600 14040
rect 0 14004 4 14036
rect 36 14004 324 14036
rect 356 14004 5044 14036
rect 5076 14004 5524 14036
rect 5556 14004 10244 14036
rect 10276 14004 10564 14036
rect 10596 14004 10600 14036
rect 0 14000 10600 14004
rect 0 13956 10600 13960
rect 0 13924 84 13956
rect 116 13924 244 13956
rect 276 13924 4484 13956
rect 4516 13924 4644 13956
rect 4676 13924 10324 13956
rect 10356 13924 10484 13956
rect 10516 13924 10600 13956
rect 0 13920 10600 13924
rect 0 13876 10600 13880
rect 0 13844 164 13876
rect 196 13844 4564 13876
rect 4596 13844 10404 13876
rect 10436 13844 10600 13876
rect 0 13840 10600 13844
rect 0 13796 10600 13800
rect 0 13764 84 13796
rect 116 13764 244 13796
rect 276 13764 4484 13796
rect 4516 13764 4644 13796
rect 4676 13764 10324 13796
rect 10356 13764 10484 13796
rect 10516 13764 10600 13796
rect 0 13760 10600 13764
rect 0 13716 10600 13720
rect 0 13684 4 13716
rect 36 13684 324 13716
rect 356 13684 5044 13716
rect 5076 13684 5524 13716
rect 5556 13684 10244 13716
rect 10276 13684 10564 13716
rect 10596 13684 10600 13716
rect 0 13680 10600 13684
rect 0 13636 10600 13640
rect 0 13600 4244 13636
rect 0 13480 1560 13600
rect 1680 13480 2520 13600
rect 2640 13480 4244 13600
rect 0 13444 4244 13480
rect 4276 13444 4404 13636
rect 4436 13600 10600 13636
rect 4436 13480 7960 13600
rect 8080 13480 8920 13600
rect 9040 13480 10600 13600
rect 4436 13444 10600 13480
rect 0 13440 10600 13444
rect 0 13396 10600 13400
rect 0 13360 4724 13396
rect 0 13240 1080 13360
rect 1200 13240 2040 13360
rect 2160 13240 3000 13360
rect 3120 13240 4724 13360
rect 0 13204 4724 13240
rect 4756 13204 4884 13396
rect 4916 13204 5044 13396
rect 5076 13204 5524 13396
rect 5556 13204 5684 13396
rect 5716 13204 5844 13396
rect 5876 13204 6164 13396
rect 6196 13204 6324 13396
rect 6356 13360 10600 13396
rect 6356 13240 7480 13360
rect 7600 13240 8440 13360
rect 8560 13240 9400 13360
rect 9520 13240 10600 13360
rect 6356 13204 10600 13240
rect 0 13200 10600 13204
rect 0 13156 10600 13160
rect 0 13120 4484 13156
rect 0 13000 600 13120
rect 720 13000 3480 13120
rect 3600 13000 4484 13120
rect 0 12964 4484 13000
rect 4516 12964 4644 13156
rect 4676 13120 10600 13156
rect 4676 13000 7000 13120
rect 7120 13000 9880 13120
rect 10000 13000 10600 13120
rect 4676 12964 10600 13000
rect 0 12960 10600 12964
rect 0 12916 10600 12920
rect 0 12880 5924 12916
rect 0 12760 120 12880
rect 240 12760 3960 12880
rect 4080 12760 5924 12880
rect 0 12724 5924 12760
rect 5956 12724 6084 12916
rect 6116 12880 10600 12916
rect 6116 12760 6520 12880
rect 6640 12760 10360 12880
rect 10480 12760 10600 12880
rect 6116 12724 10600 12760
rect 0 12720 10600 12724
rect 4240 12636 4440 12640
rect 4240 12604 4244 12636
rect 4276 12604 4404 12636
rect 4436 12604 4440 12636
rect 4240 12600 4440 12604
rect 4480 12636 4680 12640
rect 4480 12604 4484 12636
rect 4516 12604 4644 12636
rect 4676 12604 4680 12636
rect 4480 12600 4680 12604
rect 4720 12636 5080 12640
rect 4720 12604 4724 12636
rect 4756 12604 4884 12636
rect 4916 12604 5044 12636
rect 5076 12604 5080 12636
rect 4720 12600 5080 12604
rect 5120 12636 5480 12640
rect 5120 12604 5124 12636
rect 5156 12604 5284 12636
rect 5316 12604 5444 12636
rect 5476 12604 5480 12636
rect 5120 12600 5480 12604
rect 5520 12636 5880 12640
rect 5520 12604 5524 12636
rect 5556 12604 5684 12636
rect 5716 12604 5844 12636
rect 5876 12604 5880 12636
rect 5520 12600 5880 12604
rect 5920 12636 6120 12640
rect 5920 12604 5924 12636
rect 5956 12604 6084 12636
rect 6116 12604 6120 12636
rect 5920 12600 6120 12604
rect 6160 12636 6360 12640
rect 6160 12604 6164 12636
rect 6196 12604 6324 12636
rect 6356 12604 6360 12636
rect 6160 12600 6360 12604
rect 4240 12556 4440 12560
rect 4240 12524 4244 12556
rect 4276 12524 4404 12556
rect 4436 12524 4440 12556
rect 4240 12520 4440 12524
rect 4480 12556 4680 12560
rect 4480 12524 4484 12556
rect 4516 12524 4644 12556
rect 4676 12524 4680 12556
rect 4480 12520 4680 12524
rect 4720 12556 5080 12560
rect 4720 12524 4724 12556
rect 4756 12524 4884 12556
rect 4916 12524 5044 12556
rect 5076 12524 5080 12556
rect 4720 12520 5080 12524
rect 5120 12556 5480 12560
rect 5120 12524 5124 12556
rect 5156 12524 5284 12556
rect 5316 12524 5444 12556
rect 5476 12524 5480 12556
rect 5120 12520 5480 12524
rect 5520 12556 5880 12560
rect 5520 12524 5524 12556
rect 5556 12524 5684 12556
rect 5716 12524 5844 12556
rect 5876 12524 5880 12556
rect 5520 12520 5880 12524
rect 5920 12556 6120 12560
rect 5920 12524 5924 12556
rect 5956 12524 6084 12556
rect 6116 12524 6120 12556
rect 5920 12520 6120 12524
rect 6160 12556 6360 12560
rect 6160 12524 6164 12556
rect 6196 12524 6324 12556
rect 6356 12524 6360 12556
rect 6160 12520 6360 12524
rect 4240 12476 4440 12480
rect 4240 12444 4244 12476
rect 4276 12444 4404 12476
rect 4436 12444 4440 12476
rect 4240 12440 4440 12444
rect 4480 12476 4680 12480
rect 4480 12444 4484 12476
rect 4516 12444 4644 12476
rect 4676 12444 4680 12476
rect 4480 12440 4680 12444
rect 4720 12476 5080 12480
rect 4720 12444 4724 12476
rect 4756 12444 4884 12476
rect 4916 12444 5044 12476
rect 5076 12444 5080 12476
rect 4720 12440 5080 12444
rect 5120 12476 5480 12480
rect 5120 12444 5124 12476
rect 5156 12444 5284 12476
rect 5316 12444 5444 12476
rect 5476 12444 5480 12476
rect 5120 12440 5480 12444
rect 5520 12476 5880 12480
rect 5520 12444 5524 12476
rect 5556 12444 5684 12476
rect 5716 12444 5844 12476
rect 5876 12444 5880 12476
rect 5520 12440 5880 12444
rect 5920 12476 6120 12480
rect 5920 12444 5924 12476
rect 5956 12444 6084 12476
rect 6116 12444 6120 12476
rect 5920 12440 6120 12444
rect 6160 12476 6360 12480
rect 6160 12444 6164 12476
rect 6196 12444 6324 12476
rect 6356 12444 6360 12476
rect 6160 12440 6360 12444
rect 4240 12396 4440 12400
rect 4240 12364 4244 12396
rect 4276 12364 4404 12396
rect 4436 12364 4440 12396
rect 4240 12360 4440 12364
rect 4480 12396 4680 12400
rect 4480 12364 4484 12396
rect 4516 12364 4644 12396
rect 4676 12364 4680 12396
rect 4480 12360 4680 12364
rect 4720 12396 5080 12400
rect 4720 12364 4724 12396
rect 4756 12364 4884 12396
rect 4916 12364 5044 12396
rect 5076 12364 5080 12396
rect 4720 12360 5080 12364
rect 5120 12396 5480 12400
rect 5120 12364 5124 12396
rect 5156 12364 5284 12396
rect 5316 12364 5444 12396
rect 5476 12364 5480 12396
rect 5120 12360 5480 12364
rect 5520 12396 5880 12400
rect 5520 12364 5524 12396
rect 5556 12364 5684 12396
rect 5716 12364 5844 12396
rect 5876 12364 5880 12396
rect 5520 12360 5880 12364
rect 5920 12396 6120 12400
rect 5920 12364 5924 12396
rect 5956 12364 6084 12396
rect 6116 12364 6120 12396
rect 5920 12360 6120 12364
rect 6160 12396 6360 12400
rect 6160 12364 6164 12396
rect 6196 12364 6324 12396
rect 6356 12364 6360 12396
rect 6160 12360 6360 12364
rect 4240 12316 4440 12320
rect 4240 12284 4244 12316
rect 4276 12284 4404 12316
rect 4436 12284 4440 12316
rect 4240 12280 4440 12284
rect 4480 12316 4680 12320
rect 4480 12284 4484 12316
rect 4516 12284 4644 12316
rect 4676 12284 4680 12316
rect 4480 12280 4680 12284
rect 4720 12316 5080 12320
rect 4720 12284 4724 12316
rect 4756 12284 4884 12316
rect 4916 12284 5044 12316
rect 5076 12284 5080 12316
rect 4720 12280 5080 12284
rect 5120 12316 5480 12320
rect 5120 12284 5124 12316
rect 5156 12284 5284 12316
rect 5316 12284 5444 12316
rect 5476 12284 5480 12316
rect 5120 12280 5480 12284
rect 5520 12316 5880 12320
rect 5520 12284 5524 12316
rect 5556 12284 5684 12316
rect 5716 12284 5844 12316
rect 5876 12284 5880 12316
rect 5520 12280 5880 12284
rect 5920 12316 6120 12320
rect 5920 12284 5924 12316
rect 5956 12284 6084 12316
rect 6116 12284 6120 12316
rect 5920 12280 6120 12284
rect 6160 12316 6360 12320
rect 6160 12284 6164 12316
rect 6196 12284 6324 12316
rect 6356 12284 6360 12316
rect 6160 12280 6360 12284
rect 4240 12236 4440 12240
rect 4240 12204 4244 12236
rect 4276 12204 4404 12236
rect 4436 12204 4440 12236
rect 4240 12200 4440 12204
rect 4480 12236 4680 12240
rect 4480 12204 4484 12236
rect 4516 12204 4644 12236
rect 4676 12204 4680 12236
rect 4480 12200 4680 12204
rect 4720 12236 5080 12240
rect 4720 12204 4724 12236
rect 4756 12204 4884 12236
rect 4916 12204 5044 12236
rect 5076 12204 5080 12236
rect 4720 12200 5080 12204
rect 5120 12236 5480 12240
rect 5120 12204 5124 12236
rect 5156 12204 5284 12236
rect 5316 12204 5444 12236
rect 5476 12204 5480 12236
rect 5120 12200 5480 12204
rect 5520 12236 5880 12240
rect 5520 12204 5524 12236
rect 5556 12204 5684 12236
rect 5716 12204 5844 12236
rect 5876 12204 5880 12236
rect 5520 12200 5880 12204
rect 5920 12236 6120 12240
rect 5920 12204 5924 12236
rect 5956 12204 6084 12236
rect 6116 12204 6120 12236
rect 5920 12200 6120 12204
rect 6160 12236 6360 12240
rect 6160 12204 6164 12236
rect 6196 12204 6324 12236
rect 6356 12204 6360 12236
rect 6160 12200 6360 12204
rect 4240 12156 4440 12160
rect 4240 12124 4244 12156
rect 4276 12124 4404 12156
rect 4436 12124 4440 12156
rect 4240 12120 4440 12124
rect 4480 12156 4680 12160
rect 4480 12124 4484 12156
rect 4516 12124 4644 12156
rect 4676 12124 4680 12156
rect 4480 12120 4680 12124
rect 4720 12156 5080 12160
rect 4720 12124 4724 12156
rect 4756 12124 4884 12156
rect 4916 12124 5044 12156
rect 5076 12124 5080 12156
rect 4720 12120 5080 12124
rect 5120 12156 5480 12160
rect 5120 12124 5124 12156
rect 5156 12124 5284 12156
rect 5316 12124 5444 12156
rect 5476 12124 5480 12156
rect 5120 12120 5480 12124
rect 5520 12156 5880 12160
rect 5520 12124 5524 12156
rect 5556 12124 5684 12156
rect 5716 12124 5844 12156
rect 5876 12124 5880 12156
rect 5520 12120 5880 12124
rect 5920 12156 6120 12160
rect 5920 12124 5924 12156
rect 5956 12124 6084 12156
rect 6116 12124 6120 12156
rect 5920 12120 6120 12124
rect 6160 12156 6360 12160
rect 6160 12124 6164 12156
rect 6196 12124 6324 12156
rect 6356 12124 6360 12156
rect 6160 12120 6360 12124
rect 4240 11836 4440 11840
rect 4240 11804 4244 11836
rect 4276 11804 4404 11836
rect 4436 11804 4440 11836
rect 4240 11800 4440 11804
rect 4480 11836 4680 11840
rect 4480 11804 4484 11836
rect 4516 11804 4644 11836
rect 4676 11804 4680 11836
rect 4480 11800 4680 11804
rect 4720 11836 5080 11840
rect 4720 11804 4724 11836
rect 4756 11804 4884 11836
rect 4916 11804 5044 11836
rect 5076 11804 5080 11836
rect 4720 11800 5080 11804
rect 5120 11836 5480 11840
rect 5120 11804 5124 11836
rect 5156 11804 5284 11836
rect 5316 11804 5444 11836
rect 5476 11804 5480 11836
rect 5120 11800 5480 11804
rect 5520 11836 5880 11840
rect 5520 11804 5524 11836
rect 5556 11804 5684 11836
rect 5716 11804 5844 11836
rect 5876 11804 5880 11836
rect 5520 11800 5880 11804
rect 5920 11836 6120 11840
rect 5920 11804 5924 11836
rect 5956 11804 6084 11836
rect 6116 11804 6120 11836
rect 5920 11800 6120 11804
rect 6160 11836 6360 11840
rect 6160 11804 6164 11836
rect 6196 11804 6324 11836
rect 6356 11804 6360 11836
rect 6160 11800 6360 11804
rect 4240 11756 4440 11760
rect 4240 11724 4244 11756
rect 4276 11724 4404 11756
rect 4436 11724 4440 11756
rect 4240 11720 4440 11724
rect 4480 11756 4680 11760
rect 4480 11724 4484 11756
rect 4516 11724 4644 11756
rect 4676 11724 4680 11756
rect 4480 11720 4680 11724
rect 4720 11756 5080 11760
rect 4720 11724 4724 11756
rect 4756 11724 4884 11756
rect 4916 11724 5044 11756
rect 5076 11724 5080 11756
rect 4720 11720 5080 11724
rect 5120 11756 5480 11760
rect 5120 11724 5124 11756
rect 5156 11724 5284 11756
rect 5316 11724 5444 11756
rect 5476 11724 5480 11756
rect 5120 11720 5480 11724
rect 5520 11756 5880 11760
rect 5520 11724 5524 11756
rect 5556 11724 5684 11756
rect 5716 11724 5844 11756
rect 5876 11724 5880 11756
rect 5520 11720 5880 11724
rect 5920 11756 6120 11760
rect 5920 11724 5924 11756
rect 5956 11724 6084 11756
rect 6116 11724 6120 11756
rect 5920 11720 6120 11724
rect 6160 11756 6360 11760
rect 6160 11724 6164 11756
rect 6196 11724 6324 11756
rect 6356 11724 6360 11756
rect 6160 11720 6360 11724
rect 4240 11676 4440 11680
rect 4240 11644 4244 11676
rect 4276 11644 4404 11676
rect 4436 11644 4440 11676
rect 4240 11640 4440 11644
rect 4480 11676 4680 11680
rect 4480 11644 4484 11676
rect 4516 11644 4644 11676
rect 4676 11644 4680 11676
rect 4480 11640 4680 11644
rect 4720 11676 5080 11680
rect 4720 11644 4724 11676
rect 4756 11644 4884 11676
rect 4916 11644 5044 11676
rect 5076 11644 5080 11676
rect 4720 11640 5080 11644
rect 5120 11676 5480 11680
rect 5120 11644 5124 11676
rect 5156 11644 5284 11676
rect 5316 11644 5444 11676
rect 5476 11644 5480 11676
rect 5120 11640 5480 11644
rect 5520 11676 5880 11680
rect 5520 11644 5524 11676
rect 5556 11644 5684 11676
rect 5716 11644 5844 11676
rect 5876 11644 5880 11676
rect 5520 11640 5880 11644
rect 5920 11676 6120 11680
rect 5920 11644 5924 11676
rect 5956 11644 6084 11676
rect 6116 11644 6120 11676
rect 5920 11640 6120 11644
rect 6160 11676 6360 11680
rect 6160 11644 6164 11676
rect 6196 11644 6324 11676
rect 6356 11644 6360 11676
rect 6160 11640 6360 11644
rect 4240 11596 4440 11600
rect 4240 11564 4244 11596
rect 4276 11564 4404 11596
rect 4436 11564 4440 11596
rect 4240 11560 4440 11564
rect 4480 11596 4680 11600
rect 4480 11564 4484 11596
rect 4516 11564 4644 11596
rect 4676 11564 4680 11596
rect 4480 11560 4680 11564
rect 4720 11596 5080 11600
rect 4720 11564 4724 11596
rect 4756 11564 4884 11596
rect 4916 11564 5044 11596
rect 5076 11564 5080 11596
rect 4720 11560 5080 11564
rect 5120 11596 5480 11600
rect 5120 11564 5124 11596
rect 5156 11564 5284 11596
rect 5316 11564 5444 11596
rect 5476 11564 5480 11596
rect 5120 11560 5480 11564
rect 5520 11596 5880 11600
rect 5520 11564 5524 11596
rect 5556 11564 5684 11596
rect 5716 11564 5844 11596
rect 5876 11564 5880 11596
rect 5520 11560 5880 11564
rect 5920 11596 6120 11600
rect 5920 11564 5924 11596
rect 5956 11564 6084 11596
rect 6116 11564 6120 11596
rect 5920 11560 6120 11564
rect 6160 11596 6360 11600
rect 6160 11564 6164 11596
rect 6196 11564 6324 11596
rect 6356 11564 6360 11596
rect 6160 11560 6360 11564
rect 4240 11516 4440 11520
rect 4240 11484 4244 11516
rect 4276 11484 4404 11516
rect 4436 11484 4440 11516
rect 4240 11480 4440 11484
rect 4480 11516 4680 11520
rect 4480 11484 4484 11516
rect 4516 11484 4644 11516
rect 4676 11484 4680 11516
rect 4480 11480 4680 11484
rect 4720 11516 5080 11520
rect 4720 11484 4724 11516
rect 4756 11484 4884 11516
rect 4916 11484 5044 11516
rect 5076 11484 5080 11516
rect 4720 11480 5080 11484
rect 5120 11516 5480 11520
rect 5120 11484 5124 11516
rect 5156 11484 5284 11516
rect 5316 11484 5444 11516
rect 5476 11484 5480 11516
rect 5120 11480 5480 11484
rect 5520 11516 5880 11520
rect 5520 11484 5524 11516
rect 5556 11484 5684 11516
rect 5716 11484 5844 11516
rect 5876 11484 5880 11516
rect 5520 11480 5880 11484
rect 5920 11516 6120 11520
rect 5920 11484 5924 11516
rect 5956 11484 6084 11516
rect 6116 11484 6120 11516
rect 5920 11480 6120 11484
rect 6160 11516 6360 11520
rect 6160 11484 6164 11516
rect 6196 11484 6324 11516
rect 6356 11484 6360 11516
rect 6160 11480 6360 11484
rect 4240 11436 4440 11440
rect 4240 11404 4244 11436
rect 4276 11404 4404 11436
rect 4436 11404 4440 11436
rect 4240 11400 4440 11404
rect 4480 11436 4680 11440
rect 4480 11404 4484 11436
rect 4516 11404 4644 11436
rect 4676 11404 4680 11436
rect 4480 11400 4680 11404
rect 4720 11436 5080 11440
rect 4720 11404 4724 11436
rect 4756 11404 4884 11436
rect 4916 11404 5044 11436
rect 5076 11404 5080 11436
rect 4720 11400 5080 11404
rect 5120 11436 5480 11440
rect 5120 11404 5124 11436
rect 5156 11404 5284 11436
rect 5316 11404 5444 11436
rect 5476 11404 5480 11436
rect 5120 11400 5480 11404
rect 5520 11436 5880 11440
rect 5520 11404 5524 11436
rect 5556 11404 5684 11436
rect 5716 11404 5844 11436
rect 5876 11404 5880 11436
rect 5520 11400 5880 11404
rect 5920 11436 6120 11440
rect 5920 11404 5924 11436
rect 5956 11404 6084 11436
rect 6116 11404 6120 11436
rect 5920 11400 6120 11404
rect 6160 11436 6360 11440
rect 6160 11404 6164 11436
rect 6196 11404 6324 11436
rect 6356 11404 6360 11436
rect 6160 11400 6360 11404
rect 4240 10876 4440 10880
rect 4240 10844 4244 10876
rect 4276 10844 4404 10876
rect 4436 10844 4440 10876
rect 4240 10840 4440 10844
rect 4480 10876 4680 10880
rect 4480 10844 4484 10876
rect 4516 10844 4644 10876
rect 4676 10844 4680 10876
rect 4480 10840 4680 10844
rect 4720 10876 5080 10880
rect 4720 10844 4724 10876
rect 4756 10844 4884 10876
rect 4916 10844 5044 10876
rect 5076 10844 5080 10876
rect 4720 10840 5080 10844
rect 5120 10876 5480 10880
rect 5120 10844 5124 10876
rect 5156 10844 5284 10876
rect 5316 10844 5444 10876
rect 5476 10844 5480 10876
rect 5120 10840 5480 10844
rect 5520 10876 5880 10880
rect 5520 10844 5524 10876
rect 5556 10844 5684 10876
rect 5716 10844 5844 10876
rect 5876 10844 5880 10876
rect 5520 10840 5880 10844
rect 5920 10876 6120 10880
rect 5920 10844 5924 10876
rect 5956 10844 6084 10876
rect 6116 10844 6120 10876
rect 5920 10840 6120 10844
rect 6160 10876 6360 10880
rect 6160 10844 6164 10876
rect 6196 10844 6324 10876
rect 6356 10844 6360 10876
rect 6160 10840 6360 10844
rect 4240 10796 4440 10800
rect 4240 10764 4244 10796
rect 4276 10764 4404 10796
rect 4436 10764 4440 10796
rect 4240 10760 4440 10764
rect 4480 10796 4680 10800
rect 4480 10764 4484 10796
rect 4516 10764 4644 10796
rect 4676 10764 4680 10796
rect 4480 10760 4680 10764
rect 4720 10796 5080 10800
rect 4720 10764 4724 10796
rect 4756 10764 4884 10796
rect 4916 10764 5044 10796
rect 5076 10764 5080 10796
rect 4720 10760 5080 10764
rect 5120 10796 5480 10800
rect 5120 10764 5124 10796
rect 5156 10764 5284 10796
rect 5316 10764 5444 10796
rect 5476 10764 5480 10796
rect 5120 10760 5480 10764
rect 5520 10796 5880 10800
rect 5520 10764 5524 10796
rect 5556 10764 5684 10796
rect 5716 10764 5844 10796
rect 5876 10764 5880 10796
rect 5520 10760 5880 10764
rect 5920 10796 6120 10800
rect 5920 10764 5924 10796
rect 5956 10764 6084 10796
rect 6116 10764 6120 10796
rect 5920 10760 6120 10764
rect 6160 10796 6360 10800
rect 6160 10764 6164 10796
rect 6196 10764 6324 10796
rect 6356 10764 6360 10796
rect 6160 10760 6360 10764
rect 4240 10716 4440 10720
rect 4240 10684 4244 10716
rect 4276 10684 4404 10716
rect 4436 10684 4440 10716
rect 4240 10680 4440 10684
rect 4480 10716 4680 10720
rect 4480 10684 4484 10716
rect 4516 10684 4644 10716
rect 4676 10684 4680 10716
rect 4480 10680 4680 10684
rect 4720 10716 5080 10720
rect 4720 10684 4724 10716
rect 4756 10684 4884 10716
rect 4916 10684 5044 10716
rect 5076 10684 5080 10716
rect 4720 10680 5080 10684
rect 5120 10716 5480 10720
rect 5120 10684 5124 10716
rect 5156 10684 5284 10716
rect 5316 10684 5444 10716
rect 5476 10684 5480 10716
rect 5120 10680 5480 10684
rect 5520 10716 5880 10720
rect 5520 10684 5524 10716
rect 5556 10684 5684 10716
rect 5716 10684 5844 10716
rect 5876 10684 5880 10716
rect 5520 10680 5880 10684
rect 5920 10716 6120 10720
rect 5920 10684 5924 10716
rect 5956 10684 6084 10716
rect 6116 10684 6120 10716
rect 5920 10680 6120 10684
rect 6160 10716 6360 10720
rect 6160 10684 6164 10716
rect 6196 10684 6324 10716
rect 6356 10684 6360 10716
rect 6160 10680 6360 10684
rect 4240 10636 4440 10640
rect 4240 10604 4244 10636
rect 4276 10604 4404 10636
rect 4436 10604 4440 10636
rect 4240 10600 4440 10604
rect 4480 10636 4680 10640
rect 4480 10604 4484 10636
rect 4516 10604 4644 10636
rect 4676 10604 4680 10636
rect 4480 10600 4680 10604
rect 4720 10636 5080 10640
rect 4720 10604 4724 10636
rect 4756 10604 4884 10636
rect 4916 10604 5044 10636
rect 5076 10604 5080 10636
rect 4720 10600 5080 10604
rect 5120 10636 5480 10640
rect 5120 10604 5124 10636
rect 5156 10604 5284 10636
rect 5316 10604 5444 10636
rect 5476 10604 5480 10636
rect 5120 10600 5480 10604
rect 5520 10636 5880 10640
rect 5520 10604 5524 10636
rect 5556 10604 5684 10636
rect 5716 10604 5844 10636
rect 5876 10604 5880 10636
rect 5520 10600 5880 10604
rect 5920 10636 6120 10640
rect 5920 10604 5924 10636
rect 5956 10604 6084 10636
rect 6116 10604 6120 10636
rect 5920 10600 6120 10604
rect 6160 10636 6360 10640
rect 6160 10604 6164 10636
rect 6196 10604 6324 10636
rect 6356 10604 6360 10636
rect 6160 10600 6360 10604
rect 4240 10556 4440 10560
rect 4240 10524 4244 10556
rect 4276 10524 4404 10556
rect 4436 10524 4440 10556
rect 4240 10520 4440 10524
rect 4480 10556 4680 10560
rect 4480 10524 4484 10556
rect 4516 10524 4644 10556
rect 4676 10524 4680 10556
rect 4480 10520 4680 10524
rect 4720 10556 5080 10560
rect 4720 10524 4724 10556
rect 4756 10524 4884 10556
rect 4916 10524 5044 10556
rect 5076 10524 5080 10556
rect 4720 10520 5080 10524
rect 5120 10556 5480 10560
rect 5120 10524 5124 10556
rect 5156 10524 5284 10556
rect 5316 10524 5444 10556
rect 5476 10524 5480 10556
rect 5120 10520 5480 10524
rect 5520 10556 5880 10560
rect 5520 10524 5524 10556
rect 5556 10524 5684 10556
rect 5716 10524 5844 10556
rect 5876 10524 5880 10556
rect 5520 10520 5880 10524
rect 5920 10556 6120 10560
rect 5920 10524 5924 10556
rect 5956 10524 6084 10556
rect 6116 10524 6120 10556
rect 5920 10520 6120 10524
rect 6160 10556 6360 10560
rect 6160 10524 6164 10556
rect 6196 10524 6324 10556
rect 6356 10524 6360 10556
rect 6160 10520 6360 10524
rect 4240 10476 4440 10480
rect 4240 10444 4244 10476
rect 4276 10444 4404 10476
rect 4436 10444 4440 10476
rect 4240 10440 4440 10444
rect 4480 10476 4680 10480
rect 4480 10444 4484 10476
rect 4516 10444 4644 10476
rect 4676 10444 4680 10476
rect 4480 10440 4680 10444
rect 4720 10476 5080 10480
rect 4720 10444 4724 10476
rect 4756 10444 4884 10476
rect 4916 10444 5044 10476
rect 5076 10444 5080 10476
rect 4720 10440 5080 10444
rect 5120 10476 5480 10480
rect 5120 10444 5124 10476
rect 5156 10444 5284 10476
rect 5316 10444 5444 10476
rect 5476 10444 5480 10476
rect 5120 10440 5480 10444
rect 5520 10476 5880 10480
rect 5520 10444 5524 10476
rect 5556 10444 5684 10476
rect 5716 10444 5844 10476
rect 5876 10444 5880 10476
rect 5520 10440 5880 10444
rect 5920 10476 6120 10480
rect 5920 10444 5924 10476
rect 5956 10444 6084 10476
rect 6116 10444 6120 10476
rect 5920 10440 6120 10444
rect 6160 10476 6360 10480
rect 6160 10444 6164 10476
rect 6196 10444 6324 10476
rect 6356 10444 6360 10476
rect 6160 10440 6360 10444
rect 4240 10396 4440 10400
rect 4240 10364 4244 10396
rect 4276 10364 4404 10396
rect 4436 10364 4440 10396
rect 4240 10360 4440 10364
rect 4480 10396 4680 10400
rect 4480 10364 4484 10396
rect 4516 10364 4644 10396
rect 4676 10364 4680 10396
rect 4480 10360 4680 10364
rect 4720 10396 5080 10400
rect 4720 10364 4724 10396
rect 4756 10364 4884 10396
rect 4916 10364 5044 10396
rect 5076 10364 5080 10396
rect 4720 10360 5080 10364
rect 5120 10396 5480 10400
rect 5120 10364 5124 10396
rect 5156 10364 5284 10396
rect 5316 10364 5444 10396
rect 5476 10364 5480 10396
rect 5120 10360 5480 10364
rect 5520 10396 5880 10400
rect 5520 10364 5524 10396
rect 5556 10364 5684 10396
rect 5716 10364 5844 10396
rect 5876 10364 5880 10396
rect 5520 10360 5880 10364
rect 5920 10396 6120 10400
rect 5920 10364 5924 10396
rect 5956 10364 6084 10396
rect 6116 10364 6120 10396
rect 5920 10360 6120 10364
rect 6160 10396 6360 10400
rect 6160 10364 6164 10396
rect 6196 10364 6324 10396
rect 6356 10364 6360 10396
rect 6160 10360 6360 10364
rect 4240 10316 4440 10320
rect 4240 10284 4244 10316
rect 4276 10284 4404 10316
rect 4436 10284 4440 10316
rect 4240 10280 4440 10284
rect 4480 10316 4680 10320
rect 4480 10284 4484 10316
rect 4516 10284 4644 10316
rect 4676 10284 4680 10316
rect 4480 10280 4680 10284
rect 4720 10316 5080 10320
rect 4720 10284 4724 10316
rect 4756 10284 4884 10316
rect 4916 10284 5044 10316
rect 5076 10284 5080 10316
rect 4720 10280 5080 10284
rect 5120 10316 5480 10320
rect 5120 10284 5124 10316
rect 5156 10284 5284 10316
rect 5316 10284 5444 10316
rect 5476 10284 5480 10316
rect 5120 10280 5480 10284
rect 5520 10316 5880 10320
rect 5520 10284 5524 10316
rect 5556 10284 5684 10316
rect 5716 10284 5844 10316
rect 5876 10284 5880 10316
rect 5520 10280 5880 10284
rect 5920 10316 6120 10320
rect 5920 10284 5924 10316
rect 5956 10284 6084 10316
rect 6116 10284 6120 10316
rect 5920 10280 6120 10284
rect 6160 10316 6360 10320
rect 6160 10284 6164 10316
rect 6196 10284 6324 10316
rect 6356 10284 6360 10316
rect 6160 10280 6360 10284
rect 4240 10236 4440 10240
rect 4240 10204 4244 10236
rect 4276 10204 4404 10236
rect 4436 10204 4440 10236
rect 4240 10200 4440 10204
rect 4480 10236 4680 10240
rect 4480 10204 4484 10236
rect 4516 10204 4644 10236
rect 4676 10204 4680 10236
rect 4480 10200 4680 10204
rect 4720 10236 5080 10240
rect 4720 10204 4724 10236
rect 4756 10204 4884 10236
rect 4916 10204 5044 10236
rect 5076 10204 5080 10236
rect 4720 10200 5080 10204
rect 5120 10236 5480 10240
rect 5120 10204 5124 10236
rect 5156 10204 5284 10236
rect 5316 10204 5444 10236
rect 5476 10204 5480 10236
rect 5120 10200 5480 10204
rect 5520 10236 5880 10240
rect 5520 10204 5524 10236
rect 5556 10204 5684 10236
rect 5716 10204 5844 10236
rect 5876 10204 5880 10236
rect 5520 10200 5880 10204
rect 5920 10236 6120 10240
rect 5920 10204 5924 10236
rect 5956 10204 6084 10236
rect 6116 10204 6120 10236
rect 5920 10200 6120 10204
rect 6160 10236 6360 10240
rect 6160 10204 6164 10236
rect 6196 10204 6324 10236
rect 6356 10204 6360 10236
rect 6160 10200 6360 10204
rect 4240 10156 4440 10160
rect 4240 10124 4244 10156
rect 4276 10124 4404 10156
rect 4436 10124 4440 10156
rect 4240 10120 4440 10124
rect 4480 10156 4680 10160
rect 4480 10124 4484 10156
rect 4516 10124 4644 10156
rect 4676 10124 4680 10156
rect 4480 10120 4680 10124
rect 4720 10156 5080 10160
rect 4720 10124 4724 10156
rect 4756 10124 4884 10156
rect 4916 10124 5044 10156
rect 5076 10124 5080 10156
rect 4720 10120 5080 10124
rect 5120 10156 5480 10160
rect 5120 10124 5124 10156
rect 5156 10124 5284 10156
rect 5316 10124 5444 10156
rect 5476 10124 5480 10156
rect 5120 10120 5480 10124
rect 5520 10156 5880 10160
rect 5520 10124 5524 10156
rect 5556 10124 5684 10156
rect 5716 10124 5844 10156
rect 5876 10124 5880 10156
rect 5520 10120 5880 10124
rect 5920 10156 6120 10160
rect 5920 10124 5924 10156
rect 5956 10124 6084 10156
rect 6116 10124 6120 10156
rect 5920 10120 6120 10124
rect 6160 10156 6360 10160
rect 6160 10124 6164 10156
rect 6196 10124 6324 10156
rect 6356 10124 6360 10156
rect 6160 10120 6360 10124
rect 4240 10076 4440 10080
rect 4240 10044 4244 10076
rect 4276 10044 4404 10076
rect 4436 10044 4440 10076
rect 4240 10040 4440 10044
rect 4480 10076 4680 10080
rect 4480 10044 4484 10076
rect 4516 10044 4644 10076
rect 4676 10044 4680 10076
rect 4480 10040 4680 10044
rect 4720 10076 5080 10080
rect 4720 10044 4724 10076
rect 4756 10044 4884 10076
rect 4916 10044 5044 10076
rect 5076 10044 5080 10076
rect 4720 10040 5080 10044
rect 5120 10076 5480 10080
rect 5120 10044 5124 10076
rect 5156 10044 5284 10076
rect 5316 10044 5444 10076
rect 5476 10044 5480 10076
rect 5120 10040 5480 10044
rect 5520 10076 5880 10080
rect 5520 10044 5524 10076
rect 5556 10044 5684 10076
rect 5716 10044 5844 10076
rect 5876 10044 5880 10076
rect 5520 10040 5880 10044
rect 5920 10076 6120 10080
rect 5920 10044 5924 10076
rect 5956 10044 6084 10076
rect 6116 10044 6120 10076
rect 5920 10040 6120 10044
rect 6160 10076 6360 10080
rect 6160 10044 6164 10076
rect 6196 10044 6324 10076
rect 6356 10044 6360 10076
rect 6160 10040 6360 10044
rect 4240 9996 4440 10000
rect 4240 9964 4244 9996
rect 4276 9964 4404 9996
rect 4436 9964 4440 9996
rect 4240 9960 4440 9964
rect 4480 9996 4680 10000
rect 4480 9964 4484 9996
rect 4516 9964 4644 9996
rect 4676 9964 4680 9996
rect 4480 9960 4680 9964
rect 4720 9996 5080 10000
rect 4720 9964 4724 9996
rect 4756 9964 4884 9996
rect 4916 9964 5044 9996
rect 5076 9964 5080 9996
rect 4720 9960 5080 9964
rect 5120 9996 5480 10000
rect 5120 9964 5124 9996
rect 5156 9964 5284 9996
rect 5316 9964 5444 9996
rect 5476 9964 5480 9996
rect 5120 9960 5480 9964
rect 5520 9996 5880 10000
rect 5520 9964 5524 9996
rect 5556 9964 5684 9996
rect 5716 9964 5844 9996
rect 5876 9964 5880 9996
rect 5520 9960 5880 9964
rect 5920 9996 6120 10000
rect 5920 9964 5924 9996
rect 5956 9964 6084 9996
rect 6116 9964 6120 9996
rect 5920 9960 6120 9964
rect 6160 9996 6360 10000
rect 6160 9964 6164 9996
rect 6196 9964 6324 9996
rect 6356 9964 6360 9996
rect 6160 9960 6360 9964
rect 4240 9916 4440 9920
rect 4240 9884 4244 9916
rect 4276 9884 4404 9916
rect 4436 9884 4440 9916
rect 4240 9880 4440 9884
rect 4480 9916 4680 9920
rect 4480 9884 4484 9916
rect 4516 9884 4644 9916
rect 4676 9884 4680 9916
rect 4480 9880 4680 9884
rect 4720 9916 5080 9920
rect 4720 9884 4724 9916
rect 4756 9884 4884 9916
rect 4916 9884 5044 9916
rect 5076 9884 5080 9916
rect 4720 9880 5080 9884
rect 5120 9916 5480 9920
rect 5120 9884 5124 9916
rect 5156 9884 5284 9916
rect 5316 9884 5444 9916
rect 5476 9884 5480 9916
rect 5120 9880 5480 9884
rect 5520 9916 5880 9920
rect 5520 9884 5524 9916
rect 5556 9884 5684 9916
rect 5716 9884 5844 9916
rect 5876 9884 5880 9916
rect 5520 9880 5880 9884
rect 5920 9916 6120 9920
rect 5920 9884 5924 9916
rect 5956 9884 6084 9916
rect 6116 9884 6120 9916
rect 5920 9880 6120 9884
rect 6160 9916 6360 9920
rect 6160 9884 6164 9916
rect 6196 9884 6324 9916
rect 6356 9884 6360 9916
rect 6160 9880 6360 9884
rect 4240 9836 4440 9840
rect 4240 9804 4244 9836
rect 4276 9804 4404 9836
rect 4436 9804 4440 9836
rect 4240 9800 4440 9804
rect 4480 9836 4680 9840
rect 4480 9804 4484 9836
rect 4516 9804 4644 9836
rect 4676 9804 4680 9836
rect 4480 9800 4680 9804
rect 4720 9836 5080 9840
rect 4720 9804 4724 9836
rect 4756 9804 4884 9836
rect 4916 9804 5044 9836
rect 5076 9804 5080 9836
rect 4720 9800 5080 9804
rect 5120 9836 5480 9840
rect 5120 9804 5124 9836
rect 5156 9804 5284 9836
rect 5316 9804 5444 9836
rect 5476 9804 5480 9836
rect 5120 9800 5480 9804
rect 5520 9836 5880 9840
rect 5520 9804 5524 9836
rect 5556 9804 5684 9836
rect 5716 9804 5844 9836
rect 5876 9804 5880 9836
rect 5520 9800 5880 9804
rect 5920 9836 6120 9840
rect 5920 9804 5924 9836
rect 5956 9804 6084 9836
rect 6116 9804 6120 9836
rect 5920 9800 6120 9804
rect 6160 9836 6360 9840
rect 6160 9804 6164 9836
rect 6196 9804 6324 9836
rect 6356 9804 6360 9836
rect 6160 9800 6360 9804
rect 4240 9756 4440 9760
rect 4240 9724 4244 9756
rect 4276 9724 4404 9756
rect 4436 9724 4440 9756
rect 4240 9720 4440 9724
rect 4480 9756 4680 9760
rect 4480 9724 4484 9756
rect 4516 9724 4644 9756
rect 4676 9724 4680 9756
rect 4480 9720 4680 9724
rect 4720 9756 5080 9760
rect 4720 9724 4724 9756
rect 4756 9724 4884 9756
rect 4916 9724 5044 9756
rect 5076 9724 5080 9756
rect 4720 9720 5080 9724
rect 5120 9756 5480 9760
rect 5120 9724 5124 9756
rect 5156 9724 5284 9756
rect 5316 9724 5444 9756
rect 5476 9724 5480 9756
rect 5120 9720 5480 9724
rect 5520 9756 5880 9760
rect 5520 9724 5524 9756
rect 5556 9724 5684 9756
rect 5716 9724 5844 9756
rect 5876 9724 5880 9756
rect 5520 9720 5880 9724
rect 5920 9756 6120 9760
rect 5920 9724 5924 9756
rect 5956 9724 6084 9756
rect 6116 9724 6120 9756
rect 5920 9720 6120 9724
rect 6160 9756 6360 9760
rect 6160 9724 6164 9756
rect 6196 9724 6324 9756
rect 6356 9724 6360 9756
rect 6160 9720 6360 9724
rect 4240 9356 4440 9360
rect 4240 9324 4244 9356
rect 4276 9324 4404 9356
rect 4436 9324 4440 9356
rect 4240 9320 4440 9324
rect 4480 9356 4680 9360
rect 4480 9324 4484 9356
rect 4516 9324 4644 9356
rect 4676 9324 4680 9356
rect 4480 9320 4680 9324
rect 4720 9356 5080 9360
rect 4720 9324 4724 9356
rect 4756 9324 4884 9356
rect 4916 9324 5044 9356
rect 5076 9324 5080 9356
rect 4720 9320 5080 9324
rect 5120 9356 5480 9360
rect 5120 9324 5124 9356
rect 5156 9324 5284 9356
rect 5316 9324 5444 9356
rect 5476 9324 5480 9356
rect 5120 9320 5480 9324
rect 5520 9356 5880 9360
rect 5520 9324 5524 9356
rect 5556 9324 5684 9356
rect 5716 9324 5844 9356
rect 5876 9324 5880 9356
rect 5520 9320 5880 9324
rect 5920 9356 6120 9360
rect 5920 9324 5924 9356
rect 5956 9324 6084 9356
rect 6116 9324 6120 9356
rect 5920 9320 6120 9324
rect 6160 9356 6360 9360
rect 6160 9324 6164 9356
rect 6196 9324 6324 9356
rect 6356 9324 6360 9356
rect 6160 9320 6360 9324
rect 4240 9276 4440 9280
rect 4240 9244 4244 9276
rect 4276 9244 4404 9276
rect 4436 9244 4440 9276
rect 4240 9240 4440 9244
rect 4480 9276 4680 9280
rect 4480 9244 4484 9276
rect 4516 9244 4644 9276
rect 4676 9244 4680 9276
rect 4480 9240 4680 9244
rect 4720 9276 5080 9280
rect 4720 9244 4724 9276
rect 4756 9244 4884 9276
rect 4916 9244 5044 9276
rect 5076 9244 5080 9276
rect 4720 9240 5080 9244
rect 5120 9276 5480 9280
rect 5120 9244 5124 9276
rect 5156 9244 5284 9276
rect 5316 9244 5444 9276
rect 5476 9244 5480 9276
rect 5120 9240 5480 9244
rect 5520 9276 5880 9280
rect 5520 9244 5524 9276
rect 5556 9244 5684 9276
rect 5716 9244 5844 9276
rect 5876 9244 5880 9276
rect 5520 9240 5880 9244
rect 5920 9276 6120 9280
rect 5920 9244 5924 9276
rect 5956 9244 6084 9276
rect 6116 9244 6120 9276
rect 5920 9240 6120 9244
rect 6160 9276 6360 9280
rect 6160 9244 6164 9276
rect 6196 9244 6324 9276
rect 6356 9244 6360 9276
rect 6160 9240 6360 9244
rect 4240 9196 4440 9200
rect 4240 9164 4244 9196
rect 4276 9164 4404 9196
rect 4436 9164 4440 9196
rect 4240 9160 4440 9164
rect 4480 9196 4680 9200
rect 4480 9164 4484 9196
rect 4516 9164 4644 9196
rect 4676 9164 4680 9196
rect 4480 9160 4680 9164
rect 4720 9196 5080 9200
rect 4720 9164 4724 9196
rect 4756 9164 4884 9196
rect 4916 9164 5044 9196
rect 5076 9164 5080 9196
rect 4720 9160 5080 9164
rect 5120 9196 5480 9200
rect 5120 9164 5124 9196
rect 5156 9164 5284 9196
rect 5316 9164 5444 9196
rect 5476 9164 5480 9196
rect 5120 9160 5480 9164
rect 5520 9196 5880 9200
rect 5520 9164 5524 9196
rect 5556 9164 5684 9196
rect 5716 9164 5844 9196
rect 5876 9164 5880 9196
rect 5520 9160 5880 9164
rect 5920 9196 6120 9200
rect 5920 9164 5924 9196
rect 5956 9164 6084 9196
rect 6116 9164 6120 9196
rect 5920 9160 6120 9164
rect 6160 9196 6360 9200
rect 6160 9164 6164 9196
rect 6196 9164 6324 9196
rect 6356 9164 6360 9196
rect 6160 9160 6360 9164
rect 4240 8876 4440 8880
rect 4240 8844 4244 8876
rect 4276 8844 4404 8876
rect 4436 8844 4440 8876
rect 4240 8840 4440 8844
rect 4480 8876 4680 8880
rect 4480 8844 4484 8876
rect 4516 8844 4644 8876
rect 4676 8844 4680 8876
rect 4480 8840 4680 8844
rect 4720 8876 5080 8880
rect 4720 8844 4724 8876
rect 4756 8844 4884 8876
rect 4916 8844 5044 8876
rect 5076 8844 5080 8876
rect 4720 8840 5080 8844
rect 5120 8876 5480 8880
rect 5120 8844 5124 8876
rect 5156 8844 5284 8876
rect 5316 8844 5444 8876
rect 5476 8844 5480 8876
rect 5120 8840 5480 8844
rect 5520 8876 5880 8880
rect 5520 8844 5524 8876
rect 5556 8844 5684 8876
rect 5716 8844 5844 8876
rect 5876 8844 5880 8876
rect 5520 8840 5880 8844
rect 5920 8876 6120 8880
rect 5920 8844 5924 8876
rect 5956 8844 6084 8876
rect 6116 8844 6120 8876
rect 5920 8840 6120 8844
rect 6160 8876 6360 8880
rect 6160 8844 6164 8876
rect 6196 8844 6324 8876
rect 6356 8844 6360 8876
rect 6160 8840 6360 8844
rect 4240 8796 4440 8800
rect 4240 8764 4244 8796
rect 4276 8764 4404 8796
rect 4436 8764 4440 8796
rect 4240 8760 4440 8764
rect 4480 8796 4680 8800
rect 4480 8764 4484 8796
rect 4516 8764 4644 8796
rect 4676 8764 4680 8796
rect 4480 8760 4680 8764
rect 4720 8796 5080 8800
rect 4720 8764 4724 8796
rect 4756 8764 4884 8796
rect 4916 8764 5044 8796
rect 5076 8764 5080 8796
rect 4720 8760 5080 8764
rect 5120 8796 5480 8800
rect 5120 8764 5124 8796
rect 5156 8764 5284 8796
rect 5316 8764 5444 8796
rect 5476 8764 5480 8796
rect 5120 8760 5480 8764
rect 5520 8796 5880 8800
rect 5520 8764 5524 8796
rect 5556 8764 5684 8796
rect 5716 8764 5844 8796
rect 5876 8764 5880 8796
rect 5520 8760 5880 8764
rect 5920 8796 6120 8800
rect 5920 8764 5924 8796
rect 5956 8764 6084 8796
rect 6116 8764 6120 8796
rect 5920 8760 6120 8764
rect 6160 8796 6360 8800
rect 6160 8764 6164 8796
rect 6196 8764 6324 8796
rect 6356 8764 6360 8796
rect 6160 8760 6360 8764
rect 4240 8716 4440 8720
rect 4240 8684 4244 8716
rect 4276 8684 4404 8716
rect 4436 8684 4440 8716
rect 4240 8680 4440 8684
rect 4480 8716 4680 8720
rect 4480 8684 4484 8716
rect 4516 8684 4644 8716
rect 4676 8684 4680 8716
rect 4480 8680 4680 8684
rect 4720 8716 5080 8720
rect 4720 8684 4724 8716
rect 4756 8684 4884 8716
rect 4916 8684 5044 8716
rect 5076 8684 5080 8716
rect 4720 8680 5080 8684
rect 5120 8716 5480 8720
rect 5120 8684 5124 8716
rect 5156 8684 5284 8716
rect 5316 8684 5444 8716
rect 5476 8684 5480 8716
rect 5120 8680 5480 8684
rect 5520 8716 5880 8720
rect 5520 8684 5524 8716
rect 5556 8684 5684 8716
rect 5716 8684 5844 8716
rect 5876 8684 5880 8716
rect 5520 8680 5880 8684
rect 5920 8716 6120 8720
rect 5920 8684 5924 8716
rect 5956 8684 6084 8716
rect 6116 8684 6120 8716
rect 5920 8680 6120 8684
rect 6160 8716 6360 8720
rect 6160 8684 6164 8716
rect 6196 8684 6324 8716
rect 6356 8684 6360 8716
rect 6160 8680 6360 8684
rect 4240 8636 4440 8640
rect 4240 8604 4244 8636
rect 4276 8604 4404 8636
rect 4436 8604 4440 8636
rect 4240 8600 4440 8604
rect 4480 8636 4680 8640
rect 4480 8604 4484 8636
rect 4516 8604 4644 8636
rect 4676 8604 4680 8636
rect 4480 8600 4680 8604
rect 4720 8636 5080 8640
rect 4720 8604 4724 8636
rect 4756 8604 4884 8636
rect 4916 8604 5044 8636
rect 5076 8604 5080 8636
rect 4720 8600 5080 8604
rect 5120 8636 5480 8640
rect 5120 8604 5124 8636
rect 5156 8604 5284 8636
rect 5316 8604 5444 8636
rect 5476 8604 5480 8636
rect 5120 8600 5480 8604
rect 5520 8636 5880 8640
rect 5520 8604 5524 8636
rect 5556 8604 5684 8636
rect 5716 8604 5844 8636
rect 5876 8604 5880 8636
rect 5520 8600 5880 8604
rect 5920 8636 6120 8640
rect 5920 8604 5924 8636
rect 5956 8604 6084 8636
rect 6116 8604 6120 8636
rect 5920 8600 6120 8604
rect 6160 8636 6360 8640
rect 6160 8604 6164 8636
rect 6196 8604 6324 8636
rect 6356 8604 6360 8636
rect 6160 8600 6360 8604
rect 4240 8556 4440 8560
rect 4240 8524 4244 8556
rect 4276 8524 4404 8556
rect 4436 8524 4440 8556
rect 4240 8520 4440 8524
rect 4480 8556 4680 8560
rect 4480 8524 4484 8556
rect 4516 8524 4644 8556
rect 4676 8524 4680 8556
rect 4480 8520 4680 8524
rect 4720 8556 5080 8560
rect 4720 8524 4724 8556
rect 4756 8524 4884 8556
rect 4916 8524 5044 8556
rect 5076 8524 5080 8556
rect 4720 8520 5080 8524
rect 5120 8556 5480 8560
rect 5120 8524 5124 8556
rect 5156 8524 5284 8556
rect 5316 8524 5444 8556
rect 5476 8524 5480 8556
rect 5120 8520 5480 8524
rect 5520 8556 5880 8560
rect 5520 8524 5524 8556
rect 5556 8524 5684 8556
rect 5716 8524 5844 8556
rect 5876 8524 5880 8556
rect 5520 8520 5880 8524
rect 5920 8556 6120 8560
rect 5920 8524 5924 8556
rect 5956 8524 6084 8556
rect 6116 8524 6120 8556
rect 5920 8520 6120 8524
rect 6160 8556 6360 8560
rect 6160 8524 6164 8556
rect 6196 8524 6324 8556
rect 6356 8524 6360 8556
rect 6160 8520 6360 8524
rect 4240 7636 4440 7640
rect 4240 7604 4244 7636
rect 4276 7604 4404 7636
rect 4436 7604 4440 7636
rect 4240 7600 4440 7604
rect 4480 7636 4680 7640
rect 4480 7604 4484 7636
rect 4516 7604 4644 7636
rect 4676 7604 4680 7636
rect 4480 7600 4680 7604
rect 4720 7636 5080 7640
rect 4720 7604 4724 7636
rect 4756 7604 4884 7636
rect 4916 7604 5044 7636
rect 5076 7604 5080 7636
rect 4720 7600 5080 7604
rect 5120 7636 5480 7640
rect 5120 7604 5124 7636
rect 5156 7604 5284 7636
rect 5316 7604 5444 7636
rect 5476 7604 5480 7636
rect 5120 7600 5480 7604
rect 5520 7636 5880 7640
rect 5520 7604 5524 7636
rect 5556 7604 5684 7636
rect 5716 7604 5844 7636
rect 5876 7604 5880 7636
rect 5520 7600 5880 7604
rect 5920 7636 6120 7640
rect 5920 7604 5924 7636
rect 5956 7604 6084 7636
rect 6116 7604 6120 7636
rect 5920 7600 6120 7604
rect 6160 7636 6360 7640
rect 6160 7604 6164 7636
rect 6196 7604 6324 7636
rect 6356 7604 6360 7636
rect 6160 7600 6360 7604
rect 4240 7556 4440 7560
rect 4240 7524 4244 7556
rect 4276 7524 4404 7556
rect 4436 7524 4440 7556
rect 4240 7520 4440 7524
rect 4480 7556 4680 7560
rect 4480 7524 4484 7556
rect 4516 7524 4644 7556
rect 4676 7524 4680 7556
rect 4480 7520 4680 7524
rect 4720 7556 5080 7560
rect 4720 7524 4724 7556
rect 4756 7524 4884 7556
rect 4916 7524 5044 7556
rect 5076 7524 5080 7556
rect 4720 7520 5080 7524
rect 5120 7556 5480 7560
rect 5120 7524 5124 7556
rect 5156 7524 5284 7556
rect 5316 7524 5444 7556
rect 5476 7524 5480 7556
rect 5120 7520 5480 7524
rect 5520 7556 5880 7560
rect 5520 7524 5524 7556
rect 5556 7524 5684 7556
rect 5716 7524 5844 7556
rect 5876 7524 5880 7556
rect 5520 7520 5880 7524
rect 5920 7556 6120 7560
rect 5920 7524 5924 7556
rect 5956 7524 6084 7556
rect 6116 7524 6120 7556
rect 5920 7520 6120 7524
rect 6160 7556 6360 7560
rect 6160 7524 6164 7556
rect 6196 7524 6324 7556
rect 6356 7524 6360 7556
rect 6160 7520 6360 7524
rect 4240 7476 4440 7480
rect 4240 7444 4244 7476
rect 4276 7444 4404 7476
rect 4436 7444 4440 7476
rect 4240 7440 4440 7444
rect 4480 7476 4680 7480
rect 4480 7444 4484 7476
rect 4516 7444 4644 7476
rect 4676 7444 4680 7476
rect 4480 7440 4680 7444
rect 4720 7476 5080 7480
rect 4720 7444 4724 7476
rect 4756 7444 4884 7476
rect 4916 7444 5044 7476
rect 5076 7444 5080 7476
rect 4720 7440 5080 7444
rect 5120 7476 5480 7480
rect 5120 7444 5124 7476
rect 5156 7444 5284 7476
rect 5316 7444 5444 7476
rect 5476 7444 5480 7476
rect 5120 7440 5480 7444
rect 5520 7476 5880 7480
rect 5520 7444 5524 7476
rect 5556 7444 5684 7476
rect 5716 7444 5844 7476
rect 5876 7444 5880 7476
rect 5520 7440 5880 7444
rect 5920 7476 6120 7480
rect 5920 7444 5924 7476
rect 5956 7444 6084 7476
rect 6116 7444 6120 7476
rect 5920 7440 6120 7444
rect 6160 7476 6360 7480
rect 6160 7444 6164 7476
rect 6196 7444 6324 7476
rect 6356 7444 6360 7476
rect 6160 7440 6360 7444
rect 4240 7396 4440 7400
rect 4240 7364 4244 7396
rect 4276 7364 4404 7396
rect 4436 7364 4440 7396
rect 4240 7360 4440 7364
rect 4480 7396 4680 7400
rect 4480 7364 4484 7396
rect 4516 7364 4644 7396
rect 4676 7364 4680 7396
rect 4480 7360 4680 7364
rect 4720 7396 5080 7400
rect 4720 7364 4724 7396
rect 4756 7364 4884 7396
rect 4916 7364 5044 7396
rect 5076 7364 5080 7396
rect 4720 7360 5080 7364
rect 5120 7396 5480 7400
rect 5120 7364 5124 7396
rect 5156 7364 5284 7396
rect 5316 7364 5444 7396
rect 5476 7364 5480 7396
rect 5120 7360 5480 7364
rect 5520 7396 5880 7400
rect 5520 7364 5524 7396
rect 5556 7364 5684 7396
rect 5716 7364 5844 7396
rect 5876 7364 5880 7396
rect 5520 7360 5880 7364
rect 5920 7396 6120 7400
rect 5920 7364 5924 7396
rect 5956 7364 6084 7396
rect 6116 7364 6120 7396
rect 5920 7360 6120 7364
rect 6160 7396 6360 7400
rect 6160 7364 6164 7396
rect 6196 7364 6324 7396
rect 6356 7364 6360 7396
rect 6160 7360 6360 7364
rect 4240 7316 4440 7320
rect 4240 7284 4244 7316
rect 4276 7284 4404 7316
rect 4436 7284 4440 7316
rect 4240 7280 4440 7284
rect 4480 7316 4680 7320
rect 4480 7284 4484 7316
rect 4516 7284 4644 7316
rect 4676 7284 4680 7316
rect 4480 7280 4680 7284
rect 4720 7316 5080 7320
rect 4720 7284 4724 7316
rect 4756 7284 4884 7316
rect 4916 7284 5044 7316
rect 5076 7284 5080 7316
rect 4720 7280 5080 7284
rect 5120 7316 5480 7320
rect 5120 7284 5124 7316
rect 5156 7284 5284 7316
rect 5316 7284 5444 7316
rect 5476 7284 5480 7316
rect 5120 7280 5480 7284
rect 5520 7316 5880 7320
rect 5520 7284 5524 7316
rect 5556 7284 5684 7316
rect 5716 7284 5844 7316
rect 5876 7284 5880 7316
rect 5520 7280 5880 7284
rect 5920 7316 6120 7320
rect 5920 7284 5924 7316
rect 5956 7284 6084 7316
rect 6116 7284 6120 7316
rect 5920 7280 6120 7284
rect 6160 7316 6360 7320
rect 6160 7284 6164 7316
rect 6196 7284 6324 7316
rect 6356 7284 6360 7316
rect 6160 7280 6360 7284
rect 4240 7236 4440 7240
rect 4240 7204 4244 7236
rect 4276 7204 4404 7236
rect 4436 7204 4440 7236
rect 4240 7200 4440 7204
rect 4480 7236 4680 7240
rect 4480 7204 4484 7236
rect 4516 7204 4644 7236
rect 4676 7204 4680 7236
rect 4480 7200 4680 7204
rect 4720 7236 5080 7240
rect 4720 7204 4724 7236
rect 4756 7204 4884 7236
rect 4916 7204 5044 7236
rect 5076 7204 5080 7236
rect 4720 7200 5080 7204
rect 5120 7236 5480 7240
rect 5120 7204 5124 7236
rect 5156 7204 5284 7236
rect 5316 7204 5444 7236
rect 5476 7204 5480 7236
rect 5120 7200 5480 7204
rect 5520 7236 5880 7240
rect 5520 7204 5524 7236
rect 5556 7204 5684 7236
rect 5716 7204 5844 7236
rect 5876 7204 5880 7236
rect 5520 7200 5880 7204
rect 5920 7236 6120 7240
rect 5920 7204 5924 7236
rect 5956 7204 6084 7236
rect 6116 7204 6120 7236
rect 5920 7200 6120 7204
rect 6160 7236 6360 7240
rect 6160 7204 6164 7236
rect 6196 7204 6324 7236
rect 6356 7204 6360 7236
rect 6160 7200 6360 7204
rect 4240 7156 4440 7160
rect 4240 7124 4244 7156
rect 4276 7124 4404 7156
rect 4436 7124 4440 7156
rect 4240 7120 4440 7124
rect 4480 7156 4680 7160
rect 4480 7124 4484 7156
rect 4516 7124 4644 7156
rect 4676 7124 4680 7156
rect 4480 7120 4680 7124
rect 4720 7156 5080 7160
rect 4720 7124 4724 7156
rect 4756 7124 4884 7156
rect 4916 7124 5044 7156
rect 5076 7124 5080 7156
rect 4720 7120 5080 7124
rect 5120 7156 5480 7160
rect 5120 7124 5124 7156
rect 5156 7124 5284 7156
rect 5316 7124 5444 7156
rect 5476 7124 5480 7156
rect 5120 7120 5480 7124
rect 5520 7156 5880 7160
rect 5520 7124 5524 7156
rect 5556 7124 5684 7156
rect 5716 7124 5844 7156
rect 5876 7124 5880 7156
rect 5520 7120 5880 7124
rect 5920 7156 6120 7160
rect 5920 7124 5924 7156
rect 5956 7124 6084 7156
rect 6116 7124 6120 7156
rect 5920 7120 6120 7124
rect 6160 7156 6360 7160
rect 6160 7124 6164 7156
rect 6196 7124 6324 7156
rect 6356 7124 6360 7156
rect 6160 7120 6360 7124
rect 4240 7076 4440 7080
rect 4240 7044 4244 7076
rect 4276 7044 4404 7076
rect 4436 7044 4440 7076
rect 4240 7040 4440 7044
rect 4480 7076 4680 7080
rect 4480 7044 4484 7076
rect 4516 7044 4644 7076
rect 4676 7044 4680 7076
rect 4480 7040 4680 7044
rect 4720 7076 5080 7080
rect 4720 7044 4724 7076
rect 4756 7044 4884 7076
rect 4916 7044 5044 7076
rect 5076 7044 5080 7076
rect 4720 7040 5080 7044
rect 5120 7076 5480 7080
rect 5120 7044 5124 7076
rect 5156 7044 5284 7076
rect 5316 7044 5444 7076
rect 5476 7044 5480 7076
rect 5120 7040 5480 7044
rect 5520 7076 5880 7080
rect 5520 7044 5524 7076
rect 5556 7044 5684 7076
rect 5716 7044 5844 7076
rect 5876 7044 5880 7076
rect 5520 7040 5880 7044
rect 5920 7076 6120 7080
rect 5920 7044 5924 7076
rect 5956 7044 6084 7076
rect 6116 7044 6120 7076
rect 5920 7040 6120 7044
rect 6160 7076 6360 7080
rect 6160 7044 6164 7076
rect 6196 7044 6324 7076
rect 6356 7044 6360 7076
rect 6160 7040 6360 7044
rect 4240 6756 4440 6760
rect 4240 6724 4244 6756
rect 4276 6724 4404 6756
rect 4436 6724 4440 6756
rect 4240 6720 4440 6724
rect 4480 6756 4680 6760
rect 4480 6724 4484 6756
rect 4516 6724 4644 6756
rect 4676 6724 4680 6756
rect 4480 6720 4680 6724
rect 4720 6756 5080 6760
rect 4720 6724 4724 6756
rect 4756 6724 4884 6756
rect 4916 6724 5044 6756
rect 5076 6724 5080 6756
rect 4720 6720 5080 6724
rect 5120 6756 5480 6760
rect 5120 6724 5124 6756
rect 5156 6724 5284 6756
rect 5316 6724 5444 6756
rect 5476 6724 5480 6756
rect 5120 6720 5480 6724
rect 5520 6756 5880 6760
rect 5520 6724 5524 6756
rect 5556 6724 5684 6756
rect 5716 6724 5844 6756
rect 5876 6724 5880 6756
rect 5520 6720 5880 6724
rect 5920 6756 6120 6760
rect 5920 6724 5924 6756
rect 5956 6724 6084 6756
rect 6116 6724 6120 6756
rect 5920 6720 6120 6724
rect 6160 6756 6360 6760
rect 6160 6724 6164 6756
rect 6196 6724 6324 6756
rect 6356 6724 6360 6756
rect 6160 6720 6360 6724
rect 4240 6676 4440 6680
rect 4240 6644 4244 6676
rect 4276 6644 4404 6676
rect 4436 6644 4440 6676
rect 4240 6640 4440 6644
rect 4480 6676 4680 6680
rect 4480 6644 4484 6676
rect 4516 6644 4644 6676
rect 4676 6644 4680 6676
rect 4480 6640 4680 6644
rect 4720 6676 5080 6680
rect 4720 6644 4724 6676
rect 4756 6644 4884 6676
rect 4916 6644 5044 6676
rect 5076 6644 5080 6676
rect 4720 6640 5080 6644
rect 5120 6676 5480 6680
rect 5120 6644 5124 6676
rect 5156 6644 5284 6676
rect 5316 6644 5444 6676
rect 5476 6644 5480 6676
rect 5120 6640 5480 6644
rect 5520 6676 5880 6680
rect 5520 6644 5524 6676
rect 5556 6644 5684 6676
rect 5716 6644 5844 6676
rect 5876 6644 5880 6676
rect 5520 6640 5880 6644
rect 5920 6676 6120 6680
rect 5920 6644 5924 6676
rect 5956 6644 6084 6676
rect 6116 6644 6120 6676
rect 5920 6640 6120 6644
rect 6160 6676 6360 6680
rect 6160 6644 6164 6676
rect 6196 6644 6324 6676
rect 6356 6644 6360 6676
rect 6160 6640 6360 6644
rect 4240 6596 4440 6600
rect 4240 6564 4244 6596
rect 4276 6564 4404 6596
rect 4436 6564 4440 6596
rect 4240 6560 4440 6564
rect 4480 6596 4680 6600
rect 4480 6564 4484 6596
rect 4516 6564 4644 6596
rect 4676 6564 4680 6596
rect 4480 6560 4680 6564
rect 4720 6596 5080 6600
rect 4720 6564 4724 6596
rect 4756 6564 4884 6596
rect 4916 6564 5044 6596
rect 5076 6564 5080 6596
rect 4720 6560 5080 6564
rect 5120 6596 5480 6600
rect 5120 6564 5124 6596
rect 5156 6564 5284 6596
rect 5316 6564 5444 6596
rect 5476 6564 5480 6596
rect 5120 6560 5480 6564
rect 5520 6596 5880 6600
rect 5520 6564 5524 6596
rect 5556 6564 5684 6596
rect 5716 6564 5844 6596
rect 5876 6564 5880 6596
rect 5520 6560 5880 6564
rect 5920 6596 6120 6600
rect 5920 6564 5924 6596
rect 5956 6564 6084 6596
rect 6116 6564 6120 6596
rect 5920 6560 6120 6564
rect 6160 6596 6360 6600
rect 6160 6564 6164 6596
rect 6196 6564 6324 6596
rect 6356 6564 6360 6596
rect 6160 6560 6360 6564
rect 4240 6516 4440 6520
rect 4240 6484 4244 6516
rect 4276 6484 4404 6516
rect 4436 6484 4440 6516
rect 4240 6480 4440 6484
rect 4480 6516 4680 6520
rect 4480 6484 4484 6516
rect 4516 6484 4644 6516
rect 4676 6484 4680 6516
rect 4480 6480 4680 6484
rect 4720 6516 5080 6520
rect 4720 6484 4724 6516
rect 4756 6484 4884 6516
rect 4916 6484 5044 6516
rect 5076 6484 5080 6516
rect 4720 6480 5080 6484
rect 5120 6516 5480 6520
rect 5120 6484 5124 6516
rect 5156 6484 5284 6516
rect 5316 6484 5444 6516
rect 5476 6484 5480 6516
rect 5120 6480 5480 6484
rect 5520 6516 5880 6520
rect 5520 6484 5524 6516
rect 5556 6484 5684 6516
rect 5716 6484 5844 6516
rect 5876 6484 5880 6516
rect 5520 6480 5880 6484
rect 5920 6516 6120 6520
rect 5920 6484 5924 6516
rect 5956 6484 6084 6516
rect 6116 6484 6120 6516
rect 5920 6480 6120 6484
rect 6160 6516 6360 6520
rect 6160 6484 6164 6516
rect 6196 6484 6324 6516
rect 6356 6484 6360 6516
rect 6160 6480 6360 6484
rect 4240 6436 4440 6440
rect 4240 6404 4244 6436
rect 4276 6404 4404 6436
rect 4436 6404 4440 6436
rect 4240 6400 4440 6404
rect 4480 6436 4680 6440
rect 4480 6404 4484 6436
rect 4516 6404 4644 6436
rect 4676 6404 4680 6436
rect 4480 6400 4680 6404
rect 4720 6436 5080 6440
rect 4720 6404 4724 6436
rect 4756 6404 4884 6436
rect 4916 6404 5044 6436
rect 5076 6404 5080 6436
rect 4720 6400 5080 6404
rect 5120 6436 5480 6440
rect 5120 6404 5124 6436
rect 5156 6404 5284 6436
rect 5316 6404 5444 6436
rect 5476 6404 5480 6436
rect 5120 6400 5480 6404
rect 5520 6436 5880 6440
rect 5520 6404 5524 6436
rect 5556 6404 5684 6436
rect 5716 6404 5844 6436
rect 5876 6404 5880 6436
rect 5520 6400 5880 6404
rect 5920 6436 6120 6440
rect 5920 6404 5924 6436
rect 5956 6404 6084 6436
rect 6116 6404 6120 6436
rect 5920 6400 6120 6404
rect 6160 6436 6360 6440
rect 6160 6404 6164 6436
rect 6196 6404 6324 6436
rect 6356 6404 6360 6436
rect 6160 6400 6360 6404
rect 4240 6356 4440 6360
rect 4240 6324 4244 6356
rect 4276 6324 4404 6356
rect 4436 6324 4440 6356
rect 4240 6320 4440 6324
rect 4480 6356 4680 6360
rect 4480 6324 4484 6356
rect 4516 6324 4644 6356
rect 4676 6324 4680 6356
rect 4480 6320 4680 6324
rect 4720 6356 5080 6360
rect 4720 6324 4724 6356
rect 4756 6324 4884 6356
rect 4916 6324 5044 6356
rect 5076 6324 5080 6356
rect 4720 6320 5080 6324
rect 5120 6356 5480 6360
rect 5120 6324 5124 6356
rect 5156 6324 5284 6356
rect 5316 6324 5444 6356
rect 5476 6324 5480 6356
rect 5120 6320 5480 6324
rect 5520 6356 5880 6360
rect 5520 6324 5524 6356
rect 5556 6324 5684 6356
rect 5716 6324 5844 6356
rect 5876 6324 5880 6356
rect 5520 6320 5880 6324
rect 5920 6356 6120 6360
rect 5920 6324 5924 6356
rect 5956 6324 6084 6356
rect 6116 6324 6120 6356
rect 5920 6320 6120 6324
rect 6160 6356 6360 6360
rect 6160 6324 6164 6356
rect 6196 6324 6324 6356
rect 6356 6324 6360 6356
rect 6160 6320 6360 6324
rect 4240 5796 4440 5800
rect 4240 5764 4244 5796
rect 4276 5764 4404 5796
rect 4436 5764 4440 5796
rect 4240 5760 4440 5764
rect 4480 5796 4680 5800
rect 4480 5764 4484 5796
rect 4516 5764 4644 5796
rect 4676 5764 4680 5796
rect 4480 5760 4680 5764
rect 4720 5796 5080 5800
rect 4720 5764 4724 5796
rect 4756 5764 4884 5796
rect 4916 5764 5044 5796
rect 5076 5764 5080 5796
rect 4720 5760 5080 5764
rect 5120 5796 5480 5800
rect 5120 5764 5124 5796
rect 5156 5764 5284 5796
rect 5316 5764 5444 5796
rect 5476 5764 5480 5796
rect 5120 5760 5480 5764
rect 5520 5796 5880 5800
rect 5520 5764 5524 5796
rect 5556 5764 5684 5796
rect 5716 5764 5844 5796
rect 5876 5764 5880 5796
rect 5520 5760 5880 5764
rect 5920 5796 6120 5800
rect 5920 5764 5924 5796
rect 5956 5764 6084 5796
rect 6116 5764 6120 5796
rect 5920 5760 6120 5764
rect 6160 5796 6360 5800
rect 6160 5764 6164 5796
rect 6196 5764 6324 5796
rect 6356 5764 6360 5796
rect 6160 5760 6360 5764
rect 4240 5716 4440 5720
rect 4240 5684 4244 5716
rect 4276 5684 4404 5716
rect 4436 5684 4440 5716
rect 4240 5680 4440 5684
rect 4480 5716 4680 5720
rect 4480 5684 4484 5716
rect 4516 5684 4644 5716
rect 4676 5684 4680 5716
rect 4480 5680 4680 5684
rect 4720 5716 5080 5720
rect 4720 5684 4724 5716
rect 4756 5684 4884 5716
rect 4916 5684 5044 5716
rect 5076 5684 5080 5716
rect 4720 5680 5080 5684
rect 5120 5716 5480 5720
rect 5120 5684 5124 5716
rect 5156 5684 5284 5716
rect 5316 5684 5444 5716
rect 5476 5684 5480 5716
rect 5120 5680 5480 5684
rect 5520 5716 5880 5720
rect 5520 5684 5524 5716
rect 5556 5684 5684 5716
rect 5716 5684 5844 5716
rect 5876 5684 5880 5716
rect 5520 5680 5880 5684
rect 5920 5716 6120 5720
rect 5920 5684 5924 5716
rect 5956 5684 6084 5716
rect 6116 5684 6120 5716
rect 5920 5680 6120 5684
rect 6160 5716 6360 5720
rect 6160 5684 6164 5716
rect 6196 5684 6324 5716
rect 6356 5684 6360 5716
rect 6160 5680 6360 5684
rect 4240 5636 4440 5640
rect 4240 5604 4244 5636
rect 4276 5604 4404 5636
rect 4436 5604 4440 5636
rect 4240 5600 4440 5604
rect 4480 5636 4680 5640
rect 4480 5604 4484 5636
rect 4516 5604 4644 5636
rect 4676 5604 4680 5636
rect 4480 5600 4680 5604
rect 4720 5636 5080 5640
rect 4720 5604 4724 5636
rect 4756 5604 4884 5636
rect 4916 5604 5044 5636
rect 5076 5604 5080 5636
rect 4720 5600 5080 5604
rect 5120 5636 5480 5640
rect 5120 5604 5124 5636
rect 5156 5604 5284 5636
rect 5316 5604 5444 5636
rect 5476 5604 5480 5636
rect 5120 5600 5480 5604
rect 5520 5636 5880 5640
rect 5520 5604 5524 5636
rect 5556 5604 5684 5636
rect 5716 5604 5844 5636
rect 5876 5604 5880 5636
rect 5520 5600 5880 5604
rect 5920 5636 6120 5640
rect 5920 5604 5924 5636
rect 5956 5604 6084 5636
rect 6116 5604 6120 5636
rect 5920 5600 6120 5604
rect 6160 5636 6360 5640
rect 6160 5604 6164 5636
rect 6196 5604 6324 5636
rect 6356 5604 6360 5636
rect 6160 5600 6360 5604
rect 4240 5556 4440 5560
rect 4240 5524 4244 5556
rect 4276 5524 4404 5556
rect 4436 5524 4440 5556
rect 4240 5520 4440 5524
rect 4480 5556 4680 5560
rect 4480 5524 4484 5556
rect 4516 5524 4644 5556
rect 4676 5524 4680 5556
rect 4480 5520 4680 5524
rect 4720 5556 5080 5560
rect 4720 5524 4724 5556
rect 4756 5524 4884 5556
rect 4916 5524 5044 5556
rect 5076 5524 5080 5556
rect 4720 5520 5080 5524
rect 5120 5556 5480 5560
rect 5120 5524 5124 5556
rect 5156 5524 5284 5556
rect 5316 5524 5444 5556
rect 5476 5524 5480 5556
rect 5120 5520 5480 5524
rect 5520 5556 5880 5560
rect 5520 5524 5524 5556
rect 5556 5524 5684 5556
rect 5716 5524 5844 5556
rect 5876 5524 5880 5556
rect 5520 5520 5880 5524
rect 5920 5556 6120 5560
rect 5920 5524 5924 5556
rect 5956 5524 6084 5556
rect 6116 5524 6120 5556
rect 5920 5520 6120 5524
rect 6160 5556 6360 5560
rect 6160 5524 6164 5556
rect 6196 5524 6324 5556
rect 6356 5524 6360 5556
rect 6160 5520 6360 5524
rect 4240 5476 4440 5480
rect 4240 5444 4244 5476
rect 4276 5444 4404 5476
rect 4436 5444 4440 5476
rect 4240 5440 4440 5444
rect 4480 5476 4680 5480
rect 4480 5444 4484 5476
rect 4516 5444 4644 5476
rect 4676 5444 4680 5476
rect 4480 5440 4680 5444
rect 4720 5476 5080 5480
rect 4720 5444 4724 5476
rect 4756 5444 4884 5476
rect 4916 5444 5044 5476
rect 5076 5444 5080 5476
rect 4720 5440 5080 5444
rect 5120 5476 5480 5480
rect 5120 5444 5124 5476
rect 5156 5444 5284 5476
rect 5316 5444 5444 5476
rect 5476 5444 5480 5476
rect 5120 5440 5480 5444
rect 5520 5476 5880 5480
rect 5520 5444 5524 5476
rect 5556 5444 5684 5476
rect 5716 5444 5844 5476
rect 5876 5444 5880 5476
rect 5520 5440 5880 5444
rect 5920 5476 6120 5480
rect 5920 5444 5924 5476
rect 5956 5444 6084 5476
rect 6116 5444 6120 5476
rect 5920 5440 6120 5444
rect 6160 5476 6360 5480
rect 6160 5444 6164 5476
rect 6196 5444 6324 5476
rect 6356 5444 6360 5476
rect 6160 5440 6360 5444
rect 4240 5396 4440 5400
rect 4240 5364 4244 5396
rect 4276 5364 4404 5396
rect 4436 5364 4440 5396
rect 4240 5360 4440 5364
rect 4480 5396 4680 5400
rect 4480 5364 4484 5396
rect 4516 5364 4644 5396
rect 4676 5364 4680 5396
rect 4480 5360 4680 5364
rect 4720 5396 5080 5400
rect 4720 5364 4724 5396
rect 4756 5364 4884 5396
rect 4916 5364 5044 5396
rect 5076 5364 5080 5396
rect 4720 5360 5080 5364
rect 5120 5396 5480 5400
rect 5120 5364 5124 5396
rect 5156 5364 5284 5396
rect 5316 5364 5444 5396
rect 5476 5364 5480 5396
rect 5120 5360 5480 5364
rect 5520 5396 5880 5400
rect 5520 5364 5524 5396
rect 5556 5364 5684 5396
rect 5716 5364 5844 5396
rect 5876 5364 5880 5396
rect 5520 5360 5880 5364
rect 5920 5396 6120 5400
rect 5920 5364 5924 5396
rect 5956 5364 6084 5396
rect 6116 5364 6120 5396
rect 5920 5360 6120 5364
rect 6160 5396 6360 5400
rect 6160 5364 6164 5396
rect 6196 5364 6324 5396
rect 6356 5364 6360 5396
rect 6160 5360 6360 5364
rect 4240 5316 4440 5320
rect 4240 5284 4244 5316
rect 4276 5284 4404 5316
rect 4436 5284 4440 5316
rect 4240 5280 4440 5284
rect 4480 5316 4680 5320
rect 4480 5284 4484 5316
rect 4516 5284 4644 5316
rect 4676 5284 4680 5316
rect 4480 5280 4680 5284
rect 4720 5316 5080 5320
rect 4720 5284 4724 5316
rect 4756 5284 4884 5316
rect 4916 5284 5044 5316
rect 5076 5284 5080 5316
rect 4720 5280 5080 5284
rect 5120 5316 5480 5320
rect 5120 5284 5124 5316
rect 5156 5284 5284 5316
rect 5316 5284 5444 5316
rect 5476 5284 5480 5316
rect 5120 5280 5480 5284
rect 5520 5316 5880 5320
rect 5520 5284 5524 5316
rect 5556 5284 5684 5316
rect 5716 5284 5844 5316
rect 5876 5284 5880 5316
rect 5520 5280 5880 5284
rect 5920 5316 6120 5320
rect 5920 5284 5924 5316
rect 5956 5284 6084 5316
rect 6116 5284 6120 5316
rect 5920 5280 6120 5284
rect 6160 5316 6360 5320
rect 6160 5284 6164 5316
rect 6196 5284 6324 5316
rect 6356 5284 6360 5316
rect 6160 5280 6360 5284
rect 4240 5236 4440 5240
rect 4240 5204 4244 5236
rect 4276 5204 4404 5236
rect 4436 5204 4440 5236
rect 4240 5200 4440 5204
rect 4480 5236 4680 5240
rect 4480 5204 4484 5236
rect 4516 5204 4644 5236
rect 4676 5204 4680 5236
rect 4480 5200 4680 5204
rect 4720 5236 5080 5240
rect 4720 5204 4724 5236
rect 4756 5204 4884 5236
rect 4916 5204 5044 5236
rect 5076 5204 5080 5236
rect 4720 5200 5080 5204
rect 5120 5236 5480 5240
rect 5120 5204 5124 5236
rect 5156 5204 5284 5236
rect 5316 5204 5444 5236
rect 5476 5204 5480 5236
rect 5120 5200 5480 5204
rect 5520 5236 5880 5240
rect 5520 5204 5524 5236
rect 5556 5204 5684 5236
rect 5716 5204 5844 5236
rect 5876 5204 5880 5236
rect 5520 5200 5880 5204
rect 5920 5236 6120 5240
rect 5920 5204 5924 5236
rect 5956 5204 6084 5236
rect 6116 5204 6120 5236
rect 5920 5200 6120 5204
rect 6160 5236 6360 5240
rect 6160 5204 6164 5236
rect 6196 5204 6324 5236
rect 6356 5204 6360 5236
rect 6160 5200 6360 5204
rect 4240 5156 4440 5160
rect 4240 5124 4244 5156
rect 4276 5124 4404 5156
rect 4436 5124 4440 5156
rect 4240 5120 4440 5124
rect 4480 5156 4680 5160
rect 4480 5124 4484 5156
rect 4516 5124 4644 5156
rect 4676 5124 4680 5156
rect 4480 5120 4680 5124
rect 4720 5156 5080 5160
rect 4720 5124 4724 5156
rect 4756 5124 4884 5156
rect 4916 5124 5044 5156
rect 5076 5124 5080 5156
rect 4720 5120 5080 5124
rect 5120 5156 5480 5160
rect 5120 5124 5124 5156
rect 5156 5124 5284 5156
rect 5316 5124 5444 5156
rect 5476 5124 5480 5156
rect 5120 5120 5480 5124
rect 5520 5156 5880 5160
rect 5520 5124 5524 5156
rect 5556 5124 5684 5156
rect 5716 5124 5844 5156
rect 5876 5124 5880 5156
rect 5520 5120 5880 5124
rect 5920 5156 6120 5160
rect 5920 5124 5924 5156
rect 5956 5124 6084 5156
rect 6116 5124 6120 5156
rect 5920 5120 6120 5124
rect 6160 5156 6360 5160
rect 6160 5124 6164 5156
rect 6196 5124 6324 5156
rect 6356 5124 6360 5156
rect 6160 5120 6360 5124
rect 4240 5076 4440 5080
rect 4240 5044 4244 5076
rect 4276 5044 4404 5076
rect 4436 5044 4440 5076
rect 4240 5040 4440 5044
rect 4480 5076 4680 5080
rect 4480 5044 4484 5076
rect 4516 5044 4644 5076
rect 4676 5044 4680 5076
rect 4480 5040 4680 5044
rect 4720 5076 5080 5080
rect 4720 5044 4724 5076
rect 4756 5044 4884 5076
rect 4916 5044 5044 5076
rect 5076 5044 5080 5076
rect 4720 5040 5080 5044
rect 5120 5076 5480 5080
rect 5120 5044 5124 5076
rect 5156 5044 5284 5076
rect 5316 5044 5444 5076
rect 5476 5044 5480 5076
rect 5120 5040 5480 5044
rect 5520 5076 5880 5080
rect 5520 5044 5524 5076
rect 5556 5044 5684 5076
rect 5716 5044 5844 5076
rect 5876 5044 5880 5076
rect 5520 5040 5880 5044
rect 5920 5076 6120 5080
rect 5920 5044 5924 5076
rect 5956 5044 6084 5076
rect 6116 5044 6120 5076
rect 5920 5040 6120 5044
rect 6160 5076 6360 5080
rect 6160 5044 6164 5076
rect 6196 5044 6324 5076
rect 6356 5044 6360 5076
rect 6160 5040 6360 5044
rect 4240 4996 4440 5000
rect 4240 4964 4244 4996
rect 4276 4964 4404 4996
rect 4436 4964 4440 4996
rect 4240 4960 4440 4964
rect 4480 4996 4680 5000
rect 4480 4964 4484 4996
rect 4516 4964 4644 4996
rect 4676 4964 4680 4996
rect 4480 4960 4680 4964
rect 4720 4996 5080 5000
rect 4720 4964 4724 4996
rect 4756 4964 4884 4996
rect 4916 4964 5044 4996
rect 5076 4964 5080 4996
rect 4720 4960 5080 4964
rect 5120 4996 5480 5000
rect 5120 4964 5124 4996
rect 5156 4964 5284 4996
rect 5316 4964 5444 4996
rect 5476 4964 5480 4996
rect 5120 4960 5480 4964
rect 5520 4996 5880 5000
rect 5520 4964 5524 4996
rect 5556 4964 5684 4996
rect 5716 4964 5844 4996
rect 5876 4964 5880 4996
rect 5520 4960 5880 4964
rect 5920 4996 6120 5000
rect 5920 4964 5924 4996
rect 5956 4964 6084 4996
rect 6116 4964 6120 4996
rect 5920 4960 6120 4964
rect 6160 4996 6360 5000
rect 6160 4964 6164 4996
rect 6196 4964 6324 4996
rect 6356 4964 6360 4996
rect 6160 4960 6360 4964
rect 4240 4436 4440 4440
rect 4240 4404 4244 4436
rect 4276 4404 4404 4436
rect 4436 4404 4440 4436
rect 4240 4400 4440 4404
rect 4480 4436 4680 4440
rect 4480 4404 4484 4436
rect 4516 4404 4644 4436
rect 4676 4404 4680 4436
rect 4480 4400 4680 4404
rect 4720 4436 5080 4440
rect 4720 4404 4724 4436
rect 4756 4404 4884 4436
rect 4916 4404 5044 4436
rect 5076 4404 5080 4436
rect 4720 4400 5080 4404
rect 5120 4436 5480 4440
rect 5120 4404 5124 4436
rect 5156 4404 5284 4436
rect 5316 4404 5444 4436
rect 5476 4404 5480 4436
rect 5120 4400 5480 4404
rect 5520 4436 5880 4440
rect 5520 4404 5524 4436
rect 5556 4404 5684 4436
rect 5716 4404 5844 4436
rect 5876 4404 5880 4436
rect 5520 4400 5880 4404
rect 5920 4436 6120 4440
rect 5920 4404 5924 4436
rect 5956 4404 6084 4436
rect 6116 4404 6120 4436
rect 5920 4400 6120 4404
rect 6160 4436 6360 4440
rect 6160 4404 6164 4436
rect 6196 4404 6324 4436
rect 6356 4404 6360 4436
rect 6160 4400 6360 4404
rect 4240 4356 4440 4360
rect 4240 4324 4244 4356
rect 4276 4324 4404 4356
rect 4436 4324 4440 4356
rect 4240 4320 4440 4324
rect 4480 4356 4680 4360
rect 4480 4324 4484 4356
rect 4516 4324 4644 4356
rect 4676 4324 4680 4356
rect 4480 4320 4680 4324
rect 4720 4356 5080 4360
rect 4720 4324 4724 4356
rect 4756 4324 4884 4356
rect 4916 4324 5044 4356
rect 5076 4324 5080 4356
rect 4720 4320 5080 4324
rect 5120 4356 5480 4360
rect 5120 4324 5124 4356
rect 5156 4324 5284 4356
rect 5316 4324 5444 4356
rect 5476 4324 5480 4356
rect 5120 4320 5480 4324
rect 5520 4356 5880 4360
rect 5520 4324 5524 4356
rect 5556 4324 5684 4356
rect 5716 4324 5844 4356
rect 5876 4324 5880 4356
rect 5520 4320 5880 4324
rect 5920 4356 6120 4360
rect 5920 4324 5924 4356
rect 5956 4324 6084 4356
rect 6116 4324 6120 4356
rect 5920 4320 6120 4324
rect 6160 4356 6360 4360
rect 6160 4324 6164 4356
rect 6196 4324 6324 4356
rect 6356 4324 6360 4356
rect 6160 4320 6360 4324
rect 4240 4276 4440 4280
rect 4240 4244 4244 4276
rect 4276 4244 4404 4276
rect 4436 4244 4440 4276
rect 4240 4240 4440 4244
rect 4480 4276 4680 4280
rect 4480 4244 4484 4276
rect 4516 4244 4644 4276
rect 4676 4244 4680 4276
rect 4480 4240 4680 4244
rect 4720 4276 5080 4280
rect 4720 4244 4724 4276
rect 4756 4244 4884 4276
rect 4916 4244 5044 4276
rect 5076 4244 5080 4276
rect 4720 4240 5080 4244
rect 5120 4276 5480 4280
rect 5120 4244 5124 4276
rect 5156 4244 5284 4276
rect 5316 4244 5444 4276
rect 5476 4244 5480 4276
rect 5120 4240 5480 4244
rect 5520 4276 5880 4280
rect 5520 4244 5524 4276
rect 5556 4244 5684 4276
rect 5716 4244 5844 4276
rect 5876 4244 5880 4276
rect 5520 4240 5880 4244
rect 5920 4276 6120 4280
rect 5920 4244 5924 4276
rect 5956 4244 6084 4276
rect 6116 4244 6120 4276
rect 5920 4240 6120 4244
rect 6160 4276 6360 4280
rect 6160 4244 6164 4276
rect 6196 4244 6324 4276
rect 6356 4244 6360 4276
rect 6160 4240 6360 4244
rect 4240 4196 4440 4200
rect 4240 4164 4244 4196
rect 4276 4164 4404 4196
rect 4436 4164 4440 4196
rect 4240 4160 4440 4164
rect 4480 4196 4680 4200
rect 4480 4164 4484 4196
rect 4516 4164 4644 4196
rect 4676 4164 4680 4196
rect 4480 4160 4680 4164
rect 4720 4196 5080 4200
rect 4720 4164 4724 4196
rect 4756 4164 4884 4196
rect 4916 4164 5044 4196
rect 5076 4164 5080 4196
rect 4720 4160 5080 4164
rect 5120 4196 5480 4200
rect 5120 4164 5124 4196
rect 5156 4164 5284 4196
rect 5316 4164 5444 4196
rect 5476 4164 5480 4196
rect 5120 4160 5480 4164
rect 5520 4196 5880 4200
rect 5520 4164 5524 4196
rect 5556 4164 5684 4196
rect 5716 4164 5844 4196
rect 5876 4164 5880 4196
rect 5520 4160 5880 4164
rect 5920 4196 6120 4200
rect 5920 4164 5924 4196
rect 5956 4164 6084 4196
rect 6116 4164 6120 4196
rect 5920 4160 6120 4164
rect 6160 4196 6360 4200
rect 6160 4164 6164 4196
rect 6196 4164 6324 4196
rect 6356 4164 6360 4196
rect 6160 4160 6360 4164
rect 4240 4116 4440 4120
rect 4240 4084 4244 4116
rect 4276 4084 4404 4116
rect 4436 4084 4440 4116
rect 4240 4080 4440 4084
rect 4480 4116 4680 4120
rect 4480 4084 4484 4116
rect 4516 4084 4644 4116
rect 4676 4084 4680 4116
rect 4480 4080 4680 4084
rect 4720 4116 5080 4120
rect 4720 4084 4724 4116
rect 4756 4084 4884 4116
rect 4916 4084 5044 4116
rect 5076 4084 5080 4116
rect 4720 4080 5080 4084
rect 5120 4116 5480 4120
rect 5120 4084 5124 4116
rect 5156 4084 5284 4116
rect 5316 4084 5444 4116
rect 5476 4084 5480 4116
rect 5120 4080 5480 4084
rect 5520 4116 5880 4120
rect 5520 4084 5524 4116
rect 5556 4084 5684 4116
rect 5716 4084 5844 4116
rect 5876 4084 5880 4116
rect 5520 4080 5880 4084
rect 5920 4116 6120 4120
rect 5920 4084 5924 4116
rect 5956 4084 6084 4116
rect 6116 4084 6120 4116
rect 5920 4080 6120 4084
rect 6160 4116 6360 4120
rect 6160 4084 6164 4116
rect 6196 4084 6324 4116
rect 6356 4084 6360 4116
rect 6160 4080 6360 4084
rect 4240 4036 4440 4040
rect 4240 4004 4244 4036
rect 4276 4004 4404 4036
rect 4436 4004 4440 4036
rect 4240 4000 4440 4004
rect 4480 4036 4680 4040
rect 4480 4004 4484 4036
rect 4516 4004 4644 4036
rect 4676 4004 4680 4036
rect 4480 4000 4680 4004
rect 4720 4036 5080 4040
rect 4720 4004 4724 4036
rect 4756 4004 4884 4036
rect 4916 4004 5044 4036
rect 5076 4004 5080 4036
rect 4720 4000 5080 4004
rect 5120 4036 5480 4040
rect 5120 4004 5124 4036
rect 5156 4004 5284 4036
rect 5316 4004 5444 4036
rect 5476 4004 5480 4036
rect 5120 4000 5480 4004
rect 5520 4036 5880 4040
rect 5520 4004 5524 4036
rect 5556 4004 5684 4036
rect 5716 4004 5844 4036
rect 5876 4004 5880 4036
rect 5520 4000 5880 4004
rect 5920 4036 6120 4040
rect 5920 4004 5924 4036
rect 5956 4004 6084 4036
rect 6116 4004 6120 4036
rect 5920 4000 6120 4004
rect 6160 4036 6360 4040
rect 6160 4004 6164 4036
rect 6196 4004 6324 4036
rect 6356 4004 6360 4036
rect 6160 4000 6360 4004
rect 4240 3956 4440 3960
rect 4240 3924 4244 3956
rect 4276 3924 4404 3956
rect 4436 3924 4440 3956
rect 4240 3920 4440 3924
rect 4480 3956 4680 3960
rect 4480 3924 4484 3956
rect 4516 3924 4644 3956
rect 4676 3924 4680 3956
rect 4480 3920 4680 3924
rect 4720 3956 5080 3960
rect 4720 3924 4724 3956
rect 4756 3924 4884 3956
rect 4916 3924 5044 3956
rect 5076 3924 5080 3956
rect 4720 3920 5080 3924
rect 5120 3956 5480 3960
rect 5120 3924 5124 3956
rect 5156 3924 5284 3956
rect 5316 3924 5444 3956
rect 5476 3924 5480 3956
rect 5120 3920 5480 3924
rect 5520 3956 5880 3960
rect 5520 3924 5524 3956
rect 5556 3924 5684 3956
rect 5716 3924 5844 3956
rect 5876 3924 5880 3956
rect 5520 3920 5880 3924
rect 5920 3956 6120 3960
rect 5920 3924 5924 3956
rect 5956 3924 6084 3956
rect 6116 3924 6120 3956
rect 5920 3920 6120 3924
rect 6160 3956 6360 3960
rect 6160 3924 6164 3956
rect 6196 3924 6324 3956
rect 6356 3924 6360 3956
rect 6160 3920 6360 3924
rect 4240 3156 4440 3160
rect 4240 3124 4244 3156
rect 4276 3124 4404 3156
rect 4436 3124 4440 3156
rect 4240 3120 4440 3124
rect 4480 3156 4680 3160
rect 4480 3124 4484 3156
rect 4516 3124 4644 3156
rect 4676 3124 4680 3156
rect 4480 3120 4680 3124
rect 4720 3156 5080 3160
rect 4720 3124 4724 3156
rect 4756 3124 4884 3156
rect 4916 3124 5044 3156
rect 5076 3124 5080 3156
rect 4720 3120 5080 3124
rect 5120 3156 5480 3160
rect 5120 3124 5124 3156
rect 5156 3124 5284 3156
rect 5316 3124 5444 3156
rect 5476 3124 5480 3156
rect 5120 3120 5480 3124
rect 5520 3156 5880 3160
rect 5520 3124 5524 3156
rect 5556 3124 5684 3156
rect 5716 3124 5844 3156
rect 5876 3124 5880 3156
rect 5520 3120 5880 3124
rect 5920 3156 6120 3160
rect 5920 3124 5924 3156
rect 5956 3124 6084 3156
rect 6116 3124 6120 3156
rect 5920 3120 6120 3124
rect 6160 3156 6360 3160
rect 6160 3124 6164 3156
rect 6196 3124 6324 3156
rect 6356 3124 6360 3156
rect 6160 3120 6360 3124
rect 4240 3076 4440 3080
rect 4240 3044 4244 3076
rect 4276 3044 4404 3076
rect 4436 3044 4440 3076
rect 4240 3040 4440 3044
rect 4480 3076 4680 3080
rect 4480 3044 4484 3076
rect 4516 3044 4644 3076
rect 4676 3044 4680 3076
rect 4480 3040 4680 3044
rect 4720 3076 5080 3080
rect 4720 3044 4724 3076
rect 4756 3044 4884 3076
rect 4916 3044 5044 3076
rect 5076 3044 5080 3076
rect 4720 3040 5080 3044
rect 5120 3076 5480 3080
rect 5120 3044 5124 3076
rect 5156 3044 5284 3076
rect 5316 3044 5444 3076
rect 5476 3044 5480 3076
rect 5120 3040 5480 3044
rect 5520 3076 5880 3080
rect 5520 3044 5524 3076
rect 5556 3044 5684 3076
rect 5716 3044 5844 3076
rect 5876 3044 5880 3076
rect 5520 3040 5880 3044
rect 5920 3076 6120 3080
rect 5920 3044 5924 3076
rect 5956 3044 6084 3076
rect 6116 3044 6120 3076
rect 5920 3040 6120 3044
rect 6160 3076 6360 3080
rect 6160 3044 6164 3076
rect 6196 3044 6324 3076
rect 6356 3044 6360 3076
rect 6160 3040 6360 3044
rect 4240 2996 4440 3000
rect 4240 2964 4244 2996
rect 4276 2964 4404 2996
rect 4436 2964 4440 2996
rect 4240 2960 4440 2964
rect 4480 2996 4680 3000
rect 4480 2964 4484 2996
rect 4516 2964 4644 2996
rect 4676 2964 4680 2996
rect 4480 2960 4680 2964
rect 4720 2996 5080 3000
rect 4720 2964 4724 2996
rect 4756 2964 4884 2996
rect 4916 2964 5044 2996
rect 5076 2964 5080 2996
rect 4720 2960 5080 2964
rect 5120 2996 5480 3000
rect 5120 2964 5124 2996
rect 5156 2964 5284 2996
rect 5316 2964 5444 2996
rect 5476 2964 5480 2996
rect 5120 2960 5480 2964
rect 5520 2996 5880 3000
rect 5520 2964 5524 2996
rect 5556 2964 5684 2996
rect 5716 2964 5844 2996
rect 5876 2964 5880 2996
rect 5520 2960 5880 2964
rect 5920 2996 6120 3000
rect 5920 2964 5924 2996
rect 5956 2964 6084 2996
rect 6116 2964 6120 2996
rect 5920 2960 6120 2964
rect 6160 2996 6360 3000
rect 6160 2964 6164 2996
rect 6196 2964 6324 2996
rect 6356 2964 6360 2996
rect 6160 2960 6360 2964
rect 4240 2916 4440 2920
rect 4240 2884 4244 2916
rect 4276 2884 4404 2916
rect 4436 2884 4440 2916
rect 4240 2880 4440 2884
rect 4480 2916 4680 2920
rect 4480 2884 4484 2916
rect 4516 2884 4644 2916
rect 4676 2884 4680 2916
rect 4480 2880 4680 2884
rect 4720 2916 5080 2920
rect 4720 2884 4724 2916
rect 4756 2884 4884 2916
rect 4916 2884 5044 2916
rect 5076 2884 5080 2916
rect 4720 2880 5080 2884
rect 5120 2916 5480 2920
rect 5120 2884 5124 2916
rect 5156 2884 5284 2916
rect 5316 2884 5444 2916
rect 5476 2884 5480 2916
rect 5120 2880 5480 2884
rect 5520 2916 5880 2920
rect 5520 2884 5524 2916
rect 5556 2884 5684 2916
rect 5716 2884 5844 2916
rect 5876 2884 5880 2916
rect 5520 2880 5880 2884
rect 5920 2916 6120 2920
rect 5920 2884 5924 2916
rect 5956 2884 6084 2916
rect 6116 2884 6120 2916
rect 5920 2880 6120 2884
rect 6160 2916 6360 2920
rect 6160 2884 6164 2916
rect 6196 2884 6324 2916
rect 6356 2884 6360 2916
rect 6160 2880 6360 2884
rect 4240 2836 4440 2840
rect 4240 2804 4244 2836
rect 4276 2804 4404 2836
rect 4436 2804 4440 2836
rect 4240 2800 4440 2804
rect 4480 2836 4680 2840
rect 4480 2804 4484 2836
rect 4516 2804 4644 2836
rect 4676 2804 4680 2836
rect 4480 2800 4680 2804
rect 4720 2836 5080 2840
rect 4720 2804 4724 2836
rect 4756 2804 4884 2836
rect 4916 2804 5044 2836
rect 5076 2804 5080 2836
rect 4720 2800 5080 2804
rect 5120 2836 5480 2840
rect 5120 2804 5124 2836
rect 5156 2804 5284 2836
rect 5316 2804 5444 2836
rect 5476 2804 5480 2836
rect 5120 2800 5480 2804
rect 5520 2836 5880 2840
rect 5520 2804 5524 2836
rect 5556 2804 5684 2836
rect 5716 2804 5844 2836
rect 5876 2804 5880 2836
rect 5520 2800 5880 2804
rect 5920 2836 6120 2840
rect 5920 2804 5924 2836
rect 5956 2804 6084 2836
rect 6116 2804 6120 2836
rect 5920 2800 6120 2804
rect 6160 2836 6360 2840
rect 6160 2804 6164 2836
rect 6196 2804 6324 2836
rect 6356 2804 6360 2836
rect 6160 2800 6360 2804
rect 4240 2756 4440 2760
rect 4240 2724 4244 2756
rect 4276 2724 4404 2756
rect 4436 2724 4440 2756
rect 4240 2720 4440 2724
rect 4480 2756 4680 2760
rect 4480 2724 4484 2756
rect 4516 2724 4644 2756
rect 4676 2724 4680 2756
rect 4480 2720 4680 2724
rect 4720 2756 5080 2760
rect 4720 2724 4724 2756
rect 4756 2724 4884 2756
rect 4916 2724 5044 2756
rect 5076 2724 5080 2756
rect 4720 2720 5080 2724
rect 5120 2756 5480 2760
rect 5120 2724 5124 2756
rect 5156 2724 5284 2756
rect 5316 2724 5444 2756
rect 5476 2724 5480 2756
rect 5120 2720 5480 2724
rect 5520 2756 5880 2760
rect 5520 2724 5524 2756
rect 5556 2724 5684 2756
rect 5716 2724 5844 2756
rect 5876 2724 5880 2756
rect 5520 2720 5880 2724
rect 5920 2756 6120 2760
rect 5920 2724 5924 2756
rect 5956 2724 6084 2756
rect 6116 2724 6120 2756
rect 5920 2720 6120 2724
rect 6160 2756 6360 2760
rect 6160 2724 6164 2756
rect 6196 2724 6324 2756
rect 6356 2724 6360 2756
rect 6160 2720 6360 2724
rect 4240 2676 4440 2680
rect 4240 2644 4244 2676
rect 4276 2644 4404 2676
rect 4436 2644 4440 2676
rect 4240 2640 4440 2644
rect 4480 2676 4680 2680
rect 4480 2644 4484 2676
rect 4516 2644 4644 2676
rect 4676 2644 4680 2676
rect 4480 2640 4680 2644
rect 4720 2676 5080 2680
rect 4720 2644 4724 2676
rect 4756 2644 4884 2676
rect 4916 2644 5044 2676
rect 5076 2644 5080 2676
rect 4720 2640 5080 2644
rect 5120 2676 5480 2680
rect 5120 2644 5124 2676
rect 5156 2644 5284 2676
rect 5316 2644 5444 2676
rect 5476 2644 5480 2676
rect 5120 2640 5480 2644
rect 5520 2676 5880 2680
rect 5520 2644 5524 2676
rect 5556 2644 5684 2676
rect 5716 2644 5844 2676
rect 5876 2644 5880 2676
rect 5520 2640 5880 2644
rect 5920 2676 6120 2680
rect 5920 2644 5924 2676
rect 5956 2644 6084 2676
rect 6116 2644 6120 2676
rect 5920 2640 6120 2644
rect 6160 2676 6360 2680
rect 6160 2644 6164 2676
rect 6196 2644 6324 2676
rect 6356 2644 6360 2676
rect 6160 2640 6360 2644
rect 4240 2596 4440 2600
rect 4240 2564 4244 2596
rect 4276 2564 4404 2596
rect 4436 2564 4440 2596
rect 4240 2560 4440 2564
rect 4480 2596 4680 2600
rect 4480 2564 4484 2596
rect 4516 2564 4644 2596
rect 4676 2564 4680 2596
rect 4480 2560 4680 2564
rect 4720 2596 5080 2600
rect 4720 2564 4724 2596
rect 4756 2564 4884 2596
rect 4916 2564 5044 2596
rect 5076 2564 5080 2596
rect 4720 2560 5080 2564
rect 5120 2596 5480 2600
rect 5120 2564 5124 2596
rect 5156 2564 5284 2596
rect 5316 2564 5444 2596
rect 5476 2564 5480 2596
rect 5120 2560 5480 2564
rect 5520 2596 5880 2600
rect 5520 2564 5524 2596
rect 5556 2564 5684 2596
rect 5716 2564 5844 2596
rect 5876 2564 5880 2596
rect 5520 2560 5880 2564
rect 5920 2596 6120 2600
rect 5920 2564 5924 2596
rect 5956 2564 6084 2596
rect 6116 2564 6120 2596
rect 5920 2560 6120 2564
rect 6160 2596 6360 2600
rect 6160 2564 6164 2596
rect 6196 2564 6324 2596
rect 6356 2564 6360 2596
rect 6160 2560 6360 2564
rect 4240 2516 4440 2520
rect 4240 2484 4244 2516
rect 4276 2484 4404 2516
rect 4436 2484 4440 2516
rect 4240 2480 4440 2484
rect 4480 2516 4680 2520
rect 4480 2484 4484 2516
rect 4516 2484 4644 2516
rect 4676 2484 4680 2516
rect 4480 2480 4680 2484
rect 4720 2516 5080 2520
rect 4720 2484 4724 2516
rect 4756 2484 4884 2516
rect 4916 2484 5044 2516
rect 5076 2484 5080 2516
rect 4720 2480 5080 2484
rect 5120 2516 5480 2520
rect 5120 2484 5124 2516
rect 5156 2484 5284 2516
rect 5316 2484 5444 2516
rect 5476 2484 5480 2516
rect 5120 2480 5480 2484
rect 5520 2516 5880 2520
rect 5520 2484 5524 2516
rect 5556 2484 5684 2516
rect 5716 2484 5844 2516
rect 5876 2484 5880 2516
rect 5520 2480 5880 2484
rect 5920 2516 6120 2520
rect 5920 2484 5924 2516
rect 5956 2484 6084 2516
rect 6116 2484 6120 2516
rect 5920 2480 6120 2484
rect 6160 2516 6360 2520
rect 6160 2484 6164 2516
rect 6196 2484 6324 2516
rect 6356 2484 6360 2516
rect 6160 2480 6360 2484
rect 4240 2436 4440 2440
rect 4240 2404 4244 2436
rect 4276 2404 4404 2436
rect 4436 2404 4440 2436
rect 4240 2400 4440 2404
rect 4480 2436 4680 2440
rect 4480 2404 4484 2436
rect 4516 2404 4644 2436
rect 4676 2404 4680 2436
rect 4480 2400 4680 2404
rect 4720 2436 5080 2440
rect 4720 2404 4724 2436
rect 4756 2404 4884 2436
rect 4916 2404 5044 2436
rect 5076 2404 5080 2436
rect 4720 2400 5080 2404
rect 5120 2436 5480 2440
rect 5120 2404 5124 2436
rect 5156 2404 5284 2436
rect 5316 2404 5444 2436
rect 5476 2404 5480 2436
rect 5120 2400 5480 2404
rect 5520 2436 5880 2440
rect 5520 2404 5524 2436
rect 5556 2404 5684 2436
rect 5716 2404 5844 2436
rect 5876 2404 5880 2436
rect 5520 2400 5880 2404
rect 5920 2436 6120 2440
rect 5920 2404 5924 2436
rect 5956 2404 6084 2436
rect 6116 2404 6120 2436
rect 5920 2400 6120 2404
rect 6160 2436 6360 2440
rect 6160 2404 6164 2436
rect 6196 2404 6324 2436
rect 6356 2404 6360 2436
rect 6160 2400 6360 2404
rect 4240 2356 4440 2360
rect 4240 2324 4244 2356
rect 4276 2324 4404 2356
rect 4436 2324 4440 2356
rect 4240 2320 4440 2324
rect 4480 2356 4680 2360
rect 4480 2324 4484 2356
rect 4516 2324 4644 2356
rect 4676 2324 4680 2356
rect 4480 2320 4680 2324
rect 4720 2356 5080 2360
rect 4720 2324 4724 2356
rect 4756 2324 4884 2356
rect 4916 2324 5044 2356
rect 5076 2324 5080 2356
rect 4720 2320 5080 2324
rect 5120 2356 5480 2360
rect 5120 2324 5124 2356
rect 5156 2324 5284 2356
rect 5316 2324 5444 2356
rect 5476 2324 5480 2356
rect 5120 2320 5480 2324
rect 5520 2356 5880 2360
rect 5520 2324 5524 2356
rect 5556 2324 5684 2356
rect 5716 2324 5844 2356
rect 5876 2324 5880 2356
rect 5520 2320 5880 2324
rect 5920 2356 6120 2360
rect 5920 2324 5924 2356
rect 5956 2324 6084 2356
rect 6116 2324 6120 2356
rect 5920 2320 6120 2324
rect 6160 2356 6360 2360
rect 6160 2324 6164 2356
rect 6196 2324 6324 2356
rect 6356 2324 6360 2356
rect 6160 2320 6360 2324
rect 4240 2276 4440 2280
rect 4240 2244 4244 2276
rect 4276 2244 4404 2276
rect 4436 2244 4440 2276
rect 4240 2240 4440 2244
rect 4480 2276 4680 2280
rect 4480 2244 4484 2276
rect 4516 2244 4644 2276
rect 4676 2244 4680 2276
rect 4480 2240 4680 2244
rect 4720 2276 5080 2280
rect 4720 2244 4724 2276
rect 4756 2244 4884 2276
rect 4916 2244 5044 2276
rect 5076 2244 5080 2276
rect 4720 2240 5080 2244
rect 5120 2276 5480 2280
rect 5120 2244 5124 2276
rect 5156 2244 5284 2276
rect 5316 2244 5444 2276
rect 5476 2244 5480 2276
rect 5120 2240 5480 2244
rect 5520 2276 5880 2280
rect 5520 2244 5524 2276
rect 5556 2244 5684 2276
rect 5716 2244 5844 2276
rect 5876 2244 5880 2276
rect 5520 2240 5880 2244
rect 5920 2276 6120 2280
rect 5920 2244 5924 2276
rect 5956 2244 6084 2276
rect 6116 2244 6120 2276
rect 5920 2240 6120 2244
rect 6160 2276 6360 2280
rect 6160 2244 6164 2276
rect 6196 2244 6324 2276
rect 6356 2244 6360 2276
rect 6160 2240 6360 2244
rect 4240 2196 4440 2200
rect 4240 2164 4244 2196
rect 4276 2164 4404 2196
rect 4436 2164 4440 2196
rect 4240 2160 4440 2164
rect 4480 2196 4680 2200
rect 4480 2164 4484 2196
rect 4516 2164 4644 2196
rect 4676 2164 4680 2196
rect 4480 2160 4680 2164
rect 4720 2196 5080 2200
rect 4720 2164 4724 2196
rect 4756 2164 4884 2196
rect 4916 2164 5044 2196
rect 5076 2164 5080 2196
rect 4720 2160 5080 2164
rect 5120 2196 5480 2200
rect 5120 2164 5124 2196
rect 5156 2164 5284 2196
rect 5316 2164 5444 2196
rect 5476 2164 5480 2196
rect 5120 2160 5480 2164
rect 5520 2196 5880 2200
rect 5520 2164 5524 2196
rect 5556 2164 5684 2196
rect 5716 2164 5844 2196
rect 5876 2164 5880 2196
rect 5520 2160 5880 2164
rect 5920 2196 6120 2200
rect 5920 2164 5924 2196
rect 5956 2164 6084 2196
rect 6116 2164 6120 2196
rect 5920 2160 6120 2164
rect 6160 2196 6360 2200
rect 6160 2164 6164 2196
rect 6196 2164 6324 2196
rect 6356 2164 6360 2196
rect 6160 2160 6360 2164
rect 4240 2116 4440 2120
rect 4240 2084 4244 2116
rect 4276 2084 4404 2116
rect 4436 2084 4440 2116
rect 4240 2080 4440 2084
rect 4480 2116 4680 2120
rect 4480 2084 4484 2116
rect 4516 2084 4644 2116
rect 4676 2084 4680 2116
rect 4480 2080 4680 2084
rect 4720 2116 5080 2120
rect 4720 2084 4724 2116
rect 4756 2084 4884 2116
rect 4916 2084 5044 2116
rect 5076 2084 5080 2116
rect 4720 2080 5080 2084
rect 5120 2116 5480 2120
rect 5120 2084 5124 2116
rect 5156 2084 5284 2116
rect 5316 2084 5444 2116
rect 5476 2084 5480 2116
rect 5120 2080 5480 2084
rect 5520 2116 5880 2120
rect 5520 2084 5524 2116
rect 5556 2084 5684 2116
rect 5716 2084 5844 2116
rect 5876 2084 5880 2116
rect 5520 2080 5880 2084
rect 5920 2116 6120 2120
rect 5920 2084 5924 2116
rect 5956 2084 6084 2116
rect 6116 2084 6120 2116
rect 5920 2080 6120 2084
rect 6160 2116 6360 2120
rect 6160 2084 6164 2116
rect 6196 2084 6324 2116
rect 6356 2084 6360 2116
rect 6160 2080 6360 2084
rect 4240 2036 4440 2040
rect 4240 2004 4244 2036
rect 4276 2004 4404 2036
rect 4436 2004 4440 2036
rect 4240 2000 4440 2004
rect 4480 2036 4680 2040
rect 4480 2004 4484 2036
rect 4516 2004 4644 2036
rect 4676 2004 4680 2036
rect 4480 2000 4680 2004
rect 4720 2036 5080 2040
rect 4720 2004 4724 2036
rect 4756 2004 4884 2036
rect 4916 2004 5044 2036
rect 5076 2004 5080 2036
rect 4720 2000 5080 2004
rect 5120 2036 5480 2040
rect 5120 2004 5124 2036
rect 5156 2004 5284 2036
rect 5316 2004 5444 2036
rect 5476 2004 5480 2036
rect 5120 2000 5480 2004
rect 5520 2036 5880 2040
rect 5520 2004 5524 2036
rect 5556 2004 5684 2036
rect 5716 2004 5844 2036
rect 5876 2004 5880 2036
rect 5520 2000 5880 2004
rect 5920 2036 6120 2040
rect 5920 2004 5924 2036
rect 5956 2004 6084 2036
rect 6116 2004 6120 2036
rect 5920 2000 6120 2004
rect 6160 2036 6360 2040
rect 6160 2004 6164 2036
rect 6196 2004 6324 2036
rect 6356 2004 6360 2036
rect 6160 2000 6360 2004
rect 4240 1636 4440 1640
rect 4240 1604 4244 1636
rect 4276 1604 4404 1636
rect 4436 1604 4440 1636
rect 4240 1600 4440 1604
rect 4480 1636 4680 1640
rect 4480 1604 4484 1636
rect 4516 1604 4644 1636
rect 4676 1604 4680 1636
rect 4480 1600 4680 1604
rect 4720 1636 5080 1640
rect 4720 1604 4724 1636
rect 4756 1604 4884 1636
rect 4916 1604 5044 1636
rect 5076 1604 5080 1636
rect 4720 1600 5080 1604
rect 5120 1636 5480 1640
rect 5120 1604 5124 1636
rect 5156 1604 5284 1636
rect 5316 1604 5444 1636
rect 5476 1604 5480 1636
rect 5120 1600 5480 1604
rect 5520 1636 5880 1640
rect 5520 1604 5524 1636
rect 5556 1604 5684 1636
rect 5716 1604 5844 1636
rect 5876 1604 5880 1636
rect 5520 1600 5880 1604
rect 5920 1636 6120 1640
rect 5920 1604 5924 1636
rect 5956 1604 6084 1636
rect 6116 1604 6120 1636
rect 5920 1600 6120 1604
rect 6160 1636 6360 1640
rect 6160 1604 6164 1636
rect 6196 1604 6324 1636
rect 6356 1604 6360 1636
rect 6160 1600 6360 1604
rect 4240 1556 4440 1560
rect 4240 1524 4244 1556
rect 4276 1524 4404 1556
rect 4436 1524 4440 1556
rect 4240 1520 4440 1524
rect 4480 1556 4680 1560
rect 4480 1524 4484 1556
rect 4516 1524 4644 1556
rect 4676 1524 4680 1556
rect 4480 1520 4680 1524
rect 4720 1556 5080 1560
rect 4720 1524 4724 1556
rect 4756 1524 4884 1556
rect 4916 1524 5044 1556
rect 5076 1524 5080 1556
rect 4720 1520 5080 1524
rect 5120 1556 5480 1560
rect 5120 1524 5124 1556
rect 5156 1524 5284 1556
rect 5316 1524 5444 1556
rect 5476 1524 5480 1556
rect 5120 1520 5480 1524
rect 5520 1556 5880 1560
rect 5520 1524 5524 1556
rect 5556 1524 5684 1556
rect 5716 1524 5844 1556
rect 5876 1524 5880 1556
rect 5520 1520 5880 1524
rect 5920 1556 6120 1560
rect 5920 1524 5924 1556
rect 5956 1524 6084 1556
rect 6116 1524 6120 1556
rect 5920 1520 6120 1524
rect 6160 1556 6360 1560
rect 6160 1524 6164 1556
rect 6196 1524 6324 1556
rect 6356 1524 6360 1556
rect 6160 1520 6360 1524
rect 4240 1476 4440 1480
rect 4240 1444 4244 1476
rect 4276 1444 4404 1476
rect 4436 1444 4440 1476
rect 4240 1440 4440 1444
rect 4480 1476 4680 1480
rect 4480 1444 4484 1476
rect 4516 1444 4644 1476
rect 4676 1444 4680 1476
rect 4480 1440 4680 1444
rect 4720 1476 5080 1480
rect 4720 1444 4724 1476
rect 4756 1444 4884 1476
rect 4916 1444 5044 1476
rect 5076 1444 5080 1476
rect 4720 1440 5080 1444
rect 5120 1476 5480 1480
rect 5120 1444 5124 1476
rect 5156 1444 5284 1476
rect 5316 1444 5444 1476
rect 5476 1444 5480 1476
rect 5120 1440 5480 1444
rect 5520 1476 5880 1480
rect 5520 1444 5524 1476
rect 5556 1444 5684 1476
rect 5716 1444 5844 1476
rect 5876 1444 5880 1476
rect 5520 1440 5880 1444
rect 5920 1476 6120 1480
rect 5920 1444 5924 1476
rect 5956 1444 6084 1476
rect 6116 1444 6120 1476
rect 5920 1440 6120 1444
rect 6160 1476 6360 1480
rect 6160 1444 6164 1476
rect 6196 1444 6324 1476
rect 6356 1444 6360 1476
rect 6160 1440 6360 1444
rect 4240 1396 4440 1400
rect 4240 1364 4244 1396
rect 4276 1364 4404 1396
rect 4436 1364 4440 1396
rect 4240 1360 4440 1364
rect 4480 1396 4680 1400
rect 4480 1364 4484 1396
rect 4516 1364 4644 1396
rect 4676 1364 4680 1396
rect 4480 1360 4680 1364
rect 4720 1396 5080 1400
rect 4720 1364 4724 1396
rect 4756 1364 4884 1396
rect 4916 1364 5044 1396
rect 5076 1364 5080 1396
rect 4720 1360 5080 1364
rect 5120 1396 5480 1400
rect 5120 1364 5124 1396
rect 5156 1364 5284 1396
rect 5316 1364 5444 1396
rect 5476 1364 5480 1396
rect 5120 1360 5480 1364
rect 5520 1396 5880 1400
rect 5520 1364 5524 1396
rect 5556 1364 5684 1396
rect 5716 1364 5844 1396
rect 5876 1364 5880 1396
rect 5520 1360 5880 1364
rect 5920 1396 6120 1400
rect 5920 1364 5924 1396
rect 5956 1364 6084 1396
rect 6116 1364 6120 1396
rect 5920 1360 6120 1364
rect 6160 1396 6360 1400
rect 6160 1364 6164 1396
rect 6196 1364 6324 1396
rect 6356 1364 6360 1396
rect 6160 1360 6360 1364
rect 4240 1316 4440 1320
rect 4240 1284 4244 1316
rect 4276 1284 4404 1316
rect 4436 1284 4440 1316
rect 4240 1280 4440 1284
rect 4480 1316 4680 1320
rect 4480 1284 4484 1316
rect 4516 1284 4644 1316
rect 4676 1284 4680 1316
rect 4480 1280 4680 1284
rect 4720 1316 5080 1320
rect 4720 1284 4724 1316
rect 4756 1284 4884 1316
rect 4916 1284 5044 1316
rect 5076 1284 5080 1316
rect 4720 1280 5080 1284
rect 5120 1316 5480 1320
rect 5120 1284 5124 1316
rect 5156 1284 5284 1316
rect 5316 1284 5444 1316
rect 5476 1284 5480 1316
rect 5120 1280 5480 1284
rect 5520 1316 5880 1320
rect 5520 1284 5524 1316
rect 5556 1284 5684 1316
rect 5716 1284 5844 1316
rect 5876 1284 5880 1316
rect 5520 1280 5880 1284
rect 5920 1316 6120 1320
rect 5920 1284 5924 1316
rect 5956 1284 6084 1316
rect 6116 1284 6120 1316
rect 5920 1280 6120 1284
rect 6160 1316 6360 1320
rect 6160 1284 6164 1316
rect 6196 1284 6324 1316
rect 6356 1284 6360 1316
rect 6160 1280 6360 1284
rect 4240 1236 4440 1240
rect 4240 1204 4244 1236
rect 4276 1204 4404 1236
rect 4436 1204 4440 1236
rect 4240 1200 4440 1204
rect 4480 1236 4680 1240
rect 4480 1204 4484 1236
rect 4516 1204 4644 1236
rect 4676 1204 4680 1236
rect 4480 1200 4680 1204
rect 4720 1236 5080 1240
rect 4720 1204 4724 1236
rect 4756 1204 4884 1236
rect 4916 1204 5044 1236
rect 5076 1204 5080 1236
rect 4720 1200 5080 1204
rect 5120 1236 5480 1240
rect 5120 1204 5124 1236
rect 5156 1204 5284 1236
rect 5316 1204 5444 1236
rect 5476 1204 5480 1236
rect 5120 1200 5480 1204
rect 5520 1236 5880 1240
rect 5520 1204 5524 1236
rect 5556 1204 5684 1236
rect 5716 1204 5844 1236
rect 5876 1204 5880 1236
rect 5520 1200 5880 1204
rect 5920 1236 6120 1240
rect 5920 1204 5924 1236
rect 5956 1204 6084 1236
rect 6116 1204 6120 1236
rect 5920 1200 6120 1204
rect 6160 1236 6360 1240
rect 6160 1204 6164 1236
rect 6196 1204 6324 1236
rect 6356 1204 6360 1236
rect 6160 1200 6360 1204
rect 4240 1156 4440 1160
rect 4240 1124 4244 1156
rect 4276 1124 4404 1156
rect 4436 1124 4440 1156
rect 4240 1120 4440 1124
rect 4480 1156 4680 1160
rect 4480 1124 4484 1156
rect 4516 1124 4644 1156
rect 4676 1124 4680 1156
rect 4480 1120 4680 1124
rect 4720 1156 5080 1160
rect 4720 1124 4724 1156
rect 4756 1124 4884 1156
rect 4916 1124 5044 1156
rect 5076 1124 5080 1156
rect 4720 1120 5080 1124
rect 5120 1156 5480 1160
rect 5120 1124 5124 1156
rect 5156 1124 5284 1156
rect 5316 1124 5444 1156
rect 5476 1124 5480 1156
rect 5120 1120 5480 1124
rect 5520 1156 5880 1160
rect 5520 1124 5524 1156
rect 5556 1124 5684 1156
rect 5716 1124 5844 1156
rect 5876 1124 5880 1156
rect 5520 1120 5880 1124
rect 5920 1156 6120 1160
rect 5920 1124 5924 1156
rect 5956 1124 6084 1156
rect 6116 1124 6120 1156
rect 5920 1120 6120 1124
rect 6160 1156 6360 1160
rect 6160 1124 6164 1156
rect 6196 1124 6324 1156
rect 6356 1124 6360 1156
rect 6160 1120 6360 1124
rect 4240 1076 4440 1080
rect 4240 1044 4244 1076
rect 4276 1044 4404 1076
rect 4436 1044 4440 1076
rect 4240 1040 4440 1044
rect 4480 1076 4680 1080
rect 4480 1044 4484 1076
rect 4516 1044 4644 1076
rect 4676 1044 4680 1076
rect 4480 1040 4680 1044
rect 4720 1076 5080 1080
rect 4720 1044 4724 1076
rect 4756 1044 4884 1076
rect 4916 1044 5044 1076
rect 5076 1044 5080 1076
rect 4720 1040 5080 1044
rect 5120 1076 5480 1080
rect 5120 1044 5124 1076
rect 5156 1044 5284 1076
rect 5316 1044 5444 1076
rect 5476 1044 5480 1076
rect 5120 1040 5480 1044
rect 5520 1076 5880 1080
rect 5520 1044 5524 1076
rect 5556 1044 5684 1076
rect 5716 1044 5844 1076
rect 5876 1044 5880 1076
rect 5520 1040 5880 1044
rect 5920 1076 6120 1080
rect 5920 1044 5924 1076
rect 5956 1044 6084 1076
rect 6116 1044 6120 1076
rect 5920 1040 6120 1044
rect 6160 1076 6360 1080
rect 6160 1044 6164 1076
rect 6196 1044 6324 1076
rect 6356 1044 6360 1076
rect 6160 1040 6360 1044
rect 4240 756 4440 760
rect 4240 724 4244 756
rect 4276 724 4404 756
rect 4436 724 4440 756
rect 4240 720 4440 724
rect 4480 756 4680 760
rect 4480 724 4484 756
rect 4516 724 4644 756
rect 4676 724 4680 756
rect 4480 720 4680 724
rect 4720 756 5080 760
rect 4720 724 4724 756
rect 4756 724 4884 756
rect 4916 724 5044 756
rect 5076 724 5080 756
rect 4720 720 5080 724
rect 5120 756 5480 760
rect 5120 724 5124 756
rect 5156 724 5284 756
rect 5316 724 5444 756
rect 5476 724 5480 756
rect 5120 720 5480 724
rect 5520 756 5880 760
rect 5520 724 5524 756
rect 5556 724 5684 756
rect 5716 724 5844 756
rect 5876 724 5880 756
rect 5520 720 5880 724
rect 5920 756 6120 760
rect 5920 724 5924 756
rect 5956 724 6084 756
rect 6116 724 6120 756
rect 5920 720 6120 724
rect 6160 756 6360 760
rect 6160 724 6164 756
rect 6196 724 6324 756
rect 6356 724 6360 756
rect 6160 720 6360 724
rect 4240 676 4440 680
rect 4240 644 4244 676
rect 4276 644 4404 676
rect 4436 644 4440 676
rect 4240 640 4440 644
rect 4480 676 4680 680
rect 4480 644 4484 676
rect 4516 644 4644 676
rect 4676 644 4680 676
rect 4480 640 4680 644
rect 4720 676 5080 680
rect 4720 644 4724 676
rect 4756 644 4884 676
rect 4916 644 5044 676
rect 5076 644 5080 676
rect 4720 640 5080 644
rect 5120 676 5480 680
rect 5120 644 5124 676
rect 5156 644 5284 676
rect 5316 644 5444 676
rect 5476 644 5480 676
rect 5120 640 5480 644
rect 5520 676 5880 680
rect 5520 644 5524 676
rect 5556 644 5684 676
rect 5716 644 5844 676
rect 5876 644 5880 676
rect 5520 640 5880 644
rect 5920 676 6120 680
rect 5920 644 5924 676
rect 5956 644 6084 676
rect 6116 644 6120 676
rect 5920 640 6120 644
rect 6160 676 6360 680
rect 6160 644 6164 676
rect 6196 644 6324 676
rect 6356 644 6360 676
rect 6160 640 6360 644
rect 4240 596 4440 600
rect 4240 564 4244 596
rect 4276 564 4404 596
rect 4436 564 4440 596
rect 4240 560 4440 564
rect 4480 596 4680 600
rect 4480 564 4484 596
rect 4516 564 4644 596
rect 4676 564 4680 596
rect 4480 560 4680 564
rect 4720 596 5080 600
rect 4720 564 4724 596
rect 4756 564 4884 596
rect 4916 564 5044 596
rect 5076 564 5080 596
rect 4720 560 5080 564
rect 5120 596 5480 600
rect 5120 564 5124 596
rect 5156 564 5284 596
rect 5316 564 5444 596
rect 5476 564 5480 596
rect 5120 560 5480 564
rect 5520 596 5880 600
rect 5520 564 5524 596
rect 5556 564 5684 596
rect 5716 564 5844 596
rect 5876 564 5880 596
rect 5520 560 5880 564
rect 5920 596 6120 600
rect 5920 564 5924 596
rect 5956 564 6084 596
rect 6116 564 6120 596
rect 5920 560 6120 564
rect 6160 596 6360 600
rect 6160 564 6164 596
rect 6196 564 6324 596
rect 6356 564 6360 596
rect 6160 560 6360 564
rect 4240 196 4440 200
rect 4240 164 4244 196
rect 4276 164 4404 196
rect 4436 164 4440 196
rect 4240 160 4440 164
rect 4480 196 4680 200
rect 4480 164 4484 196
rect 4516 164 4644 196
rect 4676 164 4680 196
rect 4480 160 4680 164
rect 4720 196 5080 200
rect 4720 164 4724 196
rect 4756 164 4884 196
rect 4916 164 5044 196
rect 5076 164 5080 196
rect 4720 160 5080 164
rect 5120 196 5480 200
rect 5120 164 5124 196
rect 5156 164 5284 196
rect 5316 164 5444 196
rect 5476 164 5480 196
rect 5120 160 5480 164
rect 5520 196 5880 200
rect 5520 164 5524 196
rect 5556 164 5684 196
rect 5716 164 5844 196
rect 5876 164 5880 196
rect 5520 160 5880 164
rect 5920 196 6120 200
rect 5920 164 5924 196
rect 5956 164 6084 196
rect 6116 164 6120 196
rect 5920 160 6120 164
rect 6160 196 6360 200
rect 6160 164 6164 196
rect 6196 164 6324 196
rect 6356 164 6360 196
rect 6160 160 6360 164
rect 4240 116 4440 120
rect 4240 84 4244 116
rect 4276 84 4404 116
rect 4436 84 4440 116
rect 4240 80 4440 84
rect 4480 116 4680 120
rect 4480 84 4484 116
rect 4516 84 4644 116
rect 4676 84 4680 116
rect 4480 80 4680 84
rect 4720 116 5080 120
rect 4720 84 4724 116
rect 4756 84 4884 116
rect 4916 84 5044 116
rect 5076 84 5080 116
rect 4720 80 5080 84
rect 5120 116 5480 120
rect 5120 84 5124 116
rect 5156 84 5284 116
rect 5316 84 5444 116
rect 5476 84 5480 116
rect 5120 80 5480 84
rect 5520 116 5880 120
rect 5520 84 5524 116
rect 5556 84 5684 116
rect 5716 84 5844 116
rect 5876 84 5880 116
rect 5520 80 5880 84
rect 5920 116 6120 120
rect 5920 84 5924 116
rect 5956 84 6084 116
rect 6116 84 6120 116
rect 5920 80 6120 84
rect 6160 116 6360 120
rect 6160 84 6164 116
rect 6196 84 6324 116
rect 6356 84 6360 116
rect 6160 80 6360 84
rect 4240 36 4440 40
rect 4240 4 4244 36
rect 4276 4 4404 36
rect 4436 4 4440 36
rect 4240 0 4440 4
rect 4480 36 4680 40
rect 4480 4 4484 36
rect 4516 4 4644 36
rect 4676 4 4680 36
rect 4480 0 4680 4
rect 4720 36 5080 40
rect 4720 4 4724 36
rect 4756 4 4884 36
rect 4916 4 5044 36
rect 5076 4 5080 36
rect 4720 0 5080 4
rect 5120 36 5480 40
rect 5120 4 5124 36
rect 5156 4 5284 36
rect 5316 4 5444 36
rect 5476 4 5480 36
rect 5120 0 5480 4
rect 5520 36 5880 40
rect 5520 4 5524 36
rect 5556 4 5684 36
rect 5716 4 5844 36
rect 5876 4 5880 36
rect 5520 0 5880 4
rect 5920 36 6120 40
rect 5920 4 5924 36
rect 5956 4 6084 36
rect 6116 4 6120 36
rect 5920 0 6120 4
rect 6160 36 6360 40
rect 6160 4 6164 36
rect 6196 4 6324 36
rect 6356 4 6360 36
rect 6160 0 6360 4
<< via4 >>
rect 1560 13480 1680 13600
rect 2520 13480 2640 13600
rect 7960 13480 8080 13600
rect 8920 13480 9040 13600
rect 1080 13240 1200 13360
rect 2040 13240 2160 13360
rect 3000 13240 3120 13360
rect 7480 13240 7600 13360
rect 8440 13240 8560 13360
rect 9400 13240 9520 13360
rect 600 13000 720 13120
rect 3480 13000 3600 13120
rect 7000 13000 7120 13120
rect 9880 13000 10000 13120
rect 120 12760 240 12880
rect 3960 12760 4080 12880
rect 6520 12760 6640 12880
rect 10360 12760 10480 12880
<< metal5 >>
rect 80 12880 280 13640
rect 80 12760 120 12880
rect 240 12760 280 12880
rect 80 12680 280 12760
rect 560 13120 760 13640
rect 560 13000 600 13120
rect 720 13000 760 13120
rect 560 12680 760 13000
rect 1040 13360 1240 13640
rect 1040 13240 1080 13360
rect 1200 13240 1240 13360
rect 1040 12680 1240 13240
rect 1520 13600 1720 13640
rect 1520 13480 1560 13600
rect 1680 13480 1720 13600
rect 1520 12680 1720 13480
rect 2000 13360 2200 13640
rect 2000 13240 2040 13360
rect 2160 13240 2200 13360
rect 2000 12680 2200 13240
rect 2480 13600 2680 13640
rect 2480 13480 2520 13600
rect 2640 13480 2680 13600
rect 2480 12680 2680 13480
rect 2960 13360 3160 13640
rect 2960 13240 3000 13360
rect 3120 13240 3160 13360
rect 2960 12680 3160 13240
rect 3440 13120 3640 13640
rect 3440 13000 3480 13120
rect 3600 13000 3640 13120
rect 3440 12680 3640 13000
rect 3920 12880 4120 13640
rect 3920 12760 3960 12880
rect 4080 12760 4120 12880
rect 3920 12680 4120 12760
rect 6480 12880 6680 13640
rect 6480 12760 6520 12880
rect 6640 12760 6680 12880
rect 6480 12680 6680 12760
rect 6960 13120 7160 13640
rect 6960 13000 7000 13120
rect 7120 13000 7160 13120
rect 6960 12680 7160 13000
rect 7440 13360 7640 13640
rect 7440 13240 7480 13360
rect 7600 13240 7640 13360
rect 7440 12680 7640 13240
rect 7920 13600 8120 13640
rect 7920 13480 7960 13600
rect 8080 13480 8120 13600
rect 7920 12680 8120 13480
rect 8400 13360 8600 13640
rect 8400 13240 8440 13360
rect 8560 13240 8600 13360
rect 8400 12680 8600 13240
rect 8880 13600 9080 13640
rect 8880 13480 8920 13600
rect 9040 13480 9080 13600
rect 8880 12680 9080 13480
rect 9360 13360 9560 13640
rect 9360 13240 9400 13360
rect 9520 13240 9560 13360
rect 9360 12680 9560 13240
rect 9840 13120 10040 13640
rect 9840 13000 9880 13120
rect 10000 13000 10040 13120
rect 9840 12680 10040 13000
rect 10320 12880 10520 13640
rect 10320 12760 10360 12880
rect 10480 12760 10520 12880
rect 10320 12680 10520 12760
rect 80 10640 280 10680
rect 560 10640 760 10680
rect 1040 10640 1240 10680
rect 1520 10640 1720 10680
rect 2000 10640 2200 10680
rect 2480 10640 2680 10680
rect 2960 10640 3160 10680
rect 3440 10640 3640 10680
rect 3920 10640 4120 10680
rect 6480 10640 6680 10680
rect 6960 10640 7160 10680
rect 7440 10640 7640 10680
rect 7920 10640 8120 10680
rect 8400 10640 8600 10680
rect 8880 10640 9080 10680
rect 9360 10640 9560 10680
rect 9840 10640 10040 10680
rect 10320 10640 10520 10680
rect 80 7600 280 7640
rect 560 7600 760 7640
rect 1040 7600 1240 7640
rect 1520 7600 1720 7640
rect 2000 7600 2200 7640
rect 2480 7600 2680 7640
rect 2960 7600 3160 7640
rect 3440 7600 3640 7640
rect 3920 7600 4120 7640
rect 6480 7600 6680 7640
rect 6960 7600 7160 7640
rect 7440 7600 7640 7640
rect 7920 7600 8120 7640
rect 8400 7600 8600 7640
rect 8880 7600 9080 7640
rect 9360 7600 9560 7640
rect 9840 7600 10040 7640
rect 10320 7600 10520 7640
rect 80 5560 280 5600
rect 560 5560 760 5600
rect 1040 5560 1240 5600
rect 1520 5560 1720 5600
rect 2000 5560 2200 5600
rect 2480 5560 2680 5600
rect 2960 5560 3160 5600
rect 3440 5560 3640 5600
rect 3920 5560 4120 5600
rect 6480 5560 6680 5600
rect 6960 5560 7160 5600
rect 7440 5560 7640 5600
rect 7920 5560 8120 5600
rect 8400 5560 8600 5600
rect 8880 5560 9080 5600
rect 9360 5560 9560 5600
rect 9840 5560 10040 5600
rect 10320 5560 10520 5600
rect 80 -40 280 0
rect 560 -40 760 0
rect 1040 -40 1240 0
rect 1520 -40 1720 0
rect 2000 -40 2200 0
rect 2480 -40 2680 0
rect 2960 -40 3160 0
rect 3440 -40 3640 0
rect 3920 -40 4120 0
use invt  br ../../inv/mag
timestamp 1637985169
transform -1 0 10600 0 1 7640
box 0 0 4200 3000
use invt  bl
timestamp 1637985169
transform 1 0 0 0 1 7640
box 0 0 4200 3000
use inv_2_2  ar ../../inv/mag
timestamp 1637985251
transform -1 0 10600 0 1 5600
box 0 0 4200 2000
use inv_2_2  cr
timestamp 1637985251
transform -1 0 10600 0 1 10680
box 0 0 4200 2000
use inv_2_2  cl
timestamp 1637985251
transform 1 0 0 0 1 10680
box 0 0 4200 2000
use inv_2_2  al
timestamp 1637985251
transform 1 0 0 0 1 5600
box 0 0 4200 2000
use inv_bias  biasr ../../inv/mag
timestamp 1637985316
transform -1 0 10600 0 1 520
box 0 -520 4200 5040
use inv_bias  biasl
timestamp 1637985316
transform 1 0 0 0 1 520
box 0 -520 4200 5040
<< labels >>
rlabel metal3 4800 -40 4840 0 0 im
port 0 nsew
rlabel metal3 5760 -40 5800 0 0 ip
port 1 nsew
rlabel metal3 5120 -40 5160 0 0 out
port 2 nsew
rlabel metal3 4320 -40 4360 0 0 ib
port 3 nsew
rlabel metal3 6240 -40 6280 0 0 q
port 4 nsew
rlabel metal5 80 -40 280 0 0 vdda
port 5 nsew
rlabel metal3 4560 -40 4600 0 0 bp
port 6 nsew
rlabel metal5 560 -40 760 0 0 vddx
port 7 nsew
rlabel metal5 1040 -40 1240 0 0 gnda
port 8 nsew
rlabel metal5 1520 -40 1720 0 0 vssa
port 9 nsew
rlabel metal3 5200 -40 5240 0 0 xn
port 10 nsew
rlabel metal3 5360 -40 5400 0 0 xp
port 11 nsew
rlabel metal3 4960 -40 5000 0 0 x
port 12 nsew
rlabel metal3 5600 -40 5640 0 0 y
port 13 nsew
rlabel metal3 6000 -40 6040 0 0 z
port 14 nsew
<< end >>
